module top (\dcnt_reg[0]/P0001 , \dcnt_reg[1]/P0001 , \dcnt_reg[2]/P0001 , \dcnt_reg[3]/P0001 , \key[0]_pad , \key[100]_pad , \key[101]_pad , \key[102]_pad , \key[103]_pad , \key[104]_pad , \key[105]_pad , \key[106]_pad , \key[107]_pad , \key[108]_pad , \key[109]_pad , \key[10]_pad , \key[110]_pad , \key[111]_pad , \key[112]_pad , \key[113]_pad , \key[114]_pad , \key[115]_pad , \key[116]_pad , \key[117]_pad , \key[118]_pad , \key[119]_pad , \key[11]_pad , \key[120]_pad , \key[121]_pad , \key[122]_pad , \key[123]_pad , \key[124]_pad , \key[125]_pad , \key[126]_pad , \key[127]_pad , \key[12]_pad , \key[13]_pad , \key[14]_pad , \key[15]_pad , \key[16]_pad , \key[17]_pad , \key[18]_pad , \key[19]_pad , \key[1]_pad , \key[20]_pad , \key[21]_pad , \key[22]_pad , \key[23]_pad , \key[24]_pad , \key[25]_pad , \key[26]_pad , \key[27]_pad , \key[28]_pad , \key[29]_pad , \key[2]_pad , \key[30]_pad , \key[31]_pad , \key[32]_pad , \key[33]_pad , \key[34]_pad , \key[35]_pad , \key[36]_pad , \key[37]_pad , \key[38]_pad , \key[39]_pad , \key[3]_pad , \key[40]_pad , \key[41]_pad , \key[42]_pad , \key[43]_pad , \key[44]_pad , \key[45]_pad , \key[46]_pad , \key[47]_pad , \key[48]_pad , \key[49]_pad , \key[4]_pad , \key[50]_pad , \key[51]_pad , \key[52]_pad , \key[53]_pad , \key[54]_pad , \key[55]_pad , \key[56]_pad , \key[57]_pad , \key[58]_pad , \key[59]_pad , \key[5]_pad , \key[60]_pad , \key[61]_pad , \key[62]_pad , \key[63]_pad , \key[64]_pad , \key[65]_pad , \key[66]_pad , \key[67]_pad , \key[68]_pad , \key[69]_pad , \key[6]_pad , \key[70]_pad , \key[71]_pad , \key[72]_pad , \key[73]_pad , \key[74]_pad , \key[75]_pad , \key[76]_pad , \key[77]_pad , \key[78]_pad , \key[79]_pad , \key[7]_pad , \key[80]_pad , \key[81]_pad , \key[82]_pad , \key[83]_pad , \key[84]_pad , \key[85]_pad , \key[86]_pad , \key[87]_pad , \key[88]_pad , \key[89]_pad , \key[8]_pad , \key[90]_pad , \key[91]_pad , \key[92]_pad , \key[93]_pad , \key[94]_pad , \key[95]_pad , \key[96]_pad , \key[97]_pad , \key[98]_pad , \key[99]_pad , \key[9]_pad , ld_pad, \ld_r_reg/P0001 , rst_pad, \sa00_reg[0]/P0001 , \sa00_reg[1]/P0001 , \sa00_reg[2]/P0001 , \sa00_reg[3]/P0001 , \sa00_reg[4]/P0001 , \sa00_reg[5]/P0001 , \sa00_reg[6]/NET0131 , \sa00_reg[7]/NET0131 , \sa01_reg[0]/P0001 , \sa01_reg[1]/P0001 , \sa01_reg[2]/P0001 , \sa01_reg[3]/P0001 , \sa01_reg[4]/P0001 , \sa01_reg[5]/P0001 , \sa01_reg[6]/NET0131 , \sa01_reg[7]/NET0131 , \sa02_reg[0]/P0001 , \sa02_reg[1]/P0001 , \sa02_reg[2]/P0001 , \sa02_reg[3]/P0001 , \sa02_reg[4]/P0001 , \sa02_reg[5]/P0001 , \sa02_reg[6]/NET0131 , \sa02_reg[7]/NET0131 , \sa03_reg[0]/P0001 , \sa03_reg[1]/P0001 , \sa03_reg[2]/P0001 , \sa03_reg[3]/P0001 , \sa03_reg[4]/P0001 , \sa03_reg[5]/P0001 , \sa03_reg[6]/NET0131 , \sa03_reg[7]/NET0131 , \sa10_reg[0]/P0001 , \sa10_reg[1]/P0001 , \sa10_reg[2]/P0001 , \sa10_reg[3]/P0001 , \sa10_reg[4]/P0001 , \sa10_reg[5]/P0001 , \sa10_reg[6]/NET0131 , \sa10_reg[7]/NET0131 , \sa11_reg[0]/P0001 , \sa11_reg[1]/P0001 , \sa11_reg[2]/P0001 , \sa11_reg[3]/P0001 , \sa11_reg[4]/P0001 , \sa11_reg[5]/P0001 , \sa11_reg[6]/NET0131 , \sa11_reg[7]/NET0131 , \sa12_reg[0]/P0001 , \sa12_reg[1]/P0001 , \sa12_reg[2]/P0001 , \sa12_reg[3]/P0001 , \sa12_reg[4]/P0001 , \sa12_reg[5]/P0001 , \sa12_reg[6]/NET0131 , \sa12_reg[7]/NET0131 , \sa13_reg[0]/P0001 , \sa13_reg[1]/P0001 , \sa13_reg[2]/P0001 , \sa13_reg[3]/P0001 , \sa13_reg[4]/P0001 , \sa13_reg[5]/P0001 , \sa13_reg[6]/NET0131 , \sa13_reg[7]/NET0131 , \sa20_reg[0]/P0001 , \sa20_reg[1]/P0001 , \sa20_reg[2]/P0001 , \sa20_reg[3]/P0001 , \sa20_reg[4]/P0001 , \sa20_reg[5]/P0001 , \sa20_reg[6]/NET0131 , \sa20_reg[7]/NET0131 , \sa21_reg[0]/P0001 , \sa21_reg[1]/P0001 , \sa21_reg[2]/P0001 , \sa21_reg[3]/P0001 , \sa21_reg[4]/P0001 , \sa21_reg[5]/P0001 , \sa21_reg[6]/NET0131 , \sa21_reg[7]/P0001 , \sa22_reg[0]/P0001 , \sa22_reg[1]/P0001 , \sa22_reg[2]/P0001 , \sa22_reg[3]/P0001 , \sa22_reg[4]/P0001 , \sa22_reg[5]/P0001 , \sa22_reg[6]/NET0131 , \sa22_reg[7]/NET0131 , \sa23_reg[0]/P0001 , \sa23_reg[1]/P0001 , \sa23_reg[2]/P0001 , \sa23_reg[3]/P0001 , \sa23_reg[4]/P0001 , \sa23_reg[5]/P0001 , \sa23_reg[6]/NET0131 , \sa23_reg[7]/NET0131 , \sa30_reg[0]/P0002 , \sa30_reg[1]/P0001 , \sa30_reg[2]/P0001 , \sa30_reg[3]/P0001 , \sa30_reg[4]/P0001 , \sa30_reg[5]/P0001 , \sa30_reg[6]/NET0131 , \sa30_reg[7]/P0001 , \sa31_reg[0]/P0002 , \sa31_reg[1]/P0001 , \sa31_reg[2]/P0001 , \sa31_reg[3]/P0001 , \sa31_reg[4]/P0001 , \sa31_reg[5]/P0001 , \sa31_reg[6]/NET0131 , \sa31_reg[7]/P0001 , \sa32_reg[0]/P0002 , \sa32_reg[1]/P0001 , \sa32_reg[2]/P0001 , \sa32_reg[3]/P0001 , \sa32_reg[4]/P0001 , \sa32_reg[5]/P0001 , \sa32_reg[6]/NET0131 , \sa32_reg[7]/P0001 , \sa33_reg[0]/P0001 , \sa33_reg[1]/P0001 , \sa33_reg[2]/P0001 , \sa33_reg[3]/P0001 , \sa33_reg[4]/P0001 , \sa33_reg[5]/P0001 , \sa33_reg[6]/P0001 , \sa33_reg[7]/NET0131 , \text_in_r_reg[0]/P0001 , \text_in_r_reg[100]/P0001 , \text_in_r_reg[101]/P0001 , \text_in_r_reg[102]/P0001 , \text_in_r_reg[103]/P0001 , \text_in_r_reg[104]/P0001 , \text_in_r_reg[105]/P0001 , \text_in_r_reg[106]/P0001 , \text_in_r_reg[107]/P0001 , \text_in_r_reg[108]/P0001 , \text_in_r_reg[109]/P0001 , \text_in_r_reg[10]/P0001 , \text_in_r_reg[110]/P0001 , \text_in_r_reg[111]/P0001 , \text_in_r_reg[112]/P0001 , \text_in_r_reg[113]/P0001 , \text_in_r_reg[114]/P0001 , \text_in_r_reg[115]/P0001 , \text_in_r_reg[116]/P0001 , \text_in_r_reg[117]/P0001 , \text_in_r_reg[118]/P0001 , \text_in_r_reg[119]/P0001 , \text_in_r_reg[11]/P0001 , \text_in_r_reg[120]/P0001 , \text_in_r_reg[121]/P0001 , \text_in_r_reg[122]/P0001 , \text_in_r_reg[123]/P0001 , \text_in_r_reg[124]/P0001 , \text_in_r_reg[125]/P0001 , \text_in_r_reg[126]/P0001 , \text_in_r_reg[127]/P0001 , \text_in_r_reg[12]/P0001 , \text_in_r_reg[13]/P0001 , \text_in_r_reg[14]/P0001 , \text_in_r_reg[15]/P0001 , \text_in_r_reg[16]/P0001 , \text_in_r_reg[17]/P0001 , \text_in_r_reg[18]/P0001 , \text_in_r_reg[19]/P0001 , \text_in_r_reg[1]/P0001 , \text_in_r_reg[20]/P0001 , \text_in_r_reg[21]/P0001 , \text_in_r_reg[22]/P0001 , \text_in_r_reg[23]/P0001 , \text_in_r_reg[24]/P0001 , \text_in_r_reg[25]/P0001 , \text_in_r_reg[26]/P0001 , \text_in_r_reg[27]/P0001 , \text_in_r_reg[28]/P0001 , \text_in_r_reg[29]/P0001 , \text_in_r_reg[2]/P0001 , \text_in_r_reg[30]/P0001 , \text_in_r_reg[31]/P0001 , \text_in_r_reg[32]/P0001 , \text_in_r_reg[33]/P0001 , \text_in_r_reg[34]/P0001 , \text_in_r_reg[35]/P0001 , \text_in_r_reg[36]/P0001 , \text_in_r_reg[37]/P0001 , \text_in_r_reg[38]/P0001 , \text_in_r_reg[39]/P0001 , \text_in_r_reg[3]/P0001 , \text_in_r_reg[40]/P0001 , \text_in_r_reg[41]/P0001 , \text_in_r_reg[42]/P0001 , \text_in_r_reg[43]/P0001 , \text_in_r_reg[44]/P0001 , \text_in_r_reg[45]/P0001 , \text_in_r_reg[46]/P0001 , \text_in_r_reg[47]/P0001 , \text_in_r_reg[48]/P0001 , \text_in_r_reg[49]/P0001 , \text_in_r_reg[4]/P0001 , \text_in_r_reg[50]/P0001 , \text_in_r_reg[51]/P0001 , \text_in_r_reg[52]/P0001 , \text_in_r_reg[53]/P0001 , \text_in_r_reg[54]/P0001 , \text_in_r_reg[55]/P0001 , \text_in_r_reg[56]/P0001 , \text_in_r_reg[57]/P0001 , \text_in_r_reg[58]/P0001 , \text_in_r_reg[59]/P0001 , \text_in_r_reg[5]/P0001 , \text_in_r_reg[60]/P0001 , \text_in_r_reg[61]/P0001 , \text_in_r_reg[62]/P0001 , \text_in_r_reg[63]/P0001 , \text_in_r_reg[64]/P0001 , \text_in_r_reg[65]/P0001 , \text_in_r_reg[66]/P0001 , \text_in_r_reg[67]/P0001 , \text_in_r_reg[68]/P0001 , \text_in_r_reg[69]/P0001 , \text_in_r_reg[6]/P0001 , \text_in_r_reg[70]/P0001 , \text_in_r_reg[71]/P0001 , \text_in_r_reg[72]/P0001 , \text_in_r_reg[73]/P0001 , \text_in_r_reg[74]/P0001 , \text_in_r_reg[75]/P0001 , \text_in_r_reg[76]/P0001 , \text_in_r_reg[77]/P0001 , \text_in_r_reg[78]/P0001 , \text_in_r_reg[79]/P0001 , \text_in_r_reg[7]/P0001 , \text_in_r_reg[80]/P0001 , \text_in_r_reg[81]/P0001 , \text_in_r_reg[82]/P0001 , \text_in_r_reg[83]/P0001 , \text_in_r_reg[84]/P0001 , \text_in_r_reg[85]/P0001 , \text_in_r_reg[86]/P0001 , \text_in_r_reg[87]/P0001 , \text_in_r_reg[88]/P0001 , \text_in_r_reg[89]/P0001 , \text_in_r_reg[8]/P0001 , \text_in_r_reg[90]/P0001 , \text_in_r_reg[91]/P0001 , \text_in_r_reg[92]/P0001 , \text_in_r_reg[93]/P0001 , \text_in_r_reg[94]/P0001 , \text_in_r_reg[95]/P0001 , \text_in_r_reg[96]/P0001 , \text_in_r_reg[97]/P0001 , \text_in_r_reg[98]/P0001 , \text_in_r_reg[99]/P0001 , \text_in_r_reg[9]/P0001 , \u0_r0_out_reg[24]/P0001 , \u0_r0_out_reg[25]/P0001 , \u0_r0_out_reg[26]/P0001 , \u0_r0_out_reg[27]/P0001 , \u0_r0_out_reg[28]/P0001 , \u0_r0_out_reg[29]/P0001 , \u0_r0_out_reg[30]/P0001 , \u0_r0_out_reg[31]/P0001 , \u0_r0_rcnt_reg[0]/P0001 , \u0_r0_rcnt_reg[1]/P0001 , \u0_r0_rcnt_reg[2]/P0001 , \u0_r0_rcnt_reg[3]/P0001 , \u0_w_reg[0][0]/P0001 , \u0_w_reg[0][10]/P0001 , \u0_w_reg[0][11]/P0001 , \u0_w_reg[0][12]/P0001 , \u0_w_reg[0][13]/P0001 , \u0_w_reg[0][14]/P0001 , \u0_w_reg[0][15]/P0001 , \u0_w_reg[0][16]/P0001 , \u0_w_reg[0][17]/P0001 , \u0_w_reg[0][18]/P0001 , \u0_w_reg[0][19]/P0001 , \u0_w_reg[0][1]/P0001 , \u0_w_reg[0][20]/P0001 , \u0_w_reg[0][21]/P0001 , \u0_w_reg[0][22]/P0001 , \u0_w_reg[0][23]/P0001 , \u0_w_reg[0][24]/P0001 , \u0_w_reg[0][25]/P0001 , \u0_w_reg[0][26]/P0001 , \u0_w_reg[0][27]/P0001 , \u0_w_reg[0][28]/P0001 , \u0_w_reg[0][29]/P0001 , \u0_w_reg[0][2]/P0001 , \u0_w_reg[0][30]/P0001 , \u0_w_reg[0][31]/P0001 , \u0_w_reg[0][3]/P0001 , \u0_w_reg[0][4]/P0001 , \u0_w_reg[0][5]/P0001 , \u0_w_reg[0][6]/P0001 , \u0_w_reg[0][7]/P0001 , \u0_w_reg[0][8]/P0001 , \u0_w_reg[0][9]/P0001 , \u0_w_reg[1][0]/P0001 , \u0_w_reg[1][10]/P0001 , \u0_w_reg[1][11]/P0001 , \u0_w_reg[1][12]/P0001 , \u0_w_reg[1][13]/P0001 , \u0_w_reg[1][14]/P0001 , \u0_w_reg[1][15]/P0001 , \u0_w_reg[1][16]/P0001 , \u0_w_reg[1][17]/P0001 , \u0_w_reg[1][18]/P0001 , \u0_w_reg[1][19]/P0001 , \u0_w_reg[1][1]/P0001 , \u0_w_reg[1][20]/P0001 , \u0_w_reg[1][21]/P0001 , \u0_w_reg[1][22]/P0001 , \u0_w_reg[1][23]/P0001 , \u0_w_reg[1][24]/P0002 , \u0_w_reg[1][25]/P0001 , \u0_w_reg[1][26]/P0001 , \u0_w_reg[1][27]/P0001 , \u0_w_reg[1][28]/P0001 , \u0_w_reg[1][29]/P0002 , \u0_w_reg[1][2]/P0001 , \u0_w_reg[1][30]/P0001 , \u0_w_reg[1][31]/P0001 , \u0_w_reg[1][3]/P0001 , \u0_w_reg[1][4]/P0001 , \u0_w_reg[1][5]/P0001 , \u0_w_reg[1][6]/P0001 , \u0_w_reg[1][7]/P0001 , \u0_w_reg[1][8]/P0001 , \u0_w_reg[1][9]/P0001 , \u0_w_reg[2][0]/P0001 , \u0_w_reg[2][10]/P0001 , \u0_w_reg[2][11]/P0001 , \u0_w_reg[2][12]/P0001 , \u0_w_reg[2][13]/P0001 , \u0_w_reg[2][14]/P0001 , \u0_w_reg[2][15]/P0001 , \u0_w_reg[2][16]/P0001 , \u0_w_reg[2][17]/P0001 , \u0_w_reg[2][18]/P0001 , \u0_w_reg[2][19]/P0001 , \u0_w_reg[2][1]/P0001 , \u0_w_reg[2][20]/P0001 , \u0_w_reg[2][21]/P0001 , \u0_w_reg[2][22]/P0001 , \u0_w_reg[2][23]/P0001 , \u0_w_reg[2][24]/P0001 , \u0_w_reg[2][25]/P0001 , \u0_w_reg[2][26]/P0001 , \u0_w_reg[2][27]/P0001 , \u0_w_reg[2][28]/P0001 , \u0_w_reg[2][29]/P0001 , \u0_w_reg[2][2]/P0001 , \u0_w_reg[2][30]/P0001 , \u0_w_reg[2][31]/P0001 , \u0_w_reg[2][3]/P0001 , \u0_w_reg[2][4]/P0001 , \u0_w_reg[2][5]/P0001 , \u0_w_reg[2][6]/P0001 , \u0_w_reg[2][7]/P0001 , \u0_w_reg[2][8]/P0001 , \u0_w_reg[2][9]/P0001 , \u0_w_reg[3][0]/P0001 , \u0_w_reg[3][10]/P0001 , \u0_w_reg[3][11]/P0001 , \u0_w_reg[3][12]/P0001 , \u0_w_reg[3][13]/P0001 , \u0_w_reg[3][14]/P0001 , \u0_w_reg[3][15]/P0001 , \u0_w_reg[3][16]/P0001 , \u0_w_reg[3][17]/P0001 , \u0_w_reg[3][18]/P0001 , \u0_w_reg[3][19]/P0001 , \u0_w_reg[3][1]/P0001 , \u0_w_reg[3][20]/P0001 , \u0_w_reg[3][21]/P0001 , \u0_w_reg[3][22]/P0001 , \u0_w_reg[3][23]/P0001 , \u0_w_reg[3][24]/P0001 , \u0_w_reg[3][25]/P0001 , \u0_w_reg[3][26]/P0001 , \u0_w_reg[3][27]/P0001 , \u0_w_reg[3][28]/P0001 , \u0_w_reg[3][29]/P0001 , \u0_w_reg[3][2]/P0001 , \u0_w_reg[3][30]/P0001 , \u0_w_reg[3][31]/P0001 , \u0_w_reg[3][3]/P0001 , \u0_w_reg[3][4]/P0001 , \u0_w_reg[3][5]/P0001 , \u0_w_reg[3][6]/P0001 , \u0_w_reg[3][7]/P0001 , \u0_w_reg[3][8]/P0001 , \u0_w_reg[3][9]/P0001 , \_al_n0 , \_al_n1 , \g21/_0_ , \g56610/_0_ , \g56611/_0_ , \g56612/_0_ , \g56613/_0_ , \g56614/_0_ , \g56615/_0_ , \g56616/_0_ , \g56617/_0_ , \g56630/_0_ , \g56631/_0_ , \g56632/_0_ , \g56633/_0_ , \g56634/_0_ , \g56635/_0_ , \g56645/_0_ , \g56646/_0_ , \g56647/_0_ , \g56648/_0_ , \g56649/_0_ , \g56650/_0_ , \g56651/_0_ , \g56652/_0_ , \g56666/_0_ , \g56667/_0_ , \g56668/_0_ , \g56669/_0_ , \g56670/_0_ , \g56671/_0_ , \g56672/_0_ , \g56674/_0_ , \g56675/_0_ , \g56704/_0_ , \g56739/_0_ , \g56743/_0_ , \g56763/_0_ , \g56776/_0_ , \g56812/_0_ , \g56818/_0_ , \g56861/_0_ , \g56874/_0_ , \g56919/_0_ , \g56920/_0_ , \g56921/_0_ , \g56923/_0_ , \g56924/_0_ , \g56925/_0_ , \g56926/_0_ , \g56956/_0_ , \g56957/_0_ , \g56958/_0_ , \g56959/_0_ , \g56960/_0_ , \g56961/_0_ , \g56972/_0_ , \g56973/_0_ , \g56974/_0_ , \g56976/_0_ , \g56977/_0_ , \g56978/_0_ , \g56979/_0_ , \g56980/_0_ , \g57008/_0_ , \g57010/_0_ , \g57011/_0_ , \g57012/_0_ , \g57013/_0_ , \g57014/_0_ , \g57015/_0_ , \g57016/_0_ , \g57017/_0_ , \g57086/_0_ , \g57091/_0_ , \g57114/_0_ , \g57129/_0_ , \g57163/_0_ , \g57171/_0_ , \g57204/_0_ , \g57218/_0_ , \g57262/_0_ , \g57263/_0_ , \g57264/_0_ , \g57265/_0_ , \g57266/_0_ , \g57267/_0_ , \g57268/_0_ , \g57269/_0_ , \g57300/_0_ , \g57301/_0_ , \g57302/_0_ , \g57303/_0_ , \g57304/_0_ , \g57316/_0_ , \g57317/_0_ , \g57319/_0_ , \g57320/_0_ , \g57321/_0_ , \g57322/_0_ , \g57323/_0_ , \g57324/_0_ , \g57350/_0_ , \g57353/_0_ , \g57354/_0_ , \g57355/_0_ , \g57356/_0_ , \g57357/_0_ , \g57358/_0_ , \g57359/_0_ , \g57360/_0_ , \g57427/_0_ , \g57432/_0_ , \g57456/_0_ , \g57471/_0_ , \g57506/_0_ , \g57512/_0_ , \g57540/_0_ , \g57547/_0_ , \g57654/_0_ , \g57655/_0_ , \g57656/_0_ , \g57657/_0_ , \g57658/_0_ , \g57676/_0_ , \g57677/_0_ , \g57678/_0_ , \g57679/_0_ , \g57680/_0_ , \g57681/_0_ , \g57682/_0_ , \g57683/_0_ , \g57684/_0_ , \g57685/_0_ , \g57686/_0_ , \g57687/_0_ , \g57688/_0_ , \g57689/_0_ , \g57690/_0_ , \g57691/_0_ , \g57700/_0_ , \g57701/_0_ , \g57702/_0_ , \g57703/_0_ , \g57704/_0_ , \g57705/_0_ , \g57706/_0_ , \g57707/_0_ , \g57708/_0_ , \g57709/_3_ , \g57710/_3_ , \g57711/_0_ , \g57712/_3_ , \g57715/_3_ , \g57716/_3_ , \g57767/_0_ , \g57768/_3_ , \g57769/_3_ , \g57770/_3_ , \g57771/_3_ , \g57777/_3_ , \g57779/_3_ , \g57804/_3_ , \g57805/_3_ , \g57806/_3_ , \g57807/_3_ , \g57808/_3_ , \g57809/_3_ , \g57810/_3_ , \g57811/_3_ , \g57812/_3_ , \g57813/_3_ , \g57814/_3_ , \g57815/_3_ , \g57816/_0_ , \g57817/_3_ , \g57818/_3_ , \g57819/_3_ , \g57822/_3_ , \g57823/_3_ , \g57824/_3_ , \g57830/_3_ , \g57835/_3_ , \g57836/_3_ , \g57837/_3_ , \g57841/_3_ , \g57842/_3_ , \g57843/_3_ , \g57854/_3_ , \g57855/_3_ , \g57856/_3_ , \g57857/_3_ , \g57858/_3_ , \g57859/_3_ , \g57860/_3_ , \g57861/_3_ , \g57871/_3_ , \g57872/_3_ , \g57874/_3_ , \g57968/_3_ , \g57969/_3_ , \g57970/_3_ , \g57971/_3_ , \g57980/_3_ , \g57983/_3_ , \g57984/_3_ , \g57985/_3_ , \g58012/_3_ , \g58013/_3_ , \g58015/_3_ , \g58057/_3_ , \g58058/_3_ , \g58059/_3_ , \g58189/_3_ , \g58190/_3_ , \g58191/_3_ , \g58192/_3_ , \g58193/_3_ , \g58194/_3_ , \g58195/_3_ , \g58196/_3_ , \g58197/_3_ , \g58224/_3_ , \g58226/_3_ , \g58229/_3_ , \g58255/_3_ , \g58256/_3_ , \g58257/_3_ , \g58258/_3_ , \g58259/_3_ , \g58260/_3_ , \g58261/_3_ , \g58262/_3_ , \g58263/_3_ , \g58264/_3_ , \g58265/_3_ , \g58266/_3_ , \g58267/_3_ , \g58268/_3_ , \g58269/_3_ , \g58270/_0_ , \g58271/_3_ , \g58272/_3_ , \g58273/_3_ , \g58274/_3_ , \g58275/_3_ , \g58276/_3_ , \g58277/_3_ , \g58278/_3_ , \g58279/_3_ , \g58285/_3_ , \g58286/_3_ , \g58288/_3_ , \g58289/_3_ , \g58290/_3_ , \g58292/_3_ , \g58294/_3_ , \g58295/_3_ , \g58297/_3_ , \g58330/_0_ , \g58331/_0_ , \g58332/_0_ , \g58333/_0_ , \g58444/_3_ , \g58445/_3_ , \g58446/_3_ , \g58462/_0_ , \g58506/_0_ , \g58507/_0_ , \g58508/_0_ , \g58509/_0_ , \g58531/_0_ , \g58532/_0_ , \g58533/_0_ , \g58550/_0_ , \g58551/_0_ , \g58552/_0_ , \g58553/_0_ , \g58554/_0_ , \g58555/_0_ , \g58556/_0_ , \g58557/_0_ , \g58558/_0_ , \g58559/_0_ , \g58560/_0_ , \g58600/_3_ , \g58601/_3_ , \g58602/_3_ , \g58603/_3_ , \g58604/_3_ , \g58605/_3_ , \g58606/_3_ , \g58607/_3_ , \g58608/_3_ , \g58611/_0_ , \g58612/_0_ , \g58613/_0_ , \g58614/_0_ , \g58617/_0_ , \g58618/_0_ , \g58619/_0_ , \g58634/_0_ , \g58635/_0_ , \g58636/_0_ , \g58637/_0_ , \g58638/_0_ , \g58639/_0_ , \g58640/_0_ , \g58641/_0_ , \g58829/_3_ , \g58830/_3_ , \g58831/_3_ , \g58832/_3_ , \g58833/_3_ , \g58834/_3_ , \g58835/_0_ , \g58844/_0_ , \g58902/_0_ , \g58903/_0_ , \g58904/_0_ , \g58905/_0_ , \g58910/_0_ , \g58913/_0_ , \g58934/_0_ , \g58935/_0_ , \g58936/_0_ , \g58937/_0_ , \g58938/_0_ , \g58970/_0_ , \g58972/_0_ , \g58994/_0_ , \g58995/_0_ , \g58996/_0_ , \g58997/_0_ , \g58998/_0_ , \g58999/_0_ , \g59000/_0_ , \g59002/_0_ , \g59003/_0_ , \g59004/_0_ , \g59254/_0_ , \g59257/_0_ , \g59258/_0_ , \g59259/_0_ , \g59276/_0_ , \g59277/_0_ , \g59278/_0_ , \g59279/_0_ , \g59280/_0_ , \g59291/_0_ , \g59292/_0_ , \g59293/_0_ , \g59294/_0_ , \g59295/_0_ , \g59308/_0_ , \g59309/_0_ , \g59310/_0_ , \g59311/_0_ , \g59330/_0_ , \g59331/_0_ , \g59332/_0_ , \g59333/_0_ , \g59334/_0_ , \g59335/_0_ , \g59336/_0_ , \g59337/_0_ , \g59338/_0_ , \g59339/_0_ , \g59596/_0_ , \g59597/_0_ , \g59598/_0_ , \g59599/_0_ , \g59625/_0_ , \g59626/_0_ , \g59627/_0_ , \g59628/_0_ , \g59837/_0_ , \g59838/_0_ , \g59839/_0_ , \g59840/_0_ , \g60090/_0_ , \g60320/_0_ , \g60321/_0_ , \g60409/_0_ , \g60539/_0_ , \g60860/_0_ , \g60977/_0_ , \g61012/_0_ , \g61185/_0_ , \g61524/_2_ , \g61776/_0_ , \g61895/_0_ , \g61897/_0_ , \g62220/_0_ , \g65958/_0_ , \g72347/_3_ , \g77848/_0_ , \g85056/_0_ , \sa30_reg[0]/_05_ , \sa31_reg[0]/_05_ , \sa32_reg[0]/_05_ , \u0_w_reg[1][24]/_05_ , \u0_w_reg[1][29]/_05_ );
	input \dcnt_reg[0]/P0001  ;
	input \dcnt_reg[1]/P0001  ;
	input \dcnt_reg[2]/P0001  ;
	input \dcnt_reg[3]/P0001  ;
	input \key[0]_pad  ;
	input \key[100]_pad  ;
	input \key[101]_pad  ;
	input \key[102]_pad  ;
	input \key[103]_pad  ;
	input \key[104]_pad  ;
	input \key[105]_pad  ;
	input \key[106]_pad  ;
	input \key[107]_pad  ;
	input \key[108]_pad  ;
	input \key[109]_pad  ;
	input \key[10]_pad  ;
	input \key[110]_pad  ;
	input \key[111]_pad  ;
	input \key[112]_pad  ;
	input \key[113]_pad  ;
	input \key[114]_pad  ;
	input \key[115]_pad  ;
	input \key[116]_pad  ;
	input \key[117]_pad  ;
	input \key[118]_pad  ;
	input \key[119]_pad  ;
	input \key[11]_pad  ;
	input \key[120]_pad  ;
	input \key[121]_pad  ;
	input \key[122]_pad  ;
	input \key[123]_pad  ;
	input \key[124]_pad  ;
	input \key[125]_pad  ;
	input \key[126]_pad  ;
	input \key[127]_pad  ;
	input \key[12]_pad  ;
	input \key[13]_pad  ;
	input \key[14]_pad  ;
	input \key[15]_pad  ;
	input \key[16]_pad  ;
	input \key[17]_pad  ;
	input \key[18]_pad  ;
	input \key[19]_pad  ;
	input \key[1]_pad  ;
	input \key[20]_pad  ;
	input \key[21]_pad  ;
	input \key[22]_pad  ;
	input \key[23]_pad  ;
	input \key[24]_pad  ;
	input \key[25]_pad  ;
	input \key[26]_pad  ;
	input \key[27]_pad  ;
	input \key[28]_pad  ;
	input \key[29]_pad  ;
	input \key[2]_pad  ;
	input \key[30]_pad  ;
	input \key[31]_pad  ;
	input \key[32]_pad  ;
	input \key[33]_pad  ;
	input \key[34]_pad  ;
	input \key[35]_pad  ;
	input \key[36]_pad  ;
	input \key[37]_pad  ;
	input \key[38]_pad  ;
	input \key[39]_pad  ;
	input \key[3]_pad  ;
	input \key[40]_pad  ;
	input \key[41]_pad  ;
	input \key[42]_pad  ;
	input \key[43]_pad  ;
	input \key[44]_pad  ;
	input \key[45]_pad  ;
	input \key[46]_pad  ;
	input \key[47]_pad  ;
	input \key[48]_pad  ;
	input \key[49]_pad  ;
	input \key[4]_pad  ;
	input \key[50]_pad  ;
	input \key[51]_pad  ;
	input \key[52]_pad  ;
	input \key[53]_pad  ;
	input \key[54]_pad  ;
	input \key[55]_pad  ;
	input \key[56]_pad  ;
	input \key[57]_pad  ;
	input \key[58]_pad  ;
	input \key[59]_pad  ;
	input \key[5]_pad  ;
	input \key[60]_pad  ;
	input \key[61]_pad  ;
	input \key[62]_pad  ;
	input \key[63]_pad  ;
	input \key[64]_pad  ;
	input \key[65]_pad  ;
	input \key[66]_pad  ;
	input \key[67]_pad  ;
	input \key[68]_pad  ;
	input \key[69]_pad  ;
	input \key[6]_pad  ;
	input \key[70]_pad  ;
	input \key[71]_pad  ;
	input \key[72]_pad  ;
	input \key[73]_pad  ;
	input \key[74]_pad  ;
	input \key[75]_pad  ;
	input \key[76]_pad  ;
	input \key[77]_pad  ;
	input \key[78]_pad  ;
	input \key[79]_pad  ;
	input \key[7]_pad  ;
	input \key[80]_pad  ;
	input \key[81]_pad  ;
	input \key[82]_pad  ;
	input \key[83]_pad  ;
	input \key[84]_pad  ;
	input \key[85]_pad  ;
	input \key[86]_pad  ;
	input \key[87]_pad  ;
	input \key[88]_pad  ;
	input \key[89]_pad  ;
	input \key[8]_pad  ;
	input \key[90]_pad  ;
	input \key[91]_pad  ;
	input \key[92]_pad  ;
	input \key[93]_pad  ;
	input \key[94]_pad  ;
	input \key[95]_pad  ;
	input \key[96]_pad  ;
	input \key[97]_pad  ;
	input \key[98]_pad  ;
	input \key[99]_pad  ;
	input \key[9]_pad  ;
	input ld_pad ;
	input \ld_r_reg/P0001  ;
	input rst_pad ;
	input \sa00_reg[0]/P0001  ;
	input \sa00_reg[1]/P0001  ;
	input \sa00_reg[2]/P0001  ;
	input \sa00_reg[3]/P0001  ;
	input \sa00_reg[4]/P0001  ;
	input \sa00_reg[5]/P0001  ;
	input \sa00_reg[6]/NET0131  ;
	input \sa00_reg[7]/NET0131  ;
	input \sa01_reg[0]/P0001  ;
	input \sa01_reg[1]/P0001  ;
	input \sa01_reg[2]/P0001  ;
	input \sa01_reg[3]/P0001  ;
	input \sa01_reg[4]/P0001  ;
	input \sa01_reg[5]/P0001  ;
	input \sa01_reg[6]/NET0131  ;
	input \sa01_reg[7]/NET0131  ;
	input \sa02_reg[0]/P0001  ;
	input \sa02_reg[1]/P0001  ;
	input \sa02_reg[2]/P0001  ;
	input \sa02_reg[3]/P0001  ;
	input \sa02_reg[4]/P0001  ;
	input \sa02_reg[5]/P0001  ;
	input \sa02_reg[6]/NET0131  ;
	input \sa02_reg[7]/NET0131  ;
	input \sa03_reg[0]/P0001  ;
	input \sa03_reg[1]/P0001  ;
	input \sa03_reg[2]/P0001  ;
	input \sa03_reg[3]/P0001  ;
	input \sa03_reg[4]/P0001  ;
	input \sa03_reg[5]/P0001  ;
	input \sa03_reg[6]/NET0131  ;
	input \sa03_reg[7]/NET0131  ;
	input \sa10_reg[0]/P0001  ;
	input \sa10_reg[1]/P0001  ;
	input \sa10_reg[2]/P0001  ;
	input \sa10_reg[3]/P0001  ;
	input \sa10_reg[4]/P0001  ;
	input \sa10_reg[5]/P0001  ;
	input \sa10_reg[6]/NET0131  ;
	input \sa10_reg[7]/NET0131  ;
	input \sa11_reg[0]/P0001  ;
	input \sa11_reg[1]/P0001  ;
	input \sa11_reg[2]/P0001  ;
	input \sa11_reg[3]/P0001  ;
	input \sa11_reg[4]/P0001  ;
	input \sa11_reg[5]/P0001  ;
	input \sa11_reg[6]/NET0131  ;
	input \sa11_reg[7]/NET0131  ;
	input \sa12_reg[0]/P0001  ;
	input \sa12_reg[1]/P0001  ;
	input \sa12_reg[2]/P0001  ;
	input \sa12_reg[3]/P0001  ;
	input \sa12_reg[4]/P0001  ;
	input \sa12_reg[5]/P0001  ;
	input \sa12_reg[6]/NET0131  ;
	input \sa12_reg[7]/NET0131  ;
	input \sa13_reg[0]/P0001  ;
	input \sa13_reg[1]/P0001  ;
	input \sa13_reg[2]/P0001  ;
	input \sa13_reg[3]/P0001  ;
	input \sa13_reg[4]/P0001  ;
	input \sa13_reg[5]/P0001  ;
	input \sa13_reg[6]/NET0131  ;
	input \sa13_reg[7]/NET0131  ;
	input \sa20_reg[0]/P0001  ;
	input \sa20_reg[1]/P0001  ;
	input \sa20_reg[2]/P0001  ;
	input \sa20_reg[3]/P0001  ;
	input \sa20_reg[4]/P0001  ;
	input \sa20_reg[5]/P0001  ;
	input \sa20_reg[6]/NET0131  ;
	input \sa20_reg[7]/NET0131  ;
	input \sa21_reg[0]/P0001  ;
	input \sa21_reg[1]/P0001  ;
	input \sa21_reg[2]/P0001  ;
	input \sa21_reg[3]/P0001  ;
	input \sa21_reg[4]/P0001  ;
	input \sa21_reg[5]/P0001  ;
	input \sa21_reg[6]/NET0131  ;
	input \sa21_reg[7]/P0001  ;
	input \sa22_reg[0]/P0001  ;
	input \sa22_reg[1]/P0001  ;
	input \sa22_reg[2]/P0001  ;
	input \sa22_reg[3]/P0001  ;
	input \sa22_reg[4]/P0001  ;
	input \sa22_reg[5]/P0001  ;
	input \sa22_reg[6]/NET0131  ;
	input \sa22_reg[7]/NET0131  ;
	input \sa23_reg[0]/P0001  ;
	input \sa23_reg[1]/P0001  ;
	input \sa23_reg[2]/P0001  ;
	input \sa23_reg[3]/P0001  ;
	input \sa23_reg[4]/P0001  ;
	input \sa23_reg[5]/P0001  ;
	input \sa23_reg[6]/NET0131  ;
	input \sa23_reg[7]/NET0131  ;
	input \sa30_reg[0]/P0002  ;
	input \sa30_reg[1]/P0001  ;
	input \sa30_reg[2]/P0001  ;
	input \sa30_reg[3]/P0001  ;
	input \sa30_reg[4]/P0001  ;
	input \sa30_reg[5]/P0001  ;
	input \sa30_reg[6]/NET0131  ;
	input \sa30_reg[7]/P0001  ;
	input \sa31_reg[0]/P0002  ;
	input \sa31_reg[1]/P0001  ;
	input \sa31_reg[2]/P0001  ;
	input \sa31_reg[3]/P0001  ;
	input \sa31_reg[4]/P0001  ;
	input \sa31_reg[5]/P0001  ;
	input \sa31_reg[6]/NET0131  ;
	input \sa31_reg[7]/P0001  ;
	input \sa32_reg[0]/P0002  ;
	input \sa32_reg[1]/P0001  ;
	input \sa32_reg[2]/P0001  ;
	input \sa32_reg[3]/P0001  ;
	input \sa32_reg[4]/P0001  ;
	input \sa32_reg[5]/P0001  ;
	input \sa32_reg[6]/NET0131  ;
	input \sa32_reg[7]/P0001  ;
	input \sa33_reg[0]/P0001  ;
	input \sa33_reg[1]/P0001  ;
	input \sa33_reg[2]/P0001  ;
	input \sa33_reg[3]/P0001  ;
	input \sa33_reg[4]/P0001  ;
	input \sa33_reg[5]/P0001  ;
	input \sa33_reg[6]/P0001  ;
	input \sa33_reg[7]/NET0131  ;
	input \text_in_r_reg[0]/P0001  ;
	input \text_in_r_reg[100]/P0001  ;
	input \text_in_r_reg[101]/P0001  ;
	input \text_in_r_reg[102]/P0001  ;
	input \text_in_r_reg[103]/P0001  ;
	input \text_in_r_reg[104]/P0001  ;
	input \text_in_r_reg[105]/P0001  ;
	input \text_in_r_reg[106]/P0001  ;
	input \text_in_r_reg[107]/P0001  ;
	input \text_in_r_reg[108]/P0001  ;
	input \text_in_r_reg[109]/P0001  ;
	input \text_in_r_reg[10]/P0001  ;
	input \text_in_r_reg[110]/P0001  ;
	input \text_in_r_reg[111]/P0001  ;
	input \text_in_r_reg[112]/P0001  ;
	input \text_in_r_reg[113]/P0001  ;
	input \text_in_r_reg[114]/P0001  ;
	input \text_in_r_reg[115]/P0001  ;
	input \text_in_r_reg[116]/P0001  ;
	input \text_in_r_reg[117]/P0001  ;
	input \text_in_r_reg[118]/P0001  ;
	input \text_in_r_reg[119]/P0001  ;
	input \text_in_r_reg[11]/P0001  ;
	input \text_in_r_reg[120]/P0001  ;
	input \text_in_r_reg[121]/P0001  ;
	input \text_in_r_reg[122]/P0001  ;
	input \text_in_r_reg[123]/P0001  ;
	input \text_in_r_reg[124]/P0001  ;
	input \text_in_r_reg[125]/P0001  ;
	input \text_in_r_reg[126]/P0001  ;
	input \text_in_r_reg[127]/P0001  ;
	input \text_in_r_reg[12]/P0001  ;
	input \text_in_r_reg[13]/P0001  ;
	input \text_in_r_reg[14]/P0001  ;
	input \text_in_r_reg[15]/P0001  ;
	input \text_in_r_reg[16]/P0001  ;
	input \text_in_r_reg[17]/P0001  ;
	input \text_in_r_reg[18]/P0001  ;
	input \text_in_r_reg[19]/P0001  ;
	input \text_in_r_reg[1]/P0001  ;
	input \text_in_r_reg[20]/P0001  ;
	input \text_in_r_reg[21]/P0001  ;
	input \text_in_r_reg[22]/P0001  ;
	input \text_in_r_reg[23]/P0001  ;
	input \text_in_r_reg[24]/P0001  ;
	input \text_in_r_reg[25]/P0001  ;
	input \text_in_r_reg[26]/P0001  ;
	input \text_in_r_reg[27]/P0001  ;
	input \text_in_r_reg[28]/P0001  ;
	input \text_in_r_reg[29]/P0001  ;
	input \text_in_r_reg[2]/P0001  ;
	input \text_in_r_reg[30]/P0001  ;
	input \text_in_r_reg[31]/P0001  ;
	input \text_in_r_reg[32]/P0001  ;
	input \text_in_r_reg[33]/P0001  ;
	input \text_in_r_reg[34]/P0001  ;
	input \text_in_r_reg[35]/P0001  ;
	input \text_in_r_reg[36]/P0001  ;
	input \text_in_r_reg[37]/P0001  ;
	input \text_in_r_reg[38]/P0001  ;
	input \text_in_r_reg[39]/P0001  ;
	input \text_in_r_reg[3]/P0001  ;
	input \text_in_r_reg[40]/P0001  ;
	input \text_in_r_reg[41]/P0001  ;
	input \text_in_r_reg[42]/P0001  ;
	input \text_in_r_reg[43]/P0001  ;
	input \text_in_r_reg[44]/P0001  ;
	input \text_in_r_reg[45]/P0001  ;
	input \text_in_r_reg[46]/P0001  ;
	input \text_in_r_reg[47]/P0001  ;
	input \text_in_r_reg[48]/P0001  ;
	input \text_in_r_reg[49]/P0001  ;
	input \text_in_r_reg[4]/P0001  ;
	input \text_in_r_reg[50]/P0001  ;
	input \text_in_r_reg[51]/P0001  ;
	input \text_in_r_reg[52]/P0001  ;
	input \text_in_r_reg[53]/P0001  ;
	input \text_in_r_reg[54]/P0001  ;
	input \text_in_r_reg[55]/P0001  ;
	input \text_in_r_reg[56]/P0001  ;
	input \text_in_r_reg[57]/P0001  ;
	input \text_in_r_reg[58]/P0001  ;
	input \text_in_r_reg[59]/P0001  ;
	input \text_in_r_reg[5]/P0001  ;
	input \text_in_r_reg[60]/P0001  ;
	input \text_in_r_reg[61]/P0001  ;
	input \text_in_r_reg[62]/P0001  ;
	input \text_in_r_reg[63]/P0001  ;
	input \text_in_r_reg[64]/P0001  ;
	input \text_in_r_reg[65]/P0001  ;
	input \text_in_r_reg[66]/P0001  ;
	input \text_in_r_reg[67]/P0001  ;
	input \text_in_r_reg[68]/P0001  ;
	input \text_in_r_reg[69]/P0001  ;
	input \text_in_r_reg[6]/P0001  ;
	input \text_in_r_reg[70]/P0001  ;
	input \text_in_r_reg[71]/P0001  ;
	input \text_in_r_reg[72]/P0001  ;
	input \text_in_r_reg[73]/P0001  ;
	input \text_in_r_reg[74]/P0001  ;
	input \text_in_r_reg[75]/P0001  ;
	input \text_in_r_reg[76]/P0001  ;
	input \text_in_r_reg[77]/P0001  ;
	input \text_in_r_reg[78]/P0001  ;
	input \text_in_r_reg[79]/P0001  ;
	input \text_in_r_reg[7]/P0001  ;
	input \text_in_r_reg[80]/P0001  ;
	input \text_in_r_reg[81]/P0001  ;
	input \text_in_r_reg[82]/P0001  ;
	input \text_in_r_reg[83]/P0001  ;
	input \text_in_r_reg[84]/P0001  ;
	input \text_in_r_reg[85]/P0001  ;
	input \text_in_r_reg[86]/P0001  ;
	input \text_in_r_reg[87]/P0001  ;
	input \text_in_r_reg[88]/P0001  ;
	input \text_in_r_reg[89]/P0001  ;
	input \text_in_r_reg[8]/P0001  ;
	input \text_in_r_reg[90]/P0001  ;
	input \text_in_r_reg[91]/P0001  ;
	input \text_in_r_reg[92]/P0001  ;
	input \text_in_r_reg[93]/P0001  ;
	input \text_in_r_reg[94]/P0001  ;
	input \text_in_r_reg[95]/P0001  ;
	input \text_in_r_reg[96]/P0001  ;
	input \text_in_r_reg[97]/P0001  ;
	input \text_in_r_reg[98]/P0001  ;
	input \text_in_r_reg[99]/P0001  ;
	input \text_in_r_reg[9]/P0001  ;
	input \u0_r0_out_reg[24]/P0001  ;
	input \u0_r0_out_reg[25]/P0001  ;
	input \u0_r0_out_reg[26]/P0001  ;
	input \u0_r0_out_reg[27]/P0001  ;
	input \u0_r0_out_reg[28]/P0001  ;
	input \u0_r0_out_reg[29]/P0001  ;
	input \u0_r0_out_reg[30]/P0001  ;
	input \u0_r0_out_reg[31]/P0001  ;
	input \u0_r0_rcnt_reg[0]/P0001  ;
	input \u0_r0_rcnt_reg[1]/P0001  ;
	input \u0_r0_rcnt_reg[2]/P0001  ;
	input \u0_r0_rcnt_reg[3]/P0001  ;
	input \u0_w_reg[0][0]/P0001  ;
	input \u0_w_reg[0][10]/P0001  ;
	input \u0_w_reg[0][11]/P0001  ;
	input \u0_w_reg[0][12]/P0001  ;
	input \u0_w_reg[0][13]/P0001  ;
	input \u0_w_reg[0][14]/P0001  ;
	input \u0_w_reg[0][15]/P0001  ;
	input \u0_w_reg[0][16]/P0001  ;
	input \u0_w_reg[0][17]/P0001  ;
	input \u0_w_reg[0][18]/P0001  ;
	input \u0_w_reg[0][19]/P0001  ;
	input \u0_w_reg[0][1]/P0001  ;
	input \u0_w_reg[0][20]/P0001  ;
	input \u0_w_reg[0][21]/P0001  ;
	input \u0_w_reg[0][22]/P0001  ;
	input \u0_w_reg[0][23]/P0001  ;
	input \u0_w_reg[0][24]/P0001  ;
	input \u0_w_reg[0][25]/P0001  ;
	input \u0_w_reg[0][26]/P0001  ;
	input \u0_w_reg[0][27]/P0001  ;
	input \u0_w_reg[0][28]/P0001  ;
	input \u0_w_reg[0][29]/P0001  ;
	input \u0_w_reg[0][2]/P0001  ;
	input \u0_w_reg[0][30]/P0001  ;
	input \u0_w_reg[0][31]/P0001  ;
	input \u0_w_reg[0][3]/P0001  ;
	input \u0_w_reg[0][4]/P0001  ;
	input \u0_w_reg[0][5]/P0001  ;
	input \u0_w_reg[0][6]/P0001  ;
	input \u0_w_reg[0][7]/P0001  ;
	input \u0_w_reg[0][8]/P0001  ;
	input \u0_w_reg[0][9]/P0001  ;
	input \u0_w_reg[1][0]/P0001  ;
	input \u0_w_reg[1][10]/P0001  ;
	input \u0_w_reg[1][11]/P0001  ;
	input \u0_w_reg[1][12]/P0001  ;
	input \u0_w_reg[1][13]/P0001  ;
	input \u0_w_reg[1][14]/P0001  ;
	input \u0_w_reg[1][15]/P0001  ;
	input \u0_w_reg[1][16]/P0001  ;
	input \u0_w_reg[1][17]/P0001  ;
	input \u0_w_reg[1][18]/P0001  ;
	input \u0_w_reg[1][19]/P0001  ;
	input \u0_w_reg[1][1]/P0001  ;
	input \u0_w_reg[1][20]/P0001  ;
	input \u0_w_reg[1][21]/P0001  ;
	input \u0_w_reg[1][22]/P0001  ;
	input \u0_w_reg[1][23]/P0001  ;
	input \u0_w_reg[1][24]/P0002  ;
	input \u0_w_reg[1][25]/P0001  ;
	input \u0_w_reg[1][26]/P0001  ;
	input \u0_w_reg[1][27]/P0001  ;
	input \u0_w_reg[1][28]/P0001  ;
	input \u0_w_reg[1][29]/P0002  ;
	input \u0_w_reg[1][2]/P0001  ;
	input \u0_w_reg[1][30]/P0001  ;
	input \u0_w_reg[1][31]/P0001  ;
	input \u0_w_reg[1][3]/P0001  ;
	input \u0_w_reg[1][4]/P0001  ;
	input \u0_w_reg[1][5]/P0001  ;
	input \u0_w_reg[1][6]/P0001  ;
	input \u0_w_reg[1][7]/P0001  ;
	input \u0_w_reg[1][8]/P0001  ;
	input \u0_w_reg[1][9]/P0001  ;
	input \u0_w_reg[2][0]/P0001  ;
	input \u0_w_reg[2][10]/P0001  ;
	input \u0_w_reg[2][11]/P0001  ;
	input \u0_w_reg[2][12]/P0001  ;
	input \u0_w_reg[2][13]/P0001  ;
	input \u0_w_reg[2][14]/P0001  ;
	input \u0_w_reg[2][15]/P0001  ;
	input \u0_w_reg[2][16]/P0001  ;
	input \u0_w_reg[2][17]/P0001  ;
	input \u0_w_reg[2][18]/P0001  ;
	input \u0_w_reg[2][19]/P0001  ;
	input \u0_w_reg[2][1]/P0001  ;
	input \u0_w_reg[2][20]/P0001  ;
	input \u0_w_reg[2][21]/P0001  ;
	input \u0_w_reg[2][22]/P0001  ;
	input \u0_w_reg[2][23]/P0001  ;
	input \u0_w_reg[2][24]/P0001  ;
	input \u0_w_reg[2][25]/P0001  ;
	input \u0_w_reg[2][26]/P0001  ;
	input \u0_w_reg[2][27]/P0001  ;
	input \u0_w_reg[2][28]/P0001  ;
	input \u0_w_reg[2][29]/P0001  ;
	input \u0_w_reg[2][2]/P0001  ;
	input \u0_w_reg[2][30]/P0001  ;
	input \u0_w_reg[2][31]/P0001  ;
	input \u0_w_reg[2][3]/P0001  ;
	input \u0_w_reg[2][4]/P0001  ;
	input \u0_w_reg[2][5]/P0001  ;
	input \u0_w_reg[2][6]/P0001  ;
	input \u0_w_reg[2][7]/P0001  ;
	input \u0_w_reg[2][8]/P0001  ;
	input \u0_w_reg[2][9]/P0001  ;
	input \u0_w_reg[3][0]/P0001  ;
	input \u0_w_reg[3][10]/P0001  ;
	input \u0_w_reg[3][11]/P0001  ;
	input \u0_w_reg[3][12]/P0001  ;
	input \u0_w_reg[3][13]/P0001  ;
	input \u0_w_reg[3][14]/P0001  ;
	input \u0_w_reg[3][15]/P0001  ;
	input \u0_w_reg[3][16]/P0001  ;
	input \u0_w_reg[3][17]/P0001  ;
	input \u0_w_reg[3][18]/P0001  ;
	input \u0_w_reg[3][19]/P0001  ;
	input \u0_w_reg[3][1]/P0001  ;
	input \u0_w_reg[3][20]/P0001  ;
	input \u0_w_reg[3][21]/P0001  ;
	input \u0_w_reg[3][22]/P0001  ;
	input \u0_w_reg[3][23]/P0001  ;
	input \u0_w_reg[3][24]/P0001  ;
	input \u0_w_reg[3][25]/P0001  ;
	input \u0_w_reg[3][26]/P0001  ;
	input \u0_w_reg[3][27]/P0001  ;
	input \u0_w_reg[3][28]/P0001  ;
	input \u0_w_reg[3][29]/P0001  ;
	input \u0_w_reg[3][2]/P0001  ;
	input \u0_w_reg[3][30]/P0001  ;
	input \u0_w_reg[3][31]/P0001  ;
	input \u0_w_reg[3][3]/P0001  ;
	input \u0_w_reg[3][4]/P0001  ;
	input \u0_w_reg[3][5]/P0001  ;
	input \u0_w_reg[3][6]/P0001  ;
	input \u0_w_reg[3][7]/P0001  ;
	input \u0_w_reg[3][8]/P0001  ;
	input \u0_w_reg[3][9]/P0001  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g21/_0_  ;
	output \g56610/_0_  ;
	output \g56611/_0_  ;
	output \g56612/_0_  ;
	output \g56613/_0_  ;
	output \g56614/_0_  ;
	output \g56615/_0_  ;
	output \g56616/_0_  ;
	output \g56617/_0_  ;
	output \g56630/_0_  ;
	output \g56631/_0_  ;
	output \g56632/_0_  ;
	output \g56633/_0_  ;
	output \g56634/_0_  ;
	output \g56635/_0_  ;
	output \g56645/_0_  ;
	output \g56646/_0_  ;
	output \g56647/_0_  ;
	output \g56648/_0_  ;
	output \g56649/_0_  ;
	output \g56650/_0_  ;
	output \g56651/_0_  ;
	output \g56652/_0_  ;
	output \g56666/_0_  ;
	output \g56667/_0_  ;
	output \g56668/_0_  ;
	output \g56669/_0_  ;
	output \g56670/_0_  ;
	output \g56671/_0_  ;
	output \g56672/_0_  ;
	output \g56674/_0_  ;
	output \g56675/_0_  ;
	output \g56704/_0_  ;
	output \g56739/_0_  ;
	output \g56743/_0_  ;
	output \g56763/_0_  ;
	output \g56776/_0_  ;
	output \g56812/_0_  ;
	output \g56818/_0_  ;
	output \g56861/_0_  ;
	output \g56874/_0_  ;
	output \g56919/_0_  ;
	output \g56920/_0_  ;
	output \g56921/_0_  ;
	output \g56923/_0_  ;
	output \g56924/_0_  ;
	output \g56925/_0_  ;
	output \g56926/_0_  ;
	output \g56956/_0_  ;
	output \g56957/_0_  ;
	output \g56958/_0_  ;
	output \g56959/_0_  ;
	output \g56960/_0_  ;
	output \g56961/_0_  ;
	output \g56972/_0_  ;
	output \g56973/_0_  ;
	output \g56974/_0_  ;
	output \g56976/_0_  ;
	output \g56977/_0_  ;
	output \g56978/_0_  ;
	output \g56979/_0_  ;
	output \g56980/_0_  ;
	output \g57008/_0_  ;
	output \g57010/_0_  ;
	output \g57011/_0_  ;
	output \g57012/_0_  ;
	output \g57013/_0_  ;
	output \g57014/_0_  ;
	output \g57015/_0_  ;
	output \g57016/_0_  ;
	output \g57017/_0_  ;
	output \g57086/_0_  ;
	output \g57091/_0_  ;
	output \g57114/_0_  ;
	output \g57129/_0_  ;
	output \g57163/_0_  ;
	output \g57171/_0_  ;
	output \g57204/_0_  ;
	output \g57218/_0_  ;
	output \g57262/_0_  ;
	output \g57263/_0_  ;
	output \g57264/_0_  ;
	output \g57265/_0_  ;
	output \g57266/_0_  ;
	output \g57267/_0_  ;
	output \g57268/_0_  ;
	output \g57269/_0_  ;
	output \g57300/_0_  ;
	output \g57301/_0_  ;
	output \g57302/_0_  ;
	output \g57303/_0_  ;
	output \g57304/_0_  ;
	output \g57316/_0_  ;
	output \g57317/_0_  ;
	output \g57319/_0_  ;
	output \g57320/_0_  ;
	output \g57321/_0_  ;
	output \g57322/_0_  ;
	output \g57323/_0_  ;
	output \g57324/_0_  ;
	output \g57350/_0_  ;
	output \g57353/_0_  ;
	output \g57354/_0_  ;
	output \g57355/_0_  ;
	output \g57356/_0_  ;
	output \g57357/_0_  ;
	output \g57358/_0_  ;
	output \g57359/_0_  ;
	output \g57360/_0_  ;
	output \g57427/_0_  ;
	output \g57432/_0_  ;
	output \g57456/_0_  ;
	output \g57471/_0_  ;
	output \g57506/_0_  ;
	output \g57512/_0_  ;
	output \g57540/_0_  ;
	output \g57547/_0_  ;
	output \g57654/_0_  ;
	output \g57655/_0_  ;
	output \g57656/_0_  ;
	output \g57657/_0_  ;
	output \g57658/_0_  ;
	output \g57676/_0_  ;
	output \g57677/_0_  ;
	output \g57678/_0_  ;
	output \g57679/_0_  ;
	output \g57680/_0_  ;
	output \g57681/_0_  ;
	output \g57682/_0_  ;
	output \g57683/_0_  ;
	output \g57684/_0_  ;
	output \g57685/_0_  ;
	output \g57686/_0_  ;
	output \g57687/_0_  ;
	output \g57688/_0_  ;
	output \g57689/_0_  ;
	output \g57690/_0_  ;
	output \g57691/_0_  ;
	output \g57700/_0_  ;
	output \g57701/_0_  ;
	output \g57702/_0_  ;
	output \g57703/_0_  ;
	output \g57704/_0_  ;
	output \g57705/_0_  ;
	output \g57706/_0_  ;
	output \g57707/_0_  ;
	output \g57708/_0_  ;
	output \g57709/_3_  ;
	output \g57710/_3_  ;
	output \g57711/_0_  ;
	output \g57712/_3_  ;
	output \g57715/_3_  ;
	output \g57716/_3_  ;
	output \g57767/_0_  ;
	output \g57768/_3_  ;
	output \g57769/_3_  ;
	output \g57770/_3_  ;
	output \g57771/_3_  ;
	output \g57777/_3_  ;
	output \g57779/_3_  ;
	output \g57804/_3_  ;
	output \g57805/_3_  ;
	output \g57806/_3_  ;
	output \g57807/_3_  ;
	output \g57808/_3_  ;
	output \g57809/_3_  ;
	output \g57810/_3_  ;
	output \g57811/_3_  ;
	output \g57812/_3_  ;
	output \g57813/_3_  ;
	output \g57814/_3_  ;
	output \g57815/_3_  ;
	output \g57816/_0_  ;
	output \g57817/_3_  ;
	output \g57818/_3_  ;
	output \g57819/_3_  ;
	output \g57822/_3_  ;
	output \g57823/_3_  ;
	output \g57824/_3_  ;
	output \g57830/_3_  ;
	output \g57835/_3_  ;
	output \g57836/_3_  ;
	output \g57837/_3_  ;
	output \g57841/_3_  ;
	output \g57842/_3_  ;
	output \g57843/_3_  ;
	output \g57854/_3_  ;
	output \g57855/_3_  ;
	output \g57856/_3_  ;
	output \g57857/_3_  ;
	output \g57858/_3_  ;
	output \g57859/_3_  ;
	output \g57860/_3_  ;
	output \g57861/_3_  ;
	output \g57871/_3_  ;
	output \g57872/_3_  ;
	output \g57874/_3_  ;
	output \g57968/_3_  ;
	output \g57969/_3_  ;
	output \g57970/_3_  ;
	output \g57971/_3_  ;
	output \g57980/_3_  ;
	output \g57983/_3_  ;
	output \g57984/_3_  ;
	output \g57985/_3_  ;
	output \g58012/_3_  ;
	output \g58013/_3_  ;
	output \g58015/_3_  ;
	output \g58057/_3_  ;
	output \g58058/_3_  ;
	output \g58059/_3_  ;
	output \g58189/_3_  ;
	output \g58190/_3_  ;
	output \g58191/_3_  ;
	output \g58192/_3_  ;
	output \g58193/_3_  ;
	output \g58194/_3_  ;
	output \g58195/_3_  ;
	output \g58196/_3_  ;
	output \g58197/_3_  ;
	output \g58224/_3_  ;
	output \g58226/_3_  ;
	output \g58229/_3_  ;
	output \g58255/_3_  ;
	output \g58256/_3_  ;
	output \g58257/_3_  ;
	output \g58258/_3_  ;
	output \g58259/_3_  ;
	output \g58260/_3_  ;
	output \g58261/_3_  ;
	output \g58262/_3_  ;
	output \g58263/_3_  ;
	output \g58264/_3_  ;
	output \g58265/_3_  ;
	output \g58266/_3_  ;
	output \g58267/_3_  ;
	output \g58268/_3_  ;
	output \g58269/_3_  ;
	output \g58270/_0_  ;
	output \g58271/_3_  ;
	output \g58272/_3_  ;
	output \g58273/_3_  ;
	output \g58274/_3_  ;
	output \g58275/_3_  ;
	output \g58276/_3_  ;
	output \g58277/_3_  ;
	output \g58278/_3_  ;
	output \g58279/_3_  ;
	output \g58285/_3_  ;
	output \g58286/_3_  ;
	output \g58288/_3_  ;
	output \g58289/_3_  ;
	output \g58290/_3_  ;
	output \g58292/_3_  ;
	output \g58294/_3_  ;
	output \g58295/_3_  ;
	output \g58297/_3_  ;
	output \g58330/_0_  ;
	output \g58331/_0_  ;
	output \g58332/_0_  ;
	output \g58333/_0_  ;
	output \g58444/_3_  ;
	output \g58445/_3_  ;
	output \g58446/_3_  ;
	output \g58462/_0_  ;
	output \g58506/_0_  ;
	output \g58507/_0_  ;
	output \g58508/_0_  ;
	output \g58509/_0_  ;
	output \g58531/_0_  ;
	output \g58532/_0_  ;
	output \g58533/_0_  ;
	output \g58550/_0_  ;
	output \g58551/_0_  ;
	output \g58552/_0_  ;
	output \g58553/_0_  ;
	output \g58554/_0_  ;
	output \g58555/_0_  ;
	output \g58556/_0_  ;
	output \g58557/_0_  ;
	output \g58558/_0_  ;
	output \g58559/_0_  ;
	output \g58560/_0_  ;
	output \g58600/_3_  ;
	output \g58601/_3_  ;
	output \g58602/_3_  ;
	output \g58603/_3_  ;
	output \g58604/_3_  ;
	output \g58605/_3_  ;
	output \g58606/_3_  ;
	output \g58607/_3_  ;
	output \g58608/_3_  ;
	output \g58611/_0_  ;
	output \g58612/_0_  ;
	output \g58613/_0_  ;
	output \g58614/_0_  ;
	output \g58617/_0_  ;
	output \g58618/_0_  ;
	output \g58619/_0_  ;
	output \g58634/_0_  ;
	output \g58635/_0_  ;
	output \g58636/_0_  ;
	output \g58637/_0_  ;
	output \g58638/_0_  ;
	output \g58639/_0_  ;
	output \g58640/_0_  ;
	output \g58641/_0_  ;
	output \g58829/_3_  ;
	output \g58830/_3_  ;
	output \g58831/_3_  ;
	output \g58832/_3_  ;
	output \g58833/_3_  ;
	output \g58834/_3_  ;
	output \g58835/_0_  ;
	output \g58844/_0_  ;
	output \g58902/_0_  ;
	output \g58903/_0_  ;
	output \g58904/_0_  ;
	output \g58905/_0_  ;
	output \g58910/_0_  ;
	output \g58913/_0_  ;
	output \g58934/_0_  ;
	output \g58935/_0_  ;
	output \g58936/_0_  ;
	output \g58937/_0_  ;
	output \g58938/_0_  ;
	output \g58970/_0_  ;
	output \g58972/_0_  ;
	output \g58994/_0_  ;
	output \g58995/_0_  ;
	output \g58996/_0_  ;
	output \g58997/_0_  ;
	output \g58998/_0_  ;
	output \g58999/_0_  ;
	output \g59000/_0_  ;
	output \g59002/_0_  ;
	output \g59003/_0_  ;
	output \g59004/_0_  ;
	output \g59254/_0_  ;
	output \g59257/_0_  ;
	output \g59258/_0_  ;
	output \g59259/_0_  ;
	output \g59276/_0_  ;
	output \g59277/_0_  ;
	output \g59278/_0_  ;
	output \g59279/_0_  ;
	output \g59280/_0_  ;
	output \g59291/_0_  ;
	output \g59292/_0_  ;
	output \g59293/_0_  ;
	output \g59294/_0_  ;
	output \g59295/_0_  ;
	output \g59308/_0_  ;
	output \g59309/_0_  ;
	output \g59310/_0_  ;
	output \g59311/_0_  ;
	output \g59330/_0_  ;
	output \g59331/_0_  ;
	output \g59332/_0_  ;
	output \g59333/_0_  ;
	output \g59334/_0_  ;
	output \g59335/_0_  ;
	output \g59336/_0_  ;
	output \g59337/_0_  ;
	output \g59338/_0_  ;
	output \g59339/_0_  ;
	output \g59596/_0_  ;
	output \g59597/_0_  ;
	output \g59598/_0_  ;
	output \g59599/_0_  ;
	output \g59625/_0_  ;
	output \g59626/_0_  ;
	output \g59627/_0_  ;
	output \g59628/_0_  ;
	output \g59837/_0_  ;
	output \g59838/_0_  ;
	output \g59839/_0_  ;
	output \g59840/_0_  ;
	output \g60090/_0_  ;
	output \g60320/_0_  ;
	output \g60321/_0_  ;
	output \g60409/_0_  ;
	output \g60539/_0_  ;
	output \g60860/_0_  ;
	output \g60977/_0_  ;
	output \g61012/_0_  ;
	output \g61185/_0_  ;
	output \g61524/_2_  ;
	output \g61776/_0_  ;
	output \g61895/_0_  ;
	output \g61897/_0_  ;
	output \g62220/_0_  ;
	output \g65958/_0_  ;
	output \g72347/_3_  ;
	output \g77848/_0_  ;
	output \g85056/_0_  ;
	output \sa30_reg[0]/_05_  ;
	output \sa31_reg[0]/_05_  ;
	output \sa32_reg[0]/_05_  ;
	output \u0_w_reg[1][24]/_05_  ;
	output \u0_w_reg[1][29]/_05_  ;
	wire _w19967_ ;
	wire _w19966_ ;
	wire _w19965_ ;
	wire _w19964_ ;
	wire _w19963_ ;
	wire _w19962_ ;
	wire _w19961_ ;
	wire _w19960_ ;
	wire _w19959_ ;
	wire _w19958_ ;
	wire _w19957_ ;
	wire _w19956_ ;
	wire _w19955_ ;
	wire _w19954_ ;
	wire _w19953_ ;
	wire _w19952_ ;
	wire _w19951_ ;
	wire _w19950_ ;
	wire _w19949_ ;
	wire _w19948_ ;
	wire _w19947_ ;
	wire _w19946_ ;
	wire _w19945_ ;
	wire _w19944_ ;
	wire _w19943_ ;
	wire _w19942_ ;
	wire _w19941_ ;
	wire _w19940_ ;
	wire _w19939_ ;
	wire _w19938_ ;
	wire _w19937_ ;
	wire _w19936_ ;
	wire _w19935_ ;
	wire _w19934_ ;
	wire _w19933_ ;
	wire _w19932_ ;
	wire _w19931_ ;
	wire _w19930_ ;
	wire _w19929_ ;
	wire _w19928_ ;
	wire _w19927_ ;
	wire _w19926_ ;
	wire _w19925_ ;
	wire _w19924_ ;
	wire _w19923_ ;
	wire _w19922_ ;
	wire _w19921_ ;
	wire _w19920_ ;
	wire _w19919_ ;
	wire _w19918_ ;
	wire _w19917_ ;
	wire _w19916_ ;
	wire _w19915_ ;
	wire _w19914_ ;
	wire _w19913_ ;
	wire _w19912_ ;
	wire _w19911_ ;
	wire _w19910_ ;
	wire _w19909_ ;
	wire _w19908_ ;
	wire _w19907_ ;
	wire _w19906_ ;
	wire _w19905_ ;
	wire _w19904_ ;
	wire _w19903_ ;
	wire _w19902_ ;
	wire _w19901_ ;
	wire _w19900_ ;
	wire _w19899_ ;
	wire _w19898_ ;
	wire _w19897_ ;
	wire _w19896_ ;
	wire _w19895_ ;
	wire _w19894_ ;
	wire _w19893_ ;
	wire _w19892_ ;
	wire _w19891_ ;
	wire _w19890_ ;
	wire _w19889_ ;
	wire _w19888_ ;
	wire _w19887_ ;
	wire _w19886_ ;
	wire _w19885_ ;
	wire _w19884_ ;
	wire _w19883_ ;
	wire _w19882_ ;
	wire _w19881_ ;
	wire _w19880_ ;
	wire _w19879_ ;
	wire _w19878_ ;
	wire _w19877_ ;
	wire _w19876_ ;
	wire _w19875_ ;
	wire _w19874_ ;
	wire _w19873_ ;
	wire _w19872_ ;
	wire _w19871_ ;
	wire _w19870_ ;
	wire _w19869_ ;
	wire _w19868_ ;
	wire _w19867_ ;
	wire _w19866_ ;
	wire _w19865_ ;
	wire _w19864_ ;
	wire _w19863_ ;
	wire _w19862_ ;
	wire _w19861_ ;
	wire _w19860_ ;
	wire _w19859_ ;
	wire _w19858_ ;
	wire _w19857_ ;
	wire _w19856_ ;
	wire _w19855_ ;
	wire _w19854_ ;
	wire _w19853_ ;
	wire _w19852_ ;
	wire _w19851_ ;
	wire _w19850_ ;
	wire _w19849_ ;
	wire _w19848_ ;
	wire _w19847_ ;
	wire _w19846_ ;
	wire _w19845_ ;
	wire _w19844_ ;
	wire _w19843_ ;
	wire _w19842_ ;
	wire _w19841_ ;
	wire _w19840_ ;
	wire _w19839_ ;
	wire _w19838_ ;
	wire _w19837_ ;
	wire _w19836_ ;
	wire _w19835_ ;
	wire _w19834_ ;
	wire _w19833_ ;
	wire _w19832_ ;
	wire _w19831_ ;
	wire _w19830_ ;
	wire _w19829_ ;
	wire _w19828_ ;
	wire _w19827_ ;
	wire _w19826_ ;
	wire _w19825_ ;
	wire _w19824_ ;
	wire _w19823_ ;
	wire _w19822_ ;
	wire _w19821_ ;
	wire _w19820_ ;
	wire _w19819_ ;
	wire _w19818_ ;
	wire _w19817_ ;
	wire _w19816_ ;
	wire _w19815_ ;
	wire _w19814_ ;
	wire _w19813_ ;
	wire _w19812_ ;
	wire _w19811_ ;
	wire _w19810_ ;
	wire _w19809_ ;
	wire _w19808_ ;
	wire _w19807_ ;
	wire _w19806_ ;
	wire _w19805_ ;
	wire _w19804_ ;
	wire _w19803_ ;
	wire _w19802_ ;
	wire _w19801_ ;
	wire _w19800_ ;
	wire _w19799_ ;
	wire _w19798_ ;
	wire _w19797_ ;
	wire _w19796_ ;
	wire _w19795_ ;
	wire _w19794_ ;
	wire _w19793_ ;
	wire _w19792_ ;
	wire _w19791_ ;
	wire _w19790_ ;
	wire _w19789_ ;
	wire _w19788_ ;
	wire _w19787_ ;
	wire _w19786_ ;
	wire _w19785_ ;
	wire _w19784_ ;
	wire _w19783_ ;
	wire _w19782_ ;
	wire _w19781_ ;
	wire _w19780_ ;
	wire _w19779_ ;
	wire _w19778_ ;
	wire _w19777_ ;
	wire _w19776_ ;
	wire _w19775_ ;
	wire _w19774_ ;
	wire _w19773_ ;
	wire _w19772_ ;
	wire _w19771_ ;
	wire _w19770_ ;
	wire _w19769_ ;
	wire _w19768_ ;
	wire _w19767_ ;
	wire _w19766_ ;
	wire _w19765_ ;
	wire _w19764_ ;
	wire _w19763_ ;
	wire _w19762_ ;
	wire _w19761_ ;
	wire _w19760_ ;
	wire _w19759_ ;
	wire _w19758_ ;
	wire _w19757_ ;
	wire _w19756_ ;
	wire _w19755_ ;
	wire _w19754_ ;
	wire _w19753_ ;
	wire _w19752_ ;
	wire _w19751_ ;
	wire _w19750_ ;
	wire _w19749_ ;
	wire _w19748_ ;
	wire _w19747_ ;
	wire _w19746_ ;
	wire _w19745_ ;
	wire _w19744_ ;
	wire _w19743_ ;
	wire _w19742_ ;
	wire _w19741_ ;
	wire _w19740_ ;
	wire _w19739_ ;
	wire _w19738_ ;
	wire _w19737_ ;
	wire _w19736_ ;
	wire _w19735_ ;
	wire _w19734_ ;
	wire _w19733_ ;
	wire _w19732_ ;
	wire _w19731_ ;
	wire _w19730_ ;
	wire _w19729_ ;
	wire _w19728_ ;
	wire _w19727_ ;
	wire _w19726_ ;
	wire _w19725_ ;
	wire _w19724_ ;
	wire _w19723_ ;
	wire _w19722_ ;
	wire _w19721_ ;
	wire _w19720_ ;
	wire _w19719_ ;
	wire _w19718_ ;
	wire _w19717_ ;
	wire _w19716_ ;
	wire _w19715_ ;
	wire _w19714_ ;
	wire _w19713_ ;
	wire _w19712_ ;
	wire _w19711_ ;
	wire _w19710_ ;
	wire _w19709_ ;
	wire _w19708_ ;
	wire _w19707_ ;
	wire _w19706_ ;
	wire _w19705_ ;
	wire _w19704_ ;
	wire _w19703_ ;
	wire _w19702_ ;
	wire _w19701_ ;
	wire _w19700_ ;
	wire _w19699_ ;
	wire _w19698_ ;
	wire _w19697_ ;
	wire _w19696_ ;
	wire _w19695_ ;
	wire _w19694_ ;
	wire _w19693_ ;
	wire _w19692_ ;
	wire _w19691_ ;
	wire _w19690_ ;
	wire _w19689_ ;
	wire _w19688_ ;
	wire _w19687_ ;
	wire _w19686_ ;
	wire _w19685_ ;
	wire _w19684_ ;
	wire _w19683_ ;
	wire _w19682_ ;
	wire _w19681_ ;
	wire _w19680_ ;
	wire _w19679_ ;
	wire _w19678_ ;
	wire _w19677_ ;
	wire _w19676_ ;
	wire _w19675_ ;
	wire _w19674_ ;
	wire _w19673_ ;
	wire _w19672_ ;
	wire _w19671_ ;
	wire _w19670_ ;
	wire _w19669_ ;
	wire _w19668_ ;
	wire _w19667_ ;
	wire _w19666_ ;
	wire _w19665_ ;
	wire _w19664_ ;
	wire _w19663_ ;
	wire _w19662_ ;
	wire _w19661_ ;
	wire _w19660_ ;
	wire _w19659_ ;
	wire _w19658_ ;
	wire _w19657_ ;
	wire _w19656_ ;
	wire _w19655_ ;
	wire _w19654_ ;
	wire _w19653_ ;
	wire _w19652_ ;
	wire _w19651_ ;
	wire _w19650_ ;
	wire _w19649_ ;
	wire _w19648_ ;
	wire _w19647_ ;
	wire _w19646_ ;
	wire _w19645_ ;
	wire _w19644_ ;
	wire _w19643_ ;
	wire _w19642_ ;
	wire _w19641_ ;
	wire _w19640_ ;
	wire _w19639_ ;
	wire _w19638_ ;
	wire _w19637_ ;
	wire _w19636_ ;
	wire _w19635_ ;
	wire _w19634_ ;
	wire _w19633_ ;
	wire _w19632_ ;
	wire _w19631_ ;
	wire _w19630_ ;
	wire _w19629_ ;
	wire _w19628_ ;
	wire _w19627_ ;
	wire _w19626_ ;
	wire _w19625_ ;
	wire _w19624_ ;
	wire _w19623_ ;
	wire _w19622_ ;
	wire _w19621_ ;
	wire _w19620_ ;
	wire _w19619_ ;
	wire _w19618_ ;
	wire _w19617_ ;
	wire _w19616_ ;
	wire _w19615_ ;
	wire _w19614_ ;
	wire _w19613_ ;
	wire _w19612_ ;
	wire _w19611_ ;
	wire _w19610_ ;
	wire _w19609_ ;
	wire _w19608_ ;
	wire _w19607_ ;
	wire _w19606_ ;
	wire _w19605_ ;
	wire _w19604_ ;
	wire _w19603_ ;
	wire _w19602_ ;
	wire _w19601_ ;
	wire _w19600_ ;
	wire _w19599_ ;
	wire _w19598_ ;
	wire _w19597_ ;
	wire _w19596_ ;
	wire _w19595_ ;
	wire _w19594_ ;
	wire _w19593_ ;
	wire _w19592_ ;
	wire _w19591_ ;
	wire _w19590_ ;
	wire _w19589_ ;
	wire _w19588_ ;
	wire _w19587_ ;
	wire _w19586_ ;
	wire _w19585_ ;
	wire _w19584_ ;
	wire _w19583_ ;
	wire _w19582_ ;
	wire _w19581_ ;
	wire _w19580_ ;
	wire _w19579_ ;
	wire _w19578_ ;
	wire _w19577_ ;
	wire _w19576_ ;
	wire _w19575_ ;
	wire _w19574_ ;
	wire _w19573_ ;
	wire _w19572_ ;
	wire _w19571_ ;
	wire _w19570_ ;
	wire _w19569_ ;
	wire _w19568_ ;
	wire _w19567_ ;
	wire _w19566_ ;
	wire _w19565_ ;
	wire _w19564_ ;
	wire _w19563_ ;
	wire _w19562_ ;
	wire _w19561_ ;
	wire _w19560_ ;
	wire _w19559_ ;
	wire _w19558_ ;
	wire _w19557_ ;
	wire _w19556_ ;
	wire _w19555_ ;
	wire _w19554_ ;
	wire _w19553_ ;
	wire _w19552_ ;
	wire _w19551_ ;
	wire _w19550_ ;
	wire _w19549_ ;
	wire _w19548_ ;
	wire _w19547_ ;
	wire _w19546_ ;
	wire _w19545_ ;
	wire _w19544_ ;
	wire _w19543_ ;
	wire _w19542_ ;
	wire _w19541_ ;
	wire _w19540_ ;
	wire _w19539_ ;
	wire _w19538_ ;
	wire _w19537_ ;
	wire _w19536_ ;
	wire _w19535_ ;
	wire _w19534_ ;
	wire _w19533_ ;
	wire _w19532_ ;
	wire _w19531_ ;
	wire _w19530_ ;
	wire _w19529_ ;
	wire _w19528_ ;
	wire _w19527_ ;
	wire _w19526_ ;
	wire _w19525_ ;
	wire _w19524_ ;
	wire _w19523_ ;
	wire _w19522_ ;
	wire _w19521_ ;
	wire _w19520_ ;
	wire _w19519_ ;
	wire _w19518_ ;
	wire _w19517_ ;
	wire _w19516_ ;
	wire _w19515_ ;
	wire _w19514_ ;
	wire _w19513_ ;
	wire _w19512_ ;
	wire _w19511_ ;
	wire _w19510_ ;
	wire _w19509_ ;
	wire _w19508_ ;
	wire _w19507_ ;
	wire _w19506_ ;
	wire _w19505_ ;
	wire _w19504_ ;
	wire _w19503_ ;
	wire _w19502_ ;
	wire _w19501_ ;
	wire _w19500_ ;
	wire _w19499_ ;
	wire _w19498_ ;
	wire _w19497_ ;
	wire _w19496_ ;
	wire _w19495_ ;
	wire _w19494_ ;
	wire _w19493_ ;
	wire _w19492_ ;
	wire _w19491_ ;
	wire _w19490_ ;
	wire _w19489_ ;
	wire _w19488_ ;
	wire _w19487_ ;
	wire _w19486_ ;
	wire _w19485_ ;
	wire _w19484_ ;
	wire _w19483_ ;
	wire _w19482_ ;
	wire _w19481_ ;
	wire _w19480_ ;
	wire _w19479_ ;
	wire _w19478_ ;
	wire _w19477_ ;
	wire _w19476_ ;
	wire _w19475_ ;
	wire _w19474_ ;
	wire _w19473_ ;
	wire _w19472_ ;
	wire _w19471_ ;
	wire _w19470_ ;
	wire _w19469_ ;
	wire _w19468_ ;
	wire _w19467_ ;
	wire _w19466_ ;
	wire _w19465_ ;
	wire _w19464_ ;
	wire _w19463_ ;
	wire _w19462_ ;
	wire _w19461_ ;
	wire _w19460_ ;
	wire _w19459_ ;
	wire _w19458_ ;
	wire _w19457_ ;
	wire _w19456_ ;
	wire _w19455_ ;
	wire _w19454_ ;
	wire _w19453_ ;
	wire _w19452_ ;
	wire _w19451_ ;
	wire _w19450_ ;
	wire _w19449_ ;
	wire _w19448_ ;
	wire _w19447_ ;
	wire _w19446_ ;
	wire _w19445_ ;
	wire _w19444_ ;
	wire _w19443_ ;
	wire _w19442_ ;
	wire _w19441_ ;
	wire _w19440_ ;
	wire _w19439_ ;
	wire _w19438_ ;
	wire _w19437_ ;
	wire _w19436_ ;
	wire _w19435_ ;
	wire _w19434_ ;
	wire _w19433_ ;
	wire _w19432_ ;
	wire _w19431_ ;
	wire _w19430_ ;
	wire _w19429_ ;
	wire _w19428_ ;
	wire _w19427_ ;
	wire _w19426_ ;
	wire _w19425_ ;
	wire _w19424_ ;
	wire _w19423_ ;
	wire _w19422_ ;
	wire _w19421_ ;
	wire _w19420_ ;
	wire _w19419_ ;
	wire _w19418_ ;
	wire _w19417_ ;
	wire _w19416_ ;
	wire _w19415_ ;
	wire _w19414_ ;
	wire _w19413_ ;
	wire _w19412_ ;
	wire _w19411_ ;
	wire _w19410_ ;
	wire _w19409_ ;
	wire _w19408_ ;
	wire _w19407_ ;
	wire _w19406_ ;
	wire _w19405_ ;
	wire _w19404_ ;
	wire _w19403_ ;
	wire _w19402_ ;
	wire _w19401_ ;
	wire _w19400_ ;
	wire _w19399_ ;
	wire _w19398_ ;
	wire _w19397_ ;
	wire _w19396_ ;
	wire _w19395_ ;
	wire _w19394_ ;
	wire _w19393_ ;
	wire _w19392_ ;
	wire _w19391_ ;
	wire _w19390_ ;
	wire _w19389_ ;
	wire _w19388_ ;
	wire _w19387_ ;
	wire _w19386_ ;
	wire _w19385_ ;
	wire _w19384_ ;
	wire _w19383_ ;
	wire _w19382_ ;
	wire _w19381_ ;
	wire _w19380_ ;
	wire _w19379_ ;
	wire _w19378_ ;
	wire _w19377_ ;
	wire _w19376_ ;
	wire _w19375_ ;
	wire _w19374_ ;
	wire _w19373_ ;
	wire _w19372_ ;
	wire _w19371_ ;
	wire _w19370_ ;
	wire _w19369_ ;
	wire _w19368_ ;
	wire _w19367_ ;
	wire _w19366_ ;
	wire _w19365_ ;
	wire _w19364_ ;
	wire _w19363_ ;
	wire _w19362_ ;
	wire _w19361_ ;
	wire _w19360_ ;
	wire _w19359_ ;
	wire _w19358_ ;
	wire _w19357_ ;
	wire _w19356_ ;
	wire _w19355_ ;
	wire _w19354_ ;
	wire _w19353_ ;
	wire _w19352_ ;
	wire _w19351_ ;
	wire _w19350_ ;
	wire _w19349_ ;
	wire _w19348_ ;
	wire _w19347_ ;
	wire _w19346_ ;
	wire _w19345_ ;
	wire _w19344_ ;
	wire _w19343_ ;
	wire _w19342_ ;
	wire _w19341_ ;
	wire _w19340_ ;
	wire _w19339_ ;
	wire _w19338_ ;
	wire _w19337_ ;
	wire _w19336_ ;
	wire _w19335_ ;
	wire _w19334_ ;
	wire _w19333_ ;
	wire _w19332_ ;
	wire _w19331_ ;
	wire _w19330_ ;
	wire _w19329_ ;
	wire _w19328_ ;
	wire _w19327_ ;
	wire _w19326_ ;
	wire _w19325_ ;
	wire _w19324_ ;
	wire _w19323_ ;
	wire _w19322_ ;
	wire _w19321_ ;
	wire _w19320_ ;
	wire _w19319_ ;
	wire _w19318_ ;
	wire _w19317_ ;
	wire _w19316_ ;
	wire _w19315_ ;
	wire _w19314_ ;
	wire _w19313_ ;
	wire _w19312_ ;
	wire _w19311_ ;
	wire _w19310_ ;
	wire _w19309_ ;
	wire _w19308_ ;
	wire _w19307_ ;
	wire _w19306_ ;
	wire _w19305_ ;
	wire _w19304_ ;
	wire _w19303_ ;
	wire _w19302_ ;
	wire _w19301_ ;
	wire _w19300_ ;
	wire _w19299_ ;
	wire _w19298_ ;
	wire _w19297_ ;
	wire _w19296_ ;
	wire _w19295_ ;
	wire _w19294_ ;
	wire _w19293_ ;
	wire _w19292_ ;
	wire _w19291_ ;
	wire _w19290_ ;
	wire _w19289_ ;
	wire _w19288_ ;
	wire _w19287_ ;
	wire _w19286_ ;
	wire _w19285_ ;
	wire _w19284_ ;
	wire _w19283_ ;
	wire _w19282_ ;
	wire _w19281_ ;
	wire _w19280_ ;
	wire _w19279_ ;
	wire _w19278_ ;
	wire _w19277_ ;
	wire _w19276_ ;
	wire _w19275_ ;
	wire _w19274_ ;
	wire _w19273_ ;
	wire _w19272_ ;
	wire _w19271_ ;
	wire _w19270_ ;
	wire _w19269_ ;
	wire _w19268_ ;
	wire _w19267_ ;
	wire _w19266_ ;
	wire _w19265_ ;
	wire _w19264_ ;
	wire _w19263_ ;
	wire _w19262_ ;
	wire _w19261_ ;
	wire _w19260_ ;
	wire _w19259_ ;
	wire _w19258_ ;
	wire _w19257_ ;
	wire _w19256_ ;
	wire _w19255_ ;
	wire _w19254_ ;
	wire _w19253_ ;
	wire _w19252_ ;
	wire _w19251_ ;
	wire _w19250_ ;
	wire _w19249_ ;
	wire _w19248_ ;
	wire _w19247_ ;
	wire _w19246_ ;
	wire _w19245_ ;
	wire _w19244_ ;
	wire _w19243_ ;
	wire _w19242_ ;
	wire _w19241_ ;
	wire _w19240_ ;
	wire _w19239_ ;
	wire _w19238_ ;
	wire _w19237_ ;
	wire _w19236_ ;
	wire _w19235_ ;
	wire _w19234_ ;
	wire _w19233_ ;
	wire _w19232_ ;
	wire _w19231_ ;
	wire _w19230_ ;
	wire _w19229_ ;
	wire _w19228_ ;
	wire _w19227_ ;
	wire _w19226_ ;
	wire _w19225_ ;
	wire _w19224_ ;
	wire _w19223_ ;
	wire _w19222_ ;
	wire _w19221_ ;
	wire _w19220_ ;
	wire _w19219_ ;
	wire _w19218_ ;
	wire _w19217_ ;
	wire _w19216_ ;
	wire _w19215_ ;
	wire _w19214_ ;
	wire _w19213_ ;
	wire _w19212_ ;
	wire _w19211_ ;
	wire _w19210_ ;
	wire _w19209_ ;
	wire _w19208_ ;
	wire _w19207_ ;
	wire _w19206_ ;
	wire _w19205_ ;
	wire _w19204_ ;
	wire _w19203_ ;
	wire _w19202_ ;
	wire _w19201_ ;
	wire _w19200_ ;
	wire _w19199_ ;
	wire _w19198_ ;
	wire _w19197_ ;
	wire _w19196_ ;
	wire _w19195_ ;
	wire _w19194_ ;
	wire _w19193_ ;
	wire _w19192_ ;
	wire _w19191_ ;
	wire _w19190_ ;
	wire _w19189_ ;
	wire _w19188_ ;
	wire _w19187_ ;
	wire _w19186_ ;
	wire _w19185_ ;
	wire _w19184_ ;
	wire _w19183_ ;
	wire _w19182_ ;
	wire _w19181_ ;
	wire _w19180_ ;
	wire _w19179_ ;
	wire _w19178_ ;
	wire _w19177_ ;
	wire _w19176_ ;
	wire _w19175_ ;
	wire _w19174_ ;
	wire _w19173_ ;
	wire _w19172_ ;
	wire _w19171_ ;
	wire _w19170_ ;
	wire _w19169_ ;
	wire _w19168_ ;
	wire _w19167_ ;
	wire _w19166_ ;
	wire _w19165_ ;
	wire _w19164_ ;
	wire _w19163_ ;
	wire _w19162_ ;
	wire _w19161_ ;
	wire _w19160_ ;
	wire _w19159_ ;
	wire _w19158_ ;
	wire _w19157_ ;
	wire _w19156_ ;
	wire _w19155_ ;
	wire _w19154_ ;
	wire _w19153_ ;
	wire _w19152_ ;
	wire _w19151_ ;
	wire _w19150_ ;
	wire _w19149_ ;
	wire _w19148_ ;
	wire _w19147_ ;
	wire _w19146_ ;
	wire _w19145_ ;
	wire _w19144_ ;
	wire _w19143_ ;
	wire _w19142_ ;
	wire _w19141_ ;
	wire _w19140_ ;
	wire _w19139_ ;
	wire _w19138_ ;
	wire _w19137_ ;
	wire _w19136_ ;
	wire _w19135_ ;
	wire _w19134_ ;
	wire _w19133_ ;
	wire _w19132_ ;
	wire _w19131_ ;
	wire _w19130_ ;
	wire _w19129_ ;
	wire _w19128_ ;
	wire _w19127_ ;
	wire _w19126_ ;
	wire _w19125_ ;
	wire _w19124_ ;
	wire _w19123_ ;
	wire _w19122_ ;
	wire _w19121_ ;
	wire _w19120_ ;
	wire _w19119_ ;
	wire _w19118_ ;
	wire _w19117_ ;
	wire _w19116_ ;
	wire _w19115_ ;
	wire _w19114_ ;
	wire _w19113_ ;
	wire _w19112_ ;
	wire _w19111_ ;
	wire _w19110_ ;
	wire _w19109_ ;
	wire _w19108_ ;
	wire _w19107_ ;
	wire _w19106_ ;
	wire _w19105_ ;
	wire _w19104_ ;
	wire _w19103_ ;
	wire _w19102_ ;
	wire _w19101_ ;
	wire _w19100_ ;
	wire _w19099_ ;
	wire _w19098_ ;
	wire _w19097_ ;
	wire _w19096_ ;
	wire _w19095_ ;
	wire _w19094_ ;
	wire _w19093_ ;
	wire _w19092_ ;
	wire _w19091_ ;
	wire _w19090_ ;
	wire _w19089_ ;
	wire _w19088_ ;
	wire _w19087_ ;
	wire _w19086_ ;
	wire _w19085_ ;
	wire _w19084_ ;
	wire _w19083_ ;
	wire _w19082_ ;
	wire _w19081_ ;
	wire _w19080_ ;
	wire _w19079_ ;
	wire _w19078_ ;
	wire _w19077_ ;
	wire _w19076_ ;
	wire _w19075_ ;
	wire _w19074_ ;
	wire _w19073_ ;
	wire _w19072_ ;
	wire _w19071_ ;
	wire _w19070_ ;
	wire _w19069_ ;
	wire _w19068_ ;
	wire _w19067_ ;
	wire _w19066_ ;
	wire _w19065_ ;
	wire _w19064_ ;
	wire _w19063_ ;
	wire _w19062_ ;
	wire _w19061_ ;
	wire _w19060_ ;
	wire _w19059_ ;
	wire _w19058_ ;
	wire _w19057_ ;
	wire _w19056_ ;
	wire _w19055_ ;
	wire _w19054_ ;
	wire _w19053_ ;
	wire _w19052_ ;
	wire _w19051_ ;
	wire _w19050_ ;
	wire _w19049_ ;
	wire _w19048_ ;
	wire _w19047_ ;
	wire _w19046_ ;
	wire _w19045_ ;
	wire _w19044_ ;
	wire _w19043_ ;
	wire _w19042_ ;
	wire _w19041_ ;
	wire _w19040_ ;
	wire _w19039_ ;
	wire _w19038_ ;
	wire _w19037_ ;
	wire _w19036_ ;
	wire _w19035_ ;
	wire _w19034_ ;
	wire _w19033_ ;
	wire _w19032_ ;
	wire _w19031_ ;
	wire _w19030_ ;
	wire _w19029_ ;
	wire _w19028_ ;
	wire _w19027_ ;
	wire _w19026_ ;
	wire _w19025_ ;
	wire _w19024_ ;
	wire _w19023_ ;
	wire _w19022_ ;
	wire _w19021_ ;
	wire _w19020_ ;
	wire _w19019_ ;
	wire _w19018_ ;
	wire _w19017_ ;
	wire _w19016_ ;
	wire _w19015_ ;
	wire _w19014_ ;
	wire _w19013_ ;
	wire _w19012_ ;
	wire _w19011_ ;
	wire _w19010_ ;
	wire _w19009_ ;
	wire _w19008_ ;
	wire _w19007_ ;
	wire _w19006_ ;
	wire _w19005_ ;
	wire _w19004_ ;
	wire _w19003_ ;
	wire _w19002_ ;
	wire _w19001_ ;
	wire _w19000_ ;
	wire _w18999_ ;
	wire _w18998_ ;
	wire _w18997_ ;
	wire _w18996_ ;
	wire _w18995_ ;
	wire _w18994_ ;
	wire _w18993_ ;
	wire _w18992_ ;
	wire _w18991_ ;
	wire _w18990_ ;
	wire _w18989_ ;
	wire _w18988_ ;
	wire _w18987_ ;
	wire _w18986_ ;
	wire _w18985_ ;
	wire _w18984_ ;
	wire _w18983_ ;
	wire _w18982_ ;
	wire _w18981_ ;
	wire _w18980_ ;
	wire _w18979_ ;
	wire _w18978_ ;
	wire _w18977_ ;
	wire _w18976_ ;
	wire _w18975_ ;
	wire _w18974_ ;
	wire _w18973_ ;
	wire _w18972_ ;
	wire _w18971_ ;
	wire _w18970_ ;
	wire _w18969_ ;
	wire _w18968_ ;
	wire _w18967_ ;
	wire _w18966_ ;
	wire _w18965_ ;
	wire _w18964_ ;
	wire _w18963_ ;
	wire _w18962_ ;
	wire _w18961_ ;
	wire _w18960_ ;
	wire _w18959_ ;
	wire _w18958_ ;
	wire _w18957_ ;
	wire _w18956_ ;
	wire _w18955_ ;
	wire _w18954_ ;
	wire _w18953_ ;
	wire _w18952_ ;
	wire _w18951_ ;
	wire _w18950_ ;
	wire _w18949_ ;
	wire _w18948_ ;
	wire _w18947_ ;
	wire _w18946_ ;
	wire _w18945_ ;
	wire _w18944_ ;
	wire _w18943_ ;
	wire _w18942_ ;
	wire _w18941_ ;
	wire _w18940_ ;
	wire _w18939_ ;
	wire _w18938_ ;
	wire _w18937_ ;
	wire _w18936_ ;
	wire _w18935_ ;
	wire _w18934_ ;
	wire _w18933_ ;
	wire _w18932_ ;
	wire _w18931_ ;
	wire _w18930_ ;
	wire _w18929_ ;
	wire _w18928_ ;
	wire _w18927_ ;
	wire _w18926_ ;
	wire _w18925_ ;
	wire _w18924_ ;
	wire _w18923_ ;
	wire _w18922_ ;
	wire _w18921_ ;
	wire _w18920_ ;
	wire _w18919_ ;
	wire _w18918_ ;
	wire _w18917_ ;
	wire _w18916_ ;
	wire _w18915_ ;
	wire _w18914_ ;
	wire _w18913_ ;
	wire _w18912_ ;
	wire _w18911_ ;
	wire _w18910_ ;
	wire _w18909_ ;
	wire _w18908_ ;
	wire _w18907_ ;
	wire _w18906_ ;
	wire _w18905_ ;
	wire _w18904_ ;
	wire _w18903_ ;
	wire _w18902_ ;
	wire _w18901_ ;
	wire _w18900_ ;
	wire _w18899_ ;
	wire _w18898_ ;
	wire _w18897_ ;
	wire _w18896_ ;
	wire _w18895_ ;
	wire _w18894_ ;
	wire _w18893_ ;
	wire _w18892_ ;
	wire _w18891_ ;
	wire _w18890_ ;
	wire _w18889_ ;
	wire _w18888_ ;
	wire _w18887_ ;
	wire _w18886_ ;
	wire _w18885_ ;
	wire _w18884_ ;
	wire _w18883_ ;
	wire _w18882_ ;
	wire _w18881_ ;
	wire _w18880_ ;
	wire _w18879_ ;
	wire _w18878_ ;
	wire _w18877_ ;
	wire _w18876_ ;
	wire _w18875_ ;
	wire _w18874_ ;
	wire _w18873_ ;
	wire _w18872_ ;
	wire _w18871_ ;
	wire _w18870_ ;
	wire _w18869_ ;
	wire _w18868_ ;
	wire _w18867_ ;
	wire _w18866_ ;
	wire _w18865_ ;
	wire _w18864_ ;
	wire _w18863_ ;
	wire _w18862_ ;
	wire _w18861_ ;
	wire _w18860_ ;
	wire _w18859_ ;
	wire _w18858_ ;
	wire _w18857_ ;
	wire _w18856_ ;
	wire _w18855_ ;
	wire _w18854_ ;
	wire _w18853_ ;
	wire _w18852_ ;
	wire _w18851_ ;
	wire _w18850_ ;
	wire _w18849_ ;
	wire _w18848_ ;
	wire _w18847_ ;
	wire _w18846_ ;
	wire _w18845_ ;
	wire _w18844_ ;
	wire _w18843_ ;
	wire _w18842_ ;
	wire _w18841_ ;
	wire _w18840_ ;
	wire _w18839_ ;
	wire _w18838_ ;
	wire _w18837_ ;
	wire _w18836_ ;
	wire _w18835_ ;
	wire _w18834_ ;
	wire _w18833_ ;
	wire _w18832_ ;
	wire _w18831_ ;
	wire _w18830_ ;
	wire _w18829_ ;
	wire _w18828_ ;
	wire _w18827_ ;
	wire _w18826_ ;
	wire _w18825_ ;
	wire _w18824_ ;
	wire _w18823_ ;
	wire _w18822_ ;
	wire _w18821_ ;
	wire _w18820_ ;
	wire _w18819_ ;
	wire _w18818_ ;
	wire _w18817_ ;
	wire _w18816_ ;
	wire _w18815_ ;
	wire _w18814_ ;
	wire _w18813_ ;
	wire _w18812_ ;
	wire _w18811_ ;
	wire _w18810_ ;
	wire _w18809_ ;
	wire _w18808_ ;
	wire _w18807_ ;
	wire _w18806_ ;
	wire _w18805_ ;
	wire _w18804_ ;
	wire _w18803_ ;
	wire _w18802_ ;
	wire _w18801_ ;
	wire _w18800_ ;
	wire _w18799_ ;
	wire _w18798_ ;
	wire _w18797_ ;
	wire _w18796_ ;
	wire _w18795_ ;
	wire _w18794_ ;
	wire _w18793_ ;
	wire _w18792_ ;
	wire _w18791_ ;
	wire _w18790_ ;
	wire _w18789_ ;
	wire _w18788_ ;
	wire _w18787_ ;
	wire _w18786_ ;
	wire _w18785_ ;
	wire _w18784_ ;
	wire _w18783_ ;
	wire _w18782_ ;
	wire _w18781_ ;
	wire _w18780_ ;
	wire _w18779_ ;
	wire _w18778_ ;
	wire _w18777_ ;
	wire _w18776_ ;
	wire _w18775_ ;
	wire _w18774_ ;
	wire _w18773_ ;
	wire _w18772_ ;
	wire _w18771_ ;
	wire _w18770_ ;
	wire _w18769_ ;
	wire _w18768_ ;
	wire _w18767_ ;
	wire _w18766_ ;
	wire _w18765_ ;
	wire _w18764_ ;
	wire _w18763_ ;
	wire _w18762_ ;
	wire _w18761_ ;
	wire _w18760_ ;
	wire _w18759_ ;
	wire _w18758_ ;
	wire _w18757_ ;
	wire _w18756_ ;
	wire _w18755_ ;
	wire _w18754_ ;
	wire _w18753_ ;
	wire _w18752_ ;
	wire _w18751_ ;
	wire _w18750_ ;
	wire _w18749_ ;
	wire _w18748_ ;
	wire _w18747_ ;
	wire _w18746_ ;
	wire _w18745_ ;
	wire _w18744_ ;
	wire _w18743_ ;
	wire _w18742_ ;
	wire _w18741_ ;
	wire _w18740_ ;
	wire _w18739_ ;
	wire _w18738_ ;
	wire _w18737_ ;
	wire _w18736_ ;
	wire _w18735_ ;
	wire _w18734_ ;
	wire _w18733_ ;
	wire _w18732_ ;
	wire _w18731_ ;
	wire _w18730_ ;
	wire _w18729_ ;
	wire _w18728_ ;
	wire _w18727_ ;
	wire _w18726_ ;
	wire _w18725_ ;
	wire _w18724_ ;
	wire _w18723_ ;
	wire _w18722_ ;
	wire _w18721_ ;
	wire _w18720_ ;
	wire _w18719_ ;
	wire _w18718_ ;
	wire _w18717_ ;
	wire _w18716_ ;
	wire _w18715_ ;
	wire _w18714_ ;
	wire _w18713_ ;
	wire _w18712_ ;
	wire _w18711_ ;
	wire _w18710_ ;
	wire _w18709_ ;
	wire _w18708_ ;
	wire _w18707_ ;
	wire _w18706_ ;
	wire _w18705_ ;
	wire _w18704_ ;
	wire _w18703_ ;
	wire _w18702_ ;
	wire _w18701_ ;
	wire _w18700_ ;
	wire _w18699_ ;
	wire _w18698_ ;
	wire _w18697_ ;
	wire _w18696_ ;
	wire _w18695_ ;
	wire _w18694_ ;
	wire _w18693_ ;
	wire _w18692_ ;
	wire _w18691_ ;
	wire _w18690_ ;
	wire _w18689_ ;
	wire _w18688_ ;
	wire _w18687_ ;
	wire _w18686_ ;
	wire _w18685_ ;
	wire _w18684_ ;
	wire _w18683_ ;
	wire _w18682_ ;
	wire _w18681_ ;
	wire _w18680_ ;
	wire _w18679_ ;
	wire _w18678_ ;
	wire _w18677_ ;
	wire _w18676_ ;
	wire _w18675_ ;
	wire _w18674_ ;
	wire _w18673_ ;
	wire _w18672_ ;
	wire _w18671_ ;
	wire _w18670_ ;
	wire _w18669_ ;
	wire _w18668_ ;
	wire _w18667_ ;
	wire _w18666_ ;
	wire _w18665_ ;
	wire _w18664_ ;
	wire _w18663_ ;
	wire _w18662_ ;
	wire _w18661_ ;
	wire _w18660_ ;
	wire _w18659_ ;
	wire _w18658_ ;
	wire _w18657_ ;
	wire _w18656_ ;
	wire _w18655_ ;
	wire _w18654_ ;
	wire _w18653_ ;
	wire _w18652_ ;
	wire _w18651_ ;
	wire _w18650_ ;
	wire _w18649_ ;
	wire _w18648_ ;
	wire _w18647_ ;
	wire _w18646_ ;
	wire _w18645_ ;
	wire _w18644_ ;
	wire _w18643_ ;
	wire _w18642_ ;
	wire _w18641_ ;
	wire _w18640_ ;
	wire _w18639_ ;
	wire _w18638_ ;
	wire _w18637_ ;
	wire _w18636_ ;
	wire _w18635_ ;
	wire _w18634_ ;
	wire _w18633_ ;
	wire _w18632_ ;
	wire _w18631_ ;
	wire _w18630_ ;
	wire _w18629_ ;
	wire _w18628_ ;
	wire _w18627_ ;
	wire _w18626_ ;
	wire _w18625_ ;
	wire _w18624_ ;
	wire _w18623_ ;
	wire _w18622_ ;
	wire _w18621_ ;
	wire _w18620_ ;
	wire _w18619_ ;
	wire _w18618_ ;
	wire _w18617_ ;
	wire _w18616_ ;
	wire _w18615_ ;
	wire _w18614_ ;
	wire _w18613_ ;
	wire _w18612_ ;
	wire _w18611_ ;
	wire _w18610_ ;
	wire _w18609_ ;
	wire _w18608_ ;
	wire _w18607_ ;
	wire _w18606_ ;
	wire _w18605_ ;
	wire _w18604_ ;
	wire _w18603_ ;
	wire _w18602_ ;
	wire _w18601_ ;
	wire _w18600_ ;
	wire _w18599_ ;
	wire _w18598_ ;
	wire _w18597_ ;
	wire _w18596_ ;
	wire _w18595_ ;
	wire _w18594_ ;
	wire _w18593_ ;
	wire _w18592_ ;
	wire _w18591_ ;
	wire _w18590_ ;
	wire _w18589_ ;
	wire _w18588_ ;
	wire _w18587_ ;
	wire _w18586_ ;
	wire _w18585_ ;
	wire _w18584_ ;
	wire _w18583_ ;
	wire _w18582_ ;
	wire _w18581_ ;
	wire _w18580_ ;
	wire _w18579_ ;
	wire _w18578_ ;
	wire _w18577_ ;
	wire _w18576_ ;
	wire _w18575_ ;
	wire _w18574_ ;
	wire _w18573_ ;
	wire _w18572_ ;
	wire _w18571_ ;
	wire _w18570_ ;
	wire _w18569_ ;
	wire _w18568_ ;
	wire _w18567_ ;
	wire _w18566_ ;
	wire _w18565_ ;
	wire _w18564_ ;
	wire _w18563_ ;
	wire _w18562_ ;
	wire _w18561_ ;
	wire _w18560_ ;
	wire _w18559_ ;
	wire _w18558_ ;
	wire _w18557_ ;
	wire _w18556_ ;
	wire _w18555_ ;
	wire _w18554_ ;
	wire _w18553_ ;
	wire _w18552_ ;
	wire _w18551_ ;
	wire _w18550_ ;
	wire _w18549_ ;
	wire _w18548_ ;
	wire _w18547_ ;
	wire _w18546_ ;
	wire _w18545_ ;
	wire _w18544_ ;
	wire _w18543_ ;
	wire _w18542_ ;
	wire _w18541_ ;
	wire _w18540_ ;
	wire _w18539_ ;
	wire _w18538_ ;
	wire _w18537_ ;
	wire _w18536_ ;
	wire _w18535_ ;
	wire _w18534_ ;
	wire _w18533_ ;
	wire _w18532_ ;
	wire _w18531_ ;
	wire _w18530_ ;
	wire _w18529_ ;
	wire _w18528_ ;
	wire _w18527_ ;
	wire _w18526_ ;
	wire _w18525_ ;
	wire _w18524_ ;
	wire _w18523_ ;
	wire _w18522_ ;
	wire _w18521_ ;
	wire _w18520_ ;
	wire _w18519_ ;
	wire _w18518_ ;
	wire _w18517_ ;
	wire _w18516_ ;
	wire _w18515_ ;
	wire _w18514_ ;
	wire _w18513_ ;
	wire _w18512_ ;
	wire _w18511_ ;
	wire _w18510_ ;
	wire _w18509_ ;
	wire _w18508_ ;
	wire _w18507_ ;
	wire _w18506_ ;
	wire _w18505_ ;
	wire _w18504_ ;
	wire _w18503_ ;
	wire _w18502_ ;
	wire _w18501_ ;
	wire _w18500_ ;
	wire _w18499_ ;
	wire _w18498_ ;
	wire _w18497_ ;
	wire _w18496_ ;
	wire _w18495_ ;
	wire _w18494_ ;
	wire _w18493_ ;
	wire _w18492_ ;
	wire _w18491_ ;
	wire _w18490_ ;
	wire _w18489_ ;
	wire _w18488_ ;
	wire _w18487_ ;
	wire _w18486_ ;
	wire _w18485_ ;
	wire _w18484_ ;
	wire _w18483_ ;
	wire _w18482_ ;
	wire _w18481_ ;
	wire _w18480_ ;
	wire _w18479_ ;
	wire _w18478_ ;
	wire _w18477_ ;
	wire _w18476_ ;
	wire _w18475_ ;
	wire _w18474_ ;
	wire _w18473_ ;
	wire _w18472_ ;
	wire _w18471_ ;
	wire _w18470_ ;
	wire _w18469_ ;
	wire _w18468_ ;
	wire _w18467_ ;
	wire _w18466_ ;
	wire _w18465_ ;
	wire _w18464_ ;
	wire _w18463_ ;
	wire _w18462_ ;
	wire _w18461_ ;
	wire _w18460_ ;
	wire _w18459_ ;
	wire _w18458_ ;
	wire _w18457_ ;
	wire _w18456_ ;
	wire _w18455_ ;
	wire _w18454_ ;
	wire _w18453_ ;
	wire _w18452_ ;
	wire _w18451_ ;
	wire _w18450_ ;
	wire _w18449_ ;
	wire _w18448_ ;
	wire _w18447_ ;
	wire _w18446_ ;
	wire _w18445_ ;
	wire _w18444_ ;
	wire _w18443_ ;
	wire _w18442_ ;
	wire _w18441_ ;
	wire _w18440_ ;
	wire _w18439_ ;
	wire _w18438_ ;
	wire _w18437_ ;
	wire _w18436_ ;
	wire _w18435_ ;
	wire _w18434_ ;
	wire _w18433_ ;
	wire _w18432_ ;
	wire _w18431_ ;
	wire _w18430_ ;
	wire _w18429_ ;
	wire _w18428_ ;
	wire _w18427_ ;
	wire _w18426_ ;
	wire _w18425_ ;
	wire _w18424_ ;
	wire _w18423_ ;
	wire _w18422_ ;
	wire _w18421_ ;
	wire _w18420_ ;
	wire _w18419_ ;
	wire _w18418_ ;
	wire _w18417_ ;
	wire _w18416_ ;
	wire _w18415_ ;
	wire _w18414_ ;
	wire _w18413_ ;
	wire _w18412_ ;
	wire _w18411_ ;
	wire _w18410_ ;
	wire _w18409_ ;
	wire _w18408_ ;
	wire _w18407_ ;
	wire _w18406_ ;
	wire _w18405_ ;
	wire _w18404_ ;
	wire _w18403_ ;
	wire _w18402_ ;
	wire _w18401_ ;
	wire _w18400_ ;
	wire _w18399_ ;
	wire _w18398_ ;
	wire _w18397_ ;
	wire _w18396_ ;
	wire _w18395_ ;
	wire _w18394_ ;
	wire _w18393_ ;
	wire _w18392_ ;
	wire _w18391_ ;
	wire _w18390_ ;
	wire _w18389_ ;
	wire _w18388_ ;
	wire _w18387_ ;
	wire _w18386_ ;
	wire _w18385_ ;
	wire _w18384_ ;
	wire _w18383_ ;
	wire _w18382_ ;
	wire _w18381_ ;
	wire _w18380_ ;
	wire _w18379_ ;
	wire _w18378_ ;
	wire _w18377_ ;
	wire _w18376_ ;
	wire _w18375_ ;
	wire _w18374_ ;
	wire _w18373_ ;
	wire _w18372_ ;
	wire _w18371_ ;
	wire _w18370_ ;
	wire _w18369_ ;
	wire _w18368_ ;
	wire _w18367_ ;
	wire _w18366_ ;
	wire _w18365_ ;
	wire _w18364_ ;
	wire _w18363_ ;
	wire _w18362_ ;
	wire _w18361_ ;
	wire _w18360_ ;
	wire _w18359_ ;
	wire _w18358_ ;
	wire _w18357_ ;
	wire _w18356_ ;
	wire _w18355_ ;
	wire _w18354_ ;
	wire _w18353_ ;
	wire _w18352_ ;
	wire _w18351_ ;
	wire _w18350_ ;
	wire _w18349_ ;
	wire _w18348_ ;
	wire _w18347_ ;
	wire _w18346_ ;
	wire _w18345_ ;
	wire _w18344_ ;
	wire _w18343_ ;
	wire _w18342_ ;
	wire _w18341_ ;
	wire _w18340_ ;
	wire _w18339_ ;
	wire _w18338_ ;
	wire _w18337_ ;
	wire _w18336_ ;
	wire _w18335_ ;
	wire _w18334_ ;
	wire _w18333_ ;
	wire _w18332_ ;
	wire _w18331_ ;
	wire _w18330_ ;
	wire _w18329_ ;
	wire _w18328_ ;
	wire _w18327_ ;
	wire _w18326_ ;
	wire _w18325_ ;
	wire _w18324_ ;
	wire _w18323_ ;
	wire _w18322_ ;
	wire _w18321_ ;
	wire _w18320_ ;
	wire _w18319_ ;
	wire _w18318_ ;
	wire _w18317_ ;
	wire _w18316_ ;
	wire _w18315_ ;
	wire _w18314_ ;
	wire _w18313_ ;
	wire _w18312_ ;
	wire _w18311_ ;
	wire _w18310_ ;
	wire _w18309_ ;
	wire _w18308_ ;
	wire _w18307_ ;
	wire _w18306_ ;
	wire _w18305_ ;
	wire _w18304_ ;
	wire _w18303_ ;
	wire _w18302_ ;
	wire _w18301_ ;
	wire _w18300_ ;
	wire _w18299_ ;
	wire _w18298_ ;
	wire _w18297_ ;
	wire _w18296_ ;
	wire _w18295_ ;
	wire _w18294_ ;
	wire _w18293_ ;
	wire _w18292_ ;
	wire _w18291_ ;
	wire _w18290_ ;
	wire _w18289_ ;
	wire _w18288_ ;
	wire _w18287_ ;
	wire _w18286_ ;
	wire _w18285_ ;
	wire _w18284_ ;
	wire _w18283_ ;
	wire _w18282_ ;
	wire _w18281_ ;
	wire _w18280_ ;
	wire _w18279_ ;
	wire _w18278_ ;
	wire _w18277_ ;
	wire _w18276_ ;
	wire _w18275_ ;
	wire _w18274_ ;
	wire _w18273_ ;
	wire _w18272_ ;
	wire _w18271_ ;
	wire _w18270_ ;
	wire _w18269_ ;
	wire _w18268_ ;
	wire _w18267_ ;
	wire _w18266_ ;
	wire _w18265_ ;
	wire _w18264_ ;
	wire _w18263_ ;
	wire _w18262_ ;
	wire _w18261_ ;
	wire _w18260_ ;
	wire _w18259_ ;
	wire _w18258_ ;
	wire _w18257_ ;
	wire _w18256_ ;
	wire _w18255_ ;
	wire _w18254_ ;
	wire _w18253_ ;
	wire _w18252_ ;
	wire _w18251_ ;
	wire _w18250_ ;
	wire _w18249_ ;
	wire _w18248_ ;
	wire _w18247_ ;
	wire _w18246_ ;
	wire _w18245_ ;
	wire _w18244_ ;
	wire _w18243_ ;
	wire _w18242_ ;
	wire _w18241_ ;
	wire _w18240_ ;
	wire _w18239_ ;
	wire _w18238_ ;
	wire _w18237_ ;
	wire _w18236_ ;
	wire _w18235_ ;
	wire _w18234_ ;
	wire _w18233_ ;
	wire _w18232_ ;
	wire _w18231_ ;
	wire _w18230_ ;
	wire _w18229_ ;
	wire _w18228_ ;
	wire _w18227_ ;
	wire _w18226_ ;
	wire _w18225_ ;
	wire _w18224_ ;
	wire _w18223_ ;
	wire _w18222_ ;
	wire _w18221_ ;
	wire _w18220_ ;
	wire _w18219_ ;
	wire _w18218_ ;
	wire _w18217_ ;
	wire _w18216_ ;
	wire _w18215_ ;
	wire _w18214_ ;
	wire _w18213_ ;
	wire _w18212_ ;
	wire _w18211_ ;
	wire _w18210_ ;
	wire _w18209_ ;
	wire _w18208_ ;
	wire _w18207_ ;
	wire _w18206_ ;
	wire _w18205_ ;
	wire _w18204_ ;
	wire _w18203_ ;
	wire _w18202_ ;
	wire _w18201_ ;
	wire _w18200_ ;
	wire _w18199_ ;
	wire _w18198_ ;
	wire _w18197_ ;
	wire _w18196_ ;
	wire _w18195_ ;
	wire _w18194_ ;
	wire _w18193_ ;
	wire _w18192_ ;
	wire _w18191_ ;
	wire _w18190_ ;
	wire _w18189_ ;
	wire _w18188_ ;
	wire _w18187_ ;
	wire _w18186_ ;
	wire _w18185_ ;
	wire _w18184_ ;
	wire _w18183_ ;
	wire _w18182_ ;
	wire _w18181_ ;
	wire _w18180_ ;
	wire _w18179_ ;
	wire _w18178_ ;
	wire _w18177_ ;
	wire _w18176_ ;
	wire _w18175_ ;
	wire _w18174_ ;
	wire _w18173_ ;
	wire _w18172_ ;
	wire _w18171_ ;
	wire _w18170_ ;
	wire _w18169_ ;
	wire _w18168_ ;
	wire _w18167_ ;
	wire _w18166_ ;
	wire _w18165_ ;
	wire _w18164_ ;
	wire _w18163_ ;
	wire _w18162_ ;
	wire _w18161_ ;
	wire _w18160_ ;
	wire _w18159_ ;
	wire _w18158_ ;
	wire _w18157_ ;
	wire _w18156_ ;
	wire _w18155_ ;
	wire _w18154_ ;
	wire _w18153_ ;
	wire _w18152_ ;
	wire _w18151_ ;
	wire _w18150_ ;
	wire _w18149_ ;
	wire _w18148_ ;
	wire _w18147_ ;
	wire _w18146_ ;
	wire _w18145_ ;
	wire _w18144_ ;
	wire _w18143_ ;
	wire _w18142_ ;
	wire _w18141_ ;
	wire _w18140_ ;
	wire _w18139_ ;
	wire _w18138_ ;
	wire _w18137_ ;
	wire _w18136_ ;
	wire _w18135_ ;
	wire _w18134_ ;
	wire _w18133_ ;
	wire _w18132_ ;
	wire _w18131_ ;
	wire _w18130_ ;
	wire _w18129_ ;
	wire _w18128_ ;
	wire _w18127_ ;
	wire _w18126_ ;
	wire _w18125_ ;
	wire _w18124_ ;
	wire _w18123_ ;
	wire _w18122_ ;
	wire _w18121_ ;
	wire _w18120_ ;
	wire _w18119_ ;
	wire _w18118_ ;
	wire _w18117_ ;
	wire _w18116_ ;
	wire _w18115_ ;
	wire _w18114_ ;
	wire _w18113_ ;
	wire _w18112_ ;
	wire _w18111_ ;
	wire _w18110_ ;
	wire _w18109_ ;
	wire _w18108_ ;
	wire _w18107_ ;
	wire _w18106_ ;
	wire _w18105_ ;
	wire _w18104_ ;
	wire _w18103_ ;
	wire _w18102_ ;
	wire _w18101_ ;
	wire _w18100_ ;
	wire _w18099_ ;
	wire _w18098_ ;
	wire _w18097_ ;
	wire _w18096_ ;
	wire _w18095_ ;
	wire _w18094_ ;
	wire _w18093_ ;
	wire _w18092_ ;
	wire _w18091_ ;
	wire _w18090_ ;
	wire _w18089_ ;
	wire _w18088_ ;
	wire _w18087_ ;
	wire _w18086_ ;
	wire _w18085_ ;
	wire _w18084_ ;
	wire _w18083_ ;
	wire _w18082_ ;
	wire _w18081_ ;
	wire _w18080_ ;
	wire _w18079_ ;
	wire _w18078_ ;
	wire _w18077_ ;
	wire _w18076_ ;
	wire _w18075_ ;
	wire _w18074_ ;
	wire _w18073_ ;
	wire _w18072_ ;
	wire _w18071_ ;
	wire _w18070_ ;
	wire _w18069_ ;
	wire _w18068_ ;
	wire _w18067_ ;
	wire _w18066_ ;
	wire _w18065_ ;
	wire _w18064_ ;
	wire _w18063_ ;
	wire _w18062_ ;
	wire _w18061_ ;
	wire _w18060_ ;
	wire _w18059_ ;
	wire _w18058_ ;
	wire _w18057_ ;
	wire _w18056_ ;
	wire _w18055_ ;
	wire _w18054_ ;
	wire _w18053_ ;
	wire _w18052_ ;
	wire _w18051_ ;
	wire _w18050_ ;
	wire _w18049_ ;
	wire _w18048_ ;
	wire _w18047_ ;
	wire _w18046_ ;
	wire _w18045_ ;
	wire _w18044_ ;
	wire _w18043_ ;
	wire _w18042_ ;
	wire _w18041_ ;
	wire _w18040_ ;
	wire _w18039_ ;
	wire _w18038_ ;
	wire _w18037_ ;
	wire _w18036_ ;
	wire _w18035_ ;
	wire _w18034_ ;
	wire _w18033_ ;
	wire _w18032_ ;
	wire _w18031_ ;
	wire _w18030_ ;
	wire _w18029_ ;
	wire _w18028_ ;
	wire _w18027_ ;
	wire _w18026_ ;
	wire _w18025_ ;
	wire _w18024_ ;
	wire _w18023_ ;
	wire _w18022_ ;
	wire _w18021_ ;
	wire _w18020_ ;
	wire _w18019_ ;
	wire _w18018_ ;
	wire _w18017_ ;
	wire _w18016_ ;
	wire _w18015_ ;
	wire _w18014_ ;
	wire _w18013_ ;
	wire _w18012_ ;
	wire _w18011_ ;
	wire _w18010_ ;
	wire _w18009_ ;
	wire _w18008_ ;
	wire _w18007_ ;
	wire _w18006_ ;
	wire _w18005_ ;
	wire _w18004_ ;
	wire _w18003_ ;
	wire _w18002_ ;
	wire _w18001_ ;
	wire _w18000_ ;
	wire _w17999_ ;
	wire _w17998_ ;
	wire _w17997_ ;
	wire _w17996_ ;
	wire _w17995_ ;
	wire _w17994_ ;
	wire _w17993_ ;
	wire _w17992_ ;
	wire _w17991_ ;
	wire _w17990_ ;
	wire _w17989_ ;
	wire _w17988_ ;
	wire _w17987_ ;
	wire _w17986_ ;
	wire _w17985_ ;
	wire _w17984_ ;
	wire _w17983_ ;
	wire _w17982_ ;
	wire _w17981_ ;
	wire _w17980_ ;
	wire _w17979_ ;
	wire _w17978_ ;
	wire _w17977_ ;
	wire _w17976_ ;
	wire _w17975_ ;
	wire _w17974_ ;
	wire _w17973_ ;
	wire _w17972_ ;
	wire _w17971_ ;
	wire _w17970_ ;
	wire _w17969_ ;
	wire _w17968_ ;
	wire _w17967_ ;
	wire _w17966_ ;
	wire _w17965_ ;
	wire _w17964_ ;
	wire _w17963_ ;
	wire _w17962_ ;
	wire _w17961_ ;
	wire _w17960_ ;
	wire _w17959_ ;
	wire _w17958_ ;
	wire _w17957_ ;
	wire _w17956_ ;
	wire _w17955_ ;
	wire _w17954_ ;
	wire _w17953_ ;
	wire _w17952_ ;
	wire _w17951_ ;
	wire _w17950_ ;
	wire _w17949_ ;
	wire _w17948_ ;
	wire _w17947_ ;
	wire _w17946_ ;
	wire _w17945_ ;
	wire _w17944_ ;
	wire _w17943_ ;
	wire _w17942_ ;
	wire _w17941_ ;
	wire _w17940_ ;
	wire _w17939_ ;
	wire _w17938_ ;
	wire _w17937_ ;
	wire _w17936_ ;
	wire _w17935_ ;
	wire _w17934_ ;
	wire _w17933_ ;
	wire _w17932_ ;
	wire _w17931_ ;
	wire _w17930_ ;
	wire _w17929_ ;
	wire _w17928_ ;
	wire _w17927_ ;
	wire _w17926_ ;
	wire _w17925_ ;
	wire _w17924_ ;
	wire _w17923_ ;
	wire _w17922_ ;
	wire _w17921_ ;
	wire _w17920_ ;
	wire _w17919_ ;
	wire _w17918_ ;
	wire _w17917_ ;
	wire _w17916_ ;
	wire _w17915_ ;
	wire _w17914_ ;
	wire _w17913_ ;
	wire _w17912_ ;
	wire _w17911_ ;
	wire _w17910_ ;
	wire _w17909_ ;
	wire _w17908_ ;
	wire _w17907_ ;
	wire _w17906_ ;
	wire _w17905_ ;
	wire _w17904_ ;
	wire _w17903_ ;
	wire _w17902_ ;
	wire _w17901_ ;
	wire _w17900_ ;
	wire _w17899_ ;
	wire _w17898_ ;
	wire _w17897_ ;
	wire _w17896_ ;
	wire _w17895_ ;
	wire _w17894_ ;
	wire _w17893_ ;
	wire _w17892_ ;
	wire _w17891_ ;
	wire _w17890_ ;
	wire _w17889_ ;
	wire _w17888_ ;
	wire _w17887_ ;
	wire _w17886_ ;
	wire _w17885_ ;
	wire _w17884_ ;
	wire _w17883_ ;
	wire _w17882_ ;
	wire _w17881_ ;
	wire _w17880_ ;
	wire _w17879_ ;
	wire _w17878_ ;
	wire _w17877_ ;
	wire _w17876_ ;
	wire _w17875_ ;
	wire _w17874_ ;
	wire _w17873_ ;
	wire _w17872_ ;
	wire _w17871_ ;
	wire _w17870_ ;
	wire _w17869_ ;
	wire _w17868_ ;
	wire _w17867_ ;
	wire _w17866_ ;
	wire _w17865_ ;
	wire _w17864_ ;
	wire _w17863_ ;
	wire _w17862_ ;
	wire _w17861_ ;
	wire _w17860_ ;
	wire _w17859_ ;
	wire _w17858_ ;
	wire _w17857_ ;
	wire _w17856_ ;
	wire _w17855_ ;
	wire _w17854_ ;
	wire _w17853_ ;
	wire _w17852_ ;
	wire _w17851_ ;
	wire _w17850_ ;
	wire _w17849_ ;
	wire _w17848_ ;
	wire _w17847_ ;
	wire _w17846_ ;
	wire _w17845_ ;
	wire _w17844_ ;
	wire _w17843_ ;
	wire _w17842_ ;
	wire _w17841_ ;
	wire _w17840_ ;
	wire _w17839_ ;
	wire _w17838_ ;
	wire _w17837_ ;
	wire _w17836_ ;
	wire _w17835_ ;
	wire _w17834_ ;
	wire _w17833_ ;
	wire _w17832_ ;
	wire _w17831_ ;
	wire _w17830_ ;
	wire _w17829_ ;
	wire _w17828_ ;
	wire _w17827_ ;
	wire _w17826_ ;
	wire _w17825_ ;
	wire _w17824_ ;
	wire _w17823_ ;
	wire _w17822_ ;
	wire _w17821_ ;
	wire _w17820_ ;
	wire _w17819_ ;
	wire _w17818_ ;
	wire _w17817_ ;
	wire _w17816_ ;
	wire _w17815_ ;
	wire _w17814_ ;
	wire _w17813_ ;
	wire _w17812_ ;
	wire _w17811_ ;
	wire _w17810_ ;
	wire _w17809_ ;
	wire _w17808_ ;
	wire _w17807_ ;
	wire _w17806_ ;
	wire _w17805_ ;
	wire _w17804_ ;
	wire _w17803_ ;
	wire _w17802_ ;
	wire _w17801_ ;
	wire _w17800_ ;
	wire _w17799_ ;
	wire _w17798_ ;
	wire _w17797_ ;
	wire _w17796_ ;
	wire _w17795_ ;
	wire _w17794_ ;
	wire _w17793_ ;
	wire _w17792_ ;
	wire _w17791_ ;
	wire _w17790_ ;
	wire _w17789_ ;
	wire _w17788_ ;
	wire _w17787_ ;
	wire _w17786_ ;
	wire _w17785_ ;
	wire _w17784_ ;
	wire _w17783_ ;
	wire _w17782_ ;
	wire _w17781_ ;
	wire _w17780_ ;
	wire _w17779_ ;
	wire _w17778_ ;
	wire _w17777_ ;
	wire _w17776_ ;
	wire _w17775_ ;
	wire _w17774_ ;
	wire _w17773_ ;
	wire _w17772_ ;
	wire _w17771_ ;
	wire _w17770_ ;
	wire _w17769_ ;
	wire _w17768_ ;
	wire _w17767_ ;
	wire _w17766_ ;
	wire _w17765_ ;
	wire _w17764_ ;
	wire _w17763_ ;
	wire _w17762_ ;
	wire _w17761_ ;
	wire _w17760_ ;
	wire _w17759_ ;
	wire _w17758_ ;
	wire _w17757_ ;
	wire _w17756_ ;
	wire _w17755_ ;
	wire _w17754_ ;
	wire _w17753_ ;
	wire _w17752_ ;
	wire _w17751_ ;
	wire _w17750_ ;
	wire _w17749_ ;
	wire _w17748_ ;
	wire _w17747_ ;
	wire _w17746_ ;
	wire _w17745_ ;
	wire _w17744_ ;
	wire _w17743_ ;
	wire _w17742_ ;
	wire _w17741_ ;
	wire _w17740_ ;
	wire _w17739_ ;
	wire _w17738_ ;
	wire _w17737_ ;
	wire _w17736_ ;
	wire _w17735_ ;
	wire _w17734_ ;
	wire _w17733_ ;
	wire _w17732_ ;
	wire _w17731_ ;
	wire _w17730_ ;
	wire _w17729_ ;
	wire _w17728_ ;
	wire _w17727_ ;
	wire _w17726_ ;
	wire _w17725_ ;
	wire _w17724_ ;
	wire _w17723_ ;
	wire _w17722_ ;
	wire _w17721_ ;
	wire _w17720_ ;
	wire _w17719_ ;
	wire _w17718_ ;
	wire _w17717_ ;
	wire _w17716_ ;
	wire _w17715_ ;
	wire _w17714_ ;
	wire _w17713_ ;
	wire _w17712_ ;
	wire _w17711_ ;
	wire _w17710_ ;
	wire _w17709_ ;
	wire _w17708_ ;
	wire _w17707_ ;
	wire _w17706_ ;
	wire _w17705_ ;
	wire _w17704_ ;
	wire _w17703_ ;
	wire _w17702_ ;
	wire _w17701_ ;
	wire _w17700_ ;
	wire _w17699_ ;
	wire _w17698_ ;
	wire _w17697_ ;
	wire _w17696_ ;
	wire _w17695_ ;
	wire _w17694_ ;
	wire _w17693_ ;
	wire _w17692_ ;
	wire _w17691_ ;
	wire _w17690_ ;
	wire _w17689_ ;
	wire _w17688_ ;
	wire _w17687_ ;
	wire _w17686_ ;
	wire _w17685_ ;
	wire _w17684_ ;
	wire _w17683_ ;
	wire _w17682_ ;
	wire _w17681_ ;
	wire _w17680_ ;
	wire _w17679_ ;
	wire _w17678_ ;
	wire _w17677_ ;
	wire _w17676_ ;
	wire _w17675_ ;
	wire _w17674_ ;
	wire _w17673_ ;
	wire _w17672_ ;
	wire _w17671_ ;
	wire _w17670_ ;
	wire _w17669_ ;
	wire _w17668_ ;
	wire _w17667_ ;
	wire _w17666_ ;
	wire _w17665_ ;
	wire _w17664_ ;
	wire _w17663_ ;
	wire _w17662_ ;
	wire _w17661_ ;
	wire _w17660_ ;
	wire _w17659_ ;
	wire _w17658_ ;
	wire _w17657_ ;
	wire _w17656_ ;
	wire _w17655_ ;
	wire _w17654_ ;
	wire _w17653_ ;
	wire _w17652_ ;
	wire _w17651_ ;
	wire _w17650_ ;
	wire _w17649_ ;
	wire _w17648_ ;
	wire _w17647_ ;
	wire _w17646_ ;
	wire _w17645_ ;
	wire _w17644_ ;
	wire _w17643_ ;
	wire _w17642_ ;
	wire _w17641_ ;
	wire _w17640_ ;
	wire _w17639_ ;
	wire _w17638_ ;
	wire _w17637_ ;
	wire _w17636_ ;
	wire _w17635_ ;
	wire _w17634_ ;
	wire _w17633_ ;
	wire _w17632_ ;
	wire _w17631_ ;
	wire _w17630_ ;
	wire _w17629_ ;
	wire _w17628_ ;
	wire _w17627_ ;
	wire _w17626_ ;
	wire _w17625_ ;
	wire _w17624_ ;
	wire _w17623_ ;
	wire _w17622_ ;
	wire _w17621_ ;
	wire _w17620_ ;
	wire _w17619_ ;
	wire _w17618_ ;
	wire _w17617_ ;
	wire _w17616_ ;
	wire _w17615_ ;
	wire _w17614_ ;
	wire _w17613_ ;
	wire _w17612_ ;
	wire _w17611_ ;
	wire _w17610_ ;
	wire _w17609_ ;
	wire _w17608_ ;
	wire _w17607_ ;
	wire _w17606_ ;
	wire _w17605_ ;
	wire _w17604_ ;
	wire _w17603_ ;
	wire _w17602_ ;
	wire _w17601_ ;
	wire _w17600_ ;
	wire _w17599_ ;
	wire _w17598_ ;
	wire _w17597_ ;
	wire _w17596_ ;
	wire _w17595_ ;
	wire _w17594_ ;
	wire _w17593_ ;
	wire _w17592_ ;
	wire _w17591_ ;
	wire _w17590_ ;
	wire _w17589_ ;
	wire _w17588_ ;
	wire _w17587_ ;
	wire _w17586_ ;
	wire _w17585_ ;
	wire _w17584_ ;
	wire _w17583_ ;
	wire _w17582_ ;
	wire _w17581_ ;
	wire _w17580_ ;
	wire _w17579_ ;
	wire _w17578_ ;
	wire _w17577_ ;
	wire _w17576_ ;
	wire _w17575_ ;
	wire _w17574_ ;
	wire _w17573_ ;
	wire _w17572_ ;
	wire _w17571_ ;
	wire _w17570_ ;
	wire _w17569_ ;
	wire _w17568_ ;
	wire _w17567_ ;
	wire _w17566_ ;
	wire _w17565_ ;
	wire _w17564_ ;
	wire _w17563_ ;
	wire _w17562_ ;
	wire _w17561_ ;
	wire _w17560_ ;
	wire _w17559_ ;
	wire _w17558_ ;
	wire _w17557_ ;
	wire _w17556_ ;
	wire _w17555_ ;
	wire _w17554_ ;
	wire _w17553_ ;
	wire _w17552_ ;
	wire _w17551_ ;
	wire _w17550_ ;
	wire _w17549_ ;
	wire _w17548_ ;
	wire _w17547_ ;
	wire _w17546_ ;
	wire _w17545_ ;
	wire _w17544_ ;
	wire _w17543_ ;
	wire _w17542_ ;
	wire _w17541_ ;
	wire _w17540_ ;
	wire _w17539_ ;
	wire _w17538_ ;
	wire _w17537_ ;
	wire _w17536_ ;
	wire _w17535_ ;
	wire _w17534_ ;
	wire _w17533_ ;
	wire _w17532_ ;
	wire _w17531_ ;
	wire _w17530_ ;
	wire _w17529_ ;
	wire _w17528_ ;
	wire _w17527_ ;
	wire _w17526_ ;
	wire _w17525_ ;
	wire _w17524_ ;
	wire _w17523_ ;
	wire _w17522_ ;
	wire _w17521_ ;
	wire _w17520_ ;
	wire _w17519_ ;
	wire _w17518_ ;
	wire _w17517_ ;
	wire _w17516_ ;
	wire _w17515_ ;
	wire _w17514_ ;
	wire _w17513_ ;
	wire _w17512_ ;
	wire _w17511_ ;
	wire _w17510_ ;
	wire _w17509_ ;
	wire _w17508_ ;
	wire _w17507_ ;
	wire _w17506_ ;
	wire _w17505_ ;
	wire _w17504_ ;
	wire _w17503_ ;
	wire _w17502_ ;
	wire _w17501_ ;
	wire _w17500_ ;
	wire _w17499_ ;
	wire _w17498_ ;
	wire _w17497_ ;
	wire _w17496_ ;
	wire _w17495_ ;
	wire _w17494_ ;
	wire _w17493_ ;
	wire _w17492_ ;
	wire _w17491_ ;
	wire _w17490_ ;
	wire _w17489_ ;
	wire _w17488_ ;
	wire _w17487_ ;
	wire _w17486_ ;
	wire _w17485_ ;
	wire _w17484_ ;
	wire _w17483_ ;
	wire _w17482_ ;
	wire _w17481_ ;
	wire _w17480_ ;
	wire _w17479_ ;
	wire _w17478_ ;
	wire _w17477_ ;
	wire _w17476_ ;
	wire _w17475_ ;
	wire _w17474_ ;
	wire _w17473_ ;
	wire _w17472_ ;
	wire _w17471_ ;
	wire _w17470_ ;
	wire _w17469_ ;
	wire _w17468_ ;
	wire _w17467_ ;
	wire _w17466_ ;
	wire _w17465_ ;
	wire _w17464_ ;
	wire _w17463_ ;
	wire _w17462_ ;
	wire _w17461_ ;
	wire _w17460_ ;
	wire _w17459_ ;
	wire _w17458_ ;
	wire _w17457_ ;
	wire _w17456_ ;
	wire _w17455_ ;
	wire _w17454_ ;
	wire _w17453_ ;
	wire _w17452_ ;
	wire _w17451_ ;
	wire _w17450_ ;
	wire _w17449_ ;
	wire _w17448_ ;
	wire _w17447_ ;
	wire _w17446_ ;
	wire _w17445_ ;
	wire _w17444_ ;
	wire _w17443_ ;
	wire _w17442_ ;
	wire _w17441_ ;
	wire _w17440_ ;
	wire _w17439_ ;
	wire _w17438_ ;
	wire _w17437_ ;
	wire _w17436_ ;
	wire _w17435_ ;
	wire _w17434_ ;
	wire _w17433_ ;
	wire _w17432_ ;
	wire _w17431_ ;
	wire _w17430_ ;
	wire _w17429_ ;
	wire _w17428_ ;
	wire _w17427_ ;
	wire _w17426_ ;
	wire _w17425_ ;
	wire _w17424_ ;
	wire _w17423_ ;
	wire _w17422_ ;
	wire _w17421_ ;
	wire _w17420_ ;
	wire _w17419_ ;
	wire _w17418_ ;
	wire _w17417_ ;
	wire _w17416_ ;
	wire _w17415_ ;
	wire _w17414_ ;
	wire _w17413_ ;
	wire _w17412_ ;
	wire _w17411_ ;
	wire _w17410_ ;
	wire _w17409_ ;
	wire _w17408_ ;
	wire _w17407_ ;
	wire _w17406_ ;
	wire _w17405_ ;
	wire _w17404_ ;
	wire _w17403_ ;
	wire _w17402_ ;
	wire _w17401_ ;
	wire _w17400_ ;
	wire _w17399_ ;
	wire _w17398_ ;
	wire _w17397_ ;
	wire _w17396_ ;
	wire _w17395_ ;
	wire _w17394_ ;
	wire _w17393_ ;
	wire _w17392_ ;
	wire _w17391_ ;
	wire _w17390_ ;
	wire _w17389_ ;
	wire _w17388_ ;
	wire _w17387_ ;
	wire _w17386_ ;
	wire _w17385_ ;
	wire _w17384_ ;
	wire _w17383_ ;
	wire _w17382_ ;
	wire _w17381_ ;
	wire _w17380_ ;
	wire _w17379_ ;
	wire _w17378_ ;
	wire _w17377_ ;
	wire _w17376_ ;
	wire _w17375_ ;
	wire _w17374_ ;
	wire _w17373_ ;
	wire _w17372_ ;
	wire _w17371_ ;
	wire _w17370_ ;
	wire _w17369_ ;
	wire _w17368_ ;
	wire _w17367_ ;
	wire _w17366_ ;
	wire _w17365_ ;
	wire _w17364_ ;
	wire _w17363_ ;
	wire _w17362_ ;
	wire _w17361_ ;
	wire _w17360_ ;
	wire _w17359_ ;
	wire _w17358_ ;
	wire _w17357_ ;
	wire _w17356_ ;
	wire _w17355_ ;
	wire _w17354_ ;
	wire _w17353_ ;
	wire _w17352_ ;
	wire _w17351_ ;
	wire _w17350_ ;
	wire _w17349_ ;
	wire _w17348_ ;
	wire _w17347_ ;
	wire _w17346_ ;
	wire _w17345_ ;
	wire _w17344_ ;
	wire _w17343_ ;
	wire _w17342_ ;
	wire _w17341_ ;
	wire _w17340_ ;
	wire _w17339_ ;
	wire _w17338_ ;
	wire _w17337_ ;
	wire _w17336_ ;
	wire _w17335_ ;
	wire _w17334_ ;
	wire _w17333_ ;
	wire _w17332_ ;
	wire _w17331_ ;
	wire _w17330_ ;
	wire _w17329_ ;
	wire _w17328_ ;
	wire _w17327_ ;
	wire _w17326_ ;
	wire _w17325_ ;
	wire _w17324_ ;
	wire _w17323_ ;
	wire _w17322_ ;
	wire _w17321_ ;
	wire _w17320_ ;
	wire _w17319_ ;
	wire _w17318_ ;
	wire _w17317_ ;
	wire _w17316_ ;
	wire _w17315_ ;
	wire _w17314_ ;
	wire _w17313_ ;
	wire _w17312_ ;
	wire _w17311_ ;
	wire _w17310_ ;
	wire _w17309_ ;
	wire _w17308_ ;
	wire _w17307_ ;
	wire _w17306_ ;
	wire _w17305_ ;
	wire _w17304_ ;
	wire _w17303_ ;
	wire _w17302_ ;
	wire _w17301_ ;
	wire _w17300_ ;
	wire _w17299_ ;
	wire _w17298_ ;
	wire _w17297_ ;
	wire _w17296_ ;
	wire _w17295_ ;
	wire _w17294_ ;
	wire _w17293_ ;
	wire _w17292_ ;
	wire _w17291_ ;
	wire _w17290_ ;
	wire _w17289_ ;
	wire _w17288_ ;
	wire _w17287_ ;
	wire _w17286_ ;
	wire _w17285_ ;
	wire _w17284_ ;
	wire _w17283_ ;
	wire _w17282_ ;
	wire _w17281_ ;
	wire _w17280_ ;
	wire _w17279_ ;
	wire _w17278_ ;
	wire _w17277_ ;
	wire _w17276_ ;
	wire _w17275_ ;
	wire _w17274_ ;
	wire _w17273_ ;
	wire _w17272_ ;
	wire _w17271_ ;
	wire _w17270_ ;
	wire _w17269_ ;
	wire _w17268_ ;
	wire _w17267_ ;
	wire _w17266_ ;
	wire _w17265_ ;
	wire _w17264_ ;
	wire _w17263_ ;
	wire _w17262_ ;
	wire _w17261_ ;
	wire _w17260_ ;
	wire _w17259_ ;
	wire _w17258_ ;
	wire _w17257_ ;
	wire _w17256_ ;
	wire _w17255_ ;
	wire _w17254_ ;
	wire _w17253_ ;
	wire _w17252_ ;
	wire _w17251_ ;
	wire _w17250_ ;
	wire _w17249_ ;
	wire _w17248_ ;
	wire _w17247_ ;
	wire _w17246_ ;
	wire _w17245_ ;
	wire _w17244_ ;
	wire _w17243_ ;
	wire _w17242_ ;
	wire _w17241_ ;
	wire _w17240_ ;
	wire _w17239_ ;
	wire _w17238_ ;
	wire _w17237_ ;
	wire _w17236_ ;
	wire _w17235_ ;
	wire _w17234_ ;
	wire _w17233_ ;
	wire _w17232_ ;
	wire _w17231_ ;
	wire _w17230_ ;
	wire _w17229_ ;
	wire _w17228_ ;
	wire _w17227_ ;
	wire _w17226_ ;
	wire _w17225_ ;
	wire _w17224_ ;
	wire _w17223_ ;
	wire _w17222_ ;
	wire _w17221_ ;
	wire _w17220_ ;
	wire _w17219_ ;
	wire _w17218_ ;
	wire _w17217_ ;
	wire _w17216_ ;
	wire _w17215_ ;
	wire _w17214_ ;
	wire _w17213_ ;
	wire _w17212_ ;
	wire _w17211_ ;
	wire _w17210_ ;
	wire _w17209_ ;
	wire _w17208_ ;
	wire _w17207_ ;
	wire _w17206_ ;
	wire _w17205_ ;
	wire _w17204_ ;
	wire _w17203_ ;
	wire _w17202_ ;
	wire _w17201_ ;
	wire _w17200_ ;
	wire _w17199_ ;
	wire _w17198_ ;
	wire _w17197_ ;
	wire _w17196_ ;
	wire _w17195_ ;
	wire _w17194_ ;
	wire _w17193_ ;
	wire _w17192_ ;
	wire _w17191_ ;
	wire _w17190_ ;
	wire _w17189_ ;
	wire _w17188_ ;
	wire _w17187_ ;
	wire _w17186_ ;
	wire _w17185_ ;
	wire _w17184_ ;
	wire _w17183_ ;
	wire _w17182_ ;
	wire _w17181_ ;
	wire _w17180_ ;
	wire _w17179_ ;
	wire _w17178_ ;
	wire _w17177_ ;
	wire _w17176_ ;
	wire _w17175_ ;
	wire _w17174_ ;
	wire _w17173_ ;
	wire _w17172_ ;
	wire _w17171_ ;
	wire _w17170_ ;
	wire _w17169_ ;
	wire _w17168_ ;
	wire _w17167_ ;
	wire _w17166_ ;
	wire _w17165_ ;
	wire _w17164_ ;
	wire _w17163_ ;
	wire _w17162_ ;
	wire _w17161_ ;
	wire _w17160_ ;
	wire _w17159_ ;
	wire _w17158_ ;
	wire _w17157_ ;
	wire _w17156_ ;
	wire _w17155_ ;
	wire _w17154_ ;
	wire _w17153_ ;
	wire _w17152_ ;
	wire _w17151_ ;
	wire _w17150_ ;
	wire _w17149_ ;
	wire _w17148_ ;
	wire _w17147_ ;
	wire _w17146_ ;
	wire _w17145_ ;
	wire _w17144_ ;
	wire _w17143_ ;
	wire _w17142_ ;
	wire _w17141_ ;
	wire _w17140_ ;
	wire _w17139_ ;
	wire _w17138_ ;
	wire _w17137_ ;
	wire _w17136_ ;
	wire _w17135_ ;
	wire _w17134_ ;
	wire _w17133_ ;
	wire _w17132_ ;
	wire _w17131_ ;
	wire _w17130_ ;
	wire _w17129_ ;
	wire _w17128_ ;
	wire _w17127_ ;
	wire _w17126_ ;
	wire _w17125_ ;
	wire _w17124_ ;
	wire _w17123_ ;
	wire _w17122_ ;
	wire _w17121_ ;
	wire _w17120_ ;
	wire _w17119_ ;
	wire _w17118_ ;
	wire _w17117_ ;
	wire _w17116_ ;
	wire _w17115_ ;
	wire _w17114_ ;
	wire _w17113_ ;
	wire _w17112_ ;
	wire _w17111_ ;
	wire _w17110_ ;
	wire _w17109_ ;
	wire _w17108_ ;
	wire _w17107_ ;
	wire _w17106_ ;
	wire _w17105_ ;
	wire _w17104_ ;
	wire _w17103_ ;
	wire _w17102_ ;
	wire _w17101_ ;
	wire _w17100_ ;
	wire _w17099_ ;
	wire _w17098_ ;
	wire _w17097_ ;
	wire _w17096_ ;
	wire _w17095_ ;
	wire _w17094_ ;
	wire _w17093_ ;
	wire _w17092_ ;
	wire _w17091_ ;
	wire _w17090_ ;
	wire _w17089_ ;
	wire _w17088_ ;
	wire _w17087_ ;
	wire _w17086_ ;
	wire _w17085_ ;
	wire _w17084_ ;
	wire _w17083_ ;
	wire _w17082_ ;
	wire _w17081_ ;
	wire _w17080_ ;
	wire _w17079_ ;
	wire _w17078_ ;
	wire _w17077_ ;
	wire _w17076_ ;
	wire _w17075_ ;
	wire _w17074_ ;
	wire _w17073_ ;
	wire _w17072_ ;
	wire _w17071_ ;
	wire _w17070_ ;
	wire _w17069_ ;
	wire _w17068_ ;
	wire _w17067_ ;
	wire _w17066_ ;
	wire _w17065_ ;
	wire _w17064_ ;
	wire _w17063_ ;
	wire _w17062_ ;
	wire _w17061_ ;
	wire _w17060_ ;
	wire _w17059_ ;
	wire _w17058_ ;
	wire _w17057_ ;
	wire _w17056_ ;
	wire _w17055_ ;
	wire _w17054_ ;
	wire _w17053_ ;
	wire _w17052_ ;
	wire _w17051_ ;
	wire _w17050_ ;
	wire _w17049_ ;
	wire _w17048_ ;
	wire _w17047_ ;
	wire _w17046_ ;
	wire _w17045_ ;
	wire _w17044_ ;
	wire _w17043_ ;
	wire _w17042_ ;
	wire _w17041_ ;
	wire _w17040_ ;
	wire _w17039_ ;
	wire _w17038_ ;
	wire _w17037_ ;
	wire _w17036_ ;
	wire _w17035_ ;
	wire _w17034_ ;
	wire _w17033_ ;
	wire _w17032_ ;
	wire _w17031_ ;
	wire _w17030_ ;
	wire _w17029_ ;
	wire _w17028_ ;
	wire _w17027_ ;
	wire _w17026_ ;
	wire _w17025_ ;
	wire _w17024_ ;
	wire _w17023_ ;
	wire _w17022_ ;
	wire _w17021_ ;
	wire _w17020_ ;
	wire _w17019_ ;
	wire _w17018_ ;
	wire _w17017_ ;
	wire _w17016_ ;
	wire _w17015_ ;
	wire _w17014_ ;
	wire _w17013_ ;
	wire _w17012_ ;
	wire _w17011_ ;
	wire _w17010_ ;
	wire _w17009_ ;
	wire _w17008_ ;
	wire _w17007_ ;
	wire _w17006_ ;
	wire _w17005_ ;
	wire _w17004_ ;
	wire _w17003_ ;
	wire _w17002_ ;
	wire _w17001_ ;
	wire _w17000_ ;
	wire _w16999_ ;
	wire _w16998_ ;
	wire _w16997_ ;
	wire _w16996_ ;
	wire _w16995_ ;
	wire _w16994_ ;
	wire _w16993_ ;
	wire _w16992_ ;
	wire _w16991_ ;
	wire _w16990_ ;
	wire _w16989_ ;
	wire _w16988_ ;
	wire _w16987_ ;
	wire _w16986_ ;
	wire _w16985_ ;
	wire _w16984_ ;
	wire _w16983_ ;
	wire _w16982_ ;
	wire _w16981_ ;
	wire _w16980_ ;
	wire _w16979_ ;
	wire _w16978_ ;
	wire _w16977_ ;
	wire _w16976_ ;
	wire _w16975_ ;
	wire _w16974_ ;
	wire _w16973_ ;
	wire _w16972_ ;
	wire _w16971_ ;
	wire _w16970_ ;
	wire _w16969_ ;
	wire _w16968_ ;
	wire _w16967_ ;
	wire _w16966_ ;
	wire _w16965_ ;
	wire _w16964_ ;
	wire _w16963_ ;
	wire _w16962_ ;
	wire _w16961_ ;
	wire _w16960_ ;
	wire _w16959_ ;
	wire _w16958_ ;
	wire _w16957_ ;
	wire _w16956_ ;
	wire _w16955_ ;
	wire _w16954_ ;
	wire _w16953_ ;
	wire _w16952_ ;
	wire _w16951_ ;
	wire _w16950_ ;
	wire _w16949_ ;
	wire _w16948_ ;
	wire _w16947_ ;
	wire _w16946_ ;
	wire _w16945_ ;
	wire _w16944_ ;
	wire _w16943_ ;
	wire _w16942_ ;
	wire _w16941_ ;
	wire _w16940_ ;
	wire _w16939_ ;
	wire _w16938_ ;
	wire _w16937_ ;
	wire _w16936_ ;
	wire _w16935_ ;
	wire _w16934_ ;
	wire _w16933_ ;
	wire _w16932_ ;
	wire _w16931_ ;
	wire _w16930_ ;
	wire _w16929_ ;
	wire _w16928_ ;
	wire _w16927_ ;
	wire _w16926_ ;
	wire _w16925_ ;
	wire _w16924_ ;
	wire _w16923_ ;
	wire _w16922_ ;
	wire _w16921_ ;
	wire _w16920_ ;
	wire _w16919_ ;
	wire _w16918_ ;
	wire _w16917_ ;
	wire _w16916_ ;
	wire _w16915_ ;
	wire _w16914_ ;
	wire _w16913_ ;
	wire _w16912_ ;
	wire _w16911_ ;
	wire _w16910_ ;
	wire _w16909_ ;
	wire _w16908_ ;
	wire _w16907_ ;
	wire _w16906_ ;
	wire _w16905_ ;
	wire _w16904_ ;
	wire _w16903_ ;
	wire _w16902_ ;
	wire _w16901_ ;
	wire _w16900_ ;
	wire _w16899_ ;
	wire _w16898_ ;
	wire _w16897_ ;
	wire _w16896_ ;
	wire _w16895_ ;
	wire _w16894_ ;
	wire _w16893_ ;
	wire _w16892_ ;
	wire _w16891_ ;
	wire _w16890_ ;
	wire _w16889_ ;
	wire _w16888_ ;
	wire _w16887_ ;
	wire _w16886_ ;
	wire _w16885_ ;
	wire _w16884_ ;
	wire _w16883_ ;
	wire _w16882_ ;
	wire _w16881_ ;
	wire _w16880_ ;
	wire _w16879_ ;
	wire _w16878_ ;
	wire _w16877_ ;
	wire _w16876_ ;
	wire _w16875_ ;
	wire _w16874_ ;
	wire _w16873_ ;
	wire _w16872_ ;
	wire _w16871_ ;
	wire _w16870_ ;
	wire _w16869_ ;
	wire _w16868_ ;
	wire _w16867_ ;
	wire _w16866_ ;
	wire _w16865_ ;
	wire _w16864_ ;
	wire _w16863_ ;
	wire _w16862_ ;
	wire _w16861_ ;
	wire _w16860_ ;
	wire _w16859_ ;
	wire _w16858_ ;
	wire _w16857_ ;
	wire _w16856_ ;
	wire _w16855_ ;
	wire _w16854_ ;
	wire _w16853_ ;
	wire _w16852_ ;
	wire _w16851_ ;
	wire _w16850_ ;
	wire _w16849_ ;
	wire _w16848_ ;
	wire _w16847_ ;
	wire _w16846_ ;
	wire _w16845_ ;
	wire _w16844_ ;
	wire _w16843_ ;
	wire _w16842_ ;
	wire _w16841_ ;
	wire _w16840_ ;
	wire _w16839_ ;
	wire _w16838_ ;
	wire _w16837_ ;
	wire _w16836_ ;
	wire _w16835_ ;
	wire _w16834_ ;
	wire _w16833_ ;
	wire _w16832_ ;
	wire _w16831_ ;
	wire _w16830_ ;
	wire _w16829_ ;
	wire _w16828_ ;
	wire _w16827_ ;
	wire _w16826_ ;
	wire _w16825_ ;
	wire _w16824_ ;
	wire _w16823_ ;
	wire _w16822_ ;
	wire _w16821_ ;
	wire _w16820_ ;
	wire _w16819_ ;
	wire _w16818_ ;
	wire _w16817_ ;
	wire _w16816_ ;
	wire _w16815_ ;
	wire _w16814_ ;
	wire _w16813_ ;
	wire _w16812_ ;
	wire _w16811_ ;
	wire _w16810_ ;
	wire _w16809_ ;
	wire _w16808_ ;
	wire _w16807_ ;
	wire _w16806_ ;
	wire _w16805_ ;
	wire _w16804_ ;
	wire _w16803_ ;
	wire _w16802_ ;
	wire _w16801_ ;
	wire _w16800_ ;
	wire _w16799_ ;
	wire _w16798_ ;
	wire _w16797_ ;
	wire _w16796_ ;
	wire _w16795_ ;
	wire _w16794_ ;
	wire _w16793_ ;
	wire _w16792_ ;
	wire _w16791_ ;
	wire _w16790_ ;
	wire _w16789_ ;
	wire _w16788_ ;
	wire _w16787_ ;
	wire _w16786_ ;
	wire _w16785_ ;
	wire _w16784_ ;
	wire _w16783_ ;
	wire _w16782_ ;
	wire _w16781_ ;
	wire _w16780_ ;
	wire _w16779_ ;
	wire _w16778_ ;
	wire _w16777_ ;
	wire _w16776_ ;
	wire _w16775_ ;
	wire _w16774_ ;
	wire _w16773_ ;
	wire _w16772_ ;
	wire _w16771_ ;
	wire _w16770_ ;
	wire _w16769_ ;
	wire _w16768_ ;
	wire _w16767_ ;
	wire _w16766_ ;
	wire _w16765_ ;
	wire _w16764_ ;
	wire _w16763_ ;
	wire _w16762_ ;
	wire _w16761_ ;
	wire _w16760_ ;
	wire _w16759_ ;
	wire _w16758_ ;
	wire _w16757_ ;
	wire _w16756_ ;
	wire _w16755_ ;
	wire _w16754_ ;
	wire _w16753_ ;
	wire _w16752_ ;
	wire _w16751_ ;
	wire _w16750_ ;
	wire _w16749_ ;
	wire _w16748_ ;
	wire _w16747_ ;
	wire _w16746_ ;
	wire _w16745_ ;
	wire _w16744_ ;
	wire _w16743_ ;
	wire _w16742_ ;
	wire _w16741_ ;
	wire _w16740_ ;
	wire _w16739_ ;
	wire _w16738_ ;
	wire _w16737_ ;
	wire _w16736_ ;
	wire _w16735_ ;
	wire _w16734_ ;
	wire _w16733_ ;
	wire _w16732_ ;
	wire _w16731_ ;
	wire _w16730_ ;
	wire _w16729_ ;
	wire _w16728_ ;
	wire _w16727_ ;
	wire _w16726_ ;
	wire _w16725_ ;
	wire _w16724_ ;
	wire _w16723_ ;
	wire _w16722_ ;
	wire _w16721_ ;
	wire _w16720_ ;
	wire _w16719_ ;
	wire _w16718_ ;
	wire _w16717_ ;
	wire _w16716_ ;
	wire _w16715_ ;
	wire _w16714_ ;
	wire _w16713_ ;
	wire _w16712_ ;
	wire _w16711_ ;
	wire _w16710_ ;
	wire _w16709_ ;
	wire _w16708_ ;
	wire _w16707_ ;
	wire _w16706_ ;
	wire _w16705_ ;
	wire _w16704_ ;
	wire _w16703_ ;
	wire _w16702_ ;
	wire _w16701_ ;
	wire _w16700_ ;
	wire _w16699_ ;
	wire _w16698_ ;
	wire _w16697_ ;
	wire _w16696_ ;
	wire _w16695_ ;
	wire _w16694_ ;
	wire _w16693_ ;
	wire _w16692_ ;
	wire _w16691_ ;
	wire _w16690_ ;
	wire _w16689_ ;
	wire _w16688_ ;
	wire _w16687_ ;
	wire _w16686_ ;
	wire _w16685_ ;
	wire _w16684_ ;
	wire _w16683_ ;
	wire _w16682_ ;
	wire _w16681_ ;
	wire _w16680_ ;
	wire _w16679_ ;
	wire _w16678_ ;
	wire _w16677_ ;
	wire _w16676_ ;
	wire _w16675_ ;
	wire _w16674_ ;
	wire _w16673_ ;
	wire _w16672_ ;
	wire _w16671_ ;
	wire _w16670_ ;
	wire _w16669_ ;
	wire _w16668_ ;
	wire _w16667_ ;
	wire _w16666_ ;
	wire _w16665_ ;
	wire _w16664_ ;
	wire _w16663_ ;
	wire _w16662_ ;
	wire _w16661_ ;
	wire _w16660_ ;
	wire _w16659_ ;
	wire _w16658_ ;
	wire _w16657_ ;
	wire _w16656_ ;
	wire _w16655_ ;
	wire _w16654_ ;
	wire _w16653_ ;
	wire _w16652_ ;
	wire _w16651_ ;
	wire _w16650_ ;
	wire _w16649_ ;
	wire _w16648_ ;
	wire _w16647_ ;
	wire _w16646_ ;
	wire _w16645_ ;
	wire _w16644_ ;
	wire _w16643_ ;
	wire _w16642_ ;
	wire _w16641_ ;
	wire _w16640_ ;
	wire _w16639_ ;
	wire _w16638_ ;
	wire _w16637_ ;
	wire _w16636_ ;
	wire _w16635_ ;
	wire _w16634_ ;
	wire _w16633_ ;
	wire _w16632_ ;
	wire _w16631_ ;
	wire _w16630_ ;
	wire _w16629_ ;
	wire _w16628_ ;
	wire _w16627_ ;
	wire _w16626_ ;
	wire _w16625_ ;
	wire _w16624_ ;
	wire _w16623_ ;
	wire _w16622_ ;
	wire _w16621_ ;
	wire _w16620_ ;
	wire _w16619_ ;
	wire _w16618_ ;
	wire _w16617_ ;
	wire _w16616_ ;
	wire _w16615_ ;
	wire _w16614_ ;
	wire _w16613_ ;
	wire _w16612_ ;
	wire _w16611_ ;
	wire _w16610_ ;
	wire _w16609_ ;
	wire _w16608_ ;
	wire _w16607_ ;
	wire _w16606_ ;
	wire _w16605_ ;
	wire _w16604_ ;
	wire _w16603_ ;
	wire _w16602_ ;
	wire _w16601_ ;
	wire _w16600_ ;
	wire _w16599_ ;
	wire _w16598_ ;
	wire _w16597_ ;
	wire _w16596_ ;
	wire _w16595_ ;
	wire _w16594_ ;
	wire _w16593_ ;
	wire _w16592_ ;
	wire _w16591_ ;
	wire _w16590_ ;
	wire _w16589_ ;
	wire _w16588_ ;
	wire _w16587_ ;
	wire _w16586_ ;
	wire _w16585_ ;
	wire _w16584_ ;
	wire _w16583_ ;
	wire _w16582_ ;
	wire _w16581_ ;
	wire _w16580_ ;
	wire _w16579_ ;
	wire _w16578_ ;
	wire _w16577_ ;
	wire _w16576_ ;
	wire _w16575_ ;
	wire _w16574_ ;
	wire _w16573_ ;
	wire _w16572_ ;
	wire _w16571_ ;
	wire _w16570_ ;
	wire _w16569_ ;
	wire _w16568_ ;
	wire _w16567_ ;
	wire _w16566_ ;
	wire _w16565_ ;
	wire _w16564_ ;
	wire _w16563_ ;
	wire _w16562_ ;
	wire _w16561_ ;
	wire _w16560_ ;
	wire _w16559_ ;
	wire _w16558_ ;
	wire _w16557_ ;
	wire _w16556_ ;
	wire _w16555_ ;
	wire _w16554_ ;
	wire _w16553_ ;
	wire _w16552_ ;
	wire _w16551_ ;
	wire _w16550_ ;
	wire _w16549_ ;
	wire _w16548_ ;
	wire _w16547_ ;
	wire _w16546_ ;
	wire _w16545_ ;
	wire _w16544_ ;
	wire _w16543_ ;
	wire _w16542_ ;
	wire _w16541_ ;
	wire _w16540_ ;
	wire _w16539_ ;
	wire _w16538_ ;
	wire _w16537_ ;
	wire _w16536_ ;
	wire _w16535_ ;
	wire _w16534_ ;
	wire _w16533_ ;
	wire _w16532_ ;
	wire _w16531_ ;
	wire _w16530_ ;
	wire _w16529_ ;
	wire _w16528_ ;
	wire _w16527_ ;
	wire _w16526_ ;
	wire _w16525_ ;
	wire _w16524_ ;
	wire _w16523_ ;
	wire _w16522_ ;
	wire _w16521_ ;
	wire _w16520_ ;
	wire _w16519_ ;
	wire _w16518_ ;
	wire _w16517_ ;
	wire _w16516_ ;
	wire _w16515_ ;
	wire _w16514_ ;
	wire _w16513_ ;
	wire _w16512_ ;
	wire _w16511_ ;
	wire _w16510_ ;
	wire _w16509_ ;
	wire _w16508_ ;
	wire _w16507_ ;
	wire _w16506_ ;
	wire _w16505_ ;
	wire _w16504_ ;
	wire _w16503_ ;
	wire _w16502_ ;
	wire _w16501_ ;
	wire _w16500_ ;
	wire _w16499_ ;
	wire _w16498_ ;
	wire _w16497_ ;
	wire _w16496_ ;
	wire _w16495_ ;
	wire _w16494_ ;
	wire _w16493_ ;
	wire _w16492_ ;
	wire _w16491_ ;
	wire _w16490_ ;
	wire _w16489_ ;
	wire _w16488_ ;
	wire _w16487_ ;
	wire _w16486_ ;
	wire _w16485_ ;
	wire _w16484_ ;
	wire _w16483_ ;
	wire _w16482_ ;
	wire _w16481_ ;
	wire _w16480_ ;
	wire _w16479_ ;
	wire _w16478_ ;
	wire _w16477_ ;
	wire _w16476_ ;
	wire _w16475_ ;
	wire _w16474_ ;
	wire _w16473_ ;
	wire _w16472_ ;
	wire _w16471_ ;
	wire _w16470_ ;
	wire _w16469_ ;
	wire _w16468_ ;
	wire _w16467_ ;
	wire _w16466_ ;
	wire _w16465_ ;
	wire _w16464_ ;
	wire _w16463_ ;
	wire _w16462_ ;
	wire _w16461_ ;
	wire _w16460_ ;
	wire _w16459_ ;
	wire _w16458_ ;
	wire _w16457_ ;
	wire _w16456_ ;
	wire _w16455_ ;
	wire _w16454_ ;
	wire _w16453_ ;
	wire _w16452_ ;
	wire _w16451_ ;
	wire _w16450_ ;
	wire _w16449_ ;
	wire _w16448_ ;
	wire _w16447_ ;
	wire _w16446_ ;
	wire _w16445_ ;
	wire _w16444_ ;
	wire _w16443_ ;
	wire _w16442_ ;
	wire _w16441_ ;
	wire _w16440_ ;
	wire _w16439_ ;
	wire _w16438_ ;
	wire _w16437_ ;
	wire _w16436_ ;
	wire _w16435_ ;
	wire _w16434_ ;
	wire _w16433_ ;
	wire _w16432_ ;
	wire _w16431_ ;
	wire _w16430_ ;
	wire _w16429_ ;
	wire _w16428_ ;
	wire _w16427_ ;
	wire _w16426_ ;
	wire _w16425_ ;
	wire _w16424_ ;
	wire _w16423_ ;
	wire _w16422_ ;
	wire _w16421_ ;
	wire _w16420_ ;
	wire _w16419_ ;
	wire _w16418_ ;
	wire _w16417_ ;
	wire _w16416_ ;
	wire _w16415_ ;
	wire _w16414_ ;
	wire _w16413_ ;
	wire _w16412_ ;
	wire _w16411_ ;
	wire _w16410_ ;
	wire _w16409_ ;
	wire _w16408_ ;
	wire _w16407_ ;
	wire _w16406_ ;
	wire _w16405_ ;
	wire _w16404_ ;
	wire _w16403_ ;
	wire _w16402_ ;
	wire _w16401_ ;
	wire _w16400_ ;
	wire _w16399_ ;
	wire _w16398_ ;
	wire _w16397_ ;
	wire _w16396_ ;
	wire _w16395_ ;
	wire _w16394_ ;
	wire _w16393_ ;
	wire _w16392_ ;
	wire _w16391_ ;
	wire _w16390_ ;
	wire _w16389_ ;
	wire _w16388_ ;
	wire _w16387_ ;
	wire _w16386_ ;
	wire _w16385_ ;
	wire _w16384_ ;
	wire _w16383_ ;
	wire _w16382_ ;
	wire _w16381_ ;
	wire _w16380_ ;
	wire _w16379_ ;
	wire _w16378_ ;
	wire _w16377_ ;
	wire _w16376_ ;
	wire _w16375_ ;
	wire _w16374_ ;
	wire _w16373_ ;
	wire _w16372_ ;
	wire _w16371_ ;
	wire _w16370_ ;
	wire _w16369_ ;
	wire _w16368_ ;
	wire _w16367_ ;
	wire _w16366_ ;
	wire _w16365_ ;
	wire _w16364_ ;
	wire _w16363_ ;
	wire _w16362_ ;
	wire _w16361_ ;
	wire _w16360_ ;
	wire _w16359_ ;
	wire _w16358_ ;
	wire _w16357_ ;
	wire _w16356_ ;
	wire _w16355_ ;
	wire _w16354_ ;
	wire _w16353_ ;
	wire _w16352_ ;
	wire _w16351_ ;
	wire _w16350_ ;
	wire _w16349_ ;
	wire _w16348_ ;
	wire _w16347_ ;
	wire _w16346_ ;
	wire _w16345_ ;
	wire _w16344_ ;
	wire _w16343_ ;
	wire _w16342_ ;
	wire _w16341_ ;
	wire _w16340_ ;
	wire _w16339_ ;
	wire _w16338_ ;
	wire _w16337_ ;
	wire _w16336_ ;
	wire _w16335_ ;
	wire _w16334_ ;
	wire _w16333_ ;
	wire _w16332_ ;
	wire _w16331_ ;
	wire _w16330_ ;
	wire _w16329_ ;
	wire _w16328_ ;
	wire _w16327_ ;
	wire _w16326_ ;
	wire _w16325_ ;
	wire _w16324_ ;
	wire _w16323_ ;
	wire _w16322_ ;
	wire _w16321_ ;
	wire _w16320_ ;
	wire _w16319_ ;
	wire _w16318_ ;
	wire _w16317_ ;
	wire _w16316_ ;
	wire _w16315_ ;
	wire _w16314_ ;
	wire _w16313_ ;
	wire _w16312_ ;
	wire _w16311_ ;
	wire _w16310_ ;
	wire _w16309_ ;
	wire _w16308_ ;
	wire _w16307_ ;
	wire _w16306_ ;
	wire _w16305_ ;
	wire _w16304_ ;
	wire _w16303_ ;
	wire _w16302_ ;
	wire _w16301_ ;
	wire _w16300_ ;
	wire _w16299_ ;
	wire _w16298_ ;
	wire _w16297_ ;
	wire _w16296_ ;
	wire _w16295_ ;
	wire _w16294_ ;
	wire _w16293_ ;
	wire _w16292_ ;
	wire _w16291_ ;
	wire _w16290_ ;
	wire _w16289_ ;
	wire _w16288_ ;
	wire _w16287_ ;
	wire _w16286_ ;
	wire _w16285_ ;
	wire _w16284_ ;
	wire _w16283_ ;
	wire _w16282_ ;
	wire _w16281_ ;
	wire _w16280_ ;
	wire _w16279_ ;
	wire _w16278_ ;
	wire _w16277_ ;
	wire _w16276_ ;
	wire _w16275_ ;
	wire _w16274_ ;
	wire _w16273_ ;
	wire _w16272_ ;
	wire _w16271_ ;
	wire _w16270_ ;
	wire _w16269_ ;
	wire _w16268_ ;
	wire _w16267_ ;
	wire _w16266_ ;
	wire _w16265_ ;
	wire _w16264_ ;
	wire _w16263_ ;
	wire _w16262_ ;
	wire _w16261_ ;
	wire _w16260_ ;
	wire _w16259_ ;
	wire _w16258_ ;
	wire _w16257_ ;
	wire _w16256_ ;
	wire _w16255_ ;
	wire _w16254_ ;
	wire _w16253_ ;
	wire _w16252_ ;
	wire _w16251_ ;
	wire _w16250_ ;
	wire _w16249_ ;
	wire _w16248_ ;
	wire _w16247_ ;
	wire _w16246_ ;
	wire _w16245_ ;
	wire _w16244_ ;
	wire _w16243_ ;
	wire _w16242_ ;
	wire _w16241_ ;
	wire _w16240_ ;
	wire _w16239_ ;
	wire _w16238_ ;
	wire _w16237_ ;
	wire _w16236_ ;
	wire _w16235_ ;
	wire _w16234_ ;
	wire _w16233_ ;
	wire _w16232_ ;
	wire _w16231_ ;
	wire _w16230_ ;
	wire _w16229_ ;
	wire _w16228_ ;
	wire _w16227_ ;
	wire _w16226_ ;
	wire _w16225_ ;
	wire _w16224_ ;
	wire _w16223_ ;
	wire _w16222_ ;
	wire _w16221_ ;
	wire _w16220_ ;
	wire _w16219_ ;
	wire _w16218_ ;
	wire _w16217_ ;
	wire _w16216_ ;
	wire _w16215_ ;
	wire _w16214_ ;
	wire _w16213_ ;
	wire _w16212_ ;
	wire _w16211_ ;
	wire _w16210_ ;
	wire _w16209_ ;
	wire _w16208_ ;
	wire _w16207_ ;
	wire _w16206_ ;
	wire _w16205_ ;
	wire _w16204_ ;
	wire _w16203_ ;
	wire _w16202_ ;
	wire _w16201_ ;
	wire _w16200_ ;
	wire _w16199_ ;
	wire _w16198_ ;
	wire _w16197_ ;
	wire _w16196_ ;
	wire _w16195_ ;
	wire _w16194_ ;
	wire _w16193_ ;
	wire _w16192_ ;
	wire _w16191_ ;
	wire _w16190_ ;
	wire _w16189_ ;
	wire _w16188_ ;
	wire _w16187_ ;
	wire _w16186_ ;
	wire _w16185_ ;
	wire _w16184_ ;
	wire _w16183_ ;
	wire _w16182_ ;
	wire _w16181_ ;
	wire _w16180_ ;
	wire _w16179_ ;
	wire _w16178_ ;
	wire _w16177_ ;
	wire _w16176_ ;
	wire _w16175_ ;
	wire _w16174_ ;
	wire _w16173_ ;
	wire _w16172_ ;
	wire _w16171_ ;
	wire _w16170_ ;
	wire _w16169_ ;
	wire _w16168_ ;
	wire _w16167_ ;
	wire _w16166_ ;
	wire _w16165_ ;
	wire _w16164_ ;
	wire _w16163_ ;
	wire _w16162_ ;
	wire _w16161_ ;
	wire _w16160_ ;
	wire _w16159_ ;
	wire _w16158_ ;
	wire _w16157_ ;
	wire _w16156_ ;
	wire _w16155_ ;
	wire _w16154_ ;
	wire _w16153_ ;
	wire _w16152_ ;
	wire _w16151_ ;
	wire _w16150_ ;
	wire _w16149_ ;
	wire _w16148_ ;
	wire _w16147_ ;
	wire _w16146_ ;
	wire _w16145_ ;
	wire _w16144_ ;
	wire _w16143_ ;
	wire _w16142_ ;
	wire _w16141_ ;
	wire _w16140_ ;
	wire _w16139_ ;
	wire _w16138_ ;
	wire _w16137_ ;
	wire _w16136_ ;
	wire _w16135_ ;
	wire _w16134_ ;
	wire _w16133_ ;
	wire _w16132_ ;
	wire _w16131_ ;
	wire _w16130_ ;
	wire _w16129_ ;
	wire _w16128_ ;
	wire _w16127_ ;
	wire _w16126_ ;
	wire _w16125_ ;
	wire _w16124_ ;
	wire _w16123_ ;
	wire _w16122_ ;
	wire _w16121_ ;
	wire _w16120_ ;
	wire _w16119_ ;
	wire _w16118_ ;
	wire _w16117_ ;
	wire _w16116_ ;
	wire _w16115_ ;
	wire _w16114_ ;
	wire _w16113_ ;
	wire _w16112_ ;
	wire _w16111_ ;
	wire _w16110_ ;
	wire _w16109_ ;
	wire _w16108_ ;
	wire _w16107_ ;
	wire _w16106_ ;
	wire _w16105_ ;
	wire _w16104_ ;
	wire _w16103_ ;
	wire _w16102_ ;
	wire _w16101_ ;
	wire _w16100_ ;
	wire _w16099_ ;
	wire _w16098_ ;
	wire _w16097_ ;
	wire _w16096_ ;
	wire _w16095_ ;
	wire _w16094_ ;
	wire _w16093_ ;
	wire _w16092_ ;
	wire _w16091_ ;
	wire _w16090_ ;
	wire _w16089_ ;
	wire _w16088_ ;
	wire _w16087_ ;
	wire _w16086_ ;
	wire _w16085_ ;
	wire _w16084_ ;
	wire _w16083_ ;
	wire _w16082_ ;
	wire _w16081_ ;
	wire _w16080_ ;
	wire _w16079_ ;
	wire _w16078_ ;
	wire _w16077_ ;
	wire _w16076_ ;
	wire _w16075_ ;
	wire _w16074_ ;
	wire _w16073_ ;
	wire _w16072_ ;
	wire _w16071_ ;
	wire _w16070_ ;
	wire _w16069_ ;
	wire _w16068_ ;
	wire _w16067_ ;
	wire _w16066_ ;
	wire _w16065_ ;
	wire _w16064_ ;
	wire _w16063_ ;
	wire _w16062_ ;
	wire _w16061_ ;
	wire _w16060_ ;
	wire _w16059_ ;
	wire _w16058_ ;
	wire _w16057_ ;
	wire _w16056_ ;
	wire _w16055_ ;
	wire _w16054_ ;
	wire _w16053_ ;
	wire _w16052_ ;
	wire _w16051_ ;
	wire _w16050_ ;
	wire _w16049_ ;
	wire _w16048_ ;
	wire _w16047_ ;
	wire _w16046_ ;
	wire _w16045_ ;
	wire _w16044_ ;
	wire _w16043_ ;
	wire _w16042_ ;
	wire _w16041_ ;
	wire _w16040_ ;
	wire _w16039_ ;
	wire _w16038_ ;
	wire _w16037_ ;
	wire _w16036_ ;
	wire _w16035_ ;
	wire _w16034_ ;
	wire _w16033_ ;
	wire _w16032_ ;
	wire _w16031_ ;
	wire _w16030_ ;
	wire _w16029_ ;
	wire _w16028_ ;
	wire _w16027_ ;
	wire _w16026_ ;
	wire _w16025_ ;
	wire _w16024_ ;
	wire _w16023_ ;
	wire _w16022_ ;
	wire _w16021_ ;
	wire _w16020_ ;
	wire _w16019_ ;
	wire _w16018_ ;
	wire _w16017_ ;
	wire _w16016_ ;
	wire _w16015_ ;
	wire _w16014_ ;
	wire _w16013_ ;
	wire _w16012_ ;
	wire _w16011_ ;
	wire _w16010_ ;
	wire _w16009_ ;
	wire _w16008_ ;
	wire _w16007_ ;
	wire _w16006_ ;
	wire _w16005_ ;
	wire _w16004_ ;
	wire _w16003_ ;
	wire _w16002_ ;
	wire _w16001_ ;
	wire _w16000_ ;
	wire _w15999_ ;
	wire _w15998_ ;
	wire _w15997_ ;
	wire _w15996_ ;
	wire _w15995_ ;
	wire _w15994_ ;
	wire _w15993_ ;
	wire _w15992_ ;
	wire _w15991_ ;
	wire _w15990_ ;
	wire _w15989_ ;
	wire _w15988_ ;
	wire _w15987_ ;
	wire _w15986_ ;
	wire _w15985_ ;
	wire _w15984_ ;
	wire _w15983_ ;
	wire _w15982_ ;
	wire _w15981_ ;
	wire _w15980_ ;
	wire _w15979_ ;
	wire _w15978_ ;
	wire _w15977_ ;
	wire _w15976_ ;
	wire _w15975_ ;
	wire _w15974_ ;
	wire _w15973_ ;
	wire _w15972_ ;
	wire _w15971_ ;
	wire _w15970_ ;
	wire _w15969_ ;
	wire _w15968_ ;
	wire _w15967_ ;
	wire _w15966_ ;
	wire _w15965_ ;
	wire _w15964_ ;
	wire _w15963_ ;
	wire _w15962_ ;
	wire _w15961_ ;
	wire _w15960_ ;
	wire _w15959_ ;
	wire _w15958_ ;
	wire _w15957_ ;
	wire _w15956_ ;
	wire _w15955_ ;
	wire _w15954_ ;
	wire _w15953_ ;
	wire _w15952_ ;
	wire _w15951_ ;
	wire _w15950_ ;
	wire _w15949_ ;
	wire _w15948_ ;
	wire _w15947_ ;
	wire _w15946_ ;
	wire _w15945_ ;
	wire _w15944_ ;
	wire _w15943_ ;
	wire _w15942_ ;
	wire _w15941_ ;
	wire _w15940_ ;
	wire _w15939_ ;
	wire _w15938_ ;
	wire _w15937_ ;
	wire _w15936_ ;
	wire _w15935_ ;
	wire _w15934_ ;
	wire _w15933_ ;
	wire _w15932_ ;
	wire _w15931_ ;
	wire _w15930_ ;
	wire _w15929_ ;
	wire _w15928_ ;
	wire _w15927_ ;
	wire _w15926_ ;
	wire _w15925_ ;
	wire _w15924_ ;
	wire _w15923_ ;
	wire _w15922_ ;
	wire _w15921_ ;
	wire _w15920_ ;
	wire _w15919_ ;
	wire _w15918_ ;
	wire _w15917_ ;
	wire _w15916_ ;
	wire _w15915_ ;
	wire _w15914_ ;
	wire _w15913_ ;
	wire _w15912_ ;
	wire _w15911_ ;
	wire _w15910_ ;
	wire _w15909_ ;
	wire _w15908_ ;
	wire _w15907_ ;
	wire _w15906_ ;
	wire _w15905_ ;
	wire _w15904_ ;
	wire _w15903_ ;
	wire _w15902_ ;
	wire _w15901_ ;
	wire _w15900_ ;
	wire _w15899_ ;
	wire _w15898_ ;
	wire _w15897_ ;
	wire _w15896_ ;
	wire _w15895_ ;
	wire _w15894_ ;
	wire _w15893_ ;
	wire _w15892_ ;
	wire _w15891_ ;
	wire _w15890_ ;
	wire _w15889_ ;
	wire _w15888_ ;
	wire _w15887_ ;
	wire _w15886_ ;
	wire _w15885_ ;
	wire _w15884_ ;
	wire _w15883_ ;
	wire _w15882_ ;
	wire _w15881_ ;
	wire _w15880_ ;
	wire _w15879_ ;
	wire _w15878_ ;
	wire _w15877_ ;
	wire _w15876_ ;
	wire _w15875_ ;
	wire _w15874_ ;
	wire _w15873_ ;
	wire _w15872_ ;
	wire _w15871_ ;
	wire _w15870_ ;
	wire _w15869_ ;
	wire _w15868_ ;
	wire _w15867_ ;
	wire _w15866_ ;
	wire _w15865_ ;
	wire _w15864_ ;
	wire _w15863_ ;
	wire _w15862_ ;
	wire _w15861_ ;
	wire _w15860_ ;
	wire _w15859_ ;
	wire _w15858_ ;
	wire _w15857_ ;
	wire _w15856_ ;
	wire _w15855_ ;
	wire _w15854_ ;
	wire _w15853_ ;
	wire _w15852_ ;
	wire _w15851_ ;
	wire _w15850_ ;
	wire _w15849_ ;
	wire _w15848_ ;
	wire _w15847_ ;
	wire _w15846_ ;
	wire _w15845_ ;
	wire _w15844_ ;
	wire _w15843_ ;
	wire _w15842_ ;
	wire _w15841_ ;
	wire _w15840_ ;
	wire _w15839_ ;
	wire _w15838_ ;
	wire _w15837_ ;
	wire _w15836_ ;
	wire _w15835_ ;
	wire _w15834_ ;
	wire _w15833_ ;
	wire _w15832_ ;
	wire _w15831_ ;
	wire _w15830_ ;
	wire _w15829_ ;
	wire _w15828_ ;
	wire _w15827_ ;
	wire _w15826_ ;
	wire _w15825_ ;
	wire _w15824_ ;
	wire _w15823_ ;
	wire _w15822_ ;
	wire _w15821_ ;
	wire _w15820_ ;
	wire _w15819_ ;
	wire _w15818_ ;
	wire _w15817_ ;
	wire _w15816_ ;
	wire _w15815_ ;
	wire _w15814_ ;
	wire _w15813_ ;
	wire _w15812_ ;
	wire _w15811_ ;
	wire _w15810_ ;
	wire _w15809_ ;
	wire _w15808_ ;
	wire _w15807_ ;
	wire _w15806_ ;
	wire _w15805_ ;
	wire _w15804_ ;
	wire _w15803_ ;
	wire _w15802_ ;
	wire _w15801_ ;
	wire _w15800_ ;
	wire _w15799_ ;
	wire _w15798_ ;
	wire _w15797_ ;
	wire _w15796_ ;
	wire _w15795_ ;
	wire _w15794_ ;
	wire _w15793_ ;
	wire _w15792_ ;
	wire _w15791_ ;
	wire _w15790_ ;
	wire _w15789_ ;
	wire _w15788_ ;
	wire _w15787_ ;
	wire _w15786_ ;
	wire _w15785_ ;
	wire _w15784_ ;
	wire _w15783_ ;
	wire _w15782_ ;
	wire _w15781_ ;
	wire _w15780_ ;
	wire _w15779_ ;
	wire _w15778_ ;
	wire _w15777_ ;
	wire _w15776_ ;
	wire _w15775_ ;
	wire _w15774_ ;
	wire _w15773_ ;
	wire _w15772_ ;
	wire _w15771_ ;
	wire _w15770_ ;
	wire _w15769_ ;
	wire _w15768_ ;
	wire _w15767_ ;
	wire _w15766_ ;
	wire _w15765_ ;
	wire _w15764_ ;
	wire _w15763_ ;
	wire _w15762_ ;
	wire _w15761_ ;
	wire _w15760_ ;
	wire _w15759_ ;
	wire _w15758_ ;
	wire _w15757_ ;
	wire _w15756_ ;
	wire _w15755_ ;
	wire _w15754_ ;
	wire _w15753_ ;
	wire _w15752_ ;
	wire _w15751_ ;
	wire _w15750_ ;
	wire _w15749_ ;
	wire _w15748_ ;
	wire _w15747_ ;
	wire _w15746_ ;
	wire _w15745_ ;
	wire _w15744_ ;
	wire _w15743_ ;
	wire _w15742_ ;
	wire _w15741_ ;
	wire _w15740_ ;
	wire _w15739_ ;
	wire _w15738_ ;
	wire _w15737_ ;
	wire _w15736_ ;
	wire _w15735_ ;
	wire _w15734_ ;
	wire _w15733_ ;
	wire _w15732_ ;
	wire _w15731_ ;
	wire _w15730_ ;
	wire _w15729_ ;
	wire _w15728_ ;
	wire _w15727_ ;
	wire _w15726_ ;
	wire _w15725_ ;
	wire _w15724_ ;
	wire _w15723_ ;
	wire _w15722_ ;
	wire _w15721_ ;
	wire _w15720_ ;
	wire _w15719_ ;
	wire _w15718_ ;
	wire _w15717_ ;
	wire _w15716_ ;
	wire _w15715_ ;
	wire _w15714_ ;
	wire _w15713_ ;
	wire _w15712_ ;
	wire _w15711_ ;
	wire _w15710_ ;
	wire _w15709_ ;
	wire _w15708_ ;
	wire _w15707_ ;
	wire _w15706_ ;
	wire _w15705_ ;
	wire _w15704_ ;
	wire _w15703_ ;
	wire _w15702_ ;
	wire _w15701_ ;
	wire _w15700_ ;
	wire _w15699_ ;
	wire _w15698_ ;
	wire _w15697_ ;
	wire _w15696_ ;
	wire _w15695_ ;
	wire _w15694_ ;
	wire _w15693_ ;
	wire _w15692_ ;
	wire _w15691_ ;
	wire _w15690_ ;
	wire _w15689_ ;
	wire _w15688_ ;
	wire _w15687_ ;
	wire _w15686_ ;
	wire _w15685_ ;
	wire _w15684_ ;
	wire _w15683_ ;
	wire _w15682_ ;
	wire _w15681_ ;
	wire _w15680_ ;
	wire _w15679_ ;
	wire _w15678_ ;
	wire _w15677_ ;
	wire _w15676_ ;
	wire _w15675_ ;
	wire _w15674_ ;
	wire _w15673_ ;
	wire _w15672_ ;
	wire _w15671_ ;
	wire _w15670_ ;
	wire _w15669_ ;
	wire _w15668_ ;
	wire _w15667_ ;
	wire _w15666_ ;
	wire _w15665_ ;
	wire _w15664_ ;
	wire _w15663_ ;
	wire _w15662_ ;
	wire _w15661_ ;
	wire _w15660_ ;
	wire _w15659_ ;
	wire _w15658_ ;
	wire _w15657_ ;
	wire _w15656_ ;
	wire _w15655_ ;
	wire _w15654_ ;
	wire _w15653_ ;
	wire _w15652_ ;
	wire _w15651_ ;
	wire _w15650_ ;
	wire _w15649_ ;
	wire _w15648_ ;
	wire _w15647_ ;
	wire _w15646_ ;
	wire _w15645_ ;
	wire _w15644_ ;
	wire _w15643_ ;
	wire _w15642_ ;
	wire _w15641_ ;
	wire _w15640_ ;
	wire _w15639_ ;
	wire _w15638_ ;
	wire _w15637_ ;
	wire _w15636_ ;
	wire _w15635_ ;
	wire _w15634_ ;
	wire _w15633_ ;
	wire _w15632_ ;
	wire _w15631_ ;
	wire _w15630_ ;
	wire _w15629_ ;
	wire _w15628_ ;
	wire _w15627_ ;
	wire _w15626_ ;
	wire _w15625_ ;
	wire _w15624_ ;
	wire _w15623_ ;
	wire _w15622_ ;
	wire _w15621_ ;
	wire _w15620_ ;
	wire _w15619_ ;
	wire _w15618_ ;
	wire _w15617_ ;
	wire _w15616_ ;
	wire _w15615_ ;
	wire _w15614_ ;
	wire _w15613_ ;
	wire _w15612_ ;
	wire _w15611_ ;
	wire _w15610_ ;
	wire _w15609_ ;
	wire _w15608_ ;
	wire _w15607_ ;
	wire _w15606_ ;
	wire _w15605_ ;
	wire _w15604_ ;
	wire _w15603_ ;
	wire _w15602_ ;
	wire _w15601_ ;
	wire _w15600_ ;
	wire _w15599_ ;
	wire _w15598_ ;
	wire _w15597_ ;
	wire _w15596_ ;
	wire _w15595_ ;
	wire _w15594_ ;
	wire _w15593_ ;
	wire _w15592_ ;
	wire _w15591_ ;
	wire _w15590_ ;
	wire _w15589_ ;
	wire _w15588_ ;
	wire _w15587_ ;
	wire _w15586_ ;
	wire _w15585_ ;
	wire _w15584_ ;
	wire _w15583_ ;
	wire _w15582_ ;
	wire _w15581_ ;
	wire _w15580_ ;
	wire _w15579_ ;
	wire _w15578_ ;
	wire _w15577_ ;
	wire _w15576_ ;
	wire _w15575_ ;
	wire _w15574_ ;
	wire _w15573_ ;
	wire _w15572_ ;
	wire _w15571_ ;
	wire _w15570_ ;
	wire _w15569_ ;
	wire _w15568_ ;
	wire _w15567_ ;
	wire _w15566_ ;
	wire _w15565_ ;
	wire _w15564_ ;
	wire _w15563_ ;
	wire _w15562_ ;
	wire _w15561_ ;
	wire _w15560_ ;
	wire _w15559_ ;
	wire _w15558_ ;
	wire _w15557_ ;
	wire _w15556_ ;
	wire _w15555_ ;
	wire _w15554_ ;
	wire _w15553_ ;
	wire _w15552_ ;
	wire _w15551_ ;
	wire _w15550_ ;
	wire _w15549_ ;
	wire _w15548_ ;
	wire _w15547_ ;
	wire _w15546_ ;
	wire _w15545_ ;
	wire _w15544_ ;
	wire _w15543_ ;
	wire _w15542_ ;
	wire _w15541_ ;
	wire _w15540_ ;
	wire _w15539_ ;
	wire _w15538_ ;
	wire _w15537_ ;
	wire _w15536_ ;
	wire _w15535_ ;
	wire _w15534_ ;
	wire _w15533_ ;
	wire _w15532_ ;
	wire _w15531_ ;
	wire _w15530_ ;
	wire _w15529_ ;
	wire _w15528_ ;
	wire _w15527_ ;
	wire _w15526_ ;
	wire _w15525_ ;
	wire _w15524_ ;
	wire _w15523_ ;
	wire _w15522_ ;
	wire _w15521_ ;
	wire _w15520_ ;
	wire _w15519_ ;
	wire _w15518_ ;
	wire _w15517_ ;
	wire _w15516_ ;
	wire _w15515_ ;
	wire _w15514_ ;
	wire _w15513_ ;
	wire _w15512_ ;
	wire _w15511_ ;
	wire _w15510_ ;
	wire _w15509_ ;
	wire _w15508_ ;
	wire _w15507_ ;
	wire _w15506_ ;
	wire _w15505_ ;
	wire _w15504_ ;
	wire _w15503_ ;
	wire _w15502_ ;
	wire _w15501_ ;
	wire _w15500_ ;
	wire _w15499_ ;
	wire _w15498_ ;
	wire _w15497_ ;
	wire _w15496_ ;
	wire _w15495_ ;
	wire _w15494_ ;
	wire _w15493_ ;
	wire _w15492_ ;
	wire _w15491_ ;
	wire _w15490_ ;
	wire _w15489_ ;
	wire _w15488_ ;
	wire _w15487_ ;
	wire _w15486_ ;
	wire _w15485_ ;
	wire _w15484_ ;
	wire _w15483_ ;
	wire _w15482_ ;
	wire _w15481_ ;
	wire _w15480_ ;
	wire _w15479_ ;
	wire _w15478_ ;
	wire _w15477_ ;
	wire _w15476_ ;
	wire _w15475_ ;
	wire _w15474_ ;
	wire _w15473_ ;
	wire _w15472_ ;
	wire _w15471_ ;
	wire _w15470_ ;
	wire _w15469_ ;
	wire _w15468_ ;
	wire _w15467_ ;
	wire _w15466_ ;
	wire _w15465_ ;
	wire _w15464_ ;
	wire _w15463_ ;
	wire _w15462_ ;
	wire _w15461_ ;
	wire _w15460_ ;
	wire _w15459_ ;
	wire _w15458_ ;
	wire _w15457_ ;
	wire _w15456_ ;
	wire _w15455_ ;
	wire _w15454_ ;
	wire _w15453_ ;
	wire _w15452_ ;
	wire _w15451_ ;
	wire _w15450_ ;
	wire _w15449_ ;
	wire _w15448_ ;
	wire _w15447_ ;
	wire _w15446_ ;
	wire _w15445_ ;
	wire _w15444_ ;
	wire _w15443_ ;
	wire _w15442_ ;
	wire _w15441_ ;
	wire _w15440_ ;
	wire _w15439_ ;
	wire _w15438_ ;
	wire _w15437_ ;
	wire _w15436_ ;
	wire _w15435_ ;
	wire _w15434_ ;
	wire _w15433_ ;
	wire _w15432_ ;
	wire _w15431_ ;
	wire _w15430_ ;
	wire _w15429_ ;
	wire _w15428_ ;
	wire _w15427_ ;
	wire _w15426_ ;
	wire _w15425_ ;
	wire _w15424_ ;
	wire _w15423_ ;
	wire _w15422_ ;
	wire _w15421_ ;
	wire _w15420_ ;
	wire _w15419_ ;
	wire _w15418_ ;
	wire _w15417_ ;
	wire _w15416_ ;
	wire _w15415_ ;
	wire _w15414_ ;
	wire _w15413_ ;
	wire _w15412_ ;
	wire _w15411_ ;
	wire _w15410_ ;
	wire _w15409_ ;
	wire _w15408_ ;
	wire _w15407_ ;
	wire _w15406_ ;
	wire _w15405_ ;
	wire _w15404_ ;
	wire _w15403_ ;
	wire _w15402_ ;
	wire _w15401_ ;
	wire _w15400_ ;
	wire _w15399_ ;
	wire _w15398_ ;
	wire _w15397_ ;
	wire _w15396_ ;
	wire _w15395_ ;
	wire _w15394_ ;
	wire _w15393_ ;
	wire _w15392_ ;
	wire _w15391_ ;
	wire _w15390_ ;
	wire _w15389_ ;
	wire _w15388_ ;
	wire _w15387_ ;
	wire _w15386_ ;
	wire _w15385_ ;
	wire _w15384_ ;
	wire _w15383_ ;
	wire _w15382_ ;
	wire _w15381_ ;
	wire _w15380_ ;
	wire _w15379_ ;
	wire _w15378_ ;
	wire _w15377_ ;
	wire _w15376_ ;
	wire _w15375_ ;
	wire _w15374_ ;
	wire _w15373_ ;
	wire _w15372_ ;
	wire _w15371_ ;
	wire _w15370_ ;
	wire _w15369_ ;
	wire _w15368_ ;
	wire _w15367_ ;
	wire _w15366_ ;
	wire _w15365_ ;
	wire _w15364_ ;
	wire _w15363_ ;
	wire _w15362_ ;
	wire _w15361_ ;
	wire _w15360_ ;
	wire _w15359_ ;
	wire _w15358_ ;
	wire _w15357_ ;
	wire _w15356_ ;
	wire _w15355_ ;
	wire _w15354_ ;
	wire _w15353_ ;
	wire _w15352_ ;
	wire _w15351_ ;
	wire _w15350_ ;
	wire _w15349_ ;
	wire _w15348_ ;
	wire _w15347_ ;
	wire _w15346_ ;
	wire _w15345_ ;
	wire _w15344_ ;
	wire _w15343_ ;
	wire _w15342_ ;
	wire _w15341_ ;
	wire _w15340_ ;
	wire _w15339_ ;
	wire _w15338_ ;
	wire _w15337_ ;
	wire _w15336_ ;
	wire _w15335_ ;
	wire _w15334_ ;
	wire _w15333_ ;
	wire _w15332_ ;
	wire _w15331_ ;
	wire _w15330_ ;
	wire _w15329_ ;
	wire _w15328_ ;
	wire _w15327_ ;
	wire _w15326_ ;
	wire _w15325_ ;
	wire _w15324_ ;
	wire _w15323_ ;
	wire _w15322_ ;
	wire _w15321_ ;
	wire _w15320_ ;
	wire _w15319_ ;
	wire _w15318_ ;
	wire _w15317_ ;
	wire _w15316_ ;
	wire _w15315_ ;
	wire _w15314_ ;
	wire _w15313_ ;
	wire _w15312_ ;
	wire _w15311_ ;
	wire _w15310_ ;
	wire _w15309_ ;
	wire _w15308_ ;
	wire _w15307_ ;
	wire _w15306_ ;
	wire _w15305_ ;
	wire _w15304_ ;
	wire _w15303_ ;
	wire _w15302_ ;
	wire _w15301_ ;
	wire _w15300_ ;
	wire _w15299_ ;
	wire _w15298_ ;
	wire _w15297_ ;
	wire _w15296_ ;
	wire _w15295_ ;
	wire _w15294_ ;
	wire _w15293_ ;
	wire _w15292_ ;
	wire _w15291_ ;
	wire _w15290_ ;
	wire _w15289_ ;
	wire _w15288_ ;
	wire _w15287_ ;
	wire _w15286_ ;
	wire _w15285_ ;
	wire _w15284_ ;
	wire _w15283_ ;
	wire _w15282_ ;
	wire _w15281_ ;
	wire _w15280_ ;
	wire _w15279_ ;
	wire _w15278_ ;
	wire _w15277_ ;
	wire _w15276_ ;
	wire _w15275_ ;
	wire _w15274_ ;
	wire _w15273_ ;
	wire _w15272_ ;
	wire _w15271_ ;
	wire _w15270_ ;
	wire _w15269_ ;
	wire _w15268_ ;
	wire _w15267_ ;
	wire _w15266_ ;
	wire _w15265_ ;
	wire _w15264_ ;
	wire _w15263_ ;
	wire _w15262_ ;
	wire _w15261_ ;
	wire _w15260_ ;
	wire _w15259_ ;
	wire _w15258_ ;
	wire _w15257_ ;
	wire _w15256_ ;
	wire _w15255_ ;
	wire _w15254_ ;
	wire _w15253_ ;
	wire _w15252_ ;
	wire _w15251_ ;
	wire _w15250_ ;
	wire _w15249_ ;
	wire _w15248_ ;
	wire _w15247_ ;
	wire _w15246_ ;
	wire _w15245_ ;
	wire _w15244_ ;
	wire _w15243_ ;
	wire _w15242_ ;
	wire _w15241_ ;
	wire _w15240_ ;
	wire _w15239_ ;
	wire _w15238_ ;
	wire _w15237_ ;
	wire _w15236_ ;
	wire _w15235_ ;
	wire _w15234_ ;
	wire _w15233_ ;
	wire _w15232_ ;
	wire _w15231_ ;
	wire _w15230_ ;
	wire _w15229_ ;
	wire _w15228_ ;
	wire _w15227_ ;
	wire _w15226_ ;
	wire _w15225_ ;
	wire _w15224_ ;
	wire _w15223_ ;
	wire _w15222_ ;
	wire _w15221_ ;
	wire _w15220_ ;
	wire _w15219_ ;
	wire _w15218_ ;
	wire _w15217_ ;
	wire _w15216_ ;
	wire _w15215_ ;
	wire _w15214_ ;
	wire _w15213_ ;
	wire _w15212_ ;
	wire _w15211_ ;
	wire _w15210_ ;
	wire _w15209_ ;
	wire _w15208_ ;
	wire _w15207_ ;
	wire _w15206_ ;
	wire _w15205_ ;
	wire _w15204_ ;
	wire _w15203_ ;
	wire _w15202_ ;
	wire _w15201_ ;
	wire _w15200_ ;
	wire _w15199_ ;
	wire _w15198_ ;
	wire _w15197_ ;
	wire _w15196_ ;
	wire _w15195_ ;
	wire _w15194_ ;
	wire _w15193_ ;
	wire _w15192_ ;
	wire _w15191_ ;
	wire _w15190_ ;
	wire _w15189_ ;
	wire _w15188_ ;
	wire _w15187_ ;
	wire _w15186_ ;
	wire _w15185_ ;
	wire _w15184_ ;
	wire _w15183_ ;
	wire _w15182_ ;
	wire _w15181_ ;
	wire _w15180_ ;
	wire _w15179_ ;
	wire _w15178_ ;
	wire _w15177_ ;
	wire _w15176_ ;
	wire _w15175_ ;
	wire _w15174_ ;
	wire _w15173_ ;
	wire _w15172_ ;
	wire _w15171_ ;
	wire _w15170_ ;
	wire _w15169_ ;
	wire _w15168_ ;
	wire _w15167_ ;
	wire _w15166_ ;
	wire _w15165_ ;
	wire _w15164_ ;
	wire _w15163_ ;
	wire _w15162_ ;
	wire _w15161_ ;
	wire _w15160_ ;
	wire _w15159_ ;
	wire _w15158_ ;
	wire _w15157_ ;
	wire _w15156_ ;
	wire _w15155_ ;
	wire _w15154_ ;
	wire _w15153_ ;
	wire _w15152_ ;
	wire _w15151_ ;
	wire _w15150_ ;
	wire _w15149_ ;
	wire _w15148_ ;
	wire _w15147_ ;
	wire _w15146_ ;
	wire _w15145_ ;
	wire _w15144_ ;
	wire _w15143_ ;
	wire _w15142_ ;
	wire _w15141_ ;
	wire _w15140_ ;
	wire _w15139_ ;
	wire _w15138_ ;
	wire _w15137_ ;
	wire _w15136_ ;
	wire _w15135_ ;
	wire _w15134_ ;
	wire _w15133_ ;
	wire _w15132_ ;
	wire _w15131_ ;
	wire _w15130_ ;
	wire _w15129_ ;
	wire _w15128_ ;
	wire _w15127_ ;
	wire _w15126_ ;
	wire _w15125_ ;
	wire _w15124_ ;
	wire _w15123_ ;
	wire _w15122_ ;
	wire _w15121_ ;
	wire _w15120_ ;
	wire _w15119_ ;
	wire _w15118_ ;
	wire _w15117_ ;
	wire _w15116_ ;
	wire _w15115_ ;
	wire _w15114_ ;
	wire _w15113_ ;
	wire _w15112_ ;
	wire _w15111_ ;
	wire _w15110_ ;
	wire _w15109_ ;
	wire _w15108_ ;
	wire _w15107_ ;
	wire _w15106_ ;
	wire _w15105_ ;
	wire _w15104_ ;
	wire _w15103_ ;
	wire _w15102_ ;
	wire _w15101_ ;
	wire _w15100_ ;
	wire _w15099_ ;
	wire _w15098_ ;
	wire _w15097_ ;
	wire _w15096_ ;
	wire _w15095_ ;
	wire _w15094_ ;
	wire _w15093_ ;
	wire _w15092_ ;
	wire _w15091_ ;
	wire _w15090_ ;
	wire _w15089_ ;
	wire _w15088_ ;
	wire _w15087_ ;
	wire _w15086_ ;
	wire _w15085_ ;
	wire _w15084_ ;
	wire _w15083_ ;
	wire _w15082_ ;
	wire _w15081_ ;
	wire _w15080_ ;
	wire _w15079_ ;
	wire _w15078_ ;
	wire _w15077_ ;
	wire _w15076_ ;
	wire _w15075_ ;
	wire _w15074_ ;
	wire _w15073_ ;
	wire _w15072_ ;
	wire _w15071_ ;
	wire _w15070_ ;
	wire _w15069_ ;
	wire _w15068_ ;
	wire _w15067_ ;
	wire _w15066_ ;
	wire _w15065_ ;
	wire _w15064_ ;
	wire _w15063_ ;
	wire _w15062_ ;
	wire _w15061_ ;
	wire _w15060_ ;
	wire _w15059_ ;
	wire _w15058_ ;
	wire _w15057_ ;
	wire _w15056_ ;
	wire _w15055_ ;
	wire _w15054_ ;
	wire _w15053_ ;
	wire _w15052_ ;
	wire _w15051_ ;
	wire _w15050_ ;
	wire _w15049_ ;
	wire _w15048_ ;
	wire _w15047_ ;
	wire _w15046_ ;
	wire _w15045_ ;
	wire _w15044_ ;
	wire _w15043_ ;
	wire _w15042_ ;
	wire _w15041_ ;
	wire _w15040_ ;
	wire _w15039_ ;
	wire _w15038_ ;
	wire _w15037_ ;
	wire _w15036_ ;
	wire _w15035_ ;
	wire _w15034_ ;
	wire _w15033_ ;
	wire _w15032_ ;
	wire _w15031_ ;
	wire _w15030_ ;
	wire _w15029_ ;
	wire _w15028_ ;
	wire _w15027_ ;
	wire _w15026_ ;
	wire _w15025_ ;
	wire _w15024_ ;
	wire _w15023_ ;
	wire _w15022_ ;
	wire _w15021_ ;
	wire _w15020_ ;
	wire _w15019_ ;
	wire _w15018_ ;
	wire _w15017_ ;
	wire _w15016_ ;
	wire _w15015_ ;
	wire _w15014_ ;
	wire _w15013_ ;
	wire _w15012_ ;
	wire _w15011_ ;
	wire _w15010_ ;
	wire _w15009_ ;
	wire _w15008_ ;
	wire _w15007_ ;
	wire _w15006_ ;
	wire _w15005_ ;
	wire _w15004_ ;
	wire _w15003_ ;
	wire _w15002_ ;
	wire _w15001_ ;
	wire _w15000_ ;
	wire _w14999_ ;
	wire _w14998_ ;
	wire _w14997_ ;
	wire _w14996_ ;
	wire _w14995_ ;
	wire _w14994_ ;
	wire _w14993_ ;
	wire _w14992_ ;
	wire _w14991_ ;
	wire _w14990_ ;
	wire _w14989_ ;
	wire _w14988_ ;
	wire _w14987_ ;
	wire _w14986_ ;
	wire _w14985_ ;
	wire _w14984_ ;
	wire _w14983_ ;
	wire _w14982_ ;
	wire _w14981_ ;
	wire _w14980_ ;
	wire _w14979_ ;
	wire _w14978_ ;
	wire _w14977_ ;
	wire _w14976_ ;
	wire _w14975_ ;
	wire _w14974_ ;
	wire _w14973_ ;
	wire _w14972_ ;
	wire _w14971_ ;
	wire _w14970_ ;
	wire _w14969_ ;
	wire _w14968_ ;
	wire _w14967_ ;
	wire _w14966_ ;
	wire _w14965_ ;
	wire _w14964_ ;
	wire _w14963_ ;
	wire _w14962_ ;
	wire _w14961_ ;
	wire _w14960_ ;
	wire _w14959_ ;
	wire _w14958_ ;
	wire _w14957_ ;
	wire _w14956_ ;
	wire _w14955_ ;
	wire _w14954_ ;
	wire _w14953_ ;
	wire _w14952_ ;
	wire _w14951_ ;
	wire _w14950_ ;
	wire _w14949_ ;
	wire _w14948_ ;
	wire _w14947_ ;
	wire _w14946_ ;
	wire _w14945_ ;
	wire _w14944_ ;
	wire _w14943_ ;
	wire _w14942_ ;
	wire _w14941_ ;
	wire _w14940_ ;
	wire _w14939_ ;
	wire _w14938_ ;
	wire _w14937_ ;
	wire _w14936_ ;
	wire _w14935_ ;
	wire _w14934_ ;
	wire _w14933_ ;
	wire _w14932_ ;
	wire _w14931_ ;
	wire _w14930_ ;
	wire _w14929_ ;
	wire _w14928_ ;
	wire _w14927_ ;
	wire _w14926_ ;
	wire _w14925_ ;
	wire _w14924_ ;
	wire _w14923_ ;
	wire _w14922_ ;
	wire _w14921_ ;
	wire _w14920_ ;
	wire _w14919_ ;
	wire _w14918_ ;
	wire _w14917_ ;
	wire _w14916_ ;
	wire _w14915_ ;
	wire _w14914_ ;
	wire _w14913_ ;
	wire _w14912_ ;
	wire _w14911_ ;
	wire _w14910_ ;
	wire _w14909_ ;
	wire _w14908_ ;
	wire _w14907_ ;
	wire _w14906_ ;
	wire _w14905_ ;
	wire _w14904_ ;
	wire _w14903_ ;
	wire _w14902_ ;
	wire _w14901_ ;
	wire _w14900_ ;
	wire _w14899_ ;
	wire _w14898_ ;
	wire _w14897_ ;
	wire _w14896_ ;
	wire _w14895_ ;
	wire _w14894_ ;
	wire _w14893_ ;
	wire _w14892_ ;
	wire _w14891_ ;
	wire _w14890_ ;
	wire _w14889_ ;
	wire _w14888_ ;
	wire _w14887_ ;
	wire _w14886_ ;
	wire _w14885_ ;
	wire _w14884_ ;
	wire _w14883_ ;
	wire _w14882_ ;
	wire _w14881_ ;
	wire _w14880_ ;
	wire _w14879_ ;
	wire _w14878_ ;
	wire _w14877_ ;
	wire _w14876_ ;
	wire _w14875_ ;
	wire _w14874_ ;
	wire _w14873_ ;
	wire _w14872_ ;
	wire _w14871_ ;
	wire _w14870_ ;
	wire _w14869_ ;
	wire _w14868_ ;
	wire _w14867_ ;
	wire _w14866_ ;
	wire _w14865_ ;
	wire _w14864_ ;
	wire _w14863_ ;
	wire _w14862_ ;
	wire _w14861_ ;
	wire _w14860_ ;
	wire _w14859_ ;
	wire _w14858_ ;
	wire _w14857_ ;
	wire _w14856_ ;
	wire _w14855_ ;
	wire _w14854_ ;
	wire _w14853_ ;
	wire _w14852_ ;
	wire _w14851_ ;
	wire _w14850_ ;
	wire _w14849_ ;
	wire _w14848_ ;
	wire _w14847_ ;
	wire _w14846_ ;
	wire _w14845_ ;
	wire _w14844_ ;
	wire _w14843_ ;
	wire _w14842_ ;
	wire _w14841_ ;
	wire _w14840_ ;
	wire _w14839_ ;
	wire _w14838_ ;
	wire _w14837_ ;
	wire _w14836_ ;
	wire _w14835_ ;
	wire _w14834_ ;
	wire _w14833_ ;
	wire _w14832_ ;
	wire _w14831_ ;
	wire _w14830_ ;
	wire _w14829_ ;
	wire _w14828_ ;
	wire _w14827_ ;
	wire _w14826_ ;
	wire _w14825_ ;
	wire _w14824_ ;
	wire _w14823_ ;
	wire _w14822_ ;
	wire _w14821_ ;
	wire _w14820_ ;
	wire _w14819_ ;
	wire _w14818_ ;
	wire _w14817_ ;
	wire _w14816_ ;
	wire _w14815_ ;
	wire _w14814_ ;
	wire _w14813_ ;
	wire _w14812_ ;
	wire _w14811_ ;
	wire _w14810_ ;
	wire _w14809_ ;
	wire _w14808_ ;
	wire _w14807_ ;
	wire _w14806_ ;
	wire _w14805_ ;
	wire _w14804_ ;
	wire _w14803_ ;
	wire _w14802_ ;
	wire _w14801_ ;
	wire _w14800_ ;
	wire _w14799_ ;
	wire _w14798_ ;
	wire _w14797_ ;
	wire _w14796_ ;
	wire _w14795_ ;
	wire _w14794_ ;
	wire _w14793_ ;
	wire _w14792_ ;
	wire _w14791_ ;
	wire _w14790_ ;
	wire _w14789_ ;
	wire _w14788_ ;
	wire _w14787_ ;
	wire _w14786_ ;
	wire _w14785_ ;
	wire _w14784_ ;
	wire _w14783_ ;
	wire _w14782_ ;
	wire _w14781_ ;
	wire _w14780_ ;
	wire _w14779_ ;
	wire _w14778_ ;
	wire _w14777_ ;
	wire _w14776_ ;
	wire _w14775_ ;
	wire _w14774_ ;
	wire _w14773_ ;
	wire _w14772_ ;
	wire _w14771_ ;
	wire _w14770_ ;
	wire _w14769_ ;
	wire _w14768_ ;
	wire _w14767_ ;
	wire _w14766_ ;
	wire _w14765_ ;
	wire _w14764_ ;
	wire _w14763_ ;
	wire _w14762_ ;
	wire _w14761_ ;
	wire _w14760_ ;
	wire _w14759_ ;
	wire _w14758_ ;
	wire _w14757_ ;
	wire _w14756_ ;
	wire _w14755_ ;
	wire _w14754_ ;
	wire _w14753_ ;
	wire _w14752_ ;
	wire _w14751_ ;
	wire _w14750_ ;
	wire _w14749_ ;
	wire _w14748_ ;
	wire _w14747_ ;
	wire _w14746_ ;
	wire _w14745_ ;
	wire _w14744_ ;
	wire _w14743_ ;
	wire _w14742_ ;
	wire _w14741_ ;
	wire _w14740_ ;
	wire _w14739_ ;
	wire _w14738_ ;
	wire _w14737_ ;
	wire _w14736_ ;
	wire _w14735_ ;
	wire _w14734_ ;
	wire _w14733_ ;
	wire _w14732_ ;
	wire _w14731_ ;
	wire _w14730_ ;
	wire _w14729_ ;
	wire _w14728_ ;
	wire _w14727_ ;
	wire _w14726_ ;
	wire _w14725_ ;
	wire _w14724_ ;
	wire _w14723_ ;
	wire _w14722_ ;
	wire _w14721_ ;
	wire _w14720_ ;
	wire _w14719_ ;
	wire _w14718_ ;
	wire _w14717_ ;
	wire _w14716_ ;
	wire _w14715_ ;
	wire _w14714_ ;
	wire _w14713_ ;
	wire _w14712_ ;
	wire _w14711_ ;
	wire _w14710_ ;
	wire _w14709_ ;
	wire _w14708_ ;
	wire _w14707_ ;
	wire _w14706_ ;
	wire _w14705_ ;
	wire _w14704_ ;
	wire _w14703_ ;
	wire _w14702_ ;
	wire _w14701_ ;
	wire _w14700_ ;
	wire _w14699_ ;
	wire _w14698_ ;
	wire _w14697_ ;
	wire _w14696_ ;
	wire _w14695_ ;
	wire _w14694_ ;
	wire _w14693_ ;
	wire _w14692_ ;
	wire _w14691_ ;
	wire _w14690_ ;
	wire _w14689_ ;
	wire _w14688_ ;
	wire _w14687_ ;
	wire _w14686_ ;
	wire _w14685_ ;
	wire _w14684_ ;
	wire _w14683_ ;
	wire _w14682_ ;
	wire _w14681_ ;
	wire _w14680_ ;
	wire _w14679_ ;
	wire _w14678_ ;
	wire _w14677_ ;
	wire _w14676_ ;
	wire _w14675_ ;
	wire _w14674_ ;
	wire _w14673_ ;
	wire _w14672_ ;
	wire _w14671_ ;
	wire _w14670_ ;
	wire _w14669_ ;
	wire _w14668_ ;
	wire _w14667_ ;
	wire _w14666_ ;
	wire _w14665_ ;
	wire _w14664_ ;
	wire _w14663_ ;
	wire _w14662_ ;
	wire _w14661_ ;
	wire _w14660_ ;
	wire _w14659_ ;
	wire _w14658_ ;
	wire _w14657_ ;
	wire _w14656_ ;
	wire _w14655_ ;
	wire _w14654_ ;
	wire _w14653_ ;
	wire _w14652_ ;
	wire _w14651_ ;
	wire _w14650_ ;
	wire _w14649_ ;
	wire _w14648_ ;
	wire _w14647_ ;
	wire _w14646_ ;
	wire _w14645_ ;
	wire _w14644_ ;
	wire _w14643_ ;
	wire _w14642_ ;
	wire _w14641_ ;
	wire _w14640_ ;
	wire _w14639_ ;
	wire _w14638_ ;
	wire _w14637_ ;
	wire _w14636_ ;
	wire _w14635_ ;
	wire _w14634_ ;
	wire _w14633_ ;
	wire _w14632_ ;
	wire _w14631_ ;
	wire _w14630_ ;
	wire _w14629_ ;
	wire _w14628_ ;
	wire _w14627_ ;
	wire _w14626_ ;
	wire _w14625_ ;
	wire _w14624_ ;
	wire _w14623_ ;
	wire _w14622_ ;
	wire _w14621_ ;
	wire _w14620_ ;
	wire _w14619_ ;
	wire _w14618_ ;
	wire _w14617_ ;
	wire _w14616_ ;
	wire _w14615_ ;
	wire _w14614_ ;
	wire _w14613_ ;
	wire _w14612_ ;
	wire _w14611_ ;
	wire _w14610_ ;
	wire _w14609_ ;
	wire _w14608_ ;
	wire _w14607_ ;
	wire _w14606_ ;
	wire _w14605_ ;
	wire _w14604_ ;
	wire _w14603_ ;
	wire _w14602_ ;
	wire _w14601_ ;
	wire _w14600_ ;
	wire _w14599_ ;
	wire _w14598_ ;
	wire _w14597_ ;
	wire _w14596_ ;
	wire _w14595_ ;
	wire _w14594_ ;
	wire _w14593_ ;
	wire _w14592_ ;
	wire _w14591_ ;
	wire _w14590_ ;
	wire _w14589_ ;
	wire _w14588_ ;
	wire _w14587_ ;
	wire _w14586_ ;
	wire _w14585_ ;
	wire _w14584_ ;
	wire _w14583_ ;
	wire _w14582_ ;
	wire _w14581_ ;
	wire _w14580_ ;
	wire _w14579_ ;
	wire _w14578_ ;
	wire _w14577_ ;
	wire _w14576_ ;
	wire _w14575_ ;
	wire _w14574_ ;
	wire _w14573_ ;
	wire _w14572_ ;
	wire _w14571_ ;
	wire _w14570_ ;
	wire _w14569_ ;
	wire _w14568_ ;
	wire _w14567_ ;
	wire _w14566_ ;
	wire _w14565_ ;
	wire _w14564_ ;
	wire _w14563_ ;
	wire _w14562_ ;
	wire _w14561_ ;
	wire _w14560_ ;
	wire _w14559_ ;
	wire _w14558_ ;
	wire _w14557_ ;
	wire _w14556_ ;
	wire _w14555_ ;
	wire _w14554_ ;
	wire _w14553_ ;
	wire _w14552_ ;
	wire _w14551_ ;
	wire _w14550_ ;
	wire _w14549_ ;
	wire _w14548_ ;
	wire _w14547_ ;
	wire _w14546_ ;
	wire _w14545_ ;
	wire _w14544_ ;
	wire _w14543_ ;
	wire _w14542_ ;
	wire _w14541_ ;
	wire _w14540_ ;
	wire _w14539_ ;
	wire _w14538_ ;
	wire _w14537_ ;
	wire _w14536_ ;
	wire _w14535_ ;
	wire _w14534_ ;
	wire _w14533_ ;
	wire _w14532_ ;
	wire _w14531_ ;
	wire _w14530_ ;
	wire _w14529_ ;
	wire _w14528_ ;
	wire _w14527_ ;
	wire _w14526_ ;
	wire _w14525_ ;
	wire _w14524_ ;
	wire _w14523_ ;
	wire _w14522_ ;
	wire _w14521_ ;
	wire _w14520_ ;
	wire _w14519_ ;
	wire _w14518_ ;
	wire _w14517_ ;
	wire _w14516_ ;
	wire _w14515_ ;
	wire _w14514_ ;
	wire _w14513_ ;
	wire _w14512_ ;
	wire _w14511_ ;
	wire _w14510_ ;
	wire _w14509_ ;
	wire _w14508_ ;
	wire _w14507_ ;
	wire _w14506_ ;
	wire _w14505_ ;
	wire _w14504_ ;
	wire _w14503_ ;
	wire _w14502_ ;
	wire _w14501_ ;
	wire _w14500_ ;
	wire _w14499_ ;
	wire _w14498_ ;
	wire _w14497_ ;
	wire _w14496_ ;
	wire _w14495_ ;
	wire _w14494_ ;
	wire _w14493_ ;
	wire _w14492_ ;
	wire _w14491_ ;
	wire _w14490_ ;
	wire _w14489_ ;
	wire _w14488_ ;
	wire _w14487_ ;
	wire _w14486_ ;
	wire _w14485_ ;
	wire _w14484_ ;
	wire _w14483_ ;
	wire _w14482_ ;
	wire _w14481_ ;
	wire _w14480_ ;
	wire _w14479_ ;
	wire _w14478_ ;
	wire _w14477_ ;
	wire _w14476_ ;
	wire _w14475_ ;
	wire _w14474_ ;
	wire _w14473_ ;
	wire _w14472_ ;
	wire _w14471_ ;
	wire _w14470_ ;
	wire _w14469_ ;
	wire _w14468_ ;
	wire _w14467_ ;
	wire _w14466_ ;
	wire _w14465_ ;
	wire _w14464_ ;
	wire _w14463_ ;
	wire _w14462_ ;
	wire _w14461_ ;
	wire _w14460_ ;
	wire _w14459_ ;
	wire _w14458_ ;
	wire _w14457_ ;
	wire _w14456_ ;
	wire _w14455_ ;
	wire _w14454_ ;
	wire _w14453_ ;
	wire _w14452_ ;
	wire _w14451_ ;
	wire _w14450_ ;
	wire _w14449_ ;
	wire _w14448_ ;
	wire _w14447_ ;
	wire _w14446_ ;
	wire _w14445_ ;
	wire _w14444_ ;
	wire _w14443_ ;
	wire _w14442_ ;
	wire _w14441_ ;
	wire _w14440_ ;
	wire _w14439_ ;
	wire _w14438_ ;
	wire _w14437_ ;
	wire _w14436_ ;
	wire _w14435_ ;
	wire _w14434_ ;
	wire _w14433_ ;
	wire _w14432_ ;
	wire _w14431_ ;
	wire _w14430_ ;
	wire _w14429_ ;
	wire _w14428_ ;
	wire _w14427_ ;
	wire _w14426_ ;
	wire _w14425_ ;
	wire _w14424_ ;
	wire _w14423_ ;
	wire _w14422_ ;
	wire _w14421_ ;
	wire _w14420_ ;
	wire _w14419_ ;
	wire _w14418_ ;
	wire _w14417_ ;
	wire _w14416_ ;
	wire _w14415_ ;
	wire _w14414_ ;
	wire _w14413_ ;
	wire _w14412_ ;
	wire _w14411_ ;
	wire _w14410_ ;
	wire _w14409_ ;
	wire _w14408_ ;
	wire _w14407_ ;
	wire _w14406_ ;
	wire _w14405_ ;
	wire _w14404_ ;
	wire _w14403_ ;
	wire _w14402_ ;
	wire _w14401_ ;
	wire _w14400_ ;
	wire _w14399_ ;
	wire _w14398_ ;
	wire _w14397_ ;
	wire _w14396_ ;
	wire _w14395_ ;
	wire _w14394_ ;
	wire _w14393_ ;
	wire _w14392_ ;
	wire _w14391_ ;
	wire _w14390_ ;
	wire _w14389_ ;
	wire _w14388_ ;
	wire _w14387_ ;
	wire _w14386_ ;
	wire _w14385_ ;
	wire _w14384_ ;
	wire _w14383_ ;
	wire _w14382_ ;
	wire _w14381_ ;
	wire _w14380_ ;
	wire _w14379_ ;
	wire _w14378_ ;
	wire _w14377_ ;
	wire _w14376_ ;
	wire _w14375_ ;
	wire _w14374_ ;
	wire _w14373_ ;
	wire _w14372_ ;
	wire _w14371_ ;
	wire _w14370_ ;
	wire _w14369_ ;
	wire _w14368_ ;
	wire _w14367_ ;
	wire _w14366_ ;
	wire _w14365_ ;
	wire _w14364_ ;
	wire _w14363_ ;
	wire _w14362_ ;
	wire _w14361_ ;
	wire _w14360_ ;
	wire _w14359_ ;
	wire _w14358_ ;
	wire _w14357_ ;
	wire _w14356_ ;
	wire _w14355_ ;
	wire _w14354_ ;
	wire _w14353_ ;
	wire _w14352_ ;
	wire _w14351_ ;
	wire _w14350_ ;
	wire _w14349_ ;
	wire _w14348_ ;
	wire _w14347_ ;
	wire _w14346_ ;
	wire _w14345_ ;
	wire _w14344_ ;
	wire _w14343_ ;
	wire _w14342_ ;
	wire _w14341_ ;
	wire _w14340_ ;
	wire _w14339_ ;
	wire _w14338_ ;
	wire _w14337_ ;
	wire _w14336_ ;
	wire _w14335_ ;
	wire _w14334_ ;
	wire _w14333_ ;
	wire _w14332_ ;
	wire _w14331_ ;
	wire _w14330_ ;
	wire _w14329_ ;
	wire _w14328_ ;
	wire _w14327_ ;
	wire _w14326_ ;
	wire _w14325_ ;
	wire _w14324_ ;
	wire _w14323_ ;
	wire _w14322_ ;
	wire _w14321_ ;
	wire _w14320_ ;
	wire _w14319_ ;
	wire _w14318_ ;
	wire _w14317_ ;
	wire _w14316_ ;
	wire _w14315_ ;
	wire _w14314_ ;
	wire _w14313_ ;
	wire _w14312_ ;
	wire _w14311_ ;
	wire _w14310_ ;
	wire _w14309_ ;
	wire _w14308_ ;
	wire _w14307_ ;
	wire _w14306_ ;
	wire _w14305_ ;
	wire _w14304_ ;
	wire _w14303_ ;
	wire _w14302_ ;
	wire _w14301_ ;
	wire _w14300_ ;
	wire _w14299_ ;
	wire _w14298_ ;
	wire _w14297_ ;
	wire _w14296_ ;
	wire _w14295_ ;
	wire _w14294_ ;
	wire _w14293_ ;
	wire _w14292_ ;
	wire _w14291_ ;
	wire _w14290_ ;
	wire _w14289_ ;
	wire _w14288_ ;
	wire _w14287_ ;
	wire _w14286_ ;
	wire _w14285_ ;
	wire _w14284_ ;
	wire _w14283_ ;
	wire _w14282_ ;
	wire _w14281_ ;
	wire _w14280_ ;
	wire _w14279_ ;
	wire _w14278_ ;
	wire _w14277_ ;
	wire _w14276_ ;
	wire _w14275_ ;
	wire _w14274_ ;
	wire _w14273_ ;
	wire _w14272_ ;
	wire _w14271_ ;
	wire _w14270_ ;
	wire _w14269_ ;
	wire _w14268_ ;
	wire _w14267_ ;
	wire _w14266_ ;
	wire _w14265_ ;
	wire _w14264_ ;
	wire _w14263_ ;
	wire _w14262_ ;
	wire _w14261_ ;
	wire _w14260_ ;
	wire _w14259_ ;
	wire _w14258_ ;
	wire _w14257_ ;
	wire _w14256_ ;
	wire _w14255_ ;
	wire _w14254_ ;
	wire _w14253_ ;
	wire _w14252_ ;
	wire _w14251_ ;
	wire _w14250_ ;
	wire _w14249_ ;
	wire _w14248_ ;
	wire _w14247_ ;
	wire _w14246_ ;
	wire _w14245_ ;
	wire _w14244_ ;
	wire _w14243_ ;
	wire _w14242_ ;
	wire _w14241_ ;
	wire _w14240_ ;
	wire _w14239_ ;
	wire _w14238_ ;
	wire _w14237_ ;
	wire _w14236_ ;
	wire _w14235_ ;
	wire _w14234_ ;
	wire _w14233_ ;
	wire _w14232_ ;
	wire _w14231_ ;
	wire _w14230_ ;
	wire _w14229_ ;
	wire _w14228_ ;
	wire _w14227_ ;
	wire _w14226_ ;
	wire _w14225_ ;
	wire _w14224_ ;
	wire _w14223_ ;
	wire _w14222_ ;
	wire _w14221_ ;
	wire _w14220_ ;
	wire _w14219_ ;
	wire _w14218_ ;
	wire _w14217_ ;
	wire _w14216_ ;
	wire _w14215_ ;
	wire _w14214_ ;
	wire _w14213_ ;
	wire _w14212_ ;
	wire _w14211_ ;
	wire _w14210_ ;
	wire _w14209_ ;
	wire _w14208_ ;
	wire _w14207_ ;
	wire _w14206_ ;
	wire _w14205_ ;
	wire _w14204_ ;
	wire _w14203_ ;
	wire _w14202_ ;
	wire _w14201_ ;
	wire _w14200_ ;
	wire _w14199_ ;
	wire _w14198_ ;
	wire _w14197_ ;
	wire _w14196_ ;
	wire _w14195_ ;
	wire _w14194_ ;
	wire _w14193_ ;
	wire _w14192_ ;
	wire _w14191_ ;
	wire _w14190_ ;
	wire _w14189_ ;
	wire _w14188_ ;
	wire _w14187_ ;
	wire _w14186_ ;
	wire _w14185_ ;
	wire _w14184_ ;
	wire _w14183_ ;
	wire _w14182_ ;
	wire _w14181_ ;
	wire _w14180_ ;
	wire _w14179_ ;
	wire _w14178_ ;
	wire _w14177_ ;
	wire _w14176_ ;
	wire _w14175_ ;
	wire _w14174_ ;
	wire _w14173_ ;
	wire _w14172_ ;
	wire _w14171_ ;
	wire _w14170_ ;
	wire _w14169_ ;
	wire _w14168_ ;
	wire _w14167_ ;
	wire _w14166_ ;
	wire _w14165_ ;
	wire _w14164_ ;
	wire _w14163_ ;
	wire _w14162_ ;
	wire _w14161_ ;
	wire _w14160_ ;
	wire _w14159_ ;
	wire _w14158_ ;
	wire _w14157_ ;
	wire _w14156_ ;
	wire _w14155_ ;
	wire _w14154_ ;
	wire _w14153_ ;
	wire _w14152_ ;
	wire _w14151_ ;
	wire _w14150_ ;
	wire _w14149_ ;
	wire _w14148_ ;
	wire _w14147_ ;
	wire _w14146_ ;
	wire _w14145_ ;
	wire _w14144_ ;
	wire _w14143_ ;
	wire _w14142_ ;
	wire _w14141_ ;
	wire _w14140_ ;
	wire _w14139_ ;
	wire _w14138_ ;
	wire _w14137_ ;
	wire _w14136_ ;
	wire _w14135_ ;
	wire _w14134_ ;
	wire _w14133_ ;
	wire _w14132_ ;
	wire _w14131_ ;
	wire _w14130_ ;
	wire _w14129_ ;
	wire _w14128_ ;
	wire _w14127_ ;
	wire _w14126_ ;
	wire _w14125_ ;
	wire _w14124_ ;
	wire _w14123_ ;
	wire _w14122_ ;
	wire _w14121_ ;
	wire _w14120_ ;
	wire _w14119_ ;
	wire _w14118_ ;
	wire _w14117_ ;
	wire _w14116_ ;
	wire _w14115_ ;
	wire _w14114_ ;
	wire _w14113_ ;
	wire _w14112_ ;
	wire _w14111_ ;
	wire _w14110_ ;
	wire _w14109_ ;
	wire _w14108_ ;
	wire _w14107_ ;
	wire _w14106_ ;
	wire _w14105_ ;
	wire _w14104_ ;
	wire _w14103_ ;
	wire _w14102_ ;
	wire _w14101_ ;
	wire _w14100_ ;
	wire _w14099_ ;
	wire _w14098_ ;
	wire _w14097_ ;
	wire _w14096_ ;
	wire _w14095_ ;
	wire _w14094_ ;
	wire _w14093_ ;
	wire _w14092_ ;
	wire _w14091_ ;
	wire _w14090_ ;
	wire _w14089_ ;
	wire _w14088_ ;
	wire _w14087_ ;
	wire _w14086_ ;
	wire _w14085_ ;
	wire _w14084_ ;
	wire _w14083_ ;
	wire _w14082_ ;
	wire _w14081_ ;
	wire _w14080_ ;
	wire _w14079_ ;
	wire _w14078_ ;
	wire _w14077_ ;
	wire _w14076_ ;
	wire _w14075_ ;
	wire _w14074_ ;
	wire _w14073_ ;
	wire _w14072_ ;
	wire _w14071_ ;
	wire _w14070_ ;
	wire _w14069_ ;
	wire _w14068_ ;
	wire _w14067_ ;
	wire _w14066_ ;
	wire _w14065_ ;
	wire _w14064_ ;
	wire _w14063_ ;
	wire _w14062_ ;
	wire _w14061_ ;
	wire _w14060_ ;
	wire _w14059_ ;
	wire _w14058_ ;
	wire _w14057_ ;
	wire _w14056_ ;
	wire _w14055_ ;
	wire _w14054_ ;
	wire _w14053_ ;
	wire _w14052_ ;
	wire _w14051_ ;
	wire _w14050_ ;
	wire _w14049_ ;
	wire _w14048_ ;
	wire _w14047_ ;
	wire _w14046_ ;
	wire _w14045_ ;
	wire _w14044_ ;
	wire _w14043_ ;
	wire _w14042_ ;
	wire _w14041_ ;
	wire _w14040_ ;
	wire _w14039_ ;
	wire _w14038_ ;
	wire _w14037_ ;
	wire _w14036_ ;
	wire _w14035_ ;
	wire _w14034_ ;
	wire _w14033_ ;
	wire _w14032_ ;
	wire _w14031_ ;
	wire _w14030_ ;
	wire _w14029_ ;
	wire _w14028_ ;
	wire _w14027_ ;
	wire _w14026_ ;
	wire _w14025_ ;
	wire _w14024_ ;
	wire _w14023_ ;
	wire _w14022_ ;
	wire _w14021_ ;
	wire _w14020_ ;
	wire _w14019_ ;
	wire _w14018_ ;
	wire _w14017_ ;
	wire _w14016_ ;
	wire _w14015_ ;
	wire _w14014_ ;
	wire _w14013_ ;
	wire _w14012_ ;
	wire _w14011_ ;
	wire _w14010_ ;
	wire _w14009_ ;
	wire _w14008_ ;
	wire _w14007_ ;
	wire _w14006_ ;
	wire _w14005_ ;
	wire _w14004_ ;
	wire _w14003_ ;
	wire _w14002_ ;
	wire _w14001_ ;
	wire _w14000_ ;
	wire _w13999_ ;
	wire _w13998_ ;
	wire _w13997_ ;
	wire _w13996_ ;
	wire _w13995_ ;
	wire _w13994_ ;
	wire _w13993_ ;
	wire _w13992_ ;
	wire _w13991_ ;
	wire _w13990_ ;
	wire _w13989_ ;
	wire _w13988_ ;
	wire _w13987_ ;
	wire _w13986_ ;
	wire _w13985_ ;
	wire _w13984_ ;
	wire _w13983_ ;
	wire _w13982_ ;
	wire _w13981_ ;
	wire _w13980_ ;
	wire _w13979_ ;
	wire _w13978_ ;
	wire _w13977_ ;
	wire _w13976_ ;
	wire _w13975_ ;
	wire _w13974_ ;
	wire _w13973_ ;
	wire _w13972_ ;
	wire _w13971_ ;
	wire _w13970_ ;
	wire _w13969_ ;
	wire _w13968_ ;
	wire _w13967_ ;
	wire _w13966_ ;
	wire _w13965_ ;
	wire _w13964_ ;
	wire _w13963_ ;
	wire _w13962_ ;
	wire _w13961_ ;
	wire _w13960_ ;
	wire _w13959_ ;
	wire _w13958_ ;
	wire _w13957_ ;
	wire _w13956_ ;
	wire _w13955_ ;
	wire _w13954_ ;
	wire _w13953_ ;
	wire _w13952_ ;
	wire _w13951_ ;
	wire _w13950_ ;
	wire _w13949_ ;
	wire _w13948_ ;
	wire _w13947_ ;
	wire _w13946_ ;
	wire _w13945_ ;
	wire _w13944_ ;
	wire _w13943_ ;
	wire _w13942_ ;
	wire _w13941_ ;
	wire _w13940_ ;
	wire _w13939_ ;
	wire _w13938_ ;
	wire _w13937_ ;
	wire _w13936_ ;
	wire _w13935_ ;
	wire _w13934_ ;
	wire _w13933_ ;
	wire _w13932_ ;
	wire _w13931_ ;
	wire _w13930_ ;
	wire _w13929_ ;
	wire _w13928_ ;
	wire _w13927_ ;
	wire _w13926_ ;
	wire _w13925_ ;
	wire _w13924_ ;
	wire _w13923_ ;
	wire _w13922_ ;
	wire _w13921_ ;
	wire _w13920_ ;
	wire _w13919_ ;
	wire _w13918_ ;
	wire _w13917_ ;
	wire _w13916_ ;
	wire _w13915_ ;
	wire _w13914_ ;
	wire _w13913_ ;
	wire _w13912_ ;
	wire _w13911_ ;
	wire _w13910_ ;
	wire _w13909_ ;
	wire _w13908_ ;
	wire _w13907_ ;
	wire _w13906_ ;
	wire _w13905_ ;
	wire _w13904_ ;
	wire _w13903_ ;
	wire _w13902_ ;
	wire _w13901_ ;
	wire _w13900_ ;
	wire _w13899_ ;
	wire _w13898_ ;
	wire _w13897_ ;
	wire _w13896_ ;
	wire _w13895_ ;
	wire _w13894_ ;
	wire _w13893_ ;
	wire _w13892_ ;
	wire _w13891_ ;
	wire _w13890_ ;
	wire _w13889_ ;
	wire _w13888_ ;
	wire _w13887_ ;
	wire _w13886_ ;
	wire _w13885_ ;
	wire _w13884_ ;
	wire _w13883_ ;
	wire _w13882_ ;
	wire _w13881_ ;
	wire _w13880_ ;
	wire _w13879_ ;
	wire _w13878_ ;
	wire _w13877_ ;
	wire _w13876_ ;
	wire _w13875_ ;
	wire _w13874_ ;
	wire _w13873_ ;
	wire _w13872_ ;
	wire _w13871_ ;
	wire _w13870_ ;
	wire _w13869_ ;
	wire _w13868_ ;
	wire _w13867_ ;
	wire _w13866_ ;
	wire _w13865_ ;
	wire _w13864_ ;
	wire _w13863_ ;
	wire _w13862_ ;
	wire _w13861_ ;
	wire _w13860_ ;
	wire _w13859_ ;
	wire _w13858_ ;
	wire _w13857_ ;
	wire _w13856_ ;
	wire _w13855_ ;
	wire _w13854_ ;
	wire _w13853_ ;
	wire _w13852_ ;
	wire _w13851_ ;
	wire _w13850_ ;
	wire _w13849_ ;
	wire _w13848_ ;
	wire _w13847_ ;
	wire _w13846_ ;
	wire _w13845_ ;
	wire _w13844_ ;
	wire _w13843_ ;
	wire _w13842_ ;
	wire _w13841_ ;
	wire _w13840_ ;
	wire _w13839_ ;
	wire _w13838_ ;
	wire _w13837_ ;
	wire _w13836_ ;
	wire _w13835_ ;
	wire _w13834_ ;
	wire _w13833_ ;
	wire _w13832_ ;
	wire _w13831_ ;
	wire _w13830_ ;
	wire _w13829_ ;
	wire _w13828_ ;
	wire _w13827_ ;
	wire _w13826_ ;
	wire _w13825_ ;
	wire _w13824_ ;
	wire _w13823_ ;
	wire _w13822_ ;
	wire _w13821_ ;
	wire _w13820_ ;
	wire _w13819_ ;
	wire _w13818_ ;
	wire _w13817_ ;
	wire _w13816_ ;
	wire _w13815_ ;
	wire _w13814_ ;
	wire _w13813_ ;
	wire _w13812_ ;
	wire _w13811_ ;
	wire _w13810_ ;
	wire _w13809_ ;
	wire _w13808_ ;
	wire _w13807_ ;
	wire _w13806_ ;
	wire _w13805_ ;
	wire _w13804_ ;
	wire _w13803_ ;
	wire _w13802_ ;
	wire _w13801_ ;
	wire _w13800_ ;
	wire _w13799_ ;
	wire _w13798_ ;
	wire _w13797_ ;
	wire _w13796_ ;
	wire _w13795_ ;
	wire _w13794_ ;
	wire _w13793_ ;
	wire _w13792_ ;
	wire _w13791_ ;
	wire _w13790_ ;
	wire _w13789_ ;
	wire _w13788_ ;
	wire _w13787_ ;
	wire _w13786_ ;
	wire _w13785_ ;
	wire _w13784_ ;
	wire _w13783_ ;
	wire _w13782_ ;
	wire _w13781_ ;
	wire _w13780_ ;
	wire _w13779_ ;
	wire _w13778_ ;
	wire _w13777_ ;
	wire _w13776_ ;
	wire _w13775_ ;
	wire _w13774_ ;
	wire _w13773_ ;
	wire _w13772_ ;
	wire _w13771_ ;
	wire _w13770_ ;
	wire _w13769_ ;
	wire _w13768_ ;
	wire _w13767_ ;
	wire _w13766_ ;
	wire _w13765_ ;
	wire _w13764_ ;
	wire _w13763_ ;
	wire _w13762_ ;
	wire _w13761_ ;
	wire _w13760_ ;
	wire _w13759_ ;
	wire _w13758_ ;
	wire _w13757_ ;
	wire _w13756_ ;
	wire _w13755_ ;
	wire _w13754_ ;
	wire _w13753_ ;
	wire _w13752_ ;
	wire _w13751_ ;
	wire _w13750_ ;
	wire _w13749_ ;
	wire _w13748_ ;
	wire _w13747_ ;
	wire _w13746_ ;
	wire _w13745_ ;
	wire _w13744_ ;
	wire _w13743_ ;
	wire _w13742_ ;
	wire _w13741_ ;
	wire _w13740_ ;
	wire _w13739_ ;
	wire _w13738_ ;
	wire _w13737_ ;
	wire _w13736_ ;
	wire _w13735_ ;
	wire _w13734_ ;
	wire _w13733_ ;
	wire _w13732_ ;
	wire _w13731_ ;
	wire _w13730_ ;
	wire _w13729_ ;
	wire _w13728_ ;
	wire _w13727_ ;
	wire _w13726_ ;
	wire _w13725_ ;
	wire _w13724_ ;
	wire _w13723_ ;
	wire _w13722_ ;
	wire _w13721_ ;
	wire _w13720_ ;
	wire _w13719_ ;
	wire _w13718_ ;
	wire _w13717_ ;
	wire _w13716_ ;
	wire _w13715_ ;
	wire _w13714_ ;
	wire _w13713_ ;
	wire _w13712_ ;
	wire _w13711_ ;
	wire _w13710_ ;
	wire _w13709_ ;
	wire _w13708_ ;
	wire _w13707_ ;
	wire _w13706_ ;
	wire _w13705_ ;
	wire _w13704_ ;
	wire _w13703_ ;
	wire _w13702_ ;
	wire _w13701_ ;
	wire _w13700_ ;
	wire _w13699_ ;
	wire _w13698_ ;
	wire _w13697_ ;
	wire _w13696_ ;
	wire _w13695_ ;
	wire _w13694_ ;
	wire _w13693_ ;
	wire _w13692_ ;
	wire _w13691_ ;
	wire _w13690_ ;
	wire _w13689_ ;
	wire _w13688_ ;
	wire _w13687_ ;
	wire _w13686_ ;
	wire _w13685_ ;
	wire _w13684_ ;
	wire _w13683_ ;
	wire _w13682_ ;
	wire _w13681_ ;
	wire _w13680_ ;
	wire _w13679_ ;
	wire _w13678_ ;
	wire _w13677_ ;
	wire _w13676_ ;
	wire _w13675_ ;
	wire _w13674_ ;
	wire _w13673_ ;
	wire _w13672_ ;
	wire _w13671_ ;
	wire _w13670_ ;
	wire _w13669_ ;
	wire _w13668_ ;
	wire _w13667_ ;
	wire _w13666_ ;
	wire _w13665_ ;
	wire _w13664_ ;
	wire _w13663_ ;
	wire _w13662_ ;
	wire _w13661_ ;
	wire _w13660_ ;
	wire _w13659_ ;
	wire _w13658_ ;
	wire _w13657_ ;
	wire _w13656_ ;
	wire _w13655_ ;
	wire _w13654_ ;
	wire _w13653_ ;
	wire _w13652_ ;
	wire _w13651_ ;
	wire _w13650_ ;
	wire _w13649_ ;
	wire _w13648_ ;
	wire _w13647_ ;
	wire _w13646_ ;
	wire _w13645_ ;
	wire _w13644_ ;
	wire _w13643_ ;
	wire _w13642_ ;
	wire _w13641_ ;
	wire _w13640_ ;
	wire _w13639_ ;
	wire _w13638_ ;
	wire _w13637_ ;
	wire _w13636_ ;
	wire _w13635_ ;
	wire _w13634_ ;
	wire _w13633_ ;
	wire _w13632_ ;
	wire _w13631_ ;
	wire _w13630_ ;
	wire _w13629_ ;
	wire _w13628_ ;
	wire _w13627_ ;
	wire _w13626_ ;
	wire _w13625_ ;
	wire _w13624_ ;
	wire _w13623_ ;
	wire _w13622_ ;
	wire _w13621_ ;
	wire _w13620_ ;
	wire _w13619_ ;
	wire _w13618_ ;
	wire _w13617_ ;
	wire _w13616_ ;
	wire _w13615_ ;
	wire _w13614_ ;
	wire _w13613_ ;
	wire _w13612_ ;
	wire _w13611_ ;
	wire _w13610_ ;
	wire _w13609_ ;
	wire _w13608_ ;
	wire _w13607_ ;
	wire _w13606_ ;
	wire _w13605_ ;
	wire _w13604_ ;
	wire _w13603_ ;
	wire _w13602_ ;
	wire _w13601_ ;
	wire _w13600_ ;
	wire _w13599_ ;
	wire _w13598_ ;
	wire _w13597_ ;
	wire _w13596_ ;
	wire _w13595_ ;
	wire _w13594_ ;
	wire _w13593_ ;
	wire _w13592_ ;
	wire _w13591_ ;
	wire _w13590_ ;
	wire _w13589_ ;
	wire _w13588_ ;
	wire _w13587_ ;
	wire _w13586_ ;
	wire _w13585_ ;
	wire _w13584_ ;
	wire _w13583_ ;
	wire _w13582_ ;
	wire _w13581_ ;
	wire _w13580_ ;
	wire _w13579_ ;
	wire _w13578_ ;
	wire _w13577_ ;
	wire _w13576_ ;
	wire _w13575_ ;
	wire _w13574_ ;
	wire _w13573_ ;
	wire _w13572_ ;
	wire _w13571_ ;
	wire _w13570_ ;
	wire _w13569_ ;
	wire _w13568_ ;
	wire _w13567_ ;
	wire _w13566_ ;
	wire _w13565_ ;
	wire _w13564_ ;
	wire _w13563_ ;
	wire _w13562_ ;
	wire _w13561_ ;
	wire _w13560_ ;
	wire _w13559_ ;
	wire _w13558_ ;
	wire _w13557_ ;
	wire _w13556_ ;
	wire _w13555_ ;
	wire _w13554_ ;
	wire _w13553_ ;
	wire _w13552_ ;
	wire _w13551_ ;
	wire _w13550_ ;
	wire _w13549_ ;
	wire _w13548_ ;
	wire _w13547_ ;
	wire _w13546_ ;
	wire _w13545_ ;
	wire _w13544_ ;
	wire _w13543_ ;
	wire _w13542_ ;
	wire _w13541_ ;
	wire _w13540_ ;
	wire _w13539_ ;
	wire _w13538_ ;
	wire _w13537_ ;
	wire _w13536_ ;
	wire _w13535_ ;
	wire _w13534_ ;
	wire _w13533_ ;
	wire _w13532_ ;
	wire _w13531_ ;
	wire _w13530_ ;
	wire _w13529_ ;
	wire _w13528_ ;
	wire _w13527_ ;
	wire _w13526_ ;
	wire _w13525_ ;
	wire _w13524_ ;
	wire _w13523_ ;
	wire _w13522_ ;
	wire _w13521_ ;
	wire _w13520_ ;
	wire _w13519_ ;
	wire _w13518_ ;
	wire _w13517_ ;
	wire _w13516_ ;
	wire _w13515_ ;
	wire _w13514_ ;
	wire _w13513_ ;
	wire _w13512_ ;
	wire _w13511_ ;
	wire _w13510_ ;
	wire _w13509_ ;
	wire _w13508_ ;
	wire _w13507_ ;
	wire _w13506_ ;
	wire _w13505_ ;
	wire _w13504_ ;
	wire _w13503_ ;
	wire _w13502_ ;
	wire _w13501_ ;
	wire _w13500_ ;
	wire _w13499_ ;
	wire _w13498_ ;
	wire _w13497_ ;
	wire _w13496_ ;
	wire _w13495_ ;
	wire _w13494_ ;
	wire _w13493_ ;
	wire _w13492_ ;
	wire _w13491_ ;
	wire _w13490_ ;
	wire _w13489_ ;
	wire _w13488_ ;
	wire _w13487_ ;
	wire _w13486_ ;
	wire _w13485_ ;
	wire _w13484_ ;
	wire _w13483_ ;
	wire _w13482_ ;
	wire _w13481_ ;
	wire _w13480_ ;
	wire _w13479_ ;
	wire _w13478_ ;
	wire _w13477_ ;
	wire _w13476_ ;
	wire _w13475_ ;
	wire _w13474_ ;
	wire _w13473_ ;
	wire _w13472_ ;
	wire _w13471_ ;
	wire _w13470_ ;
	wire _w13469_ ;
	wire _w13468_ ;
	wire _w13467_ ;
	wire _w13466_ ;
	wire _w13465_ ;
	wire _w13464_ ;
	wire _w13463_ ;
	wire _w13462_ ;
	wire _w13461_ ;
	wire _w13460_ ;
	wire _w13459_ ;
	wire _w13458_ ;
	wire _w13457_ ;
	wire _w13456_ ;
	wire _w13455_ ;
	wire _w13454_ ;
	wire _w13453_ ;
	wire _w13452_ ;
	wire _w13451_ ;
	wire _w13450_ ;
	wire _w13449_ ;
	wire _w13448_ ;
	wire _w13447_ ;
	wire _w13446_ ;
	wire _w13445_ ;
	wire _w13444_ ;
	wire _w13443_ ;
	wire _w13442_ ;
	wire _w13441_ ;
	wire _w13440_ ;
	wire _w13439_ ;
	wire _w13438_ ;
	wire _w13437_ ;
	wire _w13436_ ;
	wire _w13435_ ;
	wire _w13434_ ;
	wire _w13433_ ;
	wire _w13432_ ;
	wire _w13431_ ;
	wire _w13430_ ;
	wire _w13429_ ;
	wire _w13428_ ;
	wire _w13427_ ;
	wire _w13426_ ;
	wire _w13425_ ;
	wire _w13424_ ;
	wire _w13423_ ;
	wire _w13422_ ;
	wire _w13421_ ;
	wire _w13420_ ;
	wire _w13419_ ;
	wire _w13418_ ;
	wire _w13417_ ;
	wire _w13416_ ;
	wire _w13415_ ;
	wire _w13414_ ;
	wire _w13413_ ;
	wire _w13412_ ;
	wire _w13411_ ;
	wire _w13410_ ;
	wire _w13409_ ;
	wire _w13408_ ;
	wire _w13407_ ;
	wire _w13406_ ;
	wire _w13405_ ;
	wire _w13404_ ;
	wire _w13403_ ;
	wire _w13402_ ;
	wire _w13401_ ;
	wire _w13400_ ;
	wire _w13399_ ;
	wire _w13398_ ;
	wire _w13397_ ;
	wire _w13396_ ;
	wire _w13395_ ;
	wire _w13394_ ;
	wire _w13393_ ;
	wire _w13392_ ;
	wire _w13391_ ;
	wire _w13390_ ;
	wire _w13389_ ;
	wire _w13388_ ;
	wire _w13387_ ;
	wire _w13386_ ;
	wire _w13385_ ;
	wire _w13384_ ;
	wire _w13383_ ;
	wire _w13382_ ;
	wire _w13381_ ;
	wire _w13380_ ;
	wire _w13379_ ;
	wire _w13378_ ;
	wire _w13377_ ;
	wire _w13376_ ;
	wire _w13375_ ;
	wire _w13374_ ;
	wire _w13373_ ;
	wire _w13372_ ;
	wire _w13371_ ;
	wire _w13370_ ;
	wire _w13369_ ;
	wire _w13368_ ;
	wire _w13367_ ;
	wire _w13366_ ;
	wire _w13365_ ;
	wire _w13364_ ;
	wire _w13363_ ;
	wire _w13362_ ;
	wire _w13361_ ;
	wire _w13360_ ;
	wire _w13359_ ;
	wire _w13358_ ;
	wire _w13357_ ;
	wire _w13356_ ;
	wire _w13355_ ;
	wire _w13354_ ;
	wire _w13353_ ;
	wire _w13352_ ;
	wire _w13351_ ;
	wire _w13350_ ;
	wire _w13349_ ;
	wire _w13348_ ;
	wire _w13347_ ;
	wire _w13346_ ;
	wire _w13345_ ;
	wire _w13344_ ;
	wire _w13343_ ;
	wire _w13342_ ;
	wire _w13341_ ;
	wire _w13340_ ;
	wire _w13339_ ;
	wire _w13338_ ;
	wire _w13337_ ;
	wire _w13336_ ;
	wire _w13335_ ;
	wire _w13334_ ;
	wire _w13333_ ;
	wire _w13332_ ;
	wire _w13331_ ;
	wire _w13330_ ;
	wire _w13329_ ;
	wire _w13328_ ;
	wire _w13327_ ;
	wire _w13326_ ;
	wire _w13325_ ;
	wire _w13324_ ;
	wire _w13323_ ;
	wire _w13322_ ;
	wire _w13321_ ;
	wire _w13320_ ;
	wire _w13319_ ;
	wire _w13318_ ;
	wire _w13317_ ;
	wire _w13316_ ;
	wire _w13315_ ;
	wire _w13314_ ;
	wire _w13313_ ;
	wire _w13312_ ;
	wire _w13311_ ;
	wire _w13310_ ;
	wire _w13309_ ;
	wire _w13308_ ;
	wire _w13307_ ;
	wire _w13306_ ;
	wire _w13305_ ;
	wire _w13304_ ;
	wire _w13303_ ;
	wire _w13302_ ;
	wire _w13301_ ;
	wire _w13300_ ;
	wire _w13299_ ;
	wire _w13298_ ;
	wire _w13297_ ;
	wire _w13296_ ;
	wire _w13295_ ;
	wire _w13294_ ;
	wire _w13293_ ;
	wire _w13292_ ;
	wire _w13291_ ;
	wire _w13290_ ;
	wire _w13289_ ;
	wire _w13288_ ;
	wire _w13287_ ;
	wire _w13286_ ;
	wire _w13285_ ;
	wire _w13284_ ;
	wire _w13283_ ;
	wire _w13282_ ;
	wire _w13281_ ;
	wire _w13280_ ;
	wire _w13279_ ;
	wire _w13278_ ;
	wire _w13277_ ;
	wire _w13276_ ;
	wire _w13275_ ;
	wire _w13274_ ;
	wire _w13273_ ;
	wire _w13272_ ;
	wire _w13271_ ;
	wire _w13270_ ;
	wire _w13269_ ;
	wire _w13268_ ;
	wire _w13267_ ;
	wire _w13266_ ;
	wire _w13265_ ;
	wire _w13264_ ;
	wire _w13263_ ;
	wire _w13262_ ;
	wire _w13261_ ;
	wire _w13260_ ;
	wire _w13259_ ;
	wire _w13258_ ;
	wire _w13257_ ;
	wire _w13256_ ;
	wire _w13255_ ;
	wire _w13254_ ;
	wire _w13253_ ;
	wire _w13252_ ;
	wire _w13251_ ;
	wire _w13250_ ;
	wire _w13249_ ;
	wire _w13248_ ;
	wire _w13247_ ;
	wire _w13246_ ;
	wire _w13245_ ;
	wire _w13244_ ;
	wire _w13243_ ;
	wire _w13242_ ;
	wire _w13241_ ;
	wire _w13240_ ;
	wire _w13239_ ;
	wire _w13238_ ;
	wire _w13237_ ;
	wire _w13236_ ;
	wire _w13235_ ;
	wire _w13234_ ;
	wire _w13233_ ;
	wire _w13232_ ;
	wire _w13231_ ;
	wire _w13230_ ;
	wire _w13229_ ;
	wire _w13228_ ;
	wire _w13227_ ;
	wire _w13226_ ;
	wire _w13225_ ;
	wire _w13224_ ;
	wire _w13223_ ;
	wire _w13222_ ;
	wire _w13221_ ;
	wire _w13220_ ;
	wire _w13219_ ;
	wire _w13218_ ;
	wire _w13217_ ;
	wire _w13216_ ;
	wire _w13215_ ;
	wire _w13214_ ;
	wire _w13213_ ;
	wire _w13212_ ;
	wire _w13211_ ;
	wire _w13210_ ;
	wire _w13209_ ;
	wire _w13208_ ;
	wire _w13207_ ;
	wire _w13206_ ;
	wire _w13205_ ;
	wire _w13204_ ;
	wire _w13203_ ;
	wire _w13202_ ;
	wire _w13201_ ;
	wire _w13200_ ;
	wire _w13199_ ;
	wire _w13198_ ;
	wire _w13197_ ;
	wire _w13196_ ;
	wire _w13195_ ;
	wire _w13194_ ;
	wire _w13193_ ;
	wire _w13192_ ;
	wire _w13191_ ;
	wire _w13190_ ;
	wire _w13189_ ;
	wire _w13188_ ;
	wire _w13187_ ;
	wire _w13186_ ;
	wire _w13185_ ;
	wire _w13184_ ;
	wire _w13183_ ;
	wire _w13182_ ;
	wire _w13181_ ;
	wire _w13180_ ;
	wire _w13179_ ;
	wire _w13178_ ;
	wire _w13177_ ;
	wire _w13176_ ;
	wire _w13175_ ;
	wire _w13174_ ;
	wire _w13173_ ;
	wire _w13172_ ;
	wire _w13171_ ;
	wire _w13170_ ;
	wire _w13169_ ;
	wire _w13168_ ;
	wire _w13167_ ;
	wire _w13166_ ;
	wire _w13165_ ;
	wire _w13164_ ;
	wire _w13163_ ;
	wire _w13162_ ;
	wire _w13161_ ;
	wire _w13160_ ;
	wire _w13159_ ;
	wire _w13158_ ;
	wire _w13157_ ;
	wire _w13156_ ;
	wire _w13155_ ;
	wire _w13154_ ;
	wire _w13153_ ;
	wire _w13152_ ;
	wire _w13151_ ;
	wire _w13150_ ;
	wire _w13149_ ;
	wire _w13148_ ;
	wire _w13147_ ;
	wire _w13146_ ;
	wire _w13145_ ;
	wire _w13144_ ;
	wire _w13143_ ;
	wire _w13142_ ;
	wire _w13141_ ;
	wire _w13140_ ;
	wire _w13139_ ;
	wire _w13138_ ;
	wire _w13137_ ;
	wire _w13136_ ;
	wire _w13135_ ;
	wire _w13134_ ;
	wire _w13133_ ;
	wire _w13132_ ;
	wire _w13131_ ;
	wire _w13130_ ;
	wire _w13129_ ;
	wire _w13128_ ;
	wire _w13127_ ;
	wire _w13126_ ;
	wire _w13125_ ;
	wire _w13124_ ;
	wire _w13123_ ;
	wire _w13122_ ;
	wire _w13121_ ;
	wire _w13120_ ;
	wire _w13119_ ;
	wire _w13118_ ;
	wire _w13117_ ;
	wire _w13116_ ;
	wire _w13115_ ;
	wire _w13114_ ;
	wire _w13113_ ;
	wire _w13112_ ;
	wire _w13111_ ;
	wire _w13110_ ;
	wire _w13109_ ;
	wire _w13108_ ;
	wire _w13107_ ;
	wire _w13106_ ;
	wire _w13105_ ;
	wire _w13104_ ;
	wire _w13103_ ;
	wire _w13102_ ;
	wire _w13101_ ;
	wire _w13100_ ;
	wire _w13099_ ;
	wire _w13098_ ;
	wire _w13097_ ;
	wire _w13096_ ;
	wire _w13095_ ;
	wire _w13094_ ;
	wire _w13093_ ;
	wire _w13092_ ;
	wire _w13091_ ;
	wire _w13090_ ;
	wire _w13089_ ;
	wire _w13088_ ;
	wire _w13087_ ;
	wire _w13086_ ;
	wire _w13085_ ;
	wire _w13084_ ;
	wire _w13083_ ;
	wire _w13082_ ;
	wire _w13081_ ;
	wire _w13080_ ;
	wire _w13079_ ;
	wire _w13078_ ;
	wire _w13077_ ;
	wire _w13076_ ;
	wire _w13075_ ;
	wire _w13074_ ;
	wire _w13073_ ;
	wire _w13072_ ;
	wire _w13071_ ;
	wire _w13070_ ;
	wire _w13069_ ;
	wire _w13068_ ;
	wire _w13067_ ;
	wire _w13066_ ;
	wire _w13065_ ;
	wire _w13064_ ;
	wire _w13063_ ;
	wire _w13062_ ;
	wire _w13061_ ;
	wire _w13060_ ;
	wire _w13059_ ;
	wire _w13058_ ;
	wire _w13057_ ;
	wire _w13056_ ;
	wire _w13055_ ;
	wire _w13054_ ;
	wire _w13053_ ;
	wire _w13052_ ;
	wire _w13051_ ;
	wire _w13050_ ;
	wire _w13049_ ;
	wire _w13048_ ;
	wire _w13047_ ;
	wire _w13046_ ;
	wire _w13045_ ;
	wire _w13044_ ;
	wire _w13043_ ;
	wire _w13042_ ;
	wire _w13041_ ;
	wire _w13040_ ;
	wire _w13039_ ;
	wire _w13038_ ;
	wire _w13037_ ;
	wire _w13036_ ;
	wire _w13035_ ;
	wire _w13034_ ;
	wire _w13033_ ;
	wire _w13032_ ;
	wire _w13031_ ;
	wire _w13030_ ;
	wire _w13029_ ;
	wire _w13028_ ;
	wire _w13027_ ;
	wire _w13026_ ;
	wire _w13025_ ;
	wire _w13024_ ;
	wire _w13023_ ;
	wire _w13022_ ;
	wire _w13021_ ;
	wire _w13020_ ;
	wire _w13019_ ;
	wire _w13018_ ;
	wire _w13017_ ;
	wire _w13016_ ;
	wire _w13015_ ;
	wire _w13014_ ;
	wire _w13013_ ;
	wire _w13012_ ;
	wire _w13011_ ;
	wire _w13010_ ;
	wire _w13009_ ;
	wire _w13008_ ;
	wire _w13007_ ;
	wire _w13006_ ;
	wire _w13005_ ;
	wire _w13004_ ;
	wire _w13003_ ;
	wire _w13002_ ;
	wire _w13001_ ;
	wire _w13000_ ;
	wire _w12999_ ;
	wire _w12998_ ;
	wire _w12997_ ;
	wire _w12996_ ;
	wire _w12995_ ;
	wire _w12994_ ;
	wire _w12993_ ;
	wire _w12992_ ;
	wire _w12991_ ;
	wire _w12990_ ;
	wire _w12989_ ;
	wire _w12988_ ;
	wire _w12987_ ;
	wire _w12986_ ;
	wire _w12985_ ;
	wire _w12984_ ;
	wire _w12983_ ;
	wire _w12982_ ;
	wire _w12981_ ;
	wire _w12980_ ;
	wire _w12979_ ;
	wire _w12978_ ;
	wire _w12977_ ;
	wire _w12976_ ;
	wire _w12975_ ;
	wire _w12974_ ;
	wire _w12973_ ;
	wire _w12972_ ;
	wire _w12971_ ;
	wire _w12970_ ;
	wire _w12969_ ;
	wire _w12968_ ;
	wire _w12967_ ;
	wire _w12966_ ;
	wire _w12965_ ;
	wire _w12964_ ;
	wire _w12963_ ;
	wire _w12962_ ;
	wire _w12961_ ;
	wire _w12960_ ;
	wire _w12959_ ;
	wire _w12958_ ;
	wire _w12957_ ;
	wire _w12956_ ;
	wire _w12955_ ;
	wire _w12954_ ;
	wire _w12953_ ;
	wire _w12952_ ;
	wire _w12951_ ;
	wire _w12950_ ;
	wire _w12949_ ;
	wire _w12948_ ;
	wire _w12947_ ;
	wire _w12946_ ;
	wire _w12945_ ;
	wire _w12944_ ;
	wire _w12943_ ;
	wire _w12942_ ;
	wire _w12941_ ;
	wire _w12940_ ;
	wire _w12939_ ;
	wire _w12938_ ;
	wire _w12937_ ;
	wire _w12936_ ;
	wire _w12935_ ;
	wire _w12934_ ;
	wire _w12933_ ;
	wire _w12932_ ;
	wire _w12931_ ;
	wire _w12930_ ;
	wire _w12929_ ;
	wire _w12928_ ;
	wire _w12927_ ;
	wire _w12926_ ;
	wire _w12925_ ;
	wire _w12924_ ;
	wire _w12923_ ;
	wire _w12922_ ;
	wire _w12921_ ;
	wire _w12920_ ;
	wire _w12919_ ;
	wire _w12918_ ;
	wire _w12917_ ;
	wire _w12916_ ;
	wire _w12915_ ;
	wire _w12914_ ;
	wire _w12913_ ;
	wire _w12912_ ;
	wire _w12911_ ;
	wire _w12910_ ;
	wire _w12909_ ;
	wire _w12908_ ;
	wire _w12907_ ;
	wire _w12906_ ;
	wire _w12905_ ;
	wire _w12904_ ;
	wire _w12903_ ;
	wire _w12902_ ;
	wire _w12901_ ;
	wire _w12900_ ;
	wire _w12899_ ;
	wire _w12898_ ;
	wire _w12897_ ;
	wire _w12896_ ;
	wire _w12895_ ;
	wire _w12894_ ;
	wire _w12893_ ;
	wire _w12892_ ;
	wire _w12891_ ;
	wire _w12890_ ;
	wire _w12889_ ;
	wire _w12888_ ;
	wire _w12887_ ;
	wire _w12886_ ;
	wire _w12885_ ;
	wire _w12884_ ;
	wire _w12883_ ;
	wire _w12882_ ;
	wire _w12881_ ;
	wire _w12880_ ;
	wire _w12879_ ;
	wire _w12878_ ;
	wire _w12877_ ;
	wire _w12876_ ;
	wire _w12875_ ;
	wire _w12874_ ;
	wire _w12873_ ;
	wire _w12872_ ;
	wire _w12871_ ;
	wire _w12870_ ;
	wire _w12869_ ;
	wire _w12868_ ;
	wire _w12867_ ;
	wire _w12866_ ;
	wire _w12865_ ;
	wire _w12864_ ;
	wire _w12863_ ;
	wire _w12862_ ;
	wire _w12861_ ;
	wire _w12860_ ;
	wire _w12859_ ;
	wire _w12858_ ;
	wire _w12857_ ;
	wire _w12856_ ;
	wire _w12855_ ;
	wire _w12854_ ;
	wire _w12853_ ;
	wire _w12852_ ;
	wire _w12851_ ;
	wire _w12850_ ;
	wire _w12849_ ;
	wire _w12848_ ;
	wire _w12847_ ;
	wire _w12846_ ;
	wire _w12845_ ;
	wire _w12844_ ;
	wire _w12843_ ;
	wire _w12842_ ;
	wire _w12841_ ;
	wire _w12840_ ;
	wire _w12839_ ;
	wire _w12838_ ;
	wire _w12837_ ;
	wire _w12836_ ;
	wire _w12835_ ;
	wire _w12834_ ;
	wire _w12833_ ;
	wire _w12832_ ;
	wire _w12831_ ;
	wire _w12830_ ;
	wire _w12829_ ;
	wire _w12828_ ;
	wire _w12827_ ;
	wire _w12826_ ;
	wire _w12825_ ;
	wire _w12824_ ;
	wire _w12823_ ;
	wire _w12822_ ;
	wire _w12821_ ;
	wire _w12820_ ;
	wire _w12819_ ;
	wire _w12818_ ;
	wire _w12817_ ;
	wire _w12816_ ;
	wire _w12815_ ;
	wire _w12814_ ;
	wire _w12813_ ;
	wire _w12812_ ;
	wire _w12811_ ;
	wire _w12810_ ;
	wire _w12809_ ;
	wire _w12808_ ;
	wire _w12807_ ;
	wire _w12806_ ;
	wire _w12805_ ;
	wire _w12804_ ;
	wire _w12803_ ;
	wire _w12802_ ;
	wire _w12801_ ;
	wire _w12800_ ;
	wire _w12799_ ;
	wire _w12798_ ;
	wire _w12797_ ;
	wire _w12796_ ;
	wire _w12795_ ;
	wire _w12794_ ;
	wire _w12793_ ;
	wire _w12792_ ;
	wire _w12791_ ;
	wire _w12790_ ;
	wire _w12789_ ;
	wire _w12788_ ;
	wire _w12787_ ;
	wire _w12786_ ;
	wire _w12785_ ;
	wire _w12784_ ;
	wire _w12783_ ;
	wire _w12782_ ;
	wire _w12781_ ;
	wire _w12780_ ;
	wire _w12779_ ;
	wire _w12778_ ;
	wire _w12777_ ;
	wire _w12776_ ;
	wire _w12775_ ;
	wire _w12774_ ;
	wire _w12773_ ;
	wire _w12772_ ;
	wire _w12771_ ;
	wire _w12770_ ;
	wire _w12769_ ;
	wire _w12768_ ;
	wire _w12767_ ;
	wire _w12766_ ;
	wire _w12765_ ;
	wire _w12764_ ;
	wire _w12763_ ;
	wire _w12762_ ;
	wire _w12761_ ;
	wire _w12760_ ;
	wire _w12759_ ;
	wire _w12758_ ;
	wire _w12757_ ;
	wire _w12756_ ;
	wire _w12755_ ;
	wire _w12754_ ;
	wire _w12753_ ;
	wire _w12752_ ;
	wire _w12751_ ;
	wire _w12750_ ;
	wire _w12749_ ;
	wire _w12748_ ;
	wire _w12747_ ;
	wire _w12746_ ;
	wire _w12745_ ;
	wire _w12744_ ;
	wire _w12743_ ;
	wire _w12742_ ;
	wire _w12741_ ;
	wire _w12740_ ;
	wire _w12739_ ;
	wire _w12738_ ;
	wire _w12737_ ;
	wire _w12736_ ;
	wire _w12735_ ;
	wire _w12734_ ;
	wire _w12733_ ;
	wire _w12732_ ;
	wire _w12731_ ;
	wire _w12730_ ;
	wire _w12729_ ;
	wire _w12728_ ;
	wire _w12727_ ;
	wire _w12726_ ;
	wire _w12725_ ;
	wire _w12724_ ;
	wire _w12723_ ;
	wire _w12722_ ;
	wire _w12721_ ;
	wire _w12720_ ;
	wire _w12719_ ;
	wire _w12718_ ;
	wire _w12717_ ;
	wire _w12716_ ;
	wire _w12715_ ;
	wire _w12714_ ;
	wire _w12713_ ;
	wire _w12712_ ;
	wire _w12711_ ;
	wire _w12710_ ;
	wire _w12709_ ;
	wire _w12708_ ;
	wire _w12707_ ;
	wire _w12706_ ;
	wire _w12705_ ;
	wire _w12704_ ;
	wire _w12703_ ;
	wire _w12702_ ;
	wire _w12701_ ;
	wire _w12700_ ;
	wire _w12699_ ;
	wire _w12698_ ;
	wire _w12697_ ;
	wire _w12696_ ;
	wire _w12695_ ;
	wire _w12694_ ;
	wire _w12693_ ;
	wire _w12692_ ;
	wire _w12691_ ;
	wire _w12690_ ;
	wire _w12689_ ;
	wire _w12688_ ;
	wire _w12687_ ;
	wire _w12686_ ;
	wire _w12685_ ;
	wire _w12684_ ;
	wire _w12683_ ;
	wire _w12682_ ;
	wire _w12681_ ;
	wire _w12680_ ;
	wire _w12679_ ;
	wire _w12678_ ;
	wire _w12677_ ;
	wire _w12676_ ;
	wire _w12675_ ;
	wire _w12674_ ;
	wire _w12673_ ;
	wire _w12672_ ;
	wire _w12671_ ;
	wire _w12670_ ;
	wire _w12669_ ;
	wire _w12668_ ;
	wire _w12667_ ;
	wire _w12666_ ;
	wire _w12665_ ;
	wire _w12664_ ;
	wire _w12663_ ;
	wire _w12662_ ;
	wire _w12661_ ;
	wire _w12660_ ;
	wire _w12659_ ;
	wire _w12658_ ;
	wire _w12657_ ;
	wire _w12656_ ;
	wire _w12655_ ;
	wire _w12654_ ;
	wire _w12653_ ;
	wire _w12652_ ;
	wire _w12651_ ;
	wire _w12650_ ;
	wire _w12649_ ;
	wire _w12648_ ;
	wire _w12647_ ;
	wire _w12646_ ;
	wire _w12645_ ;
	wire _w12644_ ;
	wire _w12643_ ;
	wire _w12642_ ;
	wire _w12641_ ;
	wire _w12640_ ;
	wire _w12639_ ;
	wire _w12638_ ;
	wire _w12637_ ;
	wire _w12636_ ;
	wire _w12635_ ;
	wire _w12634_ ;
	wire _w12633_ ;
	wire _w12632_ ;
	wire _w12631_ ;
	wire _w12630_ ;
	wire _w12629_ ;
	wire _w12628_ ;
	wire _w12627_ ;
	wire _w12626_ ;
	wire _w12625_ ;
	wire _w12624_ ;
	wire _w12623_ ;
	wire _w12622_ ;
	wire _w12621_ ;
	wire _w12620_ ;
	wire _w12619_ ;
	wire _w12618_ ;
	wire _w12617_ ;
	wire _w12616_ ;
	wire _w12615_ ;
	wire _w12614_ ;
	wire _w12613_ ;
	wire _w12612_ ;
	wire _w12611_ ;
	wire _w12610_ ;
	wire _w12609_ ;
	wire _w12608_ ;
	wire _w12607_ ;
	wire _w12606_ ;
	wire _w12605_ ;
	wire _w12604_ ;
	wire _w12603_ ;
	wire _w12602_ ;
	wire _w12601_ ;
	wire _w12600_ ;
	wire _w12599_ ;
	wire _w12598_ ;
	wire _w12597_ ;
	wire _w12596_ ;
	wire _w12595_ ;
	wire _w12594_ ;
	wire _w12593_ ;
	wire _w12592_ ;
	wire _w12591_ ;
	wire _w12590_ ;
	wire _w12589_ ;
	wire _w12588_ ;
	wire _w12587_ ;
	wire _w12586_ ;
	wire _w12585_ ;
	wire _w12584_ ;
	wire _w12583_ ;
	wire _w12582_ ;
	wire _w12581_ ;
	wire _w12580_ ;
	wire _w12579_ ;
	wire _w12578_ ;
	wire _w12577_ ;
	wire _w12576_ ;
	wire _w12575_ ;
	wire _w12574_ ;
	wire _w12573_ ;
	wire _w12572_ ;
	wire _w12571_ ;
	wire _w12570_ ;
	wire _w12569_ ;
	wire _w12568_ ;
	wire _w12567_ ;
	wire _w12566_ ;
	wire _w12565_ ;
	wire _w12564_ ;
	wire _w12563_ ;
	wire _w12562_ ;
	wire _w12561_ ;
	wire _w12560_ ;
	wire _w12559_ ;
	wire _w12558_ ;
	wire _w12557_ ;
	wire _w12556_ ;
	wire _w12555_ ;
	wire _w12554_ ;
	wire _w12553_ ;
	wire _w12552_ ;
	wire _w12551_ ;
	wire _w12550_ ;
	wire _w12549_ ;
	wire _w12548_ ;
	wire _w12547_ ;
	wire _w12546_ ;
	wire _w12545_ ;
	wire _w12544_ ;
	wire _w12543_ ;
	wire _w12542_ ;
	wire _w12541_ ;
	wire _w12540_ ;
	wire _w12539_ ;
	wire _w12538_ ;
	wire _w12537_ ;
	wire _w12536_ ;
	wire _w12535_ ;
	wire _w12534_ ;
	wire _w12533_ ;
	wire _w12532_ ;
	wire _w12531_ ;
	wire _w12530_ ;
	wire _w12529_ ;
	wire _w12528_ ;
	wire _w12527_ ;
	wire _w12526_ ;
	wire _w12525_ ;
	wire _w12524_ ;
	wire _w12523_ ;
	wire _w12522_ ;
	wire _w12521_ ;
	wire _w12520_ ;
	wire _w12519_ ;
	wire _w12518_ ;
	wire _w12517_ ;
	wire _w12516_ ;
	wire _w12515_ ;
	wire _w12514_ ;
	wire _w12513_ ;
	wire _w12512_ ;
	wire _w12511_ ;
	wire _w12510_ ;
	wire _w12509_ ;
	wire _w12508_ ;
	wire _w12507_ ;
	wire _w12506_ ;
	wire _w12505_ ;
	wire _w12504_ ;
	wire _w12503_ ;
	wire _w12502_ ;
	wire _w12501_ ;
	wire _w12500_ ;
	wire _w12499_ ;
	wire _w12498_ ;
	wire _w12497_ ;
	wire _w12496_ ;
	wire _w12495_ ;
	wire _w12494_ ;
	wire _w12493_ ;
	wire _w12492_ ;
	wire _w12491_ ;
	wire _w12490_ ;
	wire _w12489_ ;
	wire _w12488_ ;
	wire _w12487_ ;
	wire _w12486_ ;
	wire _w12485_ ;
	wire _w12484_ ;
	wire _w12483_ ;
	wire _w12482_ ;
	wire _w12481_ ;
	wire _w12480_ ;
	wire _w12479_ ;
	wire _w12478_ ;
	wire _w12477_ ;
	wire _w12476_ ;
	wire _w12475_ ;
	wire _w12474_ ;
	wire _w12473_ ;
	wire _w12472_ ;
	wire _w12471_ ;
	wire _w12470_ ;
	wire _w12469_ ;
	wire _w12468_ ;
	wire _w12467_ ;
	wire _w12466_ ;
	wire _w12465_ ;
	wire _w12464_ ;
	wire _w12463_ ;
	wire _w12462_ ;
	wire _w12461_ ;
	wire _w12460_ ;
	wire _w12459_ ;
	wire _w12458_ ;
	wire _w12457_ ;
	wire _w12456_ ;
	wire _w12455_ ;
	wire _w12454_ ;
	wire _w12453_ ;
	wire _w12452_ ;
	wire _w12451_ ;
	wire _w12450_ ;
	wire _w12449_ ;
	wire _w12448_ ;
	wire _w12447_ ;
	wire _w12446_ ;
	wire _w12445_ ;
	wire _w12444_ ;
	wire _w12443_ ;
	wire _w12442_ ;
	wire _w12441_ ;
	wire _w12440_ ;
	wire _w12439_ ;
	wire _w12438_ ;
	wire _w12437_ ;
	wire _w12436_ ;
	wire _w12435_ ;
	wire _w12434_ ;
	wire _w12433_ ;
	wire _w12432_ ;
	wire _w12431_ ;
	wire _w12430_ ;
	wire _w12429_ ;
	wire _w12428_ ;
	wire _w12427_ ;
	wire _w12426_ ;
	wire _w12425_ ;
	wire _w12424_ ;
	wire _w12423_ ;
	wire _w12422_ ;
	wire _w12421_ ;
	wire _w12420_ ;
	wire _w12419_ ;
	wire _w12418_ ;
	wire _w12417_ ;
	wire _w12416_ ;
	wire _w12415_ ;
	wire _w12414_ ;
	wire _w12413_ ;
	wire _w12412_ ;
	wire _w12411_ ;
	wire _w12410_ ;
	wire _w12409_ ;
	wire _w12408_ ;
	wire _w12407_ ;
	wire _w12406_ ;
	wire _w12405_ ;
	wire _w12404_ ;
	wire _w12403_ ;
	wire _w12402_ ;
	wire _w12401_ ;
	wire _w12400_ ;
	wire _w12399_ ;
	wire _w12398_ ;
	wire _w12397_ ;
	wire _w12396_ ;
	wire _w12395_ ;
	wire _w12394_ ;
	wire _w12393_ ;
	wire _w12392_ ;
	wire _w12391_ ;
	wire _w12390_ ;
	wire _w12389_ ;
	wire _w12388_ ;
	wire _w12387_ ;
	wire _w12386_ ;
	wire _w12385_ ;
	wire _w12384_ ;
	wire _w12383_ ;
	wire _w12382_ ;
	wire _w12381_ ;
	wire _w12380_ ;
	wire _w12379_ ;
	wire _w12378_ ;
	wire _w12377_ ;
	wire _w12376_ ;
	wire _w12375_ ;
	wire _w12374_ ;
	wire _w12373_ ;
	wire _w12372_ ;
	wire _w12371_ ;
	wire _w12370_ ;
	wire _w12369_ ;
	wire _w12368_ ;
	wire _w12367_ ;
	wire _w12366_ ;
	wire _w12365_ ;
	wire _w12364_ ;
	wire _w12363_ ;
	wire _w12362_ ;
	wire _w12361_ ;
	wire _w12360_ ;
	wire _w12359_ ;
	wire _w12358_ ;
	wire _w12357_ ;
	wire _w12356_ ;
	wire _w12355_ ;
	wire _w12354_ ;
	wire _w12353_ ;
	wire _w12352_ ;
	wire _w12351_ ;
	wire _w12350_ ;
	wire _w12349_ ;
	wire _w12348_ ;
	wire _w12347_ ;
	wire _w12346_ ;
	wire _w12345_ ;
	wire _w12344_ ;
	wire _w12343_ ;
	wire _w12342_ ;
	wire _w12341_ ;
	wire _w12340_ ;
	wire _w12339_ ;
	wire _w12338_ ;
	wire _w12337_ ;
	wire _w12336_ ;
	wire _w12335_ ;
	wire _w12334_ ;
	wire _w12333_ ;
	wire _w12332_ ;
	wire _w12331_ ;
	wire _w12330_ ;
	wire _w12329_ ;
	wire _w12328_ ;
	wire _w12327_ ;
	wire _w12326_ ;
	wire _w12325_ ;
	wire _w12324_ ;
	wire _w12323_ ;
	wire _w12322_ ;
	wire _w12321_ ;
	wire _w12320_ ;
	wire _w12319_ ;
	wire _w12318_ ;
	wire _w12317_ ;
	wire _w12316_ ;
	wire _w12315_ ;
	wire _w12314_ ;
	wire _w12313_ ;
	wire _w12312_ ;
	wire _w12311_ ;
	wire _w12310_ ;
	wire _w12309_ ;
	wire _w12308_ ;
	wire _w12307_ ;
	wire _w12306_ ;
	wire _w12305_ ;
	wire _w12304_ ;
	wire _w12303_ ;
	wire _w12302_ ;
	wire _w12301_ ;
	wire _w12300_ ;
	wire _w12299_ ;
	wire _w12298_ ;
	wire _w12297_ ;
	wire _w12296_ ;
	wire _w12295_ ;
	wire _w12294_ ;
	wire _w12293_ ;
	wire _w12292_ ;
	wire _w12291_ ;
	wire _w12290_ ;
	wire _w12289_ ;
	wire _w12288_ ;
	wire _w12287_ ;
	wire _w12286_ ;
	wire _w12285_ ;
	wire _w12284_ ;
	wire _w12283_ ;
	wire _w12282_ ;
	wire _w12281_ ;
	wire _w12280_ ;
	wire _w12279_ ;
	wire _w12278_ ;
	wire _w12277_ ;
	wire _w12276_ ;
	wire _w12275_ ;
	wire _w12274_ ;
	wire _w12273_ ;
	wire _w12272_ ;
	wire _w12271_ ;
	wire _w12270_ ;
	wire _w12269_ ;
	wire _w12268_ ;
	wire _w12267_ ;
	wire _w12266_ ;
	wire _w12265_ ;
	wire _w12264_ ;
	wire _w12263_ ;
	wire _w12262_ ;
	wire _w12261_ ;
	wire _w12260_ ;
	wire _w12259_ ;
	wire _w12258_ ;
	wire _w12257_ ;
	wire _w12256_ ;
	wire _w12255_ ;
	wire _w12254_ ;
	wire _w12253_ ;
	wire _w12252_ ;
	wire _w12251_ ;
	wire _w12250_ ;
	wire _w12249_ ;
	wire _w12248_ ;
	wire _w12247_ ;
	wire _w12246_ ;
	wire _w12245_ ;
	wire _w12244_ ;
	wire _w12243_ ;
	wire _w12242_ ;
	wire _w12241_ ;
	wire _w12240_ ;
	wire _w12239_ ;
	wire _w12238_ ;
	wire _w12237_ ;
	wire _w12236_ ;
	wire _w12235_ ;
	wire _w12234_ ;
	wire _w12233_ ;
	wire _w12232_ ;
	wire _w12231_ ;
	wire _w12230_ ;
	wire _w12229_ ;
	wire _w12228_ ;
	wire _w12227_ ;
	wire _w12226_ ;
	wire _w12225_ ;
	wire _w12224_ ;
	wire _w12223_ ;
	wire _w12222_ ;
	wire _w12221_ ;
	wire _w12220_ ;
	wire _w12219_ ;
	wire _w12218_ ;
	wire _w12217_ ;
	wire _w12216_ ;
	wire _w12215_ ;
	wire _w12214_ ;
	wire _w12213_ ;
	wire _w12212_ ;
	wire _w12211_ ;
	wire _w12210_ ;
	wire _w12209_ ;
	wire _w12208_ ;
	wire _w12207_ ;
	wire _w12206_ ;
	wire _w12205_ ;
	wire _w12204_ ;
	wire _w12203_ ;
	wire _w12202_ ;
	wire _w12201_ ;
	wire _w12200_ ;
	wire _w12199_ ;
	wire _w12198_ ;
	wire _w12197_ ;
	wire _w12196_ ;
	wire _w12195_ ;
	wire _w12194_ ;
	wire _w12193_ ;
	wire _w12192_ ;
	wire _w12191_ ;
	wire _w12190_ ;
	wire _w12189_ ;
	wire _w12188_ ;
	wire _w12187_ ;
	wire _w12186_ ;
	wire _w12185_ ;
	wire _w12184_ ;
	wire _w12183_ ;
	wire _w12182_ ;
	wire _w12181_ ;
	wire _w12180_ ;
	wire _w12179_ ;
	wire _w12178_ ;
	wire _w12177_ ;
	wire _w12176_ ;
	wire _w12175_ ;
	wire _w12174_ ;
	wire _w12173_ ;
	wire _w12172_ ;
	wire _w12171_ ;
	wire _w12170_ ;
	wire _w12169_ ;
	wire _w12168_ ;
	wire _w12167_ ;
	wire _w12166_ ;
	wire _w12165_ ;
	wire _w12164_ ;
	wire _w12163_ ;
	wire _w12162_ ;
	wire _w12161_ ;
	wire _w12160_ ;
	wire _w12159_ ;
	wire _w12158_ ;
	wire _w12157_ ;
	wire _w12156_ ;
	wire _w12155_ ;
	wire _w12154_ ;
	wire _w12153_ ;
	wire _w12152_ ;
	wire _w12151_ ;
	wire _w12150_ ;
	wire _w12149_ ;
	wire _w12148_ ;
	wire _w12147_ ;
	wire _w12146_ ;
	wire _w12145_ ;
	wire _w12144_ ;
	wire _w12143_ ;
	wire _w12142_ ;
	wire _w12141_ ;
	wire _w12140_ ;
	wire _w12139_ ;
	wire _w12138_ ;
	wire _w12137_ ;
	wire _w12136_ ;
	wire _w12135_ ;
	wire _w12134_ ;
	wire _w12133_ ;
	wire _w12132_ ;
	wire _w12131_ ;
	wire _w12130_ ;
	wire _w12129_ ;
	wire _w12128_ ;
	wire _w12127_ ;
	wire _w12126_ ;
	wire _w12125_ ;
	wire _w12124_ ;
	wire _w12123_ ;
	wire _w12122_ ;
	wire _w12121_ ;
	wire _w12120_ ;
	wire _w12119_ ;
	wire _w12118_ ;
	wire _w12117_ ;
	wire _w12116_ ;
	wire _w12115_ ;
	wire _w12114_ ;
	wire _w12113_ ;
	wire _w12112_ ;
	wire _w12111_ ;
	wire _w12110_ ;
	wire _w12109_ ;
	wire _w12108_ ;
	wire _w12107_ ;
	wire _w12106_ ;
	wire _w12105_ ;
	wire _w12104_ ;
	wire _w12103_ ;
	wire _w12102_ ;
	wire _w12101_ ;
	wire _w12100_ ;
	wire _w12099_ ;
	wire _w12098_ ;
	wire _w12097_ ;
	wire _w12096_ ;
	wire _w12095_ ;
	wire _w12094_ ;
	wire _w12093_ ;
	wire _w12092_ ;
	wire _w12091_ ;
	wire _w12090_ ;
	wire _w12089_ ;
	wire _w12088_ ;
	wire _w12087_ ;
	wire _w12086_ ;
	wire _w12085_ ;
	wire _w12084_ ;
	wire _w12083_ ;
	wire _w12082_ ;
	wire _w12081_ ;
	wire _w12080_ ;
	wire _w12079_ ;
	wire _w12078_ ;
	wire _w12077_ ;
	wire _w12076_ ;
	wire _w12075_ ;
	wire _w12074_ ;
	wire _w12073_ ;
	wire _w12072_ ;
	wire _w12071_ ;
	wire _w12070_ ;
	wire _w12069_ ;
	wire _w12068_ ;
	wire _w12067_ ;
	wire _w12066_ ;
	wire _w12065_ ;
	wire _w12064_ ;
	wire _w12063_ ;
	wire _w12062_ ;
	wire _w12061_ ;
	wire _w12060_ ;
	wire _w12059_ ;
	wire _w12058_ ;
	wire _w12057_ ;
	wire _w12056_ ;
	wire _w12055_ ;
	wire _w12054_ ;
	wire _w12053_ ;
	wire _w12052_ ;
	wire _w12051_ ;
	wire _w12050_ ;
	wire _w12049_ ;
	wire _w12048_ ;
	wire _w12047_ ;
	wire _w12046_ ;
	wire _w12045_ ;
	wire _w12044_ ;
	wire _w12043_ ;
	wire _w12042_ ;
	wire _w12041_ ;
	wire _w12040_ ;
	wire _w12039_ ;
	wire _w12038_ ;
	wire _w12037_ ;
	wire _w12036_ ;
	wire _w12035_ ;
	wire _w12034_ ;
	wire _w12033_ ;
	wire _w12032_ ;
	wire _w12031_ ;
	wire _w12030_ ;
	wire _w12029_ ;
	wire _w12028_ ;
	wire _w12027_ ;
	wire _w12026_ ;
	wire _w12025_ ;
	wire _w12024_ ;
	wire _w12023_ ;
	wire _w12022_ ;
	wire _w12021_ ;
	wire _w12020_ ;
	wire _w12019_ ;
	wire _w12018_ ;
	wire _w12017_ ;
	wire _w12016_ ;
	wire _w12015_ ;
	wire _w12014_ ;
	wire _w12013_ ;
	wire _w12012_ ;
	wire _w12011_ ;
	wire _w12010_ ;
	wire _w12009_ ;
	wire _w12008_ ;
	wire _w12007_ ;
	wire _w12006_ ;
	wire _w12005_ ;
	wire _w12004_ ;
	wire _w12003_ ;
	wire _w12002_ ;
	wire _w12001_ ;
	wire _w12000_ ;
	wire _w11999_ ;
	wire _w11998_ ;
	wire _w11997_ ;
	wire _w11996_ ;
	wire _w11995_ ;
	wire _w11994_ ;
	wire _w11993_ ;
	wire _w11992_ ;
	wire _w11991_ ;
	wire _w11990_ ;
	wire _w11989_ ;
	wire _w11988_ ;
	wire _w11987_ ;
	wire _w11986_ ;
	wire _w11985_ ;
	wire _w11984_ ;
	wire _w11983_ ;
	wire _w11982_ ;
	wire _w11981_ ;
	wire _w11980_ ;
	wire _w11979_ ;
	wire _w11978_ ;
	wire _w11977_ ;
	wire _w11976_ ;
	wire _w11975_ ;
	wire _w11974_ ;
	wire _w11973_ ;
	wire _w11972_ ;
	wire _w11971_ ;
	wire _w11970_ ;
	wire _w11969_ ;
	wire _w11968_ ;
	wire _w11967_ ;
	wire _w11966_ ;
	wire _w11965_ ;
	wire _w11964_ ;
	wire _w11963_ ;
	wire _w11962_ ;
	wire _w11961_ ;
	wire _w11960_ ;
	wire _w11959_ ;
	wire _w11958_ ;
	wire _w11957_ ;
	wire _w11956_ ;
	wire _w11955_ ;
	wire _w11954_ ;
	wire _w11953_ ;
	wire _w11952_ ;
	wire _w11951_ ;
	wire _w11950_ ;
	wire _w11949_ ;
	wire _w11948_ ;
	wire _w11947_ ;
	wire _w11946_ ;
	wire _w11945_ ;
	wire _w11944_ ;
	wire _w11943_ ;
	wire _w11942_ ;
	wire _w11941_ ;
	wire _w11940_ ;
	wire _w11939_ ;
	wire _w11938_ ;
	wire _w11937_ ;
	wire _w11936_ ;
	wire _w11935_ ;
	wire _w11934_ ;
	wire _w11933_ ;
	wire _w11932_ ;
	wire _w11931_ ;
	wire _w11930_ ;
	wire _w11929_ ;
	wire _w11928_ ;
	wire _w11927_ ;
	wire _w11926_ ;
	wire _w11925_ ;
	wire _w11924_ ;
	wire _w11923_ ;
	wire _w11922_ ;
	wire _w11921_ ;
	wire _w11920_ ;
	wire _w11919_ ;
	wire _w11918_ ;
	wire _w11917_ ;
	wire _w11916_ ;
	wire _w11915_ ;
	wire _w11914_ ;
	wire _w11913_ ;
	wire _w11912_ ;
	wire _w11911_ ;
	wire _w11910_ ;
	wire _w11909_ ;
	wire _w11908_ ;
	wire _w11907_ ;
	wire _w11906_ ;
	wire _w11905_ ;
	wire _w11904_ ;
	wire _w11903_ ;
	wire _w11902_ ;
	wire _w11901_ ;
	wire _w11900_ ;
	wire _w11899_ ;
	wire _w11898_ ;
	wire _w11897_ ;
	wire _w11896_ ;
	wire _w11895_ ;
	wire _w11894_ ;
	wire _w11893_ ;
	wire _w11892_ ;
	wire _w11891_ ;
	wire _w11890_ ;
	wire _w11889_ ;
	wire _w11888_ ;
	wire _w11887_ ;
	wire _w11886_ ;
	wire _w11885_ ;
	wire _w11884_ ;
	wire _w11883_ ;
	wire _w11882_ ;
	wire _w11881_ ;
	wire _w11880_ ;
	wire _w11879_ ;
	wire _w11878_ ;
	wire _w11877_ ;
	wire _w11876_ ;
	wire _w11875_ ;
	wire _w11874_ ;
	wire _w11873_ ;
	wire _w11872_ ;
	wire _w11871_ ;
	wire _w11870_ ;
	wire _w11869_ ;
	wire _w11868_ ;
	wire _w11867_ ;
	wire _w11866_ ;
	wire _w11865_ ;
	wire _w11864_ ;
	wire _w11863_ ;
	wire _w11862_ ;
	wire _w11861_ ;
	wire _w11860_ ;
	wire _w11859_ ;
	wire _w11858_ ;
	wire _w11857_ ;
	wire _w11856_ ;
	wire _w11855_ ;
	wire _w11854_ ;
	wire _w11853_ ;
	wire _w11852_ ;
	wire _w11851_ ;
	wire _w11850_ ;
	wire _w11849_ ;
	wire _w11848_ ;
	wire _w11847_ ;
	wire _w11846_ ;
	wire _w11845_ ;
	wire _w11844_ ;
	wire _w11843_ ;
	wire _w11842_ ;
	wire _w11841_ ;
	wire _w11840_ ;
	wire _w11839_ ;
	wire _w11838_ ;
	wire _w11837_ ;
	wire _w11836_ ;
	wire _w11835_ ;
	wire _w11834_ ;
	wire _w11833_ ;
	wire _w11832_ ;
	wire _w11831_ ;
	wire _w11830_ ;
	wire _w11829_ ;
	wire _w11828_ ;
	wire _w11827_ ;
	wire _w11826_ ;
	wire _w11825_ ;
	wire _w11824_ ;
	wire _w11823_ ;
	wire _w11822_ ;
	wire _w11821_ ;
	wire _w11820_ ;
	wire _w11819_ ;
	wire _w11818_ ;
	wire _w11817_ ;
	wire _w11816_ ;
	wire _w11815_ ;
	wire _w11814_ ;
	wire _w11813_ ;
	wire _w11812_ ;
	wire _w11811_ ;
	wire _w11810_ ;
	wire _w11809_ ;
	wire _w11808_ ;
	wire _w11807_ ;
	wire _w11806_ ;
	wire _w11805_ ;
	wire _w11804_ ;
	wire _w11803_ ;
	wire _w11802_ ;
	wire _w11801_ ;
	wire _w11800_ ;
	wire _w11799_ ;
	wire _w11798_ ;
	wire _w11797_ ;
	wire _w11796_ ;
	wire _w11795_ ;
	wire _w11794_ ;
	wire _w11793_ ;
	wire _w11792_ ;
	wire _w11791_ ;
	wire _w11790_ ;
	wire _w11789_ ;
	wire _w11788_ ;
	wire _w11787_ ;
	wire _w11786_ ;
	wire _w11785_ ;
	wire _w11784_ ;
	wire _w11783_ ;
	wire _w11782_ ;
	wire _w11781_ ;
	wire _w11780_ ;
	wire _w11779_ ;
	wire _w11778_ ;
	wire _w11777_ ;
	wire _w11776_ ;
	wire _w11775_ ;
	wire _w11774_ ;
	wire _w11773_ ;
	wire _w11772_ ;
	wire _w11771_ ;
	wire _w11770_ ;
	wire _w11769_ ;
	wire _w11768_ ;
	wire _w11767_ ;
	wire _w11766_ ;
	wire _w11765_ ;
	wire _w11764_ ;
	wire _w11763_ ;
	wire _w11762_ ;
	wire _w11761_ ;
	wire _w11760_ ;
	wire _w11759_ ;
	wire _w11758_ ;
	wire _w11757_ ;
	wire _w11756_ ;
	wire _w11755_ ;
	wire _w11754_ ;
	wire _w11753_ ;
	wire _w11752_ ;
	wire _w11751_ ;
	wire _w11750_ ;
	wire _w11749_ ;
	wire _w11748_ ;
	wire _w11747_ ;
	wire _w11746_ ;
	wire _w11745_ ;
	wire _w11744_ ;
	wire _w11743_ ;
	wire _w11742_ ;
	wire _w11741_ ;
	wire _w11740_ ;
	wire _w11739_ ;
	wire _w11738_ ;
	wire _w11737_ ;
	wire _w11736_ ;
	wire _w11735_ ;
	wire _w11734_ ;
	wire _w11733_ ;
	wire _w11732_ ;
	wire _w11731_ ;
	wire _w11730_ ;
	wire _w11729_ ;
	wire _w11728_ ;
	wire _w11727_ ;
	wire _w11726_ ;
	wire _w11725_ ;
	wire _w11724_ ;
	wire _w11723_ ;
	wire _w11722_ ;
	wire _w11721_ ;
	wire _w11720_ ;
	wire _w11719_ ;
	wire _w11718_ ;
	wire _w11717_ ;
	wire _w11716_ ;
	wire _w11715_ ;
	wire _w11714_ ;
	wire _w11713_ ;
	wire _w11712_ ;
	wire _w11711_ ;
	wire _w11710_ ;
	wire _w11709_ ;
	wire _w11708_ ;
	wire _w11707_ ;
	wire _w11706_ ;
	wire _w11705_ ;
	wire _w11704_ ;
	wire _w11703_ ;
	wire _w11702_ ;
	wire _w11701_ ;
	wire _w11700_ ;
	wire _w11699_ ;
	wire _w11698_ ;
	wire _w11697_ ;
	wire _w11696_ ;
	wire _w11695_ ;
	wire _w11694_ ;
	wire _w11693_ ;
	wire _w11692_ ;
	wire _w11691_ ;
	wire _w11690_ ;
	wire _w11689_ ;
	wire _w11688_ ;
	wire _w11687_ ;
	wire _w11686_ ;
	wire _w11685_ ;
	wire _w11684_ ;
	wire _w11683_ ;
	wire _w11682_ ;
	wire _w11681_ ;
	wire _w11680_ ;
	wire _w11679_ ;
	wire _w11678_ ;
	wire _w11677_ ;
	wire _w11676_ ;
	wire _w11675_ ;
	wire _w11674_ ;
	wire _w11673_ ;
	wire _w11672_ ;
	wire _w11671_ ;
	wire _w11670_ ;
	wire _w11669_ ;
	wire _w11668_ ;
	wire _w11667_ ;
	wire _w11666_ ;
	wire _w11665_ ;
	wire _w11664_ ;
	wire _w11663_ ;
	wire _w11662_ ;
	wire _w11661_ ;
	wire _w11660_ ;
	wire _w11659_ ;
	wire _w11658_ ;
	wire _w11657_ ;
	wire _w11656_ ;
	wire _w11655_ ;
	wire _w11654_ ;
	wire _w11653_ ;
	wire _w11652_ ;
	wire _w11651_ ;
	wire _w11650_ ;
	wire _w11649_ ;
	wire _w11648_ ;
	wire _w11647_ ;
	wire _w11646_ ;
	wire _w11645_ ;
	wire _w11644_ ;
	wire _w11643_ ;
	wire _w11642_ ;
	wire _w11641_ ;
	wire _w11640_ ;
	wire _w11639_ ;
	wire _w11638_ ;
	wire _w11637_ ;
	wire _w11636_ ;
	wire _w11635_ ;
	wire _w11634_ ;
	wire _w11633_ ;
	wire _w11632_ ;
	wire _w11631_ ;
	wire _w11630_ ;
	wire _w11629_ ;
	wire _w11628_ ;
	wire _w11627_ ;
	wire _w11626_ ;
	wire _w11625_ ;
	wire _w11624_ ;
	wire _w11623_ ;
	wire _w11622_ ;
	wire _w11621_ ;
	wire _w11620_ ;
	wire _w11619_ ;
	wire _w11618_ ;
	wire _w11617_ ;
	wire _w11616_ ;
	wire _w11615_ ;
	wire _w11614_ ;
	wire _w11613_ ;
	wire _w11612_ ;
	wire _w11611_ ;
	wire _w11610_ ;
	wire _w11609_ ;
	wire _w11608_ ;
	wire _w11607_ ;
	wire _w11606_ ;
	wire _w11605_ ;
	wire _w11604_ ;
	wire _w11603_ ;
	wire _w11602_ ;
	wire _w11601_ ;
	wire _w11600_ ;
	wire _w11599_ ;
	wire _w11598_ ;
	wire _w11597_ ;
	wire _w11596_ ;
	wire _w11595_ ;
	wire _w11594_ ;
	wire _w11593_ ;
	wire _w11592_ ;
	wire _w11591_ ;
	wire _w11590_ ;
	wire _w11589_ ;
	wire _w11588_ ;
	wire _w11587_ ;
	wire _w11586_ ;
	wire _w11585_ ;
	wire _w11584_ ;
	wire _w11583_ ;
	wire _w11582_ ;
	wire _w11581_ ;
	wire _w11580_ ;
	wire _w11579_ ;
	wire _w11578_ ;
	wire _w11577_ ;
	wire _w11576_ ;
	wire _w11575_ ;
	wire _w11574_ ;
	wire _w11573_ ;
	wire _w11572_ ;
	wire _w11571_ ;
	wire _w11570_ ;
	wire _w11569_ ;
	wire _w11568_ ;
	wire _w11567_ ;
	wire _w11566_ ;
	wire _w11565_ ;
	wire _w11564_ ;
	wire _w11563_ ;
	wire _w11562_ ;
	wire _w11561_ ;
	wire _w11560_ ;
	wire _w11559_ ;
	wire _w11558_ ;
	wire _w11557_ ;
	wire _w11556_ ;
	wire _w11555_ ;
	wire _w11554_ ;
	wire _w11553_ ;
	wire _w11552_ ;
	wire _w11551_ ;
	wire _w11550_ ;
	wire _w11549_ ;
	wire _w11548_ ;
	wire _w11547_ ;
	wire _w11546_ ;
	wire _w11545_ ;
	wire _w11544_ ;
	wire _w11543_ ;
	wire _w11542_ ;
	wire _w11541_ ;
	wire _w11540_ ;
	wire _w11539_ ;
	wire _w11538_ ;
	wire _w11537_ ;
	wire _w11536_ ;
	wire _w11535_ ;
	wire _w11534_ ;
	wire _w11533_ ;
	wire _w11532_ ;
	wire _w11531_ ;
	wire _w11530_ ;
	wire _w11529_ ;
	wire _w11528_ ;
	wire _w11527_ ;
	wire _w11526_ ;
	wire _w11525_ ;
	wire _w11524_ ;
	wire _w11523_ ;
	wire _w11522_ ;
	wire _w11521_ ;
	wire _w11520_ ;
	wire _w11519_ ;
	wire _w11518_ ;
	wire _w11517_ ;
	wire _w11516_ ;
	wire _w11515_ ;
	wire _w11514_ ;
	wire _w11513_ ;
	wire _w11512_ ;
	wire _w11511_ ;
	wire _w11510_ ;
	wire _w11509_ ;
	wire _w11508_ ;
	wire _w11507_ ;
	wire _w11506_ ;
	wire _w11505_ ;
	wire _w11504_ ;
	wire _w11503_ ;
	wire _w11502_ ;
	wire _w11501_ ;
	wire _w11500_ ;
	wire _w11499_ ;
	wire _w11498_ ;
	wire _w11497_ ;
	wire _w11496_ ;
	wire _w11495_ ;
	wire _w11494_ ;
	wire _w11493_ ;
	wire _w11492_ ;
	wire _w11491_ ;
	wire _w11490_ ;
	wire _w11489_ ;
	wire _w11488_ ;
	wire _w11487_ ;
	wire _w11486_ ;
	wire _w11485_ ;
	wire _w11484_ ;
	wire _w11483_ ;
	wire _w11482_ ;
	wire _w11481_ ;
	wire _w11480_ ;
	wire _w11479_ ;
	wire _w11478_ ;
	wire _w11477_ ;
	wire _w11476_ ;
	wire _w11475_ ;
	wire _w11474_ ;
	wire _w11473_ ;
	wire _w11472_ ;
	wire _w11471_ ;
	wire _w11470_ ;
	wire _w11469_ ;
	wire _w11468_ ;
	wire _w11467_ ;
	wire _w11466_ ;
	wire _w11465_ ;
	wire _w11464_ ;
	wire _w11463_ ;
	wire _w11462_ ;
	wire _w11461_ ;
	wire _w11460_ ;
	wire _w11459_ ;
	wire _w11458_ ;
	wire _w11457_ ;
	wire _w11456_ ;
	wire _w11455_ ;
	wire _w11454_ ;
	wire _w11453_ ;
	wire _w11452_ ;
	wire _w11451_ ;
	wire _w11450_ ;
	wire _w11449_ ;
	wire _w11448_ ;
	wire _w11447_ ;
	wire _w11446_ ;
	wire _w11445_ ;
	wire _w11444_ ;
	wire _w11443_ ;
	wire _w11442_ ;
	wire _w11441_ ;
	wire _w11440_ ;
	wire _w11439_ ;
	wire _w11438_ ;
	wire _w11437_ ;
	wire _w11436_ ;
	wire _w11435_ ;
	wire _w11434_ ;
	wire _w11433_ ;
	wire _w11432_ ;
	wire _w11431_ ;
	wire _w11430_ ;
	wire _w11429_ ;
	wire _w11428_ ;
	wire _w11427_ ;
	wire _w11426_ ;
	wire _w11425_ ;
	wire _w11424_ ;
	wire _w11423_ ;
	wire _w11422_ ;
	wire _w11421_ ;
	wire _w11420_ ;
	wire _w11419_ ;
	wire _w11418_ ;
	wire _w11417_ ;
	wire _w11416_ ;
	wire _w11415_ ;
	wire _w11414_ ;
	wire _w11413_ ;
	wire _w11412_ ;
	wire _w11411_ ;
	wire _w11410_ ;
	wire _w11409_ ;
	wire _w11408_ ;
	wire _w11407_ ;
	wire _w11406_ ;
	wire _w11405_ ;
	wire _w11404_ ;
	wire _w11403_ ;
	wire _w11402_ ;
	wire _w11401_ ;
	wire _w11400_ ;
	wire _w11399_ ;
	wire _w11398_ ;
	wire _w11397_ ;
	wire _w11396_ ;
	wire _w11395_ ;
	wire _w11394_ ;
	wire _w11393_ ;
	wire _w11392_ ;
	wire _w11391_ ;
	wire _w11390_ ;
	wire _w11389_ ;
	wire _w11388_ ;
	wire _w11387_ ;
	wire _w11386_ ;
	wire _w11385_ ;
	wire _w11384_ ;
	wire _w11383_ ;
	wire _w11382_ ;
	wire _w11381_ ;
	wire _w11380_ ;
	wire _w11379_ ;
	wire _w11378_ ;
	wire _w11377_ ;
	wire _w11376_ ;
	wire _w11375_ ;
	wire _w11374_ ;
	wire _w11373_ ;
	wire _w11372_ ;
	wire _w11371_ ;
	wire _w11370_ ;
	wire _w11369_ ;
	wire _w11368_ ;
	wire _w11367_ ;
	wire _w11366_ ;
	wire _w11365_ ;
	wire _w11364_ ;
	wire _w11363_ ;
	wire _w11362_ ;
	wire _w11361_ ;
	wire _w11360_ ;
	wire _w11359_ ;
	wire _w11358_ ;
	wire _w11357_ ;
	wire _w11356_ ;
	wire _w11355_ ;
	wire _w11354_ ;
	wire _w11353_ ;
	wire _w11352_ ;
	wire _w11351_ ;
	wire _w11350_ ;
	wire _w11349_ ;
	wire _w11348_ ;
	wire _w11347_ ;
	wire _w11346_ ;
	wire _w11345_ ;
	wire _w11344_ ;
	wire _w11343_ ;
	wire _w11342_ ;
	wire _w11341_ ;
	wire _w11340_ ;
	wire _w11339_ ;
	wire _w11338_ ;
	wire _w11337_ ;
	wire _w11336_ ;
	wire _w11335_ ;
	wire _w11334_ ;
	wire _w11333_ ;
	wire _w11332_ ;
	wire _w11331_ ;
	wire _w11330_ ;
	wire _w11329_ ;
	wire _w11328_ ;
	wire _w11327_ ;
	wire _w11326_ ;
	wire _w11325_ ;
	wire _w11324_ ;
	wire _w11323_ ;
	wire _w11322_ ;
	wire _w11321_ ;
	wire _w11320_ ;
	wire _w11319_ ;
	wire _w11318_ ;
	wire _w11317_ ;
	wire _w11316_ ;
	wire _w11315_ ;
	wire _w11314_ ;
	wire _w11313_ ;
	wire _w11312_ ;
	wire _w11311_ ;
	wire _w11310_ ;
	wire _w11309_ ;
	wire _w11308_ ;
	wire _w11307_ ;
	wire _w11306_ ;
	wire _w11305_ ;
	wire _w11304_ ;
	wire _w11303_ ;
	wire _w11302_ ;
	wire _w11301_ ;
	wire _w11300_ ;
	wire _w11299_ ;
	wire _w11298_ ;
	wire _w11297_ ;
	wire _w11296_ ;
	wire _w11295_ ;
	wire _w11294_ ;
	wire _w11293_ ;
	wire _w11292_ ;
	wire _w11291_ ;
	wire _w11290_ ;
	wire _w11289_ ;
	wire _w11288_ ;
	wire _w11287_ ;
	wire _w11286_ ;
	wire _w11285_ ;
	wire _w11284_ ;
	wire _w11283_ ;
	wire _w11282_ ;
	wire _w11281_ ;
	wire _w11280_ ;
	wire _w11279_ ;
	wire _w11278_ ;
	wire _w11277_ ;
	wire _w11276_ ;
	wire _w11275_ ;
	wire _w11274_ ;
	wire _w11273_ ;
	wire _w11272_ ;
	wire _w11271_ ;
	wire _w11270_ ;
	wire _w11269_ ;
	wire _w11268_ ;
	wire _w11267_ ;
	wire _w11266_ ;
	wire _w11265_ ;
	wire _w11264_ ;
	wire _w11263_ ;
	wire _w11262_ ;
	wire _w11261_ ;
	wire _w11260_ ;
	wire _w11259_ ;
	wire _w11258_ ;
	wire _w11257_ ;
	wire _w11256_ ;
	wire _w11255_ ;
	wire _w11254_ ;
	wire _w11253_ ;
	wire _w11252_ ;
	wire _w11251_ ;
	wire _w11250_ ;
	wire _w11249_ ;
	wire _w11248_ ;
	wire _w11247_ ;
	wire _w11246_ ;
	wire _w11245_ ;
	wire _w11244_ ;
	wire _w11243_ ;
	wire _w11242_ ;
	wire _w11241_ ;
	wire _w11240_ ;
	wire _w11239_ ;
	wire _w11238_ ;
	wire _w11237_ ;
	wire _w11236_ ;
	wire _w11235_ ;
	wire _w11234_ ;
	wire _w11233_ ;
	wire _w11232_ ;
	wire _w11231_ ;
	wire _w11230_ ;
	wire _w11229_ ;
	wire _w11228_ ;
	wire _w11227_ ;
	wire _w11226_ ;
	wire _w11225_ ;
	wire _w11224_ ;
	wire _w11223_ ;
	wire _w11222_ ;
	wire _w11221_ ;
	wire _w11220_ ;
	wire _w11219_ ;
	wire _w11218_ ;
	wire _w11217_ ;
	wire _w11216_ ;
	wire _w11215_ ;
	wire _w11214_ ;
	wire _w11213_ ;
	wire _w11212_ ;
	wire _w11211_ ;
	wire _w11210_ ;
	wire _w11209_ ;
	wire _w11208_ ;
	wire _w11207_ ;
	wire _w11206_ ;
	wire _w11205_ ;
	wire _w11204_ ;
	wire _w11203_ ;
	wire _w11202_ ;
	wire _w11201_ ;
	wire _w11200_ ;
	wire _w11199_ ;
	wire _w11198_ ;
	wire _w11197_ ;
	wire _w11196_ ;
	wire _w11195_ ;
	wire _w11194_ ;
	wire _w11193_ ;
	wire _w11192_ ;
	wire _w11191_ ;
	wire _w11190_ ;
	wire _w11189_ ;
	wire _w11188_ ;
	wire _w11187_ ;
	wire _w11186_ ;
	wire _w11185_ ;
	wire _w11184_ ;
	wire _w11183_ ;
	wire _w11182_ ;
	wire _w11181_ ;
	wire _w11180_ ;
	wire _w11179_ ;
	wire _w11178_ ;
	wire _w11177_ ;
	wire _w11176_ ;
	wire _w11175_ ;
	wire _w11174_ ;
	wire _w11173_ ;
	wire _w11172_ ;
	wire _w11171_ ;
	wire _w11170_ ;
	wire _w11169_ ;
	wire _w11168_ ;
	wire _w11167_ ;
	wire _w11166_ ;
	wire _w11165_ ;
	wire _w11164_ ;
	wire _w11163_ ;
	wire _w11162_ ;
	wire _w11161_ ;
	wire _w11160_ ;
	wire _w11159_ ;
	wire _w11158_ ;
	wire _w11157_ ;
	wire _w11156_ ;
	wire _w11155_ ;
	wire _w11154_ ;
	wire _w11153_ ;
	wire _w11152_ ;
	wire _w11151_ ;
	wire _w11150_ ;
	wire _w11149_ ;
	wire _w11148_ ;
	wire _w11147_ ;
	wire _w11146_ ;
	wire _w11145_ ;
	wire _w11144_ ;
	wire _w11143_ ;
	wire _w11142_ ;
	wire _w11141_ ;
	wire _w11140_ ;
	wire _w11139_ ;
	wire _w11138_ ;
	wire _w11137_ ;
	wire _w11136_ ;
	wire _w11135_ ;
	wire _w11134_ ;
	wire _w11133_ ;
	wire _w11132_ ;
	wire _w11131_ ;
	wire _w11130_ ;
	wire _w11129_ ;
	wire _w11128_ ;
	wire _w11127_ ;
	wire _w11126_ ;
	wire _w11125_ ;
	wire _w11124_ ;
	wire _w11123_ ;
	wire _w11122_ ;
	wire _w11121_ ;
	wire _w11120_ ;
	wire _w11119_ ;
	wire _w11118_ ;
	wire _w11117_ ;
	wire _w11116_ ;
	wire _w11115_ ;
	wire _w11114_ ;
	wire _w11113_ ;
	wire _w11112_ ;
	wire _w11111_ ;
	wire _w11110_ ;
	wire _w11109_ ;
	wire _w11108_ ;
	wire _w11107_ ;
	wire _w11106_ ;
	wire _w11105_ ;
	wire _w11104_ ;
	wire _w11103_ ;
	wire _w11102_ ;
	wire _w11101_ ;
	wire _w11100_ ;
	wire _w11099_ ;
	wire _w11098_ ;
	wire _w11097_ ;
	wire _w11096_ ;
	wire _w11095_ ;
	wire _w11094_ ;
	wire _w11093_ ;
	wire _w11092_ ;
	wire _w11091_ ;
	wire _w11090_ ;
	wire _w11089_ ;
	wire _w11088_ ;
	wire _w11087_ ;
	wire _w11086_ ;
	wire _w11085_ ;
	wire _w11084_ ;
	wire _w11083_ ;
	wire _w11082_ ;
	wire _w11081_ ;
	wire _w11080_ ;
	wire _w11079_ ;
	wire _w11078_ ;
	wire _w11077_ ;
	wire _w11076_ ;
	wire _w11075_ ;
	wire _w11074_ ;
	wire _w11073_ ;
	wire _w11072_ ;
	wire _w11071_ ;
	wire _w11070_ ;
	wire _w11069_ ;
	wire _w11068_ ;
	wire _w11067_ ;
	wire _w11066_ ;
	wire _w11065_ ;
	wire _w11064_ ;
	wire _w11063_ ;
	wire _w11062_ ;
	wire _w11061_ ;
	wire _w11060_ ;
	wire _w11059_ ;
	wire _w11058_ ;
	wire _w11057_ ;
	wire _w11056_ ;
	wire _w11055_ ;
	wire _w11054_ ;
	wire _w11053_ ;
	wire _w11052_ ;
	wire _w11051_ ;
	wire _w11050_ ;
	wire _w11049_ ;
	wire _w11048_ ;
	wire _w11047_ ;
	wire _w11046_ ;
	wire _w11045_ ;
	wire _w11044_ ;
	wire _w11043_ ;
	wire _w11042_ ;
	wire _w11041_ ;
	wire _w11040_ ;
	wire _w11039_ ;
	wire _w11038_ ;
	wire _w11037_ ;
	wire _w11036_ ;
	wire _w11035_ ;
	wire _w11034_ ;
	wire _w11033_ ;
	wire _w11032_ ;
	wire _w11031_ ;
	wire _w11030_ ;
	wire _w11029_ ;
	wire _w11028_ ;
	wire _w11027_ ;
	wire _w11026_ ;
	wire _w11025_ ;
	wire _w11024_ ;
	wire _w11023_ ;
	wire _w11022_ ;
	wire _w11021_ ;
	wire _w11020_ ;
	wire _w11019_ ;
	wire _w11018_ ;
	wire _w11017_ ;
	wire _w11016_ ;
	wire _w11015_ ;
	wire _w11014_ ;
	wire _w11013_ ;
	wire _w11012_ ;
	wire _w11011_ ;
	wire _w11010_ ;
	wire _w11009_ ;
	wire _w11008_ ;
	wire _w11007_ ;
	wire _w11006_ ;
	wire _w11005_ ;
	wire _w11004_ ;
	wire _w11003_ ;
	wire _w11002_ ;
	wire _w11001_ ;
	wire _w11000_ ;
	wire _w10999_ ;
	wire _w10998_ ;
	wire _w10997_ ;
	wire _w10996_ ;
	wire _w10995_ ;
	wire _w10994_ ;
	wire _w10993_ ;
	wire _w10992_ ;
	wire _w10991_ ;
	wire _w10990_ ;
	wire _w10989_ ;
	wire _w10988_ ;
	wire _w10987_ ;
	wire _w10986_ ;
	wire _w10985_ ;
	wire _w10984_ ;
	wire _w10983_ ;
	wire _w10982_ ;
	wire _w10981_ ;
	wire _w10980_ ;
	wire _w10979_ ;
	wire _w10978_ ;
	wire _w10977_ ;
	wire _w10976_ ;
	wire _w10975_ ;
	wire _w10974_ ;
	wire _w10973_ ;
	wire _w10972_ ;
	wire _w10971_ ;
	wire _w10970_ ;
	wire _w10969_ ;
	wire _w10968_ ;
	wire _w10967_ ;
	wire _w10966_ ;
	wire _w10965_ ;
	wire _w10964_ ;
	wire _w10963_ ;
	wire _w10962_ ;
	wire _w10961_ ;
	wire _w10960_ ;
	wire _w10959_ ;
	wire _w10958_ ;
	wire _w10957_ ;
	wire _w10956_ ;
	wire _w10955_ ;
	wire _w10954_ ;
	wire _w10953_ ;
	wire _w10952_ ;
	wire _w10951_ ;
	wire _w10950_ ;
	wire _w10949_ ;
	wire _w10948_ ;
	wire _w10947_ ;
	wire _w10946_ ;
	wire _w10945_ ;
	wire _w10944_ ;
	wire _w10943_ ;
	wire _w10942_ ;
	wire _w10941_ ;
	wire _w10940_ ;
	wire _w10939_ ;
	wire _w10938_ ;
	wire _w10937_ ;
	wire _w10936_ ;
	wire _w10935_ ;
	wire _w10934_ ;
	wire _w10933_ ;
	wire _w10932_ ;
	wire _w10931_ ;
	wire _w10930_ ;
	wire _w10929_ ;
	wire _w10928_ ;
	wire _w10927_ ;
	wire _w10926_ ;
	wire _w10925_ ;
	wire _w10924_ ;
	wire _w10923_ ;
	wire _w10922_ ;
	wire _w10921_ ;
	wire _w10920_ ;
	wire _w10919_ ;
	wire _w10918_ ;
	wire _w10917_ ;
	wire _w10916_ ;
	wire _w10915_ ;
	wire _w10914_ ;
	wire _w10913_ ;
	wire _w10912_ ;
	wire _w10911_ ;
	wire _w10910_ ;
	wire _w10909_ ;
	wire _w10908_ ;
	wire _w10907_ ;
	wire _w10906_ ;
	wire _w10905_ ;
	wire _w10904_ ;
	wire _w10903_ ;
	wire _w10902_ ;
	wire _w10901_ ;
	wire _w10900_ ;
	wire _w10899_ ;
	wire _w10898_ ;
	wire _w10897_ ;
	wire _w10896_ ;
	wire _w10895_ ;
	wire _w10894_ ;
	wire _w10893_ ;
	wire _w10892_ ;
	wire _w10891_ ;
	wire _w10890_ ;
	wire _w10889_ ;
	wire _w10888_ ;
	wire _w10887_ ;
	wire _w10886_ ;
	wire _w10885_ ;
	wire _w10884_ ;
	wire _w10883_ ;
	wire _w10882_ ;
	wire _w10881_ ;
	wire _w10880_ ;
	wire _w10879_ ;
	wire _w10878_ ;
	wire _w10877_ ;
	wire _w10876_ ;
	wire _w10875_ ;
	wire _w10874_ ;
	wire _w10873_ ;
	wire _w10872_ ;
	wire _w10871_ ;
	wire _w10870_ ;
	wire _w10869_ ;
	wire _w10868_ ;
	wire _w10867_ ;
	wire _w10866_ ;
	wire _w10865_ ;
	wire _w10864_ ;
	wire _w10863_ ;
	wire _w10862_ ;
	wire _w10861_ ;
	wire _w10860_ ;
	wire _w10859_ ;
	wire _w10858_ ;
	wire _w10857_ ;
	wire _w10856_ ;
	wire _w10855_ ;
	wire _w10854_ ;
	wire _w10853_ ;
	wire _w10852_ ;
	wire _w10851_ ;
	wire _w10850_ ;
	wire _w10849_ ;
	wire _w10848_ ;
	wire _w10847_ ;
	wire _w10846_ ;
	wire _w10845_ ;
	wire _w10844_ ;
	wire _w10843_ ;
	wire _w10842_ ;
	wire _w10841_ ;
	wire _w10840_ ;
	wire _w10839_ ;
	wire _w10838_ ;
	wire _w10837_ ;
	wire _w10836_ ;
	wire _w10835_ ;
	wire _w10834_ ;
	wire _w10833_ ;
	wire _w10832_ ;
	wire _w10831_ ;
	wire _w10830_ ;
	wire _w10829_ ;
	wire _w10828_ ;
	wire _w10827_ ;
	wire _w10826_ ;
	wire _w10825_ ;
	wire _w10824_ ;
	wire _w10823_ ;
	wire _w10822_ ;
	wire _w10821_ ;
	wire _w10820_ ;
	wire _w10819_ ;
	wire _w10818_ ;
	wire _w10817_ ;
	wire _w10816_ ;
	wire _w10815_ ;
	wire _w10814_ ;
	wire _w10813_ ;
	wire _w10812_ ;
	wire _w10811_ ;
	wire _w10810_ ;
	wire _w10809_ ;
	wire _w10808_ ;
	wire _w10807_ ;
	wire _w10806_ ;
	wire _w10805_ ;
	wire _w5618_ ;
	wire _w5617_ ;
	wire _w5616_ ;
	wire _w5615_ ;
	wire _w5614_ ;
	wire _w5613_ ;
	wire _w5612_ ;
	wire _w5611_ ;
	wire _w5610_ ;
	wire _w5609_ ;
	wire _w5608_ ;
	wire _w5607_ ;
	wire _w5606_ ;
	wire _w5605_ ;
	wire _w5604_ ;
	wire _w5603_ ;
	wire _w5602_ ;
	wire _w5601_ ;
	wire _w5600_ ;
	wire _w5599_ ;
	wire _w5598_ ;
	wire _w5597_ ;
	wire _w5596_ ;
	wire _w5595_ ;
	wire _w5594_ ;
	wire _w5593_ ;
	wire _w5592_ ;
	wire _w5591_ ;
	wire _w5590_ ;
	wire _w5589_ ;
	wire _w5588_ ;
	wire _w5587_ ;
	wire _w5586_ ;
	wire _w5585_ ;
	wire _w5584_ ;
	wire _w5583_ ;
	wire _w5582_ ;
	wire _w5581_ ;
	wire _w5580_ ;
	wire _w5579_ ;
	wire _w5578_ ;
	wire _w5577_ ;
	wire _w5576_ ;
	wire _w5575_ ;
	wire _w5574_ ;
	wire _w5573_ ;
	wire _w5572_ ;
	wire _w5571_ ;
	wire _w5570_ ;
	wire _w5569_ ;
	wire _w5568_ ;
	wire _w5567_ ;
	wire _w5566_ ;
	wire _w5565_ ;
	wire _w5564_ ;
	wire _w5563_ ;
	wire _w5562_ ;
	wire _w5561_ ;
	wire _w5560_ ;
	wire _w5559_ ;
	wire _w5558_ ;
	wire _w5557_ ;
	wire _w5556_ ;
	wire _w5555_ ;
	wire _w5554_ ;
	wire _w5553_ ;
	wire _w5552_ ;
	wire _w5551_ ;
	wire _w5550_ ;
	wire _w5549_ ;
	wire _w5548_ ;
	wire _w5547_ ;
	wire _w5546_ ;
	wire _w5545_ ;
	wire _w5544_ ;
	wire _w5543_ ;
	wire _w5542_ ;
	wire _w5541_ ;
	wire _w5540_ ;
	wire _w5539_ ;
	wire _w5538_ ;
	wire _w5537_ ;
	wire _w5536_ ;
	wire _w5535_ ;
	wire _w5534_ ;
	wire _w5533_ ;
	wire _w5532_ ;
	wire _w5531_ ;
	wire _w5530_ ;
	wire _w5529_ ;
	wire _w5528_ ;
	wire _w5527_ ;
	wire _w5526_ ;
	wire _w5525_ ;
	wire _w5524_ ;
	wire _w5523_ ;
	wire _w5522_ ;
	wire _w5521_ ;
	wire _w5520_ ;
	wire _w5519_ ;
	wire _w5518_ ;
	wire _w5517_ ;
	wire _w5516_ ;
	wire _w5515_ ;
	wire _w5514_ ;
	wire _w5513_ ;
	wire _w5512_ ;
	wire _w5511_ ;
	wire _w5510_ ;
	wire _w5509_ ;
	wire _w5508_ ;
	wire _w5507_ ;
	wire _w5506_ ;
	wire _w5505_ ;
	wire _w5504_ ;
	wire _w5503_ ;
	wire _w5502_ ;
	wire _w5501_ ;
	wire _w5500_ ;
	wire _w5499_ ;
	wire _w5498_ ;
	wire _w5497_ ;
	wire _w5496_ ;
	wire _w5495_ ;
	wire _w5494_ ;
	wire _w5493_ ;
	wire _w5492_ ;
	wire _w5491_ ;
	wire _w5490_ ;
	wire _w5489_ ;
	wire _w5488_ ;
	wire _w5487_ ;
	wire _w5486_ ;
	wire _w5485_ ;
	wire _w5484_ ;
	wire _w5483_ ;
	wire _w5482_ ;
	wire _w5481_ ;
	wire _w5480_ ;
	wire _w5479_ ;
	wire _w5478_ ;
	wire _w5477_ ;
	wire _w5476_ ;
	wire _w5475_ ;
	wire _w5474_ ;
	wire _w5473_ ;
	wire _w5472_ ;
	wire _w5471_ ;
	wire _w5470_ ;
	wire _w5469_ ;
	wire _w5468_ ;
	wire _w5467_ ;
	wire _w5466_ ;
	wire _w5465_ ;
	wire _w5464_ ;
	wire _w5463_ ;
	wire _w5462_ ;
	wire _w5461_ ;
	wire _w5460_ ;
	wire _w5459_ ;
	wire _w5458_ ;
	wire _w5457_ ;
	wire _w5456_ ;
	wire _w5455_ ;
	wire _w5454_ ;
	wire _w5453_ ;
	wire _w5452_ ;
	wire _w5451_ ;
	wire _w5450_ ;
	wire _w5449_ ;
	wire _w5448_ ;
	wire _w5447_ ;
	wire _w5446_ ;
	wire _w5445_ ;
	wire _w5444_ ;
	wire _w5443_ ;
	wire _w5442_ ;
	wire _w5441_ ;
	wire _w5440_ ;
	wire _w5439_ ;
	wire _w5438_ ;
	wire _w5437_ ;
	wire _w5436_ ;
	wire _w5435_ ;
	wire _w5434_ ;
	wire _w5433_ ;
	wire _w5432_ ;
	wire _w5431_ ;
	wire _w5430_ ;
	wire _w5429_ ;
	wire _w5428_ ;
	wire _w5427_ ;
	wire _w5426_ ;
	wire _w5425_ ;
	wire _w5424_ ;
	wire _w5423_ ;
	wire _w5422_ ;
	wire _w5421_ ;
	wire _w5420_ ;
	wire _w5419_ ;
	wire _w5418_ ;
	wire _w5417_ ;
	wire _w5416_ ;
	wire _w5415_ ;
	wire _w5414_ ;
	wire _w5413_ ;
	wire _w5412_ ;
	wire _w5411_ ;
	wire _w5410_ ;
	wire _w5409_ ;
	wire _w5408_ ;
	wire _w5407_ ;
	wire _w5406_ ;
	wire _w5405_ ;
	wire _w5404_ ;
	wire _w5403_ ;
	wire _w5402_ ;
	wire _w5401_ ;
	wire _w5400_ ;
	wire _w5399_ ;
	wire _w5398_ ;
	wire _w5397_ ;
	wire _w5396_ ;
	wire _w5395_ ;
	wire _w5394_ ;
	wire _w5393_ ;
	wire _w5392_ ;
	wire _w5391_ ;
	wire _w5390_ ;
	wire _w5389_ ;
	wire _w5388_ ;
	wire _w5387_ ;
	wire _w5386_ ;
	wire _w5385_ ;
	wire _w5384_ ;
	wire _w5383_ ;
	wire _w5382_ ;
	wire _w5381_ ;
	wire _w5380_ ;
	wire _w5379_ ;
	wire _w5378_ ;
	wire _w5377_ ;
	wire _w5376_ ;
	wire _w5375_ ;
	wire _w5374_ ;
	wire _w5373_ ;
	wire _w5372_ ;
	wire _w5371_ ;
	wire _w5370_ ;
	wire _w5369_ ;
	wire _w5368_ ;
	wire _w5367_ ;
	wire _w5366_ ;
	wire _w5365_ ;
	wire _w5364_ ;
	wire _w5363_ ;
	wire _w5362_ ;
	wire _w5361_ ;
	wire _w5360_ ;
	wire _w5359_ ;
	wire _w5358_ ;
	wire _w5357_ ;
	wire _w5356_ ;
	wire _w5355_ ;
	wire _w5354_ ;
	wire _w5353_ ;
	wire _w5352_ ;
	wire _w5351_ ;
	wire _w5350_ ;
	wire _w5349_ ;
	wire _w5348_ ;
	wire _w5347_ ;
	wire _w5346_ ;
	wire _w5345_ ;
	wire _w5344_ ;
	wire _w5343_ ;
	wire _w5342_ ;
	wire _w5341_ ;
	wire _w5340_ ;
	wire _w5339_ ;
	wire _w5338_ ;
	wire _w5337_ ;
	wire _w5336_ ;
	wire _w5335_ ;
	wire _w5334_ ;
	wire _w5333_ ;
	wire _w5332_ ;
	wire _w5331_ ;
	wire _w5330_ ;
	wire _w5329_ ;
	wire _w5328_ ;
	wire _w5327_ ;
	wire _w5326_ ;
	wire _w5325_ ;
	wire _w5324_ ;
	wire _w5323_ ;
	wire _w5322_ ;
	wire _w5321_ ;
	wire _w5320_ ;
	wire _w5319_ ;
	wire _w5318_ ;
	wire _w5317_ ;
	wire _w5316_ ;
	wire _w5315_ ;
	wire _w5314_ ;
	wire _w5313_ ;
	wire _w5312_ ;
	wire _w5311_ ;
	wire _w5310_ ;
	wire _w5309_ ;
	wire _w5308_ ;
	wire _w5307_ ;
	wire _w5306_ ;
	wire _w5305_ ;
	wire _w5304_ ;
	wire _w5303_ ;
	wire _w5302_ ;
	wire _w5301_ ;
	wire _w5300_ ;
	wire _w5299_ ;
	wire _w5298_ ;
	wire _w5297_ ;
	wire _w5296_ ;
	wire _w5295_ ;
	wire _w5294_ ;
	wire _w5293_ ;
	wire _w5292_ ;
	wire _w5291_ ;
	wire _w5290_ ;
	wire _w5289_ ;
	wire _w5288_ ;
	wire _w5287_ ;
	wire _w5286_ ;
	wire _w5285_ ;
	wire _w5284_ ;
	wire _w5283_ ;
	wire _w5282_ ;
	wire _w5281_ ;
	wire _w5280_ ;
	wire _w5279_ ;
	wire _w5278_ ;
	wire _w5277_ ;
	wire _w5276_ ;
	wire _w5275_ ;
	wire _w5274_ ;
	wire _w5273_ ;
	wire _w5272_ ;
	wire _w5271_ ;
	wire _w5270_ ;
	wire _w5269_ ;
	wire _w5268_ ;
	wire _w5267_ ;
	wire _w5266_ ;
	wire _w5265_ ;
	wire _w5264_ ;
	wire _w5263_ ;
	wire _w5262_ ;
	wire _w5261_ ;
	wire _w5260_ ;
	wire _w5259_ ;
	wire _w5258_ ;
	wire _w5257_ ;
	wire _w5256_ ;
	wire _w5255_ ;
	wire _w5254_ ;
	wire _w5253_ ;
	wire _w5252_ ;
	wire _w5251_ ;
	wire _w5250_ ;
	wire _w5249_ ;
	wire _w5248_ ;
	wire _w5247_ ;
	wire _w5246_ ;
	wire _w5245_ ;
	wire _w5244_ ;
	wire _w5243_ ;
	wire _w5242_ ;
	wire _w5241_ ;
	wire _w5240_ ;
	wire _w5239_ ;
	wire _w5238_ ;
	wire _w5237_ ;
	wire _w5236_ ;
	wire _w5235_ ;
	wire _w5234_ ;
	wire _w5233_ ;
	wire _w5232_ ;
	wire _w5231_ ;
	wire _w5230_ ;
	wire _w5229_ ;
	wire _w5228_ ;
	wire _w5227_ ;
	wire _w5226_ ;
	wire _w5225_ ;
	wire _w5224_ ;
	wire _w5223_ ;
	wire _w5222_ ;
	wire _w5221_ ;
	wire _w5220_ ;
	wire _w5219_ ;
	wire _w5218_ ;
	wire _w5217_ ;
	wire _w5216_ ;
	wire _w5215_ ;
	wire _w5214_ ;
	wire _w5213_ ;
	wire _w5212_ ;
	wire _w5211_ ;
	wire _w5210_ ;
	wire _w5209_ ;
	wire _w5208_ ;
	wire _w5207_ ;
	wire _w5206_ ;
	wire _w5205_ ;
	wire _w5204_ ;
	wire _w5203_ ;
	wire _w5202_ ;
	wire _w5201_ ;
	wire _w5200_ ;
	wire _w5199_ ;
	wire _w5198_ ;
	wire _w5197_ ;
	wire _w5196_ ;
	wire _w5195_ ;
	wire _w5194_ ;
	wire _w5193_ ;
	wire _w5192_ ;
	wire _w5191_ ;
	wire _w5190_ ;
	wire _w5189_ ;
	wire _w5188_ ;
	wire _w5187_ ;
	wire _w5186_ ;
	wire _w5185_ ;
	wire _w5184_ ;
	wire _w5183_ ;
	wire _w5182_ ;
	wire _w5181_ ;
	wire _w5180_ ;
	wire _w5179_ ;
	wire _w5178_ ;
	wire _w5177_ ;
	wire _w5176_ ;
	wire _w5175_ ;
	wire _w5174_ ;
	wire _w5173_ ;
	wire _w5172_ ;
	wire _w5171_ ;
	wire _w5170_ ;
	wire _w5169_ ;
	wire _w5168_ ;
	wire _w5167_ ;
	wire _w5166_ ;
	wire _w5165_ ;
	wire _w5164_ ;
	wire _w5163_ ;
	wire _w5162_ ;
	wire _w5161_ ;
	wire _w5160_ ;
	wire _w5159_ ;
	wire _w5158_ ;
	wire _w5157_ ;
	wire _w5156_ ;
	wire _w5155_ ;
	wire _w5154_ ;
	wire _w5153_ ;
	wire _w5152_ ;
	wire _w5151_ ;
	wire _w5150_ ;
	wire _w5149_ ;
	wire _w5148_ ;
	wire _w5147_ ;
	wire _w5146_ ;
	wire _w5145_ ;
	wire _w5144_ ;
	wire _w5143_ ;
	wire _w5142_ ;
	wire _w5141_ ;
	wire _w5140_ ;
	wire _w5139_ ;
	wire _w5138_ ;
	wire _w5137_ ;
	wire _w5136_ ;
	wire _w5135_ ;
	wire _w5134_ ;
	wire _w5133_ ;
	wire _w5132_ ;
	wire _w5131_ ;
	wire _w5130_ ;
	wire _w5129_ ;
	wire _w5128_ ;
	wire _w5127_ ;
	wire _w5126_ ;
	wire _w5125_ ;
	wire _w5124_ ;
	wire _w5123_ ;
	wire _w5122_ ;
	wire _w5121_ ;
	wire _w5120_ ;
	wire _w5119_ ;
	wire _w5118_ ;
	wire _w5117_ ;
	wire _w5116_ ;
	wire _w5115_ ;
	wire _w5114_ ;
	wire _w5113_ ;
	wire _w5112_ ;
	wire _w5111_ ;
	wire _w5110_ ;
	wire _w5109_ ;
	wire _w5108_ ;
	wire _w5107_ ;
	wire _w5106_ ;
	wire _w5105_ ;
	wire _w5104_ ;
	wire _w5103_ ;
	wire _w5102_ ;
	wire _w5101_ ;
	wire _w5100_ ;
	wire _w5099_ ;
	wire _w5098_ ;
	wire _w5097_ ;
	wire _w5096_ ;
	wire _w5095_ ;
	wire _w5094_ ;
	wire _w5093_ ;
	wire _w5092_ ;
	wire _w5091_ ;
	wire _w5090_ ;
	wire _w5089_ ;
	wire _w5088_ ;
	wire _w5087_ ;
	wire _w5086_ ;
	wire _w5085_ ;
	wire _w5084_ ;
	wire _w5083_ ;
	wire _w5082_ ;
	wire _w5081_ ;
	wire _w5080_ ;
	wire _w5079_ ;
	wire _w5078_ ;
	wire _w5077_ ;
	wire _w5076_ ;
	wire _w5075_ ;
	wire _w5074_ ;
	wire _w5073_ ;
	wire _w5072_ ;
	wire _w5071_ ;
	wire _w5070_ ;
	wire _w5069_ ;
	wire _w5068_ ;
	wire _w5067_ ;
	wire _w5066_ ;
	wire _w5065_ ;
	wire _w5064_ ;
	wire _w5063_ ;
	wire _w5062_ ;
	wire _w5061_ ;
	wire _w5060_ ;
	wire _w5059_ ;
	wire _w5058_ ;
	wire _w5057_ ;
	wire _w5056_ ;
	wire _w5055_ ;
	wire _w5054_ ;
	wire _w5053_ ;
	wire _w5052_ ;
	wire _w5051_ ;
	wire _w5050_ ;
	wire _w5049_ ;
	wire _w5048_ ;
	wire _w5047_ ;
	wire _w5046_ ;
	wire _w5045_ ;
	wire _w5044_ ;
	wire _w5043_ ;
	wire _w5042_ ;
	wire _w5041_ ;
	wire _w5040_ ;
	wire _w5039_ ;
	wire _w5038_ ;
	wire _w5037_ ;
	wire _w5036_ ;
	wire _w5035_ ;
	wire _w5034_ ;
	wire _w5033_ ;
	wire _w5032_ ;
	wire _w5031_ ;
	wire _w5030_ ;
	wire _w5029_ ;
	wire _w5028_ ;
	wire _w5027_ ;
	wire _w5026_ ;
	wire _w5025_ ;
	wire _w5024_ ;
	wire _w5023_ ;
	wire _w5022_ ;
	wire _w5021_ ;
	wire _w5020_ ;
	wire _w5019_ ;
	wire _w5018_ ;
	wire _w5017_ ;
	wire _w5016_ ;
	wire _w5015_ ;
	wire _w5014_ ;
	wire _w5013_ ;
	wire _w5012_ ;
	wire _w5011_ ;
	wire _w5010_ ;
	wire _w5009_ ;
	wire _w5008_ ;
	wire _w5007_ ;
	wire _w5006_ ;
	wire _w5005_ ;
	wire _w5004_ ;
	wire _w5003_ ;
	wire _w5002_ ;
	wire _w5001_ ;
	wire _w5000_ ;
	wire _w4999_ ;
	wire _w4998_ ;
	wire _w4997_ ;
	wire _w4996_ ;
	wire _w4995_ ;
	wire _w4994_ ;
	wire _w4993_ ;
	wire _w4992_ ;
	wire _w4991_ ;
	wire _w4990_ ;
	wire _w4989_ ;
	wire _w4988_ ;
	wire _w4987_ ;
	wire _w4986_ ;
	wire _w4985_ ;
	wire _w4984_ ;
	wire _w4983_ ;
	wire _w4982_ ;
	wire _w4981_ ;
	wire _w4980_ ;
	wire _w4979_ ;
	wire _w4978_ ;
	wire _w4977_ ;
	wire _w4976_ ;
	wire _w4975_ ;
	wire _w4974_ ;
	wire _w4973_ ;
	wire _w4972_ ;
	wire _w4971_ ;
	wire _w4970_ ;
	wire _w4969_ ;
	wire _w4968_ ;
	wire _w4967_ ;
	wire _w4966_ ;
	wire _w4965_ ;
	wire _w4964_ ;
	wire _w4963_ ;
	wire _w4962_ ;
	wire _w4961_ ;
	wire _w4960_ ;
	wire _w4959_ ;
	wire _w4958_ ;
	wire _w4957_ ;
	wire _w4956_ ;
	wire _w4955_ ;
	wire _w4954_ ;
	wire _w4953_ ;
	wire _w4952_ ;
	wire _w4951_ ;
	wire _w4950_ ;
	wire _w4949_ ;
	wire _w4948_ ;
	wire _w4947_ ;
	wire _w4946_ ;
	wire _w4945_ ;
	wire _w4944_ ;
	wire _w4943_ ;
	wire _w4942_ ;
	wire _w4941_ ;
	wire _w4940_ ;
	wire _w4939_ ;
	wire _w4938_ ;
	wire _w4937_ ;
	wire _w4936_ ;
	wire _w4935_ ;
	wire _w4934_ ;
	wire _w4933_ ;
	wire _w4932_ ;
	wire _w4931_ ;
	wire _w4930_ ;
	wire _w4929_ ;
	wire _w4928_ ;
	wire _w4927_ ;
	wire _w4926_ ;
	wire _w4925_ ;
	wire _w4924_ ;
	wire _w4923_ ;
	wire _w4922_ ;
	wire _w4921_ ;
	wire _w4920_ ;
	wire _w4919_ ;
	wire _w4918_ ;
	wire _w4917_ ;
	wire _w4916_ ;
	wire _w4915_ ;
	wire _w4914_ ;
	wire _w4913_ ;
	wire _w4912_ ;
	wire _w4911_ ;
	wire _w4910_ ;
	wire _w4909_ ;
	wire _w4908_ ;
	wire _w4907_ ;
	wire _w4906_ ;
	wire _w4905_ ;
	wire _w4904_ ;
	wire _w4903_ ;
	wire _w4902_ ;
	wire _w4901_ ;
	wire _w4900_ ;
	wire _w4899_ ;
	wire _w4898_ ;
	wire _w4897_ ;
	wire _w4896_ ;
	wire _w4895_ ;
	wire _w4894_ ;
	wire _w4893_ ;
	wire _w4892_ ;
	wire _w4891_ ;
	wire _w4890_ ;
	wire _w4889_ ;
	wire _w4888_ ;
	wire _w4887_ ;
	wire _w4886_ ;
	wire _w4885_ ;
	wire _w4884_ ;
	wire _w4883_ ;
	wire _w4882_ ;
	wire _w4881_ ;
	wire _w4880_ ;
	wire _w4879_ ;
	wire _w4878_ ;
	wire _w4877_ ;
	wire _w4876_ ;
	wire _w4875_ ;
	wire _w4874_ ;
	wire _w4873_ ;
	wire _w4872_ ;
	wire _w4871_ ;
	wire _w4870_ ;
	wire _w4869_ ;
	wire _w4868_ ;
	wire _w4867_ ;
	wire _w4866_ ;
	wire _w4865_ ;
	wire _w4864_ ;
	wire _w4863_ ;
	wire _w4862_ ;
	wire _w4861_ ;
	wire _w4860_ ;
	wire _w4859_ ;
	wire _w4858_ ;
	wire _w4857_ ;
	wire _w4856_ ;
	wire _w4855_ ;
	wire _w4854_ ;
	wire _w4853_ ;
	wire _w4852_ ;
	wire _w4851_ ;
	wire _w4850_ ;
	wire _w4849_ ;
	wire _w4848_ ;
	wire _w4847_ ;
	wire _w4846_ ;
	wire _w4845_ ;
	wire _w4844_ ;
	wire _w4843_ ;
	wire _w4842_ ;
	wire _w4841_ ;
	wire _w4840_ ;
	wire _w4839_ ;
	wire _w4838_ ;
	wire _w4837_ ;
	wire _w4836_ ;
	wire _w4835_ ;
	wire _w4834_ ;
	wire _w4833_ ;
	wire _w4832_ ;
	wire _w4831_ ;
	wire _w4830_ ;
	wire _w4829_ ;
	wire _w4828_ ;
	wire _w4827_ ;
	wire _w4826_ ;
	wire _w4825_ ;
	wire _w4824_ ;
	wire _w4823_ ;
	wire _w4822_ ;
	wire _w4821_ ;
	wire _w4820_ ;
	wire _w4819_ ;
	wire _w4818_ ;
	wire _w4817_ ;
	wire _w4816_ ;
	wire _w4815_ ;
	wire _w4814_ ;
	wire _w4813_ ;
	wire _w4812_ ;
	wire _w4811_ ;
	wire _w4810_ ;
	wire _w4809_ ;
	wire _w4808_ ;
	wire _w4807_ ;
	wire _w4806_ ;
	wire _w4805_ ;
	wire _w4804_ ;
	wire _w4803_ ;
	wire _w4802_ ;
	wire _w4801_ ;
	wire _w4800_ ;
	wire _w4799_ ;
	wire _w4798_ ;
	wire _w4797_ ;
	wire _w4796_ ;
	wire _w4795_ ;
	wire _w4794_ ;
	wire _w4793_ ;
	wire _w4792_ ;
	wire _w4791_ ;
	wire _w4790_ ;
	wire _w4789_ ;
	wire _w4788_ ;
	wire _w4787_ ;
	wire _w4786_ ;
	wire _w4785_ ;
	wire _w4784_ ;
	wire _w4783_ ;
	wire _w4782_ ;
	wire _w4781_ ;
	wire _w4780_ ;
	wire _w4779_ ;
	wire _w4778_ ;
	wire _w4777_ ;
	wire _w4776_ ;
	wire _w4775_ ;
	wire _w4774_ ;
	wire _w4773_ ;
	wire _w4772_ ;
	wire _w4771_ ;
	wire _w4770_ ;
	wire _w4769_ ;
	wire _w4768_ ;
	wire _w4767_ ;
	wire _w4766_ ;
	wire _w4765_ ;
	wire _w4764_ ;
	wire _w4763_ ;
	wire _w4762_ ;
	wire _w4761_ ;
	wire _w4760_ ;
	wire _w4759_ ;
	wire _w4758_ ;
	wire _w4757_ ;
	wire _w4756_ ;
	wire _w4755_ ;
	wire _w4754_ ;
	wire _w4753_ ;
	wire _w4752_ ;
	wire _w4751_ ;
	wire _w4750_ ;
	wire _w4749_ ;
	wire _w4748_ ;
	wire _w4747_ ;
	wire _w4746_ ;
	wire _w4745_ ;
	wire _w4744_ ;
	wire _w4743_ ;
	wire _w4742_ ;
	wire _w4741_ ;
	wire _w4740_ ;
	wire _w4739_ ;
	wire _w4738_ ;
	wire _w4737_ ;
	wire _w4736_ ;
	wire _w4735_ ;
	wire _w4734_ ;
	wire _w4733_ ;
	wire _w4732_ ;
	wire _w4731_ ;
	wire _w4730_ ;
	wire _w4729_ ;
	wire _w4728_ ;
	wire _w4727_ ;
	wire _w4726_ ;
	wire _w4725_ ;
	wire _w4724_ ;
	wire _w4723_ ;
	wire _w4722_ ;
	wire _w4721_ ;
	wire _w4720_ ;
	wire _w4719_ ;
	wire _w4718_ ;
	wire _w4717_ ;
	wire _w4716_ ;
	wire _w4715_ ;
	wire _w4714_ ;
	wire _w4713_ ;
	wire _w4712_ ;
	wire _w4711_ ;
	wire _w4710_ ;
	wire _w4709_ ;
	wire _w4708_ ;
	wire _w4707_ ;
	wire _w4706_ ;
	wire _w4705_ ;
	wire _w4704_ ;
	wire _w4703_ ;
	wire _w4702_ ;
	wire _w4701_ ;
	wire _w4700_ ;
	wire _w4699_ ;
	wire _w4698_ ;
	wire _w4697_ ;
	wire _w4696_ ;
	wire _w4695_ ;
	wire _w4694_ ;
	wire _w4693_ ;
	wire _w4692_ ;
	wire _w4691_ ;
	wire _w4690_ ;
	wire _w4689_ ;
	wire _w4688_ ;
	wire _w4687_ ;
	wire _w4686_ ;
	wire _w4685_ ;
	wire _w4684_ ;
	wire _w4683_ ;
	wire _w4682_ ;
	wire _w4681_ ;
	wire _w4680_ ;
	wire _w4679_ ;
	wire _w4678_ ;
	wire _w4677_ ;
	wire _w4676_ ;
	wire _w4675_ ;
	wire _w4674_ ;
	wire _w4673_ ;
	wire _w4672_ ;
	wire _w4671_ ;
	wire _w4670_ ;
	wire _w4669_ ;
	wire _w4668_ ;
	wire _w4667_ ;
	wire _w4666_ ;
	wire _w4665_ ;
	wire _w4664_ ;
	wire _w4663_ ;
	wire _w4662_ ;
	wire _w4661_ ;
	wire _w4660_ ;
	wire _w4659_ ;
	wire _w4658_ ;
	wire _w4657_ ;
	wire _w4656_ ;
	wire _w4655_ ;
	wire _w4654_ ;
	wire _w4653_ ;
	wire _w4652_ ;
	wire _w4651_ ;
	wire _w4650_ ;
	wire _w4649_ ;
	wire _w4648_ ;
	wire _w4647_ ;
	wire _w4646_ ;
	wire _w4645_ ;
	wire _w4644_ ;
	wire _w4643_ ;
	wire _w4642_ ;
	wire _w4641_ ;
	wire _w4640_ ;
	wire _w4639_ ;
	wire _w4638_ ;
	wire _w4637_ ;
	wire _w4636_ ;
	wire _w4635_ ;
	wire _w4634_ ;
	wire _w4633_ ;
	wire _w4632_ ;
	wire _w4631_ ;
	wire _w4630_ ;
	wire _w4629_ ;
	wire _w4628_ ;
	wire _w4627_ ;
	wire _w4626_ ;
	wire _w4625_ ;
	wire _w4624_ ;
	wire _w4623_ ;
	wire _w4622_ ;
	wire _w4621_ ;
	wire _w4620_ ;
	wire _w4619_ ;
	wire _w4618_ ;
	wire _w4617_ ;
	wire _w4616_ ;
	wire _w4615_ ;
	wire _w4614_ ;
	wire _w4613_ ;
	wire _w4612_ ;
	wire _w4611_ ;
	wire _w4610_ ;
	wire _w4609_ ;
	wire _w4608_ ;
	wire _w4607_ ;
	wire _w4606_ ;
	wire _w4605_ ;
	wire _w4604_ ;
	wire _w4603_ ;
	wire _w4602_ ;
	wire _w4601_ ;
	wire _w4600_ ;
	wire _w4599_ ;
	wire _w4598_ ;
	wire _w4597_ ;
	wire _w4596_ ;
	wire _w4595_ ;
	wire _w4594_ ;
	wire _w4593_ ;
	wire _w4592_ ;
	wire _w4591_ ;
	wire _w4590_ ;
	wire _w4589_ ;
	wire _w4588_ ;
	wire _w4587_ ;
	wire _w4586_ ;
	wire _w4585_ ;
	wire _w4584_ ;
	wire _w4583_ ;
	wire _w4582_ ;
	wire _w4581_ ;
	wire _w4580_ ;
	wire _w4579_ ;
	wire _w4578_ ;
	wire _w4577_ ;
	wire _w4576_ ;
	wire _w4575_ ;
	wire _w4574_ ;
	wire _w4573_ ;
	wire _w4572_ ;
	wire _w4571_ ;
	wire _w4570_ ;
	wire _w4569_ ;
	wire _w4568_ ;
	wire _w4567_ ;
	wire _w4566_ ;
	wire _w4565_ ;
	wire _w4564_ ;
	wire _w4563_ ;
	wire _w4562_ ;
	wire _w4561_ ;
	wire _w4560_ ;
	wire _w4559_ ;
	wire _w4558_ ;
	wire _w4557_ ;
	wire _w4556_ ;
	wire _w4555_ ;
	wire _w4554_ ;
	wire _w4553_ ;
	wire _w4552_ ;
	wire _w4551_ ;
	wire _w4550_ ;
	wire _w4549_ ;
	wire _w4548_ ;
	wire _w4547_ ;
	wire _w4546_ ;
	wire _w4545_ ;
	wire _w4544_ ;
	wire _w4543_ ;
	wire _w4542_ ;
	wire _w4541_ ;
	wire _w4540_ ;
	wire _w4539_ ;
	wire _w4538_ ;
	wire _w4537_ ;
	wire _w4536_ ;
	wire _w4535_ ;
	wire _w4534_ ;
	wire _w4533_ ;
	wire _w4532_ ;
	wire _w4531_ ;
	wire _w4530_ ;
	wire _w4529_ ;
	wire _w4528_ ;
	wire _w4527_ ;
	wire _w4526_ ;
	wire _w4525_ ;
	wire _w4524_ ;
	wire _w4523_ ;
	wire _w4522_ ;
	wire _w4521_ ;
	wire _w4520_ ;
	wire _w4519_ ;
	wire _w4518_ ;
	wire _w4517_ ;
	wire _w4516_ ;
	wire _w4515_ ;
	wire _w4514_ ;
	wire _w4513_ ;
	wire _w4512_ ;
	wire _w4511_ ;
	wire _w4510_ ;
	wire _w4509_ ;
	wire _w4508_ ;
	wire _w4507_ ;
	wire _w4506_ ;
	wire _w4505_ ;
	wire _w4504_ ;
	wire _w4503_ ;
	wire _w4502_ ;
	wire _w4501_ ;
	wire _w4500_ ;
	wire _w4499_ ;
	wire _w4498_ ;
	wire _w4497_ ;
	wire _w4496_ ;
	wire _w4495_ ;
	wire _w4494_ ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w5619_ ;
	wire _w5620_ ;
	wire _w5621_ ;
	wire _w5622_ ;
	wire _w5623_ ;
	wire _w5624_ ;
	wire _w5625_ ;
	wire _w5626_ ;
	wire _w5627_ ;
	wire _w5628_ ;
	wire _w5629_ ;
	wire _w5630_ ;
	wire _w5631_ ;
	wire _w5632_ ;
	wire _w5633_ ;
	wire _w5634_ ;
	wire _w5635_ ;
	wire _w5636_ ;
	wire _w5637_ ;
	wire _w5638_ ;
	wire _w5639_ ;
	wire _w5640_ ;
	wire _w5641_ ;
	wire _w5642_ ;
	wire _w5643_ ;
	wire _w5644_ ;
	wire _w5645_ ;
	wire _w5646_ ;
	wire _w5647_ ;
	wire _w5648_ ;
	wire _w5649_ ;
	wire _w5650_ ;
	wire _w5651_ ;
	wire _w5652_ ;
	wire _w5653_ ;
	wire _w5654_ ;
	wire _w5655_ ;
	wire _w5656_ ;
	wire _w5657_ ;
	wire _w5658_ ;
	wire _w5659_ ;
	wire _w5660_ ;
	wire _w5661_ ;
	wire _w5662_ ;
	wire _w5663_ ;
	wire _w5664_ ;
	wire _w5665_ ;
	wire _w5666_ ;
	wire _w5667_ ;
	wire _w5668_ ;
	wire _w5669_ ;
	wire _w5670_ ;
	wire _w5671_ ;
	wire _w5672_ ;
	wire _w5673_ ;
	wire _w5674_ ;
	wire _w5675_ ;
	wire _w5676_ ;
	wire _w5677_ ;
	wire _w5678_ ;
	wire _w5679_ ;
	wire _w5680_ ;
	wire _w5681_ ;
	wire _w5682_ ;
	wire _w5683_ ;
	wire _w5684_ ;
	wire _w5685_ ;
	wire _w5686_ ;
	wire _w5687_ ;
	wire _w5688_ ;
	wire _w5689_ ;
	wire _w5690_ ;
	wire _w5691_ ;
	wire _w5692_ ;
	wire _w5693_ ;
	wire _w5694_ ;
	wire _w5695_ ;
	wire _w5696_ ;
	wire _w5697_ ;
	wire _w5698_ ;
	wire _w5699_ ;
	wire _w5700_ ;
	wire _w5701_ ;
	wire _w5702_ ;
	wire _w5703_ ;
	wire _w5704_ ;
	wire _w5705_ ;
	wire _w5706_ ;
	wire _w5707_ ;
	wire _w5708_ ;
	wire _w5709_ ;
	wire _w5710_ ;
	wire _w5711_ ;
	wire _w5712_ ;
	wire _w5713_ ;
	wire _w5714_ ;
	wire _w5715_ ;
	wire _w5716_ ;
	wire _w5717_ ;
	wire _w5718_ ;
	wire _w5719_ ;
	wire _w5720_ ;
	wire _w5721_ ;
	wire _w5722_ ;
	wire _w5723_ ;
	wire _w5724_ ;
	wire _w5725_ ;
	wire _w5726_ ;
	wire _w5727_ ;
	wire _w5728_ ;
	wire _w5729_ ;
	wire _w5730_ ;
	wire _w5731_ ;
	wire _w5732_ ;
	wire _w5733_ ;
	wire _w5734_ ;
	wire _w5735_ ;
	wire _w5736_ ;
	wire _w5737_ ;
	wire _w5738_ ;
	wire _w5739_ ;
	wire _w5740_ ;
	wire _w5741_ ;
	wire _w5742_ ;
	wire _w5743_ ;
	wire _w5744_ ;
	wire _w5745_ ;
	wire _w5746_ ;
	wire _w5747_ ;
	wire _w5748_ ;
	wire _w5749_ ;
	wire _w5750_ ;
	wire _w5751_ ;
	wire _w5752_ ;
	wire _w5753_ ;
	wire _w5754_ ;
	wire _w5755_ ;
	wire _w5756_ ;
	wire _w5757_ ;
	wire _w5758_ ;
	wire _w5759_ ;
	wire _w5760_ ;
	wire _w5761_ ;
	wire _w5762_ ;
	wire _w5763_ ;
	wire _w5764_ ;
	wire _w5765_ ;
	wire _w5766_ ;
	wire _w5767_ ;
	wire _w5768_ ;
	wire _w5769_ ;
	wire _w5770_ ;
	wire _w5771_ ;
	wire _w5772_ ;
	wire _w5773_ ;
	wire _w5774_ ;
	wire _w5775_ ;
	wire _w5776_ ;
	wire _w5777_ ;
	wire _w5778_ ;
	wire _w5779_ ;
	wire _w5780_ ;
	wire _w5781_ ;
	wire _w5782_ ;
	wire _w5783_ ;
	wire _w5784_ ;
	wire _w5785_ ;
	wire _w5786_ ;
	wire _w5787_ ;
	wire _w5788_ ;
	wire _w5789_ ;
	wire _w5790_ ;
	wire _w5791_ ;
	wire _w5792_ ;
	wire _w5793_ ;
	wire _w5794_ ;
	wire _w5795_ ;
	wire _w5796_ ;
	wire _w5797_ ;
	wire _w5798_ ;
	wire _w5799_ ;
	wire _w5800_ ;
	wire _w5801_ ;
	wire _w5802_ ;
	wire _w5803_ ;
	wire _w5804_ ;
	wire _w5805_ ;
	wire _w5806_ ;
	wire _w5807_ ;
	wire _w5808_ ;
	wire _w5809_ ;
	wire _w5810_ ;
	wire _w5811_ ;
	wire _w5812_ ;
	wire _w5813_ ;
	wire _w5814_ ;
	wire _w5815_ ;
	wire _w5816_ ;
	wire _w5817_ ;
	wire _w5818_ ;
	wire _w5819_ ;
	wire _w5820_ ;
	wire _w5821_ ;
	wire _w5822_ ;
	wire _w5823_ ;
	wire _w5824_ ;
	wire _w5825_ ;
	wire _w5826_ ;
	wire _w5827_ ;
	wire _w5828_ ;
	wire _w5829_ ;
	wire _w5830_ ;
	wire _w5831_ ;
	wire _w5832_ ;
	wire _w5833_ ;
	wire _w5834_ ;
	wire _w5835_ ;
	wire _w5836_ ;
	wire _w5837_ ;
	wire _w5838_ ;
	wire _w5839_ ;
	wire _w5840_ ;
	wire _w5841_ ;
	wire _w5842_ ;
	wire _w5843_ ;
	wire _w5844_ ;
	wire _w5845_ ;
	wire _w5846_ ;
	wire _w5847_ ;
	wire _w5848_ ;
	wire _w5849_ ;
	wire _w5850_ ;
	wire _w5851_ ;
	wire _w5852_ ;
	wire _w5853_ ;
	wire _w5854_ ;
	wire _w5855_ ;
	wire _w5856_ ;
	wire _w5857_ ;
	wire _w5858_ ;
	wire _w5859_ ;
	wire _w5860_ ;
	wire _w5861_ ;
	wire _w5862_ ;
	wire _w5863_ ;
	wire _w5864_ ;
	wire _w5865_ ;
	wire _w5866_ ;
	wire _w5867_ ;
	wire _w5868_ ;
	wire _w5869_ ;
	wire _w5870_ ;
	wire _w5871_ ;
	wire _w5872_ ;
	wire _w5873_ ;
	wire _w5874_ ;
	wire _w5875_ ;
	wire _w5876_ ;
	wire _w5877_ ;
	wire _w5878_ ;
	wire _w5879_ ;
	wire _w5880_ ;
	wire _w5881_ ;
	wire _w5882_ ;
	wire _w5883_ ;
	wire _w5884_ ;
	wire _w5885_ ;
	wire _w5886_ ;
	wire _w5887_ ;
	wire _w5888_ ;
	wire _w5889_ ;
	wire _w5890_ ;
	wire _w5891_ ;
	wire _w5892_ ;
	wire _w5893_ ;
	wire _w5894_ ;
	wire _w5895_ ;
	wire _w5896_ ;
	wire _w5897_ ;
	wire _w5898_ ;
	wire _w5899_ ;
	wire _w5900_ ;
	wire _w5901_ ;
	wire _w5902_ ;
	wire _w5903_ ;
	wire _w5904_ ;
	wire _w5905_ ;
	wire _w5906_ ;
	wire _w5907_ ;
	wire _w5908_ ;
	wire _w5909_ ;
	wire _w5910_ ;
	wire _w5911_ ;
	wire _w5912_ ;
	wire _w5913_ ;
	wire _w5914_ ;
	wire _w5915_ ;
	wire _w5916_ ;
	wire _w5917_ ;
	wire _w5918_ ;
	wire _w5919_ ;
	wire _w5920_ ;
	wire _w5921_ ;
	wire _w5922_ ;
	wire _w5923_ ;
	wire _w5924_ ;
	wire _w5925_ ;
	wire _w5926_ ;
	wire _w5927_ ;
	wire _w5928_ ;
	wire _w5929_ ;
	wire _w5930_ ;
	wire _w5931_ ;
	wire _w5932_ ;
	wire _w5933_ ;
	wire _w5934_ ;
	wire _w5935_ ;
	wire _w5936_ ;
	wire _w5937_ ;
	wire _w5938_ ;
	wire _w5939_ ;
	wire _w5940_ ;
	wire _w5941_ ;
	wire _w5942_ ;
	wire _w5943_ ;
	wire _w5944_ ;
	wire _w5945_ ;
	wire _w5946_ ;
	wire _w5947_ ;
	wire _w5948_ ;
	wire _w5949_ ;
	wire _w5950_ ;
	wire _w5951_ ;
	wire _w5952_ ;
	wire _w5953_ ;
	wire _w5954_ ;
	wire _w5955_ ;
	wire _w5956_ ;
	wire _w5957_ ;
	wire _w5958_ ;
	wire _w5959_ ;
	wire _w5960_ ;
	wire _w5961_ ;
	wire _w5962_ ;
	wire _w5963_ ;
	wire _w5964_ ;
	wire _w5965_ ;
	wire _w5966_ ;
	wire _w5967_ ;
	wire _w5968_ ;
	wire _w5969_ ;
	wire _w5970_ ;
	wire _w5971_ ;
	wire _w5972_ ;
	wire _w5973_ ;
	wire _w5974_ ;
	wire _w5975_ ;
	wire _w5976_ ;
	wire _w5977_ ;
	wire _w5978_ ;
	wire _w5979_ ;
	wire _w5980_ ;
	wire _w5981_ ;
	wire _w5982_ ;
	wire _w5983_ ;
	wire _w5984_ ;
	wire _w5985_ ;
	wire _w5986_ ;
	wire _w5987_ ;
	wire _w5988_ ;
	wire _w5989_ ;
	wire _w5990_ ;
	wire _w5991_ ;
	wire _w5992_ ;
	wire _w5993_ ;
	wire _w5994_ ;
	wire _w5995_ ;
	wire _w5996_ ;
	wire _w5997_ ;
	wire _w5998_ ;
	wire _w5999_ ;
	wire _w6000_ ;
	wire _w6001_ ;
	wire _w6002_ ;
	wire _w6003_ ;
	wire _w6004_ ;
	wire _w6005_ ;
	wire _w6006_ ;
	wire _w6007_ ;
	wire _w6008_ ;
	wire _w6009_ ;
	wire _w6010_ ;
	wire _w6011_ ;
	wire _w6012_ ;
	wire _w6013_ ;
	wire _w6014_ ;
	wire _w6015_ ;
	wire _w6016_ ;
	wire _w6017_ ;
	wire _w6018_ ;
	wire _w6019_ ;
	wire _w6020_ ;
	wire _w6021_ ;
	wire _w6022_ ;
	wire _w6023_ ;
	wire _w6024_ ;
	wire _w6025_ ;
	wire _w6026_ ;
	wire _w6027_ ;
	wire _w6028_ ;
	wire _w6029_ ;
	wire _w6030_ ;
	wire _w6031_ ;
	wire _w6032_ ;
	wire _w6033_ ;
	wire _w6034_ ;
	wire _w6035_ ;
	wire _w6036_ ;
	wire _w6037_ ;
	wire _w6038_ ;
	wire _w6039_ ;
	wire _w6040_ ;
	wire _w6041_ ;
	wire _w6042_ ;
	wire _w6043_ ;
	wire _w6044_ ;
	wire _w6045_ ;
	wire _w6046_ ;
	wire _w6047_ ;
	wire _w6048_ ;
	wire _w6049_ ;
	wire _w6050_ ;
	wire _w6051_ ;
	wire _w6052_ ;
	wire _w6053_ ;
	wire _w6054_ ;
	wire _w6055_ ;
	wire _w6056_ ;
	wire _w6057_ ;
	wire _w6058_ ;
	wire _w6059_ ;
	wire _w6060_ ;
	wire _w6061_ ;
	wire _w6062_ ;
	wire _w6063_ ;
	wire _w6064_ ;
	wire _w6065_ ;
	wire _w6066_ ;
	wire _w6067_ ;
	wire _w6068_ ;
	wire _w6069_ ;
	wire _w6070_ ;
	wire _w6071_ ;
	wire _w6072_ ;
	wire _w6073_ ;
	wire _w6074_ ;
	wire _w6075_ ;
	wire _w6076_ ;
	wire _w6077_ ;
	wire _w6078_ ;
	wire _w6079_ ;
	wire _w6080_ ;
	wire _w6081_ ;
	wire _w6082_ ;
	wire _w6083_ ;
	wire _w6084_ ;
	wire _w6085_ ;
	wire _w6086_ ;
	wire _w6087_ ;
	wire _w6088_ ;
	wire _w6089_ ;
	wire _w6090_ ;
	wire _w6091_ ;
	wire _w6092_ ;
	wire _w6093_ ;
	wire _w6094_ ;
	wire _w6095_ ;
	wire _w6096_ ;
	wire _w6097_ ;
	wire _w6098_ ;
	wire _w6099_ ;
	wire _w6100_ ;
	wire _w6101_ ;
	wire _w6102_ ;
	wire _w6103_ ;
	wire _w6104_ ;
	wire _w6105_ ;
	wire _w6106_ ;
	wire _w6107_ ;
	wire _w6108_ ;
	wire _w6109_ ;
	wire _w6110_ ;
	wire _w6111_ ;
	wire _w6112_ ;
	wire _w6113_ ;
	wire _w6114_ ;
	wire _w6115_ ;
	wire _w6116_ ;
	wire _w6117_ ;
	wire _w6118_ ;
	wire _w6119_ ;
	wire _w6120_ ;
	wire _w6121_ ;
	wire _w6122_ ;
	wire _w6123_ ;
	wire _w6124_ ;
	wire _w6125_ ;
	wire _w6126_ ;
	wire _w6127_ ;
	wire _w6128_ ;
	wire _w6129_ ;
	wire _w6130_ ;
	wire _w6131_ ;
	wire _w6132_ ;
	wire _w6133_ ;
	wire _w6134_ ;
	wire _w6135_ ;
	wire _w6136_ ;
	wire _w6137_ ;
	wire _w6138_ ;
	wire _w6139_ ;
	wire _w6140_ ;
	wire _w6141_ ;
	wire _w6142_ ;
	wire _w6143_ ;
	wire _w6144_ ;
	wire _w6145_ ;
	wire _w6146_ ;
	wire _w6147_ ;
	wire _w6148_ ;
	wire _w6149_ ;
	wire _w6150_ ;
	wire _w6151_ ;
	wire _w6152_ ;
	wire _w6153_ ;
	wire _w6154_ ;
	wire _w6155_ ;
	wire _w6156_ ;
	wire _w6157_ ;
	wire _w6158_ ;
	wire _w6159_ ;
	wire _w6160_ ;
	wire _w6161_ ;
	wire _w6162_ ;
	wire _w6163_ ;
	wire _w6164_ ;
	wire _w6165_ ;
	wire _w6166_ ;
	wire _w6167_ ;
	wire _w6168_ ;
	wire _w6169_ ;
	wire _w6170_ ;
	wire _w6171_ ;
	wire _w6172_ ;
	wire _w6173_ ;
	wire _w6174_ ;
	wire _w6175_ ;
	wire _w6176_ ;
	wire _w6177_ ;
	wire _w6178_ ;
	wire _w6179_ ;
	wire _w6180_ ;
	wire _w6181_ ;
	wire _w6182_ ;
	wire _w6183_ ;
	wire _w6184_ ;
	wire _w6185_ ;
	wire _w6186_ ;
	wire _w6187_ ;
	wire _w6188_ ;
	wire _w6189_ ;
	wire _w6190_ ;
	wire _w6191_ ;
	wire _w6192_ ;
	wire _w6193_ ;
	wire _w6194_ ;
	wire _w6195_ ;
	wire _w6196_ ;
	wire _w6197_ ;
	wire _w6198_ ;
	wire _w6199_ ;
	wire _w6200_ ;
	wire _w6201_ ;
	wire _w6202_ ;
	wire _w6203_ ;
	wire _w6204_ ;
	wire _w6205_ ;
	wire _w6206_ ;
	wire _w6207_ ;
	wire _w6208_ ;
	wire _w6209_ ;
	wire _w6210_ ;
	wire _w6211_ ;
	wire _w6212_ ;
	wire _w6213_ ;
	wire _w6214_ ;
	wire _w6215_ ;
	wire _w6216_ ;
	wire _w6217_ ;
	wire _w6218_ ;
	wire _w6219_ ;
	wire _w6220_ ;
	wire _w6221_ ;
	wire _w6222_ ;
	wire _w6223_ ;
	wire _w6224_ ;
	wire _w6225_ ;
	wire _w6226_ ;
	wire _w6227_ ;
	wire _w6228_ ;
	wire _w6229_ ;
	wire _w6230_ ;
	wire _w6231_ ;
	wire _w6232_ ;
	wire _w6233_ ;
	wire _w6234_ ;
	wire _w6235_ ;
	wire _w6236_ ;
	wire _w6237_ ;
	wire _w6238_ ;
	wire _w6239_ ;
	wire _w6240_ ;
	wire _w6241_ ;
	wire _w6242_ ;
	wire _w6243_ ;
	wire _w6244_ ;
	wire _w6245_ ;
	wire _w6246_ ;
	wire _w6247_ ;
	wire _w6248_ ;
	wire _w6249_ ;
	wire _w6250_ ;
	wire _w6251_ ;
	wire _w6252_ ;
	wire _w6253_ ;
	wire _w6254_ ;
	wire _w6255_ ;
	wire _w6256_ ;
	wire _w6257_ ;
	wire _w6258_ ;
	wire _w6259_ ;
	wire _w6260_ ;
	wire _w6261_ ;
	wire _w6262_ ;
	wire _w6263_ ;
	wire _w6264_ ;
	wire _w6265_ ;
	wire _w6266_ ;
	wire _w6267_ ;
	wire _w6268_ ;
	wire _w6269_ ;
	wire _w6270_ ;
	wire _w6271_ ;
	wire _w6272_ ;
	wire _w6273_ ;
	wire _w6274_ ;
	wire _w6275_ ;
	wire _w6276_ ;
	wire _w6277_ ;
	wire _w6278_ ;
	wire _w6279_ ;
	wire _w6280_ ;
	wire _w6281_ ;
	wire _w6282_ ;
	wire _w6283_ ;
	wire _w6284_ ;
	wire _w6285_ ;
	wire _w6286_ ;
	wire _w6287_ ;
	wire _w6288_ ;
	wire _w6289_ ;
	wire _w6290_ ;
	wire _w6291_ ;
	wire _w6292_ ;
	wire _w6293_ ;
	wire _w6294_ ;
	wire _w6295_ ;
	wire _w6296_ ;
	wire _w6297_ ;
	wire _w6298_ ;
	wire _w6299_ ;
	wire _w6300_ ;
	wire _w6301_ ;
	wire _w6302_ ;
	wire _w6303_ ;
	wire _w6304_ ;
	wire _w6305_ ;
	wire _w6306_ ;
	wire _w6307_ ;
	wire _w6308_ ;
	wire _w6309_ ;
	wire _w6310_ ;
	wire _w6311_ ;
	wire _w6312_ ;
	wire _w6313_ ;
	wire _w6314_ ;
	wire _w6315_ ;
	wire _w6316_ ;
	wire _w6317_ ;
	wire _w6318_ ;
	wire _w6319_ ;
	wire _w6320_ ;
	wire _w6321_ ;
	wire _w6322_ ;
	wire _w6323_ ;
	wire _w6324_ ;
	wire _w6325_ ;
	wire _w6326_ ;
	wire _w6327_ ;
	wire _w6328_ ;
	wire _w6329_ ;
	wire _w6330_ ;
	wire _w6331_ ;
	wire _w6332_ ;
	wire _w6333_ ;
	wire _w6334_ ;
	wire _w6335_ ;
	wire _w6336_ ;
	wire _w6337_ ;
	wire _w6338_ ;
	wire _w6339_ ;
	wire _w6340_ ;
	wire _w6341_ ;
	wire _w6342_ ;
	wire _w6343_ ;
	wire _w6344_ ;
	wire _w6345_ ;
	wire _w6346_ ;
	wire _w6347_ ;
	wire _w6348_ ;
	wire _w6349_ ;
	wire _w6350_ ;
	wire _w6351_ ;
	wire _w6352_ ;
	wire _w6353_ ;
	wire _w6354_ ;
	wire _w6355_ ;
	wire _w6356_ ;
	wire _w6357_ ;
	wire _w6358_ ;
	wire _w6359_ ;
	wire _w6360_ ;
	wire _w6361_ ;
	wire _w6362_ ;
	wire _w6363_ ;
	wire _w6364_ ;
	wire _w6365_ ;
	wire _w6366_ ;
	wire _w6367_ ;
	wire _w6368_ ;
	wire _w6369_ ;
	wire _w6370_ ;
	wire _w6371_ ;
	wire _w6372_ ;
	wire _w6373_ ;
	wire _w6374_ ;
	wire _w6375_ ;
	wire _w6376_ ;
	wire _w6377_ ;
	wire _w6378_ ;
	wire _w6379_ ;
	wire _w6380_ ;
	wire _w6381_ ;
	wire _w6382_ ;
	wire _w6383_ ;
	wire _w6384_ ;
	wire _w6385_ ;
	wire _w6386_ ;
	wire _w6387_ ;
	wire _w6388_ ;
	wire _w6389_ ;
	wire _w6390_ ;
	wire _w6391_ ;
	wire _w6392_ ;
	wire _w6393_ ;
	wire _w6394_ ;
	wire _w6395_ ;
	wire _w6396_ ;
	wire _w6397_ ;
	wire _w6398_ ;
	wire _w6399_ ;
	wire _w6400_ ;
	wire _w6401_ ;
	wire _w6402_ ;
	wire _w6403_ ;
	wire _w6404_ ;
	wire _w6405_ ;
	wire _w6406_ ;
	wire _w6407_ ;
	wire _w6408_ ;
	wire _w6409_ ;
	wire _w6410_ ;
	wire _w6411_ ;
	wire _w6412_ ;
	wire _w6413_ ;
	wire _w6414_ ;
	wire _w6415_ ;
	wire _w6416_ ;
	wire _w6417_ ;
	wire _w6418_ ;
	wire _w6419_ ;
	wire _w6420_ ;
	wire _w6421_ ;
	wire _w6422_ ;
	wire _w6423_ ;
	wire _w6424_ ;
	wire _w6425_ ;
	wire _w6426_ ;
	wire _w6427_ ;
	wire _w6428_ ;
	wire _w6429_ ;
	wire _w6430_ ;
	wire _w6431_ ;
	wire _w6432_ ;
	wire _w6433_ ;
	wire _w6434_ ;
	wire _w6435_ ;
	wire _w6436_ ;
	wire _w6437_ ;
	wire _w6438_ ;
	wire _w6439_ ;
	wire _w6440_ ;
	wire _w6441_ ;
	wire _w6442_ ;
	wire _w6443_ ;
	wire _w6444_ ;
	wire _w6445_ ;
	wire _w6446_ ;
	wire _w6447_ ;
	wire _w6448_ ;
	wire _w6449_ ;
	wire _w6450_ ;
	wire _w6451_ ;
	wire _w6452_ ;
	wire _w6453_ ;
	wire _w6454_ ;
	wire _w6455_ ;
	wire _w6456_ ;
	wire _w6457_ ;
	wire _w6458_ ;
	wire _w6459_ ;
	wire _w6460_ ;
	wire _w6461_ ;
	wire _w6462_ ;
	wire _w6463_ ;
	wire _w6464_ ;
	wire _w6465_ ;
	wire _w6466_ ;
	wire _w6467_ ;
	wire _w6468_ ;
	wire _w6469_ ;
	wire _w6470_ ;
	wire _w6471_ ;
	wire _w6472_ ;
	wire _w6473_ ;
	wire _w6474_ ;
	wire _w6475_ ;
	wire _w6476_ ;
	wire _w6477_ ;
	wire _w6478_ ;
	wire _w6479_ ;
	wire _w6480_ ;
	wire _w6481_ ;
	wire _w6482_ ;
	wire _w6483_ ;
	wire _w6484_ ;
	wire _w6485_ ;
	wire _w6486_ ;
	wire _w6487_ ;
	wire _w6488_ ;
	wire _w6489_ ;
	wire _w6490_ ;
	wire _w6491_ ;
	wire _w6492_ ;
	wire _w6493_ ;
	wire _w6494_ ;
	wire _w6495_ ;
	wire _w6496_ ;
	wire _w6497_ ;
	wire _w6498_ ;
	wire _w6499_ ;
	wire _w6500_ ;
	wire _w6501_ ;
	wire _w6502_ ;
	wire _w6503_ ;
	wire _w6504_ ;
	wire _w6505_ ;
	wire _w6506_ ;
	wire _w6507_ ;
	wire _w6508_ ;
	wire _w6509_ ;
	wire _w6510_ ;
	wire _w6511_ ;
	wire _w6512_ ;
	wire _w6513_ ;
	wire _w6514_ ;
	wire _w6515_ ;
	wire _w6516_ ;
	wire _w6517_ ;
	wire _w6518_ ;
	wire _w6519_ ;
	wire _w6520_ ;
	wire _w6521_ ;
	wire _w6522_ ;
	wire _w6523_ ;
	wire _w6524_ ;
	wire _w6525_ ;
	wire _w6526_ ;
	wire _w6527_ ;
	wire _w6528_ ;
	wire _w6529_ ;
	wire _w6530_ ;
	wire _w6531_ ;
	wire _w6532_ ;
	wire _w6533_ ;
	wire _w6534_ ;
	wire _w6535_ ;
	wire _w6536_ ;
	wire _w6537_ ;
	wire _w6538_ ;
	wire _w6539_ ;
	wire _w6540_ ;
	wire _w6541_ ;
	wire _w6542_ ;
	wire _w6543_ ;
	wire _w6544_ ;
	wire _w6545_ ;
	wire _w6546_ ;
	wire _w6547_ ;
	wire _w6548_ ;
	wire _w6549_ ;
	wire _w6550_ ;
	wire _w6551_ ;
	wire _w6552_ ;
	wire _w6553_ ;
	wire _w6554_ ;
	wire _w6555_ ;
	wire _w6556_ ;
	wire _w6557_ ;
	wire _w6558_ ;
	wire _w6559_ ;
	wire _w6560_ ;
	wire _w6561_ ;
	wire _w6562_ ;
	wire _w6563_ ;
	wire _w6564_ ;
	wire _w6565_ ;
	wire _w6566_ ;
	wire _w6567_ ;
	wire _w6568_ ;
	wire _w6569_ ;
	wire _w6570_ ;
	wire _w6571_ ;
	wire _w6572_ ;
	wire _w6573_ ;
	wire _w6574_ ;
	wire _w6575_ ;
	wire _w6576_ ;
	wire _w6577_ ;
	wire _w6578_ ;
	wire _w6579_ ;
	wire _w6580_ ;
	wire _w6581_ ;
	wire _w6582_ ;
	wire _w6583_ ;
	wire _w6584_ ;
	wire _w6585_ ;
	wire _w6586_ ;
	wire _w6587_ ;
	wire _w6588_ ;
	wire _w6589_ ;
	wire _w6590_ ;
	wire _w6591_ ;
	wire _w6592_ ;
	wire _w6593_ ;
	wire _w6594_ ;
	wire _w6595_ ;
	wire _w6596_ ;
	wire _w6597_ ;
	wire _w6598_ ;
	wire _w6599_ ;
	wire _w6600_ ;
	wire _w6601_ ;
	wire _w6602_ ;
	wire _w6603_ ;
	wire _w6604_ ;
	wire _w6605_ ;
	wire _w6606_ ;
	wire _w6607_ ;
	wire _w6608_ ;
	wire _w6609_ ;
	wire _w6610_ ;
	wire _w6611_ ;
	wire _w6612_ ;
	wire _w6613_ ;
	wire _w6614_ ;
	wire _w6615_ ;
	wire _w6616_ ;
	wire _w6617_ ;
	wire _w6618_ ;
	wire _w6619_ ;
	wire _w6620_ ;
	wire _w6621_ ;
	wire _w6622_ ;
	wire _w6623_ ;
	wire _w6624_ ;
	wire _w6625_ ;
	wire _w6626_ ;
	wire _w6627_ ;
	wire _w6628_ ;
	wire _w6629_ ;
	wire _w6630_ ;
	wire _w6631_ ;
	wire _w6632_ ;
	wire _w6633_ ;
	wire _w6634_ ;
	wire _w6635_ ;
	wire _w6636_ ;
	wire _w6637_ ;
	wire _w6638_ ;
	wire _w6639_ ;
	wire _w6640_ ;
	wire _w6641_ ;
	wire _w6642_ ;
	wire _w6643_ ;
	wire _w6644_ ;
	wire _w6645_ ;
	wire _w6646_ ;
	wire _w6647_ ;
	wire _w6648_ ;
	wire _w6649_ ;
	wire _w6650_ ;
	wire _w6651_ ;
	wire _w6652_ ;
	wire _w6653_ ;
	wire _w6654_ ;
	wire _w6655_ ;
	wire _w6656_ ;
	wire _w6657_ ;
	wire _w6658_ ;
	wire _w6659_ ;
	wire _w6660_ ;
	wire _w6661_ ;
	wire _w6662_ ;
	wire _w6663_ ;
	wire _w6664_ ;
	wire _w6665_ ;
	wire _w6666_ ;
	wire _w6667_ ;
	wire _w6668_ ;
	wire _w6669_ ;
	wire _w6670_ ;
	wire _w6671_ ;
	wire _w6672_ ;
	wire _w6673_ ;
	wire _w6674_ ;
	wire _w6675_ ;
	wire _w6676_ ;
	wire _w6677_ ;
	wire _w6678_ ;
	wire _w6679_ ;
	wire _w6680_ ;
	wire _w6681_ ;
	wire _w6682_ ;
	wire _w6683_ ;
	wire _w6684_ ;
	wire _w6685_ ;
	wire _w6686_ ;
	wire _w6687_ ;
	wire _w6688_ ;
	wire _w6689_ ;
	wire _w6690_ ;
	wire _w6691_ ;
	wire _w6692_ ;
	wire _w6693_ ;
	wire _w6694_ ;
	wire _w6695_ ;
	wire _w6696_ ;
	wire _w6697_ ;
	wire _w6698_ ;
	wire _w6699_ ;
	wire _w6700_ ;
	wire _w6701_ ;
	wire _w6702_ ;
	wire _w6703_ ;
	wire _w6704_ ;
	wire _w6705_ ;
	wire _w6706_ ;
	wire _w6707_ ;
	wire _w6708_ ;
	wire _w6709_ ;
	wire _w6710_ ;
	wire _w6711_ ;
	wire _w6712_ ;
	wire _w6713_ ;
	wire _w6714_ ;
	wire _w6715_ ;
	wire _w6716_ ;
	wire _w6717_ ;
	wire _w6718_ ;
	wire _w6719_ ;
	wire _w6720_ ;
	wire _w6721_ ;
	wire _w6722_ ;
	wire _w6723_ ;
	wire _w6724_ ;
	wire _w6725_ ;
	wire _w6726_ ;
	wire _w6727_ ;
	wire _w6728_ ;
	wire _w6729_ ;
	wire _w6730_ ;
	wire _w6731_ ;
	wire _w6732_ ;
	wire _w6733_ ;
	wire _w6734_ ;
	wire _w6735_ ;
	wire _w6736_ ;
	wire _w6737_ ;
	wire _w6738_ ;
	wire _w6739_ ;
	wire _w6740_ ;
	wire _w6741_ ;
	wire _w6742_ ;
	wire _w6743_ ;
	wire _w6744_ ;
	wire _w6745_ ;
	wire _w6746_ ;
	wire _w6747_ ;
	wire _w6748_ ;
	wire _w6749_ ;
	wire _w6750_ ;
	wire _w6751_ ;
	wire _w6752_ ;
	wire _w6753_ ;
	wire _w6754_ ;
	wire _w6755_ ;
	wire _w6756_ ;
	wire _w6757_ ;
	wire _w6758_ ;
	wire _w6759_ ;
	wire _w6760_ ;
	wire _w6761_ ;
	wire _w6762_ ;
	wire _w6763_ ;
	wire _w6764_ ;
	wire _w6765_ ;
	wire _w6766_ ;
	wire _w6767_ ;
	wire _w6768_ ;
	wire _w6769_ ;
	wire _w6770_ ;
	wire _w6771_ ;
	wire _w6772_ ;
	wire _w6773_ ;
	wire _w6774_ ;
	wire _w6775_ ;
	wire _w6776_ ;
	wire _w6777_ ;
	wire _w6778_ ;
	wire _w6779_ ;
	wire _w6780_ ;
	wire _w6781_ ;
	wire _w6782_ ;
	wire _w6783_ ;
	wire _w6784_ ;
	wire _w6785_ ;
	wire _w6786_ ;
	wire _w6787_ ;
	wire _w6788_ ;
	wire _w6789_ ;
	wire _w6790_ ;
	wire _w6791_ ;
	wire _w6792_ ;
	wire _w6793_ ;
	wire _w6794_ ;
	wire _w6795_ ;
	wire _w6796_ ;
	wire _w6797_ ;
	wire _w6798_ ;
	wire _w6799_ ;
	wire _w6800_ ;
	wire _w6801_ ;
	wire _w6802_ ;
	wire _w6803_ ;
	wire _w6804_ ;
	wire _w6805_ ;
	wire _w6806_ ;
	wire _w6807_ ;
	wire _w6808_ ;
	wire _w6809_ ;
	wire _w6810_ ;
	wire _w6811_ ;
	wire _w6812_ ;
	wire _w6813_ ;
	wire _w6814_ ;
	wire _w6815_ ;
	wire _w6816_ ;
	wire _w6817_ ;
	wire _w6818_ ;
	wire _w6819_ ;
	wire _w6820_ ;
	wire _w6821_ ;
	wire _w6822_ ;
	wire _w6823_ ;
	wire _w6824_ ;
	wire _w6825_ ;
	wire _w6826_ ;
	wire _w6827_ ;
	wire _w6828_ ;
	wire _w6829_ ;
	wire _w6830_ ;
	wire _w6831_ ;
	wire _w6832_ ;
	wire _w6833_ ;
	wire _w6834_ ;
	wire _w6835_ ;
	wire _w6836_ ;
	wire _w6837_ ;
	wire _w6838_ ;
	wire _w6839_ ;
	wire _w6840_ ;
	wire _w6841_ ;
	wire _w6842_ ;
	wire _w6843_ ;
	wire _w6844_ ;
	wire _w6845_ ;
	wire _w6846_ ;
	wire _w6847_ ;
	wire _w6848_ ;
	wire _w6849_ ;
	wire _w6850_ ;
	wire _w6851_ ;
	wire _w6852_ ;
	wire _w6853_ ;
	wire _w6854_ ;
	wire _w6855_ ;
	wire _w6856_ ;
	wire _w6857_ ;
	wire _w6858_ ;
	wire _w6859_ ;
	wire _w6860_ ;
	wire _w6861_ ;
	wire _w6862_ ;
	wire _w6863_ ;
	wire _w6864_ ;
	wire _w6865_ ;
	wire _w6866_ ;
	wire _w6867_ ;
	wire _w6868_ ;
	wire _w6869_ ;
	wire _w6870_ ;
	wire _w6871_ ;
	wire _w6872_ ;
	wire _w6873_ ;
	wire _w6874_ ;
	wire _w6875_ ;
	wire _w6876_ ;
	wire _w6877_ ;
	wire _w6878_ ;
	wire _w6879_ ;
	wire _w6880_ ;
	wire _w6881_ ;
	wire _w6882_ ;
	wire _w6883_ ;
	wire _w6884_ ;
	wire _w6885_ ;
	wire _w6886_ ;
	wire _w6887_ ;
	wire _w6888_ ;
	wire _w6889_ ;
	wire _w6890_ ;
	wire _w6891_ ;
	wire _w6892_ ;
	wire _w6893_ ;
	wire _w6894_ ;
	wire _w6895_ ;
	wire _w6896_ ;
	wire _w6897_ ;
	wire _w6898_ ;
	wire _w6899_ ;
	wire _w6900_ ;
	wire _w6901_ ;
	wire _w6902_ ;
	wire _w6903_ ;
	wire _w6904_ ;
	wire _w6905_ ;
	wire _w6906_ ;
	wire _w6907_ ;
	wire _w6908_ ;
	wire _w6909_ ;
	wire _w6910_ ;
	wire _w6911_ ;
	wire _w6912_ ;
	wire _w6913_ ;
	wire _w6914_ ;
	wire _w6915_ ;
	wire _w6916_ ;
	wire _w6917_ ;
	wire _w6918_ ;
	wire _w6919_ ;
	wire _w6920_ ;
	wire _w6921_ ;
	wire _w6922_ ;
	wire _w6923_ ;
	wire _w6924_ ;
	wire _w6925_ ;
	wire _w6926_ ;
	wire _w6927_ ;
	wire _w6928_ ;
	wire _w6929_ ;
	wire _w6930_ ;
	wire _w6931_ ;
	wire _w6932_ ;
	wire _w6933_ ;
	wire _w6934_ ;
	wire _w6935_ ;
	wire _w6936_ ;
	wire _w6937_ ;
	wire _w6938_ ;
	wire _w6939_ ;
	wire _w6940_ ;
	wire _w6941_ ;
	wire _w6942_ ;
	wire _w6943_ ;
	wire _w6944_ ;
	wire _w6945_ ;
	wire _w6946_ ;
	wire _w6947_ ;
	wire _w6948_ ;
	wire _w6949_ ;
	wire _w6950_ ;
	wire _w6951_ ;
	wire _w6952_ ;
	wire _w6953_ ;
	wire _w6954_ ;
	wire _w6955_ ;
	wire _w6956_ ;
	wire _w6957_ ;
	wire _w6958_ ;
	wire _w6959_ ;
	wire _w6960_ ;
	wire _w6961_ ;
	wire _w6962_ ;
	wire _w6963_ ;
	wire _w6964_ ;
	wire _w6965_ ;
	wire _w6966_ ;
	wire _w6967_ ;
	wire _w6968_ ;
	wire _w6969_ ;
	wire _w6970_ ;
	wire _w6971_ ;
	wire _w6972_ ;
	wire _w6973_ ;
	wire _w6974_ ;
	wire _w6975_ ;
	wire _w6976_ ;
	wire _w6977_ ;
	wire _w6978_ ;
	wire _w6979_ ;
	wire _w6980_ ;
	wire _w6981_ ;
	wire _w6982_ ;
	wire _w6983_ ;
	wire _w6984_ ;
	wire _w6985_ ;
	wire _w6986_ ;
	wire _w6987_ ;
	wire _w6988_ ;
	wire _w6989_ ;
	wire _w6990_ ;
	wire _w6991_ ;
	wire _w6992_ ;
	wire _w6993_ ;
	wire _w6994_ ;
	wire _w6995_ ;
	wire _w6996_ ;
	wire _w6997_ ;
	wire _w6998_ ;
	wire _w6999_ ;
	wire _w7000_ ;
	wire _w7001_ ;
	wire _w7002_ ;
	wire _w7003_ ;
	wire _w7004_ ;
	wire _w7005_ ;
	wire _w7006_ ;
	wire _w7007_ ;
	wire _w7008_ ;
	wire _w7009_ ;
	wire _w7010_ ;
	wire _w7011_ ;
	wire _w7012_ ;
	wire _w7013_ ;
	wire _w7014_ ;
	wire _w7015_ ;
	wire _w7016_ ;
	wire _w7017_ ;
	wire _w7018_ ;
	wire _w7019_ ;
	wire _w7020_ ;
	wire _w7021_ ;
	wire _w7022_ ;
	wire _w7023_ ;
	wire _w7024_ ;
	wire _w7025_ ;
	wire _w7026_ ;
	wire _w7027_ ;
	wire _w7028_ ;
	wire _w7029_ ;
	wire _w7030_ ;
	wire _w7031_ ;
	wire _w7032_ ;
	wire _w7033_ ;
	wire _w7034_ ;
	wire _w7035_ ;
	wire _w7036_ ;
	wire _w7037_ ;
	wire _w7038_ ;
	wire _w7039_ ;
	wire _w7040_ ;
	wire _w7041_ ;
	wire _w7042_ ;
	wire _w7043_ ;
	wire _w7044_ ;
	wire _w7045_ ;
	wire _w7046_ ;
	wire _w7047_ ;
	wire _w7048_ ;
	wire _w7049_ ;
	wire _w7050_ ;
	wire _w7051_ ;
	wire _w7052_ ;
	wire _w7053_ ;
	wire _w7054_ ;
	wire _w7055_ ;
	wire _w7056_ ;
	wire _w7057_ ;
	wire _w7058_ ;
	wire _w7059_ ;
	wire _w7060_ ;
	wire _w7061_ ;
	wire _w7062_ ;
	wire _w7063_ ;
	wire _w7064_ ;
	wire _w7065_ ;
	wire _w7066_ ;
	wire _w7067_ ;
	wire _w7068_ ;
	wire _w7069_ ;
	wire _w7070_ ;
	wire _w7071_ ;
	wire _w7072_ ;
	wire _w7073_ ;
	wire _w7074_ ;
	wire _w7075_ ;
	wire _w7076_ ;
	wire _w7077_ ;
	wire _w7078_ ;
	wire _w7079_ ;
	wire _w7080_ ;
	wire _w7081_ ;
	wire _w7082_ ;
	wire _w7083_ ;
	wire _w7084_ ;
	wire _w7085_ ;
	wire _w7086_ ;
	wire _w7087_ ;
	wire _w7088_ ;
	wire _w7089_ ;
	wire _w7090_ ;
	wire _w7091_ ;
	wire _w7092_ ;
	wire _w7093_ ;
	wire _w7094_ ;
	wire _w7095_ ;
	wire _w7096_ ;
	wire _w7097_ ;
	wire _w7098_ ;
	wire _w7099_ ;
	wire _w7100_ ;
	wire _w7101_ ;
	wire _w7102_ ;
	wire _w7103_ ;
	wire _w7104_ ;
	wire _w7105_ ;
	wire _w7106_ ;
	wire _w7107_ ;
	wire _w7108_ ;
	wire _w7109_ ;
	wire _w7110_ ;
	wire _w7111_ ;
	wire _w7112_ ;
	wire _w7113_ ;
	wire _w7114_ ;
	wire _w7115_ ;
	wire _w7116_ ;
	wire _w7117_ ;
	wire _w7118_ ;
	wire _w7119_ ;
	wire _w7120_ ;
	wire _w7121_ ;
	wire _w7122_ ;
	wire _w7123_ ;
	wire _w7124_ ;
	wire _w7125_ ;
	wire _w7126_ ;
	wire _w7127_ ;
	wire _w7128_ ;
	wire _w7129_ ;
	wire _w7130_ ;
	wire _w7131_ ;
	wire _w7132_ ;
	wire _w7133_ ;
	wire _w7134_ ;
	wire _w7135_ ;
	wire _w7136_ ;
	wire _w7137_ ;
	wire _w7138_ ;
	wire _w7139_ ;
	wire _w7140_ ;
	wire _w7141_ ;
	wire _w7142_ ;
	wire _w7143_ ;
	wire _w7144_ ;
	wire _w7145_ ;
	wire _w7146_ ;
	wire _w7147_ ;
	wire _w7148_ ;
	wire _w7149_ ;
	wire _w7150_ ;
	wire _w7151_ ;
	wire _w7152_ ;
	wire _w7153_ ;
	wire _w7154_ ;
	wire _w7155_ ;
	wire _w7156_ ;
	wire _w7157_ ;
	wire _w7158_ ;
	wire _w7159_ ;
	wire _w7160_ ;
	wire _w7161_ ;
	wire _w7162_ ;
	wire _w7163_ ;
	wire _w7164_ ;
	wire _w7165_ ;
	wire _w7166_ ;
	wire _w7167_ ;
	wire _w7168_ ;
	wire _w7169_ ;
	wire _w7170_ ;
	wire _w7171_ ;
	wire _w7172_ ;
	wire _w7173_ ;
	wire _w7174_ ;
	wire _w7175_ ;
	wire _w7176_ ;
	wire _w7177_ ;
	wire _w7178_ ;
	wire _w7179_ ;
	wire _w7180_ ;
	wire _w7181_ ;
	wire _w7182_ ;
	wire _w7183_ ;
	wire _w7184_ ;
	wire _w7185_ ;
	wire _w7186_ ;
	wire _w7187_ ;
	wire _w7188_ ;
	wire _w7189_ ;
	wire _w7190_ ;
	wire _w7191_ ;
	wire _w7192_ ;
	wire _w7193_ ;
	wire _w7194_ ;
	wire _w7195_ ;
	wire _w7196_ ;
	wire _w7197_ ;
	wire _w7198_ ;
	wire _w7199_ ;
	wire _w7200_ ;
	wire _w7201_ ;
	wire _w7202_ ;
	wire _w7203_ ;
	wire _w7204_ ;
	wire _w7205_ ;
	wire _w7206_ ;
	wire _w7207_ ;
	wire _w7208_ ;
	wire _w7209_ ;
	wire _w7210_ ;
	wire _w7211_ ;
	wire _w7212_ ;
	wire _w7213_ ;
	wire _w7214_ ;
	wire _w7215_ ;
	wire _w7216_ ;
	wire _w7217_ ;
	wire _w7218_ ;
	wire _w7219_ ;
	wire _w7220_ ;
	wire _w7221_ ;
	wire _w7222_ ;
	wire _w7223_ ;
	wire _w7224_ ;
	wire _w7225_ ;
	wire _w7226_ ;
	wire _w7227_ ;
	wire _w7228_ ;
	wire _w7229_ ;
	wire _w7230_ ;
	wire _w7231_ ;
	wire _w7232_ ;
	wire _w7233_ ;
	wire _w7234_ ;
	wire _w7235_ ;
	wire _w7236_ ;
	wire _w7237_ ;
	wire _w7238_ ;
	wire _w7239_ ;
	wire _w7240_ ;
	wire _w7241_ ;
	wire _w7242_ ;
	wire _w7243_ ;
	wire _w7244_ ;
	wire _w7245_ ;
	wire _w7246_ ;
	wire _w7247_ ;
	wire _w7248_ ;
	wire _w7249_ ;
	wire _w7250_ ;
	wire _w7251_ ;
	wire _w7252_ ;
	wire _w7253_ ;
	wire _w7254_ ;
	wire _w7255_ ;
	wire _w7256_ ;
	wire _w7257_ ;
	wire _w7258_ ;
	wire _w7259_ ;
	wire _w7260_ ;
	wire _w7261_ ;
	wire _w7262_ ;
	wire _w7263_ ;
	wire _w7264_ ;
	wire _w7265_ ;
	wire _w7266_ ;
	wire _w7267_ ;
	wire _w7268_ ;
	wire _w7269_ ;
	wire _w7270_ ;
	wire _w7271_ ;
	wire _w7272_ ;
	wire _w7273_ ;
	wire _w7274_ ;
	wire _w7275_ ;
	wire _w7276_ ;
	wire _w7277_ ;
	wire _w7278_ ;
	wire _w7279_ ;
	wire _w7280_ ;
	wire _w7281_ ;
	wire _w7282_ ;
	wire _w7283_ ;
	wire _w7284_ ;
	wire _w7285_ ;
	wire _w7286_ ;
	wire _w7287_ ;
	wire _w7288_ ;
	wire _w7289_ ;
	wire _w7290_ ;
	wire _w7291_ ;
	wire _w7292_ ;
	wire _w7293_ ;
	wire _w7294_ ;
	wire _w7295_ ;
	wire _w7296_ ;
	wire _w7297_ ;
	wire _w7298_ ;
	wire _w7299_ ;
	wire _w7300_ ;
	wire _w7301_ ;
	wire _w7302_ ;
	wire _w7303_ ;
	wire _w7304_ ;
	wire _w7305_ ;
	wire _w7306_ ;
	wire _w7307_ ;
	wire _w7308_ ;
	wire _w7309_ ;
	wire _w7310_ ;
	wire _w7311_ ;
	wire _w7312_ ;
	wire _w7313_ ;
	wire _w7314_ ;
	wire _w7315_ ;
	wire _w7316_ ;
	wire _w7317_ ;
	wire _w7318_ ;
	wire _w7319_ ;
	wire _w7320_ ;
	wire _w7321_ ;
	wire _w7322_ ;
	wire _w7323_ ;
	wire _w7324_ ;
	wire _w7325_ ;
	wire _w7326_ ;
	wire _w7327_ ;
	wire _w7328_ ;
	wire _w7329_ ;
	wire _w7330_ ;
	wire _w7331_ ;
	wire _w7332_ ;
	wire _w7333_ ;
	wire _w7334_ ;
	wire _w7335_ ;
	wire _w7336_ ;
	wire _w7337_ ;
	wire _w7338_ ;
	wire _w7339_ ;
	wire _w7340_ ;
	wire _w7341_ ;
	wire _w7342_ ;
	wire _w7343_ ;
	wire _w7344_ ;
	wire _w7345_ ;
	wire _w7346_ ;
	wire _w7347_ ;
	wire _w7348_ ;
	wire _w7349_ ;
	wire _w7350_ ;
	wire _w7351_ ;
	wire _w7352_ ;
	wire _w7353_ ;
	wire _w7354_ ;
	wire _w7355_ ;
	wire _w7356_ ;
	wire _w7357_ ;
	wire _w7358_ ;
	wire _w7359_ ;
	wire _w7360_ ;
	wire _w7361_ ;
	wire _w7362_ ;
	wire _w7363_ ;
	wire _w7364_ ;
	wire _w7365_ ;
	wire _w7366_ ;
	wire _w7367_ ;
	wire _w7368_ ;
	wire _w7369_ ;
	wire _w7370_ ;
	wire _w7371_ ;
	wire _w7372_ ;
	wire _w7373_ ;
	wire _w7374_ ;
	wire _w7375_ ;
	wire _w7376_ ;
	wire _w7377_ ;
	wire _w7378_ ;
	wire _w7379_ ;
	wire _w7380_ ;
	wire _w7381_ ;
	wire _w7382_ ;
	wire _w7383_ ;
	wire _w7384_ ;
	wire _w7385_ ;
	wire _w7386_ ;
	wire _w7387_ ;
	wire _w7388_ ;
	wire _w7389_ ;
	wire _w7390_ ;
	wire _w7391_ ;
	wire _w7392_ ;
	wire _w7393_ ;
	wire _w7394_ ;
	wire _w7395_ ;
	wire _w7396_ ;
	wire _w7397_ ;
	wire _w7398_ ;
	wire _w7399_ ;
	wire _w7400_ ;
	wire _w7401_ ;
	wire _w7402_ ;
	wire _w7403_ ;
	wire _w7404_ ;
	wire _w7405_ ;
	wire _w7406_ ;
	wire _w7407_ ;
	wire _w7408_ ;
	wire _w7409_ ;
	wire _w7410_ ;
	wire _w7411_ ;
	wire _w7412_ ;
	wire _w7413_ ;
	wire _w7414_ ;
	wire _w7415_ ;
	wire _w7416_ ;
	wire _w7417_ ;
	wire _w7418_ ;
	wire _w7419_ ;
	wire _w7420_ ;
	wire _w7421_ ;
	wire _w7422_ ;
	wire _w7423_ ;
	wire _w7424_ ;
	wire _w7425_ ;
	wire _w7426_ ;
	wire _w7427_ ;
	wire _w7428_ ;
	wire _w7429_ ;
	wire _w7430_ ;
	wire _w7431_ ;
	wire _w7432_ ;
	wire _w7433_ ;
	wire _w7434_ ;
	wire _w7435_ ;
	wire _w7436_ ;
	wire _w7437_ ;
	wire _w7438_ ;
	wire _w7439_ ;
	wire _w7440_ ;
	wire _w7441_ ;
	wire _w7442_ ;
	wire _w7443_ ;
	wire _w7444_ ;
	wire _w7445_ ;
	wire _w7446_ ;
	wire _w7447_ ;
	wire _w7448_ ;
	wire _w7449_ ;
	wire _w7450_ ;
	wire _w7451_ ;
	wire _w7452_ ;
	wire _w7453_ ;
	wire _w7454_ ;
	wire _w7455_ ;
	wire _w7456_ ;
	wire _w7457_ ;
	wire _w7458_ ;
	wire _w7459_ ;
	wire _w7460_ ;
	wire _w7461_ ;
	wire _w7462_ ;
	wire _w7463_ ;
	wire _w7464_ ;
	wire _w7465_ ;
	wire _w7466_ ;
	wire _w7467_ ;
	wire _w7468_ ;
	wire _w7469_ ;
	wire _w7470_ ;
	wire _w7471_ ;
	wire _w7472_ ;
	wire _w7473_ ;
	wire _w7474_ ;
	wire _w7475_ ;
	wire _w7476_ ;
	wire _w7477_ ;
	wire _w7478_ ;
	wire _w7479_ ;
	wire _w7480_ ;
	wire _w7481_ ;
	wire _w7482_ ;
	wire _w7483_ ;
	wire _w7484_ ;
	wire _w7485_ ;
	wire _w7486_ ;
	wire _w7487_ ;
	wire _w7488_ ;
	wire _w7489_ ;
	wire _w7490_ ;
	wire _w7491_ ;
	wire _w7492_ ;
	wire _w7493_ ;
	wire _w7494_ ;
	wire _w7495_ ;
	wire _w7496_ ;
	wire _w7497_ ;
	wire _w7498_ ;
	wire _w7499_ ;
	wire _w7500_ ;
	wire _w7501_ ;
	wire _w7502_ ;
	wire _w7503_ ;
	wire _w7504_ ;
	wire _w7505_ ;
	wire _w7506_ ;
	wire _w7507_ ;
	wire _w7508_ ;
	wire _w7509_ ;
	wire _w7510_ ;
	wire _w7511_ ;
	wire _w7512_ ;
	wire _w7513_ ;
	wire _w7514_ ;
	wire _w7515_ ;
	wire _w7516_ ;
	wire _w7517_ ;
	wire _w7518_ ;
	wire _w7519_ ;
	wire _w7520_ ;
	wire _w7521_ ;
	wire _w7522_ ;
	wire _w7523_ ;
	wire _w7524_ ;
	wire _w7525_ ;
	wire _w7526_ ;
	wire _w7527_ ;
	wire _w7528_ ;
	wire _w7529_ ;
	wire _w7530_ ;
	wire _w7531_ ;
	wire _w7532_ ;
	wire _w7533_ ;
	wire _w7534_ ;
	wire _w7535_ ;
	wire _w7536_ ;
	wire _w7537_ ;
	wire _w7538_ ;
	wire _w7539_ ;
	wire _w7540_ ;
	wire _w7541_ ;
	wire _w7542_ ;
	wire _w7543_ ;
	wire _w7544_ ;
	wire _w7545_ ;
	wire _w7546_ ;
	wire _w7547_ ;
	wire _w7548_ ;
	wire _w7549_ ;
	wire _w7550_ ;
	wire _w7551_ ;
	wire _w7552_ ;
	wire _w7553_ ;
	wire _w7554_ ;
	wire _w7555_ ;
	wire _w7556_ ;
	wire _w7557_ ;
	wire _w7558_ ;
	wire _w7559_ ;
	wire _w7560_ ;
	wire _w7561_ ;
	wire _w7562_ ;
	wire _w7563_ ;
	wire _w7564_ ;
	wire _w7565_ ;
	wire _w7566_ ;
	wire _w7567_ ;
	wire _w7568_ ;
	wire _w7569_ ;
	wire _w7570_ ;
	wire _w7571_ ;
	wire _w7572_ ;
	wire _w7573_ ;
	wire _w7574_ ;
	wire _w7575_ ;
	wire _w7576_ ;
	wire _w7577_ ;
	wire _w7578_ ;
	wire _w7579_ ;
	wire _w7580_ ;
	wire _w7581_ ;
	wire _w7582_ ;
	wire _w7583_ ;
	wire _w7584_ ;
	wire _w7585_ ;
	wire _w7586_ ;
	wire _w7587_ ;
	wire _w7588_ ;
	wire _w7589_ ;
	wire _w7590_ ;
	wire _w7591_ ;
	wire _w7592_ ;
	wire _w7593_ ;
	wire _w7594_ ;
	wire _w7595_ ;
	wire _w7596_ ;
	wire _w7597_ ;
	wire _w7598_ ;
	wire _w7599_ ;
	wire _w7600_ ;
	wire _w7601_ ;
	wire _w7602_ ;
	wire _w7603_ ;
	wire _w7604_ ;
	wire _w7605_ ;
	wire _w7606_ ;
	wire _w7607_ ;
	wire _w7608_ ;
	wire _w7609_ ;
	wire _w7610_ ;
	wire _w7611_ ;
	wire _w7612_ ;
	wire _w7613_ ;
	wire _w7614_ ;
	wire _w7615_ ;
	wire _w7616_ ;
	wire _w7617_ ;
	wire _w7618_ ;
	wire _w7619_ ;
	wire _w7620_ ;
	wire _w7621_ ;
	wire _w7622_ ;
	wire _w7623_ ;
	wire _w7624_ ;
	wire _w7625_ ;
	wire _w7626_ ;
	wire _w7627_ ;
	wire _w7628_ ;
	wire _w7629_ ;
	wire _w7630_ ;
	wire _w7631_ ;
	wire _w7632_ ;
	wire _w7633_ ;
	wire _w7634_ ;
	wire _w7635_ ;
	wire _w7636_ ;
	wire _w7637_ ;
	wire _w7638_ ;
	wire _w7639_ ;
	wire _w7640_ ;
	wire _w7641_ ;
	wire _w7642_ ;
	wire _w7643_ ;
	wire _w7644_ ;
	wire _w7645_ ;
	wire _w7646_ ;
	wire _w7647_ ;
	wire _w7648_ ;
	wire _w7649_ ;
	wire _w7650_ ;
	wire _w7651_ ;
	wire _w7652_ ;
	wire _w7653_ ;
	wire _w7654_ ;
	wire _w7655_ ;
	wire _w7656_ ;
	wire _w7657_ ;
	wire _w7658_ ;
	wire _w7659_ ;
	wire _w7660_ ;
	wire _w7661_ ;
	wire _w7662_ ;
	wire _w7663_ ;
	wire _w7664_ ;
	wire _w7665_ ;
	wire _w7666_ ;
	wire _w7667_ ;
	wire _w7668_ ;
	wire _w7669_ ;
	wire _w7670_ ;
	wire _w7671_ ;
	wire _w7672_ ;
	wire _w7673_ ;
	wire _w7674_ ;
	wire _w7675_ ;
	wire _w7676_ ;
	wire _w7677_ ;
	wire _w7678_ ;
	wire _w7679_ ;
	wire _w7680_ ;
	wire _w7681_ ;
	wire _w7682_ ;
	wire _w7683_ ;
	wire _w7684_ ;
	wire _w7685_ ;
	wire _w7686_ ;
	wire _w7687_ ;
	wire _w7688_ ;
	wire _w7689_ ;
	wire _w7690_ ;
	wire _w7691_ ;
	wire _w7692_ ;
	wire _w7693_ ;
	wire _w7694_ ;
	wire _w7695_ ;
	wire _w7696_ ;
	wire _w7697_ ;
	wire _w7698_ ;
	wire _w7699_ ;
	wire _w7700_ ;
	wire _w7701_ ;
	wire _w7702_ ;
	wire _w7703_ ;
	wire _w7704_ ;
	wire _w7705_ ;
	wire _w7706_ ;
	wire _w7707_ ;
	wire _w7708_ ;
	wire _w7709_ ;
	wire _w7710_ ;
	wire _w7711_ ;
	wire _w7712_ ;
	wire _w7713_ ;
	wire _w7714_ ;
	wire _w7715_ ;
	wire _w7716_ ;
	wire _w7717_ ;
	wire _w7718_ ;
	wire _w7719_ ;
	wire _w7720_ ;
	wire _w7721_ ;
	wire _w7722_ ;
	wire _w7723_ ;
	wire _w7724_ ;
	wire _w7725_ ;
	wire _w7726_ ;
	wire _w7727_ ;
	wire _w7728_ ;
	wire _w7729_ ;
	wire _w7730_ ;
	wire _w7731_ ;
	wire _w7732_ ;
	wire _w7733_ ;
	wire _w7734_ ;
	wire _w7735_ ;
	wire _w7736_ ;
	wire _w7737_ ;
	wire _w7738_ ;
	wire _w7739_ ;
	wire _w7740_ ;
	wire _w7741_ ;
	wire _w7742_ ;
	wire _w7743_ ;
	wire _w7744_ ;
	wire _w7745_ ;
	wire _w7746_ ;
	wire _w7747_ ;
	wire _w7748_ ;
	wire _w7749_ ;
	wire _w7750_ ;
	wire _w7751_ ;
	wire _w7752_ ;
	wire _w7753_ ;
	wire _w7754_ ;
	wire _w7755_ ;
	wire _w7756_ ;
	wire _w7757_ ;
	wire _w7758_ ;
	wire _w7759_ ;
	wire _w7760_ ;
	wire _w7761_ ;
	wire _w7762_ ;
	wire _w7763_ ;
	wire _w7764_ ;
	wire _w7765_ ;
	wire _w7766_ ;
	wire _w7767_ ;
	wire _w7768_ ;
	wire _w7769_ ;
	wire _w7770_ ;
	wire _w7771_ ;
	wire _w7772_ ;
	wire _w7773_ ;
	wire _w7774_ ;
	wire _w7775_ ;
	wire _w7776_ ;
	wire _w7777_ ;
	wire _w7778_ ;
	wire _w7779_ ;
	wire _w7780_ ;
	wire _w7781_ ;
	wire _w7782_ ;
	wire _w7783_ ;
	wire _w7784_ ;
	wire _w7785_ ;
	wire _w7786_ ;
	wire _w7787_ ;
	wire _w7788_ ;
	wire _w7789_ ;
	wire _w7790_ ;
	wire _w7791_ ;
	wire _w7792_ ;
	wire _w7793_ ;
	wire _w7794_ ;
	wire _w7795_ ;
	wire _w7796_ ;
	wire _w7797_ ;
	wire _w7798_ ;
	wire _w7799_ ;
	wire _w7800_ ;
	wire _w7801_ ;
	wire _w7802_ ;
	wire _w7803_ ;
	wire _w7804_ ;
	wire _w7805_ ;
	wire _w7806_ ;
	wire _w7807_ ;
	wire _w7808_ ;
	wire _w7809_ ;
	wire _w7810_ ;
	wire _w7811_ ;
	wire _w7812_ ;
	wire _w7813_ ;
	wire _w7814_ ;
	wire _w7815_ ;
	wire _w7816_ ;
	wire _w7817_ ;
	wire _w7818_ ;
	wire _w7819_ ;
	wire _w7820_ ;
	wire _w7821_ ;
	wire _w7822_ ;
	wire _w7823_ ;
	wire _w7824_ ;
	wire _w7825_ ;
	wire _w7826_ ;
	wire _w7827_ ;
	wire _w7828_ ;
	wire _w7829_ ;
	wire _w7830_ ;
	wire _w7831_ ;
	wire _w7832_ ;
	wire _w7833_ ;
	wire _w7834_ ;
	wire _w7835_ ;
	wire _w7836_ ;
	wire _w7837_ ;
	wire _w7838_ ;
	wire _w7839_ ;
	wire _w7840_ ;
	wire _w7841_ ;
	wire _w7842_ ;
	wire _w7843_ ;
	wire _w7844_ ;
	wire _w7845_ ;
	wire _w7846_ ;
	wire _w7847_ ;
	wire _w7848_ ;
	wire _w7849_ ;
	wire _w7850_ ;
	wire _w7851_ ;
	wire _w7852_ ;
	wire _w7853_ ;
	wire _w7854_ ;
	wire _w7855_ ;
	wire _w7856_ ;
	wire _w7857_ ;
	wire _w7858_ ;
	wire _w7859_ ;
	wire _w7860_ ;
	wire _w7861_ ;
	wire _w7862_ ;
	wire _w7863_ ;
	wire _w7864_ ;
	wire _w7865_ ;
	wire _w7866_ ;
	wire _w7867_ ;
	wire _w7868_ ;
	wire _w7869_ ;
	wire _w7870_ ;
	wire _w7871_ ;
	wire _w7872_ ;
	wire _w7873_ ;
	wire _w7874_ ;
	wire _w7875_ ;
	wire _w7876_ ;
	wire _w7877_ ;
	wire _w7878_ ;
	wire _w7879_ ;
	wire _w7880_ ;
	wire _w7881_ ;
	wire _w7882_ ;
	wire _w7883_ ;
	wire _w7884_ ;
	wire _w7885_ ;
	wire _w7886_ ;
	wire _w7887_ ;
	wire _w7888_ ;
	wire _w7889_ ;
	wire _w7890_ ;
	wire _w7891_ ;
	wire _w7892_ ;
	wire _w7893_ ;
	wire _w7894_ ;
	wire _w7895_ ;
	wire _w7896_ ;
	wire _w7897_ ;
	wire _w7898_ ;
	wire _w7899_ ;
	wire _w7900_ ;
	wire _w7901_ ;
	wire _w7902_ ;
	wire _w7903_ ;
	wire _w7904_ ;
	wire _w7905_ ;
	wire _w7906_ ;
	wire _w7907_ ;
	wire _w7908_ ;
	wire _w7909_ ;
	wire _w7910_ ;
	wire _w7911_ ;
	wire _w7912_ ;
	wire _w7913_ ;
	wire _w7914_ ;
	wire _w7915_ ;
	wire _w7916_ ;
	wire _w7917_ ;
	wire _w7918_ ;
	wire _w7919_ ;
	wire _w7920_ ;
	wire _w7921_ ;
	wire _w7922_ ;
	wire _w7923_ ;
	wire _w7924_ ;
	wire _w7925_ ;
	wire _w7926_ ;
	wire _w7927_ ;
	wire _w7928_ ;
	wire _w7929_ ;
	wire _w7930_ ;
	wire _w7931_ ;
	wire _w7932_ ;
	wire _w7933_ ;
	wire _w7934_ ;
	wire _w7935_ ;
	wire _w7936_ ;
	wire _w7937_ ;
	wire _w7938_ ;
	wire _w7939_ ;
	wire _w7940_ ;
	wire _w7941_ ;
	wire _w7942_ ;
	wire _w7943_ ;
	wire _w7944_ ;
	wire _w7945_ ;
	wire _w7946_ ;
	wire _w7947_ ;
	wire _w7948_ ;
	wire _w7949_ ;
	wire _w7950_ ;
	wire _w7951_ ;
	wire _w7952_ ;
	wire _w7953_ ;
	wire _w7954_ ;
	wire _w7955_ ;
	wire _w7956_ ;
	wire _w7957_ ;
	wire _w7958_ ;
	wire _w7959_ ;
	wire _w7960_ ;
	wire _w7961_ ;
	wire _w7962_ ;
	wire _w7963_ ;
	wire _w7964_ ;
	wire _w7965_ ;
	wire _w7966_ ;
	wire _w7967_ ;
	wire _w7968_ ;
	wire _w7969_ ;
	wire _w7970_ ;
	wire _w7971_ ;
	wire _w7972_ ;
	wire _w7973_ ;
	wire _w7974_ ;
	wire _w7975_ ;
	wire _w7976_ ;
	wire _w7977_ ;
	wire _w7978_ ;
	wire _w7979_ ;
	wire _w7980_ ;
	wire _w7981_ ;
	wire _w7982_ ;
	wire _w7983_ ;
	wire _w7984_ ;
	wire _w7985_ ;
	wire _w7986_ ;
	wire _w7987_ ;
	wire _w7988_ ;
	wire _w7989_ ;
	wire _w7990_ ;
	wire _w7991_ ;
	wire _w7992_ ;
	wire _w7993_ ;
	wire _w7994_ ;
	wire _w7995_ ;
	wire _w7996_ ;
	wire _w7997_ ;
	wire _w7998_ ;
	wire _w7999_ ;
	wire _w8000_ ;
	wire _w8001_ ;
	wire _w8002_ ;
	wire _w8003_ ;
	wire _w8004_ ;
	wire _w8005_ ;
	wire _w8006_ ;
	wire _w8007_ ;
	wire _w8008_ ;
	wire _w8009_ ;
	wire _w8010_ ;
	wire _w8011_ ;
	wire _w8012_ ;
	wire _w8013_ ;
	wire _w8014_ ;
	wire _w8015_ ;
	wire _w8016_ ;
	wire _w8017_ ;
	wire _w8018_ ;
	wire _w8019_ ;
	wire _w8020_ ;
	wire _w8021_ ;
	wire _w8022_ ;
	wire _w8023_ ;
	wire _w8024_ ;
	wire _w8025_ ;
	wire _w8026_ ;
	wire _w8027_ ;
	wire _w8028_ ;
	wire _w8029_ ;
	wire _w8030_ ;
	wire _w8031_ ;
	wire _w8032_ ;
	wire _w8033_ ;
	wire _w8034_ ;
	wire _w8035_ ;
	wire _w8036_ ;
	wire _w8037_ ;
	wire _w8038_ ;
	wire _w8039_ ;
	wire _w8040_ ;
	wire _w8041_ ;
	wire _w8042_ ;
	wire _w8043_ ;
	wire _w8044_ ;
	wire _w8045_ ;
	wire _w8046_ ;
	wire _w8047_ ;
	wire _w8048_ ;
	wire _w8049_ ;
	wire _w8050_ ;
	wire _w8051_ ;
	wire _w8052_ ;
	wire _w8053_ ;
	wire _w8054_ ;
	wire _w8055_ ;
	wire _w8056_ ;
	wire _w8057_ ;
	wire _w8058_ ;
	wire _w8059_ ;
	wire _w8060_ ;
	wire _w8061_ ;
	wire _w8062_ ;
	wire _w8063_ ;
	wire _w8064_ ;
	wire _w8065_ ;
	wire _w8066_ ;
	wire _w8067_ ;
	wire _w8068_ ;
	wire _w8069_ ;
	wire _w8070_ ;
	wire _w8071_ ;
	wire _w8072_ ;
	wire _w8073_ ;
	wire _w8074_ ;
	wire _w8075_ ;
	wire _w8076_ ;
	wire _w8077_ ;
	wire _w8078_ ;
	wire _w8079_ ;
	wire _w8080_ ;
	wire _w8081_ ;
	wire _w8082_ ;
	wire _w8083_ ;
	wire _w8084_ ;
	wire _w8085_ ;
	wire _w8086_ ;
	wire _w8087_ ;
	wire _w8088_ ;
	wire _w8089_ ;
	wire _w8090_ ;
	wire _w8091_ ;
	wire _w8092_ ;
	wire _w8093_ ;
	wire _w8094_ ;
	wire _w8095_ ;
	wire _w8096_ ;
	wire _w8097_ ;
	wire _w8098_ ;
	wire _w8099_ ;
	wire _w8100_ ;
	wire _w8101_ ;
	wire _w8102_ ;
	wire _w8103_ ;
	wire _w8104_ ;
	wire _w8105_ ;
	wire _w8106_ ;
	wire _w8107_ ;
	wire _w8108_ ;
	wire _w8109_ ;
	wire _w8110_ ;
	wire _w8111_ ;
	wire _w8112_ ;
	wire _w8113_ ;
	wire _w8114_ ;
	wire _w8115_ ;
	wire _w8116_ ;
	wire _w8117_ ;
	wire _w8118_ ;
	wire _w8119_ ;
	wire _w8120_ ;
	wire _w8121_ ;
	wire _w8122_ ;
	wire _w8123_ ;
	wire _w8124_ ;
	wire _w8125_ ;
	wire _w8126_ ;
	wire _w8127_ ;
	wire _w8128_ ;
	wire _w8129_ ;
	wire _w8130_ ;
	wire _w8131_ ;
	wire _w8132_ ;
	wire _w8133_ ;
	wire _w8134_ ;
	wire _w8135_ ;
	wire _w8136_ ;
	wire _w8137_ ;
	wire _w8138_ ;
	wire _w8139_ ;
	wire _w8140_ ;
	wire _w8141_ ;
	wire _w8142_ ;
	wire _w8143_ ;
	wire _w8144_ ;
	wire _w8145_ ;
	wire _w8146_ ;
	wire _w8147_ ;
	wire _w8148_ ;
	wire _w8149_ ;
	wire _w8150_ ;
	wire _w8151_ ;
	wire _w8152_ ;
	wire _w8153_ ;
	wire _w8154_ ;
	wire _w8155_ ;
	wire _w8156_ ;
	wire _w8157_ ;
	wire _w8158_ ;
	wire _w8159_ ;
	wire _w8160_ ;
	wire _w8161_ ;
	wire _w8162_ ;
	wire _w8163_ ;
	wire _w8164_ ;
	wire _w8165_ ;
	wire _w8166_ ;
	wire _w8167_ ;
	wire _w8168_ ;
	wire _w8169_ ;
	wire _w8170_ ;
	wire _w8171_ ;
	wire _w8172_ ;
	wire _w8173_ ;
	wire _w8174_ ;
	wire _w8175_ ;
	wire _w8176_ ;
	wire _w8177_ ;
	wire _w8178_ ;
	wire _w8179_ ;
	wire _w8180_ ;
	wire _w8181_ ;
	wire _w8182_ ;
	wire _w8183_ ;
	wire _w8184_ ;
	wire _w8185_ ;
	wire _w8186_ ;
	wire _w8187_ ;
	wire _w8188_ ;
	wire _w8189_ ;
	wire _w8190_ ;
	wire _w8191_ ;
	wire _w8192_ ;
	wire _w8193_ ;
	wire _w8194_ ;
	wire _w8195_ ;
	wire _w8196_ ;
	wire _w8197_ ;
	wire _w8198_ ;
	wire _w8199_ ;
	wire _w8200_ ;
	wire _w8201_ ;
	wire _w8202_ ;
	wire _w8203_ ;
	wire _w8204_ ;
	wire _w8205_ ;
	wire _w8206_ ;
	wire _w8207_ ;
	wire _w8208_ ;
	wire _w8209_ ;
	wire _w8210_ ;
	wire _w8211_ ;
	wire _w8212_ ;
	wire _w8213_ ;
	wire _w8214_ ;
	wire _w8215_ ;
	wire _w8216_ ;
	wire _w8217_ ;
	wire _w8218_ ;
	wire _w8219_ ;
	wire _w8220_ ;
	wire _w8221_ ;
	wire _w8222_ ;
	wire _w8223_ ;
	wire _w8224_ ;
	wire _w8225_ ;
	wire _w8226_ ;
	wire _w8227_ ;
	wire _w8228_ ;
	wire _w8229_ ;
	wire _w8230_ ;
	wire _w8231_ ;
	wire _w8232_ ;
	wire _w8233_ ;
	wire _w8234_ ;
	wire _w8235_ ;
	wire _w8236_ ;
	wire _w8237_ ;
	wire _w8238_ ;
	wire _w8239_ ;
	wire _w8240_ ;
	wire _w8241_ ;
	wire _w8242_ ;
	wire _w8243_ ;
	wire _w8244_ ;
	wire _w8245_ ;
	wire _w8246_ ;
	wire _w8247_ ;
	wire _w8248_ ;
	wire _w8249_ ;
	wire _w8250_ ;
	wire _w8251_ ;
	wire _w8252_ ;
	wire _w8253_ ;
	wire _w8254_ ;
	wire _w8255_ ;
	wire _w8256_ ;
	wire _w8257_ ;
	wire _w8258_ ;
	wire _w8259_ ;
	wire _w8260_ ;
	wire _w8261_ ;
	wire _w8262_ ;
	wire _w8263_ ;
	wire _w8264_ ;
	wire _w8265_ ;
	wire _w8266_ ;
	wire _w8267_ ;
	wire _w8268_ ;
	wire _w8269_ ;
	wire _w8270_ ;
	wire _w8271_ ;
	wire _w8272_ ;
	wire _w8273_ ;
	wire _w8274_ ;
	wire _w8275_ ;
	wire _w8276_ ;
	wire _w8277_ ;
	wire _w8278_ ;
	wire _w8279_ ;
	wire _w8280_ ;
	wire _w8281_ ;
	wire _w8282_ ;
	wire _w8283_ ;
	wire _w8284_ ;
	wire _w8285_ ;
	wire _w8286_ ;
	wire _w8287_ ;
	wire _w8288_ ;
	wire _w8289_ ;
	wire _w8290_ ;
	wire _w8291_ ;
	wire _w8292_ ;
	wire _w8293_ ;
	wire _w8294_ ;
	wire _w8295_ ;
	wire _w8296_ ;
	wire _w8297_ ;
	wire _w8298_ ;
	wire _w8299_ ;
	wire _w8300_ ;
	wire _w8301_ ;
	wire _w8302_ ;
	wire _w8303_ ;
	wire _w8304_ ;
	wire _w8305_ ;
	wire _w8306_ ;
	wire _w8307_ ;
	wire _w8308_ ;
	wire _w8309_ ;
	wire _w8310_ ;
	wire _w8311_ ;
	wire _w8312_ ;
	wire _w8313_ ;
	wire _w8314_ ;
	wire _w8315_ ;
	wire _w8316_ ;
	wire _w8317_ ;
	wire _w8318_ ;
	wire _w8319_ ;
	wire _w8320_ ;
	wire _w8321_ ;
	wire _w8322_ ;
	wire _w8323_ ;
	wire _w8324_ ;
	wire _w8325_ ;
	wire _w8326_ ;
	wire _w8327_ ;
	wire _w8328_ ;
	wire _w8329_ ;
	wire _w8330_ ;
	wire _w8331_ ;
	wire _w8332_ ;
	wire _w8333_ ;
	wire _w8334_ ;
	wire _w8335_ ;
	wire _w8336_ ;
	wire _w8337_ ;
	wire _w8338_ ;
	wire _w8339_ ;
	wire _w8340_ ;
	wire _w8341_ ;
	wire _w8342_ ;
	wire _w8343_ ;
	wire _w8344_ ;
	wire _w8345_ ;
	wire _w8346_ ;
	wire _w8347_ ;
	wire _w8348_ ;
	wire _w8349_ ;
	wire _w8350_ ;
	wire _w8351_ ;
	wire _w8352_ ;
	wire _w8353_ ;
	wire _w8354_ ;
	wire _w8355_ ;
	wire _w8356_ ;
	wire _w8357_ ;
	wire _w8358_ ;
	wire _w8359_ ;
	wire _w8360_ ;
	wire _w8361_ ;
	wire _w8362_ ;
	wire _w8363_ ;
	wire _w8364_ ;
	wire _w8365_ ;
	wire _w8366_ ;
	wire _w8367_ ;
	wire _w8368_ ;
	wire _w8369_ ;
	wire _w8370_ ;
	wire _w8371_ ;
	wire _w8372_ ;
	wire _w8373_ ;
	wire _w8374_ ;
	wire _w8375_ ;
	wire _w8376_ ;
	wire _w8377_ ;
	wire _w8378_ ;
	wire _w8379_ ;
	wire _w8380_ ;
	wire _w8381_ ;
	wire _w8382_ ;
	wire _w8383_ ;
	wire _w8384_ ;
	wire _w8385_ ;
	wire _w8386_ ;
	wire _w8387_ ;
	wire _w8388_ ;
	wire _w8389_ ;
	wire _w8390_ ;
	wire _w8391_ ;
	wire _w8392_ ;
	wire _w8393_ ;
	wire _w8394_ ;
	wire _w8395_ ;
	wire _w8396_ ;
	wire _w8397_ ;
	wire _w8398_ ;
	wire _w8399_ ;
	wire _w8400_ ;
	wire _w8401_ ;
	wire _w8402_ ;
	wire _w8403_ ;
	wire _w8404_ ;
	wire _w8405_ ;
	wire _w8406_ ;
	wire _w8407_ ;
	wire _w8408_ ;
	wire _w8409_ ;
	wire _w8410_ ;
	wire _w8411_ ;
	wire _w8412_ ;
	wire _w8413_ ;
	wire _w8414_ ;
	wire _w8415_ ;
	wire _w8416_ ;
	wire _w8417_ ;
	wire _w8418_ ;
	wire _w8419_ ;
	wire _w8420_ ;
	wire _w8421_ ;
	wire _w8422_ ;
	wire _w8423_ ;
	wire _w8424_ ;
	wire _w8425_ ;
	wire _w8426_ ;
	wire _w8427_ ;
	wire _w8428_ ;
	wire _w8429_ ;
	wire _w8430_ ;
	wire _w8431_ ;
	wire _w8432_ ;
	wire _w8433_ ;
	wire _w8434_ ;
	wire _w8435_ ;
	wire _w8436_ ;
	wire _w8437_ ;
	wire _w8438_ ;
	wire _w8439_ ;
	wire _w8440_ ;
	wire _w8441_ ;
	wire _w8442_ ;
	wire _w8443_ ;
	wire _w8444_ ;
	wire _w8445_ ;
	wire _w8446_ ;
	wire _w8447_ ;
	wire _w8448_ ;
	wire _w8449_ ;
	wire _w8450_ ;
	wire _w8451_ ;
	wire _w8452_ ;
	wire _w8453_ ;
	wire _w8454_ ;
	wire _w8455_ ;
	wire _w8456_ ;
	wire _w8457_ ;
	wire _w8458_ ;
	wire _w8459_ ;
	wire _w8460_ ;
	wire _w8461_ ;
	wire _w8462_ ;
	wire _w8463_ ;
	wire _w8464_ ;
	wire _w8465_ ;
	wire _w8466_ ;
	wire _w8467_ ;
	wire _w8468_ ;
	wire _w8469_ ;
	wire _w8470_ ;
	wire _w8471_ ;
	wire _w8472_ ;
	wire _w8473_ ;
	wire _w8474_ ;
	wire _w8475_ ;
	wire _w8476_ ;
	wire _w8477_ ;
	wire _w8478_ ;
	wire _w8479_ ;
	wire _w8480_ ;
	wire _w8481_ ;
	wire _w8482_ ;
	wire _w8483_ ;
	wire _w8484_ ;
	wire _w8485_ ;
	wire _w8486_ ;
	wire _w8487_ ;
	wire _w8488_ ;
	wire _w8489_ ;
	wire _w8490_ ;
	wire _w8491_ ;
	wire _w8492_ ;
	wire _w8493_ ;
	wire _w8494_ ;
	wire _w8495_ ;
	wire _w8496_ ;
	wire _w8497_ ;
	wire _w8498_ ;
	wire _w8499_ ;
	wire _w8500_ ;
	wire _w8501_ ;
	wire _w8502_ ;
	wire _w8503_ ;
	wire _w8504_ ;
	wire _w8505_ ;
	wire _w8506_ ;
	wire _w8507_ ;
	wire _w8508_ ;
	wire _w8509_ ;
	wire _w8510_ ;
	wire _w8511_ ;
	wire _w8512_ ;
	wire _w8513_ ;
	wire _w8514_ ;
	wire _w8515_ ;
	wire _w8516_ ;
	wire _w8517_ ;
	wire _w8518_ ;
	wire _w8519_ ;
	wire _w8520_ ;
	wire _w8521_ ;
	wire _w8522_ ;
	wire _w8523_ ;
	wire _w8524_ ;
	wire _w8525_ ;
	wire _w8526_ ;
	wire _w8527_ ;
	wire _w8528_ ;
	wire _w8529_ ;
	wire _w8530_ ;
	wire _w8531_ ;
	wire _w8532_ ;
	wire _w8533_ ;
	wire _w8534_ ;
	wire _w8535_ ;
	wire _w8536_ ;
	wire _w8537_ ;
	wire _w8538_ ;
	wire _w8539_ ;
	wire _w8540_ ;
	wire _w8541_ ;
	wire _w8542_ ;
	wire _w8543_ ;
	wire _w8544_ ;
	wire _w8545_ ;
	wire _w8546_ ;
	wire _w8547_ ;
	wire _w8548_ ;
	wire _w8549_ ;
	wire _w8550_ ;
	wire _w8551_ ;
	wire _w8552_ ;
	wire _w8553_ ;
	wire _w8554_ ;
	wire _w8555_ ;
	wire _w8556_ ;
	wire _w8557_ ;
	wire _w8558_ ;
	wire _w8559_ ;
	wire _w8560_ ;
	wire _w8561_ ;
	wire _w8562_ ;
	wire _w8563_ ;
	wire _w8564_ ;
	wire _w8565_ ;
	wire _w8566_ ;
	wire _w8567_ ;
	wire _w8568_ ;
	wire _w8569_ ;
	wire _w8570_ ;
	wire _w8571_ ;
	wire _w8572_ ;
	wire _w8573_ ;
	wire _w8574_ ;
	wire _w8575_ ;
	wire _w8576_ ;
	wire _w8577_ ;
	wire _w8578_ ;
	wire _w8579_ ;
	wire _w8580_ ;
	wire _w8581_ ;
	wire _w8582_ ;
	wire _w8583_ ;
	wire _w8584_ ;
	wire _w8585_ ;
	wire _w8586_ ;
	wire _w8587_ ;
	wire _w8588_ ;
	wire _w8589_ ;
	wire _w8590_ ;
	wire _w8591_ ;
	wire _w8592_ ;
	wire _w8593_ ;
	wire _w8594_ ;
	wire _w8595_ ;
	wire _w8596_ ;
	wire _w8597_ ;
	wire _w8598_ ;
	wire _w8599_ ;
	wire _w8600_ ;
	wire _w8601_ ;
	wire _w8602_ ;
	wire _w8603_ ;
	wire _w8604_ ;
	wire _w8605_ ;
	wire _w8606_ ;
	wire _w8607_ ;
	wire _w8608_ ;
	wire _w8609_ ;
	wire _w8610_ ;
	wire _w8611_ ;
	wire _w8612_ ;
	wire _w8613_ ;
	wire _w8614_ ;
	wire _w8615_ ;
	wire _w8616_ ;
	wire _w8617_ ;
	wire _w8618_ ;
	wire _w8619_ ;
	wire _w8620_ ;
	wire _w8621_ ;
	wire _w8622_ ;
	wire _w8623_ ;
	wire _w8624_ ;
	wire _w8625_ ;
	wire _w8626_ ;
	wire _w8627_ ;
	wire _w8628_ ;
	wire _w8629_ ;
	wire _w8630_ ;
	wire _w8631_ ;
	wire _w8632_ ;
	wire _w8633_ ;
	wire _w8634_ ;
	wire _w8635_ ;
	wire _w8636_ ;
	wire _w8637_ ;
	wire _w8638_ ;
	wire _w8639_ ;
	wire _w8640_ ;
	wire _w8641_ ;
	wire _w8642_ ;
	wire _w8643_ ;
	wire _w8644_ ;
	wire _w8645_ ;
	wire _w8646_ ;
	wire _w8647_ ;
	wire _w8648_ ;
	wire _w8649_ ;
	wire _w8650_ ;
	wire _w8651_ ;
	wire _w8652_ ;
	wire _w8653_ ;
	wire _w8654_ ;
	wire _w8655_ ;
	wire _w8656_ ;
	wire _w8657_ ;
	wire _w8658_ ;
	wire _w8659_ ;
	wire _w8660_ ;
	wire _w8661_ ;
	wire _w8662_ ;
	wire _w8663_ ;
	wire _w8664_ ;
	wire _w8665_ ;
	wire _w8666_ ;
	wire _w8667_ ;
	wire _w8668_ ;
	wire _w8669_ ;
	wire _w8670_ ;
	wire _w8671_ ;
	wire _w8672_ ;
	wire _w8673_ ;
	wire _w8674_ ;
	wire _w8675_ ;
	wire _w8676_ ;
	wire _w8677_ ;
	wire _w8678_ ;
	wire _w8679_ ;
	wire _w8680_ ;
	wire _w8681_ ;
	wire _w8682_ ;
	wire _w8683_ ;
	wire _w8684_ ;
	wire _w8685_ ;
	wire _w8686_ ;
	wire _w8687_ ;
	wire _w8688_ ;
	wire _w8689_ ;
	wire _w8690_ ;
	wire _w8691_ ;
	wire _w8692_ ;
	wire _w8693_ ;
	wire _w8694_ ;
	wire _w8695_ ;
	wire _w8696_ ;
	wire _w8697_ ;
	wire _w8698_ ;
	wire _w8699_ ;
	wire _w8700_ ;
	wire _w8701_ ;
	wire _w8702_ ;
	wire _w8703_ ;
	wire _w8704_ ;
	wire _w8705_ ;
	wire _w8706_ ;
	wire _w8707_ ;
	wire _w8708_ ;
	wire _w8709_ ;
	wire _w8710_ ;
	wire _w8711_ ;
	wire _w8712_ ;
	wire _w8713_ ;
	wire _w8714_ ;
	wire _w8715_ ;
	wire _w8716_ ;
	wire _w8717_ ;
	wire _w8718_ ;
	wire _w8719_ ;
	wire _w8720_ ;
	wire _w8721_ ;
	wire _w8722_ ;
	wire _w8723_ ;
	wire _w8724_ ;
	wire _w8725_ ;
	wire _w8726_ ;
	wire _w8727_ ;
	wire _w8728_ ;
	wire _w8729_ ;
	wire _w8730_ ;
	wire _w8731_ ;
	wire _w8732_ ;
	wire _w8733_ ;
	wire _w8734_ ;
	wire _w8735_ ;
	wire _w8736_ ;
	wire _w8737_ ;
	wire _w8738_ ;
	wire _w8739_ ;
	wire _w8740_ ;
	wire _w8741_ ;
	wire _w8742_ ;
	wire _w8743_ ;
	wire _w8744_ ;
	wire _w8745_ ;
	wire _w8746_ ;
	wire _w8747_ ;
	wire _w8748_ ;
	wire _w8749_ ;
	wire _w8750_ ;
	wire _w8751_ ;
	wire _w8752_ ;
	wire _w8753_ ;
	wire _w8754_ ;
	wire _w8755_ ;
	wire _w8756_ ;
	wire _w8757_ ;
	wire _w8758_ ;
	wire _w8759_ ;
	wire _w8760_ ;
	wire _w8761_ ;
	wire _w8762_ ;
	wire _w8763_ ;
	wire _w8764_ ;
	wire _w8765_ ;
	wire _w8766_ ;
	wire _w8767_ ;
	wire _w8768_ ;
	wire _w8769_ ;
	wire _w8770_ ;
	wire _w8771_ ;
	wire _w8772_ ;
	wire _w8773_ ;
	wire _w8774_ ;
	wire _w8775_ ;
	wire _w8776_ ;
	wire _w8777_ ;
	wire _w8778_ ;
	wire _w8779_ ;
	wire _w8780_ ;
	wire _w8781_ ;
	wire _w8782_ ;
	wire _w8783_ ;
	wire _w8784_ ;
	wire _w8785_ ;
	wire _w8786_ ;
	wire _w8787_ ;
	wire _w8788_ ;
	wire _w8789_ ;
	wire _w8790_ ;
	wire _w8791_ ;
	wire _w8792_ ;
	wire _w8793_ ;
	wire _w8794_ ;
	wire _w8795_ ;
	wire _w8796_ ;
	wire _w8797_ ;
	wire _w8798_ ;
	wire _w8799_ ;
	wire _w8800_ ;
	wire _w8801_ ;
	wire _w8802_ ;
	wire _w8803_ ;
	wire _w8804_ ;
	wire _w8805_ ;
	wire _w8806_ ;
	wire _w8807_ ;
	wire _w8808_ ;
	wire _w8809_ ;
	wire _w8810_ ;
	wire _w8811_ ;
	wire _w8812_ ;
	wire _w8813_ ;
	wire _w8814_ ;
	wire _w8815_ ;
	wire _w8816_ ;
	wire _w8817_ ;
	wire _w8818_ ;
	wire _w8819_ ;
	wire _w8820_ ;
	wire _w8821_ ;
	wire _w8822_ ;
	wire _w8823_ ;
	wire _w8824_ ;
	wire _w8825_ ;
	wire _w8826_ ;
	wire _w8827_ ;
	wire _w8828_ ;
	wire _w8829_ ;
	wire _w8830_ ;
	wire _w8831_ ;
	wire _w8832_ ;
	wire _w8833_ ;
	wire _w8834_ ;
	wire _w8835_ ;
	wire _w8836_ ;
	wire _w8837_ ;
	wire _w8838_ ;
	wire _w8839_ ;
	wire _w8840_ ;
	wire _w8841_ ;
	wire _w8842_ ;
	wire _w8843_ ;
	wire _w8844_ ;
	wire _w8845_ ;
	wire _w8846_ ;
	wire _w8847_ ;
	wire _w8848_ ;
	wire _w8849_ ;
	wire _w8850_ ;
	wire _w8851_ ;
	wire _w8852_ ;
	wire _w8853_ ;
	wire _w8854_ ;
	wire _w8855_ ;
	wire _w8856_ ;
	wire _w8857_ ;
	wire _w8858_ ;
	wire _w8859_ ;
	wire _w8860_ ;
	wire _w8861_ ;
	wire _w8862_ ;
	wire _w8863_ ;
	wire _w8864_ ;
	wire _w8865_ ;
	wire _w8866_ ;
	wire _w8867_ ;
	wire _w8868_ ;
	wire _w8869_ ;
	wire _w8870_ ;
	wire _w8871_ ;
	wire _w8872_ ;
	wire _w8873_ ;
	wire _w8874_ ;
	wire _w8875_ ;
	wire _w8876_ ;
	wire _w8877_ ;
	wire _w8878_ ;
	wire _w8879_ ;
	wire _w8880_ ;
	wire _w8881_ ;
	wire _w8882_ ;
	wire _w8883_ ;
	wire _w8884_ ;
	wire _w8885_ ;
	wire _w8886_ ;
	wire _w8887_ ;
	wire _w8888_ ;
	wire _w8889_ ;
	wire _w8890_ ;
	wire _w8891_ ;
	wire _w8892_ ;
	wire _w8893_ ;
	wire _w8894_ ;
	wire _w8895_ ;
	wire _w8896_ ;
	wire _w8897_ ;
	wire _w8898_ ;
	wire _w8899_ ;
	wire _w8900_ ;
	wire _w8901_ ;
	wire _w8902_ ;
	wire _w8903_ ;
	wire _w8904_ ;
	wire _w8905_ ;
	wire _w8906_ ;
	wire _w8907_ ;
	wire _w8908_ ;
	wire _w8909_ ;
	wire _w8910_ ;
	wire _w8911_ ;
	wire _w8912_ ;
	wire _w8913_ ;
	wire _w8914_ ;
	wire _w8915_ ;
	wire _w8916_ ;
	wire _w8917_ ;
	wire _w8918_ ;
	wire _w8919_ ;
	wire _w8920_ ;
	wire _w8921_ ;
	wire _w8922_ ;
	wire _w8923_ ;
	wire _w8924_ ;
	wire _w8925_ ;
	wire _w8926_ ;
	wire _w8927_ ;
	wire _w8928_ ;
	wire _w8929_ ;
	wire _w8930_ ;
	wire _w8931_ ;
	wire _w8932_ ;
	wire _w8933_ ;
	wire _w8934_ ;
	wire _w8935_ ;
	wire _w8936_ ;
	wire _w8937_ ;
	wire _w8938_ ;
	wire _w8939_ ;
	wire _w8940_ ;
	wire _w8941_ ;
	wire _w8942_ ;
	wire _w8943_ ;
	wire _w8944_ ;
	wire _w8945_ ;
	wire _w8946_ ;
	wire _w8947_ ;
	wire _w8948_ ;
	wire _w8949_ ;
	wire _w8950_ ;
	wire _w8951_ ;
	wire _w8952_ ;
	wire _w8953_ ;
	wire _w8954_ ;
	wire _w8955_ ;
	wire _w8956_ ;
	wire _w8957_ ;
	wire _w8958_ ;
	wire _w8959_ ;
	wire _w8960_ ;
	wire _w8961_ ;
	wire _w8962_ ;
	wire _w8963_ ;
	wire _w8964_ ;
	wire _w8965_ ;
	wire _w8966_ ;
	wire _w8967_ ;
	wire _w8968_ ;
	wire _w8969_ ;
	wire _w8970_ ;
	wire _w8971_ ;
	wire _w8972_ ;
	wire _w8973_ ;
	wire _w8974_ ;
	wire _w8975_ ;
	wire _w8976_ ;
	wire _w8977_ ;
	wire _w8978_ ;
	wire _w8979_ ;
	wire _w8980_ ;
	wire _w8981_ ;
	wire _w8982_ ;
	wire _w8983_ ;
	wire _w8984_ ;
	wire _w8985_ ;
	wire _w8986_ ;
	wire _w8987_ ;
	wire _w8988_ ;
	wire _w8989_ ;
	wire _w8990_ ;
	wire _w8991_ ;
	wire _w8992_ ;
	wire _w8993_ ;
	wire _w8994_ ;
	wire _w8995_ ;
	wire _w8996_ ;
	wire _w8997_ ;
	wire _w8998_ ;
	wire _w8999_ ;
	wire _w9000_ ;
	wire _w9001_ ;
	wire _w9002_ ;
	wire _w9003_ ;
	wire _w9004_ ;
	wire _w9005_ ;
	wire _w9006_ ;
	wire _w9007_ ;
	wire _w9008_ ;
	wire _w9009_ ;
	wire _w9010_ ;
	wire _w9011_ ;
	wire _w9012_ ;
	wire _w9013_ ;
	wire _w9014_ ;
	wire _w9015_ ;
	wire _w9016_ ;
	wire _w9017_ ;
	wire _w9018_ ;
	wire _w9019_ ;
	wire _w9020_ ;
	wire _w9021_ ;
	wire _w9022_ ;
	wire _w9023_ ;
	wire _w9024_ ;
	wire _w9025_ ;
	wire _w9026_ ;
	wire _w9027_ ;
	wire _w9028_ ;
	wire _w9029_ ;
	wire _w9030_ ;
	wire _w9031_ ;
	wire _w9032_ ;
	wire _w9033_ ;
	wire _w9034_ ;
	wire _w9035_ ;
	wire _w9036_ ;
	wire _w9037_ ;
	wire _w9038_ ;
	wire _w9039_ ;
	wire _w9040_ ;
	wire _w9041_ ;
	wire _w9042_ ;
	wire _w9043_ ;
	wire _w9044_ ;
	wire _w9045_ ;
	wire _w9046_ ;
	wire _w9047_ ;
	wire _w9048_ ;
	wire _w9049_ ;
	wire _w9050_ ;
	wire _w9051_ ;
	wire _w9052_ ;
	wire _w9053_ ;
	wire _w9054_ ;
	wire _w9055_ ;
	wire _w9056_ ;
	wire _w9057_ ;
	wire _w9058_ ;
	wire _w9059_ ;
	wire _w9060_ ;
	wire _w9061_ ;
	wire _w9062_ ;
	wire _w9063_ ;
	wire _w9064_ ;
	wire _w9065_ ;
	wire _w9066_ ;
	wire _w9067_ ;
	wire _w9068_ ;
	wire _w9069_ ;
	wire _w9070_ ;
	wire _w9071_ ;
	wire _w9072_ ;
	wire _w9073_ ;
	wire _w9074_ ;
	wire _w9075_ ;
	wire _w9076_ ;
	wire _w9077_ ;
	wire _w9078_ ;
	wire _w9079_ ;
	wire _w9080_ ;
	wire _w9081_ ;
	wire _w9082_ ;
	wire _w9083_ ;
	wire _w9084_ ;
	wire _w9085_ ;
	wire _w9086_ ;
	wire _w9087_ ;
	wire _w9088_ ;
	wire _w9089_ ;
	wire _w9090_ ;
	wire _w9091_ ;
	wire _w9092_ ;
	wire _w9093_ ;
	wire _w9094_ ;
	wire _w9095_ ;
	wire _w9096_ ;
	wire _w9097_ ;
	wire _w9098_ ;
	wire _w9099_ ;
	wire _w9100_ ;
	wire _w9101_ ;
	wire _w9102_ ;
	wire _w9103_ ;
	wire _w9104_ ;
	wire _w9105_ ;
	wire _w9106_ ;
	wire _w9107_ ;
	wire _w9108_ ;
	wire _w9109_ ;
	wire _w9110_ ;
	wire _w9111_ ;
	wire _w9112_ ;
	wire _w9113_ ;
	wire _w9114_ ;
	wire _w9115_ ;
	wire _w9116_ ;
	wire _w9117_ ;
	wire _w9118_ ;
	wire _w9119_ ;
	wire _w9120_ ;
	wire _w9121_ ;
	wire _w9122_ ;
	wire _w9123_ ;
	wire _w9124_ ;
	wire _w9125_ ;
	wire _w9126_ ;
	wire _w9127_ ;
	wire _w9128_ ;
	wire _w9129_ ;
	wire _w9130_ ;
	wire _w9131_ ;
	wire _w9132_ ;
	wire _w9133_ ;
	wire _w9134_ ;
	wire _w9135_ ;
	wire _w9136_ ;
	wire _w9137_ ;
	wire _w9138_ ;
	wire _w9139_ ;
	wire _w9140_ ;
	wire _w9141_ ;
	wire _w9142_ ;
	wire _w9143_ ;
	wire _w9144_ ;
	wire _w9145_ ;
	wire _w9146_ ;
	wire _w9147_ ;
	wire _w9148_ ;
	wire _w9149_ ;
	wire _w9150_ ;
	wire _w9151_ ;
	wire _w9152_ ;
	wire _w9153_ ;
	wire _w9154_ ;
	wire _w9155_ ;
	wire _w9156_ ;
	wire _w9157_ ;
	wire _w9158_ ;
	wire _w9159_ ;
	wire _w9160_ ;
	wire _w9161_ ;
	wire _w9162_ ;
	wire _w9163_ ;
	wire _w9164_ ;
	wire _w9165_ ;
	wire _w9166_ ;
	wire _w9167_ ;
	wire _w9168_ ;
	wire _w9169_ ;
	wire _w9170_ ;
	wire _w9171_ ;
	wire _w9172_ ;
	wire _w9173_ ;
	wire _w9174_ ;
	wire _w9175_ ;
	wire _w9176_ ;
	wire _w9177_ ;
	wire _w9178_ ;
	wire _w9179_ ;
	wire _w9180_ ;
	wire _w9181_ ;
	wire _w9182_ ;
	wire _w9183_ ;
	wire _w9184_ ;
	wire _w9185_ ;
	wire _w9186_ ;
	wire _w9187_ ;
	wire _w9188_ ;
	wire _w9189_ ;
	wire _w9190_ ;
	wire _w9191_ ;
	wire _w9192_ ;
	wire _w9193_ ;
	wire _w9194_ ;
	wire _w9195_ ;
	wire _w9196_ ;
	wire _w9197_ ;
	wire _w9198_ ;
	wire _w9199_ ;
	wire _w9200_ ;
	wire _w9201_ ;
	wire _w9202_ ;
	wire _w9203_ ;
	wire _w9204_ ;
	wire _w9205_ ;
	wire _w9206_ ;
	wire _w9207_ ;
	wire _w9208_ ;
	wire _w9209_ ;
	wire _w9210_ ;
	wire _w9211_ ;
	wire _w9212_ ;
	wire _w9213_ ;
	wire _w9214_ ;
	wire _w9215_ ;
	wire _w9216_ ;
	wire _w9217_ ;
	wire _w9218_ ;
	wire _w9219_ ;
	wire _w9220_ ;
	wire _w9221_ ;
	wire _w9222_ ;
	wire _w9223_ ;
	wire _w9224_ ;
	wire _w9225_ ;
	wire _w9226_ ;
	wire _w9227_ ;
	wire _w9228_ ;
	wire _w9229_ ;
	wire _w9230_ ;
	wire _w9231_ ;
	wire _w9232_ ;
	wire _w9233_ ;
	wire _w9234_ ;
	wire _w9235_ ;
	wire _w9236_ ;
	wire _w9237_ ;
	wire _w9238_ ;
	wire _w9239_ ;
	wire _w9240_ ;
	wire _w9241_ ;
	wire _w9242_ ;
	wire _w9243_ ;
	wire _w9244_ ;
	wire _w9245_ ;
	wire _w9246_ ;
	wire _w9247_ ;
	wire _w9248_ ;
	wire _w9249_ ;
	wire _w9250_ ;
	wire _w9251_ ;
	wire _w9252_ ;
	wire _w9253_ ;
	wire _w9254_ ;
	wire _w9255_ ;
	wire _w9256_ ;
	wire _w9257_ ;
	wire _w9258_ ;
	wire _w9259_ ;
	wire _w9260_ ;
	wire _w9261_ ;
	wire _w9262_ ;
	wire _w9263_ ;
	wire _w9264_ ;
	wire _w9265_ ;
	wire _w9266_ ;
	wire _w9267_ ;
	wire _w9268_ ;
	wire _w9269_ ;
	wire _w9270_ ;
	wire _w9271_ ;
	wire _w9272_ ;
	wire _w9273_ ;
	wire _w9274_ ;
	wire _w9275_ ;
	wire _w9276_ ;
	wire _w9277_ ;
	wire _w9278_ ;
	wire _w9279_ ;
	wire _w9280_ ;
	wire _w9281_ ;
	wire _w9282_ ;
	wire _w9283_ ;
	wire _w9284_ ;
	wire _w9285_ ;
	wire _w9286_ ;
	wire _w9287_ ;
	wire _w9288_ ;
	wire _w9289_ ;
	wire _w9290_ ;
	wire _w9291_ ;
	wire _w9292_ ;
	wire _w9293_ ;
	wire _w9294_ ;
	wire _w9295_ ;
	wire _w9296_ ;
	wire _w9297_ ;
	wire _w9298_ ;
	wire _w9299_ ;
	wire _w9300_ ;
	wire _w9301_ ;
	wire _w9302_ ;
	wire _w9303_ ;
	wire _w9304_ ;
	wire _w9305_ ;
	wire _w9306_ ;
	wire _w9307_ ;
	wire _w9308_ ;
	wire _w9309_ ;
	wire _w9310_ ;
	wire _w9311_ ;
	wire _w9312_ ;
	wire _w9313_ ;
	wire _w9314_ ;
	wire _w9315_ ;
	wire _w9316_ ;
	wire _w9317_ ;
	wire _w9318_ ;
	wire _w9319_ ;
	wire _w9320_ ;
	wire _w9321_ ;
	wire _w9322_ ;
	wire _w9323_ ;
	wire _w9324_ ;
	wire _w9325_ ;
	wire _w9326_ ;
	wire _w9327_ ;
	wire _w9328_ ;
	wire _w9329_ ;
	wire _w9330_ ;
	wire _w9331_ ;
	wire _w9332_ ;
	wire _w9333_ ;
	wire _w9334_ ;
	wire _w9335_ ;
	wire _w9336_ ;
	wire _w9337_ ;
	wire _w9338_ ;
	wire _w9339_ ;
	wire _w9340_ ;
	wire _w9341_ ;
	wire _w9342_ ;
	wire _w9343_ ;
	wire _w9344_ ;
	wire _w9345_ ;
	wire _w9346_ ;
	wire _w9347_ ;
	wire _w9348_ ;
	wire _w9349_ ;
	wire _w9350_ ;
	wire _w9351_ ;
	wire _w9352_ ;
	wire _w9353_ ;
	wire _w9354_ ;
	wire _w9355_ ;
	wire _w9356_ ;
	wire _w9357_ ;
	wire _w9358_ ;
	wire _w9359_ ;
	wire _w9360_ ;
	wire _w9361_ ;
	wire _w9362_ ;
	wire _w9363_ ;
	wire _w9364_ ;
	wire _w9365_ ;
	wire _w9366_ ;
	wire _w9367_ ;
	wire _w9368_ ;
	wire _w9369_ ;
	wire _w9370_ ;
	wire _w9371_ ;
	wire _w9372_ ;
	wire _w9373_ ;
	wire _w9374_ ;
	wire _w9375_ ;
	wire _w9376_ ;
	wire _w9377_ ;
	wire _w9378_ ;
	wire _w9379_ ;
	wire _w9380_ ;
	wire _w9381_ ;
	wire _w9382_ ;
	wire _w9383_ ;
	wire _w9384_ ;
	wire _w9385_ ;
	wire _w9386_ ;
	wire _w9387_ ;
	wire _w9388_ ;
	wire _w9389_ ;
	wire _w9390_ ;
	wire _w9391_ ;
	wire _w9392_ ;
	wire _w9393_ ;
	wire _w9394_ ;
	wire _w9395_ ;
	wire _w9396_ ;
	wire _w9397_ ;
	wire _w9398_ ;
	wire _w9399_ ;
	wire _w9400_ ;
	wire _w9401_ ;
	wire _w9402_ ;
	wire _w9403_ ;
	wire _w9404_ ;
	wire _w9405_ ;
	wire _w9406_ ;
	wire _w9407_ ;
	wire _w9408_ ;
	wire _w9409_ ;
	wire _w9410_ ;
	wire _w9411_ ;
	wire _w9412_ ;
	wire _w9413_ ;
	wire _w9414_ ;
	wire _w9415_ ;
	wire _w9416_ ;
	wire _w9417_ ;
	wire _w9418_ ;
	wire _w9419_ ;
	wire _w9420_ ;
	wire _w9421_ ;
	wire _w9422_ ;
	wire _w9423_ ;
	wire _w9424_ ;
	wire _w9425_ ;
	wire _w9426_ ;
	wire _w9427_ ;
	wire _w9428_ ;
	wire _w9429_ ;
	wire _w9430_ ;
	wire _w9431_ ;
	wire _w9432_ ;
	wire _w9433_ ;
	wire _w9434_ ;
	wire _w9435_ ;
	wire _w9436_ ;
	wire _w9437_ ;
	wire _w9438_ ;
	wire _w9439_ ;
	wire _w9440_ ;
	wire _w9441_ ;
	wire _w9442_ ;
	wire _w9443_ ;
	wire _w9444_ ;
	wire _w9445_ ;
	wire _w9446_ ;
	wire _w9447_ ;
	wire _w9448_ ;
	wire _w9449_ ;
	wire _w9450_ ;
	wire _w9451_ ;
	wire _w9452_ ;
	wire _w9453_ ;
	wire _w9454_ ;
	wire _w9455_ ;
	wire _w9456_ ;
	wire _w9457_ ;
	wire _w9458_ ;
	wire _w9459_ ;
	wire _w9460_ ;
	wire _w9461_ ;
	wire _w9462_ ;
	wire _w9463_ ;
	wire _w9464_ ;
	wire _w9465_ ;
	wire _w9466_ ;
	wire _w9467_ ;
	wire _w9468_ ;
	wire _w9469_ ;
	wire _w9470_ ;
	wire _w9471_ ;
	wire _w9472_ ;
	wire _w9473_ ;
	wire _w9474_ ;
	wire _w9475_ ;
	wire _w9476_ ;
	wire _w9477_ ;
	wire _w9478_ ;
	wire _w9479_ ;
	wire _w9480_ ;
	wire _w9481_ ;
	wire _w9482_ ;
	wire _w9483_ ;
	wire _w9484_ ;
	wire _w9485_ ;
	wire _w9486_ ;
	wire _w9487_ ;
	wire _w9488_ ;
	wire _w9489_ ;
	wire _w9490_ ;
	wire _w9491_ ;
	wire _w9492_ ;
	wire _w9493_ ;
	wire _w9494_ ;
	wire _w9495_ ;
	wire _w9496_ ;
	wire _w9497_ ;
	wire _w9498_ ;
	wire _w9499_ ;
	wire _w9500_ ;
	wire _w9501_ ;
	wire _w9502_ ;
	wire _w9503_ ;
	wire _w9504_ ;
	wire _w9505_ ;
	wire _w9506_ ;
	wire _w9507_ ;
	wire _w9508_ ;
	wire _w9509_ ;
	wire _w9510_ ;
	wire _w9511_ ;
	wire _w9512_ ;
	wire _w9513_ ;
	wire _w9514_ ;
	wire _w9515_ ;
	wire _w9516_ ;
	wire _w9517_ ;
	wire _w9518_ ;
	wire _w9519_ ;
	wire _w9520_ ;
	wire _w9521_ ;
	wire _w9522_ ;
	wire _w9523_ ;
	wire _w9524_ ;
	wire _w9525_ ;
	wire _w9526_ ;
	wire _w9527_ ;
	wire _w9528_ ;
	wire _w9529_ ;
	wire _w9530_ ;
	wire _w9531_ ;
	wire _w9532_ ;
	wire _w9533_ ;
	wire _w9534_ ;
	wire _w9535_ ;
	wire _w9536_ ;
	wire _w9537_ ;
	wire _w9538_ ;
	wire _w9539_ ;
	wire _w9540_ ;
	wire _w9541_ ;
	wire _w9542_ ;
	wire _w9543_ ;
	wire _w9544_ ;
	wire _w9545_ ;
	wire _w9546_ ;
	wire _w9547_ ;
	wire _w9548_ ;
	wire _w9549_ ;
	wire _w9550_ ;
	wire _w9551_ ;
	wire _w9552_ ;
	wire _w9553_ ;
	wire _w9554_ ;
	wire _w9555_ ;
	wire _w9556_ ;
	wire _w9557_ ;
	wire _w9558_ ;
	wire _w9559_ ;
	wire _w9560_ ;
	wire _w9561_ ;
	wire _w9562_ ;
	wire _w9563_ ;
	wire _w9564_ ;
	wire _w9565_ ;
	wire _w9566_ ;
	wire _w9567_ ;
	wire _w9568_ ;
	wire _w9569_ ;
	wire _w9570_ ;
	wire _w9571_ ;
	wire _w9572_ ;
	wire _w9573_ ;
	wire _w9574_ ;
	wire _w9575_ ;
	wire _w9576_ ;
	wire _w9577_ ;
	wire _w9578_ ;
	wire _w9579_ ;
	wire _w9580_ ;
	wire _w9581_ ;
	wire _w9582_ ;
	wire _w9583_ ;
	wire _w9584_ ;
	wire _w9585_ ;
	wire _w9586_ ;
	wire _w9587_ ;
	wire _w9588_ ;
	wire _w9589_ ;
	wire _w9590_ ;
	wire _w9591_ ;
	wire _w9592_ ;
	wire _w9593_ ;
	wire _w9594_ ;
	wire _w9595_ ;
	wire _w9596_ ;
	wire _w9597_ ;
	wire _w9598_ ;
	wire _w9599_ ;
	wire _w9600_ ;
	wire _w9601_ ;
	wire _w9602_ ;
	wire _w9603_ ;
	wire _w9604_ ;
	wire _w9605_ ;
	wire _w9606_ ;
	wire _w9607_ ;
	wire _w9608_ ;
	wire _w9609_ ;
	wire _w9610_ ;
	wire _w9611_ ;
	wire _w9612_ ;
	wire _w9613_ ;
	wire _w9614_ ;
	wire _w9615_ ;
	wire _w9616_ ;
	wire _w9617_ ;
	wire _w9618_ ;
	wire _w9619_ ;
	wire _w9620_ ;
	wire _w9621_ ;
	wire _w9622_ ;
	wire _w9623_ ;
	wire _w9624_ ;
	wire _w9625_ ;
	wire _w9626_ ;
	wire _w9627_ ;
	wire _w9628_ ;
	wire _w9629_ ;
	wire _w9630_ ;
	wire _w9631_ ;
	wire _w9632_ ;
	wire _w9633_ ;
	wire _w9634_ ;
	wire _w9635_ ;
	wire _w9636_ ;
	wire _w9637_ ;
	wire _w9638_ ;
	wire _w9639_ ;
	wire _w9640_ ;
	wire _w9641_ ;
	wire _w9642_ ;
	wire _w9643_ ;
	wire _w9644_ ;
	wire _w9645_ ;
	wire _w9646_ ;
	wire _w9647_ ;
	wire _w9648_ ;
	wire _w9649_ ;
	wire _w9650_ ;
	wire _w9651_ ;
	wire _w9652_ ;
	wire _w9653_ ;
	wire _w9654_ ;
	wire _w9655_ ;
	wire _w9656_ ;
	wire _w9657_ ;
	wire _w9658_ ;
	wire _w9659_ ;
	wire _w9660_ ;
	wire _w9661_ ;
	wire _w9662_ ;
	wire _w9663_ ;
	wire _w9664_ ;
	wire _w9665_ ;
	wire _w9666_ ;
	wire _w9667_ ;
	wire _w9668_ ;
	wire _w9669_ ;
	wire _w9670_ ;
	wire _w9671_ ;
	wire _w9672_ ;
	wire _w9673_ ;
	wire _w9674_ ;
	wire _w9675_ ;
	wire _w9676_ ;
	wire _w9677_ ;
	wire _w9678_ ;
	wire _w9679_ ;
	wire _w9680_ ;
	wire _w9681_ ;
	wire _w9682_ ;
	wire _w9683_ ;
	wire _w9684_ ;
	wire _w9685_ ;
	wire _w9686_ ;
	wire _w9687_ ;
	wire _w9688_ ;
	wire _w9689_ ;
	wire _w9690_ ;
	wire _w9691_ ;
	wire _w9692_ ;
	wire _w9693_ ;
	wire _w9694_ ;
	wire _w9695_ ;
	wire _w9696_ ;
	wire _w9697_ ;
	wire _w9698_ ;
	wire _w9699_ ;
	wire _w9700_ ;
	wire _w9701_ ;
	wire _w9702_ ;
	wire _w9703_ ;
	wire _w9704_ ;
	wire _w9705_ ;
	wire _w9706_ ;
	wire _w9707_ ;
	wire _w9708_ ;
	wire _w9709_ ;
	wire _w9710_ ;
	wire _w9711_ ;
	wire _w9712_ ;
	wire _w9713_ ;
	wire _w9714_ ;
	wire _w9715_ ;
	wire _w9716_ ;
	wire _w9717_ ;
	wire _w9718_ ;
	wire _w9719_ ;
	wire _w9720_ ;
	wire _w9721_ ;
	wire _w9722_ ;
	wire _w9723_ ;
	wire _w9724_ ;
	wire _w9725_ ;
	wire _w9726_ ;
	wire _w9727_ ;
	wire _w9728_ ;
	wire _w9729_ ;
	wire _w9730_ ;
	wire _w9731_ ;
	wire _w9732_ ;
	wire _w9733_ ;
	wire _w9734_ ;
	wire _w9735_ ;
	wire _w9736_ ;
	wire _w9737_ ;
	wire _w9738_ ;
	wire _w9739_ ;
	wire _w9740_ ;
	wire _w9741_ ;
	wire _w9742_ ;
	wire _w9743_ ;
	wire _w9744_ ;
	wire _w9745_ ;
	wire _w9746_ ;
	wire _w9747_ ;
	wire _w9748_ ;
	wire _w9749_ ;
	wire _w9750_ ;
	wire _w9751_ ;
	wire _w9752_ ;
	wire _w9753_ ;
	wire _w9754_ ;
	wire _w9755_ ;
	wire _w9756_ ;
	wire _w9757_ ;
	wire _w9758_ ;
	wire _w9759_ ;
	wire _w9760_ ;
	wire _w9761_ ;
	wire _w9762_ ;
	wire _w9763_ ;
	wire _w9764_ ;
	wire _w9765_ ;
	wire _w9766_ ;
	wire _w9767_ ;
	wire _w9768_ ;
	wire _w9769_ ;
	wire _w9770_ ;
	wire _w9771_ ;
	wire _w9772_ ;
	wire _w9773_ ;
	wire _w9774_ ;
	wire _w9775_ ;
	wire _w9776_ ;
	wire _w9777_ ;
	wire _w9778_ ;
	wire _w9779_ ;
	wire _w9780_ ;
	wire _w9781_ ;
	wire _w9782_ ;
	wire _w9783_ ;
	wire _w9784_ ;
	wire _w9785_ ;
	wire _w9786_ ;
	wire _w9787_ ;
	wire _w9788_ ;
	wire _w9789_ ;
	wire _w9790_ ;
	wire _w9791_ ;
	wire _w9792_ ;
	wire _w9793_ ;
	wire _w9794_ ;
	wire _w9795_ ;
	wire _w9796_ ;
	wire _w9797_ ;
	wire _w9798_ ;
	wire _w9799_ ;
	wire _w9800_ ;
	wire _w9801_ ;
	wire _w9802_ ;
	wire _w9803_ ;
	wire _w9804_ ;
	wire _w9805_ ;
	wire _w9806_ ;
	wire _w9807_ ;
	wire _w9808_ ;
	wire _w9809_ ;
	wire _w9810_ ;
	wire _w9811_ ;
	wire _w9812_ ;
	wire _w9813_ ;
	wire _w9814_ ;
	wire _w9815_ ;
	wire _w9816_ ;
	wire _w9817_ ;
	wire _w9818_ ;
	wire _w9819_ ;
	wire _w9820_ ;
	wire _w9821_ ;
	wire _w9822_ ;
	wire _w9823_ ;
	wire _w9824_ ;
	wire _w9825_ ;
	wire _w9826_ ;
	wire _w9827_ ;
	wire _w9828_ ;
	wire _w9829_ ;
	wire _w9830_ ;
	wire _w9831_ ;
	wire _w9832_ ;
	wire _w9833_ ;
	wire _w9834_ ;
	wire _w9835_ ;
	wire _w9836_ ;
	wire _w9837_ ;
	wire _w9838_ ;
	wire _w9839_ ;
	wire _w9840_ ;
	wire _w9841_ ;
	wire _w9842_ ;
	wire _w9843_ ;
	wire _w9844_ ;
	wire _w9845_ ;
	wire _w9846_ ;
	wire _w9847_ ;
	wire _w9848_ ;
	wire _w9849_ ;
	wire _w9850_ ;
	wire _w9851_ ;
	wire _w9852_ ;
	wire _w9853_ ;
	wire _w9854_ ;
	wire _w9855_ ;
	wire _w9856_ ;
	wire _w9857_ ;
	wire _w9858_ ;
	wire _w9859_ ;
	wire _w9860_ ;
	wire _w9861_ ;
	wire _w9862_ ;
	wire _w9863_ ;
	wire _w9864_ ;
	wire _w9865_ ;
	wire _w9866_ ;
	wire _w9867_ ;
	wire _w9868_ ;
	wire _w9869_ ;
	wire _w9870_ ;
	wire _w9871_ ;
	wire _w9872_ ;
	wire _w9873_ ;
	wire _w9874_ ;
	wire _w9875_ ;
	wire _w9876_ ;
	wire _w9877_ ;
	wire _w9878_ ;
	wire _w9879_ ;
	wire _w9880_ ;
	wire _w9881_ ;
	wire _w9882_ ;
	wire _w9883_ ;
	wire _w9884_ ;
	wire _w9885_ ;
	wire _w9886_ ;
	wire _w9887_ ;
	wire _w9888_ ;
	wire _w9889_ ;
	wire _w9890_ ;
	wire _w9891_ ;
	wire _w9892_ ;
	wire _w9893_ ;
	wire _w9894_ ;
	wire _w9895_ ;
	wire _w9896_ ;
	wire _w9897_ ;
	wire _w9898_ ;
	wire _w9899_ ;
	wire _w9900_ ;
	wire _w9901_ ;
	wire _w9902_ ;
	wire _w9903_ ;
	wire _w9904_ ;
	wire _w9905_ ;
	wire _w9906_ ;
	wire _w9907_ ;
	wire _w9908_ ;
	wire _w9909_ ;
	wire _w9910_ ;
	wire _w9911_ ;
	wire _w9912_ ;
	wire _w9913_ ;
	wire _w9914_ ;
	wire _w9915_ ;
	wire _w9916_ ;
	wire _w9917_ ;
	wire _w9918_ ;
	wire _w9919_ ;
	wire _w9920_ ;
	wire _w9921_ ;
	wire _w9922_ ;
	wire _w9923_ ;
	wire _w9924_ ;
	wire _w9925_ ;
	wire _w9926_ ;
	wire _w9927_ ;
	wire _w9928_ ;
	wire _w9929_ ;
	wire _w9930_ ;
	wire _w9931_ ;
	wire _w9932_ ;
	wire _w9933_ ;
	wire _w9934_ ;
	wire _w9935_ ;
	wire _w9936_ ;
	wire _w9937_ ;
	wire _w9938_ ;
	wire _w9939_ ;
	wire _w9940_ ;
	wire _w9941_ ;
	wire _w9942_ ;
	wire _w9943_ ;
	wire _w9944_ ;
	wire _w9945_ ;
	wire _w9946_ ;
	wire _w9947_ ;
	wire _w9948_ ;
	wire _w9949_ ;
	wire _w9950_ ;
	wire _w9951_ ;
	wire _w9952_ ;
	wire _w9953_ ;
	wire _w9954_ ;
	wire _w9955_ ;
	wire _w9956_ ;
	wire _w9957_ ;
	wire _w9958_ ;
	wire _w9959_ ;
	wire _w9960_ ;
	wire _w9961_ ;
	wire _w9962_ ;
	wire _w9963_ ;
	wire _w9964_ ;
	wire _w9965_ ;
	wire _w9966_ ;
	wire _w9967_ ;
	wire _w9968_ ;
	wire _w9969_ ;
	wire _w9970_ ;
	wire _w9971_ ;
	wire _w9972_ ;
	wire _w9973_ ;
	wire _w9974_ ;
	wire _w9975_ ;
	wire _w9976_ ;
	wire _w9977_ ;
	wire _w9978_ ;
	wire _w9979_ ;
	wire _w9980_ ;
	wire _w9981_ ;
	wire _w9982_ ;
	wire _w9983_ ;
	wire _w9984_ ;
	wire _w9985_ ;
	wire _w9986_ ;
	wire _w9987_ ;
	wire _w9988_ ;
	wire _w9989_ ;
	wire _w9990_ ;
	wire _w9991_ ;
	wire _w9992_ ;
	wire _w9993_ ;
	wire _w9994_ ;
	wire _w9995_ ;
	wire _w9996_ ;
	wire _w9997_ ;
	wire _w9998_ ;
	wire _w9999_ ;
	wire _w10000_ ;
	wire _w10001_ ;
	wire _w10002_ ;
	wire _w10003_ ;
	wire _w10004_ ;
	wire _w10005_ ;
	wire _w10006_ ;
	wire _w10007_ ;
	wire _w10008_ ;
	wire _w10009_ ;
	wire _w10010_ ;
	wire _w10011_ ;
	wire _w10012_ ;
	wire _w10013_ ;
	wire _w10014_ ;
	wire _w10015_ ;
	wire _w10016_ ;
	wire _w10017_ ;
	wire _w10018_ ;
	wire _w10019_ ;
	wire _w10020_ ;
	wire _w10021_ ;
	wire _w10022_ ;
	wire _w10023_ ;
	wire _w10024_ ;
	wire _w10025_ ;
	wire _w10026_ ;
	wire _w10027_ ;
	wire _w10028_ ;
	wire _w10029_ ;
	wire _w10030_ ;
	wire _w10031_ ;
	wire _w10032_ ;
	wire _w10033_ ;
	wire _w10034_ ;
	wire _w10035_ ;
	wire _w10036_ ;
	wire _w10037_ ;
	wire _w10038_ ;
	wire _w10039_ ;
	wire _w10040_ ;
	wire _w10041_ ;
	wire _w10042_ ;
	wire _w10043_ ;
	wire _w10044_ ;
	wire _w10045_ ;
	wire _w10046_ ;
	wire _w10047_ ;
	wire _w10048_ ;
	wire _w10049_ ;
	wire _w10050_ ;
	wire _w10051_ ;
	wire _w10052_ ;
	wire _w10053_ ;
	wire _w10054_ ;
	wire _w10055_ ;
	wire _w10056_ ;
	wire _w10057_ ;
	wire _w10058_ ;
	wire _w10059_ ;
	wire _w10060_ ;
	wire _w10061_ ;
	wire _w10062_ ;
	wire _w10063_ ;
	wire _w10064_ ;
	wire _w10065_ ;
	wire _w10066_ ;
	wire _w10067_ ;
	wire _w10068_ ;
	wire _w10069_ ;
	wire _w10070_ ;
	wire _w10071_ ;
	wire _w10072_ ;
	wire _w10073_ ;
	wire _w10074_ ;
	wire _w10075_ ;
	wire _w10076_ ;
	wire _w10077_ ;
	wire _w10078_ ;
	wire _w10079_ ;
	wire _w10080_ ;
	wire _w10081_ ;
	wire _w10082_ ;
	wire _w10083_ ;
	wire _w10084_ ;
	wire _w10085_ ;
	wire _w10086_ ;
	wire _w10087_ ;
	wire _w10088_ ;
	wire _w10089_ ;
	wire _w10090_ ;
	wire _w10091_ ;
	wire _w10092_ ;
	wire _w10093_ ;
	wire _w10094_ ;
	wire _w10095_ ;
	wire _w10096_ ;
	wire _w10097_ ;
	wire _w10098_ ;
	wire _w10099_ ;
	wire _w10100_ ;
	wire _w10101_ ;
	wire _w10102_ ;
	wire _w10103_ ;
	wire _w10104_ ;
	wire _w10105_ ;
	wire _w10106_ ;
	wire _w10107_ ;
	wire _w10108_ ;
	wire _w10109_ ;
	wire _w10110_ ;
	wire _w10111_ ;
	wire _w10112_ ;
	wire _w10113_ ;
	wire _w10114_ ;
	wire _w10115_ ;
	wire _w10116_ ;
	wire _w10117_ ;
	wire _w10118_ ;
	wire _w10119_ ;
	wire _w10120_ ;
	wire _w10121_ ;
	wire _w10122_ ;
	wire _w10123_ ;
	wire _w10124_ ;
	wire _w10125_ ;
	wire _w10126_ ;
	wire _w10127_ ;
	wire _w10128_ ;
	wire _w10129_ ;
	wire _w10130_ ;
	wire _w10131_ ;
	wire _w10132_ ;
	wire _w10133_ ;
	wire _w10134_ ;
	wire _w10135_ ;
	wire _w10136_ ;
	wire _w10137_ ;
	wire _w10138_ ;
	wire _w10139_ ;
	wire _w10140_ ;
	wire _w10141_ ;
	wire _w10142_ ;
	wire _w10143_ ;
	wire _w10144_ ;
	wire _w10145_ ;
	wire _w10146_ ;
	wire _w10147_ ;
	wire _w10148_ ;
	wire _w10149_ ;
	wire _w10150_ ;
	wire _w10151_ ;
	wire _w10152_ ;
	wire _w10153_ ;
	wire _w10154_ ;
	wire _w10155_ ;
	wire _w10156_ ;
	wire _w10157_ ;
	wire _w10158_ ;
	wire _w10159_ ;
	wire _w10160_ ;
	wire _w10161_ ;
	wire _w10162_ ;
	wire _w10163_ ;
	wire _w10164_ ;
	wire _w10165_ ;
	wire _w10166_ ;
	wire _w10167_ ;
	wire _w10168_ ;
	wire _w10169_ ;
	wire _w10170_ ;
	wire _w10171_ ;
	wire _w10172_ ;
	wire _w10173_ ;
	wire _w10174_ ;
	wire _w10175_ ;
	wire _w10176_ ;
	wire _w10177_ ;
	wire _w10178_ ;
	wire _w10179_ ;
	wire _w10180_ ;
	wire _w10181_ ;
	wire _w10182_ ;
	wire _w10183_ ;
	wire _w10184_ ;
	wire _w10185_ ;
	wire _w10186_ ;
	wire _w10187_ ;
	wire _w10188_ ;
	wire _w10189_ ;
	wire _w10190_ ;
	wire _w10191_ ;
	wire _w10192_ ;
	wire _w10193_ ;
	wire _w10194_ ;
	wire _w10195_ ;
	wire _w10196_ ;
	wire _w10197_ ;
	wire _w10198_ ;
	wire _w10199_ ;
	wire _w10200_ ;
	wire _w10201_ ;
	wire _w10202_ ;
	wire _w10203_ ;
	wire _w10204_ ;
	wire _w10205_ ;
	wire _w10206_ ;
	wire _w10207_ ;
	wire _w10208_ ;
	wire _w10209_ ;
	wire _w10210_ ;
	wire _w10211_ ;
	wire _w10212_ ;
	wire _w10213_ ;
	wire _w10214_ ;
	wire _w10215_ ;
	wire _w10216_ ;
	wire _w10217_ ;
	wire _w10218_ ;
	wire _w10219_ ;
	wire _w10220_ ;
	wire _w10221_ ;
	wire _w10222_ ;
	wire _w10223_ ;
	wire _w10224_ ;
	wire _w10225_ ;
	wire _w10226_ ;
	wire _w10227_ ;
	wire _w10228_ ;
	wire _w10229_ ;
	wire _w10230_ ;
	wire _w10231_ ;
	wire _w10232_ ;
	wire _w10233_ ;
	wire _w10234_ ;
	wire _w10235_ ;
	wire _w10236_ ;
	wire _w10237_ ;
	wire _w10238_ ;
	wire _w10239_ ;
	wire _w10240_ ;
	wire _w10241_ ;
	wire _w10242_ ;
	wire _w10243_ ;
	wire _w10244_ ;
	wire _w10245_ ;
	wire _w10246_ ;
	wire _w10247_ ;
	wire _w10248_ ;
	wire _w10249_ ;
	wire _w10250_ ;
	wire _w10251_ ;
	wire _w10252_ ;
	wire _w10253_ ;
	wire _w10254_ ;
	wire _w10255_ ;
	wire _w10256_ ;
	wire _w10257_ ;
	wire _w10258_ ;
	wire _w10259_ ;
	wire _w10260_ ;
	wire _w10261_ ;
	wire _w10262_ ;
	wire _w10263_ ;
	wire _w10264_ ;
	wire _w10265_ ;
	wire _w10266_ ;
	wire _w10267_ ;
	wire _w10268_ ;
	wire _w10269_ ;
	wire _w10270_ ;
	wire _w10271_ ;
	wire _w10272_ ;
	wire _w10273_ ;
	wire _w10274_ ;
	wire _w10275_ ;
	wire _w10276_ ;
	wire _w10277_ ;
	wire _w10278_ ;
	wire _w10279_ ;
	wire _w10280_ ;
	wire _w10281_ ;
	wire _w10282_ ;
	wire _w10283_ ;
	wire _w10284_ ;
	wire _w10285_ ;
	wire _w10286_ ;
	wire _w10287_ ;
	wire _w10288_ ;
	wire _w10289_ ;
	wire _w10290_ ;
	wire _w10291_ ;
	wire _w10292_ ;
	wire _w10293_ ;
	wire _w10294_ ;
	wire _w10295_ ;
	wire _w10296_ ;
	wire _w10297_ ;
	wire _w10298_ ;
	wire _w10299_ ;
	wire _w10300_ ;
	wire _w10301_ ;
	wire _w10302_ ;
	wire _w10303_ ;
	wire _w10304_ ;
	wire _w10305_ ;
	wire _w10306_ ;
	wire _w10307_ ;
	wire _w10308_ ;
	wire _w10309_ ;
	wire _w10310_ ;
	wire _w10311_ ;
	wire _w10312_ ;
	wire _w10313_ ;
	wire _w10314_ ;
	wire _w10315_ ;
	wire _w10316_ ;
	wire _w10317_ ;
	wire _w10318_ ;
	wire _w10319_ ;
	wire _w10320_ ;
	wire _w10321_ ;
	wire _w10322_ ;
	wire _w10323_ ;
	wire _w10324_ ;
	wire _w10325_ ;
	wire _w10326_ ;
	wire _w10327_ ;
	wire _w10328_ ;
	wire _w10329_ ;
	wire _w10330_ ;
	wire _w10331_ ;
	wire _w10332_ ;
	wire _w10333_ ;
	wire _w10334_ ;
	wire _w10335_ ;
	wire _w10336_ ;
	wire _w10337_ ;
	wire _w10338_ ;
	wire _w10339_ ;
	wire _w10340_ ;
	wire _w10341_ ;
	wire _w10342_ ;
	wire _w10343_ ;
	wire _w10344_ ;
	wire _w10345_ ;
	wire _w10346_ ;
	wire _w10347_ ;
	wire _w10348_ ;
	wire _w10349_ ;
	wire _w10350_ ;
	wire _w10351_ ;
	wire _w10352_ ;
	wire _w10353_ ;
	wire _w10354_ ;
	wire _w10355_ ;
	wire _w10356_ ;
	wire _w10357_ ;
	wire _w10358_ ;
	wire _w10359_ ;
	wire _w10360_ ;
	wire _w10361_ ;
	wire _w10362_ ;
	wire _w10363_ ;
	wire _w10364_ ;
	wire _w10365_ ;
	wire _w10366_ ;
	wire _w10367_ ;
	wire _w10368_ ;
	wire _w10369_ ;
	wire _w10370_ ;
	wire _w10371_ ;
	wire _w10372_ ;
	wire _w10373_ ;
	wire _w10374_ ;
	wire _w10375_ ;
	wire _w10376_ ;
	wire _w10377_ ;
	wire _w10378_ ;
	wire _w10379_ ;
	wire _w10380_ ;
	wire _w10381_ ;
	wire _w10382_ ;
	wire _w10383_ ;
	wire _w10384_ ;
	wire _w10385_ ;
	wire _w10386_ ;
	wire _w10387_ ;
	wire _w10388_ ;
	wire _w10389_ ;
	wire _w10390_ ;
	wire _w10391_ ;
	wire _w10392_ ;
	wire _w10393_ ;
	wire _w10394_ ;
	wire _w10395_ ;
	wire _w10396_ ;
	wire _w10397_ ;
	wire _w10398_ ;
	wire _w10399_ ;
	wire _w10400_ ;
	wire _w10401_ ;
	wire _w10402_ ;
	wire _w10403_ ;
	wire _w10404_ ;
	wire _w10405_ ;
	wire _w10406_ ;
	wire _w10407_ ;
	wire _w10408_ ;
	wire _w10409_ ;
	wire _w10410_ ;
	wire _w10411_ ;
	wire _w10412_ ;
	wire _w10413_ ;
	wire _w10414_ ;
	wire _w10415_ ;
	wire _w10416_ ;
	wire _w10417_ ;
	wire _w10418_ ;
	wire _w10419_ ;
	wire _w10420_ ;
	wire _w10421_ ;
	wire _w10422_ ;
	wire _w10423_ ;
	wire _w10424_ ;
	wire _w10425_ ;
	wire _w10426_ ;
	wire _w10427_ ;
	wire _w10428_ ;
	wire _w10429_ ;
	wire _w10430_ ;
	wire _w10431_ ;
	wire _w10432_ ;
	wire _w10433_ ;
	wire _w10434_ ;
	wire _w10435_ ;
	wire _w10436_ ;
	wire _w10437_ ;
	wire _w10438_ ;
	wire _w10439_ ;
	wire _w10440_ ;
	wire _w10441_ ;
	wire _w10442_ ;
	wire _w10443_ ;
	wire _w10444_ ;
	wire _w10445_ ;
	wire _w10446_ ;
	wire _w10447_ ;
	wire _w10448_ ;
	wire _w10449_ ;
	wire _w10450_ ;
	wire _w10451_ ;
	wire _w10452_ ;
	wire _w10453_ ;
	wire _w10454_ ;
	wire _w10455_ ;
	wire _w10456_ ;
	wire _w10457_ ;
	wire _w10458_ ;
	wire _w10459_ ;
	wire _w10460_ ;
	wire _w10461_ ;
	wire _w10462_ ;
	wire _w10463_ ;
	wire _w10464_ ;
	wire _w10465_ ;
	wire _w10466_ ;
	wire _w10467_ ;
	wire _w10468_ ;
	wire _w10469_ ;
	wire _w10470_ ;
	wire _w10471_ ;
	wire _w10472_ ;
	wire _w10473_ ;
	wire _w10474_ ;
	wire _w10475_ ;
	wire _w10476_ ;
	wire _w10477_ ;
	wire _w10478_ ;
	wire _w10479_ ;
	wire _w10480_ ;
	wire _w10481_ ;
	wire _w10482_ ;
	wire _w10483_ ;
	wire _w10484_ ;
	wire _w10485_ ;
	wire _w10486_ ;
	wire _w10487_ ;
	wire _w10488_ ;
	wire _w10489_ ;
	wire _w10490_ ;
	wire _w10491_ ;
	wire _w10492_ ;
	wire _w10493_ ;
	wire _w10494_ ;
	wire _w10495_ ;
	wire _w10496_ ;
	wire _w10497_ ;
	wire _w10498_ ;
	wire _w10499_ ;
	wire _w10500_ ;
	wire _w10501_ ;
	wire _w10502_ ;
	wire _w10503_ ;
	wire _w10504_ ;
	wire _w10505_ ;
	wire _w10506_ ;
	wire _w10507_ ;
	wire _w10508_ ;
	wire _w10509_ ;
	wire _w10510_ ;
	wire _w10511_ ;
	wire _w10512_ ;
	wire _w10513_ ;
	wire _w10514_ ;
	wire _w10515_ ;
	wire _w10516_ ;
	wire _w10517_ ;
	wire _w10518_ ;
	wire _w10519_ ;
	wire _w10520_ ;
	wire _w10521_ ;
	wire _w10522_ ;
	wire _w10523_ ;
	wire _w10524_ ;
	wire _w10525_ ;
	wire _w10526_ ;
	wire _w10527_ ;
	wire _w10528_ ;
	wire _w10529_ ;
	wire _w10530_ ;
	wire _w10531_ ;
	wire _w10532_ ;
	wire _w10533_ ;
	wire _w10534_ ;
	wire _w10535_ ;
	wire _w10536_ ;
	wire _w10537_ ;
	wire _w10538_ ;
	wire _w10539_ ;
	wire _w10540_ ;
	wire _w10541_ ;
	wire _w10542_ ;
	wire _w10543_ ;
	wire _w10544_ ;
	wire _w10545_ ;
	wire _w10546_ ;
	wire _w10547_ ;
	wire _w10548_ ;
	wire _w10549_ ;
	wire _w10550_ ;
	wire _w10551_ ;
	wire _w10552_ ;
	wire _w10553_ ;
	wire _w10554_ ;
	wire _w10555_ ;
	wire _w10556_ ;
	wire _w10557_ ;
	wire _w10558_ ;
	wire _w10559_ ;
	wire _w10560_ ;
	wire _w10561_ ;
	wire _w10562_ ;
	wire _w10563_ ;
	wire _w10564_ ;
	wire _w10565_ ;
	wire _w10566_ ;
	wire _w10567_ ;
	wire _w10568_ ;
	wire _w10569_ ;
	wire _w10570_ ;
	wire _w10571_ ;
	wire _w10572_ ;
	wire _w10573_ ;
	wire _w10574_ ;
	wire _w10575_ ;
	wire _w10576_ ;
	wire _w10577_ ;
	wire _w10578_ ;
	wire _w10579_ ;
	wire _w10580_ ;
	wire _w10581_ ;
	wire _w10582_ ;
	wire _w10583_ ;
	wire _w10584_ ;
	wire _w10585_ ;
	wire _w10586_ ;
	wire _w10587_ ;
	wire _w10588_ ;
	wire _w10589_ ;
	wire _w10590_ ;
	wire _w10591_ ;
	wire _w10592_ ;
	wire _w10593_ ;
	wire _w10594_ ;
	wire _w10595_ ;
	wire _w10596_ ;
	wire _w10597_ ;
	wire _w10598_ ;
	wire _w10599_ ;
	wire _w10600_ ;
	wire _w10601_ ;
	wire _w10602_ ;
	wire _w10603_ ;
	wire _w10604_ ;
	wire _w10605_ ;
	wire _w10606_ ;
	wire _w10607_ ;
	wire _w10608_ ;
	wire _w10609_ ;
	wire _w10610_ ;
	wire _w10611_ ;
	wire _w10612_ ;
	wire _w10613_ ;
	wire _w10614_ ;
	wire _w10615_ ;
	wire _w10616_ ;
	wire _w10617_ ;
	wire _w10618_ ;
	wire _w10619_ ;
	wire _w10620_ ;
	wire _w10621_ ;
	wire _w10622_ ;
	wire _w10623_ ;
	wire _w10624_ ;
	wire _w10625_ ;
	wire _w10626_ ;
	wire _w10627_ ;
	wire _w10628_ ;
	wire _w10629_ ;
	wire _w10630_ ;
	wire _w10631_ ;
	wire _w10632_ ;
	wire _w10633_ ;
	wire _w10634_ ;
	wire _w10635_ ;
	wire _w10636_ ;
	wire _w10637_ ;
	wire _w10638_ ;
	wire _w10639_ ;
	wire _w10640_ ;
	wire _w10641_ ;
	wire _w10642_ ;
	wire _w10643_ ;
	wire _w10644_ ;
	wire _w10645_ ;
	wire _w10646_ ;
	wire _w10647_ ;
	wire _w10648_ ;
	wire _w10649_ ;
	wire _w10650_ ;
	wire _w10651_ ;
	wire _w10652_ ;
	wire _w10653_ ;
	wire _w10654_ ;
	wire _w10655_ ;
	wire _w10656_ ;
	wire _w10657_ ;
	wire _w10658_ ;
	wire _w10659_ ;
	wire _w10660_ ;
	wire _w10661_ ;
	wire _w10662_ ;
	wire _w10663_ ;
	wire _w10664_ ;
	wire _w10665_ ;
	wire _w10666_ ;
	wire _w10667_ ;
	wire _w10668_ ;
	wire _w10669_ ;
	wire _w10670_ ;
	wire _w10671_ ;
	wire _w10672_ ;
	wire _w10673_ ;
	wire _w10674_ ;
	wire _w10675_ ;
	wire _w10676_ ;
	wire _w10677_ ;
	wire _w10678_ ;
	wire _w10679_ ;
	wire _w10680_ ;
	wire _w10681_ ;
	wire _w10682_ ;
	wire _w10683_ ;
	wire _w10684_ ;
	wire _w10685_ ;
	wire _w10686_ ;
	wire _w10687_ ;
	wire _w10688_ ;
	wire _w10689_ ;
	wire _w10690_ ;
	wire _w10691_ ;
	wire _w10692_ ;
	wire _w10693_ ;
	wire _w10694_ ;
	wire _w10695_ ;
	wire _w10696_ ;
	wire _w10697_ ;
	wire _w10698_ ;
	wire _w10699_ ;
	wire _w10700_ ;
	wire _w10701_ ;
	wire _w10702_ ;
	wire _w10703_ ;
	wire _w10704_ ;
	wire _w10705_ ;
	wire _w10706_ ;
	wire _w10707_ ;
	wire _w10708_ ;
	wire _w10709_ ;
	wire _w10710_ ;
	wire _w10711_ ;
	wire _w10712_ ;
	wire _w10713_ ;
	wire _w10714_ ;
	wire _w10715_ ;
	wire _w10716_ ;
	wire _w10717_ ;
	wire _w10718_ ;
	wire _w10719_ ;
	wire _w10720_ ;
	wire _w10721_ ;
	wire _w10722_ ;
	wire _w10723_ ;
	wire _w10724_ ;
	wire _w10725_ ;
	wire _w10726_ ;
	wire _w10727_ ;
	wire _w10728_ ;
	wire _w10729_ ;
	wire _w10730_ ;
	wire _w10731_ ;
	wire _w10732_ ;
	wire _w10733_ ;
	wire _w10734_ ;
	wire _w10735_ ;
	wire _w10736_ ;
	wire _w10737_ ;
	wire _w10738_ ;
	wire _w10739_ ;
	wire _w10740_ ;
	wire _w10741_ ;
	wire _w10742_ ;
	wire _w10743_ ;
	wire _w10744_ ;
	wire _w10745_ ;
	wire _w10746_ ;
	wire _w10747_ ;
	wire _w10748_ ;
	wire _w10749_ ;
	wire _w10750_ ;
	wire _w10751_ ;
	wire _w10752_ ;
	wire _w10753_ ;
	wire _w10754_ ;
	wire _w10755_ ;
	wire _w10756_ ;
	wire _w10757_ ;
	wire _w10758_ ;
	wire _w10759_ ;
	wire _w10760_ ;
	wire _w10761_ ;
	wire _w10762_ ;
	wire _w10763_ ;
	wire _w10764_ ;
	wire _w10765_ ;
	wire _w10766_ ;
	wire _w10767_ ;
	wire _w10768_ ;
	wire _w10769_ ;
	wire _w10770_ ;
	wire _w10771_ ;
	wire _w10772_ ;
	wire _w10773_ ;
	wire _w10774_ ;
	wire _w10775_ ;
	wire _w10776_ ;
	wire _w10777_ ;
	wire _w10778_ ;
	wire _w10779_ ;
	wire _w10780_ ;
	wire _w10781_ ;
	wire _w10782_ ;
	wire _w10783_ ;
	wire _w10784_ ;
	wire _w10785_ ;
	wire _w10786_ ;
	wire _w10787_ ;
	wire _w10788_ ;
	wire _w10789_ ;
	wire _w10790_ ;
	wire _w10791_ ;
	wire _w10792_ ;
	wire _w10793_ ;
	wire _w10794_ ;
	wire _w10795_ ;
	wire _w10796_ ;
	wire _w10797_ ;
	wire _w10798_ ;
	wire _w10799_ ;
	wire _w10800_ ;
	wire _w10801_ ;
	wire _w10802_ ;
	wire _w10803_ ;
	wire _w10804_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w532_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w533_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		_w532_,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w535_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w536_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		_w535_,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		_w534_,
		_w537_,
		_w538_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\sa13_reg[2]/P0001 ,
		_w538_,
		_w539_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\sa13_reg[7]/NET0131 ,
		_w535_,
		_w540_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		\sa13_reg[3]/P0001 ,
		_w540_,
		_w541_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\sa13_reg[4]/P0001 ,
		_w541_,
		_w542_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w543_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\sa13_reg[3]/P0001 ,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\sa13_reg[4]/P0001 ,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w542_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w547_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		_w536_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w549_
	);
	LUT2 #(
		.INIT('h2)
	) name18 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		_w550_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		_w549_,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w548_,
		_w551_,
		_w552_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		_w546_,
		_w552_,
		_w553_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		\sa13_reg[2]/P0001 ,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w555_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w556_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\sa13_reg[5]/P0001 ,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		_w555_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w559_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		\sa13_reg[3]/P0001 ,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		\sa13_reg[4]/P0001 ,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w558_,
		_w561_,
		_w562_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w563_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[5]/P0001 ,
		_w564_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		\sa13_reg[3]/P0001 ,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		_w563_,
		_w565_,
		_w566_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\sa13_reg[4]/P0001 ,
		_w543_,
		_w567_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		\sa13_reg[5]/P0001 ,
		_w549_,
		_w568_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		\sa13_reg[4]/P0001 ,
		_w568_,
		_w569_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w570_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w563_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\sa13_reg[3]/P0001 ,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w567_,
		_w569_,
		_w573_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		_w572_,
		_w573_,
		_w574_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		\sa13_reg[2]/P0001 ,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		_w562_,
		_w566_,
		_w576_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		_w575_,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		\sa13_reg[1]/P0001 ,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w579_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\sa13_reg[4]/P0001 ,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w581_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w580_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w583_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		\sa13_reg[4]/P0001 ,
		_w583_,
		_w584_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w564_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		_w582_,
		_w585_,
		_w586_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w587_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		_w532_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		\sa13_reg[3]/P0001 ,
		_w557_,
		_w589_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		\sa13_reg[2]/P0001 ,
		_w589_,
		_w590_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		\sa13_reg[5]/P0001 ,
		_w543_,
		_w591_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		\sa13_reg[7]/NET0131 ,
		_w555_,
		_w592_
	);
	LUT2 #(
		.INIT('h2)
	) name61 (
		\sa13_reg[2]/P0001 ,
		_w591_,
		_w593_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		_w592_,
		_w593_,
		_w594_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w590_,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h2)
	) name64 (
		_w586_,
		_w588_,
		_w596_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		_w595_,
		_w596_,
		_w597_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\sa13_reg[1]/P0001 ,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w539_,
		_w554_,
		_w599_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		_w598_,
		_w599_,
		_w600_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		_w578_,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		\sa13_reg[0]/P0001 ,
		_w601_,
		_w602_
	);
	LUT2 #(
		.INIT('h2)
	) name71 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w603_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		\sa13_reg[4]/P0001 ,
		_w579_,
		_w604_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		\sa13_reg[4]/P0001 ,
		_w559_,
		_w605_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w604_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h2)
	) name75 (
		_w603_,
		_w606_,
		_w607_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		\sa13_reg[5]/P0001 ,
		_w555_,
		_w608_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		_w543_,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\sa13_reg[4]/P0001 ,
		_w547_,
		_w610_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w611_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		_w610_,
		_w611_,
		_w612_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		\sa13_reg[1]/P0001 ,
		_w609_,
		_w613_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		_w612_,
		_w613_,
		_w614_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		_w607_,
		_w614_,
		_w615_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		\sa13_reg[3]/P0001 ,
		_w570_,
		_w616_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\sa13_reg[3]/P0001 ,
		_w549_,
		_w617_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		_w616_,
		_w617_,
		_w618_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		\sa13_reg[4]/P0001 ,
		_w618_,
		_w619_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		\sa13_reg[6]/NET0131 ,
		_w533_,
		_w620_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		\sa13_reg[5]/P0001 ,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\sa13_reg[7]/NET0131 ,
		_w621_,
		_w622_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w623_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		_w557_,
		_w623_,
		_w624_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		_w581_,
		_w587_,
		_w625_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		\sa13_reg[1]/P0001 ,
		_w537_,
		_w626_
	);
	LUT2 #(
		.INIT('h4)
	) name95 (
		_w625_,
		_w626_,
		_w627_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		_w624_,
		_w627_,
		_w628_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w619_,
		_w622_,
		_w629_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		_w628_,
		_w629_,
		_w630_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		_w615_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		\sa13_reg[4]/P0001 ,
		_w547_,
		_w632_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		\sa13_reg[3]/P0001 ,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		_w550_,
		_w556_,
		_w634_
	);
	LUT2 #(
		.INIT('h2)
	) name103 (
		\sa13_reg[4]/P0001 ,
		_w583_,
		_w635_
	);
	LUT2 #(
		.INIT('h2)
	) name104 (
		_w634_,
		_w635_,
		_w636_
	);
	LUT2 #(
		.INIT('h4)
	) name105 (
		\sa13_reg[7]/NET0131 ,
		_w533_,
		_w637_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w535_,
		_w637_,
		_w638_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		\sa13_reg[2]/P0001 ,
		_w633_,
		_w639_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		_w636_,
		_w638_,
		_w640_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		_w639_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		\sa13_reg[3]/P0001 ,
		_w610_,
		_w642_
	);
	LUT2 #(
		.INIT('h2)
	) name111 (
		\sa13_reg[2]/P0001 ,
		_w642_,
		_w643_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		_w622_,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w641_,
		_w644_,
		_w645_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		_w631_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		\sa13_reg[0]/P0001 ,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		_w543_,
		_w550_,
		_w648_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\sa13_reg[4]/P0001 ,
		_w648_,
		_w649_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		\sa13_reg[5]/P0001 ,
		_w556_,
		_w650_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		\sa13_reg[3]/P0001 ,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		\sa13_reg[6]/NET0131 ,
		_w580_,
		_w652_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w653_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		_w556_,
		_w653_,
		_w654_
	);
	LUT2 #(
		.INIT('h2)
	) name123 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w655_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		\sa13_reg[5]/P0001 ,
		_w655_,
		_w656_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		_w549_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		_w652_,
		_w654_,
		_w658_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		_w657_,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		\sa13_reg[1]/P0001 ,
		_w659_,
		_w660_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w649_,
		_w651_,
		_w661_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		_w660_,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		\sa13_reg[2]/P0001 ,
		_w662_,
		_w663_
	);
	LUT2 #(
		.INIT('h2)
	) name132 (
		_w568_,
		_w653_,
		_w664_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		\sa13_reg[5]/P0001 ,
		_w567_,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		_w664_,
		_w665_,
		_w666_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		\sa13_reg[2]/P0001 ,
		_w666_,
		_w667_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		_w535_,
		_w653_,
		_w668_
	);
	LUT2 #(
		.INIT('h4)
	) name137 (
		\sa13_reg[6]/NET0131 ,
		_w592_,
		_w669_
	);
	LUT2 #(
		.INIT('h2)
	) name138 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w670_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		_w540_,
		_w670_,
		_w671_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		\sa13_reg[4]/P0001 ,
		_w556_,
		_w672_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		_w623_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		_w668_,
		_w669_,
		_w674_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		_w671_,
		_w673_,
		_w675_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		_w674_,
		_w675_,
		_w676_
	);
	LUT2 #(
		.INIT('h4)
	) name145 (
		_w667_,
		_w676_,
		_w677_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		\sa13_reg[1]/P0001 ,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w581_,
		_w588_,
		_w679_
	);
	LUT2 #(
		.INIT('h2)
	) name148 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[2]/P0001 ,
		_w680_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		_w557_,
		_w655_,
		_w681_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		_w680_,
		_w681_,
		_w682_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		\sa13_reg[5]/P0001 ,
		_w654_,
		_w683_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		_w679_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		_w682_,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h4)
	) name154 (
		_w678_,
		_w685_,
		_w686_
	);
	LUT2 #(
		.INIT('h4)
	) name155 (
		_w663_,
		_w686_,
		_w687_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		_w647_,
		_w687_,
		_w688_
	);
	LUT2 #(
		.INIT('h4)
	) name157 (
		_w602_,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w690_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w691_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		_w690_,
		_w691_,
		_w692_
	);
	LUT2 #(
		.INIT('h2)
	) name161 (
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w693_
	);
	LUT2 #(
		.INIT('h4)
	) name162 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		_w694_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		_w693_,
		_w694_,
		_w695_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		_w692_,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		\sa20_reg[2]/P0001 ,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w698_
	);
	LUT2 #(
		.INIT('h4)
	) name167 (
		\sa20_reg[7]/NET0131 ,
		_w698_,
		_w699_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		\sa20_reg[4]/P0001 ,
		_w699_,
		_w700_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w701_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		_w691_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		\sa20_reg[7]/NET0131 ,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		_w700_,
		_w703_,
		_w704_
	);
	LUT2 #(
		.INIT('h4)
	) name173 (
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w705_
	);
	LUT2 #(
		.INIT('h2)
	) name174 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		_w706_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		_w705_,
		_w706_,
		_w707_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w708_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w709_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		_w708_,
		_w709_,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		_w707_,
		_w710_,
		_w711_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		_w704_,
		_w711_,
		_w712_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		\sa20_reg[2]/P0001 ,
		_w712_,
		_w713_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w714_
	);
	LUT2 #(
		.INIT('h8)
	) name183 (
		_w690_,
		_w714_,
		_w715_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w716_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w717_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		_w716_,
		_w717_,
		_w718_
	);
	LUT2 #(
		.INIT('h4)
	) name187 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w719_
	);
	LUT2 #(
		.INIT('h4)
	) name188 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w720_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		_w719_,
		_w720_,
		_w721_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		_w718_,
		_w721_,
		_w722_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w723_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		\sa20_reg[5]/P0001 ,
		_w723_,
		_w724_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		\sa20_reg[3]/P0001 ,
		_w724_,
		_w725_
	);
	LUT2 #(
		.INIT('h2)
	) name194 (
		_w722_,
		_w725_,
		_w726_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		\sa20_reg[2]/P0001 ,
		_w726_,
		_w727_
	);
	LUT2 #(
		.INIT('h4)
	) name196 (
		\sa20_reg[5]/P0001 ,
		_w693_,
		_w728_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		\sa20_reg[3]/P0001 ,
		_w714_,
		_w729_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		_w728_,
		_w729_,
		_w730_
	);
	LUT2 #(
		.INIT('h2)
	) name199 (
		\sa20_reg[2]/P0001 ,
		_w730_,
		_w731_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		_w715_,
		_w731_,
		_w732_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		_w727_,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		\sa20_reg[1]/P0001 ,
		_w733_,
		_w734_
	);
	LUT2 #(
		.INIT('h4)
	) name203 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w735_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w736_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		_w735_,
		_w736_,
		_w737_
	);
	LUT2 #(
		.INIT('h4)
	) name206 (
		\sa20_reg[4]/P0001 ,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		\sa20_reg[4]/P0001 ,
		_w693_,
		_w739_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		_w694_,
		_w705_,
		_w740_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		_w739_,
		_w740_,
		_w741_
	);
	LUT2 #(
		.INIT('h4)
	) name210 (
		_w738_,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		\sa20_reg[2]/P0001 ,
		_w742_,
		_w743_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w744_
	);
	LUT2 #(
		.INIT('h2)
	) name213 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w745_
	);
	LUT2 #(
		.INIT('h8)
	) name214 (
		_w744_,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		_w747_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		\sa20_reg[5]/P0001 ,
		_w719_,
		_w748_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		_w747_,
		_w748_,
		_w749_
	);
	LUT2 #(
		.INIT('h4)
	) name218 (
		\sa20_reg[6]/NET0131 ,
		_w716_,
		_w750_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		\sa20_reg[5]/P0001 ,
		_w750_,
		_w751_
	);
	LUT2 #(
		.INIT('h4)
	) name220 (
		\sa20_reg[7]/NET0131 ,
		_w751_,
		_w752_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		_w746_,
		_w749_,
		_w753_
	);
	LUT2 #(
		.INIT('h4)
	) name222 (
		_w752_,
		_w753_,
		_w754_
	);
	LUT2 #(
		.INIT('h4)
	) name223 (
		_w743_,
		_w754_,
		_w755_
	);
	LUT2 #(
		.INIT('h2)
	) name224 (
		\sa20_reg[1]/P0001 ,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w697_,
		_w713_,
		_w757_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		_w734_,
		_w757_,
		_w758_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		_w756_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h2)
	) name228 (
		\sa20_reg[0]/P0001 ,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		_w761_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w724_,
		_w761_,
		_w762_
	);
	LUT2 #(
		.INIT('h4)
	) name231 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		_w763_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		_w714_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w765_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		_w706_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		\sa20_reg[4]/P0001 ,
		_w735_,
		_w767_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		_w736_,
		_w767_,
		_w768_
	);
	LUT2 #(
		.INIT('h4)
	) name237 (
		\sa20_reg[6]/NET0131 ,
		_w736_,
		_w769_
	);
	LUT2 #(
		.INIT('h4)
	) name238 (
		\sa20_reg[4]/P0001 ,
		_w769_,
		_w770_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		\sa20_reg[1]/P0001 ,
		_w695_,
		_w771_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		_w764_,
		_w766_,
		_w772_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w771_,
		_w772_,
		_w773_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w762_,
		_w768_,
		_w774_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		_w770_,
		_w774_,
		_w775_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		_w773_,
		_w775_,
		_w776_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w777_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		_w698_,
		_w777_,
		_w778_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		\sa20_reg[4]/P0001 ,
		_w778_,
		_w779_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		\sa20_reg[2]/P0001 ,
		_w710_,
		_w780_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		\sa20_reg[4]/P0001 ,
		_w744_,
		_w781_
	);
	LUT2 #(
		.INIT('h4)
	) name250 (
		\sa20_reg[4]/P0001 ,
		_w717_,
		_w782_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		_w781_,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		_w761_,
		_w780_,
		_w784_
	);
	LUT2 #(
		.INIT('h4)
	) name253 (
		_w783_,
		_w784_,
		_w785_
	);
	LUT2 #(
		.INIT('h2)
	) name254 (
		\sa20_reg[1]/P0001 ,
		_w779_,
		_w786_
	);
	LUT2 #(
		.INIT('h4)
	) name255 (
		_w785_,
		_w786_,
		_w787_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		_w776_,
		_w787_,
		_w788_
	);
	LUT2 #(
		.INIT('h4)
	) name257 (
		\sa20_reg[7]/NET0131 ,
		_w691_,
		_w789_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		_w701_,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		\sa20_reg[4]/P0001 ,
		_w708_,
		_w791_
	);
	LUT2 #(
		.INIT('h2)
	) name260 (
		_w706_,
		_w723_,
		_w792_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w791_,
		_w792_,
		_w793_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w716_,
		_w793_,
		_w794_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		_w698_,
		_w720_,
		_w795_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		\sa20_reg[2]/P0001 ,
		_w795_,
		_w796_
	);
	LUT2 #(
		.INIT('h4)
	) name265 (
		_w790_,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('h4)
	) name266 (
		_w794_,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w799_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		_w708_,
		_w799_,
		_w800_
	);
	LUT2 #(
		.INIT('h2)
	) name269 (
		\sa20_reg[2]/P0001 ,
		_w800_,
		_w801_
	);
	LUT2 #(
		.INIT('h4)
	) name270 (
		_w768_,
		_w801_,
		_w802_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		_w798_,
		_w802_,
		_w803_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w788_,
		_w803_,
		_w804_
	);
	LUT2 #(
		.INIT('h1)
	) name273 (
		\sa20_reg[0]/P0001 ,
		_w804_,
		_w805_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		\sa20_reg[1]/P0001 ,
		\sa20_reg[2]/P0001 ,
		_w806_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		\sa20_reg[4]/P0001 ,
		_w723_,
		_w807_
	);
	LUT2 #(
		.INIT('h4)
	) name276 (
		\sa20_reg[5]/P0001 ,
		_w807_,
		_w808_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		_w723_,
		_w799_,
		_w809_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		\sa20_reg[5]/P0001 ,
		_w745_,
		_w810_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		_w705_,
		_w810_,
		_w811_
	);
	LUT2 #(
		.INIT('h1)
	) name280 (
		_w808_,
		_w809_,
		_w812_
	);
	LUT2 #(
		.INIT('h4)
	) name281 (
		_w811_,
		_w812_,
		_w813_
	);
	LUT2 #(
		.INIT('h2)
	) name282 (
		_w806_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h2)
	) name283 (
		\sa20_reg[1]/P0001 ,
		\sa20_reg[2]/P0001 ,
		_w815_
	);
	LUT2 #(
		.INIT('h4)
	) name284 (
		\sa20_reg[6]/NET0131 ,
		_w745_,
		_w816_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		_w777_,
		_w816_,
		_w817_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		_w815_,
		_w817_,
		_w818_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		_w819_
	);
	LUT2 #(
		.INIT('h4)
	) name288 (
		\sa20_reg[5]/P0001 ,
		_w723_,
		_w820_
	);
	LUT2 #(
		.INIT('h8)
	) name289 (
		_w819_,
		_w820_,
		_w821_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		_w716_,
		_w728_,
		_w822_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		\sa20_reg[2]/P0001 ,
		_w822_,
		_w823_
	);
	LUT2 #(
		.INIT('h4)
	) name292 (
		\sa20_reg[7]/NET0131 ,
		_w800_,
		_w824_
	);
	LUT2 #(
		.INIT('h8)
	) name293 (
		_w715_,
		_w763_,
		_w825_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w826_
	);
	LUT2 #(
		.INIT('h8)
	) name295 (
		_w694_,
		_w826_,
		_w827_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		\sa20_reg[2]/P0001 ,
		_w827_,
		_w828_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		_w723_,
		_w745_,
		_w829_
	);
	LUT2 #(
		.INIT('h2)
	) name298 (
		_w828_,
		_w829_,
		_w830_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		\sa20_reg[2]/P0001 ,
		_w715_,
		_w831_
	);
	LUT2 #(
		.INIT('h4)
	) name300 (
		\sa20_reg[5]/P0001 ,
		_w739_,
		_w832_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		\sa20_reg[3]/P0001 ,
		_w744_,
		_w833_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		\sa20_reg[6]/NET0131 ,
		_w833_,
		_w834_
	);
	LUT2 #(
		.INIT('h2)
	) name303 (
		_w831_,
		_w832_,
		_w835_
	);
	LUT2 #(
		.INIT('h4)
	) name304 (
		_w834_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		_w830_,
		_w836_,
		_w837_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		_w701_,
		_w799_,
		_w838_
	);
	LUT2 #(
		.INIT('h8)
	) name307 (
		_w705_,
		_w716_,
		_w839_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		_w838_,
		_w839_,
		_w840_
	);
	LUT2 #(
		.INIT('h4)
	) name309 (
		_w837_,
		_w840_,
		_w841_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		\sa20_reg[1]/P0001 ,
		_w841_,
		_w842_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		_w821_,
		_w824_,
		_w843_
	);
	LUT2 #(
		.INIT('h4)
	) name312 (
		_w825_,
		_w843_,
		_w844_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		_w818_,
		_w823_,
		_w845_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		_w844_,
		_w845_,
		_w846_
	);
	LUT2 #(
		.INIT('h4)
	) name315 (
		_w814_,
		_w846_,
		_w847_
	);
	LUT2 #(
		.INIT('h4)
	) name316 (
		_w842_,
		_w847_,
		_w848_
	);
	LUT2 #(
		.INIT('h4)
	) name317 (
		_w805_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h4)
	) name318 (
		_w760_,
		_w849_,
		_w850_
	);
	LUT2 #(
		.INIT('h2)
	) name319 (
		_w689_,
		_w850_,
		_w851_
	);
	LUT2 #(
		.INIT('h4)
	) name320 (
		_w689_,
		_w850_,
		_w852_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		_w851_,
		_w852_,
		_w853_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		_w550_,
		_w556_,
		_w854_
	);
	LUT2 #(
		.INIT('h4)
	) name323 (
		\sa13_reg[5]/P0001 ,
		_w583_,
		_w855_
	);
	LUT2 #(
		.INIT('h4)
	) name324 (
		\sa13_reg[3]/P0001 ,
		_w855_,
		_w856_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		\sa13_reg[7]/NET0131 ,
		_w608_,
		_w857_
	);
	LUT2 #(
		.INIT('h8)
	) name326 (
		\sa13_reg[5]/P0001 ,
		_w567_,
		_w858_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		_w560_,
		_w858_,
		_w859_
	);
	LUT2 #(
		.INIT('h2)
	) name328 (
		\sa13_reg[2]/P0001 ,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		\sa13_reg[5]/P0001 ,
		_w543_,
		_w861_
	);
	LUT2 #(
		.INIT('h4)
	) name330 (
		\sa13_reg[3]/P0001 ,
		_w861_,
		_w862_
	);
	LUT2 #(
		.INIT('h4)
	) name331 (
		\sa13_reg[4]/P0001 ,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		\sa13_reg[3]/P0001 ,
		_w549_,
		_w864_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		\sa13_reg[4]/P0001 ,
		_w543_,
		_w865_
	);
	LUT2 #(
		.INIT('h4)
	) name334 (
		\sa13_reg[3]/P0001 ,
		_w865_,
		_w866_
	);
	LUT2 #(
		.INIT('h1)
	) name335 (
		_w534_,
		_w864_,
		_w867_
	);
	LUT2 #(
		.INIT('h4)
	) name336 (
		_w866_,
		_w867_,
		_w868_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		\sa13_reg[2]/P0001 ,
		_w868_,
		_w869_
	);
	LUT2 #(
		.INIT('h1)
	) name338 (
		_w569_,
		_w854_,
		_w870_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		_w856_,
		_w857_,
		_w871_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		_w870_,
		_w871_,
		_w872_
	);
	LUT2 #(
		.INIT('h4)
	) name341 (
		_w863_,
		_w872_,
		_w873_
	);
	LUT2 #(
		.INIT('h1)
	) name342 (
		_w860_,
		_w869_,
		_w874_
	);
	LUT2 #(
		.INIT('h8)
	) name343 (
		_w873_,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h2)
	) name344 (
		\sa13_reg[1]/P0001 ,
		_w875_,
		_w876_
	);
	LUT2 #(
		.INIT('h4)
	) name345 (
		\sa13_reg[3]/P0001 ,
		_w591_,
		_w877_
	);
	LUT2 #(
		.INIT('h1)
	) name346 (
		_w604_,
		_w877_,
		_w878_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		_w653_,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w672_,
		_w857_,
		_w880_
	);
	LUT2 #(
		.INIT('h4)
	) name349 (
		_w879_,
		_w880_,
		_w881_
	);
	LUT2 #(
		.INIT('h2)
	) name350 (
		\sa13_reg[2]/P0001 ,
		_w881_,
		_w882_
	);
	LUT2 #(
		.INIT('h8)
	) name351 (
		\sa13_reg[2]/P0001 ,
		_w655_,
		_w883_
	);
	LUT2 #(
		.INIT('h8)
	) name352 (
		\sa13_reg[7]/NET0131 ,
		_w533_,
		_w884_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		_w883_,
		_w884_,
		_w885_
	);
	LUT2 #(
		.INIT('h2)
	) name354 (
		_w547_,
		_w885_,
		_w886_
	);
	LUT2 #(
		.INIT('h8)
	) name355 (
		\sa13_reg[2]/P0001 ,
		_w650_,
		_w887_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		_w559_,
		_w563_,
		_w888_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		_w887_,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h1)
	) name358 (
		\sa13_reg[3]/P0001 ,
		_w889_,
		_w890_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		_w886_,
		_w890_,
		_w891_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		\sa13_reg[1]/P0001 ,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h4)
	) name361 (
		\sa13_reg[2]/P0001 ,
		_w588_,
		_w893_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w548_,
		_w893_,
		_w894_
	);
	LUT2 #(
		.INIT('h8)
	) name363 (
		_w586_,
		_w894_,
		_w895_
	);
	LUT2 #(
		.INIT('h4)
	) name364 (
		_w882_,
		_w895_,
		_w896_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w892_,
		_w896_,
		_w897_
	);
	LUT2 #(
		.INIT('h4)
	) name366 (
		_w876_,
		_w897_,
		_w898_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		\sa13_reg[0]/P0001 ,
		_w898_,
		_w899_
	);
	LUT2 #(
		.INIT('h2)
	) name368 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w900_
	);
	LUT2 #(
		.INIT('h4)
	) name369 (
		\sa13_reg[4]/P0001 ,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h8)
	) name370 (
		\sa13_reg[3]/P0001 ,
		_w861_,
		_w902_
	);
	LUT2 #(
		.INIT('h4)
	) name371 (
		\sa13_reg[4]/P0001 ,
		_w544_,
		_w903_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		_w902_,
		_w903_,
		_w904_
	);
	LUT2 #(
		.INIT('h4)
	) name373 (
		_w901_,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('h1)
	) name374 (
		\sa13_reg[2]/P0001 ,
		_w905_,
		_w906_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		_w535_,
		_w587_,
		_w907_
	);
	LUT2 #(
		.INIT('h8)
	) name376 (
		_w563_,
		_w579_,
		_w908_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		_w907_,
		_w908_,
		_w909_
	);
	LUT2 #(
		.INIT('h2)
	) name378 (
		_w603_,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h8)
	) name379 (
		\sa13_reg[3]/P0001 ,
		_w537_,
		_w911_
	);
	LUT2 #(
		.INIT('h4)
	) name380 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w912_
	);
	LUT2 #(
		.INIT('h8)
	) name381 (
		_w587_,
		_w912_,
		_w913_
	);
	LUT2 #(
		.INIT('h4)
	) name382 (
		\sa13_reg[2]/P0001 ,
		_w913_,
		_w914_
	);
	LUT2 #(
		.INIT('h1)
	) name383 (
		_w580_,
		_w610_,
		_w915_
	);
	LUT2 #(
		.INIT('h4)
	) name384 (
		_w656_,
		_w915_,
		_w916_
	);
	LUT2 #(
		.INIT('h2)
	) name385 (
		_w680_,
		_w916_,
		_w917_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		\sa13_reg[3]/P0001 ,
		_w652_,
		_w918_
	);
	LUT2 #(
		.INIT('h4)
	) name387 (
		\sa13_reg[4]/P0001 ,
		_w864_,
		_w919_
	);
	LUT2 #(
		.INIT('h4)
	) name388 (
		\sa13_reg[3]/P0001 ,
		_w532_,
		_w920_
	);
	LUT2 #(
		.INIT('h8)
	) name389 (
		_w587_,
		_w920_,
		_w921_
	);
	LUT2 #(
		.INIT('h1)
	) name390 (
		_w558_,
		_w919_,
		_w922_
	);
	LUT2 #(
		.INIT('h4)
	) name391 (
		_w921_,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('h4)
	) name392 (
		_w918_,
		_w923_,
		_w924_
	);
	LUT2 #(
		.INIT('h2)
	) name393 (
		\sa13_reg[1]/P0001 ,
		_w924_,
		_w925_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		_w551_,
		_w861_,
		_w926_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		\sa13_reg[2]/P0001 ,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h4)
	) name396 (
		\sa13_reg[4]/P0001 ,
		_w912_,
		_w928_
	);
	LUT2 #(
		.INIT('h8)
	) name397 (
		_w555_,
		_w556_,
		_w929_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		_w928_,
		_w929_,
		_w930_
	);
	LUT2 #(
		.INIT('h2)
	) name399 (
		\sa13_reg[2]/P0001 ,
		_w930_,
		_w931_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		_w542_,
		_w902_,
		_w932_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		_w927_,
		_w931_,
		_w933_
	);
	LUT2 #(
		.INIT('h8)
	) name402 (
		_w932_,
		_w933_,
		_w934_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		\sa13_reg[1]/P0001 ,
		_w934_,
		_w935_
	);
	LUT2 #(
		.INIT('h1)
	) name404 (
		_w911_,
		_w914_,
		_w936_
	);
	LUT2 #(
		.INIT('h4)
	) name405 (
		_w910_,
		_w936_,
		_w937_
	);
	LUT2 #(
		.INIT('h4)
	) name406 (
		_w917_,
		_w937_,
		_w938_
	);
	LUT2 #(
		.INIT('h4)
	) name407 (
		_w906_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h4)
	) name408 (
		_w925_,
		_w939_,
		_w940_
	);
	LUT2 #(
		.INIT('h4)
	) name409 (
		_w935_,
		_w940_,
		_w941_
	);
	LUT2 #(
		.INIT('h2)
	) name410 (
		\sa13_reg[0]/P0001 ,
		_w941_,
		_w942_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		_w543_,
		_w549_,
		_w943_
	);
	LUT2 #(
		.INIT('h1)
	) name412 (
		\sa13_reg[5]/P0001 ,
		_w943_,
		_w944_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		_w533_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h4)
	) name414 (
		\sa13_reg[6]/NET0131 ,
		_w555_,
		_w946_
	);
	LUT2 #(
		.INIT('h8)
	) name415 (
		\sa13_reg[5]/P0001 ,
		_w946_,
		_w947_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		_w542_,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h4)
	) name417 (
		_w945_,
		_w948_,
		_w949_
	);
	LUT2 #(
		.INIT('h2)
	) name418 (
		\sa13_reg[2]/P0001 ,
		_w949_,
		_w950_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		_w654_,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		\sa13_reg[1]/P0001 ,
		_w951_,
		_w952_
	);
	LUT2 #(
		.INIT('h8)
	) name421 (
		\sa13_reg[4]/P0001 ,
		_w624_,
		_w953_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		_w603_,
		_w858_,
		_w954_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		\sa13_reg[3]/P0001 ,
		_w547_,
		_w955_
	);
	LUT2 #(
		.INIT('h8)
	) name424 (
		_w536_,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		_w893_,
		_w956_,
		_w957_
	);
	LUT2 #(
		.INIT('h4)
	) name426 (
		_w954_,
		_w957_,
		_w958_
	);
	LUT2 #(
		.INIT('h2)
	) name427 (
		\sa13_reg[1]/P0001 ,
		_w958_,
		_w959_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		_w681_,
		_w856_,
		_w960_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		\sa13_reg[2]/P0001 ,
		_w960_,
		_w961_
	);
	LUT2 #(
		.INIT('h1)
	) name430 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[2]/P0001 ,
		_w962_
	);
	LUT2 #(
		.INIT('h4)
	) name431 (
		\sa13_reg[3]/P0001 ,
		_w559_,
		_w963_
	);
	LUT2 #(
		.INIT('h4)
	) name432 (
		\sa13_reg[4]/P0001 ,
		_w963_,
		_w964_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		_w609_,
		_w913_,
		_w965_
	);
	LUT2 #(
		.INIT('h4)
	) name434 (
		_w964_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h2)
	) name435 (
		_w962_,
		_w966_,
		_w967_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		_w953_,
		_w961_,
		_w968_
	);
	LUT2 #(
		.INIT('h4)
	) name437 (
		_w959_,
		_w968_,
		_w969_
	);
	LUT2 #(
		.INIT('h4)
	) name438 (
		_w967_,
		_w969_,
		_w970_
	);
	LUT2 #(
		.INIT('h4)
	) name439 (
		_w952_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h4)
	) name440 (
		_w942_,
		_w971_,
		_w972_
	);
	LUT2 #(
		.INIT('h4)
	) name441 (
		_w899_,
		_w972_,
		_w973_
	);
	LUT2 #(
		.INIT('h1)
	) name442 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w974_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w975_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		\sa02_reg[7]/NET0131 ,
		_w975_,
		_w976_
	);
	LUT2 #(
		.INIT('h8)
	) name445 (
		_w974_,
		_w976_,
		_w977_
	);
	LUT2 #(
		.INIT('h2)
	) name446 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		_w978_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w979_
	);
	LUT2 #(
		.INIT('h4)
	) name448 (
		\sa02_reg[5]/P0001 ,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h8)
	) name449 (
		_w978_,
		_w980_,
		_w981_
	);
	LUT2 #(
		.INIT('h1)
	) name450 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w982_
	);
	LUT2 #(
		.INIT('h4)
	) name451 (
		\sa02_reg[4]/P0001 ,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h8)
	) name452 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		_w984_
	);
	LUT2 #(
		.INIT('h8)
	) name453 (
		_w983_,
		_w984_,
		_w985_
	);
	LUT2 #(
		.INIT('h4)
	) name454 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w986_
	);
	LUT2 #(
		.INIT('h8)
	) name455 (
		_w982_,
		_w986_,
		_w987_
	);
	LUT2 #(
		.INIT('h8)
	) name456 (
		\sa02_reg[7]/NET0131 ,
		_w987_,
		_w988_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		_w977_,
		_w981_,
		_w989_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		_w985_,
		_w988_,
		_w990_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		_w989_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		\sa02_reg[1]/P0001 ,
		_w991_,
		_w992_
	);
	LUT2 #(
		.INIT('h8)
	) name461 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w993_
	);
	LUT2 #(
		.INIT('h8)
	) name462 (
		\sa02_reg[4]/P0001 ,
		_w993_,
		_w994_
	);
	LUT2 #(
		.INIT('h1)
	) name463 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w995_
	);
	LUT2 #(
		.INIT('h4)
	) name464 (
		\sa02_reg[4]/P0001 ,
		_w995_,
		_w996_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		_w994_,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h2)
	) name466 (
		_w984_,
		_w997_,
		_w998_
	);
	LUT2 #(
		.INIT('h2)
	) name467 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w999_
	);
	LUT2 #(
		.INIT('h8)
	) name468 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w1000_
	);
	LUT2 #(
		.INIT('h8)
	) name469 (
		_w999_,
		_w1000_,
		_w1001_
	);
	LUT2 #(
		.INIT('h4)
	) name470 (
		\sa02_reg[2]/P0001 ,
		_w1001_,
		_w1002_
	);
	LUT2 #(
		.INIT('h4)
	) name471 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w1003_
	);
	LUT2 #(
		.INIT('h4)
	) name472 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w1004_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		_w1003_,
		_w1004_,
		_w1005_
	);
	LUT2 #(
		.INIT('h2)
	) name474 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w1006_
	);
	LUT2 #(
		.INIT('h4)
	) name475 (
		\sa02_reg[5]/P0001 ,
		_w1006_,
		_w1007_
	);
	LUT2 #(
		.INIT('h8)
	) name476 (
		\sa02_reg[3]/P0001 ,
		_w1007_,
		_w1008_
	);
	LUT2 #(
		.INIT('h1)
	) name477 (
		_w1005_,
		_w1008_,
		_w1009_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		\sa02_reg[2]/P0001 ,
		_w1009_,
		_w1010_
	);
	LUT2 #(
		.INIT('h4)
	) name479 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w1011_
	);
	LUT2 #(
		.INIT('h8)
	) name480 (
		_w986_,
		_w1011_,
		_w1012_
	);
	LUT2 #(
		.INIT('h8)
	) name481 (
		\sa02_reg[2]/P0001 ,
		_w1012_,
		_w1013_
	);
	LUT2 #(
		.INIT('h4)
	) name482 (
		\sa02_reg[7]/NET0131 ,
		_w1013_,
		_w1014_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w1015_
	);
	LUT2 #(
		.INIT('h2)
	) name484 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w1016_
	);
	LUT2 #(
		.INIT('h1)
	) name485 (
		_w982_,
		_w1016_,
		_w1017_
	);
	LUT2 #(
		.INIT('h2)
	) name486 (
		_w1015_,
		_w1017_,
		_w1018_
	);
	LUT2 #(
		.INIT('h8)
	) name487 (
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w1019_
	);
	LUT2 #(
		.INIT('h4)
	) name488 (
		\sa02_reg[5]/P0001 ,
		_w1019_,
		_w1020_
	);
	LUT2 #(
		.INIT('h4)
	) name489 (
		\sa02_reg[3]/P0001 ,
		_w1020_,
		_w1021_
	);
	LUT2 #(
		.INIT('h8)
	) name490 (
		_w986_,
		_w999_,
		_w1022_
	);
	LUT2 #(
		.INIT('h4)
	) name491 (
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w1023_
	);
	LUT2 #(
		.INIT('h8)
	) name492 (
		\sa02_reg[3]/P0001 ,
		_w1023_,
		_w1024_
	);
	LUT2 #(
		.INIT('h2)
	) name493 (
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w1025_
	);
	LUT2 #(
		.INIT('h8)
	) name494 (
		_w974_,
		_w1025_,
		_w1026_
	);
	LUT2 #(
		.INIT('h1)
	) name495 (
		\sa02_reg[2]/P0001 ,
		_w1022_,
		_w1027_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w1024_,
		_w1026_,
		_w1028_
	);
	LUT2 #(
		.INIT('h8)
	) name497 (
		_w1027_,
		_w1028_,
		_w1029_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		\sa02_reg[3]/P0001 ,
		_w993_,
		_w1030_
	);
	LUT2 #(
		.INIT('h8)
	) name499 (
		_w975_,
		_w1006_,
		_w1031_
	);
	LUT2 #(
		.INIT('h2)
	) name500 (
		\sa02_reg[2]/P0001 ,
		_w1030_,
		_w1032_
	);
	LUT2 #(
		.INIT('h4)
	) name501 (
		_w1031_,
		_w1032_,
		_w1033_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		_w1029_,
		_w1033_,
		_w1034_
	);
	LUT2 #(
		.INIT('h2)
	) name503 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		_w1035_
	);
	LUT2 #(
		.INIT('h4)
	) name504 (
		\sa02_reg[6]/NET0131 ,
		_w1035_,
		_w1036_
	);
	LUT2 #(
		.INIT('h4)
	) name505 (
		\sa02_reg[7]/NET0131 ,
		_w1036_,
		_w1037_
	);
	LUT2 #(
		.INIT('h8)
	) name506 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w1038_
	);
	LUT2 #(
		.INIT('h8)
	) name507 (
		\sa02_reg[7]/NET0131 ,
		_w1038_,
		_w1039_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		_w1026_,
		_w1039_,
		_w1040_
	);
	LUT2 #(
		.INIT('h2)
	) name509 (
		\sa02_reg[5]/P0001 ,
		_w1040_,
		_w1041_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		\sa02_reg[5]/P0001 ,
		_w1023_,
		_w1042_
	);
	LUT2 #(
		.INIT('h4)
	) name511 (
		\sa02_reg[4]/P0001 ,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		_w1021_,
		_w1037_,
		_w1044_
	);
	LUT2 #(
		.INIT('h4)
	) name513 (
		_w1043_,
		_w1044_,
		_w1045_
	);
	LUT2 #(
		.INIT('h4)
	) name514 (
		_w1041_,
		_w1045_,
		_w1046_
	);
	LUT2 #(
		.INIT('h4)
	) name515 (
		_w1034_,
		_w1046_,
		_w1047_
	);
	LUT2 #(
		.INIT('h2)
	) name516 (
		\sa02_reg[1]/P0001 ,
		_w1047_,
		_w1048_
	);
	LUT2 #(
		.INIT('h1)
	) name517 (
		_w1002_,
		_w1018_,
		_w1049_
	);
	LUT2 #(
		.INIT('h4)
	) name518 (
		_w998_,
		_w1049_,
		_w1050_
	);
	LUT2 #(
		.INIT('h4)
	) name519 (
		_w1014_,
		_w1050_,
		_w1051_
	);
	LUT2 #(
		.INIT('h4)
	) name520 (
		_w1010_,
		_w1051_,
		_w1052_
	);
	LUT2 #(
		.INIT('h4)
	) name521 (
		_w992_,
		_w1052_,
		_w1053_
	);
	LUT2 #(
		.INIT('h4)
	) name522 (
		_w1048_,
		_w1053_,
		_w1054_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		\sa02_reg[0]/P0001 ,
		_w1054_,
		_w1055_
	);
	LUT2 #(
		.INIT('h2)
	) name524 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w1056_
	);
	LUT2 #(
		.INIT('h8)
	) name525 (
		_w1038_,
		_w1056_,
		_w1057_
	);
	LUT2 #(
		.INIT('h4)
	) name526 (
		\sa02_reg[6]/NET0131 ,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h2)
	) name527 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w1059_
	);
	LUT2 #(
		.INIT('h8)
	) name528 (
		_w1023_,
		_w1059_,
		_w1060_
	);
	LUT2 #(
		.INIT('h4)
	) name529 (
		\sa02_reg[7]/NET0131 ,
		_w987_,
		_w1061_
	);
	LUT2 #(
		.INIT('h4)
	) name530 (
		\sa02_reg[3]/P0001 ,
		_w999_,
		_w1062_
	);
	LUT2 #(
		.INIT('h8)
	) name531 (
		_w1000_,
		_w1062_,
		_w1063_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w1058_,
		_w1060_,
		_w1064_
	);
	LUT2 #(
		.INIT('h1)
	) name533 (
		_w1061_,
		_w1063_,
		_w1065_
	);
	LUT2 #(
		.INIT('h8)
	) name534 (
		_w1064_,
		_w1065_,
		_w1066_
	);
	LUT2 #(
		.INIT('h2)
	) name535 (
		\sa02_reg[1]/P0001 ,
		_w1066_,
		_w1067_
	);
	LUT2 #(
		.INIT('h8)
	) name536 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w1068_
	);
	LUT2 #(
		.INIT('h8)
	) name537 (
		_w1015_,
		_w1068_,
		_w1069_
	);
	LUT2 #(
		.INIT('h8)
	) name538 (
		\sa02_reg[5]/P0001 ,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h8)
	) name539 (
		_w976_,
		_w986_,
		_w1071_
	);
	LUT2 #(
		.INIT('h8)
	) name540 (
		_w995_,
		_w1004_,
		_w1072_
	);
	LUT2 #(
		.INIT('h4)
	) name541 (
		\sa02_reg[3]/P0001 ,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h1)
	) name542 (
		_w1071_,
		_w1073_,
		_w1074_
	);
	LUT2 #(
		.INIT('h2)
	) name543 (
		\sa02_reg[2]/P0001 ,
		_w1074_,
		_w1075_
	);
	LUT2 #(
		.INIT('h8)
	) name544 (
		_w1000_,
		_w1011_,
		_w1076_
	);
	LUT2 #(
		.INIT('h4)
	) name545 (
		\sa02_reg[2]/P0001 ,
		_w1076_,
		_w1077_
	);
	LUT2 #(
		.INIT('h8)
	) name546 (
		\sa02_reg[5]/P0001 ,
		_w1059_,
		_w1078_
	);
	LUT2 #(
		.INIT('h1)
	) name547 (
		_w983_,
		_w1007_,
		_w1079_
	);
	LUT2 #(
		.INIT('h4)
	) name548 (
		_w1078_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h2)
	) name549 (
		\sa02_reg[1]/P0001 ,
		_w1080_,
		_w1081_
	);
	LUT2 #(
		.INIT('h8)
	) name550 (
		_w1056_,
		_w1068_,
		_w1082_
	);
	LUT2 #(
		.INIT('h1)
	) name551 (
		_w1069_,
		_w1082_,
		_w1083_
	);
	LUT2 #(
		.INIT('h4)
	) name552 (
		\sa02_reg[4]/P0001 ,
		_w1056_,
		_w1084_
	);
	LUT2 #(
		.INIT('h2)
	) name553 (
		_w1083_,
		_w1084_,
		_w1085_
	);
	LUT2 #(
		.INIT('h4)
	) name554 (
		_w1081_,
		_w1085_,
		_w1086_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		\sa02_reg[2]/P0001 ,
		_w1086_,
		_w1087_
	);
	LUT2 #(
		.INIT('h8)
	) name556 (
		\sa02_reg[5]/P0001 ,
		_w1025_,
		_w1088_
	);
	LUT2 #(
		.INIT('h4)
	) name557 (
		_w978_,
		_w1088_,
		_w1089_
	);
	LUT2 #(
		.INIT('h4)
	) name558 (
		\sa02_reg[4]/P0001 ,
		_w1011_,
		_w1090_
	);
	LUT2 #(
		.INIT('h8)
	) name559 (
		_w979_,
		_w1038_,
		_w1091_
	);
	LUT2 #(
		.INIT('h1)
	) name560 (
		_w1090_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h2)
	) name561 (
		\sa02_reg[2]/P0001 ,
		_w1092_,
		_w1093_
	);
	LUT2 #(
		.INIT('h4)
	) name562 (
		\sa02_reg[5]/P0001 ,
		_w1023_,
		_w1094_
	);
	LUT2 #(
		.INIT('h4)
	) name563 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		_w1095_
	);
	LUT2 #(
		.INIT('h8)
	) name564 (
		_w1094_,
		_w1095_,
		_w1096_
	);
	LUT2 #(
		.INIT('h1)
	) name565 (
		_w1071_,
		_w1089_,
		_w1097_
	);
	LUT2 #(
		.INIT('h4)
	) name566 (
		_w1096_,
		_w1097_,
		_w1098_
	);
	LUT2 #(
		.INIT('h4)
	) name567 (
		_w1093_,
		_w1098_,
		_w1099_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		\sa02_reg[1]/P0001 ,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h1)
	) name569 (
		_w1070_,
		_w1077_,
		_w1101_
	);
	LUT2 #(
		.INIT('h4)
	) name570 (
		_w1075_,
		_w1101_,
		_w1102_
	);
	LUT2 #(
		.INIT('h4)
	) name571 (
		_w1067_,
		_w1102_,
		_w1103_
	);
	LUT2 #(
		.INIT('h4)
	) name572 (
		_w1087_,
		_w1103_,
		_w1104_
	);
	LUT2 #(
		.INIT('h4)
	) name573 (
		_w1100_,
		_w1104_,
		_w1105_
	);
	LUT2 #(
		.INIT('h2)
	) name574 (
		\sa02_reg[0]/P0001 ,
		_w1105_,
		_w1106_
	);
	LUT2 #(
		.INIT('h2)
	) name575 (
		\sa02_reg[2]/P0001 ,
		_w1058_,
		_w1107_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		\sa02_reg[2]/P0001 ,
		_w1021_,
		_w1108_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		\sa02_reg[6]/NET0131 ,
		_w1059_,
		_w1109_
	);
	LUT2 #(
		.INIT('h8)
	) name578 (
		_w1056_,
		_w1109_,
		_w1110_
	);
	LUT2 #(
		.INIT('h2)
	) name579 (
		_w1108_,
		_w1110_,
		_w1111_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		_w1107_,
		_w1111_,
		_w1112_
	);
	LUT2 #(
		.INIT('h8)
	) name581 (
		_w978_,
		_w1025_,
		_w1113_
	);
	LUT2 #(
		.INIT('h8)
	) name582 (
		\sa02_reg[4]/P0001 ,
		_w1113_,
		_w1114_
	);
	LUT2 #(
		.INIT('h8)
	) name583 (
		\sa02_reg[5]/P0001 ,
		_w1114_,
		_w1115_
	);
	LUT2 #(
		.INIT('h8)
	) name584 (
		_w979_,
		_w1059_,
		_w1116_
	);
	LUT2 #(
		.INIT('h4)
	) name585 (
		\sa02_reg[5]/P0001 ,
		_w1116_,
		_w1117_
	);
	LUT2 #(
		.INIT('h1)
	) name586 (
		_w1002_,
		_w1117_,
		_w1118_
	);
	LUT2 #(
		.INIT('h4)
	) name587 (
		_w1115_,
		_w1118_,
		_w1119_
	);
	LUT2 #(
		.INIT('h2)
	) name588 (
		\sa02_reg[1]/P0001 ,
		_w1119_,
		_w1120_
	);
	LUT2 #(
		.INIT('h8)
	) name589 (
		_w974_,
		_w979_,
		_w1121_
	);
	LUT2 #(
		.INIT('h8)
	) name590 (
		\sa02_reg[7]/NET0131 ,
		_w974_,
		_w1122_
	);
	LUT2 #(
		.INIT('h8)
	) name591 (
		_w1025_,
		_w1038_,
		_w1123_
	);
	LUT2 #(
		.INIT('h1)
	) name592 (
		_w1122_,
		_w1123_,
		_w1124_
	);
	LUT2 #(
		.INIT('h2)
	) name593 (
		\sa02_reg[5]/P0001 ,
		_w1124_,
		_w1125_
	);
	LUT2 #(
		.INIT('h1)
	) name594 (
		_w1076_,
		_w1125_,
		_w1126_
	);
	LUT2 #(
		.INIT('h1)
	) name595 (
		\sa02_reg[2]/P0001 ,
		_w1126_,
		_w1127_
	);
	LUT2 #(
		.INIT('h8)
	) name596 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w1128_
	);
	LUT2 #(
		.INIT('h2)
	) name597 (
		\sa02_reg[3]/P0001 ,
		_w999_,
		_w1129_
	);
	LUT2 #(
		.INIT('h4)
	) name598 (
		\sa02_reg[5]/P0001 ,
		_w1025_,
		_w1130_
	);
	LUT2 #(
		.INIT('h1)
	) name599 (
		_w1094_,
		_w1130_,
		_w1131_
	);
	LUT2 #(
		.INIT('h1)
	) name600 (
		\sa02_reg[3]/P0001 ,
		_w976_,
		_w1132_
	);
	LUT2 #(
		.INIT('h8)
	) name601 (
		_w1131_,
		_w1132_,
		_w1133_
	);
	LUT2 #(
		.INIT('h2)
	) name602 (
		_w1128_,
		_w1129_,
		_w1134_
	);
	LUT2 #(
		.INIT('h4)
	) name603 (
		_w1133_,
		_w1134_,
		_w1135_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		_w1121_,
		_w1135_,
		_w1136_
	);
	LUT2 #(
		.INIT('h4)
	) name605 (
		_w1127_,
		_w1136_,
		_w1137_
	);
	LUT2 #(
		.INIT('h1)
	) name606 (
		\sa02_reg[1]/P0001 ,
		_w1137_,
		_w1138_
	);
	LUT2 #(
		.INIT('h1)
	) name607 (
		_w1112_,
		_w1120_,
		_w1139_
	);
	LUT2 #(
		.INIT('h4)
	) name608 (
		_w1138_,
		_w1139_,
		_w1140_
	);
	LUT2 #(
		.INIT('h4)
	) name609 (
		_w1055_,
		_w1140_,
		_w1141_
	);
	LUT2 #(
		.INIT('h4)
	) name610 (
		_w1106_,
		_w1141_,
		_w1142_
	);
	LUT2 #(
		.INIT('h1)
	) name611 (
		_w973_,
		_w1142_,
		_w1143_
	);
	LUT2 #(
		.INIT('h8)
	) name612 (
		_w973_,
		_w1142_,
		_w1144_
	);
	LUT2 #(
		.INIT('h1)
	) name613 (
		_w1143_,
		_w1144_,
		_w1145_
	);
	LUT2 #(
		.INIT('h4)
	) name614 (
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w1146_
	);
	LUT2 #(
		.INIT('h8)
	) name615 (
		\sa31_reg[5]/P0001 ,
		_w1146_,
		_w1147_
	);
	LUT2 #(
		.INIT('h4)
	) name616 (
		\sa31_reg[4]/P0001 ,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h2)
	) name617 (
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w1149_
	);
	LUT2 #(
		.INIT('h8)
	) name618 (
		\sa31_reg[4]/P0001 ,
		_w1149_,
		_w1150_
	);
	LUT2 #(
		.INIT('h4)
	) name619 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w1151_
	);
	LUT2 #(
		.INIT('h1)
	) name620 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w1152_
	);
	LUT2 #(
		.INIT('h8)
	) name621 (
		\sa31_reg[7]/P0001 ,
		_w1152_,
		_w1153_
	);
	LUT2 #(
		.INIT('h8)
	) name622 (
		_w1151_,
		_w1153_,
		_w1154_
	);
	LUT2 #(
		.INIT('h1)
	) name623 (
		_w1148_,
		_w1150_,
		_w1155_
	);
	LUT2 #(
		.INIT('h4)
	) name624 (
		_w1154_,
		_w1155_,
		_w1156_
	);
	LUT2 #(
		.INIT('h2)
	) name625 (
		\sa31_reg[2]/P0001 ,
		_w1156_,
		_w1157_
	);
	LUT2 #(
		.INIT('h2)
	) name626 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w1158_
	);
	LUT2 #(
		.INIT('h8)
	) name627 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w1159_
	);
	LUT2 #(
		.INIT('h4)
	) name628 (
		\sa31_reg[6]/NET0131 ,
		_w1159_,
		_w1160_
	);
	LUT2 #(
		.INIT('h8)
	) name629 (
		_w1158_,
		_w1160_,
		_w1161_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		_w1162_
	);
	LUT2 #(
		.INIT('h4)
	) name631 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w1163_
	);
	LUT2 #(
		.INIT('h1)
	) name632 (
		\sa31_reg[5]/P0001 ,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h8)
	) name633 (
		_w1162_,
		_w1164_,
		_w1165_
	);
	LUT2 #(
		.INIT('h8)
	) name634 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w1166_
	);
	LUT2 #(
		.INIT('h8)
	) name635 (
		\sa31_reg[3]/P0001 ,
		_w1166_,
		_w1167_
	);
	LUT2 #(
		.INIT('h4)
	) name636 (
		\sa31_reg[4]/P0001 ,
		_w1167_,
		_w1168_
	);
	LUT2 #(
		.INIT('h1)
	) name637 (
		_w1161_,
		_w1165_,
		_w1169_
	);
	LUT2 #(
		.INIT('h4)
	) name638 (
		_w1168_,
		_w1169_,
		_w1170_
	);
	LUT2 #(
		.INIT('h4)
	) name639 (
		_w1157_,
		_w1170_,
		_w1171_
	);
	LUT2 #(
		.INIT('h2)
	) name640 (
		\sa31_reg[1]/P0001 ,
		_w1171_,
		_w1172_
	);
	LUT2 #(
		.INIT('h4)
	) name641 (
		\sa31_reg[5]/P0001 ,
		_w1149_,
		_w1173_
	);
	LUT2 #(
		.INIT('h8)
	) name642 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w1174_
	);
	LUT2 #(
		.INIT('h8)
	) name643 (
		\sa31_reg[3]/P0001 ,
		_w1174_,
		_w1175_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		_w1173_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h2)
	) name645 (
		\sa31_reg[2]/P0001 ,
		_w1176_,
		_w1177_
	);
	LUT2 #(
		.INIT('h2)
	) name646 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w1178_
	);
	LUT2 #(
		.INIT('h8)
	) name647 (
		_w1174_,
		_w1178_,
		_w1179_
	);
	LUT2 #(
		.INIT('h1)
	) name648 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w1180_
	);
	LUT2 #(
		.INIT('h8)
	) name649 (
		_w1159_,
		_w1180_,
		_w1181_
	);
	LUT2 #(
		.INIT('h4)
	) name650 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w1182_
	);
	LUT2 #(
		.INIT('h8)
	) name651 (
		_w1163_,
		_w1182_,
		_w1183_
	);
	LUT2 #(
		.INIT('h1)
	) name652 (
		_w1181_,
		_w1183_,
		_w1184_
	);
	LUT2 #(
		.INIT('h1)
	) name653 (
		\sa31_reg[2]/P0001 ,
		_w1184_,
		_w1185_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w1186_
	);
	LUT2 #(
		.INIT('h8)
	) name655 (
		\sa31_reg[5]/P0001 ,
		_w1186_,
		_w1187_
	);
	LUT2 #(
		.INIT('h8)
	) name656 (
		_w1162_,
		_w1187_,
		_w1188_
	);
	LUT2 #(
		.INIT('h1)
	) name657 (
		_w1179_,
		_w1188_,
		_w1189_
	);
	LUT2 #(
		.INIT('h4)
	) name658 (
		_w1177_,
		_w1189_,
		_w1190_
	);
	LUT2 #(
		.INIT('h4)
	) name659 (
		_w1185_,
		_w1190_,
		_w1191_
	);
	LUT2 #(
		.INIT('h1)
	) name660 (
		\sa31_reg[1]/P0001 ,
		_w1191_,
		_w1192_
	);
	LUT2 #(
		.INIT('h8)
	) name661 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w1193_
	);
	LUT2 #(
		.INIT('h4)
	) name662 (
		\sa31_reg[7]/P0001 ,
		_w1193_,
		_w1194_
	);
	LUT2 #(
		.INIT('h4)
	) name663 (
		\sa31_reg[4]/P0001 ,
		_w1194_,
		_w1195_
	);
	LUT2 #(
		.INIT('h4)
	) name664 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w1196_
	);
	LUT2 #(
		.INIT('h8)
	) name665 (
		_w1178_,
		_w1196_,
		_w1197_
	);
	LUT2 #(
		.INIT('h1)
	) name666 (
		_w1195_,
		_w1197_,
		_w1198_
	);
	LUT2 #(
		.INIT('h1)
	) name667 (
		\sa31_reg[2]/P0001 ,
		_w1198_,
		_w1199_
	);
	LUT2 #(
		.INIT('h8)
	) name668 (
		\sa31_reg[3]/P0001 ,
		_w1150_,
		_w1200_
	);
	LUT2 #(
		.INIT('h8)
	) name669 (
		\sa31_reg[6]/NET0131 ,
		_w1166_,
		_w1201_
	);
	LUT2 #(
		.INIT('h8)
	) name670 (
		_w1196_,
		_w1201_,
		_w1202_
	);
	LUT2 #(
		.INIT('h1)
	) name671 (
		_w1200_,
		_w1202_,
		_w1203_
	);
	LUT2 #(
		.INIT('h4)
	) name672 (
		\sa31_reg[4]/P0001 ,
		_w1180_,
		_w1204_
	);
	LUT2 #(
		.INIT('h4)
	) name673 (
		\sa31_reg[6]/NET0131 ,
		_w1204_,
		_w1205_
	);
	LUT2 #(
		.INIT('h8)
	) name674 (
		\sa31_reg[3]/P0001 ,
		_w1146_,
		_w1206_
	);
	LUT2 #(
		.INIT('h4)
	) name675 (
		\sa31_reg[5]/P0001 ,
		_w1206_,
		_w1207_
	);
	LUT2 #(
		.INIT('h1)
	) name676 (
		_w1205_,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h8)
	) name677 (
		_w1203_,
		_w1208_,
		_w1209_
	);
	LUT2 #(
		.INIT('h2)
	) name678 (
		\sa31_reg[2]/P0001 ,
		_w1209_,
		_w1210_
	);
	LUT2 #(
		.INIT('h1)
	) name679 (
		_w1199_,
		_w1210_,
		_w1211_
	);
	LUT2 #(
		.INIT('h4)
	) name680 (
		_w1192_,
		_w1211_,
		_w1212_
	);
	LUT2 #(
		.INIT('h4)
	) name681 (
		_w1172_,
		_w1212_,
		_w1213_
	);
	LUT2 #(
		.INIT('h2)
	) name682 (
		\sa31_reg[0]/P0002 ,
		_w1213_,
		_w1214_
	);
	LUT2 #(
		.INIT('h8)
	) name683 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w1215_
	);
	LUT2 #(
		.INIT('h2)
	) name684 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		_w1216_
	);
	LUT2 #(
		.INIT('h8)
	) name685 (
		_w1149_,
		_w1216_,
		_w1217_
	);
	LUT2 #(
		.INIT('h8)
	) name686 (
		_w1215_,
		_w1217_,
		_w1218_
	);
	LUT2 #(
		.INIT('h4)
	) name687 (
		\sa31_reg[5]/P0001 ,
		_w1186_,
		_w1219_
	);
	LUT2 #(
		.INIT('h4)
	) name688 (
		\sa31_reg[3]/P0001 ,
		_w1219_,
		_w1220_
	);
	LUT2 #(
		.INIT('h8)
	) name689 (
		\sa31_reg[2]/P0001 ,
		_w1220_,
		_w1221_
	);
	LUT2 #(
		.INIT('h4)
	) name690 (
		\sa31_reg[2]/P0001 ,
		_w1175_,
		_w1222_
	);
	LUT2 #(
		.INIT('h8)
	) name691 (
		_w1178_,
		_w1222_,
		_w1223_
	);
	LUT2 #(
		.INIT('h2)
	) name692 (
		\sa31_reg[1]/P0001 ,
		\sa31_reg[2]/P0001 ,
		_w1224_
	);
	LUT2 #(
		.INIT('h2)
	) name693 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w1225_
	);
	LUT2 #(
		.INIT('h4)
	) name694 (
		\sa31_reg[6]/NET0131 ,
		_w1225_,
		_w1226_
	);
	LUT2 #(
		.INIT('h8)
	) name695 (
		_w1158_,
		_w1226_,
		_w1227_
	);
	LUT2 #(
		.INIT('h8)
	) name696 (
		_w1224_,
		_w1227_,
		_w1228_
	);
	LUT2 #(
		.INIT('h1)
	) name697 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w1229_
	);
	LUT2 #(
		.INIT('h4)
	) name698 (
		\sa31_reg[7]/P0001 ,
		_w1152_,
		_w1230_
	);
	LUT2 #(
		.INIT('h8)
	) name699 (
		_w1229_,
		_w1230_,
		_w1231_
	);
	LUT2 #(
		.INIT('h8)
	) name700 (
		\sa31_reg[1]/P0001 ,
		\sa31_reg[2]/P0001 ,
		_w1232_
	);
	LUT2 #(
		.INIT('h8)
	) name701 (
		\sa31_reg[4]/P0001 ,
		_w1219_,
		_w1233_
	);
	LUT2 #(
		.INIT('h8)
	) name702 (
		_w1152_,
		_w1186_,
		_w1234_
	);
	LUT2 #(
		.INIT('h8)
	) name703 (
		\sa31_reg[3]/P0001 ,
		_w1148_,
		_w1235_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		_w1233_,
		_w1234_,
		_w1236_
	);
	LUT2 #(
		.INIT('h4)
	) name705 (
		_w1235_,
		_w1236_,
		_w1237_
	);
	LUT2 #(
		.INIT('h2)
	) name706 (
		_w1232_,
		_w1237_,
		_w1238_
	);
	LUT2 #(
		.INIT('h4)
	) name707 (
		\sa31_reg[5]/P0001 ,
		_w1150_,
		_w1239_
	);
	LUT2 #(
		.INIT('h8)
	) name708 (
		\sa31_reg[5]/P0001 ,
		_w1206_,
		_w1240_
	);
	LUT2 #(
		.INIT('h1)
	) name709 (
		_w1179_,
		_w1239_,
		_w1241_
	);
	LUT2 #(
		.INIT('h4)
	) name710 (
		_w1240_,
		_w1241_,
		_w1242_
	);
	LUT2 #(
		.INIT('h1)
	) name711 (
		\sa31_reg[2]/P0001 ,
		_w1242_,
		_w1243_
	);
	LUT2 #(
		.INIT('h2)
	) name712 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w1244_
	);
	LUT2 #(
		.INIT('h8)
	) name713 (
		_w1201_,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('h8)
	) name714 (
		_w1146_,
		_w1159_,
		_w1246_
	);
	LUT2 #(
		.INIT('h8)
	) name715 (
		_w1152_,
		_w1193_,
		_w1247_
	);
	LUT2 #(
		.INIT('h8)
	) name716 (
		\sa31_reg[3]/P0001 ,
		_w1244_,
		_w1248_
	);
	LUT2 #(
		.INIT('h8)
	) name717 (
		_w1186_,
		_w1248_,
		_w1249_
	);
	LUT2 #(
		.INIT('h1)
	) name718 (
		_w1246_,
		_w1247_,
		_w1250_
	);
	LUT2 #(
		.INIT('h4)
	) name719 (
		_w1245_,
		_w1250_,
		_w1251_
	);
	LUT2 #(
		.INIT('h4)
	) name720 (
		_w1249_,
		_w1251_,
		_w1252_
	);
	LUT2 #(
		.INIT('h4)
	) name721 (
		_w1243_,
		_w1252_,
		_w1253_
	);
	LUT2 #(
		.INIT('h1)
	) name722 (
		\sa31_reg[1]/P0001 ,
		_w1253_,
		_w1254_
	);
	LUT2 #(
		.INIT('h8)
	) name723 (
		_w1196_,
		_w1229_,
		_w1255_
	);
	LUT2 #(
		.INIT('h8)
	) name724 (
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w1256_
	);
	LUT2 #(
		.INIT('h2)
	) name725 (
		\sa31_reg[4]/P0001 ,
		_w1256_,
		_w1257_
	);
	LUT2 #(
		.INIT('h4)
	) name726 (
		_w1186_,
		_w1216_,
		_w1258_
	);
	LUT2 #(
		.INIT('h4)
	) name727 (
		_w1257_,
		_w1258_,
		_w1259_
	);
	LUT2 #(
		.INIT('h8)
	) name728 (
		\sa31_reg[6]/NET0131 ,
		_w1196_,
		_w1260_
	);
	LUT2 #(
		.INIT('h8)
	) name729 (
		_w1158_,
		_w1260_,
		_w1261_
	);
	LUT2 #(
		.INIT('h1)
	) name730 (
		_w1255_,
		_w1259_,
		_w1262_
	);
	LUT2 #(
		.INIT('h4)
	) name731 (
		_w1261_,
		_w1262_,
		_w1263_
	);
	LUT2 #(
		.INIT('h1)
	) name732 (
		\sa31_reg[2]/P0001 ,
		_w1263_,
		_w1264_
	);
	LUT2 #(
		.INIT('h8)
	) name733 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		_w1265_
	);
	LUT2 #(
		.INIT('h8)
	) name734 (
		_w1187_,
		_w1265_,
		_w1266_
	);
	LUT2 #(
		.INIT('h1)
	) name735 (
		_w1225_,
		_w1260_,
		_w1267_
	);
	LUT2 #(
		.INIT('h2)
	) name736 (
		_w1182_,
		_w1267_,
		_w1268_
	);
	LUT2 #(
		.INIT('h4)
	) name737 (
		\sa31_reg[3]/P0001 ,
		_w1146_,
		_w1269_
	);
	LUT2 #(
		.INIT('h1)
	) name738 (
		_w1194_,
		_w1269_,
		_w1270_
	);
	LUT2 #(
		.INIT('h1)
	) name739 (
		\sa31_reg[4]/P0001 ,
		_w1270_,
		_w1271_
	);
	LUT2 #(
		.INIT('h1)
	) name740 (
		\sa31_reg[1]/P0001 ,
		_w1222_,
		_w1272_
	);
	LUT2 #(
		.INIT('h4)
	) name741 (
		_w1266_,
		_w1272_,
		_w1273_
	);
	LUT2 #(
		.INIT('h1)
	) name742 (
		_w1268_,
		_w1271_,
		_w1274_
	);
	LUT2 #(
		.INIT('h8)
	) name743 (
		_w1273_,
		_w1274_,
		_w1275_
	);
	LUT2 #(
		.INIT('h2)
	) name744 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w1276_
	);
	LUT2 #(
		.INIT('h8)
	) name745 (
		\sa31_reg[4]/P0001 ,
		_w1193_,
		_w1277_
	);
	LUT2 #(
		.INIT('h8)
	) name746 (
		_w1276_,
		_w1277_,
		_w1278_
	);
	LUT2 #(
		.INIT('h2)
	) name747 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		_w1279_
	);
	LUT2 #(
		.INIT('h8)
	) name748 (
		\sa31_reg[4]/P0001 ,
		_w1166_,
		_w1280_
	);
	LUT2 #(
		.INIT('h1)
	) name749 (
		_w1204_,
		_w1280_,
		_w1281_
	);
	LUT2 #(
		.INIT('h2)
	) name750 (
		_w1279_,
		_w1281_,
		_w1282_
	);
	LUT2 #(
		.INIT('h4)
	) name751 (
		\sa31_reg[2]/P0001 ,
		_w1205_,
		_w1283_
	);
	LUT2 #(
		.INIT('h2)
	) name752 (
		\sa31_reg[1]/P0001 ,
		_w1278_,
		_w1284_
	);
	LUT2 #(
		.INIT('h4)
	) name753 (
		_w1282_,
		_w1284_,
		_w1285_
	);
	LUT2 #(
		.INIT('h4)
	) name754 (
		_w1283_,
		_w1285_,
		_w1286_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		_w1275_,
		_w1286_,
		_w1287_
	);
	LUT2 #(
		.INIT('h8)
	) name756 (
		_w1164_,
		_w1279_,
		_w1288_
	);
	LUT2 #(
		.INIT('h4)
	) name757 (
		_w1257_,
		_w1288_,
		_w1289_
	);
	LUT2 #(
		.INIT('h1)
	) name758 (
		_w1264_,
		_w1289_,
		_w1290_
	);
	LUT2 #(
		.INIT('h4)
	) name759 (
		_w1287_,
		_w1290_,
		_w1291_
	);
	LUT2 #(
		.INIT('h1)
	) name760 (
		\sa31_reg[0]/P0002 ,
		_w1291_,
		_w1292_
	);
	LUT2 #(
		.INIT('h1)
	) name761 (
		_w1218_,
		_w1231_,
		_w1293_
	);
	LUT2 #(
		.INIT('h4)
	) name762 (
		_w1221_,
		_w1293_,
		_w1294_
	);
	LUT2 #(
		.INIT('h1)
	) name763 (
		_w1223_,
		_w1228_,
		_w1295_
	);
	LUT2 #(
		.INIT('h8)
	) name764 (
		_w1294_,
		_w1295_,
		_w1296_
	);
	LUT2 #(
		.INIT('h4)
	) name765 (
		_w1238_,
		_w1296_,
		_w1297_
	);
	LUT2 #(
		.INIT('h4)
	) name766 (
		_w1254_,
		_w1297_,
		_w1298_
	);
	LUT2 #(
		.INIT('h4)
	) name767 (
		_w1292_,
		_w1298_,
		_w1299_
	);
	LUT2 #(
		.INIT('h4)
	) name768 (
		_w1214_,
		_w1299_,
		_w1300_
	);
	LUT2 #(
		.INIT('h2)
	) name769 (
		\u0_w_reg[2][30]/P0001 ,
		_w1300_,
		_w1301_
	);
	LUT2 #(
		.INIT('h4)
	) name770 (
		\u0_w_reg[2][30]/P0001 ,
		_w1300_,
		_w1302_
	);
	LUT2 #(
		.INIT('h1)
	) name771 (
		_w1301_,
		_w1302_,
		_w1303_
	);
	LUT2 #(
		.INIT('h8)
	) name772 (
		_w1145_,
		_w1303_,
		_w1304_
	);
	LUT2 #(
		.INIT('h1)
	) name773 (
		_w1145_,
		_w1303_,
		_w1305_
	);
	LUT2 #(
		.INIT('h1)
	) name774 (
		_w1304_,
		_w1305_,
		_w1306_
	);
	LUT2 #(
		.INIT('h1)
	) name775 (
		_w853_,
		_w1306_,
		_w1307_
	);
	LUT2 #(
		.INIT('h8)
	) name776 (
		_w853_,
		_w1306_,
		_w1308_
	);
	LUT2 #(
		.INIT('h1)
	) name777 (
		\ld_r_reg/P0001 ,
		_w1307_,
		_w1309_
	);
	LUT2 #(
		.INIT('h4)
	) name778 (
		_w1308_,
		_w1309_,
		_w1310_
	);
	LUT2 #(
		.INIT('h2)
	) name779 (
		\text_in_r_reg[62]/P0001 ,
		\u0_w_reg[2][30]/P0001 ,
		_w1311_
	);
	LUT2 #(
		.INIT('h4)
	) name780 (
		\text_in_r_reg[62]/P0001 ,
		\u0_w_reg[2][30]/P0001 ,
		_w1312_
	);
	LUT2 #(
		.INIT('h2)
	) name781 (
		\ld_r_reg/P0001 ,
		_w1311_,
		_w1313_
	);
	LUT2 #(
		.INIT('h4)
	) name782 (
		_w1312_,
		_w1313_,
		_w1314_
	);
	LUT2 #(
		.INIT('h1)
	) name783 (
		_w1310_,
		_w1314_,
		_w1315_
	);
	LUT2 #(
		.INIT('h8)
	) name784 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1316_
	);
	LUT2 #(
		.INIT('h8)
	) name785 (
		\sa03_reg[7]/NET0131 ,
		_w1316_,
		_w1317_
	);
	LUT2 #(
		.INIT('h2)
	) name786 (
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1318_
	);
	LUT2 #(
		.INIT('h4)
	) name787 (
		\sa03_reg[4]/P0001 ,
		_w1318_,
		_w1319_
	);
	LUT2 #(
		.INIT('h4)
	) name788 (
		\sa03_reg[3]/P0001 ,
		_w1319_,
		_w1320_
	);
	LUT2 #(
		.INIT('h1)
	) name789 (
		_w1317_,
		_w1320_,
		_w1321_
	);
	LUT2 #(
		.INIT('h2)
	) name790 (
		\sa03_reg[5]/P0001 ,
		_w1321_,
		_w1322_
	);
	LUT2 #(
		.INIT('h1)
	) name791 (
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1323_
	);
	LUT2 #(
		.INIT('h2)
	) name792 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		_w1324_
	);
	LUT2 #(
		.INIT('h8)
	) name793 (
		_w1323_,
		_w1324_,
		_w1325_
	);
	LUT2 #(
		.INIT('h4)
	) name794 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1326_
	);
	LUT2 #(
		.INIT('h4)
	) name795 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1327_
	);
	LUT2 #(
		.INIT('h8)
	) name796 (
		_w1326_,
		_w1327_,
		_w1328_
	);
	LUT2 #(
		.INIT('h2)
	) name797 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1329_
	);
	LUT2 #(
		.INIT('h4)
	) name798 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1330_
	);
	LUT2 #(
		.INIT('h8)
	) name799 (
		_w1329_,
		_w1330_,
		_w1331_
	);
	LUT2 #(
		.INIT('h4)
	) name800 (
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1332_
	);
	LUT2 #(
		.INIT('h8)
	) name801 (
		\sa03_reg[3]/P0001 ,
		_w1332_,
		_w1333_
	);
	LUT2 #(
		.INIT('h4)
	) name802 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1334_
	);
	LUT2 #(
		.INIT('h8)
	) name803 (
		_w1329_,
		_w1334_,
		_w1335_
	);
	LUT2 #(
		.INIT('h1)
	) name804 (
		\sa03_reg[2]/P0001 ,
		_w1333_,
		_w1336_
	);
	LUT2 #(
		.INIT('h4)
	) name805 (
		_w1335_,
		_w1336_,
		_w1337_
	);
	LUT2 #(
		.INIT('h4)
	) name806 (
		_w1320_,
		_w1337_,
		_w1338_
	);
	LUT2 #(
		.INIT('h8)
	) name807 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1339_
	);
	LUT2 #(
		.INIT('h8)
	) name808 (
		\sa03_reg[3]/P0001 ,
		_w1339_,
		_w1340_
	);
	LUT2 #(
		.INIT('h2)
	) name809 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1341_
	);
	LUT2 #(
		.INIT('h8)
	) name810 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1342_
	);
	LUT2 #(
		.INIT('h8)
	) name811 (
		_w1341_,
		_w1342_,
		_w1343_
	);
	LUT2 #(
		.INIT('h2)
	) name812 (
		\sa03_reg[2]/P0001 ,
		_w1340_,
		_w1344_
	);
	LUT2 #(
		.INIT('h4)
	) name813 (
		_w1343_,
		_w1344_,
		_w1345_
	);
	LUT2 #(
		.INIT('h1)
	) name814 (
		_w1338_,
		_w1345_,
		_w1346_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w1325_,
		_w1328_,
		_w1347_
	);
	LUT2 #(
		.INIT('h4)
	) name816 (
		_w1331_,
		_w1347_,
		_w1348_
	);
	LUT2 #(
		.INIT('h4)
	) name817 (
		_w1322_,
		_w1348_,
		_w1349_
	);
	LUT2 #(
		.INIT('h4)
	) name818 (
		_w1346_,
		_w1349_,
		_w1350_
	);
	LUT2 #(
		.INIT('h2)
	) name819 (
		\sa03_reg[1]/P0001 ,
		_w1350_,
		_w1351_
	);
	LUT2 #(
		.INIT('h1)
	) name820 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1352_
	);
	LUT2 #(
		.INIT('h8)
	) name821 (
		\sa03_reg[7]/NET0131 ,
		_w1342_,
		_w1353_
	);
	LUT2 #(
		.INIT('h8)
	) name822 (
		_w1352_,
		_w1353_,
		_w1354_
	);
	LUT2 #(
		.INIT('h1)
	) name823 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1355_
	);
	LUT2 #(
		.INIT('h2)
	) name824 (
		\sa03_reg[2]/P0001 ,
		_w1316_,
		_w1356_
	);
	LUT2 #(
		.INIT('h4)
	) name825 (
		_w1327_,
		_w1355_,
		_w1357_
	);
	LUT2 #(
		.INIT('h8)
	) name826 (
		_w1356_,
		_w1357_,
		_w1358_
	);
	LUT2 #(
		.INIT('h8)
	) name827 (
		_w1327_,
		_w1355_,
		_w1359_
	);
	LUT2 #(
		.INIT('h8)
	) name828 (
		\sa03_reg[4]/P0001 ,
		_w1359_,
		_w1360_
	);
	LUT2 #(
		.INIT('h1)
	) name829 (
		_w1354_,
		_w1358_,
		_w1361_
	);
	LUT2 #(
		.INIT('h4)
	) name830 (
		_w1360_,
		_w1361_,
		_w1362_
	);
	LUT2 #(
		.INIT('h1)
	) name831 (
		\sa03_reg[1]/P0001 ,
		_w1362_,
		_w1363_
	);
	LUT2 #(
		.INIT('h8)
	) name832 (
		\sa03_reg[4]/P0001 ,
		_w1329_,
		_w1364_
	);
	LUT2 #(
		.INIT('h8)
	) name833 (
		\sa03_reg[7]/NET0131 ,
		_w1364_,
		_w1365_
	);
	LUT2 #(
		.INIT('h4)
	) name834 (
		\sa03_reg[2]/P0001 ,
		_w1365_,
		_w1366_
	);
	LUT2 #(
		.INIT('h4)
	) name835 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1367_
	);
	LUT2 #(
		.INIT('h4)
	) name836 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1368_
	);
	LUT2 #(
		.INIT('h8)
	) name837 (
		_w1367_,
		_w1368_,
		_w1369_
	);
	LUT2 #(
		.INIT('h4)
	) name838 (
		\sa03_reg[5]/P0001 ,
		_w1341_,
		_w1370_
	);
	LUT2 #(
		.INIT('h8)
	) name839 (
		\sa03_reg[3]/P0001 ,
		_w1370_,
		_w1371_
	);
	LUT2 #(
		.INIT('h1)
	) name840 (
		_w1369_,
		_w1371_,
		_w1372_
	);
	LUT2 #(
		.INIT('h1)
	) name841 (
		\sa03_reg[2]/P0001 ,
		_w1372_,
		_w1373_
	);
	LUT2 #(
		.INIT('h8)
	) name842 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1374_
	);
	LUT2 #(
		.INIT('h8)
	) name843 (
		\sa03_reg[4]/P0001 ,
		_w1339_,
		_w1375_
	);
	LUT2 #(
		.INIT('h1)
	) name844 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1376_
	);
	LUT2 #(
		.INIT('h4)
	) name845 (
		\sa03_reg[4]/P0001 ,
		_w1376_,
		_w1377_
	);
	LUT2 #(
		.INIT('h1)
	) name846 (
		_w1375_,
		_w1377_,
		_w1378_
	);
	LUT2 #(
		.INIT('h2)
	) name847 (
		_w1374_,
		_w1378_,
		_w1379_
	);
	LUT2 #(
		.INIT('h4)
	) name848 (
		\sa03_reg[5]/P0001 ,
		_w1318_,
		_w1380_
	);
	LUT2 #(
		.INIT('h8)
	) name849 (
		\sa03_reg[2]/P0001 ,
		_w1334_,
		_w1381_
	);
	LUT2 #(
		.INIT('h8)
	) name850 (
		_w1380_,
		_w1381_,
		_w1382_
	);
	LUT2 #(
		.INIT('h1)
	) name851 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1383_
	);
	LUT2 #(
		.INIT('h2)
	) name852 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1384_
	);
	LUT2 #(
		.INIT('h1)
	) name853 (
		_w1355_,
		_w1384_,
		_w1385_
	);
	LUT2 #(
		.INIT('h2)
	) name854 (
		_w1383_,
		_w1385_,
		_w1386_
	);
	LUT2 #(
		.INIT('h1)
	) name855 (
		_w1382_,
		_w1386_,
		_w1387_
	);
	LUT2 #(
		.INIT('h4)
	) name856 (
		_w1366_,
		_w1387_,
		_w1388_
	);
	LUT2 #(
		.INIT('h4)
	) name857 (
		_w1379_,
		_w1388_,
		_w1389_
	);
	LUT2 #(
		.INIT('h4)
	) name858 (
		_w1373_,
		_w1389_,
		_w1390_
	);
	LUT2 #(
		.INIT('h4)
	) name859 (
		_w1363_,
		_w1390_,
		_w1391_
	);
	LUT2 #(
		.INIT('h4)
	) name860 (
		_w1351_,
		_w1391_,
		_w1392_
	);
	LUT2 #(
		.INIT('h1)
	) name861 (
		\sa03_reg[0]/P0001 ,
		_w1392_,
		_w1393_
	);
	LUT2 #(
		.INIT('h8)
	) name862 (
		_w1364_,
		_w1374_,
		_w1394_
	);
	LUT2 #(
		.INIT('h8)
	) name863 (
		_w1339_,
		_w1352_,
		_w1395_
	);
	LUT2 #(
		.INIT('h8)
	) name864 (
		\sa03_reg[4]/P0001 ,
		_w1326_,
		_w1396_
	);
	LUT2 #(
		.INIT('h8)
	) name865 (
		\sa03_reg[7]/NET0131 ,
		_w1396_,
		_w1397_
	);
	LUT2 #(
		.INIT('h8)
	) name866 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1398_
	);
	LUT2 #(
		.INIT('h8)
	) name867 (
		_w1341_,
		_w1398_,
		_w1399_
	);
	LUT2 #(
		.INIT('h8)
	) name868 (
		\sa03_reg[5]/P0001 ,
		_w1399_,
		_w1400_
	);
	LUT2 #(
		.INIT('h1)
	) name869 (
		_w1395_,
		_w1397_,
		_w1401_
	);
	LUT2 #(
		.INIT('h4)
	) name870 (
		_w1400_,
		_w1401_,
		_w1402_
	);
	LUT2 #(
		.INIT('h1)
	) name871 (
		\sa03_reg[2]/P0001 ,
		_w1402_,
		_w1403_
	);
	LUT2 #(
		.INIT('h4)
	) name872 (
		\sa03_reg[5]/P0001 ,
		_w1332_,
		_w1404_
	);
	LUT2 #(
		.INIT('h1)
	) name873 (
		_w1380_,
		_w1404_,
		_w1405_
	);
	LUT2 #(
		.INIT('h4)
	) name874 (
		_w1353_,
		_w1405_,
		_w1406_
	);
	LUT2 #(
		.INIT('h2)
	) name875 (
		_w1381_,
		_w1406_,
		_w1407_
	);
	LUT2 #(
		.INIT('h1)
	) name876 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1408_
	);
	LUT2 #(
		.INIT('h8)
	) name877 (
		_w1383_,
		_w1408_,
		_w1409_
	);
	LUT2 #(
		.INIT('h1)
	) name878 (
		_w1394_,
		_w1409_,
		_w1410_
	);
	LUT2 #(
		.INIT('h4)
	) name879 (
		_w1407_,
		_w1410_,
		_w1411_
	);
	LUT2 #(
		.INIT('h4)
	) name880 (
		_w1403_,
		_w1411_,
		_w1412_
	);
	LUT2 #(
		.INIT('h1)
	) name881 (
		\sa03_reg[1]/P0001 ,
		_w1412_,
		_w1413_
	);
	LUT2 #(
		.INIT('h8)
	) name882 (
		_w1329_,
		_w1341_,
		_w1414_
	);
	LUT2 #(
		.INIT('h8)
	) name883 (
		_w1374_,
		_w1414_,
		_w1415_
	);
	LUT2 #(
		.INIT('h8)
	) name884 (
		_w1329_,
		_w1383_,
		_w1416_
	);
	LUT2 #(
		.INIT('h8)
	) name885 (
		\sa03_reg[3]/P0001 ,
		_w1416_,
		_w1417_
	);
	LUT2 #(
		.INIT('h1)
	) name886 (
		_w1328_,
		_w1417_,
		_w1418_
	);
	LUT2 #(
		.INIT('h1)
	) name887 (
		\sa03_reg[2]/P0001 ,
		_w1418_,
		_w1419_
	);
	LUT2 #(
		.INIT('h8)
	) name888 (
		_w1334_,
		_w1342_,
		_w1420_
	);
	LUT2 #(
		.INIT('h4)
	) name889 (
		\sa03_reg[7]/NET0131 ,
		_w1420_,
		_w1421_
	);
	LUT2 #(
		.INIT('h8)
	) name890 (
		\sa03_reg[2]/P0001 ,
		_w1421_,
		_w1422_
	);
	LUT2 #(
		.INIT('h2)
	) name891 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1423_
	);
	LUT2 #(
		.INIT('h4)
	) name892 (
		\sa03_reg[6]/NET0131 ,
		_w1423_,
		_w1424_
	);
	LUT2 #(
		.INIT('h8)
	) name893 (
		_w1376_,
		_w1424_,
		_w1425_
	);
	LUT2 #(
		.INIT('h1)
	) name894 (
		_w1366_,
		_w1425_,
		_w1426_
	);
	LUT2 #(
		.INIT('h4)
	) name895 (
		_w1422_,
		_w1426_,
		_w1427_
	);
	LUT2 #(
		.INIT('h2)
	) name896 (
		\sa03_reg[1]/P0001 ,
		_w1427_,
		_w1428_
	);
	LUT2 #(
		.INIT('h4)
	) name897 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1429_
	);
	LUT2 #(
		.INIT('h8)
	) name898 (
		_w1404_,
		_w1429_,
		_w1430_
	);
	LUT2 #(
		.INIT('h4)
	) name899 (
		\sa03_reg[4]/P0001 ,
		_w1326_,
		_w1431_
	);
	LUT2 #(
		.INIT('h8)
	) name900 (
		_w1316_,
		_w1323_,
		_w1432_
	);
	LUT2 #(
		.INIT('h1)
	) name901 (
		_w1431_,
		_w1432_,
		_w1433_
	);
	LUT2 #(
		.INIT('h2)
	) name902 (
		\sa03_reg[2]/P0001 ,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('h8)
	) name903 (
		\sa03_reg[5]/P0001 ,
		_w1318_,
		_w1435_
	);
	LUT2 #(
		.INIT('h2)
	) name904 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1436_
	);
	LUT2 #(
		.INIT('h2)
	) name905 (
		_w1435_,
		_w1436_,
		_w1437_
	);
	LUT2 #(
		.INIT('h8)
	) name906 (
		_w1334_,
		_w1353_,
		_w1438_
	);
	LUT2 #(
		.INIT('h1)
	) name907 (
		_w1430_,
		_w1437_,
		_w1439_
	);
	LUT2 #(
		.INIT('h4)
	) name908 (
		_w1438_,
		_w1439_,
		_w1440_
	);
	LUT2 #(
		.INIT('h4)
	) name909 (
		_w1434_,
		_w1440_,
		_w1441_
	);
	LUT2 #(
		.INIT('h1)
	) name910 (
		\sa03_reg[1]/P0001 ,
		_w1441_,
		_w1442_
	);
	LUT2 #(
		.INIT('h4)
	) name911 (
		\sa03_reg[5]/P0001 ,
		_w1320_,
		_w1443_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		_w1438_,
		_w1443_,
		_w1444_
	);
	LUT2 #(
		.INIT('h2)
	) name913 (
		\sa03_reg[2]/P0001 ,
		_w1444_,
		_w1445_
	);
	LUT2 #(
		.INIT('h8)
	) name914 (
		\sa03_reg[3]/P0001 ,
		_w1435_,
		_w1446_
	);
	LUT2 #(
		.INIT('h8)
	) name915 (
		_w1383_,
		_w1398_,
		_w1447_
	);
	LUT2 #(
		.INIT('h1)
	) name916 (
		_w1446_,
		_w1447_,
		_w1448_
	);
	LUT2 #(
		.INIT('h2)
	) name917 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1449_
	);
	LUT2 #(
		.INIT('h4)
	) name918 (
		\sa03_reg[4]/P0001 ,
		_w1449_,
		_w1450_
	);
	LUT2 #(
		.INIT('h1)
	) name919 (
		_w1397_,
		_w1450_,
		_w1451_
	);
	LUT2 #(
		.INIT('h8)
	) name920 (
		_w1448_,
		_w1451_,
		_w1452_
	);
	LUT2 #(
		.INIT('h1)
	) name921 (
		\sa03_reg[2]/P0001 ,
		_w1452_,
		_w1453_
	);
	LUT2 #(
		.INIT('h8)
	) name922 (
		\sa03_reg[5]/P0001 ,
		_w1423_,
		_w1454_
	);
	LUT2 #(
		.INIT('h4)
	) name923 (
		\sa03_reg[4]/P0001 ,
		_w1355_,
		_w1455_
	);
	LUT2 #(
		.INIT('h1)
	) name924 (
		_w1370_,
		_w1454_,
		_w1456_
	);
	LUT2 #(
		.INIT('h4)
	) name925 (
		_w1455_,
		_w1456_,
		_w1457_
	);
	LUT2 #(
		.INIT('h1)
	) name926 (
		\sa03_reg[2]/P0001 ,
		_w1457_,
		_w1458_
	);
	LUT2 #(
		.INIT('h8)
	) name927 (
		\sa03_reg[5]/P0001 ,
		_w1432_,
		_w1459_
	);
	LUT2 #(
		.INIT('h4)
	) name928 (
		\sa03_reg[7]/NET0131 ,
		_w1355_,
		_w1460_
	);
	LUT2 #(
		.INIT('h8)
	) name929 (
		_w1334_,
		_w1460_,
		_w1461_
	);
	LUT2 #(
		.INIT('h8)
	) name930 (
		_w1375_,
		_w1408_,
		_w1462_
	);
	LUT2 #(
		.INIT('h8)
	) name931 (
		_w1332_,
		_w1423_,
		_w1463_
	);
	LUT2 #(
		.INIT('h1)
	) name932 (
		_w1459_,
		_w1463_,
		_w1464_
	);
	LUT2 #(
		.INIT('h1)
	) name933 (
		_w1461_,
		_w1462_,
		_w1465_
	);
	LUT2 #(
		.INIT('h8)
	) name934 (
		_w1464_,
		_w1465_,
		_w1466_
	);
	LUT2 #(
		.INIT('h4)
	) name935 (
		_w1458_,
		_w1466_,
		_w1467_
	);
	LUT2 #(
		.INIT('h2)
	) name936 (
		\sa03_reg[1]/P0001 ,
		_w1467_,
		_w1468_
	);
	LUT2 #(
		.INIT('h8)
	) name937 (
		_w1318_,
		_w1454_,
		_w1469_
	);
	LUT2 #(
		.INIT('h1)
	) name938 (
		_w1445_,
		_w1469_,
		_w1470_
	);
	LUT2 #(
		.INIT('h4)
	) name939 (
		_w1453_,
		_w1470_,
		_w1471_
	);
	LUT2 #(
		.INIT('h1)
	) name940 (
		_w1442_,
		_w1468_,
		_w1472_
	);
	LUT2 #(
		.INIT('h8)
	) name941 (
		_w1471_,
		_w1472_,
		_w1473_
	);
	LUT2 #(
		.INIT('h2)
	) name942 (
		\sa03_reg[0]/P0001 ,
		_w1473_,
		_w1474_
	);
	LUT2 #(
		.INIT('h1)
	) name943 (
		_w1415_,
		_w1419_,
		_w1475_
	);
	LUT2 #(
		.INIT('h4)
	) name944 (
		_w1428_,
		_w1475_,
		_w1476_
	);
	LUT2 #(
		.INIT('h4)
	) name945 (
		_w1413_,
		_w1476_,
		_w1477_
	);
	LUT2 #(
		.INIT('h4)
	) name946 (
		_w1393_,
		_w1477_,
		_w1478_
	);
	LUT2 #(
		.INIT('h4)
	) name947 (
		_w1474_,
		_w1478_,
		_w1479_
	);
	LUT2 #(
		.INIT('h8)
	) name948 (
		_w1339_,
		_w1423_,
		_w1480_
	);
	LUT2 #(
		.INIT('h1)
	) name949 (
		_w1459_,
		_w1480_,
		_w1481_
	);
	LUT2 #(
		.INIT('h8)
	) name950 (
		\sa03_reg[4]/P0001 ,
		_w1318_,
		_w1482_
	);
	LUT2 #(
		.INIT('h4)
	) name951 (
		\sa03_reg[4]/P0001 ,
		_w1328_,
		_w1483_
	);
	LUT2 #(
		.INIT('h1)
	) name952 (
		_w1331_,
		_w1482_,
		_w1484_
	);
	LUT2 #(
		.INIT('h4)
	) name953 (
		_w1483_,
		_w1484_,
		_w1485_
	);
	LUT2 #(
		.INIT('h2)
	) name954 (
		\sa03_reg[2]/P0001 ,
		_w1485_,
		_w1486_
	);
	LUT2 #(
		.INIT('h2)
	) name955 (
		_w1481_,
		_w1486_,
		_w1487_
	);
	LUT2 #(
		.INIT('h2)
	) name956 (
		\sa03_reg[1]/P0001 ,
		_w1487_,
		_w1488_
	);
	LUT2 #(
		.INIT('h1)
	) name957 (
		_w1399_,
		_w1438_,
		_w1489_
	);
	LUT2 #(
		.INIT('h8)
	) name958 (
		_w1355_,
		_w1383_,
		_w1490_
	);
	LUT2 #(
		.INIT('h2)
	) name959 (
		_w1489_,
		_w1490_,
		_w1491_
	);
	LUT2 #(
		.INIT('h2)
	) name960 (
		\sa03_reg[2]/P0001 ,
		_w1491_,
		_w1492_
	);
	LUT2 #(
		.INIT('h1)
	) name961 (
		_w1317_,
		_w1380_,
		_w1493_
	);
	LUT2 #(
		.INIT('h4)
	) name962 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[2]/P0001 ,
		_w1494_
	);
	LUT2 #(
		.INIT('h4)
	) name963 (
		_w1493_,
		_w1494_,
		_w1495_
	);
	LUT2 #(
		.INIT('h8)
	) name964 (
		_w1374_,
		_w1404_,
		_w1496_
	);
	LUT2 #(
		.INIT('h8)
	) name965 (
		_w1342_,
		_w1383_,
		_w1497_
	);
	LUT2 #(
		.INIT('h2)
	) name966 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1498_
	);
	LUT2 #(
		.INIT('h4)
	) name967 (
		\sa03_reg[5]/P0001 ,
		_w1498_,
		_w1499_
	);
	LUT2 #(
		.INIT('h4)
	) name968 (
		_w1368_,
		_w1499_,
		_w1500_
	);
	LUT2 #(
		.INIT('h1)
	) name969 (
		_w1335_,
		_w1497_,
		_w1501_
	);
	LUT2 #(
		.INIT('h4)
	) name970 (
		_w1500_,
		_w1501_,
		_w1502_
	);
	LUT2 #(
		.INIT('h1)
	) name971 (
		\sa03_reg[2]/P0001 ,
		_w1502_,
		_w1503_
	);
	LUT2 #(
		.INIT('h8)
	) name972 (
		_w1408_,
		_w1449_,
		_w1504_
	);
	LUT2 #(
		.INIT('h4)
	) name973 (
		\sa03_reg[2]/P0001 ,
		_w1504_,
		_w1505_
	);
	LUT2 #(
		.INIT('h1)
	) name974 (
		_w1365_,
		_w1505_,
		_w1506_
	);
	LUT2 #(
		.INIT('h4)
	) name975 (
		_w1373_,
		_w1506_,
		_w1507_
	);
	LUT2 #(
		.INIT('h1)
	) name976 (
		\sa03_reg[1]/P0001 ,
		_w1507_,
		_w1508_
	);
	LUT2 #(
		.INIT('h1)
	) name977 (
		_w1495_,
		_w1496_,
		_w1509_
	);
	LUT2 #(
		.INIT('h4)
	) name978 (
		_w1503_,
		_w1509_,
		_w1510_
	);
	LUT2 #(
		.INIT('h4)
	) name979 (
		_w1492_,
		_w1510_,
		_w1511_
	);
	LUT2 #(
		.INIT('h4)
	) name980 (
		_w1488_,
		_w1511_,
		_w1512_
	);
	LUT2 #(
		.INIT('h4)
	) name981 (
		_w1508_,
		_w1512_,
		_w1513_
	);
	LUT2 #(
		.INIT('h2)
	) name982 (
		\sa03_reg[0]/P0001 ,
		_w1513_,
		_w1514_
	);
	LUT2 #(
		.INIT('h1)
	) name983 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1515_
	);
	LUT2 #(
		.INIT('h8)
	) name984 (
		_w1460_,
		_w1515_,
		_w1516_
	);
	LUT2 #(
		.INIT('h4)
	) name985 (
		_w1378_,
		_w1436_,
		_w1517_
	);
	LUT2 #(
		.INIT('h2)
	) name986 (
		\sa03_reg[1]/P0001 ,
		_w1400_,
		_w1518_
	);
	LUT2 #(
		.INIT('h4)
	) name987 (
		_w1516_,
		_w1518_,
		_w1519_
	);
	LUT2 #(
		.INIT('h4)
	) name988 (
		_w1517_,
		_w1519_,
		_w1520_
	);
	LUT2 #(
		.INIT('h8)
	) name989 (
		\sa03_reg[3]/P0001 ,
		_w1384_,
		_w1521_
	);
	LUT2 #(
		.INIT('h8)
	) name990 (
		_w1449_,
		_w1521_,
		_w1522_
	);
	LUT2 #(
		.INIT('h4)
	) name991 (
		\sa03_reg[2]/P0001 ,
		_w1317_,
		_w1523_
	);
	LUT2 #(
		.INIT('h1)
	) name992 (
		_w1324_,
		_w1408_,
		_w1524_
	);
	LUT2 #(
		.INIT('h2)
	) name993 (
		_w1330_,
		_w1524_,
		_w1525_
	);
	LUT2 #(
		.INIT('h8)
	) name994 (
		\sa03_reg[4]/P0001 ,
		_w1328_,
		_w1526_
	);
	LUT2 #(
		.INIT('h1)
	) name995 (
		\sa03_reg[1]/P0001 ,
		_w1497_,
		_w1527_
	);
	LUT2 #(
		.INIT('h4)
	) name996 (
		_w1522_,
		_w1527_,
		_w1528_
	);
	LUT2 #(
		.INIT('h1)
	) name997 (
		_w1523_,
		_w1525_,
		_w1529_
	);
	LUT2 #(
		.INIT('h4)
	) name998 (
		_w1526_,
		_w1529_,
		_w1530_
	);
	LUT2 #(
		.INIT('h8)
	) name999 (
		_w1528_,
		_w1530_,
		_w1531_
	);
	LUT2 #(
		.INIT('h1)
	) name1000 (
		_w1520_,
		_w1531_,
		_w1532_
	);
	LUT2 #(
		.INIT('h8)
	) name1001 (
		\sa03_reg[4]/P0001 ,
		_w1355_,
		_w1533_
	);
	LUT2 #(
		.INIT('h4)
	) name1002 (
		_w1323_,
		_w1324_,
		_w1534_
	);
	LUT2 #(
		.INIT('h1)
	) name1003 (
		_w1533_,
		_w1534_,
		_w1535_
	);
	LUT2 #(
		.INIT('h1)
	) name1004 (
		_w1316_,
		_w1535_,
		_w1536_
	);
	LUT2 #(
		.INIT('h8)
	) name1005 (
		_w1367_,
		_w1398_,
		_w1537_
	);
	LUT2 #(
		.INIT('h1)
	) name1006 (
		\sa03_reg[2]/P0001 ,
		_w1537_,
		_w1538_
	);
	LUT2 #(
		.INIT('h4)
	) name1007 (
		_w1421_,
		_w1538_,
		_w1539_
	);
	LUT2 #(
		.INIT('h4)
	) name1008 (
		_w1536_,
		_w1539_,
		_w1540_
	);
	LUT2 #(
		.INIT('h8)
	) name1009 (
		_w1352_,
		_w1355_,
		_w1541_
	);
	LUT2 #(
		.INIT('h2)
	) name1010 (
		\sa03_reg[2]/P0001 ,
		_w1541_,
		_w1542_
	);
	LUT2 #(
		.INIT('h4)
	) name1011 (
		_w1526_,
		_w1542_,
		_w1543_
	);
	LUT2 #(
		.INIT('h1)
	) name1012 (
		_w1540_,
		_w1543_,
		_w1544_
	);
	LUT2 #(
		.INIT('h1)
	) name1013 (
		_w1532_,
		_w1544_,
		_w1545_
	);
	LUT2 #(
		.INIT('h1)
	) name1014 (
		\sa03_reg[0]/P0001 ,
		_w1545_,
		_w1546_
	);
	LUT2 #(
		.INIT('h8)
	) name1015 (
		_w1341_,
		_w1355_,
		_w1547_
	);
	LUT2 #(
		.INIT('h4)
	) name1016 (
		\sa03_reg[6]/NET0131 ,
		_w1480_,
		_w1548_
	);
	LUT2 #(
		.INIT('h1)
	) name1017 (
		_w1409_,
		_w1547_,
		_w1549_
	);
	LUT2 #(
		.INIT('h4)
	) name1018 (
		_w1548_,
		_w1549_,
		_w1550_
	);
	LUT2 #(
		.INIT('h2)
	) name1019 (
		\sa03_reg[1]/P0001 ,
		_w1550_,
		_w1551_
	);
	LUT2 #(
		.INIT('h8)
	) name1020 (
		_w1316_,
		_w1380_,
		_w1552_
	);
	LUT2 #(
		.INIT('h1)
	) name1021 (
		_w1551_,
		_w1552_,
		_w1553_
	);
	LUT2 #(
		.INIT('h2)
	) name1022 (
		\sa03_reg[2]/P0001 ,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('h4)
	) name1023 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1555_
	);
	LUT2 #(
		.INIT('h8)
	) name1024 (
		_w1376_,
		_w1408_,
		_w1556_
	);
	LUT2 #(
		.INIT('h4)
	) name1025 (
		_w1555_,
		_w1556_,
		_w1557_
	);
	LUT2 #(
		.INIT('h2)
	) name1026 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[2]/P0001 ,
		_w1558_
	);
	LUT2 #(
		.INIT('h8)
	) name1027 (
		_w1417_,
		_w1558_,
		_w1559_
	);
	LUT2 #(
		.INIT('h8)
	) name1028 (
		_w1365_,
		_w1429_,
		_w1560_
	);
	LUT2 #(
		.INIT('h8)
	) name1029 (
		_w1339_,
		_w1368_,
		_w1561_
	);
	LUT2 #(
		.INIT('h2)
	) name1030 (
		\sa03_reg[2]/P0001 ,
		_w1561_,
		_w1562_
	);
	LUT2 #(
		.INIT('h4)
	) name1031 (
		\sa03_reg[7]/NET0131 ,
		_w1424_,
		_w1563_
	);
	LUT2 #(
		.INIT('h2)
	) name1032 (
		_w1562_,
		_w1563_,
		_w1564_
	);
	LUT2 #(
		.INIT('h4)
	) name1033 (
		\sa03_reg[6]/NET0131 ,
		_w1340_,
		_w1565_
	);
	LUT2 #(
		.INIT('h4)
	) name1034 (
		\sa03_reg[7]/NET0131 ,
		_w1396_,
		_w1566_
	);
	LUT2 #(
		.INIT('h1)
	) name1035 (
		\sa03_reg[2]/P0001 ,
		_w1365_,
		_w1567_
	);
	LUT2 #(
		.INIT('h1)
	) name1036 (
		_w1565_,
		_w1566_,
		_w1568_
	);
	LUT2 #(
		.INIT('h8)
	) name1037 (
		_w1567_,
		_w1568_,
		_w1569_
	);
	LUT2 #(
		.INIT('h1)
	) name1038 (
		_w1564_,
		_w1569_,
		_w1570_
	);
	LUT2 #(
		.INIT('h8)
	) name1039 (
		_w1342_,
		_w1352_,
		_w1571_
	);
	LUT2 #(
		.INIT('h4)
	) name1040 (
		\sa03_reg[6]/NET0131 ,
		_w1317_,
		_w1572_
	);
	LUT2 #(
		.INIT('h1)
	) name1041 (
		_w1571_,
		_w1572_,
		_w1573_
	);
	LUT2 #(
		.INIT('h4)
	) name1042 (
		_w1570_,
		_w1573_,
		_w1574_
	);
	LUT2 #(
		.INIT('h1)
	) name1043 (
		\sa03_reg[1]/P0001 ,
		_w1574_,
		_w1575_
	);
	LUT2 #(
		.INIT('h1)
	) name1044 (
		_w1557_,
		_w1559_,
		_w1576_
	);
	LUT2 #(
		.INIT('h4)
	) name1045 (
		_w1560_,
		_w1576_,
		_w1577_
	);
	LUT2 #(
		.INIT('h4)
	) name1046 (
		_w1554_,
		_w1577_,
		_w1578_
	);
	LUT2 #(
		.INIT('h4)
	) name1047 (
		_w1575_,
		_w1578_,
		_w1579_
	);
	LUT2 #(
		.INIT('h4)
	) name1048 (
		_w1546_,
		_w1579_,
		_w1580_
	);
	LUT2 #(
		.INIT('h4)
	) name1049 (
		_w1514_,
		_w1580_,
		_w1581_
	);
	LUT2 #(
		.INIT('h2)
	) name1050 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1582_
	);
	LUT2 #(
		.INIT('h4)
	) name1051 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1583_
	);
	LUT2 #(
		.INIT('h8)
	) name1052 (
		_w1582_,
		_w1583_,
		_w1584_
	);
	LUT2 #(
		.INIT('h8)
	) name1053 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1585_
	);
	LUT2 #(
		.INIT('h1)
	) name1054 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1586_
	);
	LUT2 #(
		.INIT('h8)
	) name1055 (
		_w1585_,
		_w1586_,
		_w1587_
	);
	LUT2 #(
		.INIT('h1)
	) name1056 (
		_w1584_,
		_w1587_,
		_w1588_
	);
	LUT2 #(
		.INIT('h1)
	) name1057 (
		\sa10_reg[2]/P0001 ,
		_w1588_,
		_w1589_
	);
	LUT2 #(
		.INIT('h4)
	) name1058 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1590_
	);
	LUT2 #(
		.INIT('h8)
	) name1059 (
		_w1585_,
		_w1590_,
		_w1591_
	);
	LUT2 #(
		.INIT('h8)
	) name1060 (
		\sa10_reg[4]/P0001 ,
		_w1591_,
		_w1592_
	);
	LUT2 #(
		.INIT('h2)
	) name1061 (
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1593_
	);
	LUT2 #(
		.INIT('h8)
	) name1062 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1594_
	);
	LUT2 #(
		.INIT('h8)
	) name1063 (
		_w1593_,
		_w1594_,
		_w1595_
	);
	LUT2 #(
		.INIT('h1)
	) name1064 (
		_w1592_,
		_w1595_,
		_w1596_
	);
	LUT2 #(
		.INIT('h4)
	) name1065 (
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1597_
	);
	LUT2 #(
		.INIT('h2)
	) name1066 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		_w1598_
	);
	LUT2 #(
		.INIT('h8)
	) name1067 (
		_w1597_,
		_w1598_,
		_w1599_
	);
	LUT2 #(
		.INIT('h1)
	) name1068 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1600_
	);
	LUT2 #(
		.INIT('h4)
	) name1069 (
		\sa10_reg[4]/P0001 ,
		_w1600_,
		_w1601_
	);
	LUT2 #(
		.INIT('h4)
	) name1070 (
		\sa10_reg[6]/NET0131 ,
		_w1601_,
		_w1602_
	);
	LUT2 #(
		.INIT('h1)
	) name1071 (
		_w1599_,
		_w1602_,
		_w1603_
	);
	LUT2 #(
		.INIT('h8)
	) name1072 (
		_w1596_,
		_w1603_,
		_w1604_
	);
	LUT2 #(
		.INIT('h2)
	) name1073 (
		\sa10_reg[2]/P0001 ,
		_w1604_,
		_w1605_
	);
	LUT2 #(
		.INIT('h8)
	) name1074 (
		_w1594_,
		_w1600_,
		_w1606_
	);
	LUT2 #(
		.INIT('h4)
	) name1075 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1607_
	);
	LUT2 #(
		.INIT('h4)
	) name1076 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1608_
	);
	LUT2 #(
		.INIT('h8)
	) name1077 (
		_w1607_,
		_w1608_,
		_w1609_
	);
	LUT2 #(
		.INIT('h1)
	) name1078 (
		_w1606_,
		_w1609_,
		_w1610_
	);
	LUT2 #(
		.INIT('h1)
	) name1079 (
		\sa10_reg[2]/P0001 ,
		_w1610_,
		_w1611_
	);
	LUT2 #(
		.INIT('h8)
	) name1080 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1612_
	);
	LUT2 #(
		.INIT('h8)
	) name1081 (
		_w1582_,
		_w1612_,
		_w1613_
	);
	LUT2 #(
		.INIT('h1)
	) name1082 (
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1614_
	);
	LUT2 #(
		.INIT('h8)
	) name1083 (
		\sa10_reg[5]/P0001 ,
		_w1614_,
		_w1615_
	);
	LUT2 #(
		.INIT('h4)
	) name1084 (
		\sa10_reg[3]/P0001 ,
		_w1615_,
		_w1616_
	);
	LUT2 #(
		.INIT('h1)
	) name1085 (
		\sa10_reg[2]/P0001 ,
		_w1616_,
		_w1617_
	);
	LUT2 #(
		.INIT('h4)
	) name1086 (
		\sa10_reg[5]/P0001 ,
		_w1593_,
		_w1618_
	);
	LUT2 #(
		.INIT('h8)
	) name1087 (
		\sa10_reg[7]/NET0131 ,
		_w1594_,
		_w1619_
	);
	LUT2 #(
		.INIT('h2)
	) name1088 (
		\sa10_reg[2]/P0001 ,
		_w1618_,
		_w1620_
	);
	LUT2 #(
		.INIT('h4)
	) name1089 (
		_w1619_,
		_w1620_,
		_w1621_
	);
	LUT2 #(
		.INIT('h1)
	) name1090 (
		_w1617_,
		_w1621_,
		_w1622_
	);
	LUT2 #(
		.INIT('h1)
	) name1091 (
		_w1611_,
		_w1613_,
		_w1623_
	);
	LUT2 #(
		.INIT('h4)
	) name1092 (
		_w1622_,
		_w1623_,
		_w1624_
	);
	LUT2 #(
		.INIT('h1)
	) name1093 (
		\sa10_reg[1]/P0001 ,
		_w1624_,
		_w1625_
	);
	LUT2 #(
		.INIT('h8)
	) name1094 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1626_
	);
	LUT2 #(
		.INIT('h2)
	) name1095 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1627_
	);
	LUT2 #(
		.INIT('h8)
	) name1096 (
		_w1626_,
		_w1627_,
		_w1628_
	);
	LUT2 #(
		.INIT('h2)
	) name1097 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1629_
	);
	LUT2 #(
		.INIT('h4)
	) name1098 (
		\sa10_reg[6]/NET0131 ,
		_w1594_,
		_w1630_
	);
	LUT2 #(
		.INIT('h8)
	) name1099 (
		_w1629_,
		_w1630_,
		_w1631_
	);
	LUT2 #(
		.INIT('h1)
	) name1100 (
		_w1628_,
		_w1631_,
		_w1632_
	);
	LUT2 #(
		.INIT('h1)
	) name1101 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		_w1633_
	);
	LUT2 #(
		.INIT('h1)
	) name1102 (
		\sa10_reg[5]/P0001 ,
		_w1607_,
		_w1634_
	);
	LUT2 #(
		.INIT('h8)
	) name1103 (
		_w1633_,
		_w1634_,
		_w1635_
	);
	LUT2 #(
		.INIT('h8)
	) name1104 (
		\sa10_reg[4]/P0001 ,
		_w1593_,
		_w1636_
	);
	LUT2 #(
		.INIT('h4)
	) name1105 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1637_
	);
	LUT2 #(
		.INIT('h8)
	) name1106 (
		_w1582_,
		_w1637_,
		_w1638_
	);
	LUT2 #(
		.INIT('h4)
	) name1107 (
		\sa10_reg[3]/P0001 ,
		_w1609_,
		_w1639_
	);
	LUT2 #(
		.INIT('h1)
	) name1108 (
		_w1636_,
		_w1638_,
		_w1640_
	);
	LUT2 #(
		.INIT('h4)
	) name1109 (
		_w1639_,
		_w1640_,
		_w1641_
	);
	LUT2 #(
		.INIT('h2)
	) name1110 (
		\sa10_reg[2]/P0001 ,
		_w1641_,
		_w1642_
	);
	LUT2 #(
		.INIT('h2)
	) name1111 (
		_w1632_,
		_w1635_,
		_w1643_
	);
	LUT2 #(
		.INIT('h4)
	) name1112 (
		_w1642_,
		_w1643_,
		_w1644_
	);
	LUT2 #(
		.INIT('h2)
	) name1113 (
		\sa10_reg[1]/P0001 ,
		_w1644_,
		_w1645_
	);
	LUT2 #(
		.INIT('h1)
	) name1114 (
		_w1589_,
		_w1605_,
		_w1646_
	);
	LUT2 #(
		.INIT('h4)
	) name1115 (
		_w1625_,
		_w1646_,
		_w1647_
	);
	LUT2 #(
		.INIT('h4)
	) name1116 (
		_w1645_,
		_w1647_,
		_w1648_
	);
	LUT2 #(
		.INIT('h2)
	) name1117 (
		\sa10_reg[0]/P0001 ,
		_w1648_,
		_w1649_
	);
	LUT2 #(
		.INIT('h1)
	) name1118 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1650_
	);
	LUT2 #(
		.INIT('h8)
	) name1119 (
		_w1583_,
		_w1650_,
		_w1651_
	);
	LUT2 #(
		.INIT('h8)
	) name1120 (
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1652_
	);
	LUT2 #(
		.INIT('h2)
	) name1121 (
		\sa10_reg[4]/P0001 ,
		_w1652_,
		_w1653_
	);
	LUT2 #(
		.INIT('h2)
	) name1122 (
		_w1598_,
		_w1614_,
		_w1654_
	);
	LUT2 #(
		.INIT('h4)
	) name1123 (
		_w1653_,
		_w1654_,
		_w1655_
	);
	LUT2 #(
		.INIT('h4)
	) name1124 (
		\sa10_reg[7]/NET0131 ,
		_w1583_,
		_w1656_
	);
	LUT2 #(
		.INIT('h8)
	) name1125 (
		_w1585_,
		_w1656_,
		_w1657_
	);
	LUT2 #(
		.INIT('h1)
	) name1126 (
		_w1651_,
		_w1655_,
		_w1658_
	);
	LUT2 #(
		.INIT('h4)
	) name1127 (
		_w1657_,
		_w1658_,
		_w1659_
	);
	LUT2 #(
		.INIT('h1)
	) name1128 (
		\sa10_reg[2]/P0001 ,
		_w1659_,
		_w1660_
	);
	LUT2 #(
		.INIT('h2)
	) name1129 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		_w1661_
	);
	LUT2 #(
		.INIT('h8)
	) name1130 (
		_w1634_,
		_w1661_,
		_w1662_
	);
	LUT2 #(
		.INIT('h4)
	) name1131 (
		_w1653_,
		_w1662_,
		_w1663_
	);
	LUT2 #(
		.INIT('h8)
	) name1132 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		_w1664_
	);
	LUT2 #(
		.INIT('h8)
	) name1133 (
		_w1615_,
		_w1664_,
		_w1665_
	);
	LUT2 #(
		.INIT('h4)
	) name1134 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		_w1666_
	);
	LUT2 #(
		.INIT('h8)
	) name1135 (
		_w1612_,
		_w1666_,
		_w1667_
	);
	LUT2 #(
		.INIT('h1)
	) name1136 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1668_
	);
	LUT2 #(
		.INIT('h8)
	) name1137 (
		\sa10_reg[7]/NET0131 ,
		_w1668_,
		_w1669_
	);
	LUT2 #(
		.INIT('h4)
	) name1138 (
		\sa10_reg[6]/NET0131 ,
		_w1669_,
		_w1670_
	);
	LUT2 #(
		.INIT('h8)
	) name1139 (
		_w1608_,
		_w1627_,
		_w1671_
	);
	LUT2 #(
		.INIT('h4)
	) name1140 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1672_
	);
	LUT2 #(
		.INIT('h8)
	) name1141 (
		\sa10_reg[4]/P0001 ,
		_w1672_,
		_w1673_
	);
	LUT2 #(
		.INIT('h8)
	) name1142 (
		_w1590_,
		_w1673_,
		_w1674_
	);
	LUT2 #(
		.INIT('h1)
	) name1143 (
		\sa10_reg[1]/P0001 ,
		_w1587_,
		_w1675_
	);
	LUT2 #(
		.INIT('h1)
	) name1144 (
		_w1667_,
		_w1671_,
		_w1676_
	);
	LUT2 #(
		.INIT('h8)
	) name1145 (
		_w1675_,
		_w1676_,
		_w1677_
	);
	LUT2 #(
		.INIT('h1)
	) name1146 (
		_w1665_,
		_w1670_,
		_w1678_
	);
	LUT2 #(
		.INIT('h4)
	) name1147 (
		_w1674_,
		_w1678_,
		_w1679_
	);
	LUT2 #(
		.INIT('h8)
	) name1148 (
		_w1677_,
		_w1679_,
		_w1680_
	);
	LUT2 #(
		.INIT('h8)
	) name1149 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1681_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		_w1629_,
		_w1681_,
		_w1682_
	);
	LUT2 #(
		.INIT('h8)
	) name1151 (
		\sa10_reg[4]/P0001 ,
		_w1682_,
		_w1683_
	);
	LUT2 #(
		.INIT('h8)
	) name1152 (
		\sa10_reg[4]/P0001 ,
		_w1626_,
		_w1684_
	);
	LUT2 #(
		.INIT('h1)
	) name1153 (
		_w1601_,
		_w1684_,
		_w1685_
	);
	LUT2 #(
		.INIT('h2)
	) name1154 (
		_w1661_,
		_w1685_,
		_w1686_
	);
	LUT2 #(
		.INIT('h4)
	) name1155 (
		\sa10_reg[5]/P0001 ,
		_w1614_,
		_w1687_
	);
	LUT2 #(
		.INIT('h4)
	) name1156 (
		\sa10_reg[2]/P0001 ,
		_w1687_,
		_w1688_
	);
	LUT2 #(
		.INIT('h4)
	) name1157 (
		\sa10_reg[4]/P0001 ,
		_w1688_,
		_w1689_
	);
	LUT2 #(
		.INIT('h2)
	) name1158 (
		\sa10_reg[1]/P0001 ,
		_w1683_,
		_w1690_
	);
	LUT2 #(
		.INIT('h4)
	) name1159 (
		_w1686_,
		_w1690_,
		_w1691_
	);
	LUT2 #(
		.INIT('h4)
	) name1160 (
		_w1689_,
		_w1691_,
		_w1692_
	);
	LUT2 #(
		.INIT('h1)
	) name1161 (
		_w1680_,
		_w1692_,
		_w1693_
	);
	LUT2 #(
		.INIT('h1)
	) name1162 (
		_w1660_,
		_w1663_,
		_w1694_
	);
	LUT2 #(
		.INIT('h4)
	) name1163 (
		_w1693_,
		_w1694_,
		_w1695_
	);
	LUT2 #(
		.INIT('h1)
	) name1164 (
		\sa10_reg[0]/P0001 ,
		_w1695_,
		_w1696_
	);
	LUT2 #(
		.INIT('h8)
	) name1165 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[2]/P0001 ,
		_w1697_
	);
	LUT2 #(
		.INIT('h4)
	) name1166 (
		\sa10_reg[3]/P0001 ,
		_w1614_,
		_w1698_
	);
	LUT2 #(
		.INIT('h4)
	) name1167 (
		\sa10_reg[6]/NET0131 ,
		_w1626_,
		_w1699_
	);
	LUT2 #(
		.INIT('h8)
	) name1168 (
		\sa10_reg[3]/P0001 ,
		_w1699_,
		_w1700_
	);
	LUT2 #(
		.INIT('h1)
	) name1169 (
		_w1698_,
		_w1700_,
		_w1701_
	);
	LUT2 #(
		.INIT('h1)
	) name1170 (
		\sa10_reg[4]/P0001 ,
		_w1701_,
		_w1702_
	);
	LUT2 #(
		.INIT('h8)
	) name1171 (
		\sa10_reg[4]/P0001 ,
		_w1614_,
		_w1703_
	);
	LUT2 #(
		.INIT('h4)
	) name1172 (
		\sa10_reg[5]/P0001 ,
		_w1703_,
		_w1704_
	);
	LUT2 #(
		.INIT('h1)
	) name1173 (
		_w1702_,
		_w1704_,
		_w1705_
	);
	LUT2 #(
		.INIT('h2)
	) name1174 (
		_w1697_,
		_w1705_,
		_w1706_
	);
	LUT2 #(
		.INIT('h4)
	) name1175 (
		_w1668_,
		_w1699_,
		_w1707_
	);
	LUT2 #(
		.INIT('h4)
	) name1176 (
		\sa10_reg[5]/P0001 ,
		_w1636_,
		_w1708_
	);
	LUT2 #(
		.INIT('h1)
	) name1177 (
		_w1707_,
		_w1708_,
		_w1709_
	);
	LUT2 #(
		.INIT('h1)
	) name1178 (
		\sa10_reg[2]/P0001 ,
		_w1709_,
		_w1710_
	);
	LUT2 #(
		.INIT('h8)
	) name1179 (
		_w1585_,
		_w1668_,
		_w1711_
	);
	LUT2 #(
		.INIT('h4)
	) name1180 (
		\sa10_reg[6]/NET0131 ,
		_w1619_,
		_w1712_
	);
	LUT2 #(
		.INIT('h8)
	) name1181 (
		_w1607_,
		_w1626_,
		_w1713_
	);
	LUT2 #(
		.INIT('h8)
	) name1182 (
		\sa10_reg[2]/P0001 ,
		_w1713_,
		_w1714_
	);
	LUT2 #(
		.INIT('h8)
	) name1183 (
		\sa10_reg[2]/P0001 ,
		_w1627_,
		_w1715_
	);
	LUT2 #(
		.INIT('h8)
	) name1184 (
		_w1614_,
		_w1715_,
		_w1716_
	);
	LUT2 #(
		.INIT('h1)
	) name1185 (
		_w1711_,
		_w1712_,
		_w1717_
	);
	LUT2 #(
		.INIT('h1)
	) name1186 (
		_w1714_,
		_w1716_,
		_w1718_
	);
	LUT2 #(
		.INIT('h8)
	) name1187 (
		_w1717_,
		_w1718_,
		_w1719_
	);
	LUT2 #(
		.INIT('h4)
	) name1188 (
		_w1710_,
		_w1719_,
		_w1720_
	);
	LUT2 #(
		.INIT('h1)
	) name1189 (
		\sa10_reg[1]/P0001 ,
		_w1720_,
		_w1721_
	);
	LUT2 #(
		.INIT('h2)
	) name1190 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[5]/P0001 ,
		_w1722_
	);
	LUT2 #(
		.INIT('h1)
	) name1191 (
		_w1595_,
		_w1698_,
		_w1723_
	);
	LUT2 #(
		.INIT('h2)
	) name1192 (
		_w1722_,
		_w1723_,
		_w1724_
	);
	LUT2 #(
		.INIT('h8)
	) name1193 (
		_w1613_,
		_w1666_,
		_w1725_
	);
	LUT2 #(
		.INIT('h8)
	) name1194 (
		\sa10_reg[5]/P0001 ,
		_w1627_,
		_w1726_
	);
	LUT2 #(
		.INIT('h8)
	) name1195 (
		_w1614_,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('h4)
	) name1196 (
		\sa10_reg[2]/P0001 ,
		_w1727_,
		_w1728_
	);
	LUT2 #(
		.INIT('h8)
	) name1197 (
		\sa10_reg[1]/P0001 ,
		_w1728_,
		_w1729_
	);
	LUT2 #(
		.INIT('h8)
	) name1198 (
		_w1614_,
		_w1668_,
		_w1730_
	);
	LUT2 #(
		.INIT('h4)
	) name1199 (
		\sa10_reg[5]/P0001 ,
		_w1730_,
		_w1731_
	);
	LUT2 #(
		.INIT('h1)
	) name1200 (
		_w1725_,
		_w1731_,
		_w1732_
	);
	LUT2 #(
		.INIT('h4)
	) name1201 (
		_w1724_,
		_w1732_,
		_w1733_
	);
	LUT2 #(
		.INIT('h4)
	) name1202 (
		_w1729_,
		_w1733_,
		_w1734_
	);
	LUT2 #(
		.INIT('h4)
	) name1203 (
		_w1706_,
		_w1734_,
		_w1735_
	);
	LUT2 #(
		.INIT('h4)
	) name1204 (
		_w1721_,
		_w1735_,
		_w1736_
	);
	LUT2 #(
		.INIT('h4)
	) name1205 (
		_w1696_,
		_w1736_,
		_w1737_
	);
	LUT2 #(
		.INIT('h4)
	) name1206 (
		_w1649_,
		_w1737_,
		_w1738_
	);
	LUT2 #(
		.INIT('h1)
	) name1207 (
		_w1581_,
		_w1738_,
		_w1739_
	);
	LUT2 #(
		.INIT('h8)
	) name1208 (
		_w1581_,
		_w1738_,
		_w1740_
	);
	LUT2 #(
		.INIT('h1)
	) name1209 (
		_w1739_,
		_w1740_,
		_w1741_
	);
	LUT2 #(
		.INIT('h1)
	) name1210 (
		_w1479_,
		_w1741_,
		_w1742_
	);
	LUT2 #(
		.INIT('h8)
	) name1211 (
		_w1479_,
		_w1741_,
		_w1743_
	);
	LUT2 #(
		.INIT('h1)
	) name1212 (
		_w1742_,
		_w1743_,
		_w1744_
	);
	LUT2 #(
		.INIT('h2)
	) name1213 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1745_
	);
	LUT2 #(
		.INIT('h2)
	) name1214 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1746_
	);
	LUT2 #(
		.INIT('h8)
	) name1215 (
		\sa21_reg[4]/P0001 ,
		_w1746_,
		_w1747_
	);
	LUT2 #(
		.INIT('h8)
	) name1216 (
		_w1745_,
		_w1747_,
		_w1748_
	);
	LUT2 #(
		.INIT('h8)
	) name1217 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1749_
	);
	LUT2 #(
		.INIT('h8)
	) name1218 (
		\sa21_reg[3]/P0001 ,
		_w1749_,
		_w1750_
	);
	LUT2 #(
		.INIT('h4)
	) name1219 (
		\sa21_reg[4]/P0001 ,
		_w1750_,
		_w1751_
	);
	LUT2 #(
		.INIT('h1)
	) name1220 (
		_w1748_,
		_w1751_,
		_w1752_
	);
	LUT2 #(
		.INIT('h4)
	) name1221 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1753_
	);
	LUT2 #(
		.INIT('h1)
	) name1222 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		_w1754_
	);
	LUT2 #(
		.INIT('h4)
	) name1223 (
		\sa21_reg[5]/P0001 ,
		_w1754_,
		_w1755_
	);
	LUT2 #(
		.INIT('h4)
	) name1224 (
		_w1753_,
		_w1755_,
		_w1756_
	);
	LUT2 #(
		.INIT('h4)
	) name1225 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1757_
	);
	LUT2 #(
		.INIT('h4)
	) name1226 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1758_
	);
	LUT2 #(
		.INIT('h4)
	) name1227 (
		\sa21_reg[4]/P0001 ,
		_w1758_,
		_w1759_
	);
	LUT2 #(
		.INIT('h8)
	) name1228 (
		_w1757_,
		_w1759_,
		_w1760_
	);
	LUT2 #(
		.INIT('h2)
	) name1229 (
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1761_
	);
	LUT2 #(
		.INIT('h8)
	) name1230 (
		\sa21_reg[4]/P0001 ,
		_w1761_,
		_w1762_
	);
	LUT2 #(
		.INIT('h4)
	) name1231 (
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1763_
	);
	LUT2 #(
		.INIT('h8)
	) name1232 (
		\sa21_reg[5]/P0001 ,
		_w1763_,
		_w1764_
	);
	LUT2 #(
		.INIT('h4)
	) name1233 (
		\sa21_reg[4]/P0001 ,
		_w1764_,
		_w1765_
	);
	LUT2 #(
		.INIT('h1)
	) name1234 (
		_w1760_,
		_w1762_,
		_w1766_
	);
	LUT2 #(
		.INIT('h4)
	) name1235 (
		_w1765_,
		_w1766_,
		_w1767_
	);
	LUT2 #(
		.INIT('h2)
	) name1236 (
		\sa21_reg[2]/P0001 ,
		_w1767_,
		_w1768_
	);
	LUT2 #(
		.INIT('h2)
	) name1237 (
		_w1752_,
		_w1756_,
		_w1769_
	);
	LUT2 #(
		.INIT('h4)
	) name1238 (
		_w1768_,
		_w1769_,
		_w1770_
	);
	LUT2 #(
		.INIT('h2)
	) name1239 (
		\sa21_reg[1]/P0001 ,
		_w1770_,
		_w1771_
	);
	LUT2 #(
		.INIT('h2)
	) name1240 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1772_
	);
	LUT2 #(
		.INIT('h4)
	) name1241 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w1773_
	);
	LUT2 #(
		.INIT('h8)
	) name1242 (
		_w1772_,
		_w1773_,
		_w1774_
	);
	LUT2 #(
		.INIT('h4)
	) name1243 (
		\sa21_reg[4]/P0001 ,
		_w1761_,
		_w1775_
	);
	LUT2 #(
		.INIT('h8)
	) name1244 (
		\sa21_reg[5]/P0001 ,
		_w1775_,
		_w1776_
	);
	LUT2 #(
		.INIT('h1)
	) name1245 (
		_w1774_,
		_w1776_,
		_w1777_
	);
	LUT2 #(
		.INIT('h1)
	) name1246 (
		\sa21_reg[2]/P0001 ,
		_w1777_,
		_w1778_
	);
	LUT2 #(
		.INIT('h8)
	) name1247 (
		\sa21_reg[3]/P0001 ,
		_w1761_,
		_w1779_
	);
	LUT2 #(
		.INIT('h8)
	) name1248 (
		\sa21_reg[4]/P0001 ,
		_w1779_,
		_w1780_
	);
	LUT2 #(
		.INIT('h8)
	) name1249 (
		\sa21_reg[6]/NET0131 ,
		_w1749_,
		_w1781_
	);
	LUT2 #(
		.INIT('h8)
	) name1250 (
		_w1773_,
		_w1781_,
		_w1782_
	);
	LUT2 #(
		.INIT('h1)
	) name1251 (
		_w1780_,
		_w1782_,
		_w1783_
	);
	LUT2 #(
		.INIT('h1)
	) name1252 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1784_
	);
	LUT2 #(
		.INIT('h4)
	) name1253 (
		\sa21_reg[4]/P0001 ,
		_w1784_,
		_w1785_
	);
	LUT2 #(
		.INIT('h4)
	) name1254 (
		\sa21_reg[6]/NET0131 ,
		_w1785_,
		_w1786_
	);
	LUT2 #(
		.INIT('h2)
	) name1255 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		_w1787_
	);
	LUT2 #(
		.INIT('h8)
	) name1256 (
		_w1763_,
		_w1787_,
		_w1788_
	);
	LUT2 #(
		.INIT('h1)
	) name1257 (
		_w1786_,
		_w1788_,
		_w1789_
	);
	LUT2 #(
		.INIT('h8)
	) name1258 (
		_w1783_,
		_w1789_,
		_w1790_
	);
	LUT2 #(
		.INIT('h2)
	) name1259 (
		\sa21_reg[2]/P0001 ,
		_w1790_,
		_w1791_
	);
	LUT2 #(
		.INIT('h8)
	) name1260 (
		\sa21_reg[4]/P0001 ,
		_w1764_,
		_w1792_
	);
	LUT2 #(
		.INIT('h4)
	) name1261 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1793_
	);
	LUT2 #(
		.INIT('h8)
	) name1262 (
		_w1758_,
		_w1793_,
		_w1794_
	);
	LUT2 #(
		.INIT('h8)
	) name1263 (
		\sa21_reg[4]/P0001 ,
		_w1784_,
		_w1795_
	);
	LUT2 #(
		.INIT('h8)
	) name1264 (
		\sa21_reg[3]/P0001 ,
		_w1795_,
		_w1796_
	);
	LUT2 #(
		.INIT('h1)
	) name1265 (
		_w1794_,
		_w1796_,
		_w1797_
	);
	LUT2 #(
		.INIT('h1)
	) name1266 (
		\sa21_reg[2]/P0001 ,
		_w1797_,
		_w1798_
	);
	LUT2 #(
		.INIT('h1)
	) name1267 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1799_
	);
	LUT2 #(
		.INIT('h8)
	) name1268 (
		_w1772_,
		_w1799_,
		_w1800_
	);
	LUT2 #(
		.INIT('h1)
	) name1269 (
		\sa21_reg[2]/P0001 ,
		_w1800_,
		_w1801_
	);
	LUT2 #(
		.INIT('h8)
	) name1270 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w1802_
	);
	LUT2 #(
		.INIT('h8)
	) name1271 (
		\sa21_reg[7]/P0001 ,
		_w1802_,
		_w1803_
	);
	LUT2 #(
		.INIT('h4)
	) name1272 (
		\sa21_reg[5]/P0001 ,
		_w1761_,
		_w1804_
	);
	LUT2 #(
		.INIT('h2)
	) name1273 (
		\sa21_reg[2]/P0001 ,
		_w1803_,
		_w1805_
	);
	LUT2 #(
		.INIT('h4)
	) name1274 (
		_w1804_,
		_w1805_,
		_w1806_
	);
	LUT2 #(
		.INIT('h1)
	) name1275 (
		_w1801_,
		_w1806_,
		_w1807_
	);
	LUT2 #(
		.INIT('h1)
	) name1276 (
		_w1792_,
		_w1798_,
		_w1808_
	);
	LUT2 #(
		.INIT('h4)
	) name1277 (
		_w1807_,
		_w1808_,
		_w1809_
	);
	LUT2 #(
		.INIT('h1)
	) name1278 (
		\sa21_reg[1]/P0001 ,
		_w1809_,
		_w1810_
	);
	LUT2 #(
		.INIT('h1)
	) name1279 (
		_w1778_,
		_w1791_,
		_w1811_
	);
	LUT2 #(
		.INIT('h4)
	) name1280 (
		_w1771_,
		_w1811_,
		_w1812_
	);
	LUT2 #(
		.INIT('h4)
	) name1281 (
		_w1810_,
		_w1812_,
		_w1813_
	);
	LUT2 #(
		.INIT('h2)
	) name1282 (
		\sa21_reg[0]/P0001 ,
		_w1813_,
		_w1814_
	);
	LUT2 #(
		.INIT('h1)
	) name1283 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w1815_
	);
	LUT2 #(
		.INIT('h8)
	) name1284 (
		\sa21_reg[7]/P0001 ,
		_w1815_,
		_w1816_
	);
	LUT2 #(
		.INIT('h4)
	) name1285 (
		\sa21_reg[6]/NET0131 ,
		_w1816_,
		_w1817_
	);
	LUT2 #(
		.INIT('h8)
	) name1286 (
		_w1787_,
		_w1793_,
		_w1818_
	);
	LUT2 #(
		.INIT('h8)
	) name1287 (
		\sa21_reg[2]/P0001 ,
		_w1745_,
		_w1819_
	);
	LUT2 #(
		.INIT('h8)
	) name1288 (
		_w1746_,
		_w1819_,
		_w1820_
	);
	LUT2 #(
		.INIT('h4)
	) name1289 (
		\sa21_reg[2]/P0001 ,
		_w1803_,
		_w1821_
	);
	LUT2 #(
		.INIT('h8)
	) name1290 (
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1822_
	);
	LUT2 #(
		.INIT('h4)
	) name1291 (
		\sa21_reg[5]/P0001 ,
		_w1822_,
		_w1823_
	);
	LUT2 #(
		.INIT('h8)
	) name1292 (
		_w1773_,
		_w1823_,
		_w1824_
	);
	LUT2 #(
		.INIT('h1)
	) name1293 (
		_w1776_,
		_w1818_,
		_w1825_
	);
	LUT2 #(
		.INIT('h1)
	) name1294 (
		_w1817_,
		_w1820_,
		_w1826_
	);
	LUT2 #(
		.INIT('h1)
	) name1295 (
		_w1821_,
		_w1824_,
		_w1827_
	);
	LUT2 #(
		.INIT('h8)
	) name1296 (
		_w1826_,
		_w1827_,
		_w1828_
	);
	LUT2 #(
		.INIT('h8)
	) name1297 (
		_w1825_,
		_w1828_,
		_w1829_
	);
	LUT2 #(
		.INIT('h1)
	) name1298 (
		\sa21_reg[1]/P0001 ,
		_w1829_,
		_w1830_
	);
	LUT2 #(
		.INIT('h2)
	) name1299 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		_w1831_
	);
	LUT2 #(
		.INIT('h1)
	) name1300 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1832_
	);
	LUT2 #(
		.INIT('h4)
	) name1301 (
		\sa21_reg[4]/P0001 ,
		_w1832_,
		_w1833_
	);
	LUT2 #(
		.INIT('h8)
	) name1302 (
		\sa21_reg[4]/P0001 ,
		_w1823_,
		_w1834_
	);
	LUT2 #(
		.INIT('h1)
	) name1303 (
		_w1833_,
		_w1834_,
		_w1835_
	);
	LUT2 #(
		.INIT('h2)
	) name1304 (
		_w1831_,
		_w1835_,
		_w1836_
	);
	LUT2 #(
		.INIT('h8)
	) name1305 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1837_
	);
	LUT2 #(
		.INIT('h8)
	) name1306 (
		_w1799_,
		_w1837_,
		_w1838_
	);
	LUT2 #(
		.INIT('h8)
	) name1307 (
		\sa21_reg[4]/P0001 ,
		_w1838_,
		_w1839_
	);
	LUT2 #(
		.INIT('h2)
	) name1308 (
		\sa21_reg[4]/P0001 ,
		_w1822_,
		_w1840_
	);
	LUT2 #(
		.INIT('h1)
	) name1309 (
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1841_
	);
	LUT2 #(
		.INIT('h2)
	) name1310 (
		_w1787_,
		_w1841_,
		_w1842_
	);
	LUT2 #(
		.INIT('h4)
	) name1311 (
		_w1840_,
		_w1842_,
		_w1843_
	);
	LUT2 #(
		.INIT('h8)
	) name1312 (
		\sa21_reg[4]/P0001 ,
		_w1832_,
		_w1844_
	);
	LUT2 #(
		.INIT('h4)
	) name1313 (
		\sa21_reg[3]/P0001 ,
		_w1844_,
		_w1845_
	);
	LUT2 #(
		.INIT('h1)
	) name1314 (
		_w1839_,
		_w1843_,
		_w1846_
	);
	LUT2 #(
		.INIT('h4)
	) name1315 (
		_w1845_,
		_w1846_,
		_w1847_
	);
	LUT2 #(
		.INIT('h1)
	) name1316 (
		\sa21_reg[2]/P0001 ,
		_w1847_,
		_w1848_
	);
	LUT2 #(
		.INIT('h8)
	) name1317 (
		\sa21_reg[4]/P0001 ,
		_w1749_,
		_w1849_
	);
	LUT2 #(
		.INIT('h1)
	) name1318 (
		_w1785_,
		_w1849_,
		_w1850_
	);
	LUT2 #(
		.INIT('h2)
	) name1319 (
		_w1831_,
		_w1850_,
		_w1851_
	);
	LUT2 #(
		.INIT('h4)
	) name1320 (
		\sa21_reg[2]/P0001 ,
		_w1786_,
		_w1852_
	);
	LUT2 #(
		.INIT('h8)
	) name1321 (
		\sa21_reg[4]/P0001 ,
		_w1837_,
		_w1853_
	);
	LUT2 #(
		.INIT('h2)
	) name1322 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1854_
	);
	LUT2 #(
		.INIT('h8)
	) name1323 (
		_w1853_,
		_w1854_,
		_w1855_
	);
	LUT2 #(
		.INIT('h1)
	) name1324 (
		_w1851_,
		_w1855_,
		_w1856_
	);
	LUT2 #(
		.INIT('h4)
	) name1325 (
		_w1852_,
		_w1856_,
		_w1857_
	);
	LUT2 #(
		.INIT('h2)
	) name1326 (
		\sa21_reg[1]/P0001 ,
		_w1857_,
		_w1858_
	);
	LUT2 #(
		.INIT('h1)
	) name1327 (
		_w1836_,
		_w1848_,
		_w1859_
	);
	LUT2 #(
		.INIT('h4)
	) name1328 (
		_w1830_,
		_w1859_,
		_w1860_
	);
	LUT2 #(
		.INIT('h4)
	) name1329 (
		_w1858_,
		_w1860_,
		_w1861_
	);
	LUT2 #(
		.INIT('h1)
	) name1330 (
		\sa21_reg[0]/P0001 ,
		_w1861_,
		_w1862_
	);
	LUT2 #(
		.INIT('h8)
	) name1331 (
		\sa21_reg[1]/P0001 ,
		\sa21_reg[2]/P0001 ,
		_w1863_
	);
	LUT2 #(
		.INIT('h4)
	) name1332 (
		\sa21_reg[6]/NET0131 ,
		_w1795_,
		_w1864_
	);
	LUT2 #(
		.INIT('h8)
	) name1333 (
		_w1815_,
		_w1841_,
		_w1865_
	);
	LUT2 #(
		.INIT('h2)
	) name1334 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w1866_
	);
	LUT2 #(
		.INIT('h8)
	) name1335 (
		\sa21_reg[5]/P0001 ,
		_w1866_,
		_w1867_
	);
	LUT2 #(
		.INIT('h8)
	) name1336 (
		_w1763_,
		_w1867_,
		_w1868_
	);
	LUT2 #(
		.INIT('h1)
	) name1337 (
		_w1864_,
		_w1865_,
		_w1869_
	);
	LUT2 #(
		.INIT('h4)
	) name1338 (
		_w1868_,
		_w1869_,
		_w1870_
	);
	LUT2 #(
		.INIT('h2)
	) name1339 (
		_w1863_,
		_w1870_,
		_w1871_
	);
	LUT2 #(
		.INIT('h8)
	) name1340 (
		_w1799_,
		_w1832_,
		_w1872_
	);
	LUT2 #(
		.INIT('h8)
	) name1341 (
		_w1758_,
		_w1802_,
		_w1873_
	);
	LUT2 #(
		.INIT('h4)
	) name1342 (
		\sa21_reg[7]/P0001 ,
		_w1873_,
		_w1874_
	);
	LUT2 #(
		.INIT('h1)
	) name1343 (
		_w1872_,
		_w1874_,
		_w1875_
	);
	LUT2 #(
		.INIT('h2)
	) name1344 (
		\sa21_reg[2]/P0001 ,
		_w1875_,
		_w1876_
	);
	LUT2 #(
		.INIT('h4)
	) name1345 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		_w1877_
	);
	LUT2 #(
		.INIT('h8)
	) name1346 (
		_w1792_,
		_w1877_,
		_w1878_
	);
	LUT2 #(
		.INIT('h4)
	) name1347 (
		\sa21_reg[4]/P0001 ,
		_w1745_,
		_w1879_
	);
	LUT2 #(
		.INIT('h4)
	) name1348 (
		\sa21_reg[6]/NET0131 ,
		_w1879_,
		_w1880_
	);
	LUT2 #(
		.INIT('h8)
	) name1349 (
		_w1877_,
		_w1880_,
		_w1881_
	);
	LUT2 #(
		.INIT('h8)
	) name1350 (
		\sa21_reg[1]/P0001 ,
		_w1881_,
		_w1882_
	);
	LUT2 #(
		.INIT('h8)
	) name1351 (
		_w1799_,
		_w1833_,
		_w1883_
	);
	LUT2 #(
		.INIT('h4)
	) name1352 (
		\sa21_reg[5]/P0001 ,
		_w1762_,
		_w1884_
	);
	LUT2 #(
		.INIT('h4)
	) name1353 (
		\sa21_reg[6]/NET0131 ,
		_w1750_,
		_w1885_
	);
	LUT2 #(
		.INIT('h1)
	) name1354 (
		_w1792_,
		_w1884_,
		_w1886_
	);
	LUT2 #(
		.INIT('h4)
	) name1355 (
		_w1885_,
		_w1886_,
		_w1887_
	);
	LUT2 #(
		.INIT('h1)
	) name1356 (
		\sa21_reg[2]/P0001 ,
		_w1887_,
		_w1888_
	);
	LUT2 #(
		.INIT('h4)
	) name1357 (
		\sa21_reg[6]/NET0131 ,
		_w1803_,
		_w1889_
	);
	LUT2 #(
		.INIT('h4)
	) name1358 (
		\sa21_reg[3]/P0001 ,
		_w1753_,
		_w1890_
	);
	LUT2 #(
		.INIT('h8)
	) name1359 (
		\sa21_reg[5]/P0001 ,
		_w1890_,
		_w1891_
	);
	LUT2 #(
		.INIT('h8)
	) name1360 (
		_w1793_,
		_w1837_,
		_w1892_
	);
	LUT2 #(
		.INIT('h8)
	) name1361 (
		\sa21_reg[2]/P0001 ,
		_w1892_,
		_w1893_
	);
	LUT2 #(
		.INIT('h8)
	) name1362 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		_w1894_
	);
	LUT2 #(
		.INIT('h4)
	) name1363 (
		\sa21_reg[4]/P0001 ,
		_w1894_,
		_w1895_
	);
	LUT2 #(
		.INIT('h8)
	) name1364 (
		_w1841_,
		_w1895_,
		_w1896_
	);
	LUT2 #(
		.INIT('h1)
	) name1365 (
		_w1889_,
		_w1891_,
		_w1897_
	);
	LUT2 #(
		.INIT('h1)
	) name1366 (
		_w1893_,
		_w1896_,
		_w1898_
	);
	LUT2 #(
		.INIT('h8)
	) name1367 (
		_w1897_,
		_w1898_,
		_w1899_
	);
	LUT2 #(
		.INIT('h4)
	) name1368 (
		_w1888_,
		_w1899_,
		_w1900_
	);
	LUT2 #(
		.INIT('h1)
	) name1369 (
		\sa21_reg[1]/P0001 ,
		_w1900_,
		_w1901_
	);
	LUT2 #(
		.INIT('h1)
	) name1370 (
		_w1878_,
		_w1883_,
		_w1902_
	);
	LUT2 #(
		.INIT('h4)
	) name1371 (
		_w1876_,
		_w1902_,
		_w1903_
	);
	LUT2 #(
		.INIT('h4)
	) name1372 (
		_w1882_,
		_w1903_,
		_w1904_
	);
	LUT2 #(
		.INIT('h4)
	) name1373 (
		_w1871_,
		_w1904_,
		_w1905_
	);
	LUT2 #(
		.INIT('h4)
	) name1374 (
		_w1901_,
		_w1905_,
		_w1906_
	);
	LUT2 #(
		.INIT('h4)
	) name1375 (
		_w1862_,
		_w1906_,
		_w1907_
	);
	LUT2 #(
		.INIT('h4)
	) name1376 (
		_w1814_,
		_w1907_,
		_w1908_
	);
	LUT2 #(
		.INIT('h8)
	) name1377 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1909_
	);
	LUT2 #(
		.INIT('h4)
	) name1378 (
		\sa32_reg[7]/P0001 ,
		_w1909_,
		_w1910_
	);
	LUT2 #(
		.INIT('h8)
	) name1379 (
		\sa32_reg[3]/P0001 ,
		_w1910_,
		_w1911_
	);
	LUT2 #(
		.INIT('h8)
	) name1380 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w1912_
	);
	LUT2 #(
		.INIT('h1)
	) name1381 (
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1913_
	);
	LUT2 #(
		.INIT('h8)
	) name1382 (
		_w1912_,
		_w1913_,
		_w1914_
	);
	LUT2 #(
		.INIT('h4)
	) name1383 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1915_
	);
	LUT2 #(
		.INIT('h4)
	) name1384 (
		\sa32_reg[4]/P0001 ,
		_w1915_,
		_w1916_
	);
	LUT2 #(
		.INIT('h1)
	) name1385 (
		_w1914_,
		_w1916_,
		_w1917_
	);
	LUT2 #(
		.INIT('h2)
	) name1386 (
		\sa32_reg[2]/P0001 ,
		_w1917_,
		_w1918_
	);
	LUT2 #(
		.INIT('h4)
	) name1387 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w1919_
	);
	LUT2 #(
		.INIT('h8)
	) name1388 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1920_
	);
	LUT2 #(
		.INIT('h8)
	) name1389 (
		_w1919_,
		_w1920_,
		_w1921_
	);
	LUT2 #(
		.INIT('h8)
	) name1390 (
		\sa32_reg[6]/NET0131 ,
		_w1921_,
		_w1922_
	);
	LUT2 #(
		.INIT('h4)
	) name1391 (
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1923_
	);
	LUT2 #(
		.INIT('h2)
	) name1392 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		_w1924_
	);
	LUT2 #(
		.INIT('h8)
	) name1393 (
		_w1923_,
		_w1924_,
		_w1925_
	);
	LUT2 #(
		.INIT('h1)
	) name1394 (
		_w1910_,
		_w1925_,
		_w1926_
	);
	LUT2 #(
		.INIT('h1)
	) name1395 (
		\sa32_reg[2]/P0001 ,
		_w1926_,
		_w1927_
	);
	LUT2 #(
		.INIT('h1)
	) name1396 (
		\sa32_reg[1]/P0001 ,
		_w1911_,
		_w1928_
	);
	LUT2 #(
		.INIT('h4)
	) name1397 (
		_w1922_,
		_w1928_,
		_w1929_
	);
	LUT2 #(
		.INIT('h1)
	) name1398 (
		_w1918_,
		_w1927_,
		_w1930_
	);
	LUT2 #(
		.INIT('h8)
	) name1399 (
		_w1929_,
		_w1930_,
		_w1931_
	);
	LUT2 #(
		.INIT('h8)
	) name1400 (
		\sa32_reg[3]/P0001 ,
		_w1923_,
		_w1932_
	);
	LUT2 #(
		.INIT('h4)
	) name1401 (
		\sa32_reg[4]/P0001 ,
		_w1932_,
		_w1933_
	);
	LUT2 #(
		.INIT('h2)
	) name1402 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1934_
	);
	LUT2 #(
		.INIT('h8)
	) name1403 (
		_w1912_,
		_w1934_,
		_w1935_
	);
	LUT2 #(
		.INIT('h4)
	) name1404 (
		\sa32_reg[6]/NET0131 ,
		_w1935_,
		_w1936_
	);
	LUT2 #(
		.INIT('h4)
	) name1405 (
		\sa32_reg[5]/P0001 ,
		_w1913_,
		_w1937_
	);
	LUT2 #(
		.INIT('h8)
	) name1406 (
		_w1919_,
		_w1937_,
		_w1938_
	);
	LUT2 #(
		.INIT('h2)
	) name1407 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1939_
	);
	LUT2 #(
		.INIT('h8)
	) name1408 (
		_w1919_,
		_w1939_,
		_w1940_
	);
	LUT2 #(
		.INIT('h8)
	) name1409 (
		\sa32_reg[7]/P0001 ,
		_w1940_,
		_w1941_
	);
	LUT2 #(
		.INIT('h2)
	) name1410 (
		\sa32_reg[1]/P0001 ,
		_w1933_,
		_w1942_
	);
	LUT2 #(
		.INIT('h1)
	) name1411 (
		_w1936_,
		_w1938_,
		_w1943_
	);
	LUT2 #(
		.INIT('h4)
	) name1412 (
		_w1941_,
		_w1943_,
		_w1944_
	);
	LUT2 #(
		.INIT('h8)
	) name1413 (
		_w1942_,
		_w1944_,
		_w1945_
	);
	LUT2 #(
		.INIT('h1)
	) name1414 (
		_w1931_,
		_w1945_,
		_w1946_
	);
	LUT2 #(
		.INIT('h8)
	) name1415 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1947_
	);
	LUT2 #(
		.INIT('h1)
	) name1416 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1948_
	);
	LUT2 #(
		.INIT('h8)
	) name1417 (
		_w1947_,
		_w1948_,
		_w1949_
	);
	LUT2 #(
		.INIT('h1)
	) name1418 (
		_w1911_,
		_w1949_,
		_w1950_
	);
	LUT2 #(
		.INIT('h2)
	) name1419 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w1951_
	);
	LUT2 #(
		.INIT('h8)
	) name1420 (
		\sa32_reg[5]/P0001 ,
		_w1951_,
		_w1952_
	);
	LUT2 #(
		.INIT('h8)
	) name1421 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1953_
	);
	LUT2 #(
		.INIT('h4)
	) name1422 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1954_
	);
	LUT2 #(
		.INIT('h1)
	) name1423 (
		\sa32_reg[5]/P0001 ,
		_w1954_,
		_w1955_
	);
	LUT2 #(
		.INIT('h4)
	) name1424 (
		_w1953_,
		_w1955_,
		_w1956_
	);
	LUT2 #(
		.INIT('h1)
	) name1425 (
		_w1952_,
		_w1956_,
		_w1957_
	);
	LUT2 #(
		.INIT('h2)
	) name1426 (
		\sa32_reg[1]/P0001 ,
		_w1957_,
		_w1958_
	);
	LUT2 #(
		.INIT('h4)
	) name1427 (
		\sa32_reg[4]/P0001 ,
		_w1934_,
		_w1959_
	);
	LUT2 #(
		.INIT('h2)
	) name1428 (
		_w1950_,
		_w1959_,
		_w1960_
	);
	LUT2 #(
		.INIT('h4)
	) name1429 (
		_w1958_,
		_w1960_,
		_w1961_
	);
	LUT2 #(
		.INIT('h1)
	) name1430 (
		\sa32_reg[2]/P0001 ,
		_w1961_,
		_w1962_
	);
	LUT2 #(
		.INIT('h8)
	) name1431 (
		_w1915_,
		_w1953_,
		_w1963_
	);
	LUT2 #(
		.INIT('h4)
	) name1432 (
		\sa32_reg[2]/P0001 ,
		_w1963_,
		_w1964_
	);
	LUT2 #(
		.INIT('h4)
	) name1433 (
		\sa32_reg[3]/P0001 ,
		_w1915_,
		_w1965_
	);
	LUT2 #(
		.INIT('h8)
	) name1434 (
		_w1948_,
		_w1965_,
		_w1966_
	);
	LUT2 #(
		.INIT('h1)
	) name1435 (
		_w1922_,
		_w1966_,
		_w1967_
	);
	LUT2 #(
		.INIT('h2)
	) name1436 (
		\sa32_reg[2]/P0001 ,
		_w1967_,
		_w1968_
	);
	LUT2 #(
		.INIT('h4)
	) name1437 (
		\sa32_reg[7]/P0001 ,
		_w1947_,
		_w1969_
	);
	LUT2 #(
		.INIT('h4)
	) name1438 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		_w1970_
	);
	LUT2 #(
		.INIT('h8)
	) name1439 (
		_w1969_,
		_w1970_,
		_w1971_
	);
	LUT2 #(
		.INIT('h1)
	) name1440 (
		_w1964_,
		_w1971_,
		_w1972_
	);
	LUT2 #(
		.INIT('h4)
	) name1441 (
		_w1968_,
		_w1972_,
		_w1973_
	);
	LUT2 #(
		.INIT('h4)
	) name1442 (
		_w1946_,
		_w1973_,
		_w1974_
	);
	LUT2 #(
		.INIT('h4)
	) name1443 (
		_w1962_,
		_w1974_,
		_w1975_
	);
	LUT2 #(
		.INIT('h2)
	) name1444 (
		\sa32_reg[0]/P0002 ,
		_w1975_,
		_w1976_
	);
	LUT2 #(
		.INIT('h8)
	) name1445 (
		\sa32_reg[3]/P0001 ,
		_w1920_,
		_w1977_
	);
	LUT2 #(
		.INIT('h8)
	) name1446 (
		\sa32_reg[4]/P0001 ,
		_w1910_,
		_w1978_
	);
	LUT2 #(
		.INIT('h1)
	) name1447 (
		_w1977_,
		_w1978_,
		_w1979_
	);
	LUT2 #(
		.INIT('h2)
	) name1448 (
		\sa32_reg[2]/P0001 ,
		_w1979_,
		_w1980_
	);
	LUT2 #(
		.INIT('h2)
	) name1449 (
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1981_
	);
	LUT2 #(
		.INIT('h4)
	) name1450 (
		\sa32_reg[3]/P0001 ,
		_w1981_,
		_w1982_
	);
	LUT2 #(
		.INIT('h4)
	) name1451 (
		\sa32_reg[4]/P0001 ,
		_w1982_,
		_w1983_
	);
	LUT2 #(
		.INIT('h1)
	) name1452 (
		_w1932_,
		_w1940_,
		_w1984_
	);
	LUT2 #(
		.INIT('h4)
	) name1453 (
		_w1983_,
		_w1984_,
		_w1985_
	);
	LUT2 #(
		.INIT('h1)
	) name1454 (
		\sa32_reg[2]/P0001 ,
		_w1985_,
		_w1986_
	);
	LUT2 #(
		.INIT('h8)
	) name1455 (
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1987_
	);
	LUT2 #(
		.INIT('h4)
	) name1456 (
		\sa32_reg[5]/P0001 ,
		_w1987_,
		_w1988_
	);
	LUT2 #(
		.INIT('h4)
	) name1457 (
		\sa32_reg[3]/P0001 ,
		_w1988_,
		_w1989_
	);
	LUT2 #(
		.INIT('h1)
	) name1458 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1990_
	);
	LUT2 #(
		.INIT('h8)
	) name1459 (
		\sa32_reg[3]/P0001 ,
		_w1990_,
		_w1991_
	);
	LUT2 #(
		.INIT('h4)
	) name1460 (
		\sa32_reg[7]/P0001 ,
		_w1991_,
		_w1992_
	);
	LUT2 #(
		.INIT('h8)
	) name1461 (
		_w1912_,
		_w1920_,
		_w1993_
	);
	LUT2 #(
		.INIT('h8)
	) name1462 (
		_w1923_,
		_w1970_,
		_w1994_
	);
	LUT2 #(
		.INIT('h1)
	) name1463 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w1995_
	);
	LUT2 #(
		.INIT('h8)
	) name1464 (
		_w1910_,
		_w1995_,
		_w1996_
	);
	LUT2 #(
		.INIT('h1)
	) name1465 (
		_w1993_,
		_w1994_,
		_w1997_
	);
	LUT2 #(
		.INIT('h4)
	) name1466 (
		_w1989_,
		_w1997_,
		_w1998_
	);
	LUT2 #(
		.INIT('h1)
	) name1467 (
		_w1992_,
		_w1996_,
		_w1999_
	);
	LUT2 #(
		.INIT('h8)
	) name1468 (
		_w1998_,
		_w1999_,
		_w2000_
	);
	LUT2 #(
		.INIT('h4)
	) name1469 (
		_w1980_,
		_w2000_,
		_w2001_
	);
	LUT2 #(
		.INIT('h4)
	) name1470 (
		_w1986_,
		_w2001_,
		_w2002_
	);
	LUT2 #(
		.INIT('h2)
	) name1471 (
		\sa32_reg[1]/P0001 ,
		_w2002_,
		_w2003_
	);
	LUT2 #(
		.INIT('h4)
	) name1472 (
		\sa32_reg[6]/NET0131 ,
		_w1951_,
		_w2004_
	);
	LUT2 #(
		.INIT('h8)
	) name1473 (
		\sa32_reg[2]/P0001 ,
		_w2004_,
		_w2005_
	);
	LUT2 #(
		.INIT('h8)
	) name1474 (
		_w1919_,
		_w1923_,
		_w2006_
	);
	LUT2 #(
		.INIT('h1)
	) name1475 (
		_w2005_,
		_w2006_,
		_w2007_
	);
	LUT2 #(
		.INIT('h1)
	) name1476 (
		\sa32_reg[5]/P0001 ,
		_w2007_,
		_w2008_
	);
	LUT2 #(
		.INIT('h4)
	) name1477 (
		\sa32_reg[3]/P0001 ,
		_w1937_,
		_w2009_
	);
	LUT2 #(
		.INIT('h8)
	) name1478 (
		\sa32_reg[2]/P0001 ,
		_w2009_,
		_w2010_
	);
	LUT2 #(
		.INIT('h8)
	) name1479 (
		\sa32_reg[7]/P0001 ,
		_w1909_,
		_w2011_
	);
	LUT2 #(
		.INIT('h4)
	) name1480 (
		\sa32_reg[3]/P0001 ,
		_w2011_,
		_w2012_
	);
	LUT2 #(
		.INIT('h4)
	) name1481 (
		\sa32_reg[4]/P0001 ,
		_w2012_,
		_w2013_
	);
	LUT2 #(
		.INIT('h1)
	) name1482 (
		_w2010_,
		_w2013_,
		_w2014_
	);
	LUT2 #(
		.INIT('h4)
	) name1483 (
		_w2008_,
		_w2014_,
		_w2015_
	);
	LUT2 #(
		.INIT('h1)
	) name1484 (
		\sa32_reg[1]/P0001 ,
		_w2015_,
		_w2016_
	);
	LUT2 #(
		.INIT('h2)
	) name1485 (
		\sa32_reg[6]/NET0131 ,
		_w1924_,
		_w2017_
	);
	LUT2 #(
		.INIT('h2)
	) name1486 (
		_w1948_,
		_w2017_,
		_w2018_
	);
	LUT2 #(
		.INIT('h4)
	) name1487 (
		\sa32_reg[5]/P0001 ,
		_w1981_,
		_w2019_
	);
	LUT2 #(
		.INIT('h8)
	) name1488 (
		_w1919_,
		_w2019_,
		_w2020_
	);
	LUT2 #(
		.INIT('h1)
	) name1489 (
		_w1993_,
		_w2018_,
		_w2021_
	);
	LUT2 #(
		.INIT('h4)
	) name1490 (
		_w2020_,
		_w2021_,
		_w2022_
	);
	LUT2 #(
		.INIT('h2)
	) name1491 (
		\sa32_reg[2]/P0001 ,
		_w2022_,
		_w2023_
	);
	LUT2 #(
		.INIT('h8)
	) name1492 (
		_w1939_,
		_w1953_,
		_w2024_
	);
	LUT2 #(
		.INIT('h4)
	) name1493 (
		\sa32_reg[2]/P0001 ,
		_w2024_,
		_w2025_
	);
	LUT2 #(
		.INIT('h4)
	) name1494 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		_w2026_
	);
	LUT2 #(
		.INIT('h1)
	) name1495 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w2027_
	);
	LUT2 #(
		.INIT('h8)
	) name1496 (
		\sa32_reg[4]/P0001 ,
		_w2027_,
		_w2028_
	);
	LUT2 #(
		.INIT('h8)
	) name1497 (
		_w2026_,
		_w2028_,
		_w2029_
	);
	LUT2 #(
		.INIT('h1)
	) name1498 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w2030_
	);
	LUT2 #(
		.INIT('h8)
	) name1499 (
		_w1988_,
		_w2030_,
		_w2031_
	);
	LUT2 #(
		.INIT('h1)
	) name1500 (
		_w2029_,
		_w2031_,
		_w2032_
	);
	LUT2 #(
		.INIT('h8)
	) name1501 (
		_w1948_,
		_w1990_,
		_w2033_
	);
	LUT2 #(
		.INIT('h1)
	) name1502 (
		_w2025_,
		_w2033_,
		_w2034_
	);
	LUT2 #(
		.INIT('h8)
	) name1503 (
		_w2032_,
		_w2034_,
		_w2035_
	);
	LUT2 #(
		.INIT('h4)
	) name1504 (
		_w2023_,
		_w2035_,
		_w2036_
	);
	LUT2 #(
		.INIT('h4)
	) name1505 (
		_w2016_,
		_w2036_,
		_w2037_
	);
	LUT2 #(
		.INIT('h4)
	) name1506 (
		_w2003_,
		_w2037_,
		_w2038_
	);
	LUT2 #(
		.INIT('h1)
	) name1507 (
		\sa32_reg[0]/P0002 ,
		_w2038_,
		_w2039_
	);
	LUT2 #(
		.INIT('h8)
	) name1508 (
		_w1913_,
		_w1995_,
		_w2040_
	);
	LUT2 #(
		.INIT('h4)
	) name1509 (
		\sa32_reg[5]/P0001 ,
		_w1923_,
		_w2041_
	);
	LUT2 #(
		.INIT('h1)
	) name1510 (
		_w2019_,
		_w2041_,
		_w2042_
	);
	LUT2 #(
		.INIT('h1)
	) name1511 (
		\sa32_reg[3]/P0001 ,
		_w2011_,
		_w2043_
	);
	LUT2 #(
		.INIT('h8)
	) name1512 (
		_w2042_,
		_w2043_,
		_w2044_
	);
	LUT2 #(
		.INIT('h2)
	) name1513 (
		\sa32_reg[3]/P0001 ,
		_w1939_,
		_w2045_
	);
	LUT2 #(
		.INIT('h8)
	) name1514 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w2046_
	);
	LUT2 #(
		.INIT('h4)
	) name1515 (
		_w2045_,
		_w2046_,
		_w2047_
	);
	LUT2 #(
		.INIT('h4)
	) name1516 (
		_w2044_,
		_w2047_,
		_w2048_
	);
	LUT2 #(
		.INIT('h4)
	) name1517 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w2049_
	);
	LUT2 #(
		.INIT('h4)
	) name1518 (
		\sa32_reg[3]/P0001 ,
		_w2049_,
		_w2050_
	);
	LUT2 #(
		.INIT('h8)
	) name1519 (
		\sa32_reg[5]/P0001 ,
		_w2050_,
		_w2051_
	);
	LUT2 #(
		.INIT('h8)
	) name1520 (
		\sa32_reg[6]/NET0131 ,
		_w1935_,
		_w2052_
	);
	LUT2 #(
		.INIT('h1)
	) name1521 (
		_w1963_,
		_w2051_,
		_w2053_
	);
	LUT2 #(
		.INIT('h4)
	) name1522 (
		_w2052_,
		_w2053_,
		_w2054_
	);
	LUT2 #(
		.INIT('h1)
	) name1523 (
		\sa32_reg[2]/P0001 ,
		_w2054_,
		_w2055_
	);
	LUT2 #(
		.INIT('h1)
	) name1524 (
		_w2040_,
		_w2048_,
		_w2056_
	);
	LUT2 #(
		.INIT('h4)
	) name1525 (
		_w2055_,
		_w2056_,
		_w2057_
	);
	LUT2 #(
		.INIT('h1)
	) name1526 (
		\sa32_reg[1]/P0001 ,
		_w2057_,
		_w2058_
	);
	LUT2 #(
		.INIT('h8)
	) name1527 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		_w2059_
	);
	LUT2 #(
		.INIT('h8)
	) name1528 (
		\sa32_reg[5]/P0001 ,
		_w1913_,
		_w2060_
	);
	LUT2 #(
		.INIT('h8)
	) name1529 (
		_w2059_,
		_w2060_,
		_w2061_
	);
	LUT2 #(
		.INIT('h8)
	) name1530 (
		\sa32_reg[4]/P0001 ,
		_w2061_,
		_w2062_
	);
	LUT2 #(
		.INIT('h8)
	) name1531 (
		_w1934_,
		_w2004_,
		_w2063_
	);
	LUT2 #(
		.INIT('h1)
	) name1532 (
		_w1989_,
		_w2063_,
		_w2064_
	);
	LUT2 #(
		.INIT('h1)
	) name1533 (
		\sa32_reg[2]/P0001 ,
		_w2064_,
		_w2065_
	);
	LUT2 #(
		.INIT('h8)
	) name1534 (
		_w1937_,
		_w1951_,
		_w2066_
	);
	LUT2 #(
		.INIT('h8)
	) name1535 (
		\sa32_reg[2]/P0001 ,
		_w1981_,
		_w2067_
	);
	LUT2 #(
		.INIT('h8)
	) name1536 (
		\sa32_reg[5]/P0001 ,
		_w2067_,
		_w2068_
	);
	LUT2 #(
		.INIT('h8)
	) name1537 (
		_w1919_,
		_w2068_,
		_w2069_
	);
	LUT2 #(
		.INIT('h1)
	) name1538 (
		_w2025_,
		_w2066_,
		_w2070_
	);
	LUT2 #(
		.INIT('h4)
	) name1539 (
		_w2069_,
		_w2070_,
		_w2071_
	);
	LUT2 #(
		.INIT('h2)
	) name1540 (
		\sa32_reg[1]/P0001 ,
		_w2071_,
		_w2072_
	);
	LUT2 #(
		.INIT('h1)
	) name1541 (
		_w2062_,
		_w2065_,
		_w2073_
	);
	LUT2 #(
		.INIT('h4)
	) name1542 (
		_w2072_,
		_w2073_,
		_w2074_
	);
	LUT2 #(
		.INIT('h4)
	) name1543 (
		_w2058_,
		_w2074_,
		_w2075_
	);
	LUT2 #(
		.INIT('h4)
	) name1544 (
		_w1976_,
		_w2075_,
		_w2076_
	);
	LUT2 #(
		.INIT('h4)
	) name1545 (
		_w2039_,
		_w2076_,
		_w2077_
	);
	LUT2 #(
		.INIT('h2)
	) name1546 (
		\u0_w_reg[3][6]/P0001 ,
		_w2077_,
		_w2078_
	);
	LUT2 #(
		.INIT('h4)
	) name1547 (
		\u0_w_reg[3][6]/P0001 ,
		_w2077_,
		_w2079_
	);
	LUT2 #(
		.INIT('h1)
	) name1548 (
		_w2078_,
		_w2079_,
		_w2080_
	);
	LUT2 #(
		.INIT('h8)
	) name1549 (
		_w1908_,
		_w2080_,
		_w2081_
	);
	LUT2 #(
		.INIT('h1)
	) name1550 (
		_w1908_,
		_w2080_,
		_w2082_
	);
	LUT2 #(
		.INIT('h1)
	) name1551 (
		_w2081_,
		_w2082_,
		_w2083_
	);
	LUT2 #(
		.INIT('h4)
	) name1552 (
		_w1744_,
		_w2083_,
		_w2084_
	);
	LUT2 #(
		.INIT('h2)
	) name1553 (
		_w1744_,
		_w2083_,
		_w2085_
	);
	LUT2 #(
		.INIT('h1)
	) name1554 (
		\ld_r_reg/P0001 ,
		_w2084_,
		_w2086_
	);
	LUT2 #(
		.INIT('h4)
	) name1555 (
		_w2085_,
		_w2086_,
		_w2087_
	);
	LUT2 #(
		.INIT('h2)
	) name1556 (
		\text_in_r_reg[6]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w2088_
	);
	LUT2 #(
		.INIT('h4)
	) name1557 (
		\text_in_r_reg[6]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w2089_
	);
	LUT2 #(
		.INIT('h2)
	) name1558 (
		\ld_r_reg/P0001 ,
		_w2088_,
		_w2090_
	);
	LUT2 #(
		.INIT('h4)
	) name1559 (
		_w2089_,
		_w2090_,
		_w2091_
	);
	LUT2 #(
		.INIT('h1)
	) name1560 (
		_w2087_,
		_w2091_,
		_w2092_
	);
	LUT2 #(
		.INIT('h8)
	) name1561 (
		_w1600_,
		_w1607_,
		_w2093_
	);
	LUT2 #(
		.INIT('h1)
	) name1562 (
		_w1713_,
		_w2093_,
		_w2094_
	);
	LUT2 #(
		.INIT('h2)
	) name1563 (
		_w1582_,
		_w1637_,
		_w2095_
	);
	LUT2 #(
		.INIT('h2)
	) name1564 (
		_w2094_,
		_w2095_,
		_w2096_
	);
	LUT2 #(
		.INIT('h2)
	) name1565 (
		_w1666_,
		_w2096_,
		_w2097_
	);
	LUT2 #(
		.INIT('h8)
	) name1566 (
		\sa10_reg[4]/P0001 ,
		_w1650_,
		_w2098_
	);
	LUT2 #(
		.INIT('h1)
	) name1567 (
		_w1607_,
		_w2098_,
		_w2099_
	);
	LUT2 #(
		.INIT('h2)
	) name1568 (
		\sa10_reg[7]/NET0131 ,
		_w2099_,
		_w2100_
	);
	LUT2 #(
		.INIT('h8)
	) name1569 (
		_w1582_,
		_w1586_,
		_w2101_
	);
	LUT2 #(
		.INIT('h1)
	) name1570 (
		_w2100_,
		_w2101_,
		_w2102_
	);
	LUT2 #(
		.INIT('h1)
	) name1571 (
		\sa10_reg[3]/P0001 ,
		_w2102_,
		_w2103_
	);
	LUT2 #(
		.INIT('h1)
	) name1572 (
		_w1609_,
		_w1682_,
		_w2104_
	);
	LUT2 #(
		.INIT('h4)
	) name1573 (
		_w2103_,
		_w2104_,
		_w2105_
	);
	LUT2 #(
		.INIT('h2)
	) name1574 (
		\sa10_reg[2]/P0001 ,
		_w2105_,
		_w2106_
	);
	LUT2 #(
		.INIT('h1)
	) name1575 (
		_w2097_,
		_w2106_,
		_w2107_
	);
	LUT2 #(
		.INIT('h2)
	) name1576 (
		\sa10_reg[1]/P0001 ,
		_w2107_,
		_w2108_
	);
	LUT2 #(
		.INIT('h4)
	) name1577 (
		\sa10_reg[2]/P0001 ,
		_w1637_,
		_w2109_
	);
	LUT2 #(
		.INIT('h8)
	) name1578 (
		\sa10_reg[2]/P0001 ,
		_w1594_,
		_w2110_
	);
	LUT2 #(
		.INIT('h8)
	) name1579 (
		_w1608_,
		_w2110_,
		_w2111_
	);
	LUT2 #(
		.INIT('h2)
	) name1580 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w2112_
	);
	LUT2 #(
		.INIT('h8)
	) name1581 (
		_w1600_,
		_w2112_,
		_w2113_
	);
	LUT2 #(
		.INIT('h1)
	) name1582 (
		_w1628_,
		_w2109_,
		_w2114_
	);
	LUT2 #(
		.INIT('h4)
	) name1583 (
		_w2113_,
		_w2114_,
		_w2115_
	);
	LUT2 #(
		.INIT('h4)
	) name1584 (
		_w2111_,
		_w2115_,
		_w2116_
	);
	LUT2 #(
		.INIT('h1)
	) name1585 (
		\sa10_reg[1]/P0001 ,
		_w2116_,
		_w2117_
	);
	LUT2 #(
		.INIT('h8)
	) name1586 (
		_w1585_,
		_w1612_,
		_w2118_
	);
	LUT2 #(
		.INIT('h8)
	) name1587 (
		\sa10_reg[5]/P0001 ,
		_w1703_,
		_w2119_
	);
	LUT2 #(
		.INIT('h1)
	) name1588 (
		_w1602_,
		_w2118_,
		_w2120_
	);
	LUT2 #(
		.INIT('h4)
	) name1589 (
		_w2119_,
		_w2120_,
		_w2121_
	);
	LUT2 #(
		.INIT('h2)
	) name1590 (
		_w1664_,
		_w2121_,
		_w2122_
	);
	LUT2 #(
		.INIT('h8)
	) name1591 (
		_w1629_,
		_w1668_,
		_w2123_
	);
	LUT2 #(
		.INIT('h1)
	) name1592 (
		_w1591_,
		_w2123_,
		_w2124_
	);
	LUT2 #(
		.INIT('h1)
	) name1593 (
		_w1683_,
		_w1704_,
		_w2125_
	);
	LUT2 #(
		.INIT('h8)
	) name1594 (
		_w2124_,
		_w2125_,
		_w2126_
	);
	LUT2 #(
		.INIT('h1)
	) name1595 (
		\sa10_reg[2]/P0001 ,
		_w2126_,
		_w2127_
	);
	LUT2 #(
		.INIT('h8)
	) name1596 (
		_w1583_,
		_w1672_,
		_w2128_
	);
	LUT2 #(
		.INIT('h2)
	) name1597 (
		\sa10_reg[2]/P0001 ,
		_w2128_,
		_w2129_
	);
	LUT2 #(
		.INIT('h8)
	) name1598 (
		_w1593_,
		_w1598_,
		_w2130_
	);
	LUT2 #(
		.INIT('h1)
	) name1599 (
		\sa10_reg[2]/P0001 ,
		_w2130_,
		_w2131_
	);
	LUT2 #(
		.INIT('h4)
	) name1600 (
		_w1630_,
		_w2131_,
		_w2132_
	);
	LUT2 #(
		.INIT('h1)
	) name1601 (
		_w2129_,
		_w2132_,
		_w2133_
	);
	LUT2 #(
		.INIT('h1)
	) name1602 (
		_w1674_,
		_w1700_,
		_w2134_
	);
	LUT2 #(
		.INIT('h4)
	) name1603 (
		_w2133_,
		_w2134_,
		_w2135_
	);
	LUT2 #(
		.INIT('h2)
	) name1604 (
		\sa10_reg[1]/P0001 ,
		_w2135_,
		_w2136_
	);
	LUT2 #(
		.INIT('h1)
	) name1605 (
		_w2117_,
		_w2122_,
		_w2137_
	);
	LUT2 #(
		.INIT('h4)
	) name1606 (
		_w2127_,
		_w2137_,
		_w2138_
	);
	LUT2 #(
		.INIT('h4)
	) name1607 (
		_w2136_,
		_w2138_,
		_w2139_
	);
	LUT2 #(
		.INIT('h1)
	) name1608 (
		\sa10_reg[0]/P0001 ,
		_w2139_,
		_w2140_
	);
	LUT2 #(
		.INIT('h8)
	) name1609 (
		_w1669_,
		_w1722_,
		_w2141_
	);
	LUT2 #(
		.INIT('h1)
	) name1610 (
		\sa10_reg[2]/P0001 ,
		_w1582_,
		_w2142_
	);
	LUT2 #(
		.INIT('h2)
	) name1611 (
		\sa10_reg[5]/P0001 ,
		_w1637_,
		_w2143_
	);
	LUT2 #(
		.INIT('h1)
	) name1612 (
		_w1653_,
		_w2143_,
		_w2144_
	);
	LUT2 #(
		.INIT('h2)
	) name1613 (
		_w2142_,
		_w2144_,
		_w2145_
	);
	LUT2 #(
		.INIT('h8)
	) name1614 (
		_w1582_,
		_w1627_,
		_w2146_
	);
	LUT2 #(
		.INIT('h8)
	) name1615 (
		_w1593_,
		_w1633_,
		_w2147_
	);
	LUT2 #(
		.INIT('h8)
	) name1616 (
		\sa10_reg[6]/NET0131 ,
		_w1656_,
		_w2148_
	);
	LUT2 #(
		.INIT('h1)
	) name1617 (
		_w2146_,
		_w2147_,
		_w2149_
	);
	LUT2 #(
		.INIT('h4)
	) name1618 (
		_w2141_,
		_w2149_,
		_w2150_
	);
	LUT2 #(
		.INIT('h4)
	) name1619 (
		_w2148_,
		_w2150_,
		_w2151_
	);
	LUT2 #(
		.INIT('h4)
	) name1620 (
		_w2145_,
		_w2151_,
		_w2152_
	);
	LUT2 #(
		.INIT('h1)
	) name1621 (
		\sa10_reg[1]/P0001 ,
		_w2152_,
		_w2153_
	);
	LUT2 #(
		.INIT('h8)
	) name1622 (
		_w1608_,
		_w1633_,
		_w2154_
	);
	LUT2 #(
		.INIT('h4)
	) name1623 (
		\sa10_reg[6]/NET0131 ,
		_w2154_,
		_w2155_
	);
	LUT2 #(
		.INIT('h8)
	) name1624 (
		_w1619_,
		_w1672_,
		_w2156_
	);
	LUT2 #(
		.INIT('h1)
	) name1625 (
		_w2155_,
		_w2156_,
		_w2157_
	);
	LUT2 #(
		.INIT('h2)
	) name1626 (
		\sa10_reg[1]/P0001 ,
		_w2157_,
		_w2158_
	);
	LUT2 #(
		.INIT('h8)
	) name1627 (
		_w1672_,
		_w1715_,
		_w2159_
	);
	LUT2 #(
		.INIT('h8)
	) name1628 (
		\sa10_reg[5]/P0001 ,
		_w1656_,
		_w2160_
	);
	LUT2 #(
		.INIT('h8)
	) name1629 (
		\sa10_reg[4]/P0001 ,
		_w2147_,
		_w2161_
	);
	LUT2 #(
		.INIT('h2)
	) name1630 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w2162_
	);
	LUT2 #(
		.INIT('h8)
	) name1631 (
		\sa10_reg[6]/NET0131 ,
		_w2162_,
		_w2163_
	);
	LUT2 #(
		.INIT('h1)
	) name1632 (
		_w1698_,
		_w2163_,
		_w2164_
	);
	LUT2 #(
		.INIT('h8)
	) name1633 (
		_w2099_,
		_w2164_,
		_w2165_
	);
	LUT2 #(
		.INIT('h2)
	) name1634 (
		_w1697_,
		_w2165_,
		_w2166_
	);
	LUT2 #(
		.INIT('h8)
	) name1635 (
		_w1590_,
		_w1607_,
		_w2167_
	);
	LUT2 #(
		.INIT('h8)
	) name1636 (
		\sa10_reg[5]/P0001 ,
		_w1636_,
		_w2168_
	);
	LUT2 #(
		.INIT('h1)
	) name1637 (
		_w1584_,
		_w2167_,
		_w2169_
	);
	LUT2 #(
		.INIT('h4)
	) name1638 (
		_w2168_,
		_w2169_,
		_w2170_
	);
	LUT2 #(
		.INIT('h2)
	) name1639 (
		\sa10_reg[2]/P0001 ,
		_w2170_,
		_w2171_
	);
	LUT2 #(
		.INIT('h1)
	) name1640 (
		_w2159_,
		_w2160_,
		_w2172_
	);
	LUT2 #(
		.INIT('h4)
	) name1641 (
		_w2161_,
		_w2172_,
		_w2173_
	);
	LUT2 #(
		.INIT('h4)
	) name1642 (
		_w2158_,
		_w2173_,
		_w2174_
	);
	LUT2 #(
		.INIT('h1)
	) name1643 (
		_w2166_,
		_w2171_,
		_w2175_
	);
	LUT2 #(
		.INIT('h8)
	) name1644 (
		_w2174_,
		_w2175_,
		_w2176_
	);
	LUT2 #(
		.INIT('h4)
	) name1645 (
		_w2153_,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h2)
	) name1646 (
		\sa10_reg[0]/P0001 ,
		_w2177_,
		_w2178_
	);
	LUT2 #(
		.INIT('h4)
	) name1647 (
		\sa10_reg[7]/NET0131 ,
		_w1711_,
		_w2179_
	);
	LUT2 #(
		.INIT('h4)
	) name1648 (
		\sa10_reg[6]/NET0131 ,
		_w1606_,
		_w2180_
	);
	LUT2 #(
		.INIT('h1)
	) name1649 (
		_w2179_,
		_w2180_,
		_w2181_
	);
	LUT2 #(
		.INIT('h1)
	) name1650 (
		\sa10_reg[2]/P0001 ,
		_w2181_,
		_w2182_
	);
	LUT2 #(
		.INIT('h4)
	) name1651 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[2]/P0001 ,
		_w2183_
	);
	LUT2 #(
		.INIT('h8)
	) name1652 (
		_w1583_,
		_w1585_,
		_w2184_
	);
	LUT2 #(
		.INIT('h8)
	) name1653 (
		_w1598_,
		_w1614_,
		_w2185_
	);
	LUT2 #(
		.INIT('h1)
	) name1654 (
		_w2184_,
		_w2185_,
		_w2186_
	);
	LUT2 #(
		.INIT('h4)
	) name1655 (
		_w2156_,
		_w2186_,
		_w2187_
	);
	LUT2 #(
		.INIT('h2)
	) name1656 (
		_w2183_,
		_w2187_,
		_w2188_
	);
	LUT2 #(
		.INIT('h8)
	) name1657 (
		_w1583_,
		_w1626_,
		_w2189_
	);
	LUT2 #(
		.INIT('h2)
	) name1658 (
		\sa10_reg[2]/P0001 ,
		_w2189_,
		_w2190_
	);
	LUT2 #(
		.INIT('h1)
	) name1659 (
		_w1671_,
		_w2189_,
		_w2191_
	);
	LUT2 #(
		.INIT('h8)
	) name1660 (
		_w2124_,
		_w2191_,
		_w2192_
	);
	LUT2 #(
		.INIT('h1)
	) name1661 (
		\sa10_reg[1]/P0001 ,
		_w2190_,
		_w2193_
	);
	LUT2 #(
		.INIT('h4)
	) name1662 (
		_w2192_,
		_w2193_,
		_w2194_
	);
	LUT2 #(
		.INIT('h1)
	) name1663 (
		_w2182_,
		_w2188_,
		_w2195_
	);
	LUT2 #(
		.INIT('h4)
	) name1664 (
		_w2194_,
		_w2195_,
		_w2196_
	);
	LUT2 #(
		.INIT('h4)
	) name1665 (
		_w2178_,
		_w2196_,
		_w2197_
	);
	LUT2 #(
		.INIT('h4)
	) name1666 (
		_w2108_,
		_w2197_,
		_w2198_
	);
	LUT2 #(
		.INIT('h4)
	) name1667 (
		_w2140_,
		_w2198_,
		_w2199_
	);
	LUT2 #(
		.INIT('h8)
	) name1668 (
		_w1368_,
		_w1376_,
		_w2200_
	);
	LUT2 #(
		.INIT('h1)
	) name1669 (
		_w1561_,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('h2)
	) name1670 (
		_w1329_,
		_w1330_,
		_w2202_
	);
	LUT2 #(
		.INIT('h2)
	) name1671 (
		_w2201_,
		_w2202_,
		_w2203_
	);
	LUT2 #(
		.INIT('h2)
	) name1672 (
		_w1429_,
		_w2203_,
		_w2204_
	);
	LUT2 #(
		.INIT('h8)
	) name1673 (
		\sa03_reg[7]/NET0131 ,
		_w1368_,
		_w2205_
	);
	LUT2 #(
		.INIT('h8)
	) name1674 (
		\sa03_reg[4]/P0001 ,
		_w1404_,
		_w2206_
	);
	LUT2 #(
		.INIT('h1)
	) name1675 (
		_w1416_,
		_w2205_,
		_w2207_
	);
	LUT2 #(
		.INIT('h4)
	) name1676 (
		_w2206_,
		_w2207_,
		_w2208_
	);
	LUT2 #(
		.INIT('h1)
	) name1677 (
		\sa03_reg[3]/P0001 ,
		_w2208_,
		_w2209_
	);
	LUT2 #(
		.INIT('h1)
	) name1678 (
		_w1369_,
		_w1446_,
		_w2210_
	);
	LUT2 #(
		.INIT('h4)
	) name1679 (
		_w2209_,
		_w2210_,
		_w2211_
	);
	LUT2 #(
		.INIT('h2)
	) name1680 (
		\sa03_reg[2]/P0001 ,
		_w2211_,
		_w2212_
	);
	LUT2 #(
		.INIT('h1)
	) name1681 (
		_w2204_,
		_w2212_,
		_w2213_
	);
	LUT2 #(
		.INIT('h2)
	) name1682 (
		\sa03_reg[1]/P0001 ,
		_w2213_,
		_w2214_
	);
	LUT2 #(
		.INIT('h1)
	) name1683 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w2215_
	);
	LUT2 #(
		.INIT('h8)
	) name1684 (
		_w1326_,
		_w1334_,
		_w2216_
	);
	LUT2 #(
		.INIT('h4)
	) name1685 (
		_w2215_,
		_w2216_,
		_w2217_
	);
	LUT2 #(
		.INIT('h4)
	) name1686 (
		\sa03_reg[6]/NET0131 ,
		_w1316_,
		_w2218_
	);
	LUT2 #(
		.INIT('h8)
	) name1687 (
		_w1376_,
		_w1398_,
		_w2219_
	);
	LUT2 #(
		.INIT('h1)
	) name1688 (
		_w2218_,
		_w2219_,
		_w2220_
	);
	LUT2 #(
		.INIT('h1)
	) name1689 (
		\sa03_reg[2]/P0001 ,
		_w2220_,
		_w2221_
	);
	LUT2 #(
		.INIT('h1)
	) name1690 (
		_w1565_,
		_w2217_,
		_w2222_
	);
	LUT2 #(
		.INIT('h4)
	) name1691 (
		_w2221_,
		_w2222_,
		_w2223_
	);
	LUT2 #(
		.INIT('h2)
	) name1692 (
		\sa03_reg[1]/P0001 ,
		_w2223_,
		_w2224_
	);
	LUT2 #(
		.INIT('h1)
	) name1693 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w2225_
	);
	LUT2 #(
		.INIT('h2)
	) name1694 (
		\sa03_reg[5]/P0001 ,
		_w1332_,
		_w2226_
	);
	LUT2 #(
		.INIT('h4)
	) name1695 (
		_w1341_,
		_w2225_,
		_w2227_
	);
	LUT2 #(
		.INIT('h8)
	) name1696 (
		_w2226_,
		_w2227_,
		_w2228_
	);
	LUT2 #(
		.INIT('h8)
	) name1697 (
		_w1316_,
		_w1367_,
		_w2229_
	);
	LUT2 #(
		.INIT('h1)
	) name1698 (
		_w1460_,
		_w2229_,
		_w2230_
	);
	LUT2 #(
		.INIT('h2)
	) name1699 (
		_w1494_,
		_w2230_,
		_w2231_
	);
	LUT2 #(
		.INIT('h1)
	) name1700 (
		_w1454_,
		_w1515_,
		_w2232_
	);
	LUT2 #(
		.INIT('h4)
	) name1701 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w2233_
	);
	LUT2 #(
		.INIT('h4)
	) name1702 (
		_w2232_,
		_w2233_,
		_w2234_
	);
	LUT2 #(
		.INIT('h8)
	) name1703 (
		\sa03_reg[2]/P0001 ,
		_w1425_,
		_w2235_
	);
	LUT2 #(
		.INIT('h8)
	) name1704 (
		\sa03_reg[4]/P0001 ,
		_w1353_,
		_w2236_
	);
	LUT2 #(
		.INIT('h1)
	) name1705 (
		_w1414_,
		_w2236_,
		_w2237_
	);
	LUT2 #(
		.INIT('h2)
	) name1706 (
		_w1374_,
		_w2237_,
		_w2238_
	);
	LUT2 #(
		.INIT('h1)
	) name1707 (
		_w1400_,
		_w1547_,
		_w2239_
	);
	LUT2 #(
		.INIT('h1)
	) name1708 (
		\sa03_reg[2]/P0001 ,
		_w2239_,
		_w2240_
	);
	LUT2 #(
		.INIT('h1)
	) name1709 (
		\sa03_reg[0]/P0001 ,
		_w2228_,
		_w2241_
	);
	LUT2 #(
		.INIT('h4)
	) name1710 (
		_w2231_,
		_w2241_,
		_w2242_
	);
	LUT2 #(
		.INIT('h1)
	) name1711 (
		_w2234_,
		_w2235_,
		_w2243_
	);
	LUT2 #(
		.INIT('h8)
	) name1712 (
		_w2242_,
		_w2243_,
		_w2244_
	);
	LUT2 #(
		.INIT('h1)
	) name1713 (
		_w2238_,
		_w2240_,
		_w2245_
	);
	LUT2 #(
		.INIT('h8)
	) name1714 (
		_w2244_,
		_w2245_,
		_w2246_
	);
	LUT2 #(
		.INIT('h4)
	) name1715 (
		_w2224_,
		_w2246_,
		_w2247_
	);
	LUT2 #(
		.INIT('h8)
	) name1716 (
		_w1316_,
		_w1326_,
		_w2248_
	);
	LUT2 #(
		.INIT('h8)
	) name1717 (
		\sa03_reg[7]/NET0131 ,
		_w2248_,
		_w2249_
	);
	LUT2 #(
		.INIT('h8)
	) name1718 (
		_w1367_,
		_w2225_,
		_w2250_
	);
	LUT2 #(
		.INIT('h4)
	) name1719 (
		\sa03_reg[6]/NET0131 ,
		_w2250_,
		_w2251_
	);
	LUT2 #(
		.INIT('h1)
	) name1720 (
		_w1398_,
		_w1408_,
		_w2252_
	);
	LUT2 #(
		.INIT('h1)
	) name1721 (
		\sa03_reg[7]/NET0131 ,
		_w2252_,
		_w2253_
	);
	LUT2 #(
		.INIT('h1)
	) name1722 (
		_w1368_,
		_w1533_,
		_w2254_
	);
	LUT2 #(
		.INIT('h4)
	) name1723 (
		_w2253_,
		_w2254_,
		_w2255_
	);
	LUT2 #(
		.INIT('h2)
	) name1724 (
		\sa03_reg[2]/P0001 ,
		_w2255_,
		_w2256_
	);
	LUT2 #(
		.INIT('h1)
	) name1725 (
		_w2249_,
		_w2251_,
		_w2257_
	);
	LUT2 #(
		.INIT('h4)
	) name1726 (
		_w2256_,
		_w2257_,
		_w2258_
	);
	LUT2 #(
		.INIT('h2)
	) name1727 (
		\sa03_reg[1]/P0001 ,
		_w2258_,
		_w2259_
	);
	LUT2 #(
		.INIT('h8)
	) name1728 (
		\sa03_reg[4]/P0001 ,
		_w1342_,
		_w2260_
	);
	LUT2 #(
		.INIT('h1)
	) name1729 (
		_w1482_,
		_w1533_,
		_w2261_
	);
	LUT2 #(
		.INIT('h4)
	) name1730 (
		_w2260_,
		_w2261_,
		_w2262_
	);
	LUT2 #(
		.INIT('h1)
	) name1731 (
		\sa03_reg[2]/P0001 ,
		_w2262_,
		_w2263_
	);
	LUT2 #(
		.INIT('h4)
	) name1732 (
		\sa03_reg[4]/P0001 ,
		_w1367_,
		_w2264_
	);
	LUT2 #(
		.INIT('h8)
	) name1733 (
		_w1436_,
		_w2264_,
		_w2265_
	);
	LUT2 #(
		.INIT('h8)
	) name1734 (
		_w1329_,
		_w1423_,
		_w2266_
	);
	LUT2 #(
		.INIT('h2)
	) name1735 (
		\sa03_reg[2]/P0001 ,
		_w1334_,
		_w2267_
	);
	LUT2 #(
		.INIT('h2)
	) name1736 (
		_w1318_,
		_w1324_,
		_w2268_
	);
	LUT2 #(
		.INIT('h4)
	) name1737 (
		_w2267_,
		_w2268_,
		_w2269_
	);
	LUT2 #(
		.INIT('h1)
	) name1738 (
		_w2265_,
		_w2266_,
		_w2270_
	);
	LUT2 #(
		.INIT('h4)
	) name1739 (
		_w2269_,
		_w2270_,
		_w2271_
	);
	LUT2 #(
		.INIT('h4)
	) name1740 (
		_w2263_,
		_w2271_,
		_w2272_
	);
	LUT2 #(
		.INIT('h1)
	) name1741 (
		\sa03_reg[1]/P0001 ,
		_w2272_,
		_w2273_
	);
	LUT2 #(
		.INIT('h1)
	) name1742 (
		_w1364_,
		_w2205_,
		_w2274_
	);
	LUT2 #(
		.INIT('h1)
	) name1743 (
		\sa03_reg[3]/P0001 ,
		_w2274_,
		_w2275_
	);
	LUT2 #(
		.INIT('h1)
	) name1744 (
		_w1343_,
		_w2275_,
		_w2276_
	);
	LUT2 #(
		.INIT('h2)
	) name1745 (
		\sa03_reg[2]/P0001 ,
		_w2276_,
		_w2277_
	);
	LUT2 #(
		.INIT('h8)
	) name1746 (
		_w1374_,
		_w1431_,
		_w2278_
	);
	LUT2 #(
		.INIT('h8)
	) name1747 (
		_w1334_,
		_w1449_,
		_w2279_
	);
	LUT2 #(
		.INIT('h8)
	) name1748 (
		_w1482_,
		_w2225_,
		_w2280_
	);
	LUT2 #(
		.INIT('h2)
	) name1749 (
		\sa03_reg[0]/P0001 ,
		_w2279_,
		_w2281_
	);
	LUT2 #(
		.INIT('h4)
	) name1750 (
		_w2278_,
		_w2281_,
		_w2282_
	);
	LUT2 #(
		.INIT('h4)
	) name1751 (
		_w2280_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('h4)
	) name1752 (
		_w2277_,
		_w2283_,
		_w2284_
	);
	LUT2 #(
		.INIT('h4)
	) name1753 (
		_w2259_,
		_w2284_,
		_w2285_
	);
	LUT2 #(
		.INIT('h4)
	) name1754 (
		_w2273_,
		_w2285_,
		_w2286_
	);
	LUT2 #(
		.INIT('h1)
	) name1755 (
		_w2247_,
		_w2286_,
		_w2287_
	);
	LUT2 #(
		.INIT('h8)
	) name1756 (
		_w1376_,
		_w2218_,
		_w2288_
	);
	LUT2 #(
		.INIT('h4)
	) name1757 (
		\sa03_reg[3]/P0001 ,
		_w1435_,
		_w2289_
	);
	LUT2 #(
		.INIT('h4)
	) name1758 (
		\sa03_reg[4]/P0001 ,
		_w2289_,
		_w2290_
	);
	LUT2 #(
		.INIT('h1)
	) name1759 (
		_w2288_,
		_w2290_,
		_w2291_
	);
	LUT2 #(
		.INIT('h1)
	) name1760 (
		\sa03_reg[2]/P0001 ,
		_w2291_,
		_w2292_
	);
	LUT2 #(
		.INIT('h8)
	) name1761 (
		_w1334_,
		_w1339_,
		_w2293_
	);
	LUT2 #(
		.INIT('h1)
	) name1762 (
		_w1325_,
		_w1420_,
		_w2294_
	);
	LUT2 #(
		.INIT('h4)
	) name1763 (
		_w2249_,
		_w2294_,
		_w2295_
	);
	LUT2 #(
		.INIT('h2)
	) name1764 (
		\sa03_reg[2]/P0001 ,
		_w2295_,
		_w2296_
	);
	LUT2 #(
		.INIT('h8)
	) name1765 (
		_w1429_,
		_w2264_,
		_w2297_
	);
	LUT2 #(
		.INIT('h1)
	) name1766 (
		_w2228_,
		_w2293_,
		_w2298_
	);
	LUT2 #(
		.INIT('h4)
	) name1767 (
		_w2297_,
		_w2298_,
		_w2299_
	);
	LUT2 #(
		.INIT('h4)
	) name1768 (
		_w2296_,
		_w2299_,
		_w2300_
	);
	LUT2 #(
		.INIT('h1)
	) name1769 (
		\sa03_reg[1]/P0001 ,
		_w2300_,
		_w2301_
	);
	LUT2 #(
		.INIT('h1)
	) name1770 (
		_w2292_,
		_w2301_,
		_w2302_
	);
	LUT2 #(
		.INIT('h4)
	) name1771 (
		_w2214_,
		_w2302_,
		_w2303_
	);
	LUT2 #(
		.INIT('h4)
	) name1772 (
		_w2287_,
		_w2303_,
		_w2304_
	);
	LUT2 #(
		.INIT('h2)
	) name1773 (
		_w2199_,
		_w2304_,
		_w2305_
	);
	LUT2 #(
		.INIT('h4)
	) name1774 (
		_w2199_,
		_w2304_,
		_w2306_
	);
	LUT2 #(
		.INIT('h1)
	) name1775 (
		_w2305_,
		_w2306_,
		_w2307_
	);
	LUT2 #(
		.INIT('h1)
	) name1776 (
		_w1581_,
		_w2307_,
		_w2308_
	);
	LUT2 #(
		.INIT('h8)
	) name1777 (
		_w1581_,
		_w2307_,
		_w2309_
	);
	LUT2 #(
		.INIT('h1)
	) name1778 (
		_w2308_,
		_w2309_,
		_w2310_
	);
	LUT2 #(
		.INIT('h8)
	) name1779 (
		_w1920_,
		_w1951_,
		_w2311_
	);
	LUT2 #(
		.INIT('h1)
	) name1780 (
		_w1936_,
		_w2311_,
		_w2312_
	);
	LUT2 #(
		.INIT('h1)
	) name1781 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		_w2313_
	);
	LUT2 #(
		.INIT('h8)
	) name1782 (
		_w1955_,
		_w2313_,
		_w2314_
	);
	LUT2 #(
		.INIT('h8)
	) name1783 (
		\sa32_reg[4]/P0001 ,
		_w1981_,
		_w2315_
	);
	LUT2 #(
		.INIT('h8)
	) name1784 (
		_w1915_,
		_w1995_,
		_w2316_
	);
	LUT2 #(
		.INIT('h8)
	) name1785 (
		\sa32_reg[7]/P0001 ,
		_w2316_,
		_w2317_
	);
	LUT2 #(
		.INIT('h1)
	) name1786 (
		_w1994_,
		_w2315_,
		_w2318_
	);
	LUT2 #(
		.INIT('h4)
	) name1787 (
		_w2317_,
		_w2318_,
		_w2319_
	);
	LUT2 #(
		.INIT('h2)
	) name1788 (
		\sa32_reg[2]/P0001 ,
		_w2319_,
		_w2320_
	);
	LUT2 #(
		.INIT('h2)
	) name1789 (
		_w2312_,
		_w2314_,
		_w2321_
	);
	LUT2 #(
		.INIT('h4)
	) name1790 (
		_w2320_,
		_w2321_,
		_w2322_
	);
	LUT2 #(
		.INIT('h2)
	) name1791 (
		\sa32_reg[1]/P0001 ,
		_w2322_,
		_w2323_
	);
	LUT2 #(
		.INIT('h8)
	) name1792 (
		_w1970_,
		_w1981_,
		_w2324_
	);
	LUT2 #(
		.INIT('h1)
	) name1793 (
		_w1940_,
		_w2324_,
		_w2325_
	);
	LUT2 #(
		.INIT('h1)
	) name1794 (
		\sa32_reg[2]/P0001 ,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h8)
	) name1795 (
		\sa32_reg[4]/P0001 ,
		_w1969_,
		_w2327_
	);
	LUT2 #(
		.INIT('h1)
	) name1796 (
		_w1922_,
		_w2327_,
		_w2328_
	);
	LUT2 #(
		.INIT('h1)
	) name1797 (
		_w1925_,
		_w2033_,
		_w2329_
	);
	LUT2 #(
		.INIT('h8)
	) name1798 (
		_w2328_,
		_w2329_,
		_w2330_
	);
	LUT2 #(
		.INIT('h2)
	) name1799 (
		\sa32_reg[2]/P0001 ,
		_w2330_,
		_w2331_
	);
	LUT2 #(
		.INIT('h4)
	) name1800 (
		\sa32_reg[3]/P0001 ,
		_w2060_,
		_w2332_
	);
	LUT2 #(
		.INIT('h1)
	) name1801 (
		\sa32_reg[2]/P0001 ,
		_w2332_,
		_w2333_
	);
	LUT2 #(
		.INIT('h8)
	) name1802 (
		\sa32_reg[7]/P0001 ,
		_w1912_,
		_w2334_
	);
	LUT2 #(
		.INIT('h2)
	) name1803 (
		\sa32_reg[2]/P0001 ,
		_w2019_,
		_w2335_
	);
	LUT2 #(
		.INIT('h4)
	) name1804 (
		_w2334_,
		_w2335_,
		_w2336_
	);
	LUT2 #(
		.INIT('h1)
	) name1805 (
		_w2333_,
		_w2336_,
		_w2337_
	);
	LUT2 #(
		.INIT('h4)
	) name1806 (
		_w2024_,
		_w2032_,
		_w2338_
	);
	LUT2 #(
		.INIT('h4)
	) name1807 (
		_w2337_,
		_w2338_,
		_w2339_
	);
	LUT2 #(
		.INIT('h1)
	) name1808 (
		\sa32_reg[1]/P0001 ,
		_w2339_,
		_w2340_
	);
	LUT2 #(
		.INIT('h1)
	) name1809 (
		_w2326_,
		_w2331_,
		_w2341_
	);
	LUT2 #(
		.INIT('h4)
	) name1810 (
		_w2323_,
		_w2341_,
		_w2342_
	);
	LUT2 #(
		.INIT('h4)
	) name1811 (
		_w2340_,
		_w2342_,
		_w2343_
	);
	LUT2 #(
		.INIT('h2)
	) name1812 (
		\sa32_reg[0]/P0002 ,
		_w2343_,
		_w2344_
	);
	LUT2 #(
		.INIT('h8)
	) name1813 (
		_w1909_,
		_w1995_,
		_w2345_
	);
	LUT2 #(
		.INIT('h8)
	) name1814 (
		_w1970_,
		_w1987_,
		_w2346_
	);
	LUT2 #(
		.INIT('h8)
	) name1815 (
		\sa32_reg[2]/P0001 ,
		_w2346_,
		_w2347_
	);
	LUT2 #(
		.INIT('h2)
	) name1816 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w2348_
	);
	LUT2 #(
		.INIT('h8)
	) name1817 (
		_w1913_,
		_w2348_,
		_w2349_
	);
	LUT2 #(
		.INIT('h8)
	) name1818 (
		\sa32_reg[3]/P0001 ,
		_w2349_,
		_w2350_
	);
	LUT2 #(
		.INIT('h4)
	) name1819 (
		\sa32_reg[5]/P0001 ,
		_w2315_,
		_w2351_
	);
	LUT2 #(
		.INIT('h8)
	) name1820 (
		\sa32_reg[5]/P0001 ,
		_w1932_,
		_w2352_
	);
	LUT2 #(
		.INIT('h1)
	) name1821 (
		_w2024_,
		_w2351_,
		_w2353_
	);
	LUT2 #(
		.INIT('h4)
	) name1822 (
		_w2352_,
		_w2353_,
		_w2354_
	);
	LUT2 #(
		.INIT('h1)
	) name1823 (
		\sa32_reg[2]/P0001 ,
		_w2354_,
		_w2355_
	);
	LUT2 #(
		.INIT('h8)
	) name1824 (
		_w1912_,
		_w1923_,
		_w2356_
	);
	LUT2 #(
		.INIT('h1)
	) name1825 (
		_w2345_,
		_w2356_,
		_w2357_
	);
	LUT2 #(
		.INIT('h4)
	) name1826 (
		_w2347_,
		_w2357_,
		_w2358_
	);
	LUT2 #(
		.INIT('h4)
	) name1827 (
		_w2350_,
		_w2358_,
		_w2359_
	);
	LUT2 #(
		.INIT('h4)
	) name1828 (
		_w2355_,
		_w2359_,
		_w2360_
	);
	LUT2 #(
		.INIT('h1)
	) name1829 (
		\sa32_reg[1]/P0001 ,
		_w2360_,
		_w2361_
	);
	LUT2 #(
		.INIT('h4)
	) name1830 (
		\sa32_reg[7]/P0001 ,
		_w1995_,
		_w2362_
	);
	LUT2 #(
		.INIT('h8)
	) name1831 (
		_w1990_,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('h4)
	) name1832 (
		\sa32_reg[2]/P0001 ,
		_w2334_,
		_w2364_
	);
	LUT2 #(
		.INIT('h8)
	) name1833 (
		_w1939_,
		_w2364_,
		_w2365_
	);
	LUT2 #(
		.INIT('h8)
	) name1834 (
		_w1924_,
		_w1981_,
		_w2366_
	);
	LUT2 #(
		.INIT('h8)
	) name1835 (
		_w2046_,
		_w2366_,
		_w2367_
	);
	LUT2 #(
		.INIT('h4)
	) name1836 (
		\sa32_reg[2]/P0001 ,
		_w2063_,
		_w2368_
	);
	LUT2 #(
		.INIT('h8)
	) name1837 (
		\sa32_reg[1]/P0001 ,
		_w2368_,
		_w2369_
	);
	LUT2 #(
		.INIT('h8)
	) name1838 (
		\sa32_reg[1]/P0001 ,
		\sa32_reg[2]/P0001 ,
		_w2370_
	);
	LUT2 #(
		.INIT('h1)
	) name1839 (
		_w2028_,
		_w2311_,
		_w2371_
	);
	LUT2 #(
		.INIT('h4)
	) name1840 (
		_w2362_,
		_w2371_,
		_w2372_
	);
	LUT2 #(
		.INIT('h4)
	) name1841 (
		\sa32_reg[6]/NET0131 ,
		_w2370_,
		_w2373_
	);
	LUT2 #(
		.INIT('h4)
	) name1842 (
		_w2372_,
		_w2373_,
		_w2374_
	);
	LUT2 #(
		.INIT('h4)
	) name1843 (
		_w1913_,
		_w1924_,
		_w2375_
	);
	LUT2 #(
		.INIT('h2)
	) name1844 (
		\sa32_reg[4]/P0001 ,
		_w1987_,
		_w2376_
	);
	LUT2 #(
		.INIT('h2)
	) name1845 (
		_w2375_,
		_w2376_,
		_w2377_
	);
	LUT2 #(
		.INIT('h1)
	) name1846 (
		_w1910_,
		_w1990_,
		_w2378_
	);
	LUT2 #(
		.INIT('h2)
	) name1847 (
		_w1919_,
		_w2378_,
		_w2379_
	);
	LUT2 #(
		.INIT('h1)
	) name1848 (
		\sa32_reg[2]/P0001 ,
		_w2377_,
		_w2380_
	);
	LUT2 #(
		.INIT('h4)
	) name1849 (
		_w2379_,
		_w2380_,
		_w2381_
	);
	LUT2 #(
		.INIT('h8)
	) name1850 (
		_w1990_,
		_w1995_,
		_w2382_
	);
	LUT2 #(
		.INIT('h8)
	) name1851 (
		_w1953_,
		_w1965_,
		_w2383_
	);
	LUT2 #(
		.INIT('h2)
	) name1852 (
		\sa32_reg[2]/P0001 ,
		_w2382_,
		_w2384_
	);
	LUT2 #(
		.INIT('h4)
	) name1853 (
		_w2383_,
		_w2384_,
		_w2385_
	);
	LUT2 #(
		.INIT('h1)
	) name1854 (
		_w2381_,
		_w2385_,
		_w2386_
	);
	LUT2 #(
		.INIT('h4)
	) name1855 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w2387_
	);
	LUT2 #(
		.INIT('h8)
	) name1856 (
		_w1951_,
		_w2387_,
		_w2388_
	);
	LUT2 #(
		.INIT('h4)
	) name1857 (
		\sa32_reg[3]/P0001 ,
		_w1923_,
		_w2389_
	);
	LUT2 #(
		.INIT('h4)
	) name1858 (
		\sa32_reg[4]/P0001 ,
		_w2389_,
		_w2390_
	);
	LUT2 #(
		.INIT('h1)
	) name1859 (
		\sa32_reg[1]/P0001 ,
		_w2324_,
		_w2391_
	);
	LUT2 #(
		.INIT('h4)
	) name1860 (
		_w2388_,
		_w2391_,
		_w2392_
	);
	LUT2 #(
		.INIT('h1)
	) name1861 (
		_w2061_,
		_w2364_,
		_w2393_
	);
	LUT2 #(
		.INIT('h1)
	) name1862 (
		_w2383_,
		_w2390_,
		_w2394_
	);
	LUT2 #(
		.INIT('h8)
	) name1863 (
		_w2393_,
		_w2394_,
		_w2395_
	);
	LUT2 #(
		.INIT('h8)
	) name1864 (
		_w2392_,
		_w2395_,
		_w2396_
	);
	LUT2 #(
		.INIT('h2)
	) name1865 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		_w2397_
	);
	LUT2 #(
		.INIT('h8)
	) name1866 (
		\sa32_reg[4]/P0001 ,
		_w1920_,
		_w2398_
	);
	LUT2 #(
		.INIT('h4)
	) name1867 (
		\sa32_reg[4]/P0001 ,
		_w2027_,
		_w2399_
	);
	LUT2 #(
		.INIT('h1)
	) name1868 (
		_w2398_,
		_w2399_,
		_w2400_
	);
	LUT2 #(
		.INIT('h2)
	) name1869 (
		_w2397_,
		_w2400_,
		_w2401_
	);
	LUT2 #(
		.INIT('h4)
	) name1870 (
		\sa32_reg[2]/P0001 ,
		_w2033_,
		_w2402_
	);
	LUT2 #(
		.INIT('h2)
	) name1871 (
		\sa32_reg[1]/P0001 ,
		_w2052_,
		_w2403_
	);
	LUT2 #(
		.INIT('h4)
	) name1872 (
		_w2402_,
		_w2403_,
		_w2404_
	);
	LUT2 #(
		.INIT('h4)
	) name1873 (
		_w2401_,
		_w2404_,
		_w2405_
	);
	LUT2 #(
		.INIT('h1)
	) name1874 (
		_w2396_,
		_w2405_,
		_w2406_
	);
	LUT2 #(
		.INIT('h1)
	) name1875 (
		_w2386_,
		_w2406_,
		_w2407_
	);
	LUT2 #(
		.INIT('h1)
	) name1876 (
		\sa32_reg[0]/P0002 ,
		_w2407_,
		_w2408_
	);
	LUT2 #(
		.INIT('h1)
	) name1877 (
		_w2363_,
		_w2367_,
		_w2409_
	);
	LUT2 #(
		.INIT('h4)
	) name1878 (
		_w2010_,
		_w2409_,
		_w2410_
	);
	LUT2 #(
		.INIT('h4)
	) name1879 (
		_w2365_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('h1)
	) name1880 (
		_w2369_,
		_w2374_,
		_w2412_
	);
	LUT2 #(
		.INIT('h8)
	) name1881 (
		_w2411_,
		_w2412_,
		_w2413_
	);
	LUT2 #(
		.INIT('h4)
	) name1882 (
		_w2361_,
		_w2413_,
		_w2414_
	);
	LUT2 #(
		.INIT('h4)
	) name1883 (
		_w2408_,
		_w2414_,
		_w2415_
	);
	LUT2 #(
		.INIT('h4)
	) name1884 (
		_w2344_,
		_w2415_,
		_w2416_
	);
	LUT2 #(
		.INIT('h8)
	) name1885 (
		_w1753_,
		_w1784_,
		_w2417_
	);
	LUT2 #(
		.INIT('h1)
	) name1886 (
		_w1892_,
		_w2417_,
		_w2418_
	);
	LUT2 #(
		.INIT('h2)
	) name1887 (
		_w1772_,
		_w1793_,
		_w2419_
	);
	LUT2 #(
		.INIT('h2)
	) name1888 (
		_w2418_,
		_w2419_,
		_w2420_
	);
	LUT2 #(
		.INIT('h2)
	) name1889 (
		_w1877_,
		_w2420_,
		_w2421_
	);
	LUT2 #(
		.INIT('h8)
	) name1890 (
		\sa21_reg[5]/P0001 ,
		_w1841_,
		_w2422_
	);
	LUT2 #(
		.INIT('h1)
	) name1891 (
		_w1822_,
		_w2422_,
		_w2423_
	);
	LUT2 #(
		.INIT('h1)
	) name1892 (
		\sa21_reg[4]/P0001 ,
		_w2423_,
		_w2424_
	);
	LUT2 #(
		.INIT('h4)
	) name1893 (
		\sa21_reg[5]/P0001 ,
		_w1763_,
		_w2425_
	);
	LUT2 #(
		.INIT('h8)
	) name1894 (
		\sa21_reg[4]/P0001 ,
		_w2425_,
		_w2426_
	);
	LUT2 #(
		.INIT('h1)
	) name1895 (
		_w2424_,
		_w2426_,
		_w2427_
	);
	LUT2 #(
		.INIT('h1)
	) name1896 (
		\sa21_reg[3]/P0001 ,
		_w2427_,
		_w2428_
	);
	LUT2 #(
		.INIT('h8)
	) name1897 (
		_w1837_,
		_w1854_,
		_w2429_
	);
	LUT2 #(
		.INIT('h1)
	) name1898 (
		_w1794_,
		_w2429_,
		_w2430_
	);
	LUT2 #(
		.INIT('h4)
	) name1899 (
		_w2428_,
		_w2430_,
		_w2431_
	);
	LUT2 #(
		.INIT('h2)
	) name1900 (
		\sa21_reg[2]/P0001 ,
		_w2431_,
		_w2432_
	);
	LUT2 #(
		.INIT('h1)
	) name1901 (
		_w2421_,
		_w2432_,
		_w2433_
	);
	LUT2 #(
		.INIT('h2)
	) name1902 (
		\sa21_reg[1]/P0001 ,
		_w2433_,
		_w2434_
	);
	LUT2 #(
		.INIT('h8)
	) name1903 (
		\sa21_reg[7]/P0001 ,
		_w1890_,
		_w2435_
	);
	LUT2 #(
		.INIT('h8)
	) name1904 (
		\sa21_reg[5]/P0001 ,
		_w1762_,
		_w2436_
	);
	LUT2 #(
		.INIT('h4)
	) name1905 (
		\sa21_reg[3]/P0001 ,
		_w1841_,
		_w2437_
	);
	LUT2 #(
		.INIT('h1)
	) name1906 (
		_w1779_,
		_w2437_,
		_w2438_
	);
	LUT2 #(
		.INIT('h1)
	) name1907 (
		_w1753_,
		_w1844_,
		_w2439_
	);
	LUT2 #(
		.INIT('h8)
	) name1908 (
		_w2438_,
		_w2439_,
		_w2440_
	);
	LUT2 #(
		.INIT('h2)
	) name1909 (
		\sa21_reg[1]/P0001 ,
		_w2440_,
		_w2441_
	);
	LUT2 #(
		.INIT('h1)
	) name1910 (
		_w1774_,
		_w2435_,
		_w2442_
	);
	LUT2 #(
		.INIT('h4)
	) name1911 (
		_w2436_,
		_w2442_,
		_w2443_
	);
	LUT2 #(
		.INIT('h4)
	) name1912 (
		_w2441_,
		_w2443_,
		_w2444_
	);
	LUT2 #(
		.INIT('h2)
	) name1913 (
		\sa21_reg[2]/P0001 ,
		_w2444_,
		_w2445_
	);
	LUT2 #(
		.INIT('h8)
	) name1914 (
		_w1754_,
		_w1761_,
		_w2446_
	);
	LUT2 #(
		.INIT('h4)
	) name1915 (
		\sa21_reg[6]/NET0131 ,
		_w1867_,
		_w2447_
	);
	LUT2 #(
		.INIT('h1)
	) name1916 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w2448_
	);
	LUT2 #(
		.INIT('h8)
	) name1917 (
		_w1837_,
		_w2448_,
		_w2449_
	);
	LUT2 #(
		.INIT('h8)
	) name1918 (
		\sa21_reg[6]/NET0131 ,
		_w1773_,
		_w2450_
	);
	LUT2 #(
		.INIT('h4)
	) name1919 (
		\sa21_reg[7]/P0001 ,
		_w2450_,
		_w2451_
	);
	LUT2 #(
		.INIT('h4)
	) name1920 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w2452_
	);
	LUT2 #(
		.INIT('h8)
	) name1921 (
		\sa21_reg[2]/P0001 ,
		_w1815_,
		_w2453_
	);
	LUT2 #(
		.INIT('h8)
	) name1922 (
		_w2452_,
		_w2453_,
		_w2454_
	);
	LUT2 #(
		.INIT('h4)
	) name1923 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w2455_
	);
	LUT2 #(
		.INIT('h4)
	) name1924 (
		_w1772_,
		_w2455_,
		_w2456_
	);
	LUT2 #(
		.INIT('h4)
	) name1925 (
		_w1823_,
		_w2456_,
		_w2457_
	);
	LUT2 #(
		.INIT('h1)
	) name1926 (
		_w2446_,
		_w2449_,
		_w2458_
	);
	LUT2 #(
		.INIT('h4)
	) name1927 (
		_w2447_,
		_w2458_,
		_w2459_
	);
	LUT2 #(
		.INIT('h1)
	) name1928 (
		_w2451_,
		_w2454_,
		_w2460_
	);
	LUT2 #(
		.INIT('h4)
	) name1929 (
		_w2457_,
		_w2460_,
		_w2461_
	);
	LUT2 #(
		.INIT('h8)
	) name1930 (
		_w2459_,
		_w2461_,
		_w2462_
	);
	LUT2 #(
		.INIT('h1)
	) name1931 (
		\sa21_reg[1]/P0001 ,
		_w2462_,
		_w2463_
	);
	LUT2 #(
		.INIT('h8)
	) name1932 (
		_w1759_,
		_w1894_,
		_w2464_
	);
	LUT2 #(
		.INIT('h8)
	) name1933 (
		_w1802_,
		_w1823_,
		_w2465_
	);
	LUT2 #(
		.INIT('h8)
	) name1934 (
		_w1754_,
		_w2425_,
		_w2466_
	);
	LUT2 #(
		.INIT('h1)
	) name1935 (
		_w2465_,
		_w2466_,
		_w2467_
	);
	LUT2 #(
		.INIT('h2)
	) name1936 (
		\sa21_reg[1]/P0001 ,
		_w2467_,
		_w2468_
	);
	LUT2 #(
		.INIT('h8)
	) name1937 (
		_w1745_,
		_w1773_,
		_w2469_
	);
	LUT2 #(
		.INIT('h8)
	) name1938 (
		_w1754_,
		_w1762_,
		_w2470_
	);
	LUT2 #(
		.INIT('h1)
	) name1939 (
		_w2464_,
		_w2469_,
		_w2471_
	);
	LUT2 #(
		.INIT('h4)
	) name1940 (
		_w2470_,
		_w2471_,
		_w2472_
	);
	LUT2 #(
		.INIT('h4)
	) name1941 (
		_w2468_,
		_w2472_,
		_w2473_
	);
	LUT2 #(
		.INIT('h4)
	) name1942 (
		_w2445_,
		_w2473_,
		_w2474_
	);
	LUT2 #(
		.INIT('h4)
	) name1943 (
		_w2463_,
		_w2474_,
		_w2475_
	);
	LUT2 #(
		.INIT('h2)
	) name1944 (
		\sa21_reg[0]/P0001 ,
		_w2475_,
		_w2476_
	);
	LUT2 #(
		.INIT('h4)
	) name1945 (
		\sa21_reg[5]/P0001 ,
		_w1841_,
		_w2477_
	);
	LUT2 #(
		.INIT('h8)
	) name1946 (
		\sa21_reg[2]/P0001 ,
		_w2477_,
		_w2478_
	);
	LUT2 #(
		.INIT('h1)
	) name1947 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w2479_
	);
	LUT2 #(
		.INIT('h1)
	) name1948 (
		_w1867_,
		_w2479_,
		_w2480_
	);
	LUT2 #(
		.INIT('h2)
	) name1949 (
		\sa21_reg[7]/P0001 ,
		_w2480_,
		_w2481_
	);
	LUT2 #(
		.INIT('h1)
	) name1950 (
		_w2478_,
		_w2481_,
		_w2482_
	);
	LUT2 #(
		.INIT('h1)
	) name1951 (
		\sa21_reg[1]/P0001 ,
		_w2482_,
		_w2483_
	);
	LUT2 #(
		.INIT('h1)
	) name1952 (
		_w1781_,
		_w1879_,
		_w2484_
	);
	LUT2 #(
		.INIT('h2)
	) name1953 (
		_w1754_,
		_w2484_,
		_w2485_
	);
	LUT2 #(
		.INIT('h8)
	) name1954 (
		_w1786_,
		_w1894_,
		_w2486_
	);
	LUT2 #(
		.INIT('h1)
	) name1955 (
		_w1855_,
		_w1864_,
		_w2487_
	);
	LUT2 #(
		.INIT('h1)
	) name1956 (
		\sa21_reg[2]/P0001 ,
		_w2487_,
		_w2488_
	);
	LUT2 #(
		.INIT('h8)
	) name1957 (
		\sa21_reg[6]/NET0131 ,
		_w1849_,
		_w2489_
	);
	LUT2 #(
		.INIT('h8)
	) name1958 (
		\sa21_reg[4]/P0001 ,
		_w2452_,
		_w2490_
	);
	LUT2 #(
		.INIT('h4)
	) name1959 (
		\sa21_reg[1]/P0001 ,
		_w2490_,
		_w2491_
	);
	LUT2 #(
		.INIT('h8)
	) name1960 (
		\sa21_reg[4]/P0001 ,
		_w1841_,
		_w2492_
	);
	LUT2 #(
		.INIT('h8)
	) name1961 (
		\sa21_reg[5]/P0001 ,
		_w2492_,
		_w2493_
	);
	LUT2 #(
		.INIT('h1)
	) name1962 (
		_w2489_,
		_w2491_,
		_w2494_
	);
	LUT2 #(
		.INIT('h4)
	) name1963 (
		_w2493_,
		_w2494_,
		_w2495_
	);
	LUT2 #(
		.INIT('h2)
	) name1964 (
		_w1894_,
		_w2495_,
		_w2496_
	);
	LUT2 #(
		.INIT('h1)
	) name1965 (
		_w2485_,
		_w2486_,
		_w2497_
	);
	LUT2 #(
		.INIT('h4)
	) name1966 (
		_w2488_,
		_w2497_,
		_w2498_
	);
	LUT2 #(
		.INIT('h4)
	) name1967 (
		_w2483_,
		_w2498_,
		_w2499_
	);
	LUT2 #(
		.INIT('h4)
	) name1968 (
		_w2496_,
		_w2499_,
		_w2500_
	);
	LUT2 #(
		.INIT('h1)
	) name1969 (
		\sa21_reg[0]/P0001 ,
		_w2500_,
		_w2501_
	);
	LUT2 #(
		.INIT('h8)
	) name1970 (
		_w1832_,
		_w1854_,
		_w2502_
	);
	LUT2 #(
		.INIT('h8)
	) name1971 (
		\sa21_reg[5]/P0001 ,
		_w2450_,
		_w2503_
	);
	LUT2 #(
		.INIT('h1)
	) name1972 (
		_w2465_,
		_w2502_,
		_w2504_
	);
	LUT2 #(
		.INIT('h4)
	) name1973 (
		_w2503_,
		_w2504_,
		_w2505_
	);
	LUT2 #(
		.INIT('h2)
	) name1974 (
		\sa21_reg[2]/P0001 ,
		_w2505_,
		_w2506_
	);
	LUT2 #(
		.INIT('h4)
	) name1975 (
		\sa21_reg[2]/P0001 ,
		_w1818_,
		_w2507_
	);
	LUT2 #(
		.INIT('h8)
	) name1976 (
		_w1749_,
		_w1773_,
		_w2508_
	);
	LUT2 #(
		.INIT('h1)
	) name1977 (
		_w2507_,
		_w2508_,
		_w2509_
	);
	LUT2 #(
		.INIT('h4)
	) name1978 (
		_w2485_,
		_w2509_,
		_w2510_
	);
	LUT2 #(
		.INIT('h4)
	) name1979 (
		_w2506_,
		_w2510_,
		_w2511_
	);
	LUT2 #(
		.INIT('h1)
	) name1980 (
		\sa21_reg[1]/P0001 ,
		_w2511_,
		_w2512_
	);
	LUT2 #(
		.INIT('h8)
	) name1981 (
		_w1761_,
		_w1787_,
		_w2513_
	);
	LUT2 #(
		.INIT('h1)
	) name1982 (
		_w1747_,
		_w2513_,
		_w2514_
	);
	LUT2 #(
		.INIT('h1)
	) name1983 (
		\sa21_reg[2]/P0001 ,
		_w2514_,
		_w2515_
	);
	LUT2 #(
		.INIT('h4)
	) name1984 (
		\sa21_reg[5]/P0001 ,
		_w2450_,
		_w2516_
	);
	LUT2 #(
		.INIT('h4)
	) name1985 (
		_w2448_,
		_w2516_,
		_w2517_
	);
	LUT2 #(
		.INIT('h1)
	) name1986 (
		_w1885_,
		_w2515_,
		_w2518_
	);
	LUT2 #(
		.INIT('h4)
	) name1987 (
		_w2517_,
		_w2518_,
		_w2519_
	);
	LUT2 #(
		.INIT('h4)
	) name1988 (
		\sa21_reg[0]/P0001 ,
		\sa21_reg[1]/P0001 ,
		_w2520_
	);
	LUT2 #(
		.INIT('h4)
	) name1989 (
		_w2519_,
		_w2520_,
		_w2521_
	);
	LUT2 #(
		.INIT('h4)
	) name1990 (
		\sa21_reg[5]/P0001 ,
		_w1747_,
		_w2522_
	);
	LUT2 #(
		.INIT('h1)
	) name1991 (
		_w1891_,
		_w2522_,
		_w2523_
	);
	LUT2 #(
		.INIT('h2)
	) name1992 (
		_w2448_,
		_w2523_,
		_w2524_
	);
	LUT2 #(
		.INIT('h1)
	) name1993 (
		_w2521_,
		_w2524_,
		_w2525_
	);
	LUT2 #(
		.INIT('h4)
	) name1994 (
		_w2512_,
		_w2525_,
		_w2526_
	);
	LUT2 #(
		.INIT('h4)
	) name1995 (
		_w2501_,
		_w2526_,
		_w2527_
	);
	LUT2 #(
		.INIT('h4)
	) name1996 (
		_w2434_,
		_w2527_,
		_w2528_
	);
	LUT2 #(
		.INIT('h4)
	) name1997 (
		_w2476_,
		_w2528_,
		_w2529_
	);
	LUT2 #(
		.INIT('h2)
	) name1998 (
		\u0_w_reg[3][7]/P0001 ,
		_w2529_,
		_w2530_
	);
	LUT2 #(
		.INIT('h4)
	) name1999 (
		\u0_w_reg[3][7]/P0001 ,
		_w2529_,
		_w2531_
	);
	LUT2 #(
		.INIT('h1)
	) name2000 (
		_w2530_,
		_w2531_,
		_w2532_
	);
	LUT2 #(
		.INIT('h8)
	) name2001 (
		_w2416_,
		_w2532_,
		_w2533_
	);
	LUT2 #(
		.INIT('h1)
	) name2002 (
		_w2416_,
		_w2532_,
		_w2534_
	);
	LUT2 #(
		.INIT('h1)
	) name2003 (
		_w2533_,
		_w2534_,
		_w2535_
	);
	LUT2 #(
		.INIT('h1)
	) name2004 (
		_w2310_,
		_w2535_,
		_w2536_
	);
	LUT2 #(
		.INIT('h8)
	) name2005 (
		_w2310_,
		_w2535_,
		_w2537_
	);
	LUT2 #(
		.INIT('h1)
	) name2006 (
		\ld_r_reg/P0001 ,
		_w2536_,
		_w2538_
	);
	LUT2 #(
		.INIT('h4)
	) name2007 (
		_w2537_,
		_w2538_,
		_w2539_
	);
	LUT2 #(
		.INIT('h2)
	) name2008 (
		\text_in_r_reg[7]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w2540_
	);
	LUT2 #(
		.INIT('h4)
	) name2009 (
		\text_in_r_reg[7]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w2541_
	);
	LUT2 #(
		.INIT('h2)
	) name2010 (
		\ld_r_reg/P0001 ,
		_w2540_,
		_w2542_
	);
	LUT2 #(
		.INIT('h4)
	) name2011 (
		_w2541_,
		_w2542_,
		_w2543_
	);
	LUT2 #(
		.INIT('h1)
	) name2012 (
		_w2539_,
		_w2543_,
		_w2544_
	);
	LUT2 #(
		.INIT('h4)
	) name2013 (
		\sa10_reg[2]/P0001 ,
		_w2093_,
		_w2545_
	);
	LUT2 #(
		.INIT('h8)
	) name2014 (
		\sa10_reg[4]/P0001 ,
		_w1585_,
		_w2546_
	);
	LUT2 #(
		.INIT('h8)
	) name2015 (
		\sa10_reg[2]/P0001 ,
		_w2546_,
		_w2547_
	);
	LUT2 #(
		.INIT('h1)
	) name2016 (
		_w2545_,
		_w2547_,
		_w2548_
	);
	LUT2 #(
		.INIT('h2)
	) name2017 (
		\sa10_reg[3]/P0001 ,
		_w2548_,
		_w2549_
	);
	LUT2 #(
		.INIT('h4)
	) name2018 (
		\sa10_reg[4]/P0001 ,
		_w1591_,
		_w2550_
	);
	LUT2 #(
		.INIT('h1)
	) name2019 (
		_w1654_,
		_w1731_,
		_w2551_
	);
	LUT2 #(
		.INIT('h4)
	) name2020 (
		_w2550_,
		_w2551_,
		_w2552_
	);
	LUT2 #(
		.INIT('h1)
	) name2021 (
		\sa10_reg[2]/P0001 ,
		_w2552_,
		_w2553_
	);
	LUT2 #(
		.INIT('h4)
	) name2022 (
		\sa10_reg[4]/P0001 ,
		_w1599_,
		_w2554_
	);
	LUT2 #(
		.INIT('h1)
	) name2023 (
		_w2156_,
		_w2554_,
		_w2555_
	);
	LUT2 #(
		.INIT('h4)
	) name2024 (
		_w2553_,
		_w2555_,
		_w2556_
	);
	LUT2 #(
		.INIT('h2)
	) name2025 (
		\sa10_reg[1]/P0001 ,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h8)
	) name2026 (
		_w1619_,
		_w1650_,
		_w2558_
	);
	LUT2 #(
		.INIT('h8)
	) name2027 (
		_w1650_,
		_w1669_,
		_w2559_
	);
	LUT2 #(
		.INIT('h2)
	) name2028 (
		\sa10_reg[2]/P0001 ,
		_w1682_,
		_w2560_
	);
	LUT2 #(
		.INIT('h4)
	) name2029 (
		_w2146_,
		_w2560_,
		_w2561_
	);
	LUT2 #(
		.INIT('h1)
	) name2030 (
		_w1616_,
		_w2558_,
		_w2562_
	);
	LUT2 #(
		.INIT('h4)
	) name2031 (
		_w2559_,
		_w2562_,
		_w2563_
	);
	LUT2 #(
		.INIT('h8)
	) name2032 (
		_w2561_,
		_w2563_,
		_w2564_
	);
	LUT2 #(
		.INIT('h8)
	) name2033 (
		_w1590_,
		_w1672_,
		_w2565_
	);
	LUT2 #(
		.INIT('h8)
	) name2034 (
		_w1637_,
		_w1681_,
		_w2566_
	);
	LUT2 #(
		.INIT('h8)
	) name2035 (
		\sa10_reg[5]/P0001 ,
		_w2566_,
		_w2567_
	);
	LUT2 #(
		.INIT('h1)
	) name2036 (
		\sa10_reg[2]/P0001 ,
		_w2128_,
		_w2568_
	);
	LUT2 #(
		.INIT('h4)
	) name2037 (
		_w2565_,
		_w2568_,
		_w2569_
	);
	LUT2 #(
		.INIT('h4)
	) name2038 (
		_w2567_,
		_w2569_,
		_w2570_
	);
	LUT2 #(
		.INIT('h1)
	) name2039 (
		_w2564_,
		_w2570_,
		_w2571_
	);
	LUT2 #(
		.INIT('h4)
	) name2040 (
		\sa10_reg[4]/P0001 ,
		_w1616_,
		_w2572_
	);
	LUT2 #(
		.INIT('h1)
	) name2041 (
		\sa10_reg[1]/P0001 ,
		_w1683_,
		_w2573_
	);
	LUT2 #(
		.INIT('h4)
	) name2042 (
		_w2572_,
		_w2573_,
		_w2574_
	);
	LUT2 #(
		.INIT('h4)
	) name2043 (
		_w2571_,
		_w2574_,
		_w2575_
	);
	LUT2 #(
		.INIT('h8)
	) name2044 (
		_w1593_,
		_w1661_,
		_w2576_
	);
	LUT2 #(
		.INIT('h8)
	) name2045 (
		\sa10_reg[4]/P0001 ,
		_w2576_,
		_w2577_
	);
	LUT2 #(
		.INIT('h2)
	) name2046 (
		\sa10_reg[1]/P0001 ,
		_w1665_,
		_w2578_
	);
	LUT2 #(
		.INIT('h4)
	) name2047 (
		_w2577_,
		_w2578_,
		_w2579_
	);
	LUT2 #(
		.INIT('h1)
	) name2048 (
		_w2575_,
		_w2579_,
		_w2580_
	);
	LUT2 #(
		.INIT('h4)
	) name2049 (
		\sa10_reg[7]/NET0131 ,
		_w1651_,
		_w2581_
	);
	LUT2 #(
		.INIT('h4)
	) name2050 (
		\sa10_reg[4]/P0001 ,
		_w1593_,
		_w2582_
	);
	LUT2 #(
		.INIT('h8)
	) name2051 (
		\sa10_reg[7]/NET0131 ,
		_w2098_,
		_w2583_
	);
	LUT2 #(
		.INIT('h1)
	) name2052 (
		_w2582_,
		_w2583_,
		_w2584_
	);
	LUT2 #(
		.INIT('h1)
	) name2053 (
		\sa10_reg[2]/P0001 ,
		_w2584_,
		_w2585_
	);
	LUT2 #(
		.INIT('h8)
	) name2054 (
		_w1637_,
		_w2112_,
		_w2586_
	);
	LUT2 #(
		.INIT('h2)
	) name2055 (
		\sa10_reg[1]/P0001 ,
		_w2586_,
		_w2587_
	);
	LUT2 #(
		.INIT('h4)
	) name2056 (
		_w1727_,
		_w2587_,
		_w2588_
	);
	LUT2 #(
		.INIT('h4)
	) name2057 (
		_w2581_,
		_w2588_,
		_w2589_
	);
	LUT2 #(
		.INIT('h4)
	) name2058 (
		_w2585_,
		_w2589_,
		_w2590_
	);
	LUT2 #(
		.INIT('h8)
	) name2059 (
		_w1666_,
		_w1703_,
		_w2591_
	);
	LUT2 #(
		.INIT('h1)
	) name2060 (
		\sa10_reg[1]/P0001 ,
		_w2591_,
		_w2592_
	);
	LUT2 #(
		.INIT('h8)
	) name2061 (
		\sa10_reg[3]/P0001 ,
		_w1626_,
		_w2593_
	);
	LUT2 #(
		.INIT('h8)
	) name2062 (
		_w1684_,
		_w2112_,
		_w2594_
	);
	LUT2 #(
		.INIT('h1)
	) name2063 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w2595_
	);
	LUT2 #(
		.INIT('h8)
	) name2064 (
		_w1626_,
		_w2595_,
		_w2596_
	);
	LUT2 #(
		.INIT('h1)
	) name2065 (
		_w2566_,
		_w2593_,
		_w2597_
	);
	LUT2 #(
		.INIT('h4)
	) name2066 (
		_w2596_,
		_w2597_,
		_w2598_
	);
	LUT2 #(
		.INIT('h4)
	) name2067 (
		_w2594_,
		_w2598_,
		_w2599_
	);
	LUT2 #(
		.INIT('h8)
	) name2068 (
		_w2592_,
		_w2599_,
		_w2600_
	);
	LUT2 #(
		.INIT('h1)
	) name2069 (
		_w2590_,
		_w2600_,
		_w2601_
	);
	LUT2 #(
		.INIT('h2)
	) name2070 (
		\sa10_reg[2]/P0001 ,
		_w1599_,
		_w2602_
	);
	LUT2 #(
		.INIT('h4)
	) name2071 (
		\sa10_reg[6]/NET0131 ,
		_w1627_,
		_w2603_
	);
	LUT2 #(
		.INIT('h1)
	) name2072 (
		_w1656_,
		_w1713_,
		_w2604_
	);
	LUT2 #(
		.INIT('h4)
	) name2073 (
		_w2603_,
		_w2604_,
		_w2605_
	);
	LUT2 #(
		.INIT('h8)
	) name2074 (
		_w2602_,
		_w2605_,
		_w2606_
	);
	LUT2 #(
		.INIT('h8)
	) name2075 (
		_w1608_,
		_w1681_,
		_w2607_
	);
	LUT2 #(
		.INIT('h8)
	) name2076 (
		_w1593_,
		_w1627_,
		_w2608_
	);
	LUT2 #(
		.INIT('h1)
	) name2077 (
		\sa10_reg[2]/P0001 ,
		_w2607_,
		_w2609_
	);
	LUT2 #(
		.INIT('h4)
	) name2078 (
		_w2608_,
		_w2609_,
		_w2610_
	);
	LUT2 #(
		.INIT('h4)
	) name2079 (
		_w1731_,
		_w2610_,
		_w2611_
	);
	LUT2 #(
		.INIT('h1)
	) name2080 (
		_w2606_,
		_w2611_,
		_w2612_
	);
	LUT2 #(
		.INIT('h1)
	) name2081 (
		_w2601_,
		_w2612_,
		_w2613_
	);
	LUT2 #(
		.INIT('h2)
	) name2082 (
		\sa10_reg[0]/P0001 ,
		_w2613_,
		_w2614_
	);
	LUT2 #(
		.INIT('h8)
	) name2083 (
		\sa10_reg[5]/P0001 ,
		_w2147_,
		_w2615_
	);
	LUT2 #(
		.INIT('h1)
	) name2084 (
		_w1627_,
		_w1722_,
		_w2616_
	);
	LUT2 #(
		.INIT('h2)
	) name2085 (
		_w1614_,
		_w2616_,
		_w2617_
	);
	LUT2 #(
		.INIT('h1)
	) name2086 (
		\sa10_reg[1]/P0001 ,
		_w2547_,
		_w2618_
	);
	LUT2 #(
		.INIT('h1)
	) name2087 (
		_w2615_,
		_w2617_,
		_w2619_
	);
	LUT2 #(
		.INIT('h8)
	) name2088 (
		_w2618_,
		_w2619_,
		_w2620_
	);
	LUT2 #(
		.INIT('h8)
	) name2089 (
		\sa10_reg[5]/P0001 ,
		_w1593_,
		_w2621_
	);
	LUT2 #(
		.INIT('h8)
	) name2090 (
		\sa10_reg[2]/P0001 ,
		_w2621_,
		_w2622_
	);
	LUT2 #(
		.INIT('h8)
	) name2091 (
		\sa10_reg[4]/P0001 ,
		_w1608_,
		_w2623_
	);
	LUT2 #(
		.INIT('h8)
	) name2092 (
		_w1661_,
		_w2623_,
		_w2624_
	);
	LUT2 #(
		.INIT('h8)
	) name2093 (
		_w1637_,
		_w1650_,
		_w2625_
	);
	LUT2 #(
		.INIT('h4)
	) name2094 (
		_w1627_,
		_w1699_,
		_w2626_
	);
	LUT2 #(
		.INIT('h1)
	) name2095 (
		_w2625_,
		_w2626_,
		_w2627_
	);
	LUT2 #(
		.INIT('h1)
	) name2096 (
		\sa10_reg[2]/P0001 ,
		_w2627_,
		_w2628_
	);
	LUT2 #(
		.INIT('h2)
	) name2097 (
		\sa10_reg[1]/P0001 ,
		_w1595_,
		_w2629_
	);
	LUT2 #(
		.INIT('h4)
	) name2098 (
		_w2622_,
		_w2629_,
		_w2630_
	);
	LUT2 #(
		.INIT('h4)
	) name2099 (
		_w2624_,
		_w2630_,
		_w2631_
	);
	LUT2 #(
		.INIT('h4)
	) name2100 (
		_w2628_,
		_w2631_,
		_w2632_
	);
	LUT2 #(
		.INIT('h1)
	) name2101 (
		_w2620_,
		_w2632_,
		_w2633_
	);
	LUT2 #(
		.INIT('h8)
	) name2102 (
		_w1612_,
		_w1672_,
		_w2634_
	);
	LUT2 #(
		.INIT('h4)
	) name2103 (
		\sa10_reg[2]/P0001 ,
		_w2634_,
		_w2635_
	);
	LUT2 #(
		.INIT('h8)
	) name2104 (
		_w1607_,
		_w1722_,
		_w2636_
	);
	LUT2 #(
		.INIT('h1)
	) name2105 (
		_w2101_,
		_w2636_,
		_w2637_
	);
	LUT2 #(
		.INIT('h4)
	) name2106 (
		_w2635_,
		_w2637_,
		_w2638_
	);
	LUT2 #(
		.INIT('h1)
	) name2107 (
		\sa10_reg[3]/P0001 ,
		_w2638_,
		_w2639_
	);
	LUT2 #(
		.INIT('h8)
	) name2108 (
		\sa10_reg[2]/P0001 ,
		_w2180_,
		_w2640_
	);
	LUT2 #(
		.INIT('h1)
	) name2109 (
		_w2639_,
		_w2640_,
		_w2641_
	);
	LUT2 #(
		.INIT('h4)
	) name2110 (
		_w2633_,
		_w2641_,
		_w2642_
	);
	LUT2 #(
		.INIT('h1)
	) name2111 (
		\sa10_reg[0]/P0001 ,
		_w2642_,
		_w2643_
	);
	LUT2 #(
		.INIT('h1)
	) name2112 (
		_w2549_,
		_w2557_,
		_w2644_
	);
	LUT2 #(
		.INIT('h4)
	) name2113 (
		_w2580_,
		_w2644_,
		_w2645_
	);
	LUT2 #(
		.INIT('h1)
	) name2114 (
		_w2614_,
		_w2643_,
		_w2646_
	);
	LUT2 #(
		.INIT('h8)
	) name2115 (
		_w2645_,
		_w2646_,
		_w2647_
	);
	LUT2 #(
		.INIT('h1)
	) name2116 (
		_w1319_,
		_w2206_,
		_w2648_
	);
	LUT2 #(
		.INIT('h1)
	) name2117 (
		\sa03_reg[2]/P0001 ,
		_w2648_,
		_w2649_
	);
	LUT2 #(
		.INIT('h8)
	) name2118 (
		_w1330_,
		_w1384_,
		_w2650_
	);
	LUT2 #(
		.INIT('h2)
	) name2119 (
		\sa03_reg[1]/P0001 ,
		_w2650_,
		_w2651_
	);
	LUT2 #(
		.INIT('h4)
	) name2120 (
		_w1417_,
		_w2651_,
		_w2652_
	);
	LUT2 #(
		.INIT('h4)
	) name2121 (
		_w1461_,
		_w2652_,
		_w2653_
	);
	LUT2 #(
		.INIT('h4)
	) name2122 (
		_w2649_,
		_w2653_,
		_w2654_
	);
	LUT2 #(
		.INIT('h8)
	) name2123 (
		_w1330_,
		_w1398_,
		_w2655_
	);
	LUT2 #(
		.INIT('h1)
	) name2124 (
		\sa03_reg[1]/P0001 ,
		_w2655_,
		_w2656_
	);
	LUT2 #(
		.INIT('h8)
	) name2125 (
		_w2215_,
		_w2218_,
		_w2657_
	);
	LUT2 #(
		.INIT('h8)
	) name2126 (
		_w1375_,
		_w1384_,
		_w2658_
	);
	LUT2 #(
		.INIT('h1)
	) name2127 (
		\sa03_reg[3]/P0001 ,
		_w1515_,
		_w2659_
	);
	LUT2 #(
		.INIT('h2)
	) name2128 (
		_w1339_,
		_w2659_,
		_w2660_
	);
	LUT2 #(
		.INIT('h2)
	) name2129 (
		_w2656_,
		_w2657_,
		_w2661_
	);
	LUT2 #(
		.INIT('h1)
	) name2130 (
		_w2658_,
		_w2660_,
		_w2662_
	);
	LUT2 #(
		.INIT('h8)
	) name2131 (
		_w2661_,
		_w2662_,
		_w2663_
	);
	LUT2 #(
		.INIT('h1)
	) name2132 (
		_w2654_,
		_w2663_,
		_w2664_
	);
	LUT2 #(
		.INIT('h8)
	) name2133 (
		_w1324_,
		_w1332_,
		_w2665_
	);
	LUT2 #(
		.INIT('h4)
	) name2134 (
		\sa03_reg[3]/P0001 ,
		_w1341_,
		_w2666_
	);
	LUT2 #(
		.INIT('h1)
	) name2135 (
		_w1424_,
		_w2665_,
		_w2667_
	);
	LUT2 #(
		.INIT('h4)
	) name2136 (
		_w2666_,
		_w2667_,
		_w2668_
	);
	LUT2 #(
		.INIT('h8)
	) name2137 (
		_w1562_,
		_w2668_,
		_w2669_
	);
	LUT2 #(
		.INIT('h4)
	) name2138 (
		\sa03_reg[7]/NET0131 ,
		_w1541_,
		_w2670_
	);
	LUT2 #(
		.INIT('h4)
	) name2139 (
		_w1447_,
		_w1538_,
		_w2671_
	);
	LUT2 #(
		.INIT('h4)
	) name2140 (
		_w2670_,
		_w2671_,
		_w2672_
	);
	LUT2 #(
		.INIT('h1)
	) name2141 (
		_w2669_,
		_w2672_,
		_w2673_
	);
	LUT2 #(
		.INIT('h1)
	) name2142 (
		_w2664_,
		_w2673_,
		_w2674_
	);
	LUT2 #(
		.INIT('h2)
	) name2143 (
		\sa03_reg[0]/P0001 ,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h4)
	) name2144 (
		\sa03_reg[3]/P0001 ,
		_w1416_,
		_w2676_
	);
	LUT2 #(
		.INIT('h2)
	) name2145 (
		_w1449_,
		_w2252_,
		_w2677_
	);
	LUT2 #(
		.INIT('h8)
	) name2146 (
		_w1327_,
		_w1455_,
		_w2678_
	);
	LUT2 #(
		.INIT('h8)
	) name2147 (
		_w1317_,
		_w1355_,
		_w2679_
	);
	LUT2 #(
		.INIT('h2)
	) name2148 (
		\sa03_reg[2]/P0001 ,
		_w2266_,
		_w2680_
	);
	LUT2 #(
		.INIT('h4)
	) name2149 (
		_w2677_,
		_w2680_,
		_w2681_
	);
	LUT2 #(
		.INIT('h1)
	) name2150 (
		_w2678_,
		_w2679_,
		_w2682_
	);
	LUT2 #(
		.INIT('h8)
	) name2151 (
		_w2681_,
		_w2682_,
		_w2683_
	);
	LUT2 #(
		.INIT('h8)
	) name2152 (
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2684_
	);
	LUT2 #(
		.INIT('h8)
	) name2153 (
		_w1454_,
		_w2684_,
		_w2685_
	);
	LUT2 #(
		.INIT('h1)
	) name2154 (
		\sa03_reg[2]/P0001 ,
		_w1328_,
		_w2686_
	);
	LUT2 #(
		.INIT('h4)
	) name2155 (
		_w2216_,
		_w2686_,
		_w2687_
	);
	LUT2 #(
		.INIT('h4)
	) name2156 (
		_w2685_,
		_w2687_,
		_w2688_
	);
	LUT2 #(
		.INIT('h1)
	) name2157 (
		_w2683_,
		_w2688_,
		_w2689_
	);
	LUT2 #(
		.INIT('h1)
	) name2158 (
		\sa03_reg[1]/P0001 ,
		_w1400_,
		_w2690_
	);
	LUT2 #(
		.INIT('h4)
	) name2159 (
		_w2676_,
		_w2690_,
		_w2691_
	);
	LUT2 #(
		.INIT('h4)
	) name2160 (
		_w2689_,
		_w2691_,
		_w2692_
	);
	LUT2 #(
		.INIT('h8)
	) name2161 (
		_w1367_,
		_w1424_,
		_w2693_
	);
	LUT2 #(
		.INIT('h8)
	) name2162 (
		_w1436_,
		_w1482_,
		_w2694_
	);
	LUT2 #(
		.INIT('h1)
	) name2163 (
		_w1354_,
		_w1534_,
		_w2695_
	);
	LUT2 #(
		.INIT('h4)
	) name2164 (
		_w2670_,
		_w2695_,
		_w2696_
	);
	LUT2 #(
		.INIT('h1)
	) name2165 (
		\sa03_reg[2]/P0001 ,
		_w2696_,
		_w2697_
	);
	LUT2 #(
		.INIT('h2)
	) name2166 (
		\sa03_reg[1]/P0001 ,
		_w1522_,
		_w2698_
	);
	LUT2 #(
		.INIT('h1)
	) name2167 (
		_w2249_,
		_w2693_,
		_w2699_
	);
	LUT2 #(
		.INIT('h4)
	) name2168 (
		_w2694_,
		_w2699_,
		_w2700_
	);
	LUT2 #(
		.INIT('h8)
	) name2169 (
		_w2698_,
		_w2700_,
		_w2701_
	);
	LUT2 #(
		.INIT('h4)
	) name2170 (
		_w2697_,
		_w2701_,
		_w2702_
	);
	LUT2 #(
		.INIT('h1)
	) name2171 (
		_w2692_,
		_w2702_,
		_w2703_
	);
	LUT2 #(
		.INIT('h4)
	) name2172 (
		\sa03_reg[3]/P0001 ,
		_w1431_,
		_w2704_
	);
	LUT2 #(
		.INIT('h1)
	) name2173 (
		_w2288_,
		_w2704_,
		_w2705_
	);
	LUT2 #(
		.INIT('h2)
	) name2174 (
		\sa03_reg[2]/P0001 ,
		_w2705_,
		_w2706_
	);
	LUT2 #(
		.INIT('h4)
	) name2175 (
		\sa03_reg[2]/P0001 ,
		_w1397_,
		_w2707_
	);
	LUT2 #(
		.INIT('h1)
	) name2176 (
		_w1416_,
		_w2707_,
		_w2708_
	);
	LUT2 #(
		.INIT('h1)
	) name2177 (
		\sa03_reg[3]/P0001 ,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h8)
	) name2178 (
		\sa03_reg[5]/P0001 ,
		_w1332_,
		_w2710_
	);
	LUT2 #(
		.INIT('h4)
	) name2179 (
		_w1423_,
		_w2710_,
		_w2711_
	);
	LUT2 #(
		.INIT('h8)
	) name2180 (
		_w1330_,
		_w1355_,
		_w2712_
	);
	LUT2 #(
		.INIT('h1)
	) name2181 (
		_w2711_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('h1)
	) name2182 (
		\sa03_reg[2]/P0001 ,
		_w2713_,
		_w2714_
	);
	LUT2 #(
		.INIT('h8)
	) name2183 (
		\sa03_reg[2]/P0001 ,
		_w1435_,
		_w2715_
	);
	LUT2 #(
		.INIT('h8)
	) name2184 (
		_w1367_,
		_w1381_,
		_w2716_
	);
	LUT2 #(
		.INIT('h2)
	) name2185 (
		\sa03_reg[1]/P0001 ,
		_w1399_,
		_w2717_
	);
	LUT2 #(
		.INIT('h4)
	) name2186 (
		_w2715_,
		_w2717_,
		_w2718_
	);
	LUT2 #(
		.INIT('h4)
	) name2187 (
		_w2716_,
		_w2718_,
		_w2719_
	);
	LUT2 #(
		.INIT('h4)
	) name2188 (
		_w2714_,
		_w2719_,
		_w2720_
	);
	LUT2 #(
		.INIT('h1)
	) name2189 (
		\sa03_reg[2]/P0001 ,
		_w2289_,
		_w2721_
	);
	LUT2 #(
		.INIT('h2)
	) name2190 (
		\sa03_reg[2]/P0001 ,
		_w2260_,
		_w2722_
	);
	LUT2 #(
		.INIT('h4)
	) name2191 (
		_w1460_,
		_w2722_,
		_w2723_
	);
	LUT2 #(
		.INIT('h1)
	) name2192 (
		_w2721_,
		_w2723_,
		_w2724_
	);
	LUT2 #(
		.INIT('h1)
	) name2193 (
		\sa03_reg[1]/P0001 ,
		_w1563_,
		_w2725_
	);
	LUT2 #(
		.INIT('h4)
	) name2194 (
		_w2724_,
		_w2725_,
		_w2726_
	);
	LUT2 #(
		.INIT('h1)
	) name2195 (
		_w2720_,
		_w2726_,
		_w2727_
	);
	LUT2 #(
		.INIT('h1)
	) name2196 (
		_w2706_,
		_w2709_,
		_w2728_
	);
	LUT2 #(
		.INIT('h4)
	) name2197 (
		_w2727_,
		_w2728_,
		_w2729_
	);
	LUT2 #(
		.INIT('h1)
	) name2198 (
		\sa03_reg[0]/P0001 ,
		_w2729_,
		_w2730_
	);
	LUT2 #(
		.INIT('h1)
	) name2199 (
		\sa03_reg[2]/P0001 ,
		_w2200_,
		_w2731_
	);
	LUT2 #(
		.INIT('h2)
	) name2200 (
		\sa03_reg[3]/P0001 ,
		_w2722_,
		_w2732_
	);
	LUT2 #(
		.INIT('h4)
	) name2201 (
		_w2731_,
		_w2732_,
		_w2733_
	);
	LUT2 #(
		.INIT('h1)
	) name2202 (
		_w2703_,
		_w2733_,
		_w2734_
	);
	LUT2 #(
		.INIT('h4)
	) name2203 (
		_w2675_,
		_w2734_,
		_w2735_
	);
	LUT2 #(
		.INIT('h4)
	) name2204 (
		_w2730_,
		_w2735_,
		_w2736_
	);
	LUT2 #(
		.INIT('h2)
	) name2205 (
		_w2647_,
		_w2736_,
		_w2737_
	);
	LUT2 #(
		.INIT('h4)
	) name2206 (
		_w2647_,
		_w2736_,
		_w2738_
	);
	LUT2 #(
		.INIT('h1)
	) name2207 (
		_w2737_,
		_w2738_,
		_w2739_
	);
	LUT2 #(
		.INIT('h4)
	) name2208 (
		\sa10_reg[4]/P0001 ,
		_w1629_,
		_w2740_
	);
	LUT2 #(
		.INIT('h4)
	) name2209 (
		_w1612_,
		_w1634_,
		_w2741_
	);
	LUT2 #(
		.INIT('h1)
	) name2210 (
		_w1726_,
		_w2741_,
		_w2742_
	);
	LUT2 #(
		.INIT('h2)
	) name2211 (
		\sa10_reg[1]/P0001 ,
		_w2742_,
		_w2743_
	);
	LUT2 #(
		.INIT('h1)
	) name2212 (
		_w1682_,
		_w2608_,
		_w2744_
	);
	LUT2 #(
		.INIT('h4)
	) name2213 (
		_w2740_,
		_w2744_,
		_w2745_
	);
	LUT2 #(
		.INIT('h4)
	) name2214 (
		_w2743_,
		_w2745_,
		_w2746_
	);
	LUT2 #(
		.INIT('h1)
	) name2215 (
		\sa10_reg[2]/P0001 ,
		_w2746_,
		_w2747_
	);
	LUT2 #(
		.INIT('h8)
	) name2216 (
		\sa10_reg[7]/NET0131 ,
		_w1584_,
		_w2748_
	);
	LUT2 #(
		.INIT('h8)
	) name2217 (
		_w1597_,
		_w1627_,
		_w2749_
	);
	LUT2 #(
		.INIT('h1)
	) name2218 (
		_w1631_,
		_w2749_,
		_w2750_
	);
	LUT2 #(
		.INIT('h1)
	) name2219 (
		_w2581_,
		_w2748_,
		_w2751_
	);
	LUT2 #(
		.INIT('h8)
	) name2220 (
		_w2750_,
		_w2751_,
		_w2752_
	);
	LUT2 #(
		.INIT('h2)
	) name2221 (
		\sa10_reg[1]/P0001 ,
		_w2752_,
		_w2753_
	);
	LUT2 #(
		.INIT('h8)
	) name2222 (
		_w1593_,
		_w1668_,
		_w2754_
	);
	LUT2 #(
		.INIT('h4)
	) name2223 (
		\sa10_reg[5]/P0001 ,
		_w2754_,
		_w2755_
	);
	LUT2 #(
		.INIT('h1)
	) name2224 (
		_w1592_,
		_w2755_,
		_w2756_
	);
	LUT2 #(
		.INIT('h2)
	) name2225 (
		\sa10_reg[2]/P0001 ,
		_w2756_,
		_w2757_
	);
	LUT2 #(
		.INIT('h8)
	) name2226 (
		_w1627_,
		_w2621_,
		_w2758_
	);
	LUT2 #(
		.INIT('h1)
	) name2227 (
		_w1599_,
		_w2621_,
		_w2759_
	);
	LUT2 #(
		.INIT('h1)
	) name2228 (
		\sa10_reg[2]/P0001 ,
		_w2759_,
		_w2760_
	);
	LUT2 #(
		.INIT('h8)
	) name2229 (
		_w1664_,
		_w1703_,
		_w2761_
	);
	LUT2 #(
		.INIT('h1)
	) name2230 (
		_w1682_,
		_w2636_,
		_w2762_
	);
	LUT2 #(
		.INIT('h4)
	) name2231 (
		_w1592_,
		_w2762_,
		_w2763_
	);
	LUT2 #(
		.INIT('h4)
	) name2232 (
		_w2761_,
		_w2763_,
		_w2764_
	);
	LUT2 #(
		.INIT('h4)
	) name2233 (
		_w2760_,
		_w2764_,
		_w2765_
	);
	LUT2 #(
		.INIT('h1)
	) name2234 (
		\sa10_reg[1]/P0001 ,
		_w2765_,
		_w2766_
	);
	LUT2 #(
		.INIT('h1)
	) name2235 (
		_w2635_,
		_w2758_,
		_w2767_
	);
	LUT2 #(
		.INIT('h4)
	) name2236 (
		_w2757_,
		_w2767_,
		_w2768_
	);
	LUT2 #(
		.INIT('h4)
	) name2237 (
		_w2753_,
		_w2768_,
		_w2769_
	);
	LUT2 #(
		.INIT('h4)
	) name2238 (
		_w2747_,
		_w2769_,
		_w2770_
	);
	LUT2 #(
		.INIT('h4)
	) name2239 (
		_w2766_,
		_w2770_,
		_w2771_
	);
	LUT2 #(
		.INIT('h2)
	) name2240 (
		\sa10_reg[0]/P0001 ,
		_w2771_,
		_w2772_
	);
	LUT2 #(
		.INIT('h1)
	) name2241 (
		_w2168_,
		_w2593_,
		_w2773_
	);
	LUT2 #(
		.INIT('h2)
	) name2242 (
		\sa10_reg[2]/P0001 ,
		_w2773_,
		_w2774_
	);
	LUT2 #(
		.INIT('h1)
	) name2243 (
		_w1584_,
		_w2754_,
		_w2775_
	);
	LUT2 #(
		.INIT('h1)
	) name2244 (
		\sa10_reg[2]/P0001 ,
		_w2775_,
		_w2776_
	);
	LUT2 #(
		.INIT('h8)
	) name2245 (
		_w1594_,
		_w1626_,
		_w2777_
	);
	LUT2 #(
		.INIT('h8)
	) name2246 (
		_w1597_,
		_w1666_,
		_w2778_
	);
	LUT2 #(
		.INIT('h1)
	) name2247 (
		_w1638_,
		_w2185_,
		_w2779_
	);
	LUT2 #(
		.INIT('h1)
	) name2248 (
		_w2565_,
		_w2777_,
		_w2780_
	);
	LUT2 #(
		.INIT('h4)
	) name2249 (
		_w2778_,
		_w2780_,
		_w2781_
	);
	LUT2 #(
		.INIT('h4)
	) name2250 (
		_w2179_,
		_w2779_,
		_w2782_
	);
	LUT2 #(
		.INIT('h8)
	) name2251 (
		_w2781_,
		_w2782_,
		_w2783_
	);
	LUT2 #(
		.INIT('h4)
	) name2252 (
		_w2776_,
		_w2783_,
		_w2784_
	);
	LUT2 #(
		.INIT('h4)
	) name2253 (
		_w2774_,
		_w2784_,
		_w2785_
	);
	LUT2 #(
		.INIT('h2)
	) name2254 (
		\sa10_reg[1]/P0001 ,
		_w2785_,
		_w2786_
	);
	LUT2 #(
		.INIT('h4)
	) name2255 (
		\sa10_reg[3]/P0001 ,
		_w1618_,
		_w2787_
	);
	LUT2 #(
		.INIT('h1)
	) name2256 (
		_w1601_,
		_w2787_,
		_w2788_
	);
	LUT2 #(
		.INIT('h1)
	) name2257 (
		_w1668_,
		_w2788_,
		_w2789_
	);
	LUT2 #(
		.INIT('h4)
	) name2258 (
		\sa10_reg[4]/P0001 ,
		_w1614_,
		_w2790_
	);
	LUT2 #(
		.INIT('h1)
	) name2259 (
		_w2777_,
		_w2790_,
		_w2791_
	);
	LUT2 #(
		.INIT('h4)
	) name2260 (
		_w2789_,
		_w2791_,
		_w2792_
	);
	LUT2 #(
		.INIT('h2)
	) name2261 (
		\sa10_reg[2]/P0001 ,
		_w2792_,
		_w2793_
	);
	LUT2 #(
		.INIT('h1)
	) name2262 (
		_w1651_,
		_w1711_,
		_w2794_
	);
	LUT2 #(
		.INIT('h2)
	) name2263 (
		\sa10_reg[7]/NET0131 ,
		_w2794_,
		_w2795_
	);
	LUT2 #(
		.INIT('h1)
	) name2264 (
		_w1698_,
		_w2603_,
		_w2796_
	);
	LUT2 #(
		.INIT('h2)
	) name2265 (
		_w1722_,
		_w2796_,
		_w2797_
	);
	LUT2 #(
		.INIT('h1)
	) name2266 (
		_w2795_,
		_w2797_,
		_w2798_
	);
	LUT2 #(
		.INIT('h1)
	) name2267 (
		\sa10_reg[1]/P0001 ,
		_w2798_,
		_w2799_
	);
	LUT2 #(
		.INIT('h4)
	) name2268 (
		\sa10_reg[2]/P0001 ,
		_w1613_,
		_w2800_
	);
	LUT2 #(
		.INIT('h1)
	) name2269 (
		_w1602_,
		_w2800_,
		_w2801_
	);
	LUT2 #(
		.INIT('h4)
	) name2270 (
		_w1611_,
		_w2801_,
		_w2802_
	);
	LUT2 #(
		.INIT('h4)
	) name2271 (
		_w2799_,
		_w2802_,
		_w2803_
	);
	LUT2 #(
		.INIT('h4)
	) name2272 (
		_w2793_,
		_w2803_,
		_w2804_
	);
	LUT2 #(
		.INIT('h4)
	) name2273 (
		_w2786_,
		_w2804_,
		_w2805_
	);
	LUT2 #(
		.INIT('h1)
	) name2274 (
		\sa10_reg[0]/P0001 ,
		_w2805_,
		_w2806_
	);
	LUT2 #(
		.INIT('h8)
	) name2275 (
		\sa10_reg[5]/P0001 ,
		_w2761_,
		_w2807_
	);
	LUT2 #(
		.INIT('h8)
	) name2276 (
		_w1582_,
		_w2110_,
		_w2808_
	);
	LUT2 #(
		.INIT('h8)
	) name2277 (
		\sa10_reg[6]/NET0131 ,
		_w1626_,
		_w2809_
	);
	LUT2 #(
		.INIT('h1)
	) name2278 (
		_w1593_,
		_w1597_,
		_w2810_
	);
	LUT2 #(
		.INIT('h1)
	) name2279 (
		\sa10_reg[5]/P0001 ,
		_w2810_,
		_w2811_
	);
	LUT2 #(
		.INIT('h1)
	) name2280 (
		_w2809_,
		_w2811_,
		_w2812_
	);
	LUT2 #(
		.INIT('h8)
	) name2281 (
		\sa10_reg[2]/P0001 ,
		_w1583_,
		_w2813_
	);
	LUT2 #(
		.INIT('h4)
	) name2282 (
		_w2812_,
		_w2813_,
		_w2814_
	);
	LUT2 #(
		.INIT('h1)
	) name2283 (
		_w1730_,
		_w2808_,
		_w2815_
	);
	LUT2 #(
		.INIT('h4)
	) name2284 (
		_w2814_,
		_w2815_,
		_w2816_
	);
	LUT2 #(
		.INIT('h1)
	) name2285 (
		\sa10_reg[1]/P0001 ,
		_w2816_,
		_w2817_
	);
	LUT2 #(
		.INIT('h8)
	) name2286 (
		_w1661_,
		_w2168_,
		_w2818_
	);
	LUT2 #(
		.INIT('h8)
	) name2287 (
		_w1598_,
		_w2790_,
		_w2819_
	);
	LUT2 #(
		.INIT('h1)
	) name2288 (
		_w2800_,
		_w2819_,
		_w2820_
	);
	LUT2 #(
		.INIT('h4)
	) name2289 (
		_w2818_,
		_w2820_,
		_w2821_
	);
	LUT2 #(
		.INIT('h2)
	) name2290 (
		\sa10_reg[1]/P0001 ,
		_w2821_,
		_w2822_
	);
	LUT2 #(
		.INIT('h1)
	) name2291 (
		_w1727_,
		_w2565_,
		_w2823_
	);
	LUT2 #(
		.INIT('h1)
	) name2292 (
		\sa10_reg[2]/P0001 ,
		_w2823_,
		_w2824_
	);
	LUT2 #(
		.INIT('h1)
	) name2293 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[2]/P0001 ,
		_w2825_
	);
	LUT2 #(
		.INIT('h8)
	) name2294 (
		_w1626_,
		_w1668_,
		_w2826_
	);
	LUT2 #(
		.INIT('h1)
	) name2295 (
		_w2634_,
		_w2826_,
		_w2827_
	);
	LUT2 #(
		.INIT('h4)
	) name2296 (
		_w1683_,
		_w2827_,
		_w2828_
	);
	LUT2 #(
		.INIT('h2)
	) name2297 (
		_w2825_,
		_w2828_,
		_w2829_
	);
	LUT2 #(
		.INIT('h1)
	) name2298 (
		_w2807_,
		_w2824_,
		_w2830_
	);
	LUT2 #(
		.INIT('h4)
	) name2299 (
		_w2829_,
		_w2830_,
		_w2831_
	);
	LUT2 #(
		.INIT('h4)
	) name2300 (
		_w2822_,
		_w2831_,
		_w2832_
	);
	LUT2 #(
		.INIT('h4)
	) name2301 (
		_w2817_,
		_w2832_,
		_w2833_
	);
	LUT2 #(
		.INIT('h4)
	) name2302 (
		_w2772_,
		_w2833_,
		_w2834_
	);
	LUT2 #(
		.INIT('h4)
	) name2303 (
		_w2806_,
		_w2834_,
		_w2835_
	);
	LUT2 #(
		.INIT('h1)
	) name2304 (
		_w1750_,
		_w2436_,
		_w2836_
	);
	LUT2 #(
		.INIT('h2)
	) name2305 (
		\sa21_reg[2]/P0001 ,
		_w2836_,
		_w2837_
	);
	LUT2 #(
		.INIT('h8)
	) name2306 (
		_w1757_,
		_w1758_,
		_w2838_
	);
	LUT2 #(
		.INIT('h8)
	) name2307 (
		\sa21_reg[4]/P0001 ,
		_w1750_,
		_w2839_
	);
	LUT2 #(
		.INIT('h1)
	) name2308 (
		_w1764_,
		_w1838_,
		_w2840_
	);
	LUT2 #(
		.INIT('h1)
	) name2309 (
		\sa21_reg[4]/P0001 ,
		_w2840_,
		_w2841_
	);
	LUT2 #(
		.INIT('h8)
	) name2310 (
		\sa21_reg[3]/P0001 ,
		_w1763_,
		_w2842_
	);
	LUT2 #(
		.INIT('h4)
	) name2311 (
		\sa21_reg[3]/P0001 ,
		_w1775_,
		_w2843_
	);
	LUT2 #(
		.INIT('h1)
	) name2312 (
		_w1774_,
		_w2842_,
		_w2844_
	);
	LUT2 #(
		.INIT('h4)
	) name2313 (
		_w2843_,
		_w2844_,
		_w2845_
	);
	LUT2 #(
		.INIT('h1)
	) name2314 (
		\sa21_reg[2]/P0001 ,
		_w2845_,
		_w2846_
	);
	LUT2 #(
		.INIT('h1)
	) name2315 (
		_w2502_,
		_w2838_,
		_w2847_
	);
	LUT2 #(
		.INIT('h4)
	) name2316 (
		_w2839_,
		_w2847_,
		_w2848_
	);
	LUT2 #(
		.INIT('h4)
	) name2317 (
		_w2841_,
		_w2848_,
		_w2849_
	);
	LUT2 #(
		.INIT('h4)
	) name2318 (
		_w2837_,
		_w2849_,
		_w2850_
	);
	LUT2 #(
		.INIT('h4)
	) name2319 (
		_w2846_,
		_w2850_,
		_w2851_
	);
	LUT2 #(
		.INIT('h2)
	) name2320 (
		\sa21_reg[1]/P0001 ,
		_w2851_,
		_w2852_
	);
	LUT2 #(
		.INIT('h8)
	) name2321 (
		_w1816_,
		_w1837_,
		_w2853_
	);
	LUT2 #(
		.INIT('h1)
	) name2322 (
		_w2426_,
		_w2478_,
		_w2854_
	);
	LUT2 #(
		.INIT('h1)
	) name2323 (
		\sa21_reg[3]/P0001 ,
		_w2854_,
		_w2855_
	);
	LUT2 #(
		.INIT('h2)
	) name2324 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w2856_
	);
	LUT2 #(
		.INIT('h8)
	) name2325 (
		\sa21_reg[3]/P0001 ,
		_w1832_,
		_w2857_
	);
	LUT2 #(
		.INIT('h8)
	) name2326 (
		_w2856_,
		_w2857_,
		_w2858_
	);
	LUT2 #(
		.INIT('h1)
	) name2327 (
		_w2853_,
		_w2858_,
		_w2859_
	);
	LUT2 #(
		.INIT('h4)
	) name2328 (
		_w2855_,
		_w2859_,
		_w2860_
	);
	LUT2 #(
		.INIT('h1)
	) name2329 (
		\sa21_reg[1]/P0001 ,
		_w2860_,
		_w2861_
	);
	LUT2 #(
		.INIT('h4)
	) name2330 (
		\sa21_reg[4]/P0001 ,
		_w1841_,
		_w2862_
	);
	LUT2 #(
		.INIT('h2)
	) name2331 (
		\sa21_reg[3]/P0001 ,
		_w1850_,
		_w2863_
	);
	LUT2 #(
		.INIT('h8)
	) name2332 (
		\sa21_reg[4]/P0001 ,
		_w1799_,
		_w2864_
	);
	LUT2 #(
		.INIT('h8)
	) name2333 (
		_w1758_,
		_w2864_,
		_w2865_
	);
	LUT2 #(
		.INIT('h1)
	) name2334 (
		_w2862_,
		_w2865_,
		_w2866_
	);
	LUT2 #(
		.INIT('h4)
	) name2335 (
		_w2863_,
		_w2866_,
		_w2867_
	);
	LUT2 #(
		.INIT('h2)
	) name2336 (
		\sa21_reg[2]/P0001 ,
		_w2867_,
		_w2868_
	);
	LUT2 #(
		.INIT('h8)
	) name2337 (
		_w1764_,
		_w2455_,
		_w2869_
	);
	LUT2 #(
		.INIT('h1)
	) name2338 (
		_w1786_,
		_w2869_,
		_w2870_
	);
	LUT2 #(
		.INIT('h4)
	) name2339 (
		_w1798_,
		_w2870_,
		_w2871_
	);
	LUT2 #(
		.INIT('h4)
	) name2340 (
		_w2868_,
		_w2871_,
		_w2872_
	);
	LUT2 #(
		.INIT('h4)
	) name2341 (
		_w2861_,
		_w2872_,
		_w2873_
	);
	LUT2 #(
		.INIT('h4)
	) name2342 (
		_w2852_,
		_w2873_,
		_w2874_
	);
	LUT2 #(
		.INIT('h1)
	) name2343 (
		\sa21_reg[0]/P0001 ,
		_w2874_,
		_w2875_
	);
	LUT2 #(
		.INIT('h8)
	) name2344 (
		_w1753_,
		_w1854_,
		_w2876_
	);
	LUT2 #(
		.INIT('h1)
	) name2345 (
		_w2429_,
		_w2876_,
		_w2877_
	);
	LUT2 #(
		.INIT('h1)
	) name2346 (
		_w1795_,
		_w1833_,
		_w2878_
	);
	LUT2 #(
		.INIT('h4)
	) name2347 (
		_w1867_,
		_w2878_,
		_w2879_
	);
	LUT2 #(
		.INIT('h2)
	) name2348 (
		\sa21_reg[1]/P0001 ,
		_w2879_,
		_w2880_
	);
	LUT2 #(
		.INIT('h4)
	) name2349 (
		_w1879_,
		_w2877_,
		_w2881_
	);
	LUT2 #(
		.INIT('h4)
	) name2350 (
		_w2880_,
		_w2881_,
		_w2882_
	);
	LUT2 #(
		.INIT('h1)
	) name2351 (
		\sa21_reg[2]/P0001 ,
		_w2882_,
		_w2883_
	);
	LUT2 #(
		.INIT('h8)
	) name2352 (
		\sa21_reg[3]/P0001 ,
		_w2492_,
		_w2884_
	);
	LUT2 #(
		.INIT('h1)
	) name2353 (
		_w1759_,
		_w2884_,
		_w2885_
	);
	LUT2 #(
		.INIT('h2)
	) name2354 (
		\sa21_reg[2]/P0001 ,
		_w2885_,
		_w2886_
	);
	LUT2 #(
		.INIT('h8)
	) name2355 (
		_w1877_,
		_w2425_,
		_w2887_
	);
	LUT2 #(
		.INIT('h1)
	) name2356 (
		_w2429_,
		_w2449_,
		_w2888_
	);
	LUT2 #(
		.INIT('h4)
	) name2357 (
		_w1782_,
		_w2888_,
		_w2889_
	);
	LUT2 #(
		.INIT('h4)
	) name2358 (
		_w2887_,
		_w2889_,
		_w2890_
	);
	LUT2 #(
		.INIT('h4)
	) name2359 (
		_w2886_,
		_w2890_,
		_w2891_
	);
	LUT2 #(
		.INIT('h1)
	) name2360 (
		\sa21_reg[1]/P0001 ,
		_w2891_,
		_w2892_
	);
	LUT2 #(
		.INIT('h8)
	) name2361 (
		_w1764_,
		_w1773_,
		_w2893_
	);
	LUT2 #(
		.INIT('h8)
	) name2362 (
		_w1799_,
		_w1844_,
		_w2894_
	);
	LUT2 #(
		.INIT('h4)
	) name2363 (
		\sa21_reg[4]/P0001 ,
		_w2842_,
		_w2895_
	);
	LUT2 #(
		.INIT('h1)
	) name2364 (
		_w1748_,
		_w2893_,
		_w2896_
	);
	LUT2 #(
		.INIT('h1)
	) name2365 (
		_w2894_,
		_w2895_,
		_w2897_
	);
	LUT2 #(
		.INIT('h8)
	) name2366 (
		_w2896_,
		_w2897_,
		_w2898_
	);
	LUT2 #(
		.INIT('h2)
	) name2367 (
		\sa21_reg[1]/P0001 ,
		_w2898_,
		_w2899_
	);
	LUT2 #(
		.INIT('h8)
	) name2368 (
		_w1823_,
		_w2455_,
		_w2900_
	);
	LUT2 #(
		.INIT('h8)
	) name2369 (
		_w1758_,
		_w1799_,
		_w2901_
	);
	LUT2 #(
		.INIT('h4)
	) name2370 (
		\sa21_reg[4]/P0001 ,
		_w2901_,
		_w2902_
	);
	LUT2 #(
		.INIT('h1)
	) name2371 (
		_w1782_,
		_w2902_,
		_w2903_
	);
	LUT2 #(
		.INIT('h2)
	) name2372 (
		\sa21_reg[2]/P0001 ,
		_w2903_,
		_w2904_
	);
	LUT2 #(
		.INIT('h4)
	) name2373 (
		\sa21_reg[4]/P0001 ,
		_w1854_,
		_w2905_
	);
	LUT2 #(
		.INIT('h8)
	) name2374 (
		_w1837_,
		_w2905_,
		_w2906_
	);
	LUT2 #(
		.INIT('h1)
	) name2375 (
		_w2900_,
		_w2906_,
		_w2907_
	);
	LUT2 #(
		.INIT('h4)
	) name2376 (
		_w2904_,
		_w2907_,
		_w2908_
	);
	LUT2 #(
		.INIT('h4)
	) name2377 (
		_w2899_,
		_w2908_,
		_w2909_
	);
	LUT2 #(
		.INIT('h4)
	) name2378 (
		_w2883_,
		_w2909_,
		_w2910_
	);
	LUT2 #(
		.INIT('h4)
	) name2379 (
		_w2892_,
		_w2910_,
		_w2911_
	);
	LUT2 #(
		.INIT('h2)
	) name2380 (
		\sa21_reg[0]/P0001 ,
		_w2911_,
		_w2912_
	);
	LUT2 #(
		.INIT('h1)
	) name2381 (
		_w1780_,
		_w1816_,
		_w2913_
	);
	LUT2 #(
		.INIT('h2)
	) name2382 (
		\sa21_reg[5]/P0001 ,
		_w2913_,
		_w2914_
	);
	LUT2 #(
		.INIT('h1)
	) name2383 (
		_w1834_,
		_w2914_,
		_w2915_
	);
	LUT2 #(
		.INIT('h1)
	) name2384 (
		\sa21_reg[2]/P0001 ,
		_w2915_,
		_w2916_
	);
	LUT2 #(
		.INIT('h8)
	) name2385 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w2917_
	);
	LUT2 #(
		.INIT('h2)
	) name2386 (
		\sa21_reg[3]/P0001 ,
		_w1772_,
		_w2918_
	);
	LUT2 #(
		.INIT('h1)
	) name2387 (
		_w1804_,
		_w2425_,
		_w2919_
	);
	LUT2 #(
		.INIT('h1)
	) name2388 (
		\sa21_reg[3]/P0001 ,
		_w1781_,
		_w2920_
	);
	LUT2 #(
		.INIT('h8)
	) name2389 (
		_w2919_,
		_w2920_,
		_w2921_
	);
	LUT2 #(
		.INIT('h2)
	) name2390 (
		_w2917_,
		_w2918_,
		_w2922_
	);
	LUT2 #(
		.INIT('h4)
	) name2391 (
		_w2921_,
		_w2922_,
		_w2923_
	);
	LUT2 #(
		.INIT('h1)
	) name2392 (
		_w1865_,
		_w2923_,
		_w2924_
	);
	LUT2 #(
		.INIT('h4)
	) name2393 (
		_w2916_,
		_w2924_,
		_w2925_
	);
	LUT2 #(
		.INIT('h1)
	) name2394 (
		\sa21_reg[1]/P0001 ,
		_w2925_,
		_w2926_
	);
	LUT2 #(
		.INIT('h8)
	) name2395 (
		_w1755_,
		_w1822_,
		_w2927_
	);
	LUT2 #(
		.INIT('h8)
	) name2396 (
		_w1747_,
		_w1819_,
		_w2928_
	);
	LUT2 #(
		.INIT('h8)
	) name2397 (
		_w1833_,
		_w1854_,
		_w2929_
	);
	LUT2 #(
		.INIT('h8)
	) name2398 (
		_w1831_,
		_w2436_,
		_w2930_
	);
	LUT2 #(
		.INIT('h1)
	) name2399 (
		_w2869_,
		_w2929_,
		_w2931_
	);
	LUT2 #(
		.INIT('h4)
	) name2400 (
		_w2930_,
		_w2931_,
		_w2932_
	);
	LUT2 #(
		.INIT('h2)
	) name2401 (
		\sa21_reg[1]/P0001 ,
		_w2932_,
		_w2933_
	);
	LUT2 #(
		.INIT('h1)
	) name2402 (
		_w2927_,
		_w2928_,
		_w2934_
	);
	LUT2 #(
		.INIT('h4)
	) name2403 (
		_w1881_,
		_w2934_,
		_w2935_
	);
	LUT2 #(
		.INIT('h4)
	) name2404 (
		_w2933_,
		_w2935_,
		_w2936_
	);
	LUT2 #(
		.INIT('h4)
	) name2405 (
		_w2926_,
		_w2936_,
		_w2937_
	);
	LUT2 #(
		.INIT('h4)
	) name2406 (
		_w2875_,
		_w2937_,
		_w2938_
	);
	LUT2 #(
		.INIT('h4)
	) name2407 (
		_w2912_,
		_w2938_,
		_w2939_
	);
	LUT2 #(
		.INIT('h2)
	) name2408 (
		_w2835_,
		_w2939_,
		_w2940_
	);
	LUT2 #(
		.INIT('h4)
	) name2409 (
		_w2835_,
		_w2939_,
		_w2941_
	);
	LUT2 #(
		.INIT('h1)
	) name2410 (
		_w2940_,
		_w2941_,
		_w2942_
	);
	LUT2 #(
		.INIT('h2)
	) name2411 (
		\u0_w_reg[3][29]/P0001 ,
		_w2077_,
		_w2943_
	);
	LUT2 #(
		.INIT('h4)
	) name2412 (
		\u0_w_reg[3][29]/P0001 ,
		_w2077_,
		_w2944_
	);
	LUT2 #(
		.INIT('h1)
	) name2413 (
		_w2943_,
		_w2944_,
		_w2945_
	);
	LUT2 #(
		.INIT('h8)
	) name2414 (
		_w2942_,
		_w2945_,
		_w2946_
	);
	LUT2 #(
		.INIT('h1)
	) name2415 (
		_w2942_,
		_w2945_,
		_w2947_
	);
	LUT2 #(
		.INIT('h1)
	) name2416 (
		_w2946_,
		_w2947_,
		_w2948_
	);
	LUT2 #(
		.INIT('h1)
	) name2417 (
		_w2739_,
		_w2948_,
		_w2949_
	);
	LUT2 #(
		.INIT('h8)
	) name2418 (
		_w2739_,
		_w2948_,
		_w2950_
	);
	LUT2 #(
		.INIT('h1)
	) name2419 (
		\ld_r_reg/P0001 ,
		_w2949_,
		_w2951_
	);
	LUT2 #(
		.INIT('h4)
	) name2420 (
		_w2950_,
		_w2951_,
		_w2952_
	);
	LUT2 #(
		.INIT('h1)
	) name2421 (
		\text_in_r_reg[29]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		_w2953_
	);
	LUT2 #(
		.INIT('h8)
	) name2422 (
		\text_in_r_reg[29]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		_w2954_
	);
	LUT2 #(
		.INIT('h2)
	) name2423 (
		\ld_r_reg/P0001 ,
		_w2953_,
		_w2955_
	);
	LUT2 #(
		.INIT('h4)
	) name2424 (
		_w2954_,
		_w2955_,
		_w2956_
	);
	LUT2 #(
		.INIT('h1)
	) name2425 (
		_w2952_,
		_w2956_,
		_w2957_
	);
	LUT2 #(
		.INIT('h2)
	) name2426 (
		_w1738_,
		_w1908_,
		_w2958_
	);
	LUT2 #(
		.INIT('h4)
	) name2427 (
		_w1738_,
		_w1908_,
		_w2959_
	);
	LUT2 #(
		.INIT('h1)
	) name2428 (
		_w2958_,
		_w2959_,
		_w2960_
	);
	LUT2 #(
		.INIT('h1)
	) name2429 (
		_w1479_,
		_w2835_,
		_w2961_
	);
	LUT2 #(
		.INIT('h8)
	) name2430 (
		_w1479_,
		_w2835_,
		_w2962_
	);
	LUT2 #(
		.INIT('h1)
	) name2431 (
		_w2961_,
		_w2962_,
		_w2963_
	);
	LUT2 #(
		.INIT('h2)
	) name2432 (
		\u0_w_reg[3][30]/P0001 ,
		_w2416_,
		_w2964_
	);
	LUT2 #(
		.INIT('h4)
	) name2433 (
		\u0_w_reg[3][30]/P0001 ,
		_w2416_,
		_w2965_
	);
	LUT2 #(
		.INIT('h1)
	) name2434 (
		_w2964_,
		_w2965_,
		_w2966_
	);
	LUT2 #(
		.INIT('h8)
	) name2435 (
		_w2963_,
		_w2966_,
		_w2967_
	);
	LUT2 #(
		.INIT('h1)
	) name2436 (
		_w2963_,
		_w2966_,
		_w2968_
	);
	LUT2 #(
		.INIT('h1)
	) name2437 (
		_w2967_,
		_w2968_,
		_w2969_
	);
	LUT2 #(
		.INIT('h1)
	) name2438 (
		_w2960_,
		_w2969_,
		_w2970_
	);
	LUT2 #(
		.INIT('h8)
	) name2439 (
		_w2960_,
		_w2969_,
		_w2971_
	);
	LUT2 #(
		.INIT('h1)
	) name2440 (
		\ld_r_reg/P0001 ,
		_w2970_,
		_w2972_
	);
	LUT2 #(
		.INIT('h4)
	) name2441 (
		_w2971_,
		_w2972_,
		_w2973_
	);
	LUT2 #(
		.INIT('h2)
	) name2442 (
		\text_in_r_reg[30]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w2974_
	);
	LUT2 #(
		.INIT('h4)
	) name2443 (
		\text_in_r_reg[30]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w2975_
	);
	LUT2 #(
		.INIT('h2)
	) name2444 (
		\ld_r_reg/P0001 ,
		_w2974_,
		_w2976_
	);
	LUT2 #(
		.INIT('h4)
	) name2445 (
		_w2975_,
		_w2976_,
		_w2977_
	);
	LUT2 #(
		.INIT('h1)
	) name2446 (
		_w2973_,
		_w2977_,
		_w2978_
	);
	LUT2 #(
		.INIT('h8)
	) name2447 (
		\sa21_reg[5]/P0001 ,
		_w2446_,
		_w2979_
	);
	LUT2 #(
		.INIT('h8)
	) name2448 (
		\sa21_reg[3]/P0001 ,
		_w2862_,
		_w2980_
	);
	LUT2 #(
		.INIT('h1)
	) name2449 (
		_w2979_,
		_w2980_,
		_w2981_
	);
	LUT2 #(
		.INIT('h1)
	) name2450 (
		\sa21_reg[1]/P0001 ,
		_w2981_,
		_w2982_
	);
	LUT2 #(
		.INIT('h1)
	) name2451 (
		_w1853_,
		_w2477_,
		_w2983_
	);
	LUT2 #(
		.INIT('h1)
	) name2452 (
		\sa21_reg[1]/P0001 ,
		_w2983_,
		_w2984_
	);
	LUT2 #(
		.INIT('h8)
	) name2453 (
		_w1802_,
		_w2477_,
		_w2985_
	);
	LUT2 #(
		.INIT('h1)
	) name2454 (
		_w2984_,
		_w2985_,
		_w2986_
	);
	LUT2 #(
		.INIT('h2)
	) name2455 (
		\sa21_reg[2]/P0001 ,
		_w2986_,
		_w2987_
	);
	LUT2 #(
		.INIT('h8)
	) name2456 (
		\sa21_reg[2]/P0001 ,
		_w1759_,
		_w2988_
	);
	LUT2 #(
		.INIT('h1)
	) name2457 (
		_w1880_,
		_w2900_,
		_w2989_
	);
	LUT2 #(
		.INIT('h4)
	) name2458 (
		_w2988_,
		_w2989_,
		_w2990_
	);
	LUT2 #(
		.INIT('h1)
	) name2459 (
		\sa21_reg[3]/P0001 ,
		_w2990_,
		_w2991_
	);
	LUT2 #(
		.INIT('h2)
	) name2460 (
		_w1764_,
		_w1866_,
		_w2992_
	);
	LUT2 #(
		.INIT('h8)
	) name2461 (
		_w1793_,
		_w1832_,
		_w2993_
	);
	LUT2 #(
		.INIT('h1)
	) name2462 (
		_w2992_,
		_w2993_,
		_w2994_
	);
	LUT2 #(
		.INIT('h1)
	) name2463 (
		\sa21_reg[2]/P0001 ,
		_w2994_,
		_w2995_
	);
	LUT2 #(
		.INIT('h8)
	) name2464 (
		_w1831_,
		_w2490_,
		_w2996_
	);
	LUT2 #(
		.INIT('h8)
	) name2465 (
		\sa21_reg[6]/NET0131 ,
		_w1819_,
		_w2997_
	);
	LUT2 #(
		.INIT('h1)
	) name2466 (
		_w1780_,
		_w2996_,
		_w2998_
	);
	LUT2 #(
		.INIT('h4)
	) name2467 (
		_w2997_,
		_w2998_,
		_w2999_
	);
	LUT2 #(
		.INIT('h4)
	) name2468 (
		_w2995_,
		_w2999_,
		_w3000_
	);
	LUT2 #(
		.INIT('h2)
	) name2469 (
		\sa21_reg[1]/P0001 ,
		_w3000_,
		_w3001_
	);
	LUT2 #(
		.INIT('h1)
	) name2470 (
		_w2982_,
		_w2987_,
		_w3002_
	);
	LUT2 #(
		.INIT('h4)
	) name2471 (
		_w2991_,
		_w3002_,
		_w3003_
	);
	LUT2 #(
		.INIT('h4)
	) name2472 (
		_w3001_,
		_w3003_,
		_w3004_
	);
	LUT2 #(
		.INIT('h1)
	) name2473 (
		\sa21_reg[0]/P0001 ,
		_w3004_,
		_w3005_
	);
	LUT2 #(
		.INIT('h8)
	) name2474 (
		_w1762_,
		_w1831_,
		_w3006_
	);
	LUT2 #(
		.INIT('h1)
	) name2475 (
		_w1842_,
		_w1883_,
		_w3007_
	);
	LUT2 #(
		.INIT('h4)
	) name2476 (
		_w2853_,
		_w3007_,
		_w3008_
	);
	LUT2 #(
		.INIT('h1)
	) name2477 (
		\sa21_reg[2]/P0001 ,
		_w3008_,
		_w3009_
	);
	LUT2 #(
		.INIT('h4)
	) name2478 (
		\sa21_reg[5]/P0001 ,
		_w2895_,
		_w3010_
	);
	LUT2 #(
		.INIT('h1)
	) name2479 (
		_w1820_,
		_w2465_,
		_w3011_
	);
	LUT2 #(
		.INIT('h4)
	) name2480 (
		_w3006_,
		_w3011_,
		_w3012_
	);
	LUT2 #(
		.INIT('h4)
	) name2481 (
		_w3010_,
		_w3012_,
		_w3013_
	);
	LUT2 #(
		.INIT('h4)
	) name2482 (
		_w3009_,
		_w3013_,
		_w3014_
	);
	LUT2 #(
		.INIT('h2)
	) name2483 (
		\sa21_reg[1]/P0001 ,
		_w3014_,
		_w3015_
	);
	LUT2 #(
		.INIT('h8)
	) name2484 (
		_w1853_,
		_w1894_,
		_w3016_
	);
	LUT2 #(
		.INIT('h8)
	) name2485 (
		_w1877_,
		_w2417_,
		_w3017_
	);
	LUT2 #(
		.INIT('h1)
	) name2486 (
		_w1775_,
		_w2426_,
		_w3018_
	);
	LUT2 #(
		.INIT('h1)
	) name2487 (
		\sa21_reg[2]/P0001 ,
		_w3018_,
		_w3019_
	);
	LUT2 #(
		.INIT('h8)
	) name2488 (
		_w1841_,
		_w1867_,
		_w3020_
	);
	LUT2 #(
		.INIT('h8)
	) name2489 (
		_w1763_,
		_w2856_,
		_w3021_
	);
	LUT2 #(
		.INIT('h1)
	) name2490 (
		_w2894_,
		_w3021_,
		_w3022_
	);
	LUT2 #(
		.INIT('h4)
	) name2491 (
		_w3020_,
		_w3022_,
		_w3023_
	);
	LUT2 #(
		.INIT('h4)
	) name2492 (
		_w3019_,
		_w3023_,
		_w3024_
	);
	LUT2 #(
		.INIT('h2)
	) name2493 (
		\sa21_reg[1]/P0001 ,
		_w3024_,
		_w3025_
	);
	LUT2 #(
		.INIT('h1)
	) name2494 (
		\sa21_reg[3]/P0001 ,
		_w2479_,
		_w3026_
	);
	LUT2 #(
		.INIT('h2)
	) name2495 (
		_w1749_,
		_w3026_,
		_w3027_
	);
	LUT2 #(
		.INIT('h4)
	) name2496 (
		\sa21_reg[2]/P0001 ,
		_w2884_,
		_w3028_
	);
	LUT2 #(
		.INIT('h8)
	) name2497 (
		_w1822_,
		_w1866_,
		_w3029_
	);
	LUT2 #(
		.INIT('h8)
	) name2498 (
		_w1764_,
		_w2917_,
		_w3030_
	);
	LUT2 #(
		.INIT('h1)
	) name2499 (
		_w3027_,
		_w3029_,
		_w3031_
	);
	LUT2 #(
		.INIT('h4)
	) name2500 (
		_w3030_,
		_w3031_,
		_w3032_
	);
	LUT2 #(
		.INIT('h4)
	) name2501 (
		_w3028_,
		_w3032_,
		_w3033_
	);
	LUT2 #(
		.INIT('h1)
	) name2502 (
		\sa21_reg[1]/P0001 ,
		_w3033_,
		_w3034_
	);
	LUT2 #(
		.INIT('h1)
	) name2503 (
		_w1746_,
		_w1781_,
		_w3035_
	);
	LUT2 #(
		.INIT('h1)
	) name2504 (
		\sa21_reg[4]/P0001 ,
		_w3035_,
		_w3036_
	);
	LUT2 #(
		.INIT('h2)
	) name2505 (
		\sa21_reg[2]/P0001 ,
		_w1788_,
		_w3037_
	);
	LUT2 #(
		.INIT('h4)
	) name2506 (
		_w2864_,
		_w3037_,
		_w3038_
	);
	LUT2 #(
		.INIT('h4)
	) name2507 (
		_w3036_,
		_w3038_,
		_w3039_
	);
	LUT2 #(
		.INIT('h8)
	) name2508 (
		_w1787_,
		_w1822_,
		_w3040_
	);
	LUT2 #(
		.INIT('h1)
	) name2509 (
		\sa21_reg[2]/P0001 ,
		_w2876_,
		_w3041_
	);
	LUT2 #(
		.INIT('h4)
	) name2510 (
		_w3040_,
		_w3041_,
		_w3042_
	);
	LUT2 #(
		.INIT('h4)
	) name2511 (
		_w1883_,
		_w3042_,
		_w3043_
	);
	LUT2 #(
		.INIT('h1)
	) name2512 (
		_w3039_,
		_w3043_,
		_w3044_
	);
	LUT2 #(
		.INIT('h1)
	) name2513 (
		_w3025_,
		_w3044_,
		_w3045_
	);
	LUT2 #(
		.INIT('h4)
	) name2514 (
		_w3034_,
		_w3045_,
		_w3046_
	);
	LUT2 #(
		.INIT('h2)
	) name2515 (
		\sa21_reg[0]/P0001 ,
		_w3046_,
		_w3047_
	);
	LUT2 #(
		.INIT('h4)
	) name2516 (
		\sa21_reg[7]/P0001 ,
		_w1815_,
		_w3048_
	);
	LUT2 #(
		.INIT('h8)
	) name2517 (
		_w1772_,
		_w3048_,
		_w3049_
	);
	LUT2 #(
		.INIT('h8)
	) name2518 (
		_w1822_,
		_w1867_,
		_w3050_
	);
	LUT2 #(
		.INIT('h1)
	) name2519 (
		_w2516_,
		_w2838_,
		_w3051_
	);
	LUT2 #(
		.INIT('h4)
	) name2520 (
		_w3050_,
		_w3051_,
		_w3052_
	);
	LUT2 #(
		.INIT('h1)
	) name2521 (
		\sa21_reg[2]/P0001 ,
		_w3052_,
		_w3053_
	);
	LUT2 #(
		.INIT('h2)
	) name2522 (
		\sa21_reg[5]/P0001 ,
		_w2438_,
		_w3054_
	);
	LUT2 #(
		.INIT('h8)
	) name2523 (
		_w1757_,
		_w1833_,
		_w3055_
	);
	LUT2 #(
		.INIT('h8)
	) name2524 (
		_w1802_,
		_w2425_,
		_w3056_
	);
	LUT2 #(
		.INIT('h1)
	) name2525 (
		_w2447_,
		_w3055_,
		_w3057_
	);
	LUT2 #(
		.INIT('h4)
	) name2526 (
		_w3056_,
		_w3057_,
		_w3058_
	);
	LUT2 #(
		.INIT('h4)
	) name2527 (
		_w3054_,
		_w3058_,
		_w3059_
	);
	LUT2 #(
		.INIT('h2)
	) name2528 (
		\sa21_reg[2]/P0001 ,
		_w3059_,
		_w3060_
	);
	LUT2 #(
		.INIT('h1)
	) name2529 (
		_w1855_,
		_w3049_,
		_w3061_
	);
	LUT2 #(
		.INIT('h4)
	) name2530 (
		_w3053_,
		_w3061_,
		_w3062_
	);
	LUT2 #(
		.INIT('h4)
	) name2531 (
		_w3060_,
		_w3062_,
		_w3063_
	);
	LUT2 #(
		.INIT('h1)
	) name2532 (
		\sa21_reg[1]/P0001 ,
		_w3063_,
		_w3064_
	);
	LUT2 #(
		.INIT('h1)
	) name2533 (
		_w3016_,
		_w3017_,
		_w3065_
	);
	LUT2 #(
		.INIT('h4)
	) name2534 (
		_w3015_,
		_w3065_,
		_w3066_
	);
	LUT2 #(
		.INIT('h4)
	) name2535 (
		_w3064_,
		_w3066_,
		_w3067_
	);
	LUT2 #(
		.INIT('h4)
	) name2536 (
		_w3005_,
		_w3067_,
		_w3068_
	);
	LUT2 #(
		.INIT('h4)
	) name2537 (
		_w3047_,
		_w3068_,
		_w3069_
	);
	LUT2 #(
		.INIT('h2)
	) name2538 (
		_w2647_,
		_w3069_,
		_w3070_
	);
	LUT2 #(
		.INIT('h4)
	) name2539 (
		_w2647_,
		_w3069_,
		_w3071_
	);
	LUT2 #(
		.INIT('h1)
	) name2540 (
		_w3070_,
		_w3071_,
		_w3072_
	);
	LUT2 #(
		.INIT('h1)
	) name2541 (
		_w1479_,
		_w3072_,
		_w3073_
	);
	LUT2 #(
		.INIT('h8)
	) name2542 (
		_w1479_,
		_w3072_,
		_w3074_
	);
	LUT2 #(
		.INIT('h1)
	) name2543 (
		_w3073_,
		_w3074_,
		_w3075_
	);
	LUT2 #(
		.INIT('h2)
	) name2544 (
		\u0_w_reg[3][21]/P0001 ,
		_w2077_,
		_w3076_
	);
	LUT2 #(
		.INIT('h4)
	) name2545 (
		\u0_w_reg[3][21]/P0001 ,
		_w2077_,
		_w3077_
	);
	LUT2 #(
		.INIT('h1)
	) name2546 (
		_w3076_,
		_w3077_,
		_w3078_
	);
	LUT2 #(
		.INIT('h8)
	) name2547 (
		_w2939_,
		_w3078_,
		_w3079_
	);
	LUT2 #(
		.INIT('h1)
	) name2548 (
		_w2939_,
		_w3078_,
		_w3080_
	);
	LUT2 #(
		.INIT('h1)
	) name2549 (
		_w3079_,
		_w3080_,
		_w3081_
	);
	LUT2 #(
		.INIT('h1)
	) name2550 (
		_w3075_,
		_w3081_,
		_w3082_
	);
	LUT2 #(
		.INIT('h8)
	) name2551 (
		_w3075_,
		_w3081_,
		_w3083_
	);
	LUT2 #(
		.INIT('h1)
	) name2552 (
		\ld_r_reg/P0001 ,
		_w3082_,
		_w3084_
	);
	LUT2 #(
		.INIT('h4)
	) name2553 (
		_w3083_,
		_w3084_,
		_w3085_
	);
	LUT2 #(
		.INIT('h2)
	) name2554 (
		\text_in_r_reg[21]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		_w3086_
	);
	LUT2 #(
		.INIT('h4)
	) name2555 (
		\text_in_r_reg[21]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		_w3087_
	);
	LUT2 #(
		.INIT('h2)
	) name2556 (
		\ld_r_reg/P0001 ,
		_w3086_,
		_w3088_
	);
	LUT2 #(
		.INIT('h4)
	) name2557 (
		_w3087_,
		_w3088_,
		_w3089_
	);
	LUT2 #(
		.INIT('h1)
	) name2558 (
		_w3085_,
		_w3089_,
		_w3090_
	);
	LUT2 #(
		.INIT('h1)
	) name2559 (
		_w1581_,
		_w2942_,
		_w3091_
	);
	LUT2 #(
		.INIT('h8)
	) name2560 (
		_w1581_,
		_w2942_,
		_w3092_
	);
	LUT2 #(
		.INIT('h1)
	) name2561 (
		_w3091_,
		_w3092_,
		_w3093_
	);
	LUT2 #(
		.INIT('h2)
	) name2562 (
		\u0_w_reg[3][22]/P0001 ,
		_w2416_,
		_w3094_
	);
	LUT2 #(
		.INIT('h4)
	) name2563 (
		\u0_w_reg[3][22]/P0001 ,
		_w2416_,
		_w3095_
	);
	LUT2 #(
		.INIT('h1)
	) name2564 (
		_w3094_,
		_w3095_,
		_w3096_
	);
	LUT2 #(
		.INIT('h8)
	) name2565 (
		_w1908_,
		_w3096_,
		_w3097_
	);
	LUT2 #(
		.INIT('h1)
	) name2566 (
		_w1908_,
		_w3096_,
		_w3098_
	);
	LUT2 #(
		.INIT('h1)
	) name2567 (
		_w3097_,
		_w3098_,
		_w3099_
	);
	LUT2 #(
		.INIT('h1)
	) name2568 (
		_w3093_,
		_w3099_,
		_w3100_
	);
	LUT2 #(
		.INIT('h8)
	) name2569 (
		_w3093_,
		_w3099_,
		_w3101_
	);
	LUT2 #(
		.INIT('h1)
	) name2570 (
		\ld_r_reg/P0001 ,
		_w3100_,
		_w3102_
	);
	LUT2 #(
		.INIT('h4)
	) name2571 (
		_w3101_,
		_w3102_,
		_w3103_
	);
	LUT2 #(
		.INIT('h2)
	) name2572 (
		\text_in_r_reg[22]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w3104_
	);
	LUT2 #(
		.INIT('h4)
	) name2573 (
		\text_in_r_reg[22]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w3105_
	);
	LUT2 #(
		.INIT('h2)
	) name2574 (
		\ld_r_reg/P0001 ,
		_w3104_,
		_w3106_
	);
	LUT2 #(
		.INIT('h4)
	) name2575 (
		_w3105_,
		_w3106_,
		_w3107_
	);
	LUT2 #(
		.INIT('h1)
	) name2576 (
		_w3103_,
		_w3107_,
		_w3108_
	);
	LUT2 #(
		.INIT('h1)
	) name2577 (
		_w2963_,
		_w3069_,
		_w3109_
	);
	LUT2 #(
		.INIT('h8)
	) name2578 (
		_w2963_,
		_w3069_,
		_w3110_
	);
	LUT2 #(
		.INIT('h1)
	) name2579 (
		_w3109_,
		_w3110_,
		_w3111_
	);
	LUT2 #(
		.INIT('h1)
	) name2580 (
		_w2363_,
		_w2375_,
		_w3112_
	);
	LUT2 #(
		.INIT('h4)
	) name2581 (
		_w2013_,
		_w3112_,
		_w3113_
	);
	LUT2 #(
		.INIT('h1)
	) name2582 (
		\sa32_reg[2]/P0001 ,
		_w3113_,
		_w3114_
	);
	LUT2 #(
		.INIT('h8)
	) name2583 (
		_w2315_,
		_w2397_,
		_w3115_
	);
	LUT2 #(
		.INIT('h4)
	) name2584 (
		\sa32_reg[5]/P0001 ,
		_w1933_,
		_w3116_
	);
	LUT2 #(
		.INIT('h8)
	) name2585 (
		\sa32_reg[3]/P0001 ,
		_w1963_,
		_w3117_
	);
	LUT2 #(
		.INIT('h1)
	) name2586 (
		_w2061_,
		_w3115_,
		_w3118_
	);
	LUT2 #(
		.INIT('h4)
	) name2587 (
		_w3117_,
		_w3118_,
		_w3119_
	);
	LUT2 #(
		.INIT('h4)
	) name2588 (
		_w3116_,
		_w3119_,
		_w3120_
	);
	LUT2 #(
		.INIT('h4)
	) name2589 (
		_w3114_,
		_w3120_,
		_w3121_
	);
	LUT2 #(
		.INIT('h2)
	) name2590 (
		\sa32_reg[1]/P0001 ,
		_w3121_,
		_w3122_
	);
	LUT2 #(
		.INIT('h8)
	) name2591 (
		_w2030_,
		_w2366_,
		_w3123_
	);
	LUT2 #(
		.INIT('h8)
	) name2592 (
		\sa32_reg[4]/P0001 ,
		_w1909_,
		_w3124_
	);
	LUT2 #(
		.INIT('h8)
	) name2593 (
		_w2059_,
		_w3124_,
		_w3125_
	);
	LUT2 #(
		.INIT('h8)
	) name2594 (
		_w1939_,
		_w2362_,
		_w3126_
	);
	LUT2 #(
		.INIT('h1)
	) name2595 (
		_w1919_,
		_w1951_,
		_w3127_
	);
	LUT2 #(
		.INIT('h8)
	) name2596 (
		_w2041_,
		_w3127_,
		_w3128_
	);
	LUT2 #(
		.INIT('h8)
	) name2597 (
		_w1939_,
		_w1951_,
		_w3129_
	);
	LUT2 #(
		.INIT('h2)
	) name2598 (
		\sa32_reg[2]/P0001 ,
		_w3129_,
		_w3130_
	);
	LUT2 #(
		.INIT('h4)
	) name2599 (
		_w1911_,
		_w3130_,
		_w3131_
	);
	LUT2 #(
		.INIT('h1)
	) name2600 (
		_w2332_,
		_w3128_,
		_w3132_
	);
	LUT2 #(
		.INIT('h8)
	) name2601 (
		_w3131_,
		_w3132_,
		_w3133_
	);
	LUT2 #(
		.INIT('h8)
	) name2602 (
		_w1951_,
		_w2011_,
		_w3134_
	);
	LUT2 #(
		.INIT('h4)
	) name2603 (
		_w1948_,
		_w1965_,
		_w3135_
	);
	LUT2 #(
		.INIT('h1)
	) name2604 (
		\sa32_reg[2]/P0001 ,
		_w3134_,
		_w3136_
	);
	LUT2 #(
		.INIT('h4)
	) name2605 (
		_w3135_,
		_w3136_,
		_w3137_
	);
	LUT2 #(
		.INIT('h1)
	) name2606 (
		_w3133_,
		_w3137_,
		_w3138_
	);
	LUT2 #(
		.INIT('h1)
	) name2607 (
		_w2052_,
		_w3126_,
		_w3139_
	);
	LUT2 #(
		.INIT('h4)
	) name2608 (
		_w3138_,
		_w3139_,
		_w3140_
	);
	LUT2 #(
		.INIT('h1)
	) name2609 (
		\sa32_reg[1]/P0001 ,
		_w3140_,
		_w3141_
	);
	LUT2 #(
		.INIT('h4)
	) name2610 (
		\sa32_reg[3]/P0001 ,
		_w1964_,
		_w3142_
	);
	LUT2 #(
		.INIT('h8)
	) name2611 (
		\sa32_reg[5]/P0001 ,
		_w1923_,
		_w3143_
	);
	LUT2 #(
		.INIT('h4)
	) name2612 (
		_w1951_,
		_w3143_,
		_w3144_
	);
	LUT2 #(
		.INIT('h4)
	) name2613 (
		\sa32_reg[5]/P0001 ,
		_w2049_,
		_w3145_
	);
	LUT2 #(
		.INIT('h4)
	) name2614 (
		\sa32_reg[6]/NET0131 ,
		_w3145_,
		_w3146_
	);
	LUT2 #(
		.INIT('h1)
	) name2615 (
		_w3144_,
		_w3146_,
		_w3147_
	);
	LUT2 #(
		.INIT('h1)
	) name2616 (
		\sa32_reg[2]/P0001 ,
		_w3147_,
		_w3148_
	);
	LUT2 #(
		.INIT('h8)
	) name2617 (
		\sa32_reg[4]/P0001 ,
		_w2387_,
		_w3149_
	);
	LUT2 #(
		.INIT('h8)
	) name2618 (
		_w2397_,
		_w3149_,
		_w3150_
	);
	LUT2 #(
		.INIT('h1)
	) name2619 (
		_w2068_,
		_w2327_,
		_w3151_
	);
	LUT2 #(
		.INIT('h4)
	) name2620 (
		_w3150_,
		_w3151_,
		_w3152_
	);
	LUT2 #(
		.INIT('h4)
	) name2621 (
		_w3148_,
		_w3152_,
		_w3153_
	);
	LUT2 #(
		.INIT('h2)
	) name2622 (
		\sa32_reg[1]/P0001 ,
		_w3153_,
		_w3154_
	);
	LUT2 #(
		.INIT('h8)
	) name2623 (
		_w1909_,
		_w2313_,
		_w3155_
	);
	LUT2 #(
		.INIT('h1)
	) name2624 (
		_w2004_,
		_w3155_,
		_w3156_
	);
	LUT2 #(
		.INIT('h1)
	) name2625 (
		\sa32_reg[7]/P0001 ,
		_w3156_,
		_w3157_
	);
	LUT2 #(
		.INIT('h1)
	) name2626 (
		_w1937_,
		_w3124_,
		_w3158_
	);
	LUT2 #(
		.INIT('h2)
	) name2627 (
		\sa32_reg[2]/P0001 ,
		_w3158_,
		_w3159_
	);
	LUT2 #(
		.INIT('h1)
	) name2628 (
		_w3157_,
		_w3159_,
		_w3160_
	);
	LUT2 #(
		.INIT('h1)
	) name2629 (
		\sa32_reg[1]/P0001 ,
		_w3160_,
		_w3161_
	);
	LUT2 #(
		.INIT('h4)
	) name2630 (
		\sa32_reg[5]/P0001 ,
		_w1914_,
		_w3162_
	);
	LUT2 #(
		.INIT('h1)
	) name2631 (
		_w2316_,
		_w3162_,
		_w3163_
	);
	LUT2 #(
		.INIT('h2)
	) name2632 (
		\sa32_reg[2]/P0001 ,
		_w3163_,
		_w3164_
	);
	LUT2 #(
		.INIT('h1)
	) name2633 (
		_w3126_,
		_w3142_,
		_w3165_
	);
	LUT2 #(
		.INIT('h4)
	) name2634 (
		_w3164_,
		_w3165_,
		_w3166_
	);
	LUT2 #(
		.INIT('h4)
	) name2635 (
		_w3161_,
		_w3166_,
		_w3167_
	);
	LUT2 #(
		.INIT('h4)
	) name2636 (
		_w3154_,
		_w3167_,
		_w3168_
	);
	LUT2 #(
		.INIT('h1)
	) name2637 (
		\sa32_reg[0]/P0002 ,
		_w3168_,
		_w3169_
	);
	LUT2 #(
		.INIT('h1)
	) name2638 (
		\sa32_reg[3]/P0001 ,
		_w2030_,
		_w3170_
	);
	LUT2 #(
		.INIT('h2)
	) name2639 (
		_w1920_,
		_w3170_,
		_w3171_
	);
	LUT2 #(
		.INIT('h8)
	) name2640 (
		_w1947_,
		_w2049_,
		_w3172_
	);
	LUT2 #(
		.INIT('h1)
	) name2641 (
		\sa32_reg[1]/P0001 ,
		_w3172_,
		_w3173_
	);
	LUT2 #(
		.INIT('h8)
	) name2642 (
		\sa32_reg[2]/P0001 ,
		_w2024_,
		_w3174_
	);
	LUT2 #(
		.INIT('h4)
	) name2643 (
		\sa32_reg[2]/P0001 ,
		_w1914_,
		_w3175_
	);
	LUT2 #(
		.INIT('h4)
	) name2644 (
		_w3171_,
		_w3173_,
		_w3176_
	);
	LUT2 #(
		.INIT('h1)
	) name2645 (
		_w3174_,
		_w3175_,
		_w3177_
	);
	LUT2 #(
		.INIT('h8)
	) name2646 (
		_w3176_,
		_w3177_,
		_w3178_
	);
	LUT2 #(
		.INIT('h2)
	) name2647 (
		\sa32_reg[1]/P0001 ,
		_w2063_,
		_w3179_
	);
	LUT2 #(
		.INIT('h4)
	) name2648 (
		\sa32_reg[4]/P0001 ,
		_w1981_,
		_w3180_
	);
	LUT2 #(
		.INIT('h8)
	) name2649 (
		_w1953_,
		_w1990_,
		_w3181_
	);
	LUT2 #(
		.INIT('h1)
	) name2650 (
		_w3180_,
		_w3181_,
		_w3182_
	);
	LUT2 #(
		.INIT('h1)
	) name2651 (
		\sa32_reg[2]/P0001 ,
		_w3182_,
		_w3183_
	);
	LUT2 #(
		.INIT('h8)
	) name2652 (
		_w1923_,
		_w2348_,
		_w3184_
	);
	LUT2 #(
		.INIT('h1)
	) name2653 (
		_w1938_,
		_w3184_,
		_w3185_
	);
	LUT2 #(
		.INIT('h8)
	) name2654 (
		_w3179_,
		_w3185_,
		_w3186_
	);
	LUT2 #(
		.INIT('h4)
	) name2655 (
		_w3183_,
		_w3186_,
		_w3187_
	);
	LUT2 #(
		.INIT('h1)
	) name2656 (
		_w3178_,
		_w3187_,
		_w3188_
	);
	LUT2 #(
		.INIT('h4)
	) name2657 (
		\sa32_reg[7]/P0001 ,
		_w1919_,
		_w3189_
	);
	LUT2 #(
		.INIT('h2)
	) name2658 (
		\sa32_reg[2]/P0001 ,
		_w1925_,
		_w3190_
	);
	LUT2 #(
		.INIT('h1)
	) name2659 (
		_w2004_,
		_w2346_,
		_w3191_
	);
	LUT2 #(
		.INIT('h4)
	) name2660 (
		_w3189_,
		_w3191_,
		_w3192_
	);
	LUT2 #(
		.INIT('h8)
	) name2661 (
		_w3190_,
		_w3192_,
		_w3193_
	);
	LUT2 #(
		.INIT('h8)
	) name2662 (
		_w1924_,
		_w1987_,
		_w3194_
	);
	LUT2 #(
		.INIT('h1)
	) name2663 (
		\sa32_reg[2]/P0001 ,
		_w1949_,
		_w3195_
	);
	LUT2 #(
		.INIT('h4)
	) name2664 (
		_w3194_,
		_w3195_,
		_w3196_
	);
	LUT2 #(
		.INIT('h4)
	) name2665 (
		_w2363_,
		_w3196_,
		_w3197_
	);
	LUT2 #(
		.INIT('h1)
	) name2666 (
		_w3193_,
		_w3197_,
		_w3198_
	);
	LUT2 #(
		.INIT('h1)
	) name2667 (
		_w3188_,
		_w3198_,
		_w3199_
	);
	LUT2 #(
		.INIT('h2)
	) name2668 (
		\sa32_reg[0]/P0002 ,
		_w3199_,
		_w3200_
	);
	LUT2 #(
		.INIT('h1)
	) name2669 (
		_w3123_,
		_w3125_,
		_w3201_
	);
	LUT2 #(
		.INIT('h4)
	) name2670 (
		_w3122_,
		_w3201_,
		_w3202_
	);
	LUT2 #(
		.INIT('h4)
	) name2671 (
		_w3141_,
		_w3202_,
		_w3203_
	);
	LUT2 #(
		.INIT('h1)
	) name2672 (
		_w3169_,
		_w3200_,
		_w3204_
	);
	LUT2 #(
		.INIT('h8)
	) name2673 (
		_w3203_,
		_w3204_,
		_w3205_
	);
	LUT2 #(
		.INIT('h2)
	) name2674 (
		\u0_w_reg[3][13]/P0001 ,
		_w3205_,
		_w3206_
	);
	LUT2 #(
		.INIT('h4)
	) name2675 (
		\u0_w_reg[3][13]/P0001 ,
		_w3205_,
		_w3207_
	);
	LUT2 #(
		.INIT('h1)
	) name2676 (
		_w3206_,
		_w3207_,
		_w3208_
	);
	LUT2 #(
		.INIT('h8)
	) name2677 (
		_w2077_,
		_w3208_,
		_w3209_
	);
	LUT2 #(
		.INIT('h1)
	) name2678 (
		_w2077_,
		_w3208_,
		_w3210_
	);
	LUT2 #(
		.INIT('h1)
	) name2679 (
		_w3209_,
		_w3210_,
		_w3211_
	);
	LUT2 #(
		.INIT('h1)
	) name2680 (
		_w3111_,
		_w3211_,
		_w3212_
	);
	LUT2 #(
		.INIT('h8)
	) name2681 (
		_w3111_,
		_w3211_,
		_w3213_
	);
	LUT2 #(
		.INIT('h1)
	) name2682 (
		\ld_r_reg/P0001 ,
		_w3212_,
		_w3214_
	);
	LUT2 #(
		.INIT('h4)
	) name2683 (
		_w3213_,
		_w3214_,
		_w3215_
	);
	LUT2 #(
		.INIT('h1)
	) name2684 (
		\text_in_r_reg[13]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		_w3216_
	);
	LUT2 #(
		.INIT('h8)
	) name2685 (
		\text_in_r_reg[13]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		_w3217_
	);
	LUT2 #(
		.INIT('h2)
	) name2686 (
		\ld_r_reg/P0001 ,
		_w3216_,
		_w3218_
	);
	LUT2 #(
		.INIT('h4)
	) name2687 (
		_w3217_,
		_w3218_,
		_w3219_
	);
	LUT2 #(
		.INIT('h1)
	) name2688 (
		_w3215_,
		_w3219_,
		_w3220_
	);
	LUT2 #(
		.INIT('h1)
	) name2689 (
		_w1741_,
		_w2939_,
		_w3221_
	);
	LUT2 #(
		.INIT('h8)
	) name2690 (
		_w1741_,
		_w2939_,
		_w3222_
	);
	LUT2 #(
		.INIT('h1)
	) name2691 (
		_w3221_,
		_w3222_,
		_w3223_
	);
	LUT2 #(
		.INIT('h2)
	) name2692 (
		\u0_w_reg[3][14]/P0001 ,
		_w2416_,
		_w3224_
	);
	LUT2 #(
		.INIT('h4)
	) name2693 (
		\u0_w_reg[3][14]/P0001 ,
		_w2416_,
		_w3225_
	);
	LUT2 #(
		.INIT('h1)
	) name2694 (
		_w3224_,
		_w3225_,
		_w3226_
	);
	LUT2 #(
		.INIT('h8)
	) name2695 (
		_w2077_,
		_w3226_,
		_w3227_
	);
	LUT2 #(
		.INIT('h1)
	) name2696 (
		_w2077_,
		_w3226_,
		_w3228_
	);
	LUT2 #(
		.INIT('h1)
	) name2697 (
		_w3227_,
		_w3228_,
		_w3229_
	);
	LUT2 #(
		.INIT('h1)
	) name2698 (
		_w3223_,
		_w3229_,
		_w3230_
	);
	LUT2 #(
		.INIT('h8)
	) name2699 (
		_w3223_,
		_w3229_,
		_w3231_
	);
	LUT2 #(
		.INIT('h1)
	) name2700 (
		\ld_r_reg/P0001 ,
		_w3230_,
		_w3232_
	);
	LUT2 #(
		.INIT('h4)
	) name2701 (
		_w3231_,
		_w3232_,
		_w3233_
	);
	LUT2 #(
		.INIT('h1)
	) name2702 (
		\text_in_r_reg[14]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w3234_
	);
	LUT2 #(
		.INIT('h8)
	) name2703 (
		\text_in_r_reg[14]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w3235_
	);
	LUT2 #(
		.INIT('h2)
	) name2704 (
		\ld_r_reg/P0001 ,
		_w3234_,
		_w3236_
	);
	LUT2 #(
		.INIT('h4)
	) name2705 (
		_w3235_,
		_w3236_,
		_w3237_
	);
	LUT2 #(
		.INIT('h1)
	) name2706 (
		_w3233_,
		_w3237_,
		_w3238_
	);
	LUT2 #(
		.INIT('h1)
	) name2707 (
		_w1909_,
		_w1937_,
		_w3239_
	);
	LUT2 #(
		.INIT('h1)
	) name2708 (
		\sa32_reg[2]/P0001 ,
		_w3239_,
		_w3240_
	);
	LUT2 #(
		.INIT('h1)
	) name2709 (
		_w2351_,
		_w3240_,
		_w3241_
	);
	LUT2 #(
		.INIT('h2)
	) name2710 (
		\sa32_reg[1]/P0001 ,
		_w3241_,
		_w3242_
	);
	LUT2 #(
		.INIT('h1)
	) name2711 (
		_w1915_,
		_w1948_,
		_w3243_
	);
	LUT2 #(
		.INIT('h2)
	) name2712 (
		_w2026_,
		_w3243_,
		_w3244_
	);
	LUT2 #(
		.INIT('h8)
	) name2713 (
		_w1909_,
		_w1953_,
		_w3245_
	);
	LUT2 #(
		.INIT('h8)
	) name2714 (
		_w1919_,
		_w1934_,
		_w3246_
	);
	LUT2 #(
		.INIT('h1)
	) name2715 (
		_w3245_,
		_w3246_,
		_w3247_
	);
	LUT2 #(
		.INIT('h1)
	) name2716 (
		\sa32_reg[2]/P0001 ,
		_w3247_,
		_w3248_
	);
	LUT2 #(
		.INIT('h4)
	) name2717 (
		\sa32_reg[3]/P0001 ,
		_w1910_,
		_w3249_
	);
	LUT2 #(
		.INIT('h1)
	) name2718 (
		_w1941_,
		_w3146_,
		_w3250_
	);
	LUT2 #(
		.INIT('h8)
	) name2719 (
		_w2312_,
		_w3250_,
		_w3251_
	);
	LUT2 #(
		.INIT('h2)
	) name2720 (
		\sa32_reg[2]/P0001 ,
		_w3251_,
		_w3252_
	);
	LUT2 #(
		.INIT('h8)
	) name2721 (
		_w2041_,
		_w2313_,
		_w3253_
	);
	LUT2 #(
		.INIT('h8)
	) name2722 (
		\sa32_reg[4]/P0001 ,
		_w3253_,
		_w3254_
	);
	LUT2 #(
		.INIT('h2)
	) name2723 (
		\sa32_reg[5]/P0001 ,
		_w1923_,
		_w3255_
	);
	LUT2 #(
		.INIT('h2)
	) name2724 (
		_w1951_,
		_w3255_,
		_w3256_
	);
	LUT2 #(
		.INIT('h8)
	) name2725 (
		_w1934_,
		_w1995_,
		_w3257_
	);
	LUT2 #(
		.INIT('h1)
	) name2726 (
		_w1963_,
		_w1978_,
		_w3258_
	);
	LUT2 #(
		.INIT('h4)
	) name2727 (
		_w2009_,
		_w3258_,
		_w3259_
	);
	LUT2 #(
		.INIT('h2)
	) name2728 (
		\sa32_reg[2]/P0001 ,
		_w3259_,
		_w3260_
	);
	LUT2 #(
		.INIT('h1)
	) name2729 (
		_w3256_,
		_w3257_,
		_w3261_
	);
	LUT2 #(
		.INIT('h4)
	) name2730 (
		_w3254_,
		_w3261_,
		_w3262_
	);
	LUT2 #(
		.INIT('h4)
	) name2731 (
		_w3260_,
		_w3262_,
		_w3263_
	);
	LUT2 #(
		.INIT('h1)
	) name2732 (
		\sa32_reg[1]/P0001 ,
		_w3263_,
		_w3264_
	);
	LUT2 #(
		.INIT('h1)
	) name2733 (
		_w3244_,
		_w3249_,
		_w3265_
	);
	LUT2 #(
		.INIT('h4)
	) name2734 (
		_w3116_,
		_w3265_,
		_w3266_
	);
	LUT2 #(
		.INIT('h4)
	) name2735 (
		_w3248_,
		_w3266_,
		_w3267_
	);
	LUT2 #(
		.INIT('h4)
	) name2736 (
		_w3242_,
		_w3267_,
		_w3268_
	);
	LUT2 #(
		.INIT('h4)
	) name2737 (
		_w3252_,
		_w3268_,
		_w3269_
	);
	LUT2 #(
		.INIT('h4)
	) name2738 (
		_w3264_,
		_w3269_,
		_w3270_
	);
	LUT2 #(
		.INIT('h2)
	) name2739 (
		\sa32_reg[0]/P0002 ,
		_w3270_,
		_w3271_
	);
	LUT2 #(
		.INIT('h4)
	) name2740 (
		\sa32_reg[1]/P0001 ,
		_w1920_,
		_w3272_
	);
	LUT2 #(
		.INIT('h4)
	) name2741 (
		_w1947_,
		_w3272_,
		_w3273_
	);
	LUT2 #(
		.INIT('h1)
	) name2742 (
		_w1915_,
		_w2060_,
		_w3274_
	);
	LUT2 #(
		.INIT('h2)
	) name2743 (
		_w1951_,
		_w3274_,
		_w3275_
	);
	LUT2 #(
		.INIT('h2)
	) name2744 (
		\sa32_reg[2]/P0001 ,
		_w3273_,
		_w3276_
	);
	LUT2 #(
		.INIT('h4)
	) name2745 (
		_w3275_,
		_w3276_,
		_w3277_
	);
	LUT2 #(
		.INIT('h8)
	) name2746 (
		\sa32_reg[7]/P0001 ,
		_w1947_,
		_w3278_
	);
	LUT2 #(
		.INIT('h8)
	) name2747 (
		\sa32_reg[5]/P0001 ,
		_w3278_,
		_w3279_
	);
	LUT2 #(
		.INIT('h1)
	) name2748 (
		_w1941_,
		_w3279_,
		_w3280_
	);
	LUT2 #(
		.INIT('h1)
	) name2749 (
		\sa32_reg[2]/P0001 ,
		_w2382_,
		_w3281_
	);
	LUT2 #(
		.INIT('h8)
	) name2750 (
		_w3280_,
		_w3281_,
		_w3282_
	);
	LUT2 #(
		.INIT('h1)
	) name2751 (
		_w3277_,
		_w3282_,
		_w3283_
	);
	LUT2 #(
		.INIT('h8)
	) name2752 (
		_w1947_,
		_w1953_,
		_w3284_
	);
	LUT2 #(
		.INIT('h8)
	) name2753 (
		_w2313_,
		_w2387_,
		_w3285_
	);
	LUT2 #(
		.INIT('h8)
	) name2754 (
		\sa32_reg[3]/P0001 ,
		_w2068_,
		_w3286_
	);
	LUT2 #(
		.INIT('h4)
	) name2755 (
		_w1912_,
		_w1913_,
		_w3287_
	);
	LUT2 #(
		.INIT('h2)
	) name2756 (
		\sa32_reg[1]/P0001 ,
		_w3284_,
		_w3288_
	);
	LUT2 #(
		.INIT('h1)
	) name2757 (
		_w3285_,
		_w3287_,
		_w3289_
	);
	LUT2 #(
		.INIT('h8)
	) name2758 (
		_w3288_,
		_w3289_,
		_w3290_
	);
	LUT2 #(
		.INIT('h4)
	) name2759 (
		_w3286_,
		_w3290_,
		_w3291_
	);
	LUT2 #(
		.INIT('h8)
	) name2760 (
		_w1915_,
		_w1948_,
		_w3292_
	);
	LUT2 #(
		.INIT('h1)
	) name2761 (
		_w2346_,
		_w3292_,
		_w3293_
	);
	LUT2 #(
		.INIT('h1)
	) name2762 (
		\sa32_reg[3]/P0001 ,
		_w3293_,
		_w3294_
	);
	LUT2 #(
		.INIT('h1)
	) name2763 (
		\sa32_reg[1]/P0001 ,
		_w3175_,
		_w3295_
	);
	LUT2 #(
		.INIT('h4)
	) name2764 (
		_w3294_,
		_w3295_,
		_w3296_
	);
	LUT2 #(
		.INIT('h1)
	) name2765 (
		_w3291_,
		_w3296_,
		_w3297_
	);
	LUT2 #(
		.INIT('h1)
	) name2766 (
		_w3283_,
		_w3297_,
		_w3298_
	);
	LUT2 #(
		.INIT('h1)
	) name2767 (
		\sa32_reg[0]/P0002 ,
		_w3298_,
		_w3299_
	);
	LUT2 #(
		.INIT('h8)
	) name2768 (
		_w1995_,
		_w2068_,
		_w3300_
	);
	LUT2 #(
		.INIT('h4)
	) name2769 (
		\sa32_reg[2]/P0001 ,
		_w3284_,
		_w3301_
	);
	LUT2 #(
		.INIT('h8)
	) name2770 (
		\sa32_reg[7]/P0001 ,
		_w2382_,
		_w3302_
	);
	LUT2 #(
		.INIT('h1)
	) name2771 (
		_w2345_,
		_w3302_,
		_w3303_
	);
	LUT2 #(
		.INIT('h2)
	) name2772 (
		\sa32_reg[2]/P0001 ,
		_w3303_,
		_w3304_
	);
	LUT2 #(
		.INIT('h4)
	) name2773 (
		_w1970_,
		_w1982_,
		_w3305_
	);
	LUT2 #(
		.INIT('h1)
	) name2774 (
		_w3126_,
		_w3305_,
		_w3306_
	);
	LUT2 #(
		.INIT('h1)
	) name2775 (
		\sa32_reg[2]/P0001 ,
		_w3306_,
		_w3307_
	);
	LUT2 #(
		.INIT('h8)
	) name2776 (
		_w1934_,
		_w2026_,
		_w3308_
	);
	LUT2 #(
		.INIT('h8)
	) name2777 (
		_w1954_,
		_w3308_,
		_w3309_
	);
	LUT2 #(
		.INIT('h1)
	) name2778 (
		\sa32_reg[1]/P0001 ,
		_w3309_,
		_w3310_
	);
	LUT2 #(
		.INIT('h4)
	) name2779 (
		_w2062_,
		_w3310_,
		_w3311_
	);
	LUT2 #(
		.INIT('h4)
	) name2780 (
		_w3304_,
		_w3311_,
		_w3312_
	);
	LUT2 #(
		.INIT('h4)
	) name2781 (
		_w3307_,
		_w3312_,
		_w3313_
	);
	LUT2 #(
		.INIT('h1)
	) name2782 (
		_w2040_,
		_w3115_,
		_w3314_
	);
	LUT2 #(
		.INIT('h1)
	) name2783 (
		\sa32_reg[5]/P0001 ,
		_w3314_,
		_w3315_
	);
	LUT2 #(
		.INIT('h8)
	) name2784 (
		_w2041_,
		_w2059_,
		_w3316_
	);
	LUT2 #(
		.INIT('h4)
	) name2785 (
		\sa32_reg[2]/P0001 ,
		_w1921_,
		_w3317_
	);
	LUT2 #(
		.INIT('h1)
	) name2786 (
		_w3316_,
		_w3317_,
		_w3318_
	);
	LUT2 #(
		.INIT('h8)
	) name2787 (
		_w3179_,
		_w3318_,
		_w3319_
	);
	LUT2 #(
		.INIT('h4)
	) name2788 (
		_w3315_,
		_w3319_,
		_w3320_
	);
	LUT2 #(
		.INIT('h1)
	) name2789 (
		_w3313_,
		_w3320_,
		_w3321_
	);
	LUT2 #(
		.INIT('h1)
	) name2790 (
		_w3300_,
		_w3301_,
		_w3322_
	);
	LUT2 #(
		.INIT('h4)
	) name2791 (
		_w3299_,
		_w3322_,
		_w3323_
	);
	LUT2 #(
		.INIT('h4)
	) name2792 (
		_w3321_,
		_w3323_,
		_w3324_
	);
	LUT2 #(
		.INIT('h4)
	) name2793 (
		_w3271_,
		_w3324_,
		_w3325_
	);
	LUT2 #(
		.INIT('h8)
	) name2794 (
		_w2059_,
		_w3149_,
		_w3326_
	);
	LUT2 #(
		.INIT('h1)
	) name2795 (
		_w1952_,
		_w2030_,
		_w3327_
	);
	LUT2 #(
		.INIT('h2)
	) name2796 (
		\sa32_reg[7]/P0001 ,
		_w3327_,
		_w3328_
	);
	LUT2 #(
		.INIT('h1)
	) name2797 (
		_w3326_,
		_w3328_,
		_w3329_
	);
	LUT2 #(
		.INIT('h1)
	) name2798 (
		\sa32_reg[1]/P0001 ,
		_w3329_,
		_w3330_
	);
	LUT2 #(
		.INIT('h8)
	) name2799 (
		\sa32_reg[4]/P0001 ,
		_w2060_,
		_w3331_
	);
	LUT2 #(
		.INIT('h1)
	) name2800 (
		_w3245_,
		_w3331_,
		_w3332_
	);
	LUT2 #(
		.INIT('h2)
	) name2801 (
		_w2059_,
		_w3332_,
		_w3333_
	);
	LUT2 #(
		.INIT('h2)
	) name2802 (
		\sa32_reg[1]/P0001 ,
		_w1951_,
		_w3334_
	);
	LUT2 #(
		.INIT('h8)
	) name2803 (
		\sa32_reg[2]/P0001 ,
		_w1937_,
		_w3335_
	);
	LUT2 #(
		.INIT('h4)
	) name2804 (
		_w3334_,
		_w3335_,
		_w3336_
	);
	LUT2 #(
		.INIT('h1)
	) name2805 (
		_w2012_,
		_w3257_,
		_w3337_
	);
	LUT2 #(
		.INIT('h4)
	) name2806 (
		\sa32_reg[6]/NET0131 ,
		_w2028_,
		_w3338_
	);
	LUT2 #(
		.INIT('h1)
	) name2807 (
		_w2052_,
		_w3338_,
		_w3339_
	);
	LUT2 #(
		.INIT('h8)
	) name2808 (
		_w3337_,
		_w3339_,
		_w3340_
	);
	LUT2 #(
		.INIT('h1)
	) name2809 (
		\sa32_reg[2]/P0001 ,
		_w3340_,
		_w3341_
	);
	LUT2 #(
		.INIT('h4)
	) name2810 (
		\sa32_reg[6]/NET0131 ,
		_w1912_,
		_w3342_
	);
	LUT2 #(
		.INIT('h1)
	) name2811 (
		_w2366_,
		_w3342_,
		_w3343_
	);
	LUT2 #(
		.INIT('h1)
	) name2812 (
		\sa32_reg[2]/P0001 ,
		_w3343_,
		_w3344_
	);
	LUT2 #(
		.INIT('h8)
	) name2813 (
		\sa32_reg[4]/P0001 ,
		_w1915_,
		_w3345_
	);
	LUT2 #(
		.INIT('h8)
	) name2814 (
		_w2397_,
		_w3345_,
		_w3346_
	);
	LUT2 #(
		.INIT('h1)
	) name2815 (
		_w2352_,
		_w2383_,
		_w3347_
	);
	LUT2 #(
		.INIT('h4)
	) name2816 (
		_w3346_,
		_w3347_,
		_w3348_
	);
	LUT2 #(
		.INIT('h4)
	) name2817 (
		_w3344_,
		_w3348_,
		_w3349_
	);
	LUT2 #(
		.INIT('h2)
	) name2818 (
		\sa32_reg[1]/P0001 ,
		_w3349_,
		_w3350_
	);
	LUT2 #(
		.INIT('h1)
	) name2819 (
		_w3333_,
		_w3336_,
		_w3351_
	);
	LUT2 #(
		.INIT('h4)
	) name2820 (
		_w3330_,
		_w3351_,
		_w3352_
	);
	LUT2 #(
		.INIT('h4)
	) name2821 (
		_w3341_,
		_w3352_,
		_w3353_
	);
	LUT2 #(
		.INIT('h4)
	) name2822 (
		_w3350_,
		_w3353_,
		_w3354_
	);
	LUT2 #(
		.INIT('h1)
	) name2823 (
		\sa32_reg[0]/P0002 ,
		_w3354_,
		_w3355_
	);
	LUT2 #(
		.INIT('h4)
	) name2824 (
		\sa32_reg[5]/P0001 ,
		_w1951_,
		_w3356_
	);
	LUT2 #(
		.INIT('h1)
	) name2825 (
		_w2050_,
		_w3356_,
		_w3357_
	);
	LUT2 #(
		.INIT('h2)
	) name2826 (
		\sa32_reg[6]/NET0131 ,
		_w3357_,
		_w3358_
	);
	LUT2 #(
		.INIT('h1)
	) name2827 (
		_w1940_,
		_w1978_,
		_w3359_
	);
	LUT2 #(
		.INIT('h4)
	) name2828 (
		_w3358_,
		_w3359_,
		_w3360_
	);
	LUT2 #(
		.INIT('h2)
	) name2829 (
		\sa32_reg[2]/P0001 ,
		_w3360_,
		_w3361_
	);
	LUT2 #(
		.INIT('h8)
	) name2830 (
		_w2313_,
		_w2315_,
		_w3362_
	);
	LUT2 #(
		.INIT('h2)
	) name2831 (
		\sa32_reg[4]/P0001 ,
		_w1939_,
		_w3363_
	);
	LUT2 #(
		.INIT('h4)
	) name2832 (
		_w1988_,
		_w3363_,
		_w3364_
	);
	LUT2 #(
		.INIT('h1)
	) name2833 (
		_w1910_,
		_w3364_,
		_w3365_
	);
	LUT2 #(
		.INIT('h1)
	) name2834 (
		\sa32_reg[2]/P0001 ,
		_w3365_,
		_w3366_
	);
	LUT2 #(
		.INIT('h4)
	) name2835 (
		\sa32_reg[5]/P0001 ,
		_w2050_,
		_w3367_
	);
	LUT2 #(
		.INIT('h8)
	) name2836 (
		\sa32_reg[2]/P0001 ,
		_w3367_,
		_w3368_
	);
	LUT2 #(
		.INIT('h2)
	) name2837 (
		_w1982_,
		_w2348_,
		_w3369_
	);
	LUT2 #(
		.INIT('h1)
	) name2838 (
		_w3129_,
		_w3369_,
		_w3370_
	);
	LUT2 #(
		.INIT('h4)
	) name2839 (
		_w3368_,
		_w3370_,
		_w3371_
	);
	LUT2 #(
		.INIT('h4)
	) name2840 (
		_w3366_,
		_w3371_,
		_w3372_
	);
	LUT2 #(
		.INIT('h1)
	) name2841 (
		\sa32_reg[1]/P0001 ,
		_w3372_,
		_w3373_
	);
	LUT2 #(
		.INIT('h8)
	) name2842 (
		\sa32_reg[4]/P0001 ,
		_w1990_,
		_w3374_
	);
	LUT2 #(
		.INIT('h1)
	) name2843 (
		_w1954_,
		_w3374_,
		_w3375_
	);
	LUT2 #(
		.INIT('h4)
	) name2844 (
		\sa32_reg[3]/P0001 ,
		_w1913_,
		_w3376_
	);
	LUT2 #(
		.INIT('h1)
	) name2845 (
		_w1969_,
		_w3376_,
		_w3377_
	);
	LUT2 #(
		.INIT('h8)
	) name2846 (
		_w3375_,
		_w3377_,
		_w3378_
	);
	LUT2 #(
		.INIT('h2)
	) name2847 (
		\sa32_reg[2]/P0001 ,
		_w3378_,
		_w3379_
	);
	LUT2 #(
		.INIT('h1)
	) name2848 (
		_w3117_,
		_w3253_,
		_w3380_
	);
	LUT2 #(
		.INIT('h4)
	) name2849 (
		_w3379_,
		_w3380_,
		_w3381_
	);
	LUT2 #(
		.INIT('h2)
	) name2850 (
		\sa32_reg[1]/P0001 ,
		_w3381_,
		_w3382_
	);
	LUT2 #(
		.INIT('h1)
	) name2851 (
		_w3246_,
		_w3362_,
		_w3383_
	);
	LUT2 #(
		.INIT('h4)
	) name2852 (
		_w3361_,
		_w3383_,
		_w3384_
	);
	LUT2 #(
		.INIT('h4)
	) name2853 (
		_w3373_,
		_w3384_,
		_w3385_
	);
	LUT2 #(
		.INIT('h4)
	) name2854 (
		_w3382_,
		_w3385_,
		_w3386_
	);
	LUT2 #(
		.INIT('h2)
	) name2855 (
		\sa32_reg[0]/P0002 ,
		_w3386_,
		_w3387_
	);
	LUT2 #(
		.INIT('h2)
	) name2856 (
		\sa32_reg[2]/P0001 ,
		_w1921_,
		_w3388_
	);
	LUT2 #(
		.INIT('h1)
	) name2857 (
		_w1921_,
		_w2388_,
		_w3389_
	);
	LUT2 #(
		.INIT('h8)
	) name2858 (
		_w3337_,
		_w3389_,
		_w3390_
	);
	LUT2 #(
		.INIT('h1)
	) name2859 (
		_w3388_,
		_w3390_,
		_w3391_
	);
	LUT2 #(
		.INIT('h4)
	) name2860 (
		\sa32_reg[3]/P0001 ,
		_w3124_,
		_w3392_
	);
	LUT2 #(
		.INIT('h1)
	) name2861 (
		_w1992_,
		_w3117_,
		_w3393_
	);
	LUT2 #(
		.INIT('h4)
	) name2862 (
		_w3392_,
		_w3393_,
		_w3394_
	);
	LUT2 #(
		.INIT('h2)
	) name2863 (
		\sa32_reg[2]/P0001 ,
		_w3394_,
		_w3395_
	);
	LUT2 #(
		.INIT('h1)
	) name2864 (
		_w3391_,
		_w3395_,
		_w3396_
	);
	LUT2 #(
		.INIT('h1)
	) name2865 (
		\sa32_reg[1]/P0001 ,
		_w3396_,
		_w3397_
	);
	LUT2 #(
		.INIT('h1)
	) name2866 (
		_w1996_,
		_w3162_,
		_w3398_
	);
	LUT2 #(
		.INIT('h1)
	) name2867 (
		\sa32_reg[2]/P0001 ,
		_w3398_,
		_w3399_
	);
	LUT2 #(
		.INIT('h2)
	) name2868 (
		_w1939_,
		_w2049_,
		_w3400_
	);
	LUT2 #(
		.INIT('h2)
	) name2869 (
		_w3293_,
		_w3400_,
		_w3401_
	);
	LUT2 #(
		.INIT('h8)
	) name2870 (
		\sa32_reg[1]/P0001 ,
		_w2026_,
		_w3402_
	);
	LUT2 #(
		.INIT('h4)
	) name2871 (
		_w3401_,
		_w3402_,
		_w3403_
	);
	LUT2 #(
		.INIT('h2)
	) name2872 (
		\sa32_reg[7]/P0001 ,
		_w3375_,
		_w3404_
	);
	LUT2 #(
		.INIT('h8)
	) name2873 (
		_w1913_,
		_w1970_,
		_w3405_
	);
	LUT2 #(
		.INIT('h1)
	) name2874 (
		_w3404_,
		_w3405_,
		_w3406_
	);
	LUT2 #(
		.INIT('h1)
	) name2875 (
		\sa32_reg[3]/P0001 ,
		_w3406_,
		_w3407_
	);
	LUT2 #(
		.INIT('h8)
	) name2876 (
		_w1954_,
		_w2387_,
		_w3408_
	);
	LUT2 #(
		.INIT('h1)
	) name2877 (
		_w1911_,
		_w3408_,
		_w3409_
	);
	LUT2 #(
		.INIT('h4)
	) name2878 (
		_w3407_,
		_w3409_,
		_w3410_
	);
	LUT2 #(
		.INIT('h2)
	) name2879 (
		_w2370_,
		_w3410_,
		_w3411_
	);
	LUT2 #(
		.INIT('h1)
	) name2880 (
		_w3399_,
		_w3403_,
		_w3412_
	);
	LUT2 #(
		.INIT('h4)
	) name2881 (
		_w3397_,
		_w3412_,
		_w3413_
	);
	LUT2 #(
		.INIT('h4)
	) name2882 (
		_w3411_,
		_w3413_,
		_w3414_
	);
	LUT2 #(
		.INIT('h4)
	) name2883 (
		_w3355_,
		_w3414_,
		_w3415_
	);
	LUT2 #(
		.INIT('h4)
	) name2884 (
		_w3387_,
		_w3415_,
		_w3416_
	);
	LUT2 #(
		.INIT('h2)
	) name2885 (
		_w3325_,
		_w3416_,
		_w3417_
	);
	LUT2 #(
		.INIT('h4)
	) name2886 (
		_w3325_,
		_w3416_,
		_w3418_
	);
	LUT2 #(
		.INIT('h1)
	) name2887 (
		_w3417_,
		_w3418_,
		_w3419_
	);
	LUT2 #(
		.INIT('h1)
	) name2888 (
		_w2012_,
		_w2398_,
		_w3420_
	);
	LUT2 #(
		.INIT('h2)
	) name2889 (
		\sa32_reg[2]/P0001 ,
		_w3420_,
		_w3421_
	);
	LUT2 #(
		.INIT('h4)
	) name2890 (
		\sa32_reg[4]/P0001 ,
		_w1990_,
		_w3422_
	);
	LUT2 #(
		.INIT('h8)
	) name2891 (
		\sa32_reg[3]/P0001 ,
		_w3345_,
		_w3423_
	);
	LUT2 #(
		.INIT('h1)
	) name2892 (
		_w2389_,
		_w3422_,
		_w3424_
	);
	LUT2 #(
		.INIT('h4)
	) name2893 (
		_w3423_,
		_w3424_,
		_w3425_
	);
	LUT2 #(
		.INIT('h1)
	) name2894 (
		\sa32_reg[2]/P0001 ,
		_w3425_,
		_w3426_
	);
	LUT2 #(
		.INIT('h2)
	) name2895 (
		_w1950_,
		_w1992_,
		_w3427_
	);
	LUT2 #(
		.INIT('h4)
	) name2896 (
		_w3421_,
		_w3427_,
		_w3428_
	);
	LUT2 #(
		.INIT('h4)
	) name2897 (
		_w3426_,
		_w3428_,
		_w3429_
	);
	LUT2 #(
		.INIT('h2)
	) name2898 (
		\sa32_reg[1]/P0001 ,
		_w3429_,
		_w3430_
	);
	LUT2 #(
		.INIT('h1)
	) name2899 (
		_w2009_,
		_w2362_,
		_w3431_
	);
	LUT2 #(
		.INIT('h2)
	) name2900 (
		\sa32_reg[2]/P0001 ,
		_w3431_,
		_w3432_
	);
	LUT2 #(
		.INIT('h1)
	) name2901 (
		_w1941_,
		_w3134_,
		_w3433_
	);
	LUT2 #(
		.INIT('h1)
	) name2902 (
		\sa32_reg[2]/P0001 ,
		_w3433_,
		_w3434_
	);
	LUT2 #(
		.INIT('h1)
	) name2903 (
		_w3194_,
		_w3249_,
		_w3435_
	);
	LUT2 #(
		.INIT('h2)
	) name2904 (
		\sa32_reg[2]/P0001 ,
		_w3435_,
		_w3436_
	);
	LUT2 #(
		.INIT('h8)
	) name2905 (
		_w1924_,
		_w2315_,
		_w3437_
	);
	LUT2 #(
		.INIT('h1)
	) name2906 (
		_w2317_,
		_w2351_,
		_w3438_
	);
	LUT2 #(
		.INIT('h1)
	) name2907 (
		\sa32_reg[2]/P0001 ,
		_w3438_,
		_w3439_
	);
	LUT2 #(
		.INIT('h1)
	) name2908 (
		_w3134_,
		_w3437_,
		_w3440_
	);
	LUT2 #(
		.INIT('h4)
	) name2909 (
		_w3436_,
		_w3440_,
		_w3441_
	);
	LUT2 #(
		.INIT('h4)
	) name2910 (
		_w3439_,
		_w3441_,
		_w3442_
	);
	LUT2 #(
		.INIT('h1)
	) name2911 (
		\sa32_reg[1]/P0001 ,
		_w3442_,
		_w3443_
	);
	LUT2 #(
		.INIT('h1)
	) name2912 (
		_w2040_,
		_w2062_,
		_w3444_
	);
	LUT2 #(
		.INIT('h4)
	) name2913 (
		_w3432_,
		_w3444_,
		_w3445_
	);
	LUT2 #(
		.INIT('h4)
	) name2914 (
		_w3434_,
		_w3445_,
		_w3446_
	);
	LUT2 #(
		.INIT('h4)
	) name2915 (
		_w3430_,
		_w3446_,
		_w3447_
	);
	LUT2 #(
		.INIT('h4)
	) name2916 (
		_w3443_,
		_w3447_,
		_w3448_
	);
	LUT2 #(
		.INIT('h1)
	) name2917 (
		\sa32_reg[0]/P0002 ,
		_w3448_,
		_w3449_
	);
	LUT2 #(
		.INIT('h8)
	) name2918 (
		_w1909_,
		_w2334_,
		_w3450_
	);
	LUT2 #(
		.INIT('h1)
	) name2919 (
		_w3408_,
		_w3450_,
		_w3451_
	);
	LUT2 #(
		.INIT('h1)
	) name2920 (
		_w3145_,
		_w3278_,
		_w3452_
	);
	LUT2 #(
		.INIT('h4)
	) name2921 (
		_w3345_,
		_w3452_,
		_w3453_
	);
	LUT2 #(
		.INIT('h2)
	) name2922 (
		\sa32_reg[2]/P0001 ,
		_w3453_,
		_w3454_
	);
	LUT2 #(
		.INIT('h2)
	) name2923 (
		_w3451_,
		_w3454_,
		_w3455_
	);
	LUT2 #(
		.INIT('h2)
	) name2924 (
		\sa32_reg[0]/P0002 ,
		_w3455_,
		_w3456_
	);
	LUT2 #(
		.INIT('h4)
	) name2925 (
		\sa32_reg[3]/P0001 ,
		_w1939_,
		_w3457_
	);
	LUT2 #(
		.INIT('h1)
	) name2926 (
		_w2033_,
		_w3457_,
		_w3458_
	);
	LUT2 #(
		.INIT('h1)
	) name2927 (
		_w1953_,
		_w3458_,
		_w3459_
	);
	LUT2 #(
		.INIT('h1)
	) name2928 (
		_w1992_,
		_w2324_,
		_w3460_
	);
	LUT2 #(
		.INIT('h4)
	) name2929 (
		_w3459_,
		_w3460_,
		_w3461_
	);
	LUT2 #(
		.INIT('h1)
	) name2930 (
		\sa32_reg[2]/P0001 ,
		_w3461_,
		_w3462_
	);
	LUT2 #(
		.INIT('h1)
	) name2931 (
		_w3456_,
		_w3462_,
		_w3463_
	);
	LUT2 #(
		.INIT('h2)
	) name2932 (
		\sa32_reg[1]/P0001 ,
		_w3463_,
		_w3464_
	);
	LUT2 #(
		.INIT('h1)
	) name2933 (
		_w2352_,
		_w3292_,
		_w3465_
	);
	LUT2 #(
		.INIT('h1)
	) name2934 (
		_w3249_,
		_w3331_,
		_w3466_
	);
	LUT2 #(
		.INIT('h8)
	) name2935 (
		_w3465_,
		_w3466_,
		_w3467_
	);
	LUT2 #(
		.INIT('h1)
	) name2936 (
		\sa32_reg[2]/P0001 ,
		_w3467_,
		_w3468_
	);
	LUT2 #(
		.INIT('h2)
	) name2937 (
		_w1988_,
		_w2030_,
		_w3469_
	);
	LUT2 #(
		.INIT('h4)
	) name2938 (
		\sa32_reg[1]/P0001 ,
		_w1994_,
		_w3470_
	);
	LUT2 #(
		.INIT('h1)
	) name2939 (
		_w3331_,
		_w3469_,
		_w3471_
	);
	LUT2 #(
		.INIT('h4)
	) name2940 (
		_w3470_,
		_w3471_,
		_w3472_
	);
	LUT2 #(
		.INIT('h1)
	) name2941 (
		\sa32_reg[3]/P0001 ,
		_w3472_,
		_w3473_
	);
	LUT2 #(
		.INIT('h2)
	) name2942 (
		_w1932_,
		_w2348_,
		_w3474_
	);
	LUT2 #(
		.INIT('h1)
	) name2943 (
		_w1935_,
		_w3292_,
		_w3475_
	);
	LUT2 #(
		.INIT('h4)
	) name2944 (
		_w3474_,
		_w3475_,
		_w3476_
	);
	LUT2 #(
		.INIT('h1)
	) name2945 (
		\sa32_reg[1]/P0001 ,
		_w3476_,
		_w3477_
	);
	LUT2 #(
		.INIT('h1)
	) name2946 (
		_w3468_,
		_w3477_,
		_w3478_
	);
	LUT2 #(
		.INIT('h4)
	) name2947 (
		_w3473_,
		_w3478_,
		_w3479_
	);
	LUT2 #(
		.INIT('h2)
	) name2948 (
		\sa32_reg[0]/P0002 ,
		_w3479_,
		_w3480_
	);
	LUT2 #(
		.INIT('h2)
	) name2949 (
		_w1988_,
		_w3127_,
		_w3481_
	);
	LUT2 #(
		.INIT('h8)
	) name2950 (
		\sa32_reg[3]/P0001 ,
		_w3124_,
		_w3482_
	);
	LUT2 #(
		.INIT('h1)
	) name2951 (
		_w3481_,
		_w3482_,
		_w3483_
	);
	LUT2 #(
		.INIT('h2)
	) name2952 (
		_w2370_,
		_w3483_,
		_w3484_
	);
	LUT2 #(
		.INIT('h1)
	) name2953 (
		_w2033_,
		_w3181_,
		_w3485_
	);
	LUT2 #(
		.INIT('h2)
	) name2954 (
		_w2059_,
		_w3485_,
		_w3486_
	);
	LUT2 #(
		.INIT('h1)
	) name2955 (
		_w2311_,
		_w2366_,
		_w3487_
	);
	LUT2 #(
		.INIT('h4)
	) name2956 (
		_w1938_,
		_w3487_,
		_w3488_
	);
	LUT2 #(
		.INIT('h1)
	) name2957 (
		\sa32_reg[2]/P0001 ,
		_w3488_,
		_w3489_
	);
	LUT2 #(
		.INIT('h8)
	) name2958 (
		_w1990_,
		_w2334_,
		_w3490_
	);
	LUT2 #(
		.INIT('h4)
	) name2959 (
		\sa32_reg[3]/P0001 ,
		_w2041_,
		_w3491_
	);
	LUT2 #(
		.INIT('h1)
	) name2960 (
		_w1922_,
		_w2040_,
		_w3492_
	);
	LUT2 #(
		.INIT('h4)
	) name2961 (
		_w3491_,
		_w3492_,
		_w3493_
	);
	LUT2 #(
		.INIT('h2)
	) name2962 (
		\sa32_reg[2]/P0001 ,
		_w3493_,
		_w3494_
	);
	LUT2 #(
		.INIT('h1)
	) name2963 (
		_w1936_,
		_w3490_,
		_w3495_
	);
	LUT2 #(
		.INIT('h4)
	) name2964 (
		_w3489_,
		_w3495_,
		_w3496_
	);
	LUT2 #(
		.INIT('h4)
	) name2965 (
		_w3494_,
		_w3496_,
		_w3497_
	);
	LUT2 #(
		.INIT('h1)
	) name2966 (
		\sa32_reg[1]/P0001 ,
		_w3497_,
		_w3498_
	);
	LUT2 #(
		.INIT('h1)
	) name2967 (
		_w3484_,
		_w3486_,
		_w3499_
	);
	LUT2 #(
		.INIT('h4)
	) name2968 (
		_w3498_,
		_w3499_,
		_w3500_
	);
	LUT2 #(
		.INIT('h4)
	) name2969 (
		_w3464_,
		_w3500_,
		_w3501_
	);
	LUT2 #(
		.INIT('h4)
	) name2970 (
		_w3480_,
		_w3501_,
		_w3502_
	);
	LUT2 #(
		.INIT('h4)
	) name2971 (
		_w3449_,
		_w3502_,
		_w3503_
	);
	LUT2 #(
		.INIT('h2)
	) name2972 (
		\u0_w_reg[3][9]/P0001 ,
		_w3503_,
		_w3504_
	);
	LUT2 #(
		.INIT('h4)
	) name2973 (
		\u0_w_reg[3][9]/P0001 ,
		_w3503_,
		_w3505_
	);
	LUT2 #(
		.INIT('h1)
	) name2974 (
		_w3504_,
		_w3505_,
		_w3506_
	);
	LUT2 #(
		.INIT('h8)
	) name2975 (
		_w3419_,
		_w3506_,
		_w3507_
	);
	LUT2 #(
		.INIT('h1)
	) name2976 (
		_w3419_,
		_w3506_,
		_w3508_
	);
	LUT2 #(
		.INIT('h1)
	) name2977 (
		_w3507_,
		_w3508_,
		_w3509_
	);
	LUT2 #(
		.INIT('h8)
	) name2978 (
		\sa21_reg[6]/NET0131 ,
		_w1750_,
		_w3510_
	);
	LUT2 #(
		.INIT('h1)
	) name2979 (
		_w2893_,
		_w3510_,
		_w3511_
	);
	LUT2 #(
		.INIT('h4)
	) name2980 (
		\sa21_reg[3]/P0001 ,
		_w1833_,
		_w3512_
	);
	LUT2 #(
		.INIT('h2)
	) name2981 (
		_w3511_,
		_w3512_,
		_w3513_
	);
	LUT2 #(
		.INIT('h1)
	) name2982 (
		\sa21_reg[2]/P0001 ,
		_w3513_,
		_w3514_
	);
	LUT2 #(
		.INIT('h8)
	) name2983 (
		_w1754_,
		_w2452_,
		_w3515_
	);
	LUT2 #(
		.INIT('h8)
	) name2984 (
		\sa21_reg[2]/P0001 ,
		_w2429_,
		_w3516_
	);
	LUT2 #(
		.INIT('h1)
	) name2985 (
		_w1802_,
		_w1841_,
		_w3517_
	);
	LUT2 #(
		.INIT('h8)
	) name2986 (
		\sa21_reg[3]/P0001 ,
		_w1840_,
		_w3518_
	);
	LUT2 #(
		.INIT('h1)
	) name2987 (
		_w3517_,
		_w3518_,
		_w3519_
	);
	LUT2 #(
		.INIT('h1)
	) name2988 (
		_w3515_,
		_w3516_,
		_w3520_
	);
	LUT2 #(
		.INIT('h4)
	) name2989 (
		_w3519_,
		_w3520_,
		_w3521_
	);
	LUT2 #(
		.INIT('h2)
	) name2990 (
		\sa21_reg[1]/P0001 ,
		_w3521_,
		_w3522_
	);
	LUT2 #(
		.INIT('h1)
	) name2991 (
		\sa21_reg[3]/P0001 ,
		_w2418_,
		_w3523_
	);
	LUT2 #(
		.INIT('h1)
	) name2992 (
		_w3028_,
		_w3523_,
		_w3524_
	);
	LUT2 #(
		.INIT('h1)
	) name2993 (
		\sa21_reg[1]/P0001 ,
		_w3524_,
		_w3525_
	);
	LUT2 #(
		.INIT('h1)
	) name2994 (
		_w1758_,
		_w2422_,
		_w3526_
	);
	LUT2 #(
		.INIT('h2)
	) name2995 (
		_w1895_,
		_w3526_,
		_w3527_
	);
	LUT2 #(
		.INIT('h1)
	) name2996 (
		_w1757_,
		_w1763_,
		_w3528_
	);
	LUT2 #(
		.INIT('h4)
	) name2997 (
		\sa21_reg[1]/P0001 ,
		\sa21_reg[2]/P0001 ,
		_w3529_
	);
	LUT2 #(
		.INIT('h8)
	) name2998 (
		\sa21_reg[5]/P0001 ,
		_w3529_,
		_w3530_
	);
	LUT2 #(
		.INIT('h4)
	) name2999 (
		_w3528_,
		_w3530_,
		_w3531_
	);
	LUT2 #(
		.INIT('h1)
	) name3000 (
		_w3527_,
		_w3531_,
		_w3532_
	);
	LUT2 #(
		.INIT('h4)
	) name3001 (
		_w3514_,
		_w3532_,
		_w3533_
	);
	LUT2 #(
		.INIT('h1)
	) name3002 (
		_w3522_,
		_w3525_,
		_w3534_
	);
	LUT2 #(
		.INIT('h8)
	) name3003 (
		_w3533_,
		_w3534_,
		_w3535_
	);
	LUT2 #(
		.INIT('h1)
	) name3004 (
		\sa21_reg[0]/P0001 ,
		_w3535_,
		_w3536_
	);
	LUT2 #(
		.INIT('h1)
	) name3005 (
		_w1834_,
		_w1872_,
		_w3537_
	);
	LUT2 #(
		.INIT('h4)
	) name3006 (
		_w2436_,
		_w3537_,
		_w3538_
	);
	LUT2 #(
		.INIT('h2)
	) name3007 (
		\sa21_reg[2]/P0001 ,
		_w3538_,
		_w3539_
	);
	LUT2 #(
		.INIT('h2)
	) name3008 (
		\sa21_reg[5]/P0001 ,
		_w1763_,
		_w3540_
	);
	LUT2 #(
		.INIT('h2)
	) name3009 (
		_w1866_,
		_w3540_,
		_w3541_
	);
	LUT2 #(
		.INIT('h4)
	) name3010 (
		\sa21_reg[6]/NET0131 ,
		_w1757_,
		_w3542_
	);
	LUT2 #(
		.INIT('h4)
	) name3011 (
		\sa21_reg[5]/P0001 ,
		_w3542_,
		_w3543_
	);
	LUT2 #(
		.INIT('h8)
	) name3012 (
		_w2455_,
		_w3543_,
		_w3544_
	);
	LUT2 #(
		.INIT('h8)
	) name3013 (
		_w1745_,
		_w1815_,
		_w3545_
	);
	LUT2 #(
		.INIT('h1)
	) name3014 (
		_w3541_,
		_w3545_,
		_w3546_
	);
	LUT2 #(
		.INIT('h4)
	) name3015 (
		_w3544_,
		_w3546_,
		_w3547_
	);
	LUT2 #(
		.INIT('h4)
	) name3016 (
		_w3539_,
		_w3547_,
		_w3548_
	);
	LUT2 #(
		.INIT('h1)
	) name3017 (
		\sa21_reg[1]/P0001 ,
		_w3548_,
		_w3549_
	);
	LUT2 #(
		.INIT('h1)
	) name3018 (
		_w1837_,
		_w2477_,
		_w3550_
	);
	LUT2 #(
		.INIT('h1)
	) name3019 (
		\sa21_reg[2]/P0001 ,
		_w3550_,
		_w3551_
	);
	LUT2 #(
		.INIT('h1)
	) name3020 (
		_w1884_,
		_w3551_,
		_w3552_
	);
	LUT2 #(
		.INIT('h2)
	) name3021 (
		\sa21_reg[1]/P0001 ,
		_w3552_,
		_w3553_
	);
	LUT2 #(
		.INIT('h8)
	) name3022 (
		\sa21_reg[3]/P0001 ,
		_w1758_,
		_w3554_
	);
	LUT2 #(
		.INIT('h1)
	) name3023 (
		\sa21_reg[2]/P0001 ,
		_w3554_,
		_w3555_
	);
	LUT2 #(
		.INIT('h1)
	) name3024 (
		_w2469_,
		_w2905_,
		_w3556_
	);
	LUT2 #(
		.INIT('h4)
	) name3025 (
		_w2489_,
		_w3556_,
		_w3557_
	);
	LUT2 #(
		.INIT('h8)
	) name3026 (
		_w3555_,
		_w3557_,
		_w3558_
	);
	LUT2 #(
		.INIT('h2)
	) name3027 (
		\sa21_reg[2]/P0001 ,
		_w2993_,
		_w3559_
	);
	LUT2 #(
		.INIT('h4)
	) name3028 (
		_w2893_,
		_w3559_,
		_w3560_
	);
	LUT2 #(
		.INIT('h8)
	) name3029 (
		_w1752_,
		_w3560_,
		_w3561_
	);
	LUT2 #(
		.INIT('h1)
	) name3030 (
		_w3558_,
		_w3561_,
		_w3562_
	);
	LUT2 #(
		.INIT('h1)
	) name3031 (
		_w1838_,
		_w3010_,
		_w3563_
	);
	LUT2 #(
		.INIT('h4)
	) name3032 (
		_w3553_,
		_w3563_,
		_w3564_
	);
	LUT2 #(
		.INIT('h4)
	) name3033 (
		_w3562_,
		_w3564_,
		_w3565_
	);
	LUT2 #(
		.INIT('h4)
	) name3034 (
		_w3549_,
		_w3565_,
		_w3566_
	);
	LUT2 #(
		.INIT('h2)
	) name3035 (
		\sa21_reg[0]/P0001 ,
		_w3566_,
		_w3567_
	);
	LUT2 #(
		.INIT('h8)
	) name3036 (
		_w1831_,
		_w1879_,
		_w3568_
	);
	LUT2 #(
		.INIT('h1)
	) name3037 (
		_w1821_,
		_w3568_,
		_w3569_
	);
	LUT2 #(
		.INIT('h2)
	) name3038 (
		\sa21_reg[6]/NET0131 ,
		_w3569_,
		_w3570_
	);
	LUT2 #(
		.INIT('h8)
	) name3039 (
		_w1745_,
		_w1877_,
		_w3571_
	);
	LUT2 #(
		.INIT('h8)
	) name3040 (
		_w1753_,
		_w3571_,
		_w3572_
	);
	LUT2 #(
		.INIT('h1)
	) name3041 (
		\sa21_reg[2]/P0001 ,
		_w2901_,
		_w3573_
	);
	LUT2 #(
		.INIT('h4)
	) name3042 (
		_w2451_,
		_w3573_,
		_w3574_
	);
	LUT2 #(
		.INIT('h4)
	) name3043 (
		_w3049_,
		_w3574_,
		_w3575_
	);
	LUT2 #(
		.INIT('h2)
	) name3044 (
		\sa21_reg[2]/P0001 ,
		_w1891_,
		_w3576_
	);
	LUT2 #(
		.INIT('h4)
	) name3045 (
		_w3055_,
		_w3576_,
		_w3577_
	);
	LUT2 #(
		.INIT('h1)
	) name3046 (
		_w3575_,
		_w3577_,
		_w3578_
	);
	LUT2 #(
		.INIT('h1)
	) name3047 (
		_w2928_,
		_w3572_,
		_w3579_
	);
	LUT2 #(
		.INIT('h4)
	) name3048 (
		_w3578_,
		_w3579_,
		_w3580_
	);
	LUT2 #(
		.INIT('h1)
	) name3049 (
		\sa21_reg[1]/P0001 ,
		_w3580_,
		_w3581_
	);
	LUT2 #(
		.INIT('h1)
	) name3050 (
		_w1788_,
		_w2865_,
		_w3582_
	);
	LUT2 #(
		.INIT('h2)
	) name3051 (
		\sa21_reg[2]/P0001 ,
		_w3582_,
		_w3583_
	);
	LUT2 #(
		.INIT('h8)
	) name3052 (
		_w1754_,
		_w1849_,
		_w3584_
	);
	LUT2 #(
		.INIT('h1)
	) name3053 (
		_w1883_,
		_w3020_,
		_w3585_
	);
	LUT2 #(
		.INIT('h4)
	) name3054 (
		_w3584_,
		_w3585_,
		_w3586_
	);
	LUT2 #(
		.INIT('h4)
	) name3055 (
		_w3583_,
		_w3586_,
		_w3587_
	);
	LUT2 #(
		.INIT('h2)
	) name3056 (
		\sa21_reg[1]/P0001 ,
		_w3587_,
		_w3588_
	);
	LUT2 #(
		.INIT('h1)
	) name3057 (
		_w3570_,
		_w3588_,
		_w3589_
	);
	LUT2 #(
		.INIT('h4)
	) name3058 (
		_w3581_,
		_w3589_,
		_w3590_
	);
	LUT2 #(
		.INIT('h4)
	) name3059 (
		_w3536_,
		_w3590_,
		_w3591_
	);
	LUT2 #(
		.INIT('h4)
	) name3060 (
		_w3567_,
		_w3591_,
		_w3592_
	);
	LUT2 #(
		.INIT('h2)
	) name3061 (
		_w2529_,
		_w3592_,
		_w3593_
	);
	LUT2 #(
		.INIT('h4)
	) name3062 (
		_w2529_,
		_w3592_,
		_w3594_
	);
	LUT2 #(
		.INIT('h1)
	) name3063 (
		_w3593_,
		_w3594_,
		_w3595_
	);
	LUT2 #(
		.INIT('h1)
	) name3064 (
		_w1639_,
		_w1708_,
		_w3596_
	);
	LUT2 #(
		.INIT('h1)
	) name3065 (
		\sa10_reg[2]/P0001 ,
		_w3596_,
		_w3597_
	);
	LUT2 #(
		.INIT('h8)
	) name3066 (
		_w1598_,
		_w1636_,
		_w3598_
	);
	LUT2 #(
		.INIT('h4)
	) name3067 (
		\sa10_reg[3]/P0001 ,
		_w2621_,
		_w3599_
	);
	LUT2 #(
		.INIT('h1)
	) name3068 (
		_w2607_,
		_w3599_,
		_w3600_
	);
	LUT2 #(
		.INIT('h2)
	) name3069 (
		\sa10_reg[2]/P0001 ,
		_w3600_,
		_w3601_
	);
	LUT2 #(
		.INIT('h1)
	) name3070 (
		_w2567_,
		_w3598_,
		_w3602_
	);
	LUT2 #(
		.INIT('h4)
	) name3071 (
		_w3597_,
		_w3602_,
		_w3603_
	);
	LUT2 #(
		.INIT('h4)
	) name3072 (
		_w3601_,
		_w3603_,
		_w3604_
	);
	LUT2 #(
		.INIT('h1)
	) name3073 (
		\sa10_reg[0]/P0001 ,
		_w3604_,
		_w3605_
	);
	LUT2 #(
		.INIT('h1)
	) name3074 (
		_w1628_,
		_w2130_,
		_w3606_
	);
	LUT2 #(
		.INIT('h4)
	) name3075 (
		_w2581_,
		_w3606_,
		_w3607_
	);
	LUT2 #(
		.INIT('h1)
	) name3076 (
		\sa10_reg[2]/P0001 ,
		_w3607_,
		_w3608_
	);
	LUT2 #(
		.INIT('h1)
	) name3077 (
		_w1631_,
		_w2558_,
		_w3609_
	);
	LUT2 #(
		.INIT('h4)
	) name3078 (
		_w3608_,
		_w3609_,
		_w3610_
	);
	LUT2 #(
		.INIT('h4)
	) name3079 (
		_w3605_,
		_w3610_,
		_w3611_
	);
	LUT2 #(
		.INIT('h1)
	) name3080 (
		\sa10_reg[1]/P0001 ,
		_w3611_,
		_w3612_
	);
	LUT2 #(
		.INIT('h8)
	) name3081 (
		_w1585_,
		_w1619_,
		_w3613_
	);
	LUT2 #(
		.INIT('h1)
	) name3082 (
		_w1609_,
		_w3613_,
		_w3614_
	);
	LUT2 #(
		.INIT('h2)
	) name3083 (
		\sa10_reg[5]/P0001 ,
		_w1681_,
		_w3615_
	);
	LUT2 #(
		.INIT('h2)
	) name3084 (
		\sa10_reg[4]/P0001 ,
		_w1681_,
		_w3616_
	);
	LUT2 #(
		.INIT('h2)
	) name3085 (
		\sa10_reg[7]/NET0131 ,
		_w3615_,
		_w3617_
	);
	LUT2 #(
		.INIT('h4)
	) name3086 (
		_w3616_,
		_w3617_,
		_w3618_
	);
	LUT2 #(
		.INIT('h1)
	) name3087 (
		_w1673_,
		_w3618_,
		_w3619_
	);
	LUT2 #(
		.INIT('h2)
	) name3088 (
		\sa10_reg[2]/P0001 ,
		_w3619_,
		_w3620_
	);
	LUT2 #(
		.INIT('h2)
	) name3089 (
		_w3614_,
		_w3620_,
		_w3621_
	);
	LUT2 #(
		.INIT('h2)
	) name3090 (
		\sa10_reg[1]/P0001 ,
		_w3621_,
		_w3622_
	);
	LUT2 #(
		.INIT('h4)
	) name3091 (
		\sa10_reg[6]/NET0131 ,
		_w2826_,
		_w3623_
	);
	LUT2 #(
		.INIT('h2)
	) name3092 (
		_w1594_,
		_w1652_,
		_w3624_
	);
	LUT2 #(
		.INIT('h4)
	) name3093 (
		_w1600_,
		_w3624_,
		_w3625_
	);
	LUT2 #(
		.INIT('h1)
	) name3094 (
		_w2093_,
		_w2778_,
		_w3626_
	);
	LUT2 #(
		.INIT('h4)
	) name3095 (
		_w3623_,
		_w3626_,
		_w3627_
	);
	LUT2 #(
		.INIT('h4)
	) name3096 (
		_w3625_,
		_w3627_,
		_w3628_
	);
	LUT2 #(
		.INIT('h1)
	) name3097 (
		\sa10_reg[1]/P0001 ,
		_w3628_,
		_w3629_
	);
	LUT2 #(
		.INIT('h1)
	) name3098 (
		_w1700_,
		_w2093_,
		_w3630_
	);
	LUT2 #(
		.INIT('h1)
	) name3099 (
		_w2119_,
		_w3599_,
		_w3631_
	);
	LUT2 #(
		.INIT('h8)
	) name3100 (
		_w3630_,
		_w3631_,
		_w3632_
	);
	LUT2 #(
		.INIT('h1)
	) name3101 (
		\sa10_reg[2]/P0001 ,
		_w3632_,
		_w3633_
	);
	LUT2 #(
		.INIT('h2)
	) name3102 (
		_w2565_,
		_w2595_,
		_w3634_
	);
	LUT2 #(
		.INIT('h8)
	) name3103 (
		\sa10_reg[4]/P0001 ,
		_w1616_,
		_w3635_
	);
	LUT2 #(
		.INIT('h1)
	) name3104 (
		_w3634_,
		_w3635_,
		_w3636_
	);
	LUT2 #(
		.INIT('h4)
	) name3105 (
		_w3629_,
		_w3636_,
		_w3637_
	);
	LUT2 #(
		.INIT('h4)
	) name3106 (
		_w3633_,
		_w3637_,
		_w3638_
	);
	LUT2 #(
		.INIT('h4)
	) name3107 (
		_w3622_,
		_w3638_,
		_w3639_
	);
	LUT2 #(
		.INIT('h2)
	) name3108 (
		\sa10_reg[0]/P0001 ,
		_w3639_,
		_w3640_
	);
	LUT2 #(
		.INIT('h4)
	) name3109 (
		\sa10_reg[6]/NET0131 ,
		_w1590_,
		_w3641_
	);
	LUT2 #(
		.INIT('h2)
	) name3110 (
		_w1634_,
		_w3616_,
		_w3642_
	);
	LUT2 #(
		.INIT('h1)
	) name3111 (
		_w3641_,
		_w3642_,
		_w3643_
	);
	LUT2 #(
		.INIT('h1)
	) name3112 (
		\sa10_reg[2]/P0001 ,
		_w3643_,
		_w3644_
	);
	LUT2 #(
		.INIT('h1)
	) name3113 (
		_w1591_,
		_w1684_,
		_w3645_
	);
	LUT2 #(
		.INIT('h2)
	) name3114 (
		\sa10_reg[2]/P0001 ,
		_w3645_,
		_w3646_
	);
	LUT2 #(
		.INIT('h4)
	) name3115 (
		_w2185_,
		_w2744_,
		_w3647_
	);
	LUT2 #(
		.INIT('h4)
	) name3116 (
		_w3646_,
		_w3647_,
		_w3648_
	);
	LUT2 #(
		.INIT('h4)
	) name3117 (
		_w3644_,
		_w3648_,
		_w3649_
	);
	LUT2 #(
		.INIT('h2)
	) name3118 (
		\sa10_reg[1]/P0001 ,
		_w3649_,
		_w3650_
	);
	LUT2 #(
		.INIT('h1)
	) name3119 (
		_w1586_,
		_w1687_,
		_w3651_
	);
	LUT2 #(
		.INIT('h2)
	) name3120 (
		_w1661_,
		_w3651_,
		_w3652_
	);
	LUT2 #(
		.INIT('h1)
	) name3121 (
		_w2567_,
		_w2748_,
		_w3653_
	);
	LUT2 #(
		.INIT('h1)
	) name3122 (
		\sa10_reg[2]/P0001 ,
		_w3653_,
		_w3654_
	);
	LUT2 #(
		.INIT('h1)
	) name3123 (
		_w1730_,
		_w2807_,
		_w3655_
	);
	LUT2 #(
		.INIT('h4)
	) name3124 (
		_w3652_,
		_w3655_,
		_w3656_
	);
	LUT2 #(
		.INIT('h4)
	) name3125 (
		_w3654_,
		_w3656_,
		_w3657_
	);
	LUT2 #(
		.INIT('h4)
	) name3126 (
		_w3650_,
		_w3657_,
		_w3658_
	);
	LUT2 #(
		.INIT('h1)
	) name3127 (
		\sa10_reg[0]/P0001 ,
		_w3658_,
		_w3659_
	);
	LUT2 #(
		.INIT('h8)
	) name3128 (
		_w1582_,
		_w1668_,
		_w3660_
	);
	LUT2 #(
		.INIT('h1)
	) name3129 (
		_w1587_,
		_w2185_,
		_w3661_
	);
	LUT2 #(
		.INIT('h4)
	) name3130 (
		_w3660_,
		_w3661_,
		_w3662_
	);
	LUT2 #(
		.INIT('h1)
	) name3131 (
		_w1602_,
		_w1616_,
		_w3663_
	);
	LUT2 #(
		.INIT('h8)
	) name3132 (
		_w3662_,
		_w3663_,
		_w3664_
	);
	LUT2 #(
		.INIT('h2)
	) name3133 (
		\sa10_reg[1]/P0001 ,
		_w3664_,
		_w3665_
	);
	LUT2 #(
		.INIT('h1)
	) name3134 (
		\sa10_reg[2]/P0001 ,
		_w3665_,
		_w3666_
	);
	LUT2 #(
		.INIT('h4)
	) name3135 (
		\sa10_reg[5]/P0001 ,
		_w3641_,
		_w3667_
	);
	LUT2 #(
		.INIT('h1)
	) name3136 (
		\sa10_reg[1]/P0001 ,
		_w1730_,
		_w3668_
	);
	LUT2 #(
		.INIT('h4)
	) name3137 (
		_w1592_,
		_w3668_,
		_w3669_
	);
	LUT2 #(
		.INIT('h4)
	) name3138 (
		_w3667_,
		_w3669_,
		_w3670_
	);
	LUT2 #(
		.INIT('h1)
	) name3139 (
		_w1609_,
		_w2546_,
		_w3671_
	);
	LUT2 #(
		.INIT('h2)
	) name3140 (
		\sa10_reg[3]/P0001 ,
		_w3671_,
		_w3672_
	);
	LUT2 #(
		.INIT('h4)
	) name3141 (
		_w1674_,
		_w1697_,
		_w3673_
	);
	LUT2 #(
		.INIT('h4)
	) name3142 (
		_w3672_,
		_w3673_,
		_w3674_
	);
	LUT2 #(
		.INIT('h1)
	) name3143 (
		_w3670_,
		_w3674_,
		_w3675_
	);
	LUT2 #(
		.INIT('h1)
	) name3144 (
		_w2558_,
		_w2819_,
		_w3676_
	);
	LUT2 #(
		.INIT('h4)
	) name3145 (
		_w3675_,
		_w3676_,
		_w3677_
	);
	LUT2 #(
		.INIT('h1)
	) name3146 (
		_w3666_,
		_w3677_,
		_w3678_
	);
	LUT2 #(
		.INIT('h1)
	) name3147 (
		_w3659_,
		_w3678_,
		_w3679_
	);
	LUT2 #(
		.INIT('h4)
	) name3148 (
		_w3612_,
		_w3679_,
		_w3680_
	);
	LUT2 #(
		.INIT('h4)
	) name3149 (
		_w3640_,
		_w3680_,
		_w3681_
	);
	LUT2 #(
		.INIT('h1)
	) name3150 (
		_w1462_,
		_w2685_,
		_w3682_
	);
	LUT2 #(
		.INIT('h1)
	) name3151 (
		\sa03_reg[2]/P0001 ,
		_w3682_,
		_w3683_
	);
	LUT2 #(
		.INIT('h1)
	) name3152 (
		_w1537_,
		_w2289_,
		_w3684_
	);
	LUT2 #(
		.INIT('h2)
	) name3153 (
		_w1494_,
		_w3684_,
		_w3685_
	);
	LUT2 #(
		.INIT('h8)
	) name3154 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[2]/P0001 ,
		_w3686_
	);
	LUT2 #(
		.INIT('h8)
	) name3155 (
		_w1327_,
		_w1342_,
		_w3687_
	);
	LUT2 #(
		.INIT('h1)
	) name3156 (
		_w1375_,
		_w3687_,
		_w3688_
	);
	LUT2 #(
		.INIT('h2)
	) name3157 (
		_w3686_,
		_w3688_,
		_w3689_
	);
	LUT2 #(
		.INIT('h1)
	) name3158 (
		_w1383_,
		_w1460_,
		_w3690_
	);
	LUT2 #(
		.INIT('h2)
	) name3159 (
		_w1436_,
		_w3690_,
		_w3691_
	);
	LUT2 #(
		.INIT('h8)
	) name3160 (
		\sa03_reg[7]/NET0131 ,
		_w1408_,
		_w3692_
	);
	LUT2 #(
		.INIT('h1)
	) name3161 (
		_w1455_,
		_w2248_,
		_w3693_
	);
	LUT2 #(
		.INIT('h4)
	) name3162 (
		_w3692_,
		_w3693_,
		_w3694_
	);
	LUT2 #(
		.INIT('h1)
	) name3163 (
		\sa03_reg[2]/P0001 ,
		_w3694_,
		_w3695_
	);
	LUT2 #(
		.INIT('h4)
	) name3164 (
		_w1325_,
		_w1448_,
		_w3696_
	);
	LUT2 #(
		.INIT('h4)
	) name3165 (
		_w3695_,
		_w3696_,
		_w3697_
	);
	LUT2 #(
		.INIT('h2)
	) name3166 (
		\sa03_reg[1]/P0001 ,
		_w3697_,
		_w3698_
	);
	LUT2 #(
		.INIT('h1)
	) name3167 (
		_w1483_,
		_w1566_,
		_w3699_
	);
	LUT2 #(
		.INIT('h1)
	) name3168 (
		\sa03_reg[2]/P0001 ,
		_w3699_,
		_w3700_
	);
	LUT2 #(
		.INIT('h1)
	) name3169 (
		_w1552_,
		_w2685_,
		_w3701_
	);
	LUT2 #(
		.INIT('h4)
	) name3170 (
		_w3700_,
		_w3701_,
		_w3702_
	);
	LUT2 #(
		.INIT('h1)
	) name3171 (
		\sa03_reg[1]/P0001 ,
		_w3702_,
		_w3703_
	);
	LUT2 #(
		.INIT('h1)
	) name3172 (
		_w1409_,
		_w1415_,
		_w3704_
	);
	LUT2 #(
		.INIT('h4)
	) name3173 (
		_w3689_,
		_w3704_,
		_w3705_
	);
	LUT2 #(
		.INIT('h4)
	) name3174 (
		_w3691_,
		_w3705_,
		_w3706_
	);
	LUT2 #(
		.INIT('h1)
	) name3175 (
		_w3683_,
		_w3685_,
		_w3707_
	);
	LUT2 #(
		.INIT('h8)
	) name3176 (
		_w3706_,
		_w3707_,
		_w3708_
	);
	LUT2 #(
		.INIT('h4)
	) name3177 (
		_w3698_,
		_w3708_,
		_w3709_
	);
	LUT2 #(
		.INIT('h4)
	) name3178 (
		_w3703_,
		_w3709_,
		_w3710_
	);
	LUT2 #(
		.INIT('h1)
	) name3179 (
		\sa03_reg[0]/P0001 ,
		_w3710_,
		_w3711_
	);
	LUT2 #(
		.INIT('h8)
	) name3180 (
		_w1316_,
		_w1353_,
		_w3712_
	);
	LUT2 #(
		.INIT('h1)
	) name3181 (
		_w1369_,
		_w3712_,
		_w3713_
	);
	LUT2 #(
		.INIT('h8)
	) name3182 (
		\sa03_reg[3]/P0001 ,
		_w2684_,
		_w3714_
	);
	LUT2 #(
		.INIT('h1)
	) name3183 (
		_w1396_,
		_w2264_,
		_w3715_
	);
	LUT2 #(
		.INIT('h4)
	) name3184 (
		_w3714_,
		_w3715_,
		_w3716_
	);
	LUT2 #(
		.INIT('h2)
	) name3185 (
		\sa03_reg[2]/P0001 ,
		_w3716_,
		_w3717_
	);
	LUT2 #(
		.INIT('h2)
	) name3186 (
		_w3713_,
		_w3717_,
		_w3718_
	);
	LUT2 #(
		.INIT('h2)
	) name3187 (
		\sa03_reg[1]/P0001 ,
		_w3718_,
		_w3719_
	);
	LUT2 #(
		.INIT('h2)
	) name3188 (
		_w1316_,
		_w2684_,
		_w3720_
	);
	LUT2 #(
		.INIT('h4)
	) name3189 (
		_w1376_,
		_w3720_,
		_w3721_
	);
	LUT2 #(
		.INIT('h8)
	) name3190 (
		_w1332_,
		_w1429_,
		_w3722_
	);
	LUT2 #(
		.INIT('h1)
	) name3191 (
		_w3721_,
		_w3722_,
		_w3723_
	);
	LUT2 #(
		.INIT('h1)
	) name3192 (
		\sa03_reg[1]/P0001 ,
		_w3723_,
		_w3724_
	);
	LUT2 #(
		.INIT('h2)
	) name3193 (
		_w1328_,
		_w1515_,
		_w3725_
	);
	LUT2 #(
		.INIT('h4)
	) name3194 (
		\sa03_reg[3]/P0001 ,
		_w1329_,
		_w3726_
	);
	LUT2 #(
		.INIT('h4)
	) name3195 (
		\sa03_reg[1]/P0001 ,
		_w1330_,
		_w3727_
	);
	LUT2 #(
		.INIT('h1)
	) name3196 (
		_w1341_,
		_w3727_,
		_w3728_
	);
	LUT2 #(
		.INIT('h2)
	) name3197 (
		_w3726_,
		_w3728_,
		_w3729_
	);
	LUT2 #(
		.INIT('h2)
	) name3198 (
		_w2200_,
		_w3686_,
		_w3730_
	);
	LUT2 #(
		.INIT('h1)
	) name3199 (
		_w1414_,
		_w1565_,
		_w3731_
	);
	LUT2 #(
		.INIT('h4)
	) name3200 (
		_w2289_,
		_w3731_,
		_w3732_
	);
	LUT2 #(
		.INIT('h1)
	) name3201 (
		\sa03_reg[2]/P0001 ,
		_w3732_,
		_w3733_
	);
	LUT2 #(
		.INIT('h1)
	) name3202 (
		_w3725_,
		_w3730_,
		_w3734_
	);
	LUT2 #(
		.INIT('h4)
	) name3203 (
		_w3729_,
		_w3734_,
		_w3735_
	);
	LUT2 #(
		.INIT('h4)
	) name3204 (
		_w3724_,
		_w3735_,
		_w3736_
	);
	LUT2 #(
		.INIT('h4)
	) name3205 (
		_w3733_,
		_w3736_,
		_w3737_
	);
	LUT2 #(
		.INIT('h4)
	) name3206 (
		_w3719_,
		_w3737_,
		_w3738_
	);
	LUT2 #(
		.INIT('h2)
	) name3207 (
		\sa03_reg[0]/P0001 ,
		_w3738_,
		_w3739_
	);
	LUT2 #(
		.INIT('h1)
	) name3208 (
		_w1359_,
		_w1409_,
		_w3740_
	);
	LUT2 #(
		.INIT('h4)
	) name3209 (
		_w1438_,
		_w3740_,
		_w3741_
	);
	LUT2 #(
		.INIT('h2)
	) name3210 (
		\sa03_reg[2]/P0001 ,
		_w3741_,
		_w3742_
	);
	LUT2 #(
		.INIT('h1)
	) name3211 (
		_w1459_,
		_w2679_,
		_w3743_
	);
	LUT2 #(
		.INIT('h4)
	) name3212 (
		_w3742_,
		_w3743_,
		_w3744_
	);
	LUT2 #(
		.INIT('h1)
	) name3213 (
		\sa03_reg[1]/P0001 ,
		_w3744_,
		_w3745_
	);
	LUT2 #(
		.INIT('h4)
	) name3214 (
		_w1334_,
		_w1355_,
		_w3746_
	);
	LUT2 #(
		.INIT('h1)
	) name3215 (
		_w3726_,
		_w3746_,
		_w3747_
	);
	LUT2 #(
		.INIT('h1)
	) name3216 (
		\sa03_reg[7]/NET0131 ,
		_w3747_,
		_w3748_
	);
	LUT2 #(
		.INIT('h4)
	) name3217 (
		\sa03_reg[4]/P0001 ,
		_w3726_,
		_w3749_
	);
	LUT2 #(
		.INIT('h1)
	) name3218 (
		_w1497_,
		_w3749_,
		_w3750_
	);
	LUT2 #(
		.INIT('h4)
	) name3219 (
		_w3748_,
		_w3750_,
		_w3751_
	);
	LUT2 #(
		.INIT('h2)
	) name3220 (
		_w1558_,
		_w3751_,
		_w3752_
	);
	LUT2 #(
		.INIT('h1)
	) name3221 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[2]/P0001 ,
		_w3753_
	);
	LUT2 #(
		.INIT('h1)
	) name3222 (
		_w1480_,
		_w2219_,
		_w3754_
	);
	LUT2 #(
		.INIT('h4)
	) name3223 (
		_w1461_,
		_w3754_,
		_w3755_
	);
	LUT2 #(
		.INIT('h2)
	) name3224 (
		_w3753_,
		_w3755_,
		_w3756_
	);
	LUT2 #(
		.INIT('h1)
	) name3225 (
		_w1369_,
		_w2260_,
		_w3757_
	);
	LUT2 #(
		.INIT('h2)
	) name3226 (
		\sa03_reg[3]/P0001 ,
		_w3757_,
		_w3758_
	);
	LUT2 #(
		.INIT('h1)
	) name3227 (
		_w1526_,
		_w3758_,
		_w3759_
	);
	LUT2 #(
		.INIT('h2)
	) name3228 (
		_w3686_,
		_w3759_,
		_w3760_
	);
	LUT2 #(
		.INIT('h8)
	) name3229 (
		_w1384_,
		_w2229_,
		_w3761_
	);
	LUT2 #(
		.INIT('h1)
	) name3230 (
		_w2235_,
		_w3761_,
		_w3762_
	);
	LUT2 #(
		.INIT('h4)
	) name3231 (
		_w3756_,
		_w3762_,
		_w3763_
	);
	LUT2 #(
		.INIT('h4)
	) name3232 (
		_w3752_,
		_w3763_,
		_w3764_
	);
	LUT2 #(
		.INIT('h4)
	) name3233 (
		_w3760_,
		_w3764_,
		_w3765_
	);
	LUT2 #(
		.INIT('h4)
	) name3234 (
		_w3745_,
		_w3765_,
		_w3766_
	);
	LUT2 #(
		.INIT('h4)
	) name3235 (
		_w3739_,
		_w3766_,
		_w3767_
	);
	LUT2 #(
		.INIT('h4)
	) name3236 (
		_w3711_,
		_w3767_,
		_w3768_
	);
	LUT2 #(
		.INIT('h1)
	) name3237 (
		_w3681_,
		_w3768_,
		_w3769_
	);
	LUT2 #(
		.INIT('h8)
	) name3238 (
		_w3681_,
		_w3768_,
		_w3770_
	);
	LUT2 #(
		.INIT('h1)
	) name3239 (
		_w3769_,
		_w3770_,
		_w3771_
	);
	LUT2 #(
		.INIT('h8)
	) name3240 (
		_w3595_,
		_w3771_,
		_w3772_
	);
	LUT2 #(
		.INIT('h1)
	) name3241 (
		_w3595_,
		_w3771_,
		_w3773_
	);
	LUT2 #(
		.INIT('h1)
	) name3242 (
		_w3772_,
		_w3773_,
		_w3774_
	);
	LUT2 #(
		.INIT('h1)
	) name3243 (
		_w3509_,
		_w3774_,
		_w3775_
	);
	LUT2 #(
		.INIT('h8)
	) name3244 (
		_w3509_,
		_w3774_,
		_w3776_
	);
	LUT2 #(
		.INIT('h1)
	) name3245 (
		\ld_r_reg/P0001 ,
		_w3775_,
		_w3777_
	);
	LUT2 #(
		.INIT('h4)
	) name3246 (
		_w3776_,
		_w3777_,
		_w3778_
	);
	LUT2 #(
		.INIT('h1)
	) name3247 (
		\text_in_r_reg[9]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w3779_
	);
	LUT2 #(
		.INIT('h8)
	) name3248 (
		\text_in_r_reg[9]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w3780_
	);
	LUT2 #(
		.INIT('h2)
	) name3249 (
		\ld_r_reg/P0001 ,
		_w3779_,
		_w3781_
	);
	LUT2 #(
		.INIT('h4)
	) name3250 (
		_w3780_,
		_w3781_,
		_w3782_
	);
	LUT2 #(
		.INIT('h1)
	) name3251 (
		_w3778_,
		_w3782_,
		_w3783_
	);
	LUT2 #(
		.INIT('h1)
	) name3252 (
		_w2736_,
		_w2963_,
		_w3784_
	);
	LUT2 #(
		.INIT('h8)
	) name3253 (
		_w2736_,
		_w2963_,
		_w3785_
	);
	LUT2 #(
		.INIT('h1)
	) name3254 (
		_w3784_,
		_w3785_,
		_w3786_
	);
	LUT2 #(
		.INIT('h2)
	) name3255 (
		\u0_w_reg[3][5]/P0001 ,
		_w3205_,
		_w3787_
	);
	LUT2 #(
		.INIT('h4)
	) name3256 (
		\u0_w_reg[3][5]/P0001 ,
		_w3205_,
		_w3788_
	);
	LUT2 #(
		.INIT('h1)
	) name3257 (
		_w3787_,
		_w3788_,
		_w3789_
	);
	LUT2 #(
		.INIT('h8)
	) name3258 (
		_w2939_,
		_w3789_,
		_w3790_
	);
	LUT2 #(
		.INIT('h1)
	) name3259 (
		_w2939_,
		_w3789_,
		_w3791_
	);
	LUT2 #(
		.INIT('h1)
	) name3260 (
		_w3790_,
		_w3791_,
		_w3792_
	);
	LUT2 #(
		.INIT('h1)
	) name3261 (
		_w3786_,
		_w3792_,
		_w3793_
	);
	LUT2 #(
		.INIT('h8)
	) name3262 (
		_w3786_,
		_w3792_,
		_w3794_
	);
	LUT2 #(
		.INIT('h1)
	) name3263 (
		\ld_r_reg/P0001 ,
		_w3793_,
		_w3795_
	);
	LUT2 #(
		.INIT('h4)
	) name3264 (
		_w3794_,
		_w3795_,
		_w3796_
	);
	LUT2 #(
		.INIT('h1)
	) name3265 (
		\text_in_r_reg[5]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		_w3797_
	);
	LUT2 #(
		.INIT('h8)
	) name3266 (
		\text_in_r_reg[5]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		_w3798_
	);
	LUT2 #(
		.INIT('h2)
	) name3267 (
		\ld_r_reg/P0001 ,
		_w3797_,
		_w3799_
	);
	LUT2 #(
		.INIT('h4)
	) name3268 (
		_w3798_,
		_w3799_,
		_w3800_
	);
	LUT2 #(
		.INIT('h1)
	) name3269 (
		_w3796_,
		_w3800_,
		_w3801_
	);
	LUT2 #(
		.INIT('h2)
	) name3270 (
		\u0_w_reg[3][28]/P0001 ,
		_w3205_,
		_w3802_
	);
	LUT2 #(
		.INIT('h4)
	) name3271 (
		\u0_w_reg[3][28]/P0001 ,
		_w3205_,
		_w3803_
	);
	LUT2 #(
		.INIT('h1)
	) name3272 (
		_w3802_,
		_w3803_,
		_w3804_
	);
	LUT2 #(
		.INIT('h8)
	) name3273 (
		_w3072_,
		_w3804_,
		_w3805_
	);
	LUT2 #(
		.INIT('h1)
	) name3274 (
		_w3072_,
		_w3804_,
		_w3806_
	);
	LUT2 #(
		.INIT('h1)
	) name3275 (
		_w3805_,
		_w3806_,
		_w3807_
	);
	LUT2 #(
		.INIT('h1)
	) name3276 (
		_w1328_,
		_w2219_,
		_w3808_
	);
	LUT2 #(
		.INIT('h1)
	) name3277 (
		\sa03_reg[2]/P0001 ,
		_w3808_,
		_w3809_
	);
	LUT2 #(
		.INIT('h8)
	) name3278 (
		\sa03_reg[2]/P0001 ,
		_w1450_,
		_w3810_
	);
	LUT2 #(
		.INIT('h1)
	) name3279 (
		_w1409_,
		_w1571_,
		_w3811_
	);
	LUT2 #(
		.INIT('h4)
	) name3280 (
		_w1496_,
		_w3811_,
		_w3812_
	);
	LUT2 #(
		.INIT('h1)
	) name3281 (
		_w2679_,
		_w2715_,
		_w3813_
	);
	LUT2 #(
		.INIT('h4)
	) name3282 (
		_w3810_,
		_w3813_,
		_w3814_
	);
	LUT2 #(
		.INIT('h4)
	) name3283 (
		_w3809_,
		_w3812_,
		_w3815_
	);
	LUT2 #(
		.INIT('h8)
	) name3284 (
		_w3814_,
		_w3815_,
		_w3816_
	);
	LUT2 #(
		.INIT('h1)
	) name3285 (
		\sa03_reg[1]/P0001 ,
		_w3816_,
		_w3817_
	);
	LUT2 #(
		.INIT('h1)
	) name3286 (
		_w1329_,
		_w1398_,
		_w3818_
	);
	LUT2 #(
		.INIT('h4)
	) name3287 (
		\sa03_reg[7]/NET0131 ,
		_w3818_,
		_w3819_
	);
	LUT2 #(
		.INIT('h1)
	) name3288 (
		\sa03_reg[2]/P0001 ,
		_w3819_,
		_w3820_
	);
	LUT2 #(
		.INIT('h8)
	) name3289 (
		\sa03_reg[4]/P0001 ,
		_w1367_,
		_w3821_
	);
	LUT2 #(
		.INIT('h2)
	) name3290 (
		\sa03_reg[2]/P0001 ,
		_w2710_,
		_w3822_
	);
	LUT2 #(
		.INIT('h1)
	) name3291 (
		_w3726_,
		_w3821_,
		_w3823_
	);
	LUT2 #(
		.INIT('h8)
	) name3292 (
		_w3822_,
		_w3823_,
		_w3824_
	);
	LUT2 #(
		.INIT('h1)
	) name3293 (
		_w3820_,
		_w3824_,
		_w3825_
	);
	LUT2 #(
		.INIT('h1)
	) name3294 (
		_w1537_,
		_w2293_,
		_w3826_
	);
	LUT2 #(
		.INIT('h4)
	) name3295 (
		_w1365_,
		_w3826_,
		_w3827_
	);
	LUT2 #(
		.INIT('h4)
	) name3296 (
		_w3825_,
		_w3827_,
		_w3828_
	);
	LUT2 #(
		.INIT('h2)
	) name3297 (
		\sa03_reg[1]/P0001 ,
		_w3828_,
		_w3829_
	);
	LUT2 #(
		.INIT('h4)
	) name3298 (
		\sa03_reg[3]/P0001 ,
		_w1330_,
		_w3830_
	);
	LUT2 #(
		.INIT('h4)
	) name3299 (
		\sa03_reg[5]/P0001 ,
		_w3830_,
		_w3831_
	);
	LUT2 #(
		.INIT('h8)
	) name3300 (
		\sa03_reg[6]/NET0131 ,
		_w1340_,
		_w3832_
	);
	LUT2 #(
		.INIT('h1)
	) name3301 (
		_w1462_,
		_w3832_,
		_w3833_
	);
	LUT2 #(
		.INIT('h4)
	) name3302 (
		_w3831_,
		_w3833_,
		_w3834_
	);
	LUT2 #(
		.INIT('h1)
	) name3303 (
		\sa03_reg[2]/P0001 ,
		_w3834_,
		_w3835_
	);
	LUT2 #(
		.INIT('h4)
	) name3304 (
		_w1333_,
		_w1405_,
		_w3836_
	);
	LUT2 #(
		.INIT('h8)
	) name3305 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w3837_
	);
	LUT2 #(
		.INIT('h4)
	) name3306 (
		_w3836_,
		_w3837_,
		_w3838_
	);
	LUT2 #(
		.INIT('h1)
	) name3307 (
		_w1469_,
		_w3838_,
		_w3839_
	);
	LUT2 #(
		.INIT('h4)
	) name3308 (
		_w3835_,
		_w3839_,
		_w3840_
	);
	LUT2 #(
		.INIT('h4)
	) name3309 (
		_w3817_,
		_w3840_,
		_w3841_
	);
	LUT2 #(
		.INIT('h4)
	) name3310 (
		_w3829_,
		_w3841_,
		_w3842_
	);
	LUT2 #(
		.INIT('h2)
	) name3311 (
		\sa03_reg[0]/P0001 ,
		_w3842_,
		_w3843_
	);
	LUT2 #(
		.INIT('h8)
	) name3312 (
		_w1369_,
		_w1374_,
		_w3844_
	);
	LUT2 #(
		.INIT('h4)
	) name3313 (
		\sa03_reg[2]/P0001 ,
		_w2693_,
		_w3845_
	);
	LUT2 #(
		.INIT('h1)
	) name3314 (
		_w1319_,
		_w1331_,
		_w3846_
	);
	LUT2 #(
		.INIT('h4)
	) name3315 (
		_w1533_,
		_w3846_,
		_w3847_
	);
	LUT2 #(
		.INIT('h2)
	) name3316 (
		_w2225_,
		_w3847_,
		_w3848_
	);
	LUT2 #(
		.INIT('h1)
	) name3317 (
		_w2658_,
		_w3845_,
		_w3849_
	);
	LUT2 #(
		.INIT('h4)
	) name3318 (
		_w3848_,
		_w3849_,
		_w3850_
	);
	LUT2 #(
		.INIT('h2)
	) name3319 (
		\sa03_reg[1]/P0001 ,
		_w3850_,
		_w3851_
	);
	LUT2 #(
		.INIT('h8)
	) name3320 (
		\sa03_reg[6]/NET0131 ,
		_w1454_,
		_w3852_
	);
	LUT2 #(
		.INIT('h1)
	) name3321 (
		_w1537_,
		_w3852_,
		_w3853_
	);
	LUT2 #(
		.INIT('h2)
	) name3322 (
		_w3686_,
		_w3853_,
		_w3854_
	);
	LUT2 #(
		.INIT('h1)
	) name3323 (
		_w1443_,
		_w1461_,
		_w3855_
	);
	LUT2 #(
		.INIT('h2)
	) name3324 (
		_w1494_,
		_w3855_,
		_w3856_
	);
	LUT2 #(
		.INIT('h8)
	) name3325 (
		_w2655_,
		_w3753_,
		_w3857_
	);
	LUT2 #(
		.INIT('h4)
	) name3326 (
		\sa03_reg[2]/P0001 ,
		_w1489_,
		_w3858_
	);
	LUT2 #(
		.INIT('h8)
	) name3327 (
		_w1324_,
		_w1383_,
		_w3859_
	);
	LUT2 #(
		.INIT('h2)
	) name3328 (
		_w1562_,
		_w3859_,
		_w3860_
	);
	LUT2 #(
		.INIT('h1)
	) name3329 (
		_w3858_,
		_w3860_,
		_w3861_
	);
	LUT2 #(
		.INIT('h1)
	) name3330 (
		_w1377_,
		_w1421_,
		_w3862_
	);
	LUT2 #(
		.INIT('h2)
	) name3331 (
		\sa03_reg[2]/P0001 ,
		_w3862_,
		_w3863_
	);
	LUT2 #(
		.INIT('h4)
	) name3332 (
		\sa03_reg[2]/P0001 ,
		_w1331_,
		_w3864_
	);
	LUT2 #(
		.INIT('h2)
	) name3333 (
		\sa03_reg[1]/P0001 ,
		_w2665_,
		_w3865_
	);
	LUT2 #(
		.INIT('h4)
	) name3334 (
		_w1354_,
		_w3865_,
		_w3866_
	);
	LUT2 #(
		.INIT('h1)
	) name3335 (
		_w3712_,
		_w3864_,
		_w3867_
	);
	LUT2 #(
		.INIT('h8)
	) name3336 (
		_w3866_,
		_w3867_,
		_w3868_
	);
	LUT2 #(
		.INIT('h4)
	) name3337 (
		_w3863_,
		_w3868_,
		_w3869_
	);
	LUT2 #(
		.INIT('h2)
	) name3338 (
		_w1341_,
		_w1385_,
		_w3870_
	);
	LUT2 #(
		.INIT('h2)
	) name3339 (
		\sa03_reg[2]/P0001 ,
		_w1355_,
		_w3871_
	);
	LUT2 #(
		.INIT('h8)
	) name3340 (
		_w1327_,
		_w3871_,
		_w3872_
	);
	LUT2 #(
		.INIT('h1)
	) name3341 (
		\sa03_reg[1]/P0001 ,
		_w3831_,
		_w3873_
	);
	LUT2 #(
		.INIT('h1)
	) name3342 (
		_w3870_,
		_w3872_,
		_w3874_
	);
	LUT2 #(
		.INIT('h8)
	) name3343 (
		_w3873_,
		_w3874_,
		_w3875_
	);
	LUT2 #(
		.INIT('h4)
	) name3344 (
		_w1560_,
		_w3875_,
		_w3876_
	);
	LUT2 #(
		.INIT('h1)
	) name3345 (
		_w3869_,
		_w3876_,
		_w3877_
	);
	LUT2 #(
		.INIT('h1)
	) name3346 (
		_w1443_,
		_w3861_,
		_w3878_
	);
	LUT2 #(
		.INIT('h4)
	) name3347 (
		_w3877_,
		_w3878_,
		_w3879_
	);
	LUT2 #(
		.INIT('h1)
	) name3348 (
		\sa03_reg[0]/P0001 ,
		_w3879_,
		_w3880_
	);
	LUT2 #(
		.INIT('h1)
	) name3349 (
		_w1552_,
		_w3761_,
		_w3881_
	);
	LUT2 #(
		.INIT('h1)
	) name3350 (
		_w3844_,
		_w3857_,
		_w3882_
	);
	LUT2 #(
		.INIT('h8)
	) name3351 (
		_w3881_,
		_w3882_,
		_w3883_
	);
	LUT2 #(
		.INIT('h4)
	) name3352 (
		_w3854_,
		_w3883_,
		_w3884_
	);
	LUT2 #(
		.INIT('h4)
	) name3353 (
		_w3856_,
		_w3884_,
		_w3885_
	);
	LUT2 #(
		.INIT('h4)
	) name3354 (
		_w3851_,
		_w3885_,
		_w3886_
	);
	LUT2 #(
		.INIT('h4)
	) name3355 (
		_w3880_,
		_w3886_,
		_w3887_
	);
	LUT2 #(
		.INIT('h4)
	) name3356 (
		_w3843_,
		_w3887_,
		_w3888_
	);
	LUT2 #(
		.INIT('h1)
	) name3357 (
		_w1601_,
		_w1657_,
		_w3889_
	);
	LUT2 #(
		.INIT('h2)
	) name3358 (
		\sa10_reg[2]/P0001 ,
		_w3889_,
		_w3890_
	);
	LUT2 #(
		.INIT('h8)
	) name3359 (
		_w1582_,
		_w2109_,
		_w3891_
	);
	LUT2 #(
		.INIT('h1)
	) name3360 (
		_w1599_,
		_w2550_,
		_w3892_
	);
	LUT2 #(
		.INIT('h1)
	) name3361 (
		_w3613_,
		_w3891_,
		_w3893_
	);
	LUT2 #(
		.INIT('h8)
	) name3362 (
		_w3892_,
		_w3893_,
		_w3894_
	);
	LUT2 #(
		.INIT('h4)
	) name3363 (
		_w3890_,
		_w3894_,
		_w3895_
	);
	LUT2 #(
		.INIT('h2)
	) name3364 (
		\sa10_reg[1]/P0001 ,
		_w3895_,
		_w3896_
	);
	LUT2 #(
		.INIT('h8)
	) name3365 (
		_w1601_,
		_w1664_,
		_w3897_
	);
	LUT2 #(
		.INIT('h1)
	) name3366 (
		\sa10_reg[2]/P0001 ,
		_w1596_,
		_w3898_
	);
	LUT2 #(
		.INIT('h2)
	) name3367 (
		_w1590_,
		_w1650_,
		_w3899_
	);
	LUT2 #(
		.INIT('h1)
	) name3368 (
		_w1703_,
		_w3899_,
		_w3900_
	);
	LUT2 #(
		.INIT('h2)
	) name3369 (
		\sa10_reg[2]/P0001 ,
		_w3900_,
		_w3901_
	);
	LUT2 #(
		.INIT('h8)
	) name3370 (
		_w1608_,
		_w1668_,
		_w3902_
	);
	LUT2 #(
		.INIT('h1)
	) name3371 (
		_w1704_,
		_w3902_,
		_w3903_
	);
	LUT2 #(
		.INIT('h4)
	) name3372 (
		_w1725_,
		_w3903_,
		_w3904_
	);
	LUT2 #(
		.INIT('h4)
	) name3373 (
		_w3901_,
		_w3904_,
		_w3905_
	);
	LUT2 #(
		.INIT('h1)
	) name3374 (
		\sa10_reg[1]/P0001 ,
		_w3905_,
		_w3906_
	);
	LUT2 #(
		.INIT('h1)
	) name3375 (
		_w1714_,
		_w2755_,
		_w3907_
	);
	LUT2 #(
		.INIT('h4)
	) name3376 (
		_w3897_,
		_w3907_,
		_w3908_
	);
	LUT2 #(
		.INIT('h4)
	) name3377 (
		_w3898_,
		_w3908_,
		_w3909_
	);
	LUT2 #(
		.INIT('h4)
	) name3378 (
		_w3896_,
		_w3909_,
		_w3910_
	);
	LUT2 #(
		.INIT('h4)
	) name3379 (
		_w3906_,
		_w3910_,
		_w3911_
	);
	LUT2 #(
		.INIT('h1)
	) name3380 (
		\sa10_reg[0]/P0001 ,
		_w3911_,
		_w3912_
	);
	LUT2 #(
		.INIT('h8)
	) name3381 (
		_w1609_,
		_w1664_,
		_w3913_
	);
	LUT2 #(
		.INIT('h8)
	) name3382 (
		\sa10_reg[6]/NET0131 ,
		_w1726_,
		_w3914_
	);
	LUT2 #(
		.INIT('h1)
	) name3383 (
		_w2607_,
		_w3914_,
		_w3915_
	);
	LUT2 #(
		.INIT('h2)
	) name3384 (
		\sa10_reg[1]/P0001 ,
		_w3915_,
		_w3916_
	);
	LUT2 #(
		.INIT('h1)
	) name3385 (
		_w2558_,
		_w3916_,
		_w3917_
	);
	LUT2 #(
		.INIT('h2)
	) name3386 (
		\sa10_reg[2]/P0001 ,
		_w3917_,
		_w3918_
	);
	LUT2 #(
		.INIT('h1)
	) name3387 (
		_w1638_,
		_w2098_,
		_w3919_
	);
	LUT2 #(
		.INIT('h4)
	) name3388 (
		_w2582_,
		_w3919_,
		_w3920_
	);
	LUT2 #(
		.INIT('h2)
	) name3389 (
		_w1633_,
		_w3920_,
		_w3921_
	);
	LUT2 #(
		.INIT('h8)
	) name3390 (
		\sa10_reg[3]/P0001 ,
		_w1650_,
		_w3922_
	);
	LUT2 #(
		.INIT('h8)
	) name3391 (
		_w2109_,
		_w3922_,
		_w3923_
	);
	LUT2 #(
		.INIT('h1)
	) name3392 (
		_w2594_,
		_w3923_,
		_w3924_
	);
	LUT2 #(
		.INIT('h4)
	) name3393 (
		_w3921_,
		_w3924_,
		_w3925_
	);
	LUT2 #(
		.INIT('h2)
	) name3394 (
		\sa10_reg[1]/P0001 ,
		_w3925_,
		_w3926_
	);
	LUT2 #(
		.INIT('h1)
	) name3395 (
		_w2581_,
		_w2755_,
		_w3927_
	);
	LUT2 #(
		.INIT('h2)
	) name3396 (
		_w2183_,
		_w3927_,
		_w3928_
	);
	LUT2 #(
		.INIT('h8)
	) name3397 (
		_w2566_,
		_w2825_,
		_w3929_
	);
	LUT2 #(
		.INIT('h8)
	) name3398 (
		_w1626_,
		_w3616_,
		_w3930_
	);
	LUT2 #(
		.INIT('h2)
	) name3399 (
		_w1582_,
		_w2162_,
		_w3931_
	);
	LUT2 #(
		.INIT('h1)
	) name3400 (
		_w2623_,
		_w3931_,
		_w3932_
	);
	LUT2 #(
		.INIT('h2)
	) name3401 (
		\sa10_reg[2]/P0001 ,
		_w3932_,
		_w3933_
	);
	LUT2 #(
		.INIT('h1)
	) name3402 (
		_w2147_,
		_w2607_,
		_w3934_
	);
	LUT2 #(
		.INIT('h4)
	) name3403 (
		_w1688_,
		_w3934_,
		_w3935_
	);
	LUT2 #(
		.INIT('h4)
	) name3404 (
		_w3930_,
		_w3935_,
		_w3936_
	);
	LUT2 #(
		.INIT('h4)
	) name3405 (
		_w3933_,
		_w3936_,
		_w3937_
	);
	LUT2 #(
		.INIT('h2)
	) name3406 (
		\sa10_reg[1]/P0001 ,
		_w3937_,
		_w3938_
	);
	LUT2 #(
		.INIT('h8)
	) name3407 (
		\sa10_reg[6]/NET0131 ,
		_w2593_,
		_w3939_
	);
	LUT2 #(
		.INIT('h1)
	) name3408 (
		_w2748_,
		_w3939_,
		_w3940_
	);
	LUT2 #(
		.INIT('h4)
	) name3409 (
		_w3902_,
		_w3940_,
		_w3941_
	);
	LUT2 #(
		.INIT('h1)
	) name3410 (
		\sa10_reg[2]/P0001 ,
		_w3941_,
		_w3942_
	);
	LUT2 #(
		.INIT('h8)
	) name3411 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w3943_
	);
	LUT2 #(
		.INIT('h8)
	) name3412 (
		\sa10_reg[3]/P0001 ,
		_w1597_,
		_w3944_
	);
	LUT2 #(
		.INIT('h1)
	) name3413 (
		_w2811_,
		_w3944_,
		_w3945_
	);
	LUT2 #(
		.INIT('h2)
	) name3414 (
		_w3943_,
		_w3945_,
		_w3946_
	);
	LUT2 #(
		.INIT('h2)
	) name3415 (
		_w2131_,
		_w2565_,
		_w3947_
	);
	LUT2 #(
		.INIT('h1)
	) name3416 (
		_w2621_,
		_w2740_,
		_w3948_
	);
	LUT2 #(
		.INIT('h8)
	) name3417 (
		_w2602_,
		_w3948_,
		_w3949_
	);
	LUT2 #(
		.INIT('h1)
	) name3418 (
		_w3947_,
		_w3949_,
		_w3950_
	);
	LUT2 #(
		.INIT('h1)
	) name3419 (
		_w1711_,
		_w1730_,
		_w3951_
	);
	LUT2 #(
		.INIT('h4)
	) name3420 (
		_w2558_,
		_w3951_,
		_w3952_
	);
	LUT2 #(
		.INIT('h4)
	) name3421 (
		_w3950_,
		_w3952_,
		_w3953_
	);
	LUT2 #(
		.INIT('h1)
	) name3422 (
		\sa10_reg[1]/P0001 ,
		_w3953_,
		_w3954_
	);
	LUT2 #(
		.INIT('h1)
	) name3423 (
		_w2758_,
		_w3946_,
		_w3955_
	);
	LUT2 #(
		.INIT('h4)
	) name3424 (
		_w3942_,
		_w3955_,
		_w3956_
	);
	LUT2 #(
		.INIT('h4)
	) name3425 (
		_w3938_,
		_w3956_,
		_w3957_
	);
	LUT2 #(
		.INIT('h4)
	) name3426 (
		_w3954_,
		_w3957_,
		_w3958_
	);
	LUT2 #(
		.INIT('h2)
	) name3427 (
		\sa10_reg[0]/P0001 ,
		_w3958_,
		_w3959_
	);
	LUT2 #(
		.INIT('h1)
	) name3428 (
		_w3598_,
		_w3913_,
		_w3960_
	);
	LUT2 #(
		.INIT('h4)
	) name3429 (
		_w3929_,
		_w3960_,
		_w3961_
	);
	LUT2 #(
		.INIT('h4)
	) name3430 (
		_w3928_,
		_w3961_,
		_w3962_
	);
	LUT2 #(
		.INIT('h4)
	) name3431 (
		_w3918_,
		_w3962_,
		_w3963_
	);
	LUT2 #(
		.INIT('h4)
	) name3432 (
		_w3926_,
		_w3963_,
		_w3964_
	);
	LUT2 #(
		.INIT('h4)
	) name3433 (
		_w3912_,
		_w3964_,
		_w3965_
	);
	LUT2 #(
		.INIT('h4)
	) name3434 (
		_w3959_,
		_w3965_,
		_w3966_
	);
	LUT2 #(
		.INIT('h2)
	) name3435 (
		_w3888_,
		_w3966_,
		_w3967_
	);
	LUT2 #(
		.INIT('h4)
	) name3436 (
		_w3888_,
		_w3966_,
		_w3968_
	);
	LUT2 #(
		.INIT('h1)
	) name3437 (
		_w3967_,
		_w3968_,
		_w3969_
	);
	LUT2 #(
		.INIT('h4)
	) name3438 (
		_w2307_,
		_w3969_,
		_w3970_
	);
	LUT2 #(
		.INIT('h2)
	) name3439 (
		_w2307_,
		_w3969_,
		_w3971_
	);
	LUT2 #(
		.INIT('h1)
	) name3440 (
		_w3970_,
		_w3971_,
		_w3972_
	);
	LUT2 #(
		.INIT('h2)
	) name3441 (
		_w3807_,
		_w3972_,
		_w3973_
	);
	LUT2 #(
		.INIT('h4)
	) name3442 (
		_w3807_,
		_w3972_,
		_w3974_
	);
	LUT2 #(
		.INIT('h1)
	) name3443 (
		\ld_r_reg/P0001 ,
		_w3973_,
		_w3975_
	);
	LUT2 #(
		.INIT('h4)
	) name3444 (
		_w3974_,
		_w3975_,
		_w3976_
	);
	LUT2 #(
		.INIT('h2)
	) name3445 (
		\text_in_r_reg[28]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w3977_
	);
	LUT2 #(
		.INIT('h4)
	) name3446 (
		\text_in_r_reg[28]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w3978_
	);
	LUT2 #(
		.INIT('h2)
	) name3447 (
		\ld_r_reg/P0001 ,
		_w3977_,
		_w3979_
	);
	LUT2 #(
		.INIT('h4)
	) name3448 (
		_w3978_,
		_w3979_,
		_w3980_
	);
	LUT2 #(
		.INIT('h1)
	) name3449 (
		_w3976_,
		_w3980_,
		_w3981_
	);
	LUT2 #(
		.INIT('h8)
	) name3450 (
		_w1781_,
		_w1802_,
		_w3982_
	);
	LUT2 #(
		.INIT('h8)
	) name3451 (
		_w1764_,
		_w2479_,
		_w3983_
	);
	LUT2 #(
		.INIT('h1)
	) name3452 (
		_w1785_,
		_w1839_,
		_w3984_
	);
	LUT2 #(
		.INIT('h2)
	) name3453 (
		\sa21_reg[2]/P0001 ,
		_w3984_,
		_w3985_
	);
	LUT2 #(
		.INIT('h2)
	) name3454 (
		\sa21_reg[1]/P0001 ,
		_w1788_,
		_w3986_
	);
	LUT2 #(
		.INIT('h4)
	) name3455 (
		_w2853_,
		_w3986_,
		_w3987_
	);
	LUT2 #(
		.INIT('h1)
	) name3456 (
		_w3982_,
		_w3983_,
		_w3988_
	);
	LUT2 #(
		.INIT('h8)
	) name3457 (
		_w3987_,
		_w3988_,
		_w3989_
	);
	LUT2 #(
		.INIT('h4)
	) name3458 (
		_w3985_,
		_w3989_,
		_w3990_
	);
	LUT2 #(
		.INIT('h2)
	) name3459 (
		_w1757_,
		_w1832_,
		_w3991_
	);
	LUT2 #(
		.INIT('h1)
	) name3460 (
		_w2492_,
		_w3991_,
		_w3992_
	);
	LUT2 #(
		.INIT('h2)
	) name3461 (
		\sa21_reg[2]/P0001 ,
		_w3992_,
		_w3993_
	);
	LUT2 #(
		.INIT('h4)
	) name3462 (
		\sa21_reg[5]/P0001 ,
		_w1816_,
		_w3994_
	);
	LUT2 #(
		.INIT('h1)
	) name3463 (
		\sa21_reg[1]/P0001 ,
		_w1864_,
		_w3995_
	);
	LUT2 #(
		.INIT('h4)
	) name3464 (
		_w3994_,
		_w3995_,
		_w3996_
	);
	LUT2 #(
		.INIT('h1)
	) name3465 (
		_w1878_,
		_w3993_,
		_w3997_
	);
	LUT2 #(
		.INIT('h8)
	) name3466 (
		_w3996_,
		_w3997_,
		_w3998_
	);
	LUT2 #(
		.INIT('h1)
	) name3467 (
		_w3990_,
		_w3998_,
		_w3999_
	);
	LUT2 #(
		.INIT('h1)
	) name3468 (
		\sa21_reg[2]/P0001 ,
		_w1783_,
		_w4000_
	);
	LUT2 #(
		.INIT('h1)
	) name3469 (
		_w1890_,
		_w1895_,
		_w4001_
	);
	LUT2 #(
		.INIT('h2)
	) name3470 (
		_w1784_,
		_w4001_,
		_w4002_
	);
	LUT2 #(
		.INIT('h1)
	) name3471 (
		_w1893_,
		_w4002_,
		_w4003_
	);
	LUT2 #(
		.INIT('h4)
	) name3472 (
		_w4000_,
		_w4003_,
		_w4004_
	);
	LUT2 #(
		.INIT('h4)
	) name3473 (
		_w3999_,
		_w4004_,
		_w4005_
	);
	LUT2 #(
		.INIT('h1)
	) name3474 (
		\sa21_reg[0]/P0001 ,
		_w4005_,
		_w4006_
	);
	LUT2 #(
		.INIT('h8)
	) name3475 (
		\sa21_reg[2]/P0001 ,
		_w3040_,
		_w4007_
	);
	LUT2 #(
		.INIT('h1)
	) name3476 (
		_w1775_,
		_w1844_,
		_w4008_
	);
	LUT2 #(
		.INIT('h4)
	) name3477 (
		_w1765_,
		_w4008_,
		_w4009_
	);
	LUT2 #(
		.INIT('h2)
	) name3478 (
		_w1754_,
		_w4009_,
		_w4010_
	);
	LUT2 #(
		.INIT('h8)
	) name3479 (
		\sa21_reg[6]/NET0131 ,
		_w1867_,
		_w4011_
	);
	LUT2 #(
		.INIT('h1)
	) name3480 (
		_w1792_,
		_w4011_,
		_w4012_
	);
	LUT2 #(
		.INIT('h2)
	) name3481 (
		\sa21_reg[2]/P0001 ,
		_w4012_,
		_w4013_
	);
	LUT2 #(
		.INIT('h8)
	) name3482 (
		_w1877_,
		_w2993_,
		_w4014_
	);
	LUT2 #(
		.INIT('h2)
	) name3483 (
		\sa21_reg[1]/P0001 ,
		_w4007_,
		_w4015_
	);
	LUT2 #(
		.INIT('h4)
	) name3484 (
		_w4014_,
		_w4015_,
		_w4016_
	);
	LUT2 #(
		.INIT('h4)
	) name3485 (
		_w4010_,
		_w4016_,
		_w4017_
	);
	LUT2 #(
		.INIT('h4)
	) name3486 (
		_w4013_,
		_w4017_,
		_w4018_
	);
	LUT2 #(
		.INIT('h8)
	) name3487 (
		\sa21_reg[3]/P0001 ,
		_w1822_,
		_w4019_
	);
	LUT2 #(
		.INIT('h8)
	) name3488 (
		_w2479_,
		_w4019_,
		_w4020_
	);
	LUT2 #(
		.INIT('h1)
	) name3489 (
		_w1864_,
		_w2417_,
		_w4021_
	);
	LUT2 #(
		.INIT('h2)
	) name3490 (
		_w1831_,
		_w4021_,
		_w4022_
	);
	LUT2 #(
		.INIT('h1)
	) name3491 (
		\sa21_reg[1]/P0001 ,
		_w4020_,
		_w4023_
	);
	LUT2 #(
		.INIT('h4)
	) name3492 (
		_w4022_,
		_w4023_,
		_w4024_
	);
	LUT2 #(
		.INIT('h1)
	) name3493 (
		_w4018_,
		_w4024_,
		_w4025_
	);
	LUT2 #(
		.INIT('h1)
	) name3494 (
		_w1794_,
		_w2426_,
		_w4026_
	);
	LUT2 #(
		.INIT('h2)
	) name3495 (
		_w1894_,
		_w4026_,
		_w4027_
	);
	LUT2 #(
		.INIT('h2)
	) name3496 (
		_w3511_,
		_w3994_,
		_w4028_
	);
	LUT2 #(
		.INIT('h1)
	) name3497 (
		\sa21_reg[2]/P0001 ,
		_w4028_,
		_w4029_
	);
	LUT2 #(
		.INIT('h4)
	) name3498 (
		_w2842_,
		_w2919_,
		_w4030_
	);
	LUT2 #(
		.INIT('h2)
	) name3499 (
		_w2917_,
		_w4030_,
		_w4031_
	);
	LUT2 #(
		.INIT('h8)
	) name3500 (
		_w1832_,
		_w2448_,
		_w4032_
	);
	LUT2 #(
		.INIT('h2)
	) name3501 (
		_w1772_,
		_w1854_,
		_w4033_
	);
	LUT2 #(
		.INIT('h1)
	) name3502 (
		_w2490_,
		_w4033_,
		_w4034_
	);
	LUT2 #(
		.INIT('h2)
	) name3503 (
		\sa21_reg[2]/P0001 ,
		_w4034_,
		_w4035_
	);
	LUT2 #(
		.INIT('h2)
	) name3504 (
		\sa21_reg[1]/P0001 ,
		_w2446_,
		_w4036_
	);
	LUT2 #(
		.INIT('h1)
	) name3505 (
		_w2508_,
		_w3040_,
		_w4037_
	);
	LUT2 #(
		.INIT('h4)
	) name3506 (
		_w4032_,
		_w4037_,
		_w4038_
	);
	LUT2 #(
		.INIT('h4)
	) name3507 (
		_w1792_,
		_w4036_,
		_w4039_
	);
	LUT2 #(
		.INIT('h8)
	) name3508 (
		_w4038_,
		_w4039_,
		_w4040_
	);
	LUT2 #(
		.INIT('h4)
	) name3509 (
		_w4035_,
		_w4040_,
		_w4041_
	);
	LUT2 #(
		.INIT('h1)
	) name3510 (
		_w2513_,
		_w2838_,
		_w4042_
	);
	LUT2 #(
		.INIT('h1)
	) name3511 (
		\sa21_reg[2]/P0001 ,
		_w4042_,
		_w4043_
	);
	LUT2 #(
		.INIT('h1)
	) name3512 (
		_w1788_,
		_w1879_,
		_w4044_
	);
	LUT2 #(
		.INIT('h1)
	) name3513 (
		_w2479_,
		_w4044_,
		_w4045_
	);
	LUT2 #(
		.INIT('h1)
	) name3514 (
		\sa21_reg[1]/P0001 ,
		_w1865_,
		_w4046_
	);
	LUT2 #(
		.INIT('h4)
	) name3515 (
		_w1891_,
		_w4046_,
		_w4047_
	);
	LUT2 #(
		.INIT('h4)
	) name3516 (
		_w2997_,
		_w4047_,
		_w4048_
	);
	LUT2 #(
		.INIT('h1)
	) name3517 (
		_w4043_,
		_w4045_,
		_w4049_
	);
	LUT2 #(
		.INIT('h8)
	) name3518 (
		_w4048_,
		_w4049_,
		_w4050_
	);
	LUT2 #(
		.INIT('h1)
	) name3519 (
		_w4041_,
		_w4050_,
		_w4051_
	);
	LUT2 #(
		.INIT('h1)
	) name3520 (
		_w2906_,
		_w4031_,
		_w4052_
	);
	LUT2 #(
		.INIT('h4)
	) name3521 (
		_w4029_,
		_w4052_,
		_w4053_
	);
	LUT2 #(
		.INIT('h4)
	) name3522 (
		_w4051_,
		_w4053_,
		_w4054_
	);
	LUT2 #(
		.INIT('h2)
	) name3523 (
		\sa21_reg[0]/P0001 ,
		_w4054_,
		_w4055_
	);
	LUT2 #(
		.INIT('h1)
	) name3524 (
		_w1874_,
		_w4027_,
		_w4056_
	);
	LUT2 #(
		.INIT('h4)
	) name3525 (
		_w4025_,
		_w4056_,
		_w4057_
	);
	LUT2 #(
		.INIT('h4)
	) name3526 (
		_w4006_,
		_w4057_,
		_w4058_
	);
	LUT2 #(
		.INIT('h4)
	) name3527 (
		_w4055_,
		_w4058_,
		_w4059_
	);
	LUT2 #(
		.INIT('h2)
	) name3528 (
		_w3966_,
		_w4059_,
		_w4060_
	);
	LUT2 #(
		.INIT('h4)
	) name3529 (
		_w3966_,
		_w4059_,
		_w4061_
	);
	LUT2 #(
		.INIT('h1)
	) name3530 (
		_w4060_,
		_w4061_,
		_w4062_
	);
	LUT2 #(
		.INIT('h2)
	) name3531 (
		_w2199_,
		_w2736_,
		_w4063_
	);
	LUT2 #(
		.INIT('h4)
	) name3532 (
		_w2199_,
		_w2736_,
		_w4064_
	);
	LUT2 #(
		.INIT('h1)
	) name3533 (
		_w4063_,
		_w4064_,
		_w4065_
	);
	LUT2 #(
		.INIT('h8)
	) name3534 (
		_w4062_,
		_w4065_,
		_w4066_
	);
	LUT2 #(
		.INIT('h1)
	) name3535 (
		_w4062_,
		_w4065_,
		_w4067_
	);
	LUT2 #(
		.INIT('h1)
	) name3536 (
		_w4066_,
		_w4067_,
		_w4068_
	);
	LUT2 #(
		.INIT('h1)
	) name3537 (
		\u0_w_reg[3][20]/P0001 ,
		_w3205_,
		_w4069_
	);
	LUT2 #(
		.INIT('h8)
	) name3538 (
		\u0_w_reg[3][20]/P0001 ,
		_w3205_,
		_w4070_
	);
	LUT2 #(
		.INIT('h1)
	) name3539 (
		_w4069_,
		_w4070_,
		_w4071_
	);
	LUT2 #(
		.INIT('h2)
	) name3540 (
		_w2529_,
		_w3069_,
		_w4072_
	);
	LUT2 #(
		.INIT('h4)
	) name3541 (
		_w2529_,
		_w3069_,
		_w4073_
	);
	LUT2 #(
		.INIT('h1)
	) name3542 (
		_w4072_,
		_w4073_,
		_w4074_
	);
	LUT2 #(
		.INIT('h8)
	) name3543 (
		_w4071_,
		_w4074_,
		_w4075_
	);
	LUT2 #(
		.INIT('h1)
	) name3544 (
		_w4071_,
		_w4074_,
		_w4076_
	);
	LUT2 #(
		.INIT('h1)
	) name3545 (
		_w4075_,
		_w4076_,
		_w4077_
	);
	LUT2 #(
		.INIT('h2)
	) name3546 (
		_w4068_,
		_w4077_,
		_w4078_
	);
	LUT2 #(
		.INIT('h4)
	) name3547 (
		_w4068_,
		_w4077_,
		_w4079_
	);
	LUT2 #(
		.INIT('h1)
	) name3548 (
		\ld_r_reg/P0001 ,
		_w4078_,
		_w4080_
	);
	LUT2 #(
		.INIT('h4)
	) name3549 (
		_w4079_,
		_w4080_,
		_w4081_
	);
	LUT2 #(
		.INIT('h2)
	) name3550 (
		\text_in_r_reg[20]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w4082_
	);
	LUT2 #(
		.INIT('h4)
	) name3551 (
		\text_in_r_reg[20]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w4083_
	);
	LUT2 #(
		.INIT('h2)
	) name3552 (
		\ld_r_reg/P0001 ,
		_w4082_,
		_w4084_
	);
	LUT2 #(
		.INIT('h4)
	) name3553 (
		_w4083_,
		_w4084_,
		_w4085_
	);
	LUT2 #(
		.INIT('h1)
	) name3554 (
		_w4081_,
		_w4085_,
		_w4086_
	);
	LUT2 #(
		.INIT('h1)
	) name3555 (
		_w1462_,
		_w2712_,
		_w4087_
	);
	LUT2 #(
		.INIT('h8)
	) name3556 (
		_w1481_,
		_w4087_,
		_w4088_
	);
	LUT2 #(
		.INIT('h2)
	) name3557 (
		\sa03_reg[2]/P0001 ,
		_w4088_,
		_w4089_
	);
	LUT2 #(
		.INIT('h1)
	) name3558 (
		_w1326_,
		_w1383_,
		_w4090_
	);
	LUT2 #(
		.INIT('h2)
	) name3559 (
		\sa03_reg[3]/P0001 ,
		_w4090_,
		_w4091_
	);
	LUT2 #(
		.INIT('h1)
	) name3560 (
		_w2236_,
		_w2279_,
		_w4092_
	);
	LUT2 #(
		.INIT('h4)
	) name3561 (
		_w4091_,
		_w4092_,
		_w4093_
	);
	LUT2 #(
		.INIT('h1)
	) name3562 (
		\sa03_reg[2]/P0001 ,
		_w4093_,
		_w4094_
	);
	LUT2 #(
		.INIT('h1)
	) name3563 (
		_w1326_,
		_w1329_,
		_w4095_
	);
	LUT2 #(
		.INIT('h1)
	) name3564 (
		\sa03_reg[2]/P0001 ,
		_w1332_,
		_w4096_
	);
	LUT2 #(
		.INIT('h8)
	) name3565 (
		_w4095_,
		_w4096_,
		_w4097_
	);
	LUT2 #(
		.INIT('h1)
	) name3566 (
		_w1566_,
		_w4097_,
		_w4098_
	);
	LUT2 #(
		.INIT('h2)
	) name3567 (
		\sa03_reg[1]/P0001 ,
		_w4098_,
		_w4099_
	);
	LUT2 #(
		.INIT('h8)
	) name3568 (
		_w2206_,
		_w2225_,
		_w4100_
	);
	LUT2 #(
		.INIT('h2)
	) name3569 (
		_w1423_,
		_w2226_,
		_w4101_
	);
	LUT2 #(
		.INIT('h8)
	) name3570 (
		_w1352_,
		_w1449_,
		_w4102_
	);
	LUT2 #(
		.INIT('h1)
	) name3571 (
		_w1343_,
		_w1556_,
		_w4103_
	);
	LUT2 #(
		.INIT('h4)
	) name3572 (
		_w1397_,
		_w4103_,
		_w4104_
	);
	LUT2 #(
		.INIT('h2)
	) name3573 (
		\sa03_reg[2]/P0001 ,
		_w4104_,
		_w4105_
	);
	LUT2 #(
		.INIT('h1)
	) name3574 (
		_w4101_,
		_w4102_,
		_w4106_
	);
	LUT2 #(
		.INIT('h4)
	) name3575 (
		_w4100_,
		_w4106_,
		_w4107_
	);
	LUT2 #(
		.INIT('h4)
	) name3576 (
		_w4105_,
		_w4107_,
		_w4108_
	);
	LUT2 #(
		.INIT('h1)
	) name3577 (
		\sa03_reg[1]/P0001 ,
		_w4108_,
		_w4109_
	);
	LUT2 #(
		.INIT('h1)
	) name3578 (
		_w2289_,
		_w2693_,
		_w4110_
	);
	LUT2 #(
		.INIT('h4)
	) name3579 (
		_w4099_,
		_w4110_,
		_w4111_
	);
	LUT2 #(
		.INIT('h4)
	) name3580 (
		_w4089_,
		_w4111_,
		_w4112_
	);
	LUT2 #(
		.INIT('h4)
	) name3581 (
		_w4094_,
		_w4112_,
		_w4113_
	);
	LUT2 #(
		.INIT('h4)
	) name3582 (
		_w4109_,
		_w4113_,
		_w4114_
	);
	LUT2 #(
		.INIT('h2)
	) name3583 (
		\sa03_reg[0]/P0001 ,
		_w4114_,
		_w4115_
	);
	LUT2 #(
		.INIT('h4)
	) name3584 (
		_w1541_,
		_w3833_,
		_w4116_
	);
	LUT2 #(
		.INIT('h1)
	) name3585 (
		\sa03_reg[2]/P0001 ,
		_w4116_,
		_w4117_
	);
	LUT2 #(
		.INIT('h2)
	) name3586 (
		\sa03_reg[5]/P0001 ,
		_w1323_,
		_w4118_
	);
	LUT2 #(
		.INIT('h8)
	) name3587 (
		_w1423_,
		_w3871_,
		_w4119_
	);
	LUT2 #(
		.INIT('h4)
	) name3588 (
		_w4118_,
		_w4119_,
		_w4120_
	);
	LUT2 #(
		.INIT('h2)
	) name3589 (
		_w1339_,
		_w1398_,
		_w4121_
	);
	LUT2 #(
		.INIT('h8)
	) name3590 (
		_w1494_,
		_w4121_,
		_w4122_
	);
	LUT2 #(
		.INIT('h1)
	) name3591 (
		\sa03_reg[3]/P0001 ,
		_w2201_,
		_w4123_
	);
	LUT2 #(
		.INIT('h1)
	) name3592 (
		_w2657_,
		_w4123_,
		_w4124_
	);
	LUT2 #(
		.INIT('h1)
	) name3593 (
		\sa03_reg[1]/P0001 ,
		_w4124_,
		_w4125_
	);
	LUT2 #(
		.INIT('h1)
	) name3594 (
		_w1316_,
		_w1323_,
		_w4126_
	);
	LUT2 #(
		.INIT('h1)
	) name3595 (
		_w3720_,
		_w4126_,
		_w4127_
	);
	LUT2 #(
		.INIT('h8)
	) name3596 (
		\sa03_reg[3]/P0001 ,
		_w2715_,
		_w4128_
	);
	LUT2 #(
		.INIT('h1)
	) name3597 (
		_w2250_,
		_w4127_,
		_w4129_
	);
	LUT2 #(
		.INIT('h4)
	) name3598 (
		_w4128_,
		_w4129_,
		_w4130_
	);
	LUT2 #(
		.INIT('h2)
	) name3599 (
		\sa03_reg[1]/P0001 ,
		_w4130_,
		_w4131_
	);
	LUT2 #(
		.INIT('h1)
	) name3600 (
		_w4120_,
		_w4122_,
		_w4132_
	);
	LUT2 #(
		.INIT('h4)
	) name3601 (
		_w4117_,
		_w4132_,
		_w4133_
	);
	LUT2 #(
		.INIT('h1)
	) name3602 (
		_w4125_,
		_w4131_,
		_w4134_
	);
	LUT2 #(
		.INIT('h8)
	) name3603 (
		_w4133_,
		_w4134_,
		_w4135_
	);
	LUT2 #(
		.INIT('h1)
	) name3604 (
		\sa03_reg[0]/P0001 ,
		_w4135_,
		_w4136_
	);
	LUT2 #(
		.INIT('h8)
	) name3605 (
		\sa03_reg[2]/P0001 ,
		_w1352_,
		_w4137_
	);
	LUT2 #(
		.INIT('h4)
	) name3606 (
		_w1376_,
		_w4137_,
		_w4138_
	);
	LUT2 #(
		.INIT('h8)
	) name3607 (
		_w4095_,
		_w4138_,
		_w4139_
	);
	LUT2 #(
		.INIT('h8)
	) name3608 (
		_w1446_,
		_w1515_,
		_w4140_
	);
	LUT2 #(
		.INIT('h1)
	) name3609 (
		_w1380_,
		_w1416_,
		_w4141_
	);
	LUT2 #(
		.INIT('h4)
	) name3610 (
		_w1482_,
		_w4141_,
		_w4142_
	);
	LUT2 #(
		.INIT('h2)
	) name3611 (
		_w2225_,
		_w4142_,
		_w4143_
	);
	LUT2 #(
		.INIT('h1)
	) name3612 (
		_w1415_,
		_w4139_,
		_w4144_
	);
	LUT2 #(
		.INIT('h4)
	) name3613 (
		_w4140_,
		_w4144_,
		_w4145_
	);
	LUT2 #(
		.INIT('h4)
	) name3614 (
		_w4143_,
		_w4145_,
		_w4146_
	);
	LUT2 #(
		.INIT('h1)
	) name3615 (
		\sa03_reg[1]/P0001 ,
		_w4146_,
		_w4147_
	);
	LUT2 #(
		.INIT('h8)
	) name3616 (
		_w1435_,
		_w4137_,
		_w4148_
	);
	LUT2 #(
		.INIT('h8)
	) name3617 (
		\sa03_reg[6]/NET0131 ,
		_w1523_,
		_w4149_
	);
	LUT2 #(
		.INIT('h8)
	) name3618 (
		_w1436_,
		_w1566_,
		_w4150_
	);
	LUT2 #(
		.INIT('h4)
	) name3619 (
		\sa03_reg[2]/P0001 ,
		_w2293_,
		_w4151_
	);
	LUT2 #(
		.INIT('h1)
	) name3620 (
		_w1417_,
		_w1496_,
		_w4152_
	);
	LUT2 #(
		.INIT('h1)
	) name3621 (
		_w2670_,
		_w4151_,
		_w4153_
	);
	LUT2 #(
		.INIT('h8)
	) name3622 (
		_w4152_,
		_w4153_,
		_w4154_
	);
	LUT2 #(
		.INIT('h4)
	) name3623 (
		_w4150_,
		_w4154_,
		_w4155_
	);
	LUT2 #(
		.INIT('h2)
	) name3624 (
		\sa03_reg[1]/P0001 ,
		_w4155_,
		_w4156_
	);
	LUT2 #(
		.INIT('h1)
	) name3625 (
		_w4148_,
		_w4149_,
		_w4157_
	);
	LUT2 #(
		.INIT('h4)
	) name3626 (
		_w4156_,
		_w4157_,
		_w4158_
	);
	LUT2 #(
		.INIT('h4)
	) name3627 (
		_w4147_,
		_w4158_,
		_w4159_
	);
	LUT2 #(
		.INIT('h4)
	) name3628 (
		_w4136_,
		_w4159_,
		_w4160_
	);
	LUT2 #(
		.INIT('h4)
	) name3629 (
		_w4115_,
		_w4160_,
		_w4161_
	);
	LUT2 #(
		.INIT('h1)
	) name3630 (
		_w2304_,
		_w4161_,
		_w4162_
	);
	LUT2 #(
		.INIT('h8)
	) name3631 (
		_w2304_,
		_w4161_,
		_w4163_
	);
	LUT2 #(
		.INIT('h1)
	) name3632 (
		_w4162_,
		_w4163_,
		_w4164_
	);
	LUT2 #(
		.INIT('h2)
	) name3633 (
		_w3771_,
		_w4164_,
		_w4165_
	);
	LUT2 #(
		.INIT('h4)
	) name3634 (
		_w3771_,
		_w4164_,
		_w4166_
	);
	LUT2 #(
		.INIT('h1)
	) name3635 (
		_w4165_,
		_w4166_,
		_w4167_
	);
	LUT2 #(
		.INIT('h2)
	) name3636 (
		\sa21_reg[2]/P0001 ,
		_w1872_,
		_w4168_
	);
	LUT2 #(
		.INIT('h4)
	) name3637 (
		_w3048_,
		_w4168_,
		_w4169_
	);
	LUT2 #(
		.INIT('h1)
	) name3638 (
		\sa21_reg[2]/P0001 ,
		_w1865_,
		_w4170_
	);
	LUT2 #(
		.INIT('h4)
	) name3639 (
		_w2893_,
		_w4170_,
		_w4171_
	);
	LUT2 #(
		.INIT('h4)
	) name3640 (
		_w3050_,
		_w4171_,
		_w4172_
	);
	LUT2 #(
		.INIT('h1)
	) name3641 (
		_w4169_,
		_w4172_,
		_w4173_
	);
	LUT2 #(
		.INIT('h1)
	) name3642 (
		_w1760_,
		_w1884_,
		_w4174_
	);
	LUT2 #(
		.INIT('h1)
	) name3643 (
		\sa21_reg[2]/P0001 ,
		_w4174_,
		_w4175_
	);
	LUT2 #(
		.INIT('h8)
	) name3644 (
		\sa21_reg[2]/P0001 ,
		_w1838_,
		_w4176_
	);
	LUT2 #(
		.INIT('h1)
	) name3645 (
		\sa21_reg[1]/P0001 ,
		_w1874_,
		_w4177_
	);
	LUT2 #(
		.INIT('h1)
	) name3646 (
		_w3050_,
		_w4007_,
		_w4178_
	);
	LUT2 #(
		.INIT('h4)
	) name3647 (
		_w4176_,
		_w4178_,
		_w4179_
	);
	LUT2 #(
		.INIT('h8)
	) name3648 (
		_w4177_,
		_w4179_,
		_w4180_
	);
	LUT2 #(
		.INIT('h4)
	) name3649 (
		_w4175_,
		_w4180_,
		_w4181_
	);
	LUT2 #(
		.INIT('h1)
	) name3650 (
		\sa21_reg[2]/P0001 ,
		_w1833_,
		_w4182_
	);
	LUT2 #(
		.INIT('h1)
	) name3651 (
		_w1873_,
		_w3542_,
		_w4183_
	);
	LUT2 #(
		.INIT('h8)
	) name3652 (
		_w4182_,
		_w4183_,
		_w4184_
	);
	LUT2 #(
		.INIT('h4)
	) name3653 (
		\sa21_reg[3]/P0001 ,
		_w1781_,
		_w4185_
	);
	LUT2 #(
		.INIT('h2)
	) name3654 (
		\sa21_reg[2]/P0001 ,
		_w1849_,
		_w4186_
	);
	LUT2 #(
		.INIT('h4)
	) name3655 (
		_w4185_,
		_w4186_,
		_w4187_
	);
	LUT2 #(
		.INIT('h1)
	) name3656 (
		_w4184_,
		_w4187_,
		_w4188_
	);
	LUT2 #(
		.INIT('h2)
	) name3657 (
		\sa21_reg[1]/P0001 ,
		_w2502_,
		_w4189_
	);
	LUT2 #(
		.INIT('h8)
	) name3658 (
		_w2877_,
		_w4189_,
		_w4190_
	);
	LUT2 #(
		.INIT('h4)
	) name3659 (
		_w4188_,
		_w4190_,
		_w4191_
	);
	LUT2 #(
		.INIT('h1)
	) name3660 (
		_w4181_,
		_w4191_,
		_w4192_
	);
	LUT2 #(
		.INIT('h1)
	) name3661 (
		_w2928_,
		_w4173_,
		_w4193_
	);
	LUT2 #(
		.INIT('h4)
	) name3662 (
		_w4192_,
		_w4193_,
		_w4194_
	);
	LUT2 #(
		.INIT('h1)
	) name3663 (
		\sa21_reg[0]/P0001 ,
		_w4194_,
		_w4195_
	);
	LUT2 #(
		.INIT('h1)
	) name3664 (
		_w1794_,
		_w3982_,
		_w4196_
	);
	LUT2 #(
		.INIT('h8)
	) name3665 (
		\sa21_reg[4]/P0001 ,
		_w1758_,
		_w4197_
	);
	LUT2 #(
		.INIT('h4)
	) name3666 (
		\sa21_reg[5]/P0001 ,
		_w1793_,
		_w4198_
	);
	LUT2 #(
		.INIT('h1)
	) name3667 (
		_w4019_,
		_w4197_,
		_w4199_
	);
	LUT2 #(
		.INIT('h4)
	) name3668 (
		_w4198_,
		_w4199_,
		_w4200_
	);
	LUT2 #(
		.INIT('h2)
	) name3669 (
		\sa21_reg[2]/P0001 ,
		_w4200_,
		_w4201_
	);
	LUT2 #(
		.INIT('h2)
	) name3670 (
		_w4196_,
		_w4201_,
		_w4202_
	);
	LUT2 #(
		.INIT('h2)
	) name3671 (
		\sa21_reg[1]/P0001 ,
		_w4202_,
		_w4203_
	);
	LUT2 #(
		.INIT('h4)
	) name3672 (
		\sa21_reg[2]/P0001 ,
		_w2842_,
		_w4204_
	);
	LUT2 #(
		.INIT('h4)
	) name3673 (
		_w1784_,
		_w3518_,
		_w4205_
	);
	LUT2 #(
		.INIT('h8)
	) name3674 (
		_w1772_,
		_w1816_,
		_w4206_
	);
	LUT2 #(
		.INIT('h1)
	) name3675 (
		_w2417_,
		_w4204_,
		_w4207_
	);
	LUT2 #(
		.INIT('h4)
	) name3676 (
		_w4206_,
		_w4207_,
		_w4208_
	);
	LUT2 #(
		.INIT('h4)
	) name3677 (
		_w4205_,
		_w4208_,
		_w4209_
	);
	LUT2 #(
		.INIT('h1)
	) name3678 (
		\sa21_reg[1]/P0001 ,
		_w4209_,
		_w4210_
	);
	LUT2 #(
		.INIT('h8)
	) name3679 (
		_w1823_,
		_w3026_,
		_w4211_
	);
	LUT2 #(
		.INIT('h4)
	) name3680 (
		_w1894_,
		_w2493_,
		_w4212_
	);
	LUT2 #(
		.INIT('h1)
	) name3681 (
		_w1838_,
		_w2417_,
		_w4213_
	);
	LUT2 #(
		.INIT('h4)
	) name3682 (
		_w1885_,
		_w4213_,
		_w4214_
	);
	LUT2 #(
		.INIT('h1)
	) name3683 (
		\sa21_reg[2]/P0001 ,
		_w4214_,
		_w4215_
	);
	LUT2 #(
		.INIT('h1)
	) name3684 (
		_w4211_,
		_w4212_,
		_w4216_
	);
	LUT2 #(
		.INIT('h4)
	) name3685 (
		_w4215_,
		_w4216_,
		_w4217_
	);
	LUT2 #(
		.INIT('h4)
	) name3686 (
		_w4203_,
		_w4217_,
		_w4218_
	);
	LUT2 #(
		.INIT('h4)
	) name3687 (
		_w4210_,
		_w4218_,
		_w4219_
	);
	LUT2 #(
		.INIT('h2)
	) name3688 (
		\sa21_reg[0]/P0001 ,
		_w4219_,
		_w4220_
	);
	LUT2 #(
		.INIT('h1)
	) name3689 (
		_w1794_,
		_w1853_,
		_w4221_
	);
	LUT2 #(
		.INIT('h2)
	) name3690 (
		\sa21_reg[3]/P0001 ,
		_w4221_,
		_w4222_
	);
	LUT2 #(
		.INIT('h1)
	) name3691 (
		_w1824_,
		_w4222_,
		_w4223_
	);
	LUT2 #(
		.INIT('h2)
	) name3692 (
		_w1863_,
		_w4223_,
		_w4224_
	);
	LUT2 #(
		.INIT('h1)
	) name3693 (
		_w1786_,
		_w2426_,
		_w4225_
	);
	LUT2 #(
		.INIT('h2)
	) name3694 (
		_w1894_,
		_w4225_,
		_w4226_
	);
	LUT2 #(
		.INIT('h8)
	) name3695 (
		_w1772_,
		_w1815_,
		_w4227_
	);
	LUT2 #(
		.INIT('h1)
	) name3696 (
		_w1800_,
		_w2502_,
		_w4228_
	);
	LUT2 #(
		.INIT('h4)
	) name3697 (
		_w4227_,
		_w4228_,
		_w4229_
	);
	LUT2 #(
		.INIT('h1)
	) name3698 (
		_w1776_,
		_w1786_,
		_w4230_
	);
	LUT2 #(
		.INIT('h8)
	) name3699 (
		_w4229_,
		_w4230_,
		_w4231_
	);
	LUT2 #(
		.INIT('h2)
	) name3700 (
		\sa21_reg[1]/P0001 ,
		\sa21_reg[2]/P0001 ,
		_w4232_
	);
	LUT2 #(
		.INIT('h4)
	) name3701 (
		_w4231_,
		_w4232_,
		_w4233_
	);
	LUT2 #(
		.INIT('h1)
	) name3702 (
		_w1782_,
		_w1865_,
		_w4234_
	);
	LUT2 #(
		.INIT('h4)
	) name3703 (
		_w3543_,
		_w4234_,
		_w4235_
	);
	LUT2 #(
		.INIT('h2)
	) name3704 (
		_w3529_,
		_w4235_,
		_w4236_
	);
	LUT2 #(
		.INIT('h1)
	) name3705 (
		_w1751_,
		_w2513_,
		_w4237_
	);
	LUT2 #(
		.INIT('h4)
	) name3706 (
		_w2894_,
		_w4237_,
		_w4238_
	);
	LUT2 #(
		.INIT('h1)
	) name3707 (
		\sa21_reg[2]/P0001 ,
		_w4238_,
		_w4239_
	);
	LUT2 #(
		.INIT('h1)
	) name3708 (
		_w1748_,
		_w3056_,
		_w4240_
	);
	LUT2 #(
		.INIT('h4)
	) name3709 (
		_w4239_,
		_w4240_,
		_w4241_
	);
	LUT2 #(
		.INIT('h1)
	) name3710 (
		\sa21_reg[1]/P0001 ,
		_w4241_,
		_w4242_
	);
	LUT2 #(
		.INIT('h1)
	) name3711 (
		_w4224_,
		_w4226_,
		_w4243_
	);
	LUT2 #(
		.INIT('h1)
	) name3712 (
		_w4233_,
		_w4236_,
		_w4244_
	);
	LUT2 #(
		.INIT('h8)
	) name3713 (
		_w4243_,
		_w4244_,
		_w4245_
	);
	LUT2 #(
		.INIT('h4)
	) name3714 (
		_w4242_,
		_w4245_,
		_w4246_
	);
	LUT2 #(
		.INIT('h4)
	) name3715 (
		_w4195_,
		_w4246_,
		_w4247_
	);
	LUT2 #(
		.INIT('h4)
	) name3716 (
		_w4220_,
		_w4247_,
		_w4248_
	);
	LUT2 #(
		.INIT('h2)
	) name3717 (
		\u0_w_reg[3][1]/P0001 ,
		_w4248_,
		_w4249_
	);
	LUT2 #(
		.INIT('h4)
	) name3718 (
		\u0_w_reg[3][1]/P0001 ,
		_w4248_,
		_w4250_
	);
	LUT2 #(
		.INIT('h1)
	) name3719 (
		_w4249_,
		_w4250_,
		_w4251_
	);
	LUT2 #(
		.INIT('h8)
	) name3720 (
		_w3419_,
		_w4251_,
		_w4252_
	);
	LUT2 #(
		.INIT('h1)
	) name3721 (
		_w3419_,
		_w4251_,
		_w4253_
	);
	LUT2 #(
		.INIT('h1)
	) name3722 (
		_w4252_,
		_w4253_,
		_w4254_
	);
	LUT2 #(
		.INIT('h1)
	) name3723 (
		_w4167_,
		_w4254_,
		_w4255_
	);
	LUT2 #(
		.INIT('h8)
	) name3724 (
		_w4167_,
		_w4254_,
		_w4256_
	);
	LUT2 #(
		.INIT('h1)
	) name3725 (
		\ld_r_reg/P0001 ,
		_w4255_,
		_w4257_
	);
	LUT2 #(
		.INIT('h4)
	) name3726 (
		_w4256_,
		_w4257_,
		_w4258_
	);
	LUT2 #(
		.INIT('h1)
	) name3727 (
		\text_in_r_reg[1]/P0001 ,
		\u0_w_reg[3][1]/P0001 ,
		_w4259_
	);
	LUT2 #(
		.INIT('h8)
	) name3728 (
		\text_in_r_reg[1]/P0001 ,
		\u0_w_reg[3][1]/P0001 ,
		_w4260_
	);
	LUT2 #(
		.INIT('h2)
	) name3729 (
		\ld_r_reg/P0001 ,
		_w4259_,
		_w4261_
	);
	LUT2 #(
		.INIT('h4)
	) name3730 (
		_w4260_,
		_w4261_,
		_w4262_
	);
	LUT2 #(
		.INIT('h1)
	) name3731 (
		_w4258_,
		_w4262_,
		_w4263_
	);
	LUT2 #(
		.INIT('h1)
	) name3732 (
		_w1989_,
		_w2366_,
		_w4264_
	);
	LUT2 #(
		.INIT('h1)
	) name3733 (
		\sa32_reg[2]/P0001 ,
		_w4264_,
		_w4265_
	);
	LUT2 #(
		.INIT('h2)
	) name3734 (
		_w1926_,
		_w1959_,
		_w4266_
	);
	LUT2 #(
		.INIT('h2)
	) name3735 (
		\sa32_reg[2]/P0001 ,
		_w4266_,
		_w4267_
	);
	LUT2 #(
		.INIT('h1)
	) name3736 (
		_w2040_,
		_w2345_,
		_w4268_
	);
	LUT2 #(
		.INIT('h4)
	) name3737 (
		_w3490_,
		_w4268_,
		_w4269_
	);
	LUT2 #(
		.INIT('h4)
	) name3738 (
		_w4265_,
		_w4269_,
		_w4270_
	);
	LUT2 #(
		.INIT('h4)
	) name3739 (
		_w4267_,
		_w4270_,
		_w4271_
	);
	LUT2 #(
		.INIT('h1)
	) name3740 (
		\sa32_reg[1]/P0001 ,
		_w4271_,
		_w4272_
	);
	LUT2 #(
		.INIT('h2)
	) name3741 (
		_w3280_,
		_w3367_,
		_w4273_
	);
	LUT2 #(
		.INIT('h1)
	) name3742 (
		\sa32_reg[2]/P0001 ,
		_w4273_,
		_w4274_
	);
	LUT2 #(
		.INIT('h4)
	) name3743 (
		_w1932_,
		_w2042_,
		_w4275_
	);
	LUT2 #(
		.INIT('h2)
	) name3744 (
		_w2046_,
		_w4275_,
		_w4276_
	);
	LUT2 #(
		.INIT('h1)
	) name3745 (
		_w2024_,
		_w3194_,
		_w4277_
	);
	LUT2 #(
		.INIT('h1)
	) name3746 (
		_w3143_,
		_w3149_,
		_w4278_
	);
	LUT2 #(
		.INIT('h4)
	) name3747 (
		_w3457_,
		_w4278_,
		_w4279_
	);
	LUT2 #(
		.INIT('h2)
	) name3748 (
		\sa32_reg[2]/P0001 ,
		_w4279_,
		_w4280_
	);
	LUT2 #(
		.INIT('h1)
	) name3749 (
		_w1937_,
		_w1982_,
		_w4281_
	);
	LUT2 #(
		.INIT('h1)
	) name3750 (
		\sa32_reg[2]/P0001 ,
		_w4281_,
		_w4282_
	);
	LUT2 #(
		.INIT('h4)
	) name3751 (
		_w1921_,
		_w4277_,
		_w4283_
	);
	LUT2 #(
		.INIT('h4)
	) name3752 (
		_w4282_,
		_w4283_,
		_w4284_
	);
	LUT2 #(
		.INIT('h4)
	) name3753 (
		_w4280_,
		_w4284_,
		_w4285_
	);
	LUT2 #(
		.INIT('h2)
	) name3754 (
		\sa32_reg[1]/P0001 ,
		_w4285_,
		_w4286_
	);
	LUT2 #(
		.INIT('h1)
	) name3755 (
		_w1971_,
		_w4276_,
		_w4287_
	);
	LUT2 #(
		.INIT('h4)
	) name3756 (
		_w4274_,
		_w4287_,
		_w4288_
	);
	LUT2 #(
		.INIT('h4)
	) name3757 (
		_w4286_,
		_w4288_,
		_w4289_
	);
	LUT2 #(
		.INIT('h4)
	) name3758 (
		_w4272_,
		_w4289_,
		_w4290_
	);
	LUT2 #(
		.INIT('h2)
	) name3759 (
		\sa32_reg[0]/P0002 ,
		_w4290_,
		_w4291_
	);
	LUT2 #(
		.INIT('h4)
	) name3760 (
		\sa32_reg[2]/P0001 ,
		_w1994_,
		_w4292_
	);
	LUT2 #(
		.INIT('h8)
	) name3761 (
		_w1910_,
		_w1919_,
		_w4293_
	);
	LUT2 #(
		.INIT('h1)
	) name3762 (
		_w2399_,
		_w4293_,
		_w4294_
	);
	LUT2 #(
		.INIT('h2)
	) name3763 (
		\sa32_reg[2]/P0001 ,
		_w4294_,
		_w4295_
	);
	LUT2 #(
		.INIT('h2)
	) name3764 (
		\sa32_reg[1]/P0001 ,
		_w1925_,
		_w4296_
	);
	LUT2 #(
		.INIT('h4)
	) name3765 (
		_w3450_,
		_w4296_,
		_w4297_
	);
	LUT2 #(
		.INIT('h4)
	) name3766 (
		_w4292_,
		_w4297_,
		_w4298_
	);
	LUT2 #(
		.INIT('h4)
	) name3767 (
		_w2013_,
		_w4298_,
		_w4299_
	);
	LUT2 #(
		.INIT('h4)
	) name3768 (
		_w4295_,
		_w4299_,
		_w4300_
	);
	LUT2 #(
		.INIT('h8)
	) name3769 (
		_w1913_,
		_w2046_,
		_w4301_
	);
	LUT2 #(
		.INIT('h2)
	) name3770 (
		\sa32_reg[7]/P0001 ,
		_w1990_,
		_w4302_
	);
	LUT2 #(
		.INIT('h8)
	) name3771 (
		_w2397_,
		_w4302_,
		_w4303_
	);
	LUT2 #(
		.INIT('h1)
	) name3772 (
		\sa32_reg[1]/P0001 ,
		_w4301_,
		_w4304_
	);
	LUT2 #(
		.INIT('h4)
	) name3773 (
		_w3338_,
		_w4304_,
		_w4305_
	);
	LUT2 #(
		.INIT('h1)
	) name3774 (
		_w3367_,
		_w4303_,
		_w4306_
	);
	LUT2 #(
		.INIT('h8)
	) name3775 (
		_w4305_,
		_w4306_,
		_w4307_
	);
	LUT2 #(
		.INIT('h4)
	) name3776 (
		_w2365_,
		_w4307_,
		_w4308_
	);
	LUT2 #(
		.INIT('h1)
	) name3777 (
		_w4300_,
		_w4308_,
		_w4309_
	);
	LUT2 #(
		.INIT('h1)
	) name3778 (
		\sa32_reg[2]/P0001 ,
		_w2328_,
		_w4310_
	);
	LUT2 #(
		.INIT('h8)
	) name3779 (
		_w2059_,
		_w2399_,
		_w4311_
	);
	LUT2 #(
		.INIT('h1)
	) name3780 (
		_w1966_,
		_w2347_,
		_w4312_
	);
	LUT2 #(
		.INIT('h4)
	) name3781 (
		_w4311_,
		_w4312_,
		_w4313_
	);
	LUT2 #(
		.INIT('h4)
	) name3782 (
		_w4310_,
		_w4313_,
		_w4314_
	);
	LUT2 #(
		.INIT('h4)
	) name3783 (
		_w4309_,
		_w4314_,
		_w4315_
	);
	LUT2 #(
		.INIT('h1)
	) name3784 (
		\sa32_reg[0]/P0002 ,
		_w4315_,
		_w4316_
	);
	LUT2 #(
		.INIT('h8)
	) name3785 (
		_w1925_,
		_w2030_,
		_w4317_
	);
	LUT2 #(
		.INIT('h8)
	) name3786 (
		\sa32_reg[6]/NET0131 ,
		_w1952_,
		_w4318_
	);
	LUT2 #(
		.INIT('h2)
	) name3787 (
		_w4277_,
		_w4318_,
		_w4319_
	);
	LUT2 #(
		.INIT('h2)
	) name3788 (
		\sa32_reg[2]/P0001 ,
		_w4319_,
		_w4320_
	);
	LUT2 #(
		.INIT('h1)
	) name3789 (
		_w1994_,
		_w3180_,
		_w4321_
	);
	LUT2 #(
		.INIT('h4)
	) name3790 (
		_w3374_,
		_w4321_,
		_w4322_
	);
	LUT2 #(
		.INIT('h2)
	) name3791 (
		_w2313_,
		_w4322_,
		_w4323_
	);
	LUT2 #(
		.INIT('h1)
	) name3792 (
		_w4317_,
		_w4320_,
		_w4324_
	);
	LUT2 #(
		.INIT('h4)
	) name3793 (
		_w4323_,
		_w4324_,
		_w4325_
	);
	LUT2 #(
		.INIT('h2)
	) name3794 (
		\sa32_reg[1]/P0001 ,
		_w4325_,
		_w4326_
	);
	LUT2 #(
		.INIT('h1)
	) name3795 (
		_w3181_,
		_w3408_,
		_w4327_
	);
	LUT2 #(
		.INIT('h2)
	) name3796 (
		_w2059_,
		_w4327_,
		_w4328_
	);
	LUT2 #(
		.INIT('h2)
	) name3797 (
		\sa32_reg[2]/P0001 ,
		_w1938_,
		_w4329_
	);
	LUT2 #(
		.INIT('h4)
	) name3798 (
		_w1966_,
		_w4329_,
		_w4330_
	);
	LUT2 #(
		.INIT('h1)
	) name3799 (
		\sa32_reg[2]/P0001 ,
		_w3172_,
		_w4331_
	);
	LUT2 #(
		.INIT('h1)
	) name3800 (
		\sa32_reg[1]/P0001 ,
		_w4331_,
		_w4332_
	);
	LUT2 #(
		.INIT('h4)
	) name3801 (
		_w4330_,
		_w4332_,
		_w4333_
	);
	LUT2 #(
		.INIT('h1)
	) name3802 (
		_w3437_,
		_w4328_,
		_w4334_
	);
	LUT2 #(
		.INIT('h4)
	) name3803 (
		_w4333_,
		_w4334_,
		_w4335_
	);
	LUT2 #(
		.INIT('h4)
	) name3804 (
		_w4326_,
		_w4335_,
		_w4336_
	);
	LUT2 #(
		.INIT('h4)
	) name3805 (
		_w4291_,
		_w4336_,
		_w4337_
	);
	LUT2 #(
		.INIT('h4)
	) name3806 (
		_w4316_,
		_w4337_,
		_w4338_
	);
	LUT2 #(
		.INIT('h2)
	) name3807 (
		_w3416_,
		_w4338_,
		_w4339_
	);
	LUT2 #(
		.INIT('h4)
	) name3808 (
		_w3416_,
		_w4338_,
		_w4340_
	);
	LUT2 #(
		.INIT('h1)
	) name3809 (
		_w4339_,
		_w4340_,
		_w4341_
	);
	LUT2 #(
		.INIT('h2)
	) name3810 (
		\u0_w_reg[3][12]/P0001 ,
		_w3205_,
		_w4342_
	);
	LUT2 #(
		.INIT('h4)
	) name3811 (
		\u0_w_reg[3][12]/P0001 ,
		_w3205_,
		_w4343_
	);
	LUT2 #(
		.INIT('h1)
	) name3812 (
		_w4342_,
		_w4343_,
		_w4344_
	);
	LUT2 #(
		.INIT('h8)
	) name3813 (
		_w4341_,
		_w4344_,
		_w4345_
	);
	LUT2 #(
		.INIT('h1)
	) name3814 (
		_w4341_,
		_w4344_,
		_w4346_
	);
	LUT2 #(
		.INIT('h1)
	) name3815 (
		_w4345_,
		_w4346_,
		_w4347_
	);
	LUT2 #(
		.INIT('h2)
	) name3816 (
		_w2529_,
		_w4059_,
		_w4348_
	);
	LUT2 #(
		.INIT('h4)
	) name3817 (
		_w2529_,
		_w4059_,
		_w4349_
	);
	LUT2 #(
		.INIT('h1)
	) name3818 (
		_w4348_,
		_w4349_,
		_w4350_
	);
	LUT2 #(
		.INIT('h4)
	) name3819 (
		_w2739_,
		_w4350_,
		_w4351_
	);
	LUT2 #(
		.INIT('h2)
	) name3820 (
		_w2739_,
		_w4350_,
		_w4352_
	);
	LUT2 #(
		.INIT('h1)
	) name3821 (
		_w4351_,
		_w4352_,
		_w4353_
	);
	LUT2 #(
		.INIT('h2)
	) name3822 (
		_w4347_,
		_w4353_,
		_w4354_
	);
	LUT2 #(
		.INIT('h4)
	) name3823 (
		_w4347_,
		_w4353_,
		_w4355_
	);
	LUT2 #(
		.INIT('h1)
	) name3824 (
		\ld_r_reg/P0001 ,
		_w4354_,
		_w4356_
	);
	LUT2 #(
		.INIT('h4)
	) name3825 (
		_w4355_,
		_w4356_,
		_w4357_
	);
	LUT2 #(
		.INIT('h2)
	) name3826 (
		\text_in_r_reg[12]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		_w4358_
	);
	LUT2 #(
		.INIT('h4)
	) name3827 (
		\text_in_r_reg[12]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		_w4359_
	);
	LUT2 #(
		.INIT('h2)
	) name3828 (
		\ld_r_reg/P0001 ,
		_w4358_,
		_w4360_
	);
	LUT2 #(
		.INIT('h4)
	) name3829 (
		_w4359_,
		_w4360_,
		_w4361_
	);
	LUT2 #(
		.INIT('h1)
	) name3830 (
		_w4357_,
		_w4361_,
		_w4362_
	);
	LUT2 #(
		.INIT('h8)
	) name3831 (
		_w1698_,
		_w2595_,
		_w4363_
	);
	LUT2 #(
		.INIT('h1)
	) name3832 (
		_w2123_,
		_w2566_,
		_w4364_
	);
	LUT2 #(
		.INIT('h1)
	) name3833 (
		_w2576_,
		_w2586_,
		_w4365_
	);
	LUT2 #(
		.INIT('h8)
	) name3834 (
		_w4364_,
		_w4365_,
		_w4366_
	);
	LUT2 #(
		.INIT('h1)
	) name3835 (
		_w1616_,
		_w2622_,
		_w4367_
	);
	LUT2 #(
		.INIT('h1)
	) name3836 (
		_w2635_,
		_w4363_,
		_w4368_
	);
	LUT2 #(
		.INIT('h8)
	) name3837 (
		_w4367_,
		_w4368_,
		_w4369_
	);
	LUT2 #(
		.INIT('h8)
	) name3838 (
		_w4366_,
		_w4369_,
		_w4370_
	);
	LUT2 #(
		.INIT('h1)
	) name3839 (
		\sa10_reg[1]/P0001 ,
		_w4370_,
		_w4371_
	);
	LUT2 #(
		.INIT('h8)
	) name3840 (
		\sa10_reg[5]/P0001 ,
		_w2576_,
		_w4372_
	);
	LUT2 #(
		.INIT('h1)
	) name3841 (
		_w1708_,
		_w2809_,
		_w4373_
	);
	LUT2 #(
		.INIT('h4)
	) name3842 (
		_w2119_,
		_w4373_,
		_w4374_
	);
	LUT2 #(
		.INIT('h2)
	) name3843 (
		_w1664_,
		_w4374_,
		_w4375_
	);
	LUT2 #(
		.INIT('h8)
	) name3844 (
		_w2142_,
		_w3616_,
		_w4376_
	);
	LUT2 #(
		.INIT('h8)
	) name3845 (
		_w1629_,
		_w1666_,
		_w4377_
	);
	LUT2 #(
		.INIT('h8)
	) name3846 (
		_w1607_,
		_w4377_,
		_w4378_
	);
	LUT2 #(
		.INIT('h8)
	) name3847 (
		_w1586_,
		_w2112_,
		_w4379_
	);
	LUT2 #(
		.INIT('h1)
	) name3848 (
		_w4376_,
		_w4379_,
		_w4380_
	);
	LUT2 #(
		.INIT('h4)
	) name3849 (
		_w4378_,
		_w4380_,
		_w4381_
	);
	LUT2 #(
		.INIT('h2)
	) name3850 (
		\sa10_reg[1]/P0001 ,
		_w4381_,
		_w4382_
	);
	LUT2 #(
		.INIT('h1)
	) name3851 (
		_w2559_,
		_w4372_,
		_w4383_
	);
	LUT2 #(
		.INIT('h4)
	) name3852 (
		_w2572_,
		_w4383_,
		_w4384_
	);
	LUT2 #(
		.INIT('h4)
	) name3853 (
		_w4375_,
		_w4384_,
		_w4385_
	);
	LUT2 #(
		.INIT('h4)
	) name3854 (
		_w4382_,
		_w4385_,
		_w4386_
	);
	LUT2 #(
		.INIT('h4)
	) name3855 (
		_w4371_,
		_w4386_,
		_w4387_
	);
	LUT2 #(
		.INIT('h2)
	) name3856 (
		\sa10_reg[0]/P0001 ,
		_w4387_,
		_w4388_
	);
	LUT2 #(
		.INIT('h2)
	) name3857 (
		_w2190_,
		_w3922_,
		_w4389_
	);
	LUT2 #(
		.INIT('h4)
	) name3858 (
		_w2567_,
		_w4389_,
		_w4390_
	);
	LUT2 #(
		.INIT('h1)
	) name3859 (
		_w1683_,
		_w2101_,
		_w4391_
	);
	LUT2 #(
		.INIT('h4)
	) name3860 (
		_w1712_,
		_w4391_,
		_w4392_
	);
	LUT2 #(
		.INIT('h8)
	) name3861 (
		_w1617_,
		_w4392_,
		_w4393_
	);
	LUT2 #(
		.INIT('h1)
	) name3862 (
		_w4390_,
		_w4393_,
		_w4394_
	);
	LUT2 #(
		.INIT('h1)
	) name3863 (
		_w1583_,
		_w1586_,
		_w4395_
	);
	LUT2 #(
		.INIT('h8)
	) name3864 (
		_w1650_,
		_w4395_,
		_w4396_
	);
	LUT2 #(
		.INIT('h1)
	) name3865 (
		_w4394_,
		_w4396_,
		_w4397_
	);
	LUT2 #(
		.INIT('h1)
	) name3866 (
		\sa10_reg[1]/P0001 ,
		_w4397_,
		_w4398_
	);
	LUT2 #(
		.INIT('h1)
	) name3867 (
		_w1608_,
		_w1615_,
		_w4399_
	);
	LUT2 #(
		.INIT('h2)
	) name3868 (
		_w1668_,
		_w4399_,
		_w4400_
	);
	LUT2 #(
		.INIT('h1)
	) name3869 (
		_w1669_,
		_w2634_,
		_w4401_
	);
	LUT2 #(
		.INIT('h2)
	) name3870 (
		\sa10_reg[1]/P0001 ,
		_w4401_,
		_w4402_
	);
	LUT2 #(
		.INIT('h1)
	) name3871 (
		_w4400_,
		_w4402_,
		_w4403_
	);
	LUT2 #(
		.INIT('h2)
	) name3872 (
		\sa10_reg[2]/P0001 ,
		_w4403_,
		_w4404_
	);
	LUT2 #(
		.INIT('h1)
	) name3873 (
		_w2189_,
		_w4377_,
		_w4405_
	);
	LUT2 #(
		.INIT('h1)
	) name3874 (
		\sa10_reg[1]/P0001 ,
		_w4405_,
		_w4406_
	);
	LUT2 #(
		.INIT('h8)
	) name3875 (
		_w2607_,
		_w3943_,
		_w4407_
	);
	LUT2 #(
		.INIT('h1)
	) name3876 (
		_w1613_,
		_w4407_,
		_w4408_
	);
	LUT2 #(
		.INIT('h4)
	) name3877 (
		_w1728_,
		_w4408_,
		_w4409_
	);
	LUT2 #(
		.INIT('h4)
	) name3878 (
		_w4406_,
		_w4409_,
		_w4410_
	);
	LUT2 #(
		.INIT('h1)
	) name3879 (
		\sa10_reg[0]/P0001 ,
		_w4410_,
		_w4411_
	);
	LUT2 #(
		.INIT('h8)
	) name3880 (
		\sa10_reg[1]/P0001 ,
		_w1664_,
		_w4412_
	);
	LUT2 #(
		.INIT('h8)
	) name3881 (
		_w2093_,
		_w4412_,
		_w4413_
	);
	LUT2 #(
		.INIT('h8)
	) name3882 (
		\sa10_reg[4]/P0001 ,
		_w3641_,
		_w4414_
	);
	LUT2 #(
		.INIT('h2)
	) name3883 (
		_w3614_,
		_w4414_,
		_w4415_
	);
	LUT2 #(
		.INIT('h1)
	) name3884 (
		\sa10_reg[2]/P0001 ,
		_w4415_,
		_w4416_
	);
	LUT2 #(
		.INIT('h1)
	) name3885 (
		_w1698_,
		_w2608_,
		_w4417_
	);
	LUT2 #(
		.INIT('h2)
	) name3886 (
		\sa10_reg[2]/P0001 ,
		_w4417_,
		_w4418_
	);
	LUT2 #(
		.INIT('h1)
	) name3887 (
		_w1586_,
		_w1681_,
		_w4419_
	);
	LUT2 #(
		.INIT('h1)
	) name3888 (
		\sa10_reg[2]/P0001 ,
		_w1629_,
		_w4420_
	);
	LUT2 #(
		.INIT('h4)
	) name3889 (
		_w4419_,
		_w4420_,
		_w4421_
	);
	LUT2 #(
		.INIT('h1)
	) name3890 (
		_w1700_,
		_w4421_,
		_w4422_
	);
	LUT2 #(
		.INIT('h4)
	) name3891 (
		_w4418_,
		_w4422_,
		_w4423_
	);
	LUT2 #(
		.INIT('h1)
	) name3892 (
		\sa10_reg[0]/P0001 ,
		_w4423_,
		_w4424_
	);
	LUT2 #(
		.INIT('h1)
	) name3893 (
		_w2565_,
		_w4416_,
		_w4425_
	);
	LUT2 #(
		.INIT('h4)
	) name3894 (
		_w4424_,
		_w4425_,
		_w4426_
	);
	LUT2 #(
		.INIT('h2)
	) name3895 (
		\sa10_reg[1]/P0001 ,
		_w4426_,
		_w4427_
	);
	LUT2 #(
		.INIT('h1)
	) name3896 (
		_w3923_,
		_w4413_,
		_w4428_
	);
	LUT2 #(
		.INIT('h4)
	) name3897 (
		_w4404_,
		_w4428_,
		_w4429_
	);
	LUT2 #(
		.INIT('h4)
	) name3898 (
		_w4411_,
		_w4429_,
		_w4430_
	);
	LUT2 #(
		.INIT('h4)
	) name3899 (
		_w4398_,
		_w4430_,
		_w4431_
	);
	LUT2 #(
		.INIT('h4)
	) name3900 (
		_w4427_,
		_w4431_,
		_w4432_
	);
	LUT2 #(
		.INIT('h4)
	) name3901 (
		_w4388_,
		_w4432_,
		_w4433_
	);
	LUT2 #(
		.INIT('h4)
	) name3902 (
		_w1383_,
		_w3746_,
		_w4434_
	);
	LUT2 #(
		.INIT('h4)
	) name3903 (
		\sa03_reg[6]/NET0131 ,
		_w1324_,
		_w4435_
	);
	LUT2 #(
		.INIT('h2)
	) name3904 (
		\sa03_reg[2]/P0001 ,
		_w2293_,
		_w4436_
	);
	LUT2 #(
		.INIT('h4)
	) name3905 (
		_w4435_,
		_w4436_,
		_w4437_
	);
	LUT2 #(
		.INIT('h4)
	) name3906 (
		_w2685_,
		_w4437_,
		_w4438_
	);
	LUT2 #(
		.INIT('h1)
	) name3907 (
		\sa03_reg[2]/P0001 ,
		_w1416_,
		_w4439_
	);
	LUT2 #(
		.INIT('h4)
	) name3908 (
		_w1504_,
		_w4439_,
		_w4440_
	);
	LUT2 #(
		.INIT('h1)
	) name3909 (
		_w1400_,
		_w1572_,
		_w4441_
	);
	LUT2 #(
		.INIT('h8)
	) name3910 (
		_w4440_,
		_w4441_,
		_w4442_
	);
	LUT2 #(
		.INIT('h1)
	) name3911 (
		_w4438_,
		_w4442_,
		_w4443_
	);
	LUT2 #(
		.INIT('h1)
	) name3912 (
		_w4434_,
		_w4443_,
		_w4444_
	);
	LUT2 #(
		.INIT('h1)
	) name3913 (
		\sa03_reg[1]/P0001 ,
		_w4444_,
		_w4445_
	);
	LUT2 #(
		.INIT('h8)
	) name3914 (
		\sa03_reg[1]/P0001 ,
		_w1374_,
		_w4446_
	);
	LUT2 #(
		.INIT('h8)
	) name3915 (
		_w2200_,
		_w4446_,
		_w4447_
	);
	LUT2 #(
		.INIT('h4)
	) name3916 (
		_w4118_,
		_w4138_,
		_w4448_
	);
	LUT2 #(
		.INIT('h1)
	) name3917 (
		_w1397_,
		_w3830_,
		_w4449_
	);
	LUT2 #(
		.INIT('h2)
	) name3918 (
		\sa03_reg[2]/P0001 ,
		_w4449_,
		_w4450_
	);
	LUT2 #(
		.INIT('h8)
	) name3919 (
		\sa03_reg[4]/P0001 ,
		_w3692_,
		_w4451_
	);
	LUT2 #(
		.INIT('h2)
	) name3920 (
		_w3713_,
		_w4451_,
		_w4452_
	);
	LUT2 #(
		.INIT('h1)
	) name3921 (
		\sa03_reg[2]/P0001 ,
		_w4452_,
		_w4453_
	);
	LUT2 #(
		.INIT('h1)
	) name3922 (
		_w1328_,
		_w4450_,
		_w4454_
	);
	LUT2 #(
		.INIT('h4)
	) name3923 (
		_w4453_,
		_w4454_,
		_w4455_
	);
	LUT2 #(
		.INIT('h2)
	) name3924 (
		\sa03_reg[1]/P0001 ,
		_w4455_,
		_w4456_
	);
	LUT2 #(
		.INIT('h1)
	) name3925 (
		_w1383_,
		_w1398_,
		_w4457_
	);
	LUT2 #(
		.INIT('h1)
	) name3926 (
		\sa03_reg[2]/P0001 ,
		_w1449_,
		_w4458_
	);
	LUT2 #(
		.INIT('h4)
	) name3927 (
		_w4457_,
		_w4458_,
		_w4459_
	);
	LUT2 #(
		.INIT('h4)
	) name3928 (
		\sa03_reg[7]/NET0131 ,
		_w1408_,
		_w4460_
	);
	LUT2 #(
		.INIT('h1)
	) name3929 (
		_w1447_,
		_w4460_,
		_w4461_
	);
	LUT2 #(
		.INIT('h2)
	) name3930 (
		\sa03_reg[2]/P0001 ,
		_w4461_,
		_w4462_
	);
	LUT2 #(
		.INIT('h2)
	) name3931 (
		\sa03_reg[1]/P0001 ,
		_w1565_,
		_w4463_
	);
	LUT2 #(
		.INIT('h4)
	) name3932 (
		_w4459_,
		_w4463_,
		_w4464_
	);
	LUT2 #(
		.INIT('h4)
	) name3933 (
		_w4462_,
		_w4464_,
		_w4465_
	);
	LUT2 #(
		.INIT('h8)
	) name3934 (
		_w1429_,
		_w1449_,
		_w4466_
	);
	LUT2 #(
		.INIT('h1)
	) name3935 (
		\sa03_reg[1]/P0001 ,
		_w2293_,
		_w4467_
	);
	LUT2 #(
		.INIT('h4)
	) name3936 (
		_w4466_,
		_w4467_,
		_w4468_
	);
	LUT2 #(
		.INIT('h1)
	) name3937 (
		_w4465_,
		_w4468_,
		_w4469_
	);
	LUT2 #(
		.INIT('h4)
	) name3938 (
		\sa03_reg[2]/P0001 ,
		_w1417_,
		_w4470_
	);
	LUT2 #(
		.INIT('h8)
	) name3939 (
		\sa03_reg[2]/P0001 ,
		_w2249_,
		_w4471_
	);
	LUT2 #(
		.INIT('h1)
	) name3940 (
		\sa03_reg[0]/P0001 ,
		_w1365_,
		_w4472_
	);
	LUT2 #(
		.INIT('h4)
	) name3941 (
		_w4470_,
		_w4472_,
		_w4473_
	);
	LUT2 #(
		.INIT('h4)
	) name3942 (
		_w4471_,
		_w4473_,
		_w4474_
	);
	LUT2 #(
		.INIT('h4)
	) name3943 (
		_w4469_,
		_w4474_,
		_w4475_
	);
	LUT2 #(
		.INIT('h4)
	) name3944 (
		\sa03_reg[2]/P0001 ,
		_w1409_,
		_w4476_
	);
	LUT2 #(
		.INIT('h8)
	) name3945 (
		_w1318_,
		_w1436_,
		_w4477_
	);
	LUT2 #(
		.INIT('h1)
	) name3946 (
		_w1504_,
		_w2650_,
		_w4478_
	);
	LUT2 #(
		.INIT('h1)
	) name3947 (
		_w4102_,
		_w4477_,
		_w4479_
	);
	LUT2 #(
		.INIT('h8)
	) name3948 (
		_w4478_,
		_w4479_,
		_w4480_
	);
	LUT2 #(
		.INIT('h2)
	) name3949 (
		_w2656_,
		_w2715_,
		_w4481_
	);
	LUT2 #(
		.INIT('h4)
	) name3950 (
		_w4476_,
		_w4481_,
		_w4482_
	);
	LUT2 #(
		.INIT('h4)
	) name3951 (
		_w2707_,
		_w4480_,
		_w4483_
	);
	LUT2 #(
		.INIT('h8)
	) name3952 (
		_w4482_,
		_w4483_,
		_w4484_
	);
	LUT2 #(
		.INIT('h8)
	) name3953 (
		_w1383_,
		_w1384_,
		_w4485_
	);
	LUT2 #(
		.INIT('h8)
	) name3954 (
		_w1555_,
		_w3818_,
		_w4486_
	);
	LUT2 #(
		.INIT('h2)
	) name3955 (
		\sa03_reg[1]/P0001 ,
		_w4485_,
		_w4487_
	);
	LUT2 #(
		.INIT('h4)
	) name3956 (
		_w4486_,
		_w4487_,
		_w4488_
	);
	LUT2 #(
		.INIT('h4)
	) name3957 (
		_w4140_,
		_w4488_,
		_w4489_
	);
	LUT2 #(
		.INIT('h1)
	) name3958 (
		_w4484_,
		_w4489_,
		_w4490_
	);
	LUT2 #(
		.INIT('h8)
	) name3959 (
		_w1435_,
		_w1436_,
		_w4491_
	);
	LUT2 #(
		.INIT('h1)
	) name3960 (
		_w1353_,
		_w1414_,
		_w4492_
	);
	LUT2 #(
		.INIT('h4)
	) name3961 (
		_w1566_,
		_w4492_,
		_w4493_
	);
	LUT2 #(
		.INIT('h2)
	) name3962 (
		_w1374_,
		_w4493_,
		_w4494_
	);
	LUT2 #(
		.INIT('h2)
	) name3963 (
		\sa03_reg[0]/P0001 ,
		_w2676_,
		_w4495_
	);
	LUT2 #(
		.INIT('h1)
	) name3964 (
		_w2678_,
		_w4491_,
		_w4496_
	);
	LUT2 #(
		.INIT('h8)
	) name3965 (
		_w4495_,
		_w4496_,
		_w4497_
	);
	LUT2 #(
		.INIT('h4)
	) name3966 (
		_w4494_,
		_w4497_,
		_w4498_
	);
	LUT2 #(
		.INIT('h4)
	) name3967 (
		_w4490_,
		_w4498_,
		_w4499_
	);
	LUT2 #(
		.INIT('h1)
	) name3968 (
		_w4475_,
		_w4499_,
		_w4500_
	);
	LUT2 #(
		.INIT('h1)
	) name3969 (
		_w3845_,
		_w4447_,
		_w4501_
	);
	LUT2 #(
		.INIT('h4)
	) name3970 (
		_w4448_,
		_w4501_,
		_w4502_
	);
	LUT2 #(
		.INIT('h4)
	) name3971 (
		_w4445_,
		_w4502_,
		_w4503_
	);
	LUT2 #(
		.INIT('h4)
	) name3972 (
		_w4456_,
		_w4503_,
		_w4504_
	);
	LUT2 #(
		.INIT('h4)
	) name3973 (
		_w4500_,
		_w4504_,
		_w4505_
	);
	LUT2 #(
		.INIT('h2)
	) name3974 (
		_w4433_,
		_w4505_,
		_w4506_
	);
	LUT2 #(
		.INIT('h4)
	) name3975 (
		_w4433_,
		_w4505_,
		_w4507_
	);
	LUT2 #(
		.INIT('h1)
	) name3976 (
		_w4506_,
		_w4507_,
		_w4508_
	);
	LUT2 #(
		.INIT('h1)
	) name3977 (
		_w3768_,
		_w4508_,
		_w4509_
	);
	LUT2 #(
		.INIT('h8)
	) name3978 (
		_w3768_,
		_w4508_,
		_w4510_
	);
	LUT2 #(
		.INIT('h1)
	) name3979 (
		_w4509_,
		_w4510_,
		_w4511_
	);
	LUT2 #(
		.INIT('h1)
	) name3980 (
		_w2422_,
		_w2452_,
		_w4512_
	);
	LUT2 #(
		.INIT('h2)
	) name3981 (
		_w2453_,
		_w4512_,
		_w4513_
	);
	LUT2 #(
		.INIT('h2)
	) name3982 (
		_w1801_,
		_w1855_,
		_w4514_
	);
	LUT2 #(
		.INIT('h1)
	) name3983 (
		_w1880_,
		_w1889_,
		_w4515_
	);
	LUT2 #(
		.INIT('h8)
	) name3984 (
		_w4514_,
		_w4515_,
		_w4516_
	);
	LUT2 #(
		.INIT('h2)
	) name3985 (
		\sa21_reg[2]/P0001 ,
		_w2508_,
		_w4517_
	);
	LUT2 #(
		.INIT('h4)
	) name3986 (
		_w2857_,
		_w4517_,
		_w4518_
	);
	LUT2 #(
		.INIT('h4)
	) name3987 (
		_w3050_,
		_w4518_,
		_w4519_
	);
	LUT2 #(
		.INIT('h1)
	) name3988 (
		_w4516_,
		_w4519_,
		_w4520_
	);
	LUT2 #(
		.INIT('h1)
	) name3989 (
		\sa21_reg[1]/P0001 ,
		_w2993_,
		_w4521_
	);
	LUT2 #(
		.INIT('h4)
	) name3990 (
		_w2522_,
		_w4521_,
		_w4522_
	);
	LUT2 #(
		.INIT('h4)
	) name3991 (
		_w4520_,
		_w4522_,
		_w4523_
	);
	LUT2 #(
		.INIT('h8)
	) name3992 (
		_w1759_,
		_w1854_,
		_w4524_
	);
	LUT2 #(
		.INIT('h2)
	) name3993 (
		\sa21_reg[2]/P0001 ,
		_w1816_,
		_w4525_
	);
	LUT2 #(
		.INIT('h4)
	) name3994 (
		_w1834_,
		_w4525_,
		_w4526_
	);
	LUT2 #(
		.INIT('h4)
	) name3995 (
		_w4524_,
		_w4526_,
		_w4527_
	);
	LUT2 #(
		.INIT('h8)
	) name3996 (
		\sa21_reg[4]/P0001 ,
		_w3542_,
		_w4528_
	);
	LUT2 #(
		.INIT('h1)
	) name3997 (
		\sa21_reg[2]/P0001 ,
		_w4528_,
		_w4529_
	);
	LUT2 #(
		.INIT('h8)
	) name3998 (
		_w4196_,
		_w4529_,
		_w4530_
	);
	LUT2 #(
		.INIT('h1)
	) name3999 (
		_w4527_,
		_w4530_,
		_w4531_
	);
	LUT2 #(
		.INIT('h2)
	) name4000 (
		\sa21_reg[1]/P0001 ,
		_w2838_,
		_w4532_
	);
	LUT2 #(
		.INIT('h4)
	) name4001 (
		_w4531_,
		_w4532_,
		_w4533_
	);
	LUT2 #(
		.INIT('h1)
	) name4002 (
		_w4523_,
		_w4533_,
		_w4534_
	);
	LUT2 #(
		.INIT('h1)
	) name4003 (
		_w1781_,
		_w1884_,
		_w4535_
	);
	LUT2 #(
		.INIT('h4)
	) name4004 (
		_w2493_,
		_w4535_,
		_w4536_
	);
	LUT2 #(
		.INIT('h2)
	) name4005 (
		_w1894_,
		_w4536_,
		_w4537_
	);
	LUT2 #(
		.INIT('h8)
	) name4006 (
		_w1761_,
		_w1831_,
		_w4538_
	);
	LUT2 #(
		.INIT('h8)
	) name4007 (
		_w2437_,
		_w2479_,
		_w4539_
	);
	LUT2 #(
		.INIT('h1)
	) name4008 (
		\sa21_reg[1]/P0001 ,
		_w1800_,
		_w4540_
	);
	LUT2 #(
		.INIT('h1)
	) name4009 (
		_w3021_,
		_w3029_,
		_w4541_
	);
	LUT2 #(
		.INIT('h1)
	) name4010 (
		_w3545_,
		_w4538_,
		_w4542_
	);
	LUT2 #(
		.INIT('h8)
	) name4011 (
		_w4541_,
		_w4542_,
		_w4543_
	);
	LUT2 #(
		.INIT('h4)
	) name4012 (
		_w2900_,
		_w4540_,
		_w4544_
	);
	LUT2 #(
		.INIT('h1)
	) name4013 (
		_w2997_,
		_w4539_,
		_w4545_
	);
	LUT2 #(
		.INIT('h8)
	) name4014 (
		_w4544_,
		_w4545_,
		_w4546_
	);
	LUT2 #(
		.INIT('h8)
	) name4015 (
		_w4543_,
		_w4546_,
		_w4547_
	);
	LUT2 #(
		.INIT('h8)
	) name4016 (
		\sa21_reg[2]/P0001 ,
		_w2862_,
		_w4548_
	);
	LUT2 #(
		.INIT('h1)
	) name4017 (
		_w1844_,
		_w2450_,
		_w4549_
	);
	LUT2 #(
		.INIT('h1)
	) name4018 (
		\sa21_reg[2]/P0001 ,
		_w4549_,
		_w4550_
	);
	LUT2 #(
		.INIT('h2)
	) name4019 (
		\sa21_reg[1]/P0001 ,
		_w3572_,
		_w4551_
	);
	LUT2 #(
		.INIT('h4)
	) name4020 (
		_w4548_,
		_w4551_,
		_w4552_
	);
	LUT2 #(
		.INIT('h4)
	) name4021 (
		_w4550_,
		_w4552_,
		_w4553_
	);
	LUT2 #(
		.INIT('h1)
	) name4022 (
		_w4547_,
		_w4553_,
		_w4554_
	);
	LUT2 #(
		.INIT('h2)
	) name4023 (
		\sa21_reg[0]/P0001 ,
		_w3049_,
		_w4555_
	);
	LUT2 #(
		.INIT('h1)
	) name4024 (
		_w3055_,
		_w4176_,
		_w4556_
	);
	LUT2 #(
		.INIT('h8)
	) name4025 (
		_w4555_,
		_w4556_,
		_w4557_
	);
	LUT2 #(
		.INIT('h4)
	) name4026 (
		_w4537_,
		_w4557_,
		_w4558_
	);
	LUT2 #(
		.INIT('h4)
	) name4027 (
		_w4554_,
		_w4558_,
		_w4559_
	);
	LUT2 #(
		.INIT('h1)
	) name4028 (
		\sa21_reg[1]/P0001 ,
		_w2508_,
		_w4560_
	);
	LUT2 #(
		.INIT('h4)
	) name4029 (
		_w3571_,
		_w4560_,
		_w4561_
	);
	LUT2 #(
		.INIT('h1)
	) name4030 (
		_w1785_,
		_w4019_,
		_w4562_
	);
	LUT2 #(
		.INIT('h8)
	) name4031 (
		_w3555_,
		_w4562_,
		_w4563_
	);
	LUT2 #(
		.INIT('h2)
	) name4032 (
		\sa21_reg[2]/P0001 ,
		_w2437_,
		_w4564_
	);
	LUT2 #(
		.INIT('h4)
	) name4033 (
		_w2876_,
		_w4564_,
		_w4565_
	);
	LUT2 #(
		.INIT('h1)
	) name4034 (
		_w4563_,
		_w4565_,
		_w4566_
	);
	LUT2 #(
		.INIT('h2)
	) name4035 (
		\sa21_reg[1]/P0001 ,
		_w1885_,
		_w4567_
	);
	LUT2 #(
		.INIT('h4)
	) name4036 (
		_w4566_,
		_w4567_,
		_w4568_
	);
	LUT2 #(
		.INIT('h1)
	) name4037 (
		_w4561_,
		_w4568_,
		_w4569_
	);
	LUT2 #(
		.INIT('h8)
	) name4038 (
		\sa21_reg[2]/P0001 ,
		_w2465_,
		_w4570_
	);
	LUT2 #(
		.INIT('h1)
	) name4039 (
		\sa21_reg[0]/P0001 ,
		_w1792_,
		_w4571_
	);
	LUT2 #(
		.INIT('h4)
	) name4040 (
		_w1881_,
		_w4571_,
		_w4572_
	);
	LUT2 #(
		.INIT('h4)
	) name4041 (
		_w4570_,
		_w4572_,
		_w4573_
	);
	LUT2 #(
		.INIT('h4)
	) name4042 (
		_w4569_,
		_w4573_,
		_w4574_
	);
	LUT2 #(
		.INIT('h1)
	) name4043 (
		_w4559_,
		_w4574_,
		_w4575_
	);
	LUT2 #(
		.INIT('h1)
	) name4044 (
		_w4014_,
		_w4513_,
		_w4576_
	);
	LUT2 #(
		.INIT('h4)
	) name4045 (
		_w4534_,
		_w4576_,
		_w4577_
	);
	LUT2 #(
		.INIT('h4)
	) name4046 (
		_w4575_,
		_w4577_,
		_w4578_
	);
	LUT2 #(
		.INIT('h2)
	) name4047 (
		\u0_w_reg[3][2]/P0001 ,
		_w4578_,
		_w4579_
	);
	LUT2 #(
		.INIT('h4)
	) name4048 (
		\u0_w_reg[3][2]/P0001 ,
		_w4578_,
		_w4580_
	);
	LUT2 #(
		.INIT('h1)
	) name4049 (
		_w4579_,
		_w4580_,
		_w4581_
	);
	LUT2 #(
		.INIT('h8)
	) name4050 (
		_w3503_,
		_w4581_,
		_w4582_
	);
	LUT2 #(
		.INIT('h1)
	) name4051 (
		_w3503_,
		_w4581_,
		_w4583_
	);
	LUT2 #(
		.INIT('h1)
	) name4052 (
		_w4582_,
		_w4583_,
		_w4584_
	);
	LUT2 #(
		.INIT('h4)
	) name4053 (
		_w4511_,
		_w4584_,
		_w4585_
	);
	LUT2 #(
		.INIT('h2)
	) name4054 (
		_w4511_,
		_w4584_,
		_w4586_
	);
	LUT2 #(
		.INIT('h1)
	) name4055 (
		\ld_r_reg/P0001 ,
		_w4585_,
		_w4587_
	);
	LUT2 #(
		.INIT('h4)
	) name4056 (
		_w4586_,
		_w4587_,
		_w4588_
	);
	LUT2 #(
		.INIT('h1)
	) name4057 (
		\text_in_r_reg[2]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		_w4589_
	);
	LUT2 #(
		.INIT('h8)
	) name4058 (
		\text_in_r_reg[2]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		_w4590_
	);
	LUT2 #(
		.INIT('h2)
	) name4059 (
		\ld_r_reg/P0001 ,
		_w4589_,
		_w4591_
	);
	LUT2 #(
		.INIT('h4)
	) name4060 (
		_w4590_,
		_w4591_,
		_w4592_
	);
	LUT2 #(
		.INIT('h1)
	) name4061 (
		_w4588_,
		_w4592_,
		_w4593_
	);
	LUT2 #(
		.INIT('h2)
	) name4062 (
		_w3681_,
		_w4248_,
		_w4594_
	);
	LUT2 #(
		.INIT('h4)
	) name4063 (
		_w3681_,
		_w4248_,
		_w4595_
	);
	LUT2 #(
		.INIT('h1)
	) name4064 (
		_w4594_,
		_w4595_,
		_w4596_
	);
	LUT2 #(
		.INIT('h2)
	) name4065 (
		\u0_w_reg[3][25]/P0001 ,
		_w3503_,
		_w4597_
	);
	LUT2 #(
		.INIT('h4)
	) name4066 (
		\u0_w_reg[3][25]/P0001 ,
		_w3503_,
		_w4598_
	);
	LUT2 #(
		.INIT('h1)
	) name4067 (
		_w4597_,
		_w4598_,
		_w4599_
	);
	LUT2 #(
		.INIT('h8)
	) name4068 (
		_w4596_,
		_w4599_,
		_w4600_
	);
	LUT2 #(
		.INIT('h1)
	) name4069 (
		_w4596_,
		_w4599_,
		_w4601_
	);
	LUT2 #(
		.INIT('h1)
	) name4070 (
		_w4600_,
		_w4601_,
		_w4602_
	);
	LUT2 #(
		.INIT('h1)
	) name4071 (
		\sa10_reg[5]/P0001 ,
		_w1614_,
		_w4603_
	);
	LUT2 #(
		.INIT('h2)
	) name4072 (
		_w2142_,
		_w4603_,
		_w4604_
	);
	LUT2 #(
		.INIT('h1)
	) name4073 (
		_w1708_,
		_w4604_,
		_w4605_
	);
	LUT2 #(
		.INIT('h2)
	) name4074 (
		\sa10_reg[1]/P0001 ,
		_w4605_,
		_w4606_
	);
	LUT2 #(
		.INIT('h1)
	) name4075 (
		_w1586_,
		_w1672_,
		_w4607_
	);
	LUT2 #(
		.INIT('h2)
	) name4076 (
		\sa10_reg[3]/P0001 ,
		_w4607_,
		_w4608_
	);
	LUT2 #(
		.INIT('h1)
	) name4077 (
		_w2118_,
		_w2160_,
		_w4609_
	);
	LUT2 #(
		.INIT('h4)
	) name4078 (
		_w4608_,
		_w4609_,
		_w4610_
	);
	LUT2 #(
		.INIT('h1)
	) name4079 (
		\sa10_reg[2]/P0001 ,
		_w4610_,
		_w4611_
	);
	LUT2 #(
		.INIT('h1)
	) name4080 (
		_w2625_,
		_w2748_,
		_w4612_
	);
	LUT2 #(
		.INIT('h8)
	) name4081 (
		_w1632_,
		_w4612_,
		_w4613_
	);
	LUT2 #(
		.INIT('h2)
	) name4082 (
		\sa10_reg[2]/P0001 ,
		_w4613_,
		_w4614_
	);
	LUT2 #(
		.INIT('h8)
	) name4083 (
		\sa10_reg[4]/P0001 ,
		_w2155_,
		_w4615_
	);
	LUT2 #(
		.INIT('h1)
	) name4084 (
		_w2168_,
		_w2634_,
		_w4616_
	);
	LUT2 #(
		.INIT('h2)
	) name4085 (
		\sa10_reg[2]/P0001 ,
		_w4616_,
		_w4617_
	);
	LUT2 #(
		.INIT('h1)
	) name4086 (
		_w2113_,
		_w2740_,
		_w4618_
	);
	LUT2 #(
		.INIT('h1)
	) name4087 (
		\sa10_reg[3]/P0001 ,
		_w4618_,
		_w4619_
	);
	LUT2 #(
		.INIT('h2)
	) name4088 (
		\sa10_reg[5]/P0001 ,
		_w1597_,
		_w4620_
	);
	LUT2 #(
		.INIT('h2)
	) name4089 (
		_w1627_,
		_w4620_,
		_w4621_
	);
	LUT2 #(
		.INIT('h1)
	) name4090 (
		_w4615_,
		_w4621_,
		_w4622_
	);
	LUT2 #(
		.INIT('h4)
	) name4091 (
		_w4619_,
		_w4622_,
		_w4623_
	);
	LUT2 #(
		.INIT('h4)
	) name4092 (
		_w4617_,
		_w4623_,
		_w4624_
	);
	LUT2 #(
		.INIT('h1)
	) name4093 (
		\sa10_reg[1]/P0001 ,
		_w4624_,
		_w4625_
	);
	LUT2 #(
		.INIT('h1)
	) name4094 (
		_w2554_,
		_w3599_,
		_w4626_
	);
	LUT2 #(
		.INIT('h4)
	) name4095 (
		_w4606_,
		_w4626_,
		_w4627_
	);
	LUT2 #(
		.INIT('h4)
	) name4096 (
		_w4611_,
		_w4627_,
		_w4628_
	);
	LUT2 #(
		.INIT('h4)
	) name4097 (
		_w4614_,
		_w4628_,
		_w4629_
	);
	LUT2 #(
		.INIT('h4)
	) name4098 (
		_w4625_,
		_w4629_,
		_w4630_
	);
	LUT2 #(
		.INIT('h2)
	) name4099 (
		\sa10_reg[0]/P0001 ,
		_w4630_,
		_w4631_
	);
	LUT2 #(
		.INIT('h1)
	) name4100 (
		\sa10_reg[3]/P0001 ,
		_w2094_,
		_w4632_
	);
	LUT2 #(
		.INIT('h2)
	) name4101 (
		_w2592_,
		_w4632_,
		_w4633_
	);
	LUT2 #(
		.INIT('h8)
	) name4102 (
		_w1664_,
		_w2621_,
		_w4634_
	);
	LUT2 #(
		.INIT('h1)
	) name4103 (
		_w1594_,
		_w1614_,
		_w4635_
	);
	LUT2 #(
		.INIT('h1)
	) name4104 (
		_w3624_,
		_w4635_,
		_w4636_
	);
	LUT2 #(
		.INIT('h2)
	) name4105 (
		\sa10_reg[1]/P0001 ,
		_w2154_,
		_w4637_
	);
	LUT2 #(
		.INIT('h4)
	) name4106 (
		_w4634_,
		_w4637_,
		_w4638_
	);
	LUT2 #(
		.INIT('h4)
	) name4107 (
		_w4636_,
		_w4638_,
		_w4639_
	);
	LUT2 #(
		.INIT('h1)
	) name4108 (
		_w4633_,
		_w4639_,
		_w4640_
	);
	LUT2 #(
		.INIT('h8)
	) name4109 (
		_w1650_,
		_w1668_,
		_w4641_
	);
	LUT2 #(
		.INIT('h2)
	) name4110 (
		_w3940_,
		_w4641_,
		_w4642_
	);
	LUT2 #(
		.INIT('h1)
	) name4111 (
		\sa10_reg[2]/P0001 ,
		_w4642_,
		_w4643_
	);
	LUT2 #(
		.INIT('h1)
	) name4112 (
		_w1615_,
		_w1672_,
		_w4644_
	);
	LUT2 #(
		.INIT('h2)
	) name4113 (
		_w1715_,
		_w4644_,
		_w4645_
	);
	LUT2 #(
		.INIT('h8)
	) name4114 (
		\sa10_reg[7]/NET0131 ,
		_w2183_,
		_w4646_
	);
	LUT2 #(
		.INIT('h8)
	) name4115 (
		_w3615_,
		_w4646_,
		_w4647_
	);
	LUT2 #(
		.INIT('h1)
	) name4116 (
		_w4645_,
		_w4647_,
		_w4648_
	);
	LUT2 #(
		.INIT('h4)
	) name4117 (
		_w4640_,
		_w4648_,
		_w4649_
	);
	LUT2 #(
		.INIT('h4)
	) name4118 (
		_w4643_,
		_w4649_,
		_w4650_
	);
	LUT2 #(
		.INIT('h1)
	) name4119 (
		\sa10_reg[0]/P0001 ,
		_w4650_,
		_w4651_
	);
	LUT2 #(
		.INIT('h1)
	) name4120 (
		_w2148_,
		_w2787_,
		_w4652_
	);
	LUT2 #(
		.INIT('h4)
	) name4121 (
		_w2572_,
		_w4652_,
		_w4653_
	);
	LUT2 #(
		.INIT('h1)
	) name4122 (
		\sa10_reg[2]/P0001 ,
		_w4653_,
		_w4654_
	);
	LUT2 #(
		.INIT('h1)
	) name4123 (
		_w2807_,
		_w4378_,
		_w4655_
	);
	LUT2 #(
		.INIT('h4)
	) name4124 (
		_w4654_,
		_w4655_,
		_w4656_
	);
	LUT2 #(
		.INIT('h1)
	) name4125 (
		\sa10_reg[1]/P0001 ,
		_w4656_,
		_w4657_
	);
	LUT2 #(
		.INIT('h8)
	) name4126 (
		\sa10_reg[6]/NET0131 ,
		_w1667_,
		_w4658_
	);
	LUT2 #(
		.INIT('h1)
	) name4127 (
		_w1730_,
		_w2577_,
		_w4659_
	);
	LUT2 #(
		.INIT('h1)
	) name4128 (
		\sa10_reg[5]/P0001 ,
		_w4659_,
		_w4660_
	);
	LUT2 #(
		.INIT('h1)
	) name4129 (
		\sa10_reg[2]/P0001 ,
		_w2189_,
		_w4661_
	);
	LUT2 #(
		.INIT('h1)
	) name4130 (
		_w2602_,
		_w4661_,
		_w4662_
	);
	LUT2 #(
		.INIT('h1)
	) name4131 (
		_w1727_,
		_w4662_,
		_w4663_
	);
	LUT2 #(
		.INIT('h4)
	) name4132 (
		_w4660_,
		_w4663_,
		_w4664_
	);
	LUT2 #(
		.INIT('h2)
	) name4133 (
		\sa10_reg[1]/P0001 ,
		_w4664_,
		_w4665_
	);
	LUT2 #(
		.INIT('h1)
	) name4134 (
		_w1711_,
		_w2559_,
		_w4666_
	);
	LUT2 #(
		.INIT('h2)
	) name4135 (
		\sa10_reg[1]/P0001 ,
		_w2179_,
		_w4667_
	);
	LUT2 #(
		.INIT('h2)
	) name4136 (
		\sa10_reg[2]/P0001 ,
		_w4666_,
		_w4668_
	);
	LUT2 #(
		.INIT('h4)
	) name4137 (
		_w4667_,
		_w4668_,
		_w4669_
	);
	LUT2 #(
		.INIT('h1)
	) name4138 (
		_w4658_,
		_w4669_,
		_w4670_
	);
	LUT2 #(
		.INIT('h4)
	) name4139 (
		_w4665_,
		_w4670_,
		_w4671_
	);
	LUT2 #(
		.INIT('h4)
	) name4140 (
		_w4657_,
		_w4671_,
		_w4672_
	);
	LUT2 #(
		.INIT('h4)
	) name4141 (
		_w4651_,
		_w4672_,
		_w4673_
	);
	LUT2 #(
		.INIT('h4)
	) name4142 (
		_w4631_,
		_w4673_,
		_w4674_
	);
	LUT2 #(
		.INIT('h2)
	) name4143 (
		_w4161_,
		_w4674_,
		_w4675_
	);
	LUT2 #(
		.INIT('h4)
	) name4144 (
		_w4161_,
		_w4674_,
		_w4676_
	);
	LUT2 #(
		.INIT('h1)
	) name4145 (
		_w4675_,
		_w4676_,
		_w4677_
	);
	LUT2 #(
		.INIT('h4)
	) name4146 (
		_w2307_,
		_w4677_,
		_w4678_
	);
	LUT2 #(
		.INIT('h2)
	) name4147 (
		_w2307_,
		_w4677_,
		_w4679_
	);
	LUT2 #(
		.INIT('h1)
	) name4148 (
		_w4678_,
		_w4679_,
		_w4680_
	);
	LUT2 #(
		.INIT('h1)
	) name4149 (
		_w4602_,
		_w4680_,
		_w4681_
	);
	LUT2 #(
		.INIT('h8)
	) name4150 (
		_w4602_,
		_w4680_,
		_w4682_
	);
	LUT2 #(
		.INIT('h1)
	) name4151 (
		\ld_r_reg/P0001 ,
		_w4681_,
		_w4683_
	);
	LUT2 #(
		.INIT('h4)
	) name4152 (
		_w4682_,
		_w4683_,
		_w4684_
	);
	LUT2 #(
		.INIT('h1)
	) name4153 (
		\text_in_r_reg[25]/P0001 ,
		\u0_w_reg[3][25]/P0001 ,
		_w4685_
	);
	LUT2 #(
		.INIT('h8)
	) name4154 (
		\text_in_r_reg[25]/P0001 ,
		\u0_w_reg[3][25]/P0001 ,
		_w4686_
	);
	LUT2 #(
		.INIT('h2)
	) name4155 (
		\ld_r_reg/P0001 ,
		_w4685_,
		_w4687_
	);
	LUT2 #(
		.INIT('h4)
	) name4156 (
		_w4686_,
		_w4687_,
		_w4688_
	);
	LUT2 #(
		.INIT('h1)
	) name4157 (
		_w4684_,
		_w4688_,
		_w4689_
	);
	LUT2 #(
		.INIT('h1)
	) name4158 (
		_w1908_,
		_w2307_,
		_w4690_
	);
	LUT2 #(
		.INIT('h8)
	) name4159 (
		_w1908_,
		_w2307_,
		_w4691_
	);
	LUT2 #(
		.INIT('h1)
	) name4160 (
		_w4690_,
		_w4691_,
		_w4692_
	);
	LUT2 #(
		.INIT('h2)
	) name4161 (
		\u0_w_reg[3][15]/P0001 ,
		_w3416_,
		_w4693_
	);
	LUT2 #(
		.INIT('h4)
	) name4162 (
		\u0_w_reg[3][15]/P0001 ,
		_w3416_,
		_w4694_
	);
	LUT2 #(
		.INIT('h1)
	) name4163 (
		_w4693_,
		_w4694_,
		_w4695_
	);
	LUT2 #(
		.INIT('h8)
	) name4164 (
		_w2416_,
		_w4695_,
		_w4696_
	);
	LUT2 #(
		.INIT('h1)
	) name4165 (
		_w2416_,
		_w4695_,
		_w4697_
	);
	LUT2 #(
		.INIT('h1)
	) name4166 (
		_w4696_,
		_w4697_,
		_w4698_
	);
	LUT2 #(
		.INIT('h1)
	) name4167 (
		_w4692_,
		_w4698_,
		_w4699_
	);
	LUT2 #(
		.INIT('h8)
	) name4168 (
		_w4692_,
		_w4698_,
		_w4700_
	);
	LUT2 #(
		.INIT('h1)
	) name4169 (
		\ld_r_reg/P0001 ,
		_w4699_,
		_w4701_
	);
	LUT2 #(
		.INIT('h4)
	) name4170 (
		_w4700_,
		_w4701_,
		_w4702_
	);
	LUT2 #(
		.INIT('h2)
	) name4171 (
		\text_in_r_reg[15]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w4703_
	);
	LUT2 #(
		.INIT('h4)
	) name4172 (
		\text_in_r_reg[15]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w4704_
	);
	LUT2 #(
		.INIT('h2)
	) name4173 (
		\ld_r_reg/P0001 ,
		_w4703_,
		_w4705_
	);
	LUT2 #(
		.INIT('h4)
	) name4174 (
		_w4704_,
		_w4705_,
		_w4706_
	);
	LUT2 #(
		.INIT('h1)
	) name4175 (
		_w4702_,
		_w4706_,
		_w4707_
	);
	LUT2 #(
		.INIT('h2)
	) name4176 (
		_w2304_,
		_w3888_,
		_w4708_
	);
	LUT2 #(
		.INIT('h4)
	) name4177 (
		_w2304_,
		_w3888_,
		_w4709_
	);
	LUT2 #(
		.INIT('h1)
	) name4178 (
		_w4708_,
		_w4709_,
		_w4710_
	);
	LUT2 #(
		.INIT('h8)
	) name4179 (
		_w2739_,
		_w4710_,
		_w4711_
	);
	LUT2 #(
		.INIT('h1)
	) name4180 (
		_w2739_,
		_w4710_,
		_w4712_
	);
	LUT2 #(
		.INIT('h1)
	) name4181 (
		_w4711_,
		_w4712_,
		_w4713_
	);
	LUT2 #(
		.INIT('h2)
	) name4182 (
		\u0_w_reg[3][4]/P0001 ,
		_w3069_,
		_w4714_
	);
	LUT2 #(
		.INIT('h4)
	) name4183 (
		\u0_w_reg[3][4]/P0001 ,
		_w3069_,
		_w4715_
	);
	LUT2 #(
		.INIT('h1)
	) name4184 (
		_w4714_,
		_w4715_,
		_w4716_
	);
	LUT2 #(
		.INIT('h8)
	) name4185 (
		_w4341_,
		_w4716_,
		_w4717_
	);
	LUT2 #(
		.INIT('h1)
	) name4186 (
		_w4341_,
		_w4716_,
		_w4718_
	);
	LUT2 #(
		.INIT('h1)
	) name4187 (
		_w4717_,
		_w4718_,
		_w4719_
	);
	LUT2 #(
		.INIT('h1)
	) name4188 (
		_w4713_,
		_w4719_,
		_w4720_
	);
	LUT2 #(
		.INIT('h8)
	) name4189 (
		_w4713_,
		_w4719_,
		_w4721_
	);
	LUT2 #(
		.INIT('h1)
	) name4190 (
		\ld_r_reg/P0001 ,
		_w4720_,
		_w4722_
	);
	LUT2 #(
		.INIT('h4)
	) name4191 (
		_w4721_,
		_w4722_,
		_w4723_
	);
	LUT2 #(
		.INIT('h2)
	) name4192 (
		\text_in_r_reg[4]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w4724_
	);
	LUT2 #(
		.INIT('h4)
	) name4193 (
		\text_in_r_reg[4]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w4725_
	);
	LUT2 #(
		.INIT('h2)
	) name4194 (
		\ld_r_reg/P0001 ,
		_w4724_,
		_w4726_
	);
	LUT2 #(
		.INIT('h4)
	) name4195 (
		_w4725_,
		_w4726_,
		_w4727_
	);
	LUT2 #(
		.INIT('h1)
	) name4196 (
		_w4723_,
		_w4727_,
		_w4728_
	);
	LUT2 #(
		.INIT('h2)
	) name4197 (
		\u0_w_reg[3][27]/P0001 ,
		_w4338_,
		_w4729_
	);
	LUT2 #(
		.INIT('h4)
	) name4198 (
		\u0_w_reg[3][27]/P0001 ,
		_w4338_,
		_w4730_
	);
	LUT2 #(
		.INIT('h1)
	) name4199 (
		_w4729_,
		_w4730_,
		_w4731_
	);
	LUT2 #(
		.INIT('h8)
	) name4200 (
		_w4062_,
		_w4731_,
		_w4732_
	);
	LUT2 #(
		.INIT('h1)
	) name4201 (
		_w4062_,
		_w4731_,
		_w4733_
	);
	LUT2 #(
		.INIT('h1)
	) name4202 (
		_w4732_,
		_w4733_,
		_w4734_
	);
	LUT2 #(
		.INIT('h4)
	) name4203 (
		_w2307_,
		_w4508_,
		_w4735_
	);
	LUT2 #(
		.INIT('h2)
	) name4204 (
		_w2307_,
		_w4508_,
		_w4736_
	);
	LUT2 #(
		.INIT('h1)
	) name4205 (
		_w4735_,
		_w4736_,
		_w4737_
	);
	LUT2 #(
		.INIT('h2)
	) name4206 (
		_w4734_,
		_w4737_,
		_w4738_
	);
	LUT2 #(
		.INIT('h4)
	) name4207 (
		_w4734_,
		_w4737_,
		_w4739_
	);
	LUT2 #(
		.INIT('h1)
	) name4208 (
		\ld_r_reg/P0001 ,
		_w4738_,
		_w4740_
	);
	LUT2 #(
		.INIT('h4)
	) name4209 (
		_w4739_,
		_w4740_,
		_w4741_
	);
	LUT2 #(
		.INIT('h2)
	) name4210 (
		\text_in_r_reg[27]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w4742_
	);
	LUT2 #(
		.INIT('h4)
	) name4211 (
		\text_in_r_reg[27]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w4743_
	);
	LUT2 #(
		.INIT('h2)
	) name4212 (
		\ld_r_reg/P0001 ,
		_w4742_,
		_w4744_
	);
	LUT2 #(
		.INIT('h4)
	) name4213 (
		_w4743_,
		_w4744_,
		_w4745_
	);
	LUT2 #(
		.INIT('h1)
	) name4214 (
		_w4741_,
		_w4745_,
		_w4746_
	);
	LUT2 #(
		.INIT('h2)
	) name4215 (
		\u0_w_reg[3][19]/P0001 ,
		_w4338_,
		_w4747_
	);
	LUT2 #(
		.INIT('h4)
	) name4216 (
		\u0_w_reg[3][19]/P0001 ,
		_w4338_,
		_w4748_
	);
	LUT2 #(
		.INIT('h1)
	) name4217 (
		_w4747_,
		_w4748_,
		_w4749_
	);
	LUT2 #(
		.INIT('h8)
	) name4218 (
		_w4350_,
		_w4749_,
		_w4750_
	);
	LUT2 #(
		.INIT('h1)
	) name4219 (
		_w4350_,
		_w4749_,
		_w4751_
	);
	LUT2 #(
		.INIT('h1)
	) name4220 (
		_w4750_,
		_w4751_,
		_w4752_
	);
	LUT2 #(
		.INIT('h2)
	) name4221 (
		_w4433_,
		_w4578_,
		_w4753_
	);
	LUT2 #(
		.INIT('h4)
	) name4222 (
		_w4433_,
		_w4578_,
		_w4754_
	);
	LUT2 #(
		.INIT('h1)
	) name4223 (
		_w4753_,
		_w4754_,
		_w4755_
	);
	LUT2 #(
		.INIT('h2)
	) name4224 (
		_w2199_,
		_w3888_,
		_w4756_
	);
	LUT2 #(
		.INIT('h4)
	) name4225 (
		_w2199_,
		_w3888_,
		_w4757_
	);
	LUT2 #(
		.INIT('h1)
	) name4226 (
		_w4756_,
		_w4757_,
		_w4758_
	);
	LUT2 #(
		.INIT('h8)
	) name4227 (
		_w4755_,
		_w4758_,
		_w4759_
	);
	LUT2 #(
		.INIT('h1)
	) name4228 (
		_w4755_,
		_w4758_,
		_w4760_
	);
	LUT2 #(
		.INIT('h1)
	) name4229 (
		_w4759_,
		_w4760_,
		_w4761_
	);
	LUT2 #(
		.INIT('h1)
	) name4230 (
		_w4752_,
		_w4761_,
		_w4762_
	);
	LUT2 #(
		.INIT('h8)
	) name4231 (
		_w4752_,
		_w4761_,
		_w4763_
	);
	LUT2 #(
		.INIT('h1)
	) name4232 (
		\ld_r_reg/P0001 ,
		_w4762_,
		_w4764_
	);
	LUT2 #(
		.INIT('h4)
	) name4233 (
		_w4763_,
		_w4764_,
		_w4765_
	);
	LUT2 #(
		.INIT('h2)
	) name4234 (
		\text_in_r_reg[19]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w4766_
	);
	LUT2 #(
		.INIT('h4)
	) name4235 (
		\text_in_r_reg[19]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w4767_
	);
	LUT2 #(
		.INIT('h2)
	) name4236 (
		\ld_r_reg/P0001 ,
		_w4766_,
		_w4768_
	);
	LUT2 #(
		.INIT('h4)
	) name4237 (
		_w4767_,
		_w4768_,
		_w4769_
	);
	LUT2 #(
		.INIT('h1)
	) name4238 (
		_w4765_,
		_w4769_,
		_w4770_
	);
	LUT2 #(
		.INIT('h2)
	) name4239 (
		_w3592_,
		_w4674_,
		_w4771_
	);
	LUT2 #(
		.INIT('h4)
	) name4240 (
		_w3592_,
		_w4674_,
		_w4772_
	);
	LUT2 #(
		.INIT('h1)
	) name4241 (
		_w4771_,
		_w4772_,
		_w4773_
	);
	LUT2 #(
		.INIT('h2)
	) name4242 (
		_w2199_,
		_w3768_,
		_w4774_
	);
	LUT2 #(
		.INIT('h4)
	) name4243 (
		_w2199_,
		_w3768_,
		_w4775_
	);
	LUT2 #(
		.INIT('h1)
	) name4244 (
		_w4774_,
		_w4775_,
		_w4776_
	);
	LUT2 #(
		.INIT('h8)
	) name4245 (
		_w4773_,
		_w4776_,
		_w4777_
	);
	LUT2 #(
		.INIT('h1)
	) name4246 (
		_w4773_,
		_w4776_,
		_w4778_
	);
	LUT2 #(
		.INIT('h1)
	) name4247 (
		_w4777_,
		_w4778_,
		_w4779_
	);
	LUT2 #(
		.INIT('h1)
	) name4248 (
		_w2529_,
		_w3503_,
		_w4780_
	);
	LUT2 #(
		.INIT('h8)
	) name4249 (
		_w2529_,
		_w3503_,
		_w4781_
	);
	LUT2 #(
		.INIT('h1)
	) name4250 (
		_w4780_,
		_w4781_,
		_w4782_
	);
	LUT2 #(
		.INIT('h2)
	) name4251 (
		\u0_w_reg[3][17]/P0001 ,
		_w4248_,
		_w4783_
	);
	LUT2 #(
		.INIT('h4)
	) name4252 (
		\u0_w_reg[3][17]/P0001 ,
		_w4248_,
		_w4784_
	);
	LUT2 #(
		.INIT('h1)
	) name4253 (
		_w4783_,
		_w4784_,
		_w4785_
	);
	LUT2 #(
		.INIT('h8)
	) name4254 (
		_w4782_,
		_w4785_,
		_w4786_
	);
	LUT2 #(
		.INIT('h1)
	) name4255 (
		_w4782_,
		_w4785_,
		_w4787_
	);
	LUT2 #(
		.INIT('h1)
	) name4256 (
		_w4786_,
		_w4787_,
		_w4788_
	);
	LUT2 #(
		.INIT('h1)
	) name4257 (
		_w4779_,
		_w4788_,
		_w4789_
	);
	LUT2 #(
		.INIT('h8)
	) name4258 (
		_w4779_,
		_w4788_,
		_w4790_
	);
	LUT2 #(
		.INIT('h1)
	) name4259 (
		\ld_r_reg/P0001 ,
		_w4789_,
		_w4791_
	);
	LUT2 #(
		.INIT('h4)
	) name4260 (
		_w4790_,
		_w4791_,
		_w4792_
	);
	LUT2 #(
		.INIT('h1)
	) name4261 (
		\text_in_r_reg[17]/P0001 ,
		\u0_w_reg[3][17]/P0001 ,
		_w4793_
	);
	LUT2 #(
		.INIT('h8)
	) name4262 (
		\text_in_r_reg[17]/P0001 ,
		\u0_w_reg[3][17]/P0001 ,
		_w4794_
	);
	LUT2 #(
		.INIT('h2)
	) name4263 (
		\ld_r_reg/P0001 ,
		_w4793_,
		_w4795_
	);
	LUT2 #(
		.INIT('h4)
	) name4264 (
		_w4794_,
		_w4795_,
		_w4796_
	);
	LUT2 #(
		.INIT('h1)
	) name4265 (
		_w4792_,
		_w4796_,
		_w4797_
	);
	LUT2 #(
		.INIT('h2)
	) name4266 (
		_w2529_,
		_w4578_,
		_w4798_
	);
	LUT2 #(
		.INIT('h4)
	) name4267 (
		_w2529_,
		_w4578_,
		_w4799_
	);
	LUT2 #(
		.INIT('h1)
	) name4268 (
		_w4798_,
		_w4799_,
		_w4800_
	);
	LUT2 #(
		.INIT('h8)
	) name4269 (
		_w3969_,
		_w4800_,
		_w4801_
	);
	LUT2 #(
		.INIT('h1)
	) name4270 (
		_w3969_,
		_w4800_,
		_w4802_
	);
	LUT2 #(
		.INIT('h1)
	) name4271 (
		_w4801_,
		_w4802_,
		_w4803_
	);
	LUT2 #(
		.INIT('h4)
	) name4272 (
		\sa32_reg[4]/P0001 ,
		_w2366_,
		_w4804_
	);
	LUT2 #(
		.INIT('h1)
	) name4273 (
		_w1963_,
		_w2050_,
		_w4805_
	);
	LUT2 #(
		.INIT('h4)
	) name4274 (
		_w4804_,
		_w4805_,
		_w4806_
	);
	LUT2 #(
		.INIT('h2)
	) name4275 (
		\sa32_reg[2]/P0001 ,
		_w4806_,
		_w4807_
	);
	LUT2 #(
		.INIT('h4)
	) name4276 (
		_w2006_,
		_w3451_,
		_w4808_
	);
	LUT2 #(
		.INIT('h1)
	) name4277 (
		\sa32_reg[2]/P0001 ,
		_w4808_,
		_w4809_
	);
	LUT2 #(
		.INIT('h2)
	) name4278 (
		\sa32_reg[1]/P0001 ,
		_w1989_,
		_w4810_
	);
	LUT2 #(
		.INIT('h4)
	) name4279 (
		_w4807_,
		_w4810_,
		_w4811_
	);
	LUT2 #(
		.INIT('h4)
	) name4280 (
		_w4809_,
		_w4811_,
		_w4812_
	);
	LUT2 #(
		.INIT('h1)
	) name4281 (
		_w1919_,
		_w1948_,
		_w4813_
	);
	LUT2 #(
		.INIT('h8)
	) name4282 (
		_w1990_,
		_w4813_,
		_w4814_
	);
	LUT2 #(
		.INIT('h1)
	) name4283 (
		_w2356_,
		_w3405_,
		_w4815_
	);
	LUT2 #(
		.INIT('h4)
	) name4284 (
		_w2052_,
		_w4815_,
		_w4816_
	);
	LUT2 #(
		.INIT('h8)
	) name4285 (
		_w2333_,
		_w4816_,
		_w4817_
	);
	LUT2 #(
		.INIT('h1)
	) name4286 (
		_w1991_,
		_w3134_,
		_w4818_
	);
	LUT2 #(
		.INIT('h8)
	) name4287 (
		_w3388_,
		_w4818_,
		_w4819_
	);
	LUT2 #(
		.INIT('h1)
	) name4288 (
		_w4817_,
		_w4819_,
		_w4820_
	);
	LUT2 #(
		.INIT('h1)
	) name4289 (
		\sa32_reg[1]/P0001 ,
		_w4814_,
		_w4821_
	);
	LUT2 #(
		.INIT('h4)
	) name4290 (
		_w4820_,
		_w4821_,
		_w4822_
	);
	LUT2 #(
		.INIT('h1)
	) name4291 (
		_w4812_,
		_w4822_,
		_w4823_
	);
	LUT2 #(
		.INIT('h1)
	) name4292 (
		_w2060_,
		_w2387_,
		_w4824_
	);
	LUT2 #(
		.INIT('h4)
	) name4293 (
		\sa32_reg[3]/P0001 ,
		_w2348_,
		_w4825_
	);
	LUT2 #(
		.INIT('h4)
	) name4294 (
		_w4824_,
		_w4825_,
		_w4826_
	);
	LUT2 #(
		.INIT('h1)
	) name4295 (
		_w2011_,
		_w2351_,
		_w4827_
	);
	LUT2 #(
		.INIT('h4)
	) name4296 (
		_w3331_,
		_w4827_,
		_w4828_
	);
	LUT2 #(
		.INIT('h2)
	) name4297 (
		_w2059_,
		_w4828_,
		_w4829_
	);
	LUT2 #(
		.INIT('h4)
	) name4298 (
		_w1924_,
		_w2067_,
		_w4830_
	);
	LUT2 #(
		.INIT('h4)
	) name4299 (
		\sa32_reg[2]/P0001 ,
		_w2040_,
		_w4831_
	);
	LUT2 #(
		.INIT('h1)
	) name4300 (
		_w3184_,
		_w3257_,
		_w4832_
	);
	LUT2 #(
		.INIT('h4)
	) name4301 (
		_w1964_,
		_w4832_,
		_w4833_
	);
	LUT2 #(
		.INIT('h4)
	) name4302 (
		_w2332_,
		_w3173_,
		_w4834_
	);
	LUT2 #(
		.INIT('h1)
	) name4303 (
		_w4830_,
		_w4831_,
		_w4835_
	);
	LUT2 #(
		.INIT('h8)
	) name4304 (
		_w4834_,
		_w4835_,
		_w4836_
	);
	LUT2 #(
		.INIT('h8)
	) name4305 (
		_w4833_,
		_w4836_,
		_w4837_
	);
	LUT2 #(
		.INIT('h1)
	) name4306 (
		\sa32_reg[2]/P0001 ,
		_w1947_,
		_w4838_
	);
	LUT2 #(
		.INIT('h8)
	) name4307 (
		_w3363_,
		_w4838_,
		_w4839_
	);
	LUT2 #(
		.INIT('h2)
	) name4308 (
		\sa32_reg[1]/P0001 ,
		_w2349_,
		_w4840_
	);
	LUT2 #(
		.INIT('h4)
	) name4309 (
		_w3309_,
		_w4840_,
		_w4841_
	);
	LUT2 #(
		.INIT('h4)
	) name4310 (
		_w4839_,
		_w4841_,
		_w4842_
	);
	LUT2 #(
		.INIT('h1)
	) name4311 (
		_w4837_,
		_w4842_,
		_w4843_
	);
	LUT2 #(
		.INIT('h1)
	) name4312 (
		_w2068_,
		_w3146_,
		_w4844_
	);
	LUT2 #(
		.INIT('h1)
	) name4313 (
		\sa32_reg[3]/P0001 ,
		_w4844_,
		_w4845_
	);
	LUT2 #(
		.INIT('h2)
	) name4314 (
		\sa32_reg[0]/P0002 ,
		_w3126_,
		_w4846_
	);
	LUT2 #(
		.INIT('h4)
	) name4315 (
		_w4845_,
		_w4846_,
		_w4847_
	);
	LUT2 #(
		.INIT('h4)
	) name4316 (
		_w4829_,
		_w4847_,
		_w4848_
	);
	LUT2 #(
		.INIT('h4)
	) name4317 (
		_w4843_,
		_w4848_,
		_w4849_
	);
	LUT2 #(
		.INIT('h1)
	) name4318 (
		_w1947_,
		_w1948_,
		_w4850_
	);
	LUT2 #(
		.INIT('h1)
	) name4319 (
		\sa32_reg[2]/P0001 ,
		_w1934_,
		_w4851_
	);
	LUT2 #(
		.INIT('h4)
	) name4320 (
		_w4850_,
		_w4851_,
		_w4852_
	);
	LUT2 #(
		.INIT('h1)
	) name4321 (
		_w1949_,
		_w3376_,
		_w4853_
	);
	LUT2 #(
		.INIT('h2)
	) name4322 (
		\sa32_reg[2]/P0001 ,
		_w4853_,
		_w4854_
	);
	LUT2 #(
		.INIT('h2)
	) name4323 (
		\sa32_reg[1]/P0001 ,
		_w2352_,
		_w4855_
	);
	LUT2 #(
		.INIT('h4)
	) name4324 (
		_w4852_,
		_w4855_,
		_w4856_
	);
	LUT2 #(
		.INIT('h4)
	) name4325 (
		_w4854_,
		_w4856_,
		_w4857_
	);
	LUT2 #(
		.INIT('h1)
	) name4326 (
		\sa32_reg[1]/P0001 ,
		_w1921_,
		_w4858_
	);
	LUT2 #(
		.INIT('h4)
	) name4327 (
		_w3308_,
		_w4858_,
		_w4859_
	);
	LUT2 #(
		.INIT('h1)
	) name4328 (
		_w4857_,
		_w4859_,
		_w4860_
	);
	LUT2 #(
		.INIT('h8)
	) name4329 (
		\sa32_reg[6]/NET0131 ,
		_w3326_,
		_w4861_
	);
	LUT2 #(
		.INIT('h1)
	) name4330 (
		\sa32_reg[0]/P0002 ,
		_w2024_,
		_w4862_
	);
	LUT2 #(
		.INIT('h4)
	) name4331 (
		_w2368_,
		_w4862_,
		_w4863_
	);
	LUT2 #(
		.INIT('h4)
	) name4332 (
		_w4861_,
		_w4863_,
		_w4864_
	);
	LUT2 #(
		.INIT('h4)
	) name4333 (
		_w4860_,
		_w4864_,
		_w4865_
	);
	LUT2 #(
		.INIT('h1)
	) name4334 (
		_w4849_,
		_w4865_,
		_w4866_
	);
	LUT2 #(
		.INIT('h1)
	) name4335 (
		_w4317_,
		_w4826_,
		_w4867_
	);
	LUT2 #(
		.INIT('h4)
	) name4336 (
		_w4823_,
		_w4867_,
		_w4868_
	);
	LUT2 #(
		.INIT('h4)
	) name4337 (
		_w4866_,
		_w4868_,
		_w4869_
	);
	LUT2 #(
		.INIT('h2)
	) name4338 (
		\u0_w_reg[3][11]/P0001 ,
		_w4869_,
		_w4870_
	);
	LUT2 #(
		.INIT('h4)
	) name4339 (
		\u0_w_reg[3][11]/P0001 ,
		_w4869_,
		_w4871_
	);
	LUT2 #(
		.INIT('h1)
	) name4340 (
		_w4870_,
		_w4871_,
		_w4872_
	);
	LUT2 #(
		.INIT('h8)
	) name4341 (
		_w4341_,
		_w4872_,
		_w4873_
	);
	LUT2 #(
		.INIT('h1)
	) name4342 (
		_w4341_,
		_w4872_,
		_w4874_
	);
	LUT2 #(
		.INIT('h1)
	) name4343 (
		_w4873_,
		_w4874_,
		_w4875_
	);
	LUT2 #(
		.INIT('h1)
	) name4344 (
		_w4803_,
		_w4875_,
		_w4876_
	);
	LUT2 #(
		.INIT('h8)
	) name4345 (
		_w4803_,
		_w4875_,
		_w4877_
	);
	LUT2 #(
		.INIT('h1)
	) name4346 (
		\ld_r_reg/P0001 ,
		_w4876_,
		_w4878_
	);
	LUT2 #(
		.INIT('h4)
	) name4347 (
		_w4877_,
		_w4878_,
		_w4879_
	);
	LUT2 #(
		.INIT('h2)
	) name4348 (
		\text_in_r_reg[11]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w4880_
	);
	LUT2 #(
		.INIT('h4)
	) name4349 (
		\text_in_r_reg[11]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w4881_
	);
	LUT2 #(
		.INIT('h2)
	) name4350 (
		\ld_r_reg/P0001 ,
		_w4880_,
		_w4882_
	);
	LUT2 #(
		.INIT('h4)
	) name4351 (
		_w4881_,
		_w4882_,
		_w4883_
	);
	LUT2 #(
		.INIT('h1)
	) name4352 (
		_w4879_,
		_w4883_,
		_w4884_
	);
	LUT2 #(
		.INIT('h2)
	) name4353 (
		\u0_w_reg[3][26]/P0001 ,
		_w4869_,
		_w4885_
	);
	LUT2 #(
		.INIT('h4)
	) name4354 (
		\u0_w_reg[3][26]/P0001 ,
		_w4869_,
		_w4886_
	);
	LUT2 #(
		.INIT('h1)
	) name4355 (
		_w4885_,
		_w4886_,
		_w4887_
	);
	LUT2 #(
		.INIT('h8)
	) name4356 (
		_w4755_,
		_w4887_,
		_w4888_
	);
	LUT2 #(
		.INIT('h1)
	) name4357 (
		_w4755_,
		_w4887_,
		_w4889_
	);
	LUT2 #(
		.INIT('h1)
	) name4358 (
		_w4888_,
		_w4889_,
		_w4890_
	);
	LUT2 #(
		.INIT('h1)
	) name4359 (
		_w3771_,
		_w4890_,
		_w4891_
	);
	LUT2 #(
		.INIT('h8)
	) name4360 (
		_w3771_,
		_w4890_,
		_w4892_
	);
	LUT2 #(
		.INIT('h1)
	) name4361 (
		\ld_r_reg/P0001 ,
		_w4891_,
		_w4893_
	);
	LUT2 #(
		.INIT('h4)
	) name4362 (
		_w4892_,
		_w4893_,
		_w4894_
	);
	LUT2 #(
		.INIT('h2)
	) name4363 (
		\text_in_r_reg[26]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		_w4895_
	);
	LUT2 #(
		.INIT('h4)
	) name4364 (
		\text_in_r_reg[26]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		_w4896_
	);
	LUT2 #(
		.INIT('h2)
	) name4365 (
		\ld_r_reg/P0001 ,
		_w4895_,
		_w4897_
	);
	LUT2 #(
		.INIT('h4)
	) name4366 (
		_w4896_,
		_w4897_,
		_w4898_
	);
	LUT2 #(
		.INIT('h1)
	) name4367 (
		_w4894_,
		_w4898_,
		_w4899_
	);
	LUT2 #(
		.INIT('h2)
	) name4368 (
		_w2304_,
		_w4505_,
		_w4900_
	);
	LUT2 #(
		.INIT('h4)
	) name4369 (
		_w2304_,
		_w4505_,
		_w4901_
	);
	LUT2 #(
		.INIT('h1)
	) name4370 (
		_w4900_,
		_w4901_,
		_w4902_
	);
	LUT2 #(
		.INIT('h8)
	) name4371 (
		_w3969_,
		_w4902_,
		_w4903_
	);
	LUT2 #(
		.INIT('h1)
	) name4372 (
		_w3969_,
		_w4902_,
		_w4904_
	);
	LUT2 #(
		.INIT('h1)
	) name4373 (
		_w4903_,
		_w4904_,
		_w4905_
	);
	LUT2 #(
		.INIT('h1)
	) name4374 (
		_w3416_,
		_w4059_,
		_w4906_
	);
	LUT2 #(
		.INIT('h8)
	) name4375 (
		_w3416_,
		_w4059_,
		_w4907_
	);
	LUT2 #(
		.INIT('h1)
	) name4376 (
		_w4906_,
		_w4907_,
		_w4908_
	);
	LUT2 #(
		.INIT('h2)
	) name4377 (
		\u0_w_reg[3][3]/P0001 ,
		_w4869_,
		_w4909_
	);
	LUT2 #(
		.INIT('h4)
	) name4378 (
		\u0_w_reg[3][3]/P0001 ,
		_w4869_,
		_w4910_
	);
	LUT2 #(
		.INIT('h1)
	) name4379 (
		_w4909_,
		_w4910_,
		_w4911_
	);
	LUT2 #(
		.INIT('h8)
	) name4380 (
		_w4908_,
		_w4911_,
		_w4912_
	);
	LUT2 #(
		.INIT('h1)
	) name4381 (
		_w4908_,
		_w4911_,
		_w4913_
	);
	LUT2 #(
		.INIT('h1)
	) name4382 (
		_w4912_,
		_w4913_,
		_w4914_
	);
	LUT2 #(
		.INIT('h2)
	) name4383 (
		_w4905_,
		_w4914_,
		_w4915_
	);
	LUT2 #(
		.INIT('h4)
	) name4384 (
		_w4905_,
		_w4914_,
		_w4916_
	);
	LUT2 #(
		.INIT('h1)
	) name4385 (
		\ld_r_reg/P0001 ,
		_w4915_,
		_w4917_
	);
	LUT2 #(
		.INIT('h4)
	) name4386 (
		_w4916_,
		_w4917_,
		_w4918_
	);
	LUT2 #(
		.INIT('h2)
	) name4387 (
		\text_in_r_reg[3]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w4919_
	);
	LUT2 #(
		.INIT('h4)
	) name4388 (
		\text_in_r_reg[3]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w4920_
	);
	LUT2 #(
		.INIT('h2)
	) name4389 (
		\ld_r_reg/P0001 ,
		_w4919_,
		_w4921_
	);
	LUT2 #(
		.INIT('h4)
	) name4390 (
		_w4920_,
		_w4921_,
		_w4922_
	);
	LUT2 #(
		.INIT('h1)
	) name4391 (
		_w4918_,
		_w4922_,
		_w4923_
	);
	LUT2 #(
		.INIT('h1)
	) name4392 (
		\u0_w_reg[3][24]/P0001 ,
		_w3325_,
		_w4924_
	);
	LUT2 #(
		.INIT('h8)
	) name4393 (
		\u0_w_reg[3][24]/P0001 ,
		_w3325_,
		_w4925_
	);
	LUT2 #(
		.INIT('h1)
	) name4394 (
		_w4924_,
		_w4925_,
		_w4926_
	);
	LUT2 #(
		.INIT('h4)
	) name4395 (
		_w2307_,
		_w4773_,
		_w4927_
	);
	LUT2 #(
		.INIT('h2)
	) name4396 (
		_w2307_,
		_w4773_,
		_w4928_
	);
	LUT2 #(
		.INIT('h1)
	) name4397 (
		_w4927_,
		_w4928_,
		_w4929_
	);
	LUT2 #(
		.INIT('h1)
	) name4398 (
		_w4926_,
		_w4929_,
		_w4930_
	);
	LUT2 #(
		.INIT('h8)
	) name4399 (
		_w4926_,
		_w4929_,
		_w4931_
	);
	LUT2 #(
		.INIT('h1)
	) name4400 (
		\ld_r_reg/P0001 ,
		_w4930_,
		_w4932_
	);
	LUT2 #(
		.INIT('h4)
	) name4401 (
		_w4931_,
		_w4932_,
		_w4933_
	);
	LUT2 #(
		.INIT('h1)
	) name4402 (
		\text_in_r_reg[24]/P0001 ,
		\u0_w_reg[3][24]/P0001 ,
		_w4934_
	);
	LUT2 #(
		.INIT('h8)
	) name4403 (
		\text_in_r_reg[24]/P0001 ,
		\u0_w_reg[3][24]/P0001 ,
		_w4935_
	);
	LUT2 #(
		.INIT('h2)
	) name4404 (
		\ld_r_reg/P0001 ,
		_w4934_,
		_w4936_
	);
	LUT2 #(
		.INIT('h4)
	) name4405 (
		_w4935_,
		_w4936_,
		_w4937_
	);
	LUT2 #(
		.INIT('h1)
	) name4406 (
		_w4933_,
		_w4937_,
		_w4938_
	);
	LUT2 #(
		.INIT('h2)
	) name4407 (
		_w2529_,
		_w3416_,
		_w4939_
	);
	LUT2 #(
		.INIT('h4)
	) name4408 (
		_w2529_,
		_w3416_,
		_w4940_
	);
	LUT2 #(
		.INIT('h1)
	) name4409 (
		_w4939_,
		_w4940_,
		_w4941_
	);
	LUT2 #(
		.INIT('h2)
	) name4410 (
		\u0_w_reg[3][31]/P0001 ,
		_w2199_,
		_w4942_
	);
	LUT2 #(
		.INIT('h4)
	) name4411 (
		\u0_w_reg[3][31]/P0001 ,
		_w2199_,
		_w4943_
	);
	LUT2 #(
		.INIT('h1)
	) name4412 (
		_w4942_,
		_w4943_,
		_w4944_
	);
	LUT2 #(
		.INIT('h8)
	) name4413 (
		_w4941_,
		_w4944_,
		_w4945_
	);
	LUT2 #(
		.INIT('h1)
	) name4414 (
		_w4941_,
		_w4944_,
		_w4946_
	);
	LUT2 #(
		.INIT('h1)
	) name4415 (
		_w4945_,
		_w4946_,
		_w4947_
	);
	LUT2 #(
		.INIT('h4)
	) name4416 (
		_w1741_,
		_w4947_,
		_w4948_
	);
	LUT2 #(
		.INIT('h2)
	) name4417 (
		_w1741_,
		_w4947_,
		_w4949_
	);
	LUT2 #(
		.INIT('h1)
	) name4418 (
		\ld_r_reg/P0001 ,
		_w4948_,
		_w4950_
	);
	LUT2 #(
		.INIT('h4)
	) name4419 (
		_w4949_,
		_w4950_,
		_w4951_
	);
	LUT2 #(
		.INIT('h1)
	) name4420 (
		\text_in_r_reg[31]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w4952_
	);
	LUT2 #(
		.INIT('h8)
	) name4421 (
		\text_in_r_reg[31]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w4953_
	);
	LUT2 #(
		.INIT('h2)
	) name4422 (
		\ld_r_reg/P0001 ,
		_w4952_,
		_w4954_
	);
	LUT2 #(
		.INIT('h4)
	) name4423 (
		_w4953_,
		_w4954_,
		_w4955_
	);
	LUT2 #(
		.INIT('h1)
	) name4424 (
		_w4951_,
		_w4955_,
		_w4956_
	);
	LUT2 #(
		.INIT('h1)
	) name4425 (
		\u0_w_reg[3][16]/P0001 ,
		_w3325_,
		_w4957_
	);
	LUT2 #(
		.INIT('h8)
	) name4426 (
		\u0_w_reg[3][16]/P0001 ,
		_w3325_,
		_w4958_
	);
	LUT2 #(
		.INIT('h1)
	) name4427 (
		_w4957_,
		_w4958_,
		_w4959_
	);
	LUT2 #(
		.INIT('h2)
	) name4428 (
		_w2199_,
		_w4161_,
		_w4960_
	);
	LUT2 #(
		.INIT('h4)
	) name4429 (
		_w2199_,
		_w4161_,
		_w4961_
	);
	LUT2 #(
		.INIT('h1)
	) name4430 (
		_w4960_,
		_w4961_,
		_w4962_
	);
	LUT2 #(
		.INIT('h8)
	) name4431 (
		_w3595_,
		_w4962_,
		_w4963_
	);
	LUT2 #(
		.INIT('h1)
	) name4432 (
		_w3595_,
		_w4962_,
		_w4964_
	);
	LUT2 #(
		.INIT('h1)
	) name4433 (
		_w4963_,
		_w4964_,
		_w4965_
	);
	LUT2 #(
		.INIT('h4)
	) name4434 (
		_w4959_,
		_w4965_,
		_w4966_
	);
	LUT2 #(
		.INIT('h2)
	) name4435 (
		_w4959_,
		_w4965_,
		_w4967_
	);
	LUT2 #(
		.INIT('h1)
	) name4436 (
		\ld_r_reg/P0001 ,
		_w4966_,
		_w4968_
	);
	LUT2 #(
		.INIT('h4)
	) name4437 (
		_w4967_,
		_w4968_,
		_w4969_
	);
	LUT2 #(
		.INIT('h1)
	) name4438 (
		\text_in_r_reg[16]/P0001 ,
		\u0_w_reg[3][16]/P0001 ,
		_w4970_
	);
	LUT2 #(
		.INIT('h8)
	) name4439 (
		\text_in_r_reg[16]/P0001 ,
		\u0_w_reg[3][16]/P0001 ,
		_w4971_
	);
	LUT2 #(
		.INIT('h2)
	) name4440 (
		\ld_r_reg/P0001 ,
		_w4970_,
		_w4972_
	);
	LUT2 #(
		.INIT('h4)
	) name4441 (
		_w4971_,
		_w4972_,
		_w4973_
	);
	LUT2 #(
		.INIT('h1)
	) name4442 (
		_w4969_,
		_w4973_,
		_w4974_
	);
	LUT2 #(
		.INIT('h1)
	) name4443 (
		_w4505_,
		_w4596_,
		_w4975_
	);
	LUT2 #(
		.INIT('h8)
	) name4444 (
		_w4505_,
		_w4596_,
		_w4976_
	);
	LUT2 #(
		.INIT('h1)
	) name4445 (
		_w4975_,
		_w4976_,
		_w4977_
	);
	LUT2 #(
		.INIT('h2)
	) name4446 (
		\u0_w_reg[3][18]/P0001 ,
		_w4869_,
		_w4978_
	);
	LUT2 #(
		.INIT('h4)
	) name4447 (
		\u0_w_reg[3][18]/P0001 ,
		_w4869_,
		_w4979_
	);
	LUT2 #(
		.INIT('h1)
	) name4448 (
		_w4978_,
		_w4979_,
		_w4980_
	);
	LUT2 #(
		.INIT('h8)
	) name4449 (
		_w4578_,
		_w4980_,
		_w4981_
	);
	LUT2 #(
		.INIT('h1)
	) name4450 (
		_w4578_,
		_w4980_,
		_w4982_
	);
	LUT2 #(
		.INIT('h1)
	) name4451 (
		_w4981_,
		_w4982_,
		_w4983_
	);
	LUT2 #(
		.INIT('h1)
	) name4452 (
		_w4977_,
		_w4983_,
		_w4984_
	);
	LUT2 #(
		.INIT('h8)
	) name4453 (
		_w4977_,
		_w4983_,
		_w4985_
	);
	LUT2 #(
		.INIT('h1)
	) name4454 (
		\ld_r_reg/P0001 ,
		_w4984_,
		_w4986_
	);
	LUT2 #(
		.INIT('h4)
	) name4455 (
		_w4985_,
		_w4986_,
		_w4987_
	);
	LUT2 #(
		.INIT('h2)
	) name4456 (
		\text_in_r_reg[18]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		_w4988_
	);
	LUT2 #(
		.INIT('h4)
	) name4457 (
		\text_in_r_reg[18]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		_w4989_
	);
	LUT2 #(
		.INIT('h2)
	) name4458 (
		\ld_r_reg/P0001 ,
		_w4988_,
		_w4990_
	);
	LUT2 #(
		.INIT('h4)
	) name4459 (
		_w4989_,
		_w4990_,
		_w4991_
	);
	LUT2 #(
		.INIT('h1)
	) name4460 (
		_w4987_,
		_w4991_,
		_w4992_
	);
	LUT2 #(
		.INIT('h1)
	) name4461 (
		_w2304_,
		_w2960_,
		_w4993_
	);
	LUT2 #(
		.INIT('h8)
	) name4462 (
		_w2304_,
		_w2960_,
		_w4994_
	);
	LUT2 #(
		.INIT('h1)
	) name4463 (
		_w4993_,
		_w4994_,
		_w4995_
	);
	LUT2 #(
		.INIT('h1)
	) name4464 (
		\u0_w_reg[3][23]/P0001 ,
		_w4941_,
		_w4996_
	);
	LUT2 #(
		.INIT('h8)
	) name4465 (
		\u0_w_reg[3][23]/P0001 ,
		_w4941_,
		_w4997_
	);
	LUT2 #(
		.INIT('h1)
	) name4466 (
		_w4996_,
		_w4997_,
		_w4998_
	);
	LUT2 #(
		.INIT('h1)
	) name4467 (
		_w4995_,
		_w4998_,
		_w4999_
	);
	LUT2 #(
		.INIT('h8)
	) name4468 (
		_w4995_,
		_w4998_,
		_w5000_
	);
	LUT2 #(
		.INIT('h1)
	) name4469 (
		\ld_r_reg/P0001 ,
		_w4999_,
		_w5001_
	);
	LUT2 #(
		.INIT('h4)
	) name4470 (
		_w5000_,
		_w5001_,
		_w5002_
	);
	LUT2 #(
		.INIT('h2)
	) name4471 (
		\text_in_r_reg[23]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w5003_
	);
	LUT2 #(
		.INIT('h4)
	) name4472 (
		\text_in_r_reg[23]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w5004_
	);
	LUT2 #(
		.INIT('h2)
	) name4473 (
		\ld_r_reg/P0001 ,
		_w5003_,
		_w5005_
	);
	LUT2 #(
		.INIT('h4)
	) name4474 (
		_w5004_,
		_w5005_,
		_w5006_
	);
	LUT2 #(
		.INIT('h1)
	) name4475 (
		_w5002_,
		_w5006_,
		_w5007_
	);
	LUT2 #(
		.INIT('h1)
	) name4476 (
		_w4248_,
		_w4508_,
		_w5008_
	);
	LUT2 #(
		.INIT('h8)
	) name4477 (
		_w4248_,
		_w4508_,
		_w5009_
	);
	LUT2 #(
		.INIT('h1)
	) name4478 (
		_w5008_,
		_w5009_,
		_w5010_
	);
	LUT2 #(
		.INIT('h2)
	) name4479 (
		\u0_w_reg[3][10]/P0001 ,
		_w4869_,
		_w5011_
	);
	LUT2 #(
		.INIT('h4)
	) name4480 (
		\u0_w_reg[3][10]/P0001 ,
		_w4869_,
		_w5012_
	);
	LUT2 #(
		.INIT('h1)
	) name4481 (
		_w5011_,
		_w5012_,
		_w5013_
	);
	LUT2 #(
		.INIT('h8)
	) name4482 (
		_w3503_,
		_w5013_,
		_w5014_
	);
	LUT2 #(
		.INIT('h1)
	) name4483 (
		_w3503_,
		_w5013_,
		_w5015_
	);
	LUT2 #(
		.INIT('h1)
	) name4484 (
		_w5014_,
		_w5015_,
		_w5016_
	);
	LUT2 #(
		.INIT('h1)
	) name4485 (
		_w5010_,
		_w5016_,
		_w5017_
	);
	LUT2 #(
		.INIT('h8)
	) name4486 (
		_w5010_,
		_w5016_,
		_w5018_
	);
	LUT2 #(
		.INIT('h1)
	) name4487 (
		\ld_r_reg/P0001 ,
		_w5017_,
		_w5019_
	);
	LUT2 #(
		.INIT('h4)
	) name4488 (
		_w5018_,
		_w5019_,
		_w5020_
	);
	LUT2 #(
		.INIT('h2)
	) name4489 (
		\text_in_r_reg[10]/P0001 ,
		\u0_w_reg[3][10]/P0001 ,
		_w5021_
	);
	LUT2 #(
		.INIT('h4)
	) name4490 (
		\text_in_r_reg[10]/P0001 ,
		\u0_w_reg[3][10]/P0001 ,
		_w5022_
	);
	LUT2 #(
		.INIT('h2)
	) name4491 (
		\ld_r_reg/P0001 ,
		_w5021_,
		_w5023_
	);
	LUT2 #(
		.INIT('h4)
	) name4492 (
		_w5022_,
		_w5023_,
		_w5024_
	);
	LUT2 #(
		.INIT('h1)
	) name4493 (
		_w5020_,
		_w5024_,
		_w5025_
	);
	LUT2 #(
		.INIT('h1)
	) name4494 (
		\u0_w_reg[3][8]/P0001 ,
		_w3325_,
		_w5026_
	);
	LUT2 #(
		.INIT('h8)
	) name4495 (
		\u0_w_reg[3][8]/P0001 ,
		_w3325_,
		_w5027_
	);
	LUT2 #(
		.INIT('h1)
	) name4496 (
		_w5026_,
		_w5027_,
		_w5028_
	);
	LUT2 #(
		.INIT('h2)
	) name4497 (
		_w4677_,
		_w4941_,
		_w5029_
	);
	LUT2 #(
		.INIT('h4)
	) name4498 (
		_w4677_,
		_w4941_,
		_w5030_
	);
	LUT2 #(
		.INIT('h1)
	) name4499 (
		_w5029_,
		_w5030_,
		_w5031_
	);
	LUT2 #(
		.INIT('h4)
	) name4500 (
		_w5028_,
		_w5031_,
		_w5032_
	);
	LUT2 #(
		.INIT('h2)
	) name4501 (
		_w5028_,
		_w5031_,
		_w5033_
	);
	LUT2 #(
		.INIT('h1)
	) name4502 (
		\ld_r_reg/P0001 ,
		_w5032_,
		_w5034_
	);
	LUT2 #(
		.INIT('h4)
	) name4503 (
		_w5033_,
		_w5034_,
		_w5035_
	);
	LUT2 #(
		.INIT('h2)
	) name4504 (
		\text_in_r_reg[8]/P0001 ,
		\u0_w_reg[3][8]/P0001 ,
		_w5036_
	);
	LUT2 #(
		.INIT('h4)
	) name4505 (
		\text_in_r_reg[8]/P0001 ,
		\u0_w_reg[3][8]/P0001 ,
		_w5037_
	);
	LUT2 #(
		.INIT('h2)
	) name4506 (
		\ld_r_reg/P0001 ,
		_w5036_,
		_w5038_
	);
	LUT2 #(
		.INIT('h4)
	) name4507 (
		_w5037_,
		_w5038_,
		_w5039_
	);
	LUT2 #(
		.INIT('h1)
	) name4508 (
		_w5035_,
		_w5039_,
		_w5040_
	);
	LUT2 #(
		.INIT('h1)
	) name4509 (
		\u0_w_reg[3][0]/P0001 ,
		_w3416_,
		_w5041_
	);
	LUT2 #(
		.INIT('h8)
	) name4510 (
		\u0_w_reg[3][0]/P0001 ,
		_w3416_,
		_w5042_
	);
	LUT2 #(
		.INIT('h1)
	) name4511 (
		_w5041_,
		_w5042_,
		_w5043_
	);
	LUT2 #(
		.INIT('h8)
	) name4512 (
		_w4164_,
		_w4773_,
		_w5044_
	);
	LUT2 #(
		.INIT('h1)
	) name4513 (
		_w4164_,
		_w4773_,
		_w5045_
	);
	LUT2 #(
		.INIT('h1)
	) name4514 (
		_w5044_,
		_w5045_,
		_w5046_
	);
	LUT2 #(
		.INIT('h1)
	) name4515 (
		_w5043_,
		_w5046_,
		_w5047_
	);
	LUT2 #(
		.INIT('h8)
	) name4516 (
		_w5043_,
		_w5046_,
		_w5048_
	);
	LUT2 #(
		.INIT('h1)
	) name4517 (
		\ld_r_reg/P0001 ,
		_w5047_,
		_w5049_
	);
	LUT2 #(
		.INIT('h4)
	) name4518 (
		_w5048_,
		_w5049_,
		_w5050_
	);
	LUT2 #(
		.INIT('h1)
	) name4519 (
		\text_in_r_reg[0]/P0001 ,
		\u0_w_reg[3][0]/P0001 ,
		_w5051_
	);
	LUT2 #(
		.INIT('h8)
	) name4520 (
		\text_in_r_reg[0]/P0001 ,
		\u0_w_reg[3][0]/P0001 ,
		_w5052_
	);
	LUT2 #(
		.INIT('h2)
	) name4521 (
		\ld_r_reg/P0001 ,
		_w5051_,
		_w5053_
	);
	LUT2 #(
		.INIT('h4)
	) name4522 (
		_w5052_,
		_w5053_,
		_w5054_
	);
	LUT2 #(
		.INIT('h1)
	) name4523 (
		_w5050_,
		_w5054_,
		_w5055_
	);
	LUT2 #(
		.INIT('h1)
	) name4524 (
		\u0_w_reg[3][5]/P0001 ,
		_w2077_,
		_w5056_
	);
	LUT2 #(
		.INIT('h8)
	) name4525 (
		\u0_w_reg[3][5]/P0001 ,
		_w2077_,
		_w5057_
	);
	LUT2 #(
		.INIT('h1)
	) name4526 (
		_w5056_,
		_w5057_,
		_w5058_
	);
	LUT2 #(
		.INIT('h1)
	) name4527 (
		\u0_w_reg[3][6]/P0001 ,
		_w2416_,
		_w5059_
	);
	LUT2 #(
		.INIT('h8)
	) name4528 (
		\u0_w_reg[3][6]/P0001 ,
		_w2416_,
		_w5060_
	);
	LUT2 #(
		.INIT('h1)
	) name4529 (
		_w5059_,
		_w5060_,
		_w5061_
	);
	LUT2 #(
		.INIT('h1)
	) name4530 (
		\u0_w_reg[3][4]/P0001 ,
		_w3205_,
		_w5062_
	);
	LUT2 #(
		.INIT('h8)
	) name4531 (
		\u0_w_reg[3][4]/P0001 ,
		_w3205_,
		_w5063_
	);
	LUT2 #(
		.INIT('h1)
	) name4532 (
		_w5062_,
		_w5063_,
		_w5064_
	);
	LUT2 #(
		.INIT('h1)
	) name4533 (
		\u0_w_reg[3][0]/P0001 ,
		_w3325_,
		_w5065_
	);
	LUT2 #(
		.INIT('h8)
	) name4534 (
		\u0_w_reg[3][0]/P0001 ,
		_w3325_,
		_w5066_
	);
	LUT2 #(
		.INIT('h1)
	) name4535 (
		_w5065_,
		_w5066_,
		_w5067_
	);
	LUT2 #(
		.INIT('h1)
	) name4536 (
		\u0_w_reg[3][3]/P0001 ,
		_w4338_,
		_w5068_
	);
	LUT2 #(
		.INIT('h8)
	) name4537 (
		\u0_w_reg[3][3]/P0001 ,
		_w4338_,
		_w5069_
	);
	LUT2 #(
		.INIT('h1)
	) name4538 (
		_w5068_,
		_w5069_,
		_w5070_
	);
	LUT2 #(
		.INIT('h1)
	) name4539 (
		\u0_w_reg[3][1]/P0001 ,
		_w3503_,
		_w5071_
	);
	LUT2 #(
		.INIT('h8)
	) name4540 (
		\u0_w_reg[3][1]/P0001 ,
		_w3503_,
		_w5072_
	);
	LUT2 #(
		.INIT('h1)
	) name4541 (
		_w5071_,
		_w5072_,
		_w5073_
	);
	LUT2 #(
		.INIT('h1)
	) name4542 (
		\u0_w_reg[3][2]/P0001 ,
		_w4869_,
		_w5074_
	);
	LUT2 #(
		.INIT('h8)
	) name4543 (
		\u0_w_reg[3][2]/P0001 ,
		_w4869_,
		_w5075_
	);
	LUT2 #(
		.INIT('h1)
	) name4544 (
		_w5074_,
		_w5075_,
		_w5076_
	);
	LUT2 #(
		.INIT('h1)
	) name4545 (
		\u0_w_reg[3][7]/P0001 ,
		_w3416_,
		_w5077_
	);
	LUT2 #(
		.INIT('h8)
	) name4546 (
		\u0_w_reg[3][7]/P0001 ,
		_w3416_,
		_w5078_
	);
	LUT2 #(
		.INIT('h1)
	) name4547 (
		_w5077_,
		_w5078_,
		_w5079_
	);
	LUT2 #(
		.INIT('h1)
	) name4548 (
		_w1071_,
		_w1123_,
		_w5080_
	);
	LUT2 #(
		.INIT('h8)
	) name4549 (
		_w982_,
		_w1015_,
		_w5081_
	);
	LUT2 #(
		.INIT('h8)
	) name4550 (
		\sa02_reg[4]/P0001 ,
		_w1025_,
		_w5082_
	);
	LUT2 #(
		.INIT('h4)
	) name4551 (
		\sa02_reg[3]/P0001 ,
		_w1090_,
		_w5083_
	);
	LUT2 #(
		.INIT('h8)
	) name4552 (
		\sa02_reg[7]/NET0131 ,
		_w5083_,
		_w5084_
	);
	LUT2 #(
		.INIT('h1)
	) name4553 (
		_w1043_,
		_w5082_,
		_w5085_
	);
	LUT2 #(
		.INIT('h4)
	) name4554 (
		_w5084_,
		_w5085_,
		_w5086_
	);
	LUT2 #(
		.INIT('h2)
	) name4555 (
		\sa02_reg[1]/P0001 ,
		_w5086_,
		_w5087_
	);
	LUT2 #(
		.INIT('h2)
	) name4556 (
		_w5080_,
		_w5081_,
		_w5088_
	);
	LUT2 #(
		.INIT('h4)
	) name4557 (
		_w5087_,
		_w5088_,
		_w5089_
	);
	LUT2 #(
		.INIT('h2)
	) name4558 (
		\sa02_reg[2]/P0001 ,
		_w5089_,
		_w5090_
	);
	LUT2 #(
		.INIT('h8)
	) name4559 (
		\sa02_reg[5]/P0001 ,
		_w979_,
		_w5091_
	);
	LUT2 #(
		.INIT('h4)
	) name4560 (
		\sa02_reg[3]/P0001 ,
		_w5091_,
		_w5092_
	);
	LUT2 #(
		.INIT('h2)
	) name4561 (
		_w1009_,
		_w5092_,
		_w5093_
	);
	LUT2 #(
		.INIT('h1)
	) name4562 (
		\sa02_reg[2]/P0001 ,
		_w5093_,
		_w5094_
	);
	LUT2 #(
		.INIT('h1)
	) name4563 (
		_w1001_,
		_w5094_,
		_w5095_
	);
	LUT2 #(
		.INIT('h1)
	) name4564 (
		\sa02_reg[1]/P0001 ,
		_w5095_,
		_w5096_
	);
	LUT2 #(
		.INIT('h2)
	) name4565 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		_w5097_
	);
	LUT2 #(
		.INIT('h8)
	) name4566 (
		_w1024_,
		_w5097_,
		_w5098_
	);
	LUT2 #(
		.INIT('h8)
	) name4567 (
		_w975_,
		_w1015_,
		_w5099_
	);
	LUT2 #(
		.INIT('h1)
	) name4568 (
		_w1022_,
		_w5099_,
		_w5100_
	);
	LUT2 #(
		.INIT('h1)
	) name4569 (
		\sa02_reg[2]/P0001 ,
		_w5100_,
		_w5101_
	);
	LUT2 #(
		.INIT('h8)
	) name4570 (
		_w993_,
		_w1059_,
		_w5102_
	);
	LUT2 #(
		.INIT('h1)
	) name4571 (
		_w1058_,
		_w5102_,
		_w5103_
	);
	LUT2 #(
		.INIT('h2)
	) name4572 (
		\sa02_reg[1]/P0001 ,
		_w5103_,
		_w5104_
	);
	LUT2 #(
		.INIT('h1)
	) name4573 (
		_w1039_,
		_w1130_,
		_w5105_
	);
	LUT2 #(
		.INIT('h4)
	) name4574 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		_w5106_
	);
	LUT2 #(
		.INIT('h4)
	) name4575 (
		_w5105_,
		_w5106_,
		_w5107_
	);
	LUT2 #(
		.INIT('h1)
	) name4576 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		_w5108_
	);
	LUT2 #(
		.INIT('h2)
	) name4577 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[5]/P0001 ,
		_w5109_
	);
	LUT2 #(
		.INIT('h4)
	) name4578 (
		_w1004_,
		_w5109_,
		_w5110_
	);
	LUT2 #(
		.INIT('h8)
	) name4579 (
		_w5108_,
		_w5110_,
		_w5111_
	);
	LUT2 #(
		.INIT('h1)
	) name4580 (
		_w5098_,
		_w5111_,
		_w5112_
	);
	LUT2 #(
		.INIT('h4)
	) name4581 (
		_w5101_,
		_w5112_,
		_w5113_
	);
	LUT2 #(
		.INIT('h4)
	) name4582 (
		_w5107_,
		_w5113_,
		_w5114_
	);
	LUT2 #(
		.INIT('h4)
	) name4583 (
		_w5104_,
		_w5114_,
		_w5115_
	);
	LUT2 #(
		.INIT('h4)
	) name4584 (
		_w5090_,
		_w5115_,
		_w5116_
	);
	LUT2 #(
		.INIT('h4)
	) name4585 (
		_w5096_,
		_w5116_,
		_w5117_
	);
	LUT2 #(
		.INIT('h2)
	) name4586 (
		\sa02_reg[0]/P0001 ,
		_w5117_,
		_w5118_
	);
	LUT2 #(
		.INIT('h4)
	) name4587 (
		\sa02_reg[2]/P0001 ,
		_w980_,
		_w5119_
	);
	LUT2 #(
		.INIT('h4)
	) name4588 (
		\sa02_reg[4]/P0001 ,
		_w5119_,
		_w5120_
	);
	LUT2 #(
		.INIT('h2)
	) name4589 (
		_w978_,
		_w997_,
		_w5121_
	);
	LUT2 #(
		.INIT('h8)
	) name4590 (
		\sa02_reg[6]/NET0131 ,
		_w1057_,
		_w5122_
	);
	LUT2 #(
		.INIT('h2)
	) name4591 (
		\sa02_reg[1]/P0001 ,
		_w5122_,
		_w5123_
	);
	LUT2 #(
		.INIT('h4)
	) name4592 (
		_w5120_,
		_w5123_,
		_w5124_
	);
	LUT2 #(
		.INIT('h4)
	) name4593 (
		_w5121_,
		_w5124_,
		_w5125_
	);
	LUT2 #(
		.INIT('h8)
	) name4594 (
		\sa02_reg[4]/P0001 ,
		_w1021_,
		_w5126_
	);
	LUT2 #(
		.INIT('h8)
	) name4595 (
		\sa02_reg[3]/P0001 ,
		_w1056_,
		_w5127_
	);
	LUT2 #(
		.INIT('h8)
	) name4596 (
		_w1016_,
		_w5127_,
		_w5128_
	);
	LUT2 #(
		.INIT('h8)
	) name4597 (
		_w974_,
		_w1023_,
		_w5129_
	);
	LUT2 #(
		.INIT('h4)
	) name4598 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w5130_
	);
	LUT2 #(
		.INIT('h8)
	) name4599 (
		_w1035_,
		_w5130_,
		_w5131_
	);
	LUT2 #(
		.INIT('h8)
	) name4600 (
		_w1000_,
		_w1095_,
		_w5132_
	);
	LUT2 #(
		.INIT('h1)
	) name4601 (
		\sa02_reg[1]/P0001 ,
		_w5099_,
		_w5133_
	);
	LUT2 #(
		.INIT('h1)
	) name4602 (
		_w5129_,
		_w5131_,
		_w5134_
	);
	LUT2 #(
		.INIT('h4)
	) name4603 (
		_w5132_,
		_w5134_,
		_w5135_
	);
	LUT2 #(
		.INIT('h4)
	) name4604 (
		_w5128_,
		_w5133_,
		_w5136_
	);
	LUT2 #(
		.INIT('h8)
	) name4605 (
		_w5135_,
		_w5136_,
		_w5137_
	);
	LUT2 #(
		.INIT('h4)
	) name4606 (
		_w5126_,
		_w5137_,
		_w5138_
	);
	LUT2 #(
		.INIT('h1)
	) name4607 (
		_w5125_,
		_w5138_,
		_w5139_
	);
	LUT2 #(
		.INIT('h8)
	) name4608 (
		_w975_,
		_w986_,
		_w5140_
	);
	LUT2 #(
		.INIT('h4)
	) name4609 (
		\sa02_reg[7]/NET0131 ,
		_w5140_,
		_w5141_
	);
	LUT2 #(
		.INIT('h4)
	) name4610 (
		_w979_,
		_w1035_,
		_w5142_
	);
	LUT2 #(
		.INIT('h2)
	) name4611 (
		\sa02_reg[4]/P0001 ,
		_w1019_,
		_w5143_
	);
	LUT2 #(
		.INIT('h2)
	) name4612 (
		_w5142_,
		_w5143_,
		_w5144_
	);
	LUT2 #(
		.INIT('h1)
	) name4613 (
		\sa02_reg[2]/P0001 ,
		_w987_,
		_w5145_
	);
	LUT2 #(
		.INIT('h4)
	) name4614 (
		_w5141_,
		_w5145_,
		_w5146_
	);
	LUT2 #(
		.INIT('h4)
	) name4615 (
		_w5144_,
		_w5146_,
		_w5147_
	);
	LUT2 #(
		.INIT('h8)
	) name4616 (
		_w974_,
		_w982_,
		_w5148_
	);
	LUT2 #(
		.INIT('h2)
	) name4617 (
		\sa02_reg[2]/P0001 ,
		_w5148_,
		_w5149_
	);
	LUT2 #(
		.INIT('h4)
	) name4618 (
		_w5126_,
		_w5149_,
		_w5150_
	);
	LUT2 #(
		.INIT('h1)
	) name4619 (
		_w5147_,
		_w5150_,
		_w5151_
	);
	LUT2 #(
		.INIT('h1)
	) name4620 (
		_w5139_,
		_w5151_,
		_w5152_
	);
	LUT2 #(
		.INIT('h1)
	) name4621 (
		\sa02_reg[0]/P0001 ,
		_w5152_,
		_w5153_
	);
	LUT2 #(
		.INIT('h8)
	) name4622 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		_w5154_
	);
	LUT2 #(
		.INIT('h4)
	) name4623 (
		\sa02_reg[3]/P0001 ,
		_w979_,
		_w5155_
	);
	LUT2 #(
		.INIT('h4)
	) name4624 (
		\sa02_reg[6]/NET0131 ,
		_w1030_,
		_w5156_
	);
	LUT2 #(
		.INIT('h1)
	) name4625 (
		_w5155_,
		_w5156_,
		_w5157_
	);
	LUT2 #(
		.INIT('h1)
	) name4626 (
		\sa02_reg[4]/P0001 ,
		_w5157_,
		_w5158_
	);
	LUT2 #(
		.INIT('h2)
	) name4627 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w5159_
	);
	LUT2 #(
		.INIT('h8)
	) name4628 (
		_w995_,
		_w5159_,
		_w5160_
	);
	LUT2 #(
		.INIT('h1)
	) name4629 (
		_w5158_,
		_w5160_,
		_w5161_
	);
	LUT2 #(
		.INIT('h2)
	) name4630 (
		_w5154_,
		_w5161_,
		_w5162_
	);
	LUT2 #(
		.INIT('h8)
	) name4631 (
		\sa02_reg[6]/NET0131 ,
		_w1007_,
		_w5163_
	);
	LUT2 #(
		.INIT('h1)
	) name4632 (
		_w1001_,
		_w5156_,
		_w5164_
	);
	LUT2 #(
		.INIT('h4)
	) name4633 (
		_w5163_,
		_w5164_,
		_w5165_
	);
	LUT2 #(
		.INIT('h1)
	) name4634 (
		\sa02_reg[2]/P0001 ,
		_w5165_,
		_w5166_
	);
	LUT2 #(
		.INIT('h8)
	) name4635 (
		_w1023_,
		_w1038_,
		_w5167_
	);
	LUT2 #(
		.INIT('h2)
	) name4636 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w5168_
	);
	LUT2 #(
		.INIT('h8)
	) name4637 (
		_w979_,
		_w5168_,
		_w5169_
	);
	LUT2 #(
		.INIT('h8)
	) name4638 (
		\sa02_reg[3]/P0001 ,
		_w5169_,
		_w5170_
	);
	LUT2 #(
		.INIT('h8)
	) name4639 (
		_w974_,
		_w975_,
		_w5171_
	);
	LUT2 #(
		.INIT('h8)
	) name4640 (
		_w993_,
		_w1004_,
		_w5172_
	);
	LUT2 #(
		.INIT('h8)
	) name4641 (
		\sa02_reg[2]/P0001 ,
		_w5172_,
		_w5173_
	);
	LUT2 #(
		.INIT('h1)
	) name4642 (
		_w5167_,
		_w5171_,
		_w5174_
	);
	LUT2 #(
		.INIT('h4)
	) name4643 (
		_w5170_,
		_w5174_,
		_w5175_
	);
	LUT2 #(
		.INIT('h4)
	) name4644 (
		_w5173_,
		_w5175_,
		_w5176_
	);
	LUT2 #(
		.INIT('h4)
	) name4645 (
		_w5166_,
		_w5176_,
		_w5177_
	);
	LUT2 #(
		.INIT('h1)
	) name4646 (
		\sa02_reg[1]/P0001 ,
		_w5177_,
		_w5178_
	);
	LUT2 #(
		.INIT('h2)
	) name4647 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		_w5179_
	);
	LUT2 #(
		.INIT('h8)
	) name4648 (
		_w1110_,
		_w5179_,
		_w5180_
	);
	LUT2 #(
		.INIT('h4)
	) name4649 (
		\sa02_reg[7]/NET0131 ,
		_w5148_,
		_w5181_
	);
	LUT2 #(
		.INIT('h8)
	) name4650 (
		_w1001_,
		_w1095_,
		_w5182_
	);
	LUT2 #(
		.INIT('h8)
	) name4651 (
		_w984_,
		_w5163_,
		_w5183_
	);
	LUT2 #(
		.INIT('h1)
	) name4652 (
		_w981_,
		_w5181_,
		_w5184_
	);
	LUT2 #(
		.INIT('h4)
	) name4653 (
		_w5182_,
		_w5184_,
		_w5185_
	);
	LUT2 #(
		.INIT('h1)
	) name4654 (
		_w5180_,
		_w5183_,
		_w5186_
	);
	LUT2 #(
		.INIT('h8)
	) name4655 (
		_w5185_,
		_w5186_,
		_w5187_
	);
	LUT2 #(
		.INIT('h4)
	) name4656 (
		_w5162_,
		_w5187_,
		_w5188_
	);
	LUT2 #(
		.INIT('h4)
	) name4657 (
		_w5178_,
		_w5188_,
		_w5189_
	);
	LUT2 #(
		.INIT('h4)
	) name4658 (
		_w5153_,
		_w5189_,
		_w5190_
	);
	LUT2 #(
		.INIT('h4)
	) name4659 (
		_w5118_,
		_w5190_,
		_w5191_
	);
	LUT2 #(
		.INIT('h2)
	) name4660 (
		_w689_,
		_w5191_,
		_w5192_
	);
	LUT2 #(
		.INIT('h4)
	) name4661 (
		_w689_,
		_w5191_,
		_w5193_
	);
	LUT2 #(
		.INIT('h1)
	) name4662 (
		_w5192_,
		_w5193_,
		_w5194_
	);
	LUT2 #(
		.INIT('h1)
	) name4663 (
		_w1142_,
		_w5194_,
		_w5195_
	);
	LUT2 #(
		.INIT('h8)
	) name4664 (
		_w1142_,
		_w5194_,
		_w5196_
	);
	LUT2 #(
		.INIT('h1)
	) name4665 (
		_w5195_,
		_w5196_,
		_w5197_
	);
	LUT2 #(
		.INIT('h8)
	) name4666 (
		\sa31_reg[4]/P0001 ,
		_w1178_,
		_w5198_
	);
	LUT2 #(
		.INIT('h4)
	) name4667 (
		\sa31_reg[4]/P0001 ,
		_w1149_,
		_w5199_
	);
	LUT2 #(
		.INIT('h1)
	) name4668 (
		_w5198_,
		_w5199_,
		_w5200_
	);
	LUT2 #(
		.INIT('h1)
	) name4669 (
		\sa31_reg[3]/P0001 ,
		_w5200_,
		_w5201_
	);
	LUT2 #(
		.INIT('h1)
	) name4670 (
		_w1206_,
		_w5201_,
		_w5202_
	);
	LUT2 #(
		.INIT('h1)
	) name4671 (
		\sa31_reg[2]/P0001 ,
		_w5202_,
		_w5203_
	);
	LUT2 #(
		.INIT('h8)
	) name4672 (
		_w1186_,
		_w1216_,
		_w5204_
	);
	LUT2 #(
		.INIT('h4)
	) name4673 (
		\sa31_reg[5]/P0001 ,
		_w1256_,
		_w5205_
	);
	LUT2 #(
		.INIT('h4)
	) name4674 (
		\sa31_reg[3]/P0001 ,
		_w5205_,
		_w5206_
	);
	LUT2 #(
		.INIT('h8)
	) name4675 (
		_w1152_,
		_w1194_,
		_w5207_
	);
	LUT2 #(
		.INIT('h8)
	) name4676 (
		\sa31_reg[4]/P0001 ,
		_w1167_,
		_w5208_
	);
	LUT2 #(
		.INIT('h8)
	) name4677 (
		\sa31_reg[4]/P0001 ,
		_w1194_,
		_w5209_
	);
	LUT2 #(
		.INIT('h1)
	) name4678 (
		_w1167_,
		_w5209_,
		_w5210_
	);
	LUT2 #(
		.INIT('h2)
	) name4679 (
		\sa31_reg[2]/P0001 ,
		_w5210_,
		_w5211_
	);
	LUT2 #(
		.INIT('h1)
	) name4680 (
		_w1148_,
		_w5204_,
		_w5212_
	);
	LUT2 #(
		.INIT('h1)
	) name4681 (
		_w5206_,
		_w5207_,
		_w5213_
	);
	LUT2 #(
		.INIT('h4)
	) name4682 (
		_w5208_,
		_w5213_,
		_w5214_
	);
	LUT2 #(
		.INIT('h8)
	) name4683 (
		_w5212_,
		_w5214_,
		_w5215_
	);
	LUT2 #(
		.INIT('h4)
	) name4684 (
		_w5211_,
		_w5215_,
		_w5216_
	);
	LUT2 #(
		.INIT('h4)
	) name4685 (
		_w5203_,
		_w5216_,
		_w5217_
	);
	LUT2 #(
		.INIT('h2)
	) name4686 (
		\sa31_reg[1]/P0001 ,
		_w5217_,
		_w5218_
	);
	LUT2 #(
		.INIT('h2)
	) name4687 (
		\sa31_reg[3]/P0001 ,
		_w1281_,
		_w5219_
	);
	LUT2 #(
		.INIT('h4)
	) name4688 (
		\sa31_reg[4]/P0001 ,
		_w1186_,
		_w5220_
	);
	LUT2 #(
		.INIT('h4)
	) name4689 (
		\sa31_reg[3]/P0001 ,
		_w1239_,
		_w5221_
	);
	LUT2 #(
		.INIT('h1)
	) name4690 (
		_w5219_,
		_w5220_,
		_w5222_
	);
	LUT2 #(
		.INIT('h4)
	) name4691 (
		_w5221_,
		_w5222_,
		_w5223_
	);
	LUT2 #(
		.INIT('h2)
	) name4692 (
		\sa31_reg[2]/P0001 ,
		_w5223_,
		_w5224_
	);
	LUT2 #(
		.INIT('h1)
	) name4693 (
		_w1247_,
		_w1255_,
		_w5225_
	);
	LUT2 #(
		.INIT('h2)
	) name4694 (
		\sa31_reg[7]/P0001 ,
		_w5225_,
		_w5226_
	);
	LUT2 #(
		.INIT('h8)
	) name4695 (
		_w1229_,
		_w1248_,
		_w5227_
	);
	LUT2 #(
		.INIT('h1)
	) name4696 (
		_w1221_,
		_w5227_,
		_w5228_
	);
	LUT2 #(
		.INIT('h4)
	) name4697 (
		_w5226_,
		_w5228_,
		_w5229_
	);
	LUT2 #(
		.INIT('h1)
	) name4698 (
		\sa31_reg[1]/P0001 ,
		_w5229_,
		_w5230_
	);
	LUT2 #(
		.INIT('h4)
	) name4699 (
		\sa31_reg[2]/P0001 ,
		_w1179_,
		_w5231_
	);
	LUT2 #(
		.INIT('h1)
	) name4700 (
		_w1205_,
		_w5231_,
		_w5232_
	);
	LUT2 #(
		.INIT('h4)
	) name4701 (
		_w1185_,
		_w5232_,
		_w5233_
	);
	LUT2 #(
		.INIT('h4)
	) name4702 (
		_w5224_,
		_w5233_,
		_w5234_
	);
	LUT2 #(
		.INIT('h4)
	) name4703 (
		_w5230_,
		_w5234_,
		_w5235_
	);
	LUT2 #(
		.INIT('h4)
	) name4704 (
		_w5218_,
		_w5235_,
		_w5236_
	);
	LUT2 #(
		.INIT('h1)
	) name4705 (
		\sa31_reg[0]/P0002 ,
		_w5236_,
		_w5237_
	);
	LUT2 #(
		.INIT('h4)
	) name4706 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		_w5238_
	);
	LUT2 #(
		.INIT('h4)
	) name4707 (
		\sa31_reg[5]/P0001 ,
		_w1146_,
		_w5239_
	);
	LUT2 #(
		.INIT('h8)
	) name4708 (
		_w5238_,
		_w5239_,
		_w5240_
	);
	LUT2 #(
		.INIT('h4)
	) name4709 (
		\sa31_reg[4]/P0001 ,
		_w1151_,
		_w5241_
	);
	LUT2 #(
		.INIT('h8)
	) name4710 (
		_w1159_,
		_w1186_,
		_w5242_
	);
	LUT2 #(
		.INIT('h1)
	) name4711 (
		_w5241_,
		_w5242_,
		_w5243_
	);
	LUT2 #(
		.INIT('h2)
	) name4712 (
		\sa31_reg[2]/P0001 ,
		_w5243_,
		_w5244_
	);
	LUT2 #(
		.INIT('h2)
	) name4713 (
		_w1194_,
		_w1279_,
		_w5245_
	);
	LUT2 #(
		.INIT('h1)
	) name4714 (
		_w1202_,
		_w5240_,
		_w5246_
	);
	LUT2 #(
		.INIT('h4)
	) name4715 (
		_w5245_,
		_w5246_,
		_w5247_
	);
	LUT2 #(
		.INIT('h4)
	) name4716 (
		_w5244_,
		_w5247_,
		_w5248_
	);
	LUT2 #(
		.INIT('h1)
	) name4717 (
		\sa31_reg[1]/P0001 ,
		_w5248_,
		_w5249_
	);
	LUT2 #(
		.INIT('h8)
	) name4718 (
		\sa31_reg[7]/P0001 ,
		_w1197_,
		_w5250_
	);
	LUT2 #(
		.INIT('h1)
	) name4719 (
		_w1161_,
		_w5250_,
		_w5251_
	);
	LUT2 #(
		.INIT('h4)
	) name4720 (
		\sa31_reg[7]/P0001 ,
		_w1196_,
		_w5252_
	);
	LUT2 #(
		.INIT('h8)
	) name4721 (
		_w1229_,
		_w5252_,
		_w5253_
	);
	LUT2 #(
		.INIT('h4)
	) name4722 (
		\sa31_reg[4]/P0001 ,
		_w1206_,
		_w5254_
	);
	LUT2 #(
		.INIT('h1)
	) name4723 (
		_w5253_,
		_w5254_,
		_w5255_
	);
	LUT2 #(
		.INIT('h8)
	) name4724 (
		_w5251_,
		_w5255_,
		_w5256_
	);
	LUT2 #(
		.INIT('h2)
	) name4725 (
		\sa31_reg[1]/P0001 ,
		_w5256_,
		_w5257_
	);
	LUT2 #(
		.INIT('h8)
	) name4726 (
		_w1151_,
		_w1230_,
		_w5258_
	);
	LUT2 #(
		.INIT('h1)
	) name4727 (
		_w1202_,
		_w5258_,
		_w5259_
	);
	LUT2 #(
		.INIT('h2)
	) name4728 (
		\sa31_reg[2]/P0001 ,
		_w5259_,
		_w5260_
	);
	LUT2 #(
		.INIT('h8)
	) name4729 (
		_w1151_,
		_w1174_,
		_w5261_
	);
	LUT2 #(
		.INIT('h4)
	) name4730 (
		\sa31_reg[2]/P0001 ,
		_w5261_,
		_w5262_
	);
	LUT2 #(
		.INIT('h8)
	) name4731 (
		\sa31_reg[5]/P0001 ,
		_w1225_,
		_w5263_
	);
	LUT2 #(
		.INIT('h8)
	) name4732 (
		_w1149_,
		_w5263_,
		_w5264_
	);
	LUT2 #(
		.INIT('h2)
	) name4733 (
		_w1164_,
		_w1174_,
		_w5265_
	);
	LUT2 #(
		.INIT('h1)
	) name4734 (
		_w5263_,
		_w5265_,
		_w5266_
	);
	LUT2 #(
		.INIT('h2)
	) name4735 (
		\sa31_reg[1]/P0001 ,
		_w5266_,
		_w5267_
	);
	LUT2 #(
		.INIT('h4)
	) name4736 (
		\sa31_reg[4]/P0001 ,
		_w1158_,
		_w5268_
	);
	LUT2 #(
		.INIT('h8)
	) name4737 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w5269_
	);
	LUT2 #(
		.INIT('h8)
	) name4738 (
		_w1158_,
		_w5269_,
		_w5270_
	);
	LUT2 #(
		.INIT('h8)
	) name4739 (
		_w1149_,
		_w1225_,
		_w5271_
	);
	LUT2 #(
		.INIT('h1)
	) name4740 (
		_w5270_,
		_w5271_,
		_w5272_
	);
	LUT2 #(
		.INIT('h4)
	) name4741 (
		_w5268_,
		_w5272_,
		_w5273_
	);
	LUT2 #(
		.INIT('h4)
	) name4742 (
		_w5267_,
		_w5273_,
		_w5274_
	);
	LUT2 #(
		.INIT('h1)
	) name4743 (
		\sa31_reg[2]/P0001 ,
		_w5274_,
		_w5275_
	);
	LUT2 #(
		.INIT('h1)
	) name4744 (
		_w5262_,
		_w5264_,
		_w5276_
	);
	LUT2 #(
		.INIT('h4)
	) name4745 (
		_w5260_,
		_w5276_,
		_w5277_
	);
	LUT2 #(
		.INIT('h4)
	) name4746 (
		_w5257_,
		_w5277_,
		_w5278_
	);
	LUT2 #(
		.INIT('h4)
	) name4747 (
		_w5249_,
		_w5278_,
		_w5279_
	);
	LUT2 #(
		.INIT('h4)
	) name4748 (
		_w5275_,
		_w5279_,
		_w5280_
	);
	LUT2 #(
		.INIT('h2)
	) name4749 (
		\sa31_reg[0]/P0002 ,
		_w5280_,
		_w5281_
	);
	LUT2 #(
		.INIT('h1)
	) name4750 (
		_w1153_,
		_w1200_,
		_w5282_
	);
	LUT2 #(
		.INIT('h2)
	) name4751 (
		\sa31_reg[5]/P0001 ,
		_w5282_,
		_w5283_
	);
	LUT2 #(
		.INIT('h1)
	) name4752 (
		_w5261_,
		_w5283_,
		_w5284_
	);
	LUT2 #(
		.INIT('h1)
	) name4753 (
		\sa31_reg[2]/P0001 ,
		_w5284_,
		_w5285_
	);
	LUT2 #(
		.INIT('h2)
	) name4754 (
		\sa31_reg[3]/P0001 ,
		_w1178_,
		_w5286_
	);
	LUT2 #(
		.INIT('h1)
	) name4755 (
		_w1173_,
		_w5239_,
		_w5287_
	);
	LUT2 #(
		.INIT('h1)
	) name4756 (
		\sa31_reg[3]/P0001 ,
		_w1201_,
		_w5288_
	);
	LUT2 #(
		.INIT('h8)
	) name4757 (
		_w5287_,
		_w5288_,
		_w5289_
	);
	LUT2 #(
		.INIT('h2)
	) name4758 (
		_w1215_,
		_w5286_,
		_w5290_
	);
	LUT2 #(
		.INIT('h4)
	) name4759 (
		_w5289_,
		_w5290_,
		_w5291_
	);
	LUT2 #(
		.INIT('h1)
	) name4760 (
		_w1234_,
		_w5291_,
		_w5292_
	);
	LUT2 #(
		.INIT('h4)
	) name4761 (
		_w5285_,
		_w5292_,
		_w5293_
	);
	LUT2 #(
		.INIT('h1)
	) name4762 (
		\sa31_reg[1]/P0001 ,
		_w5293_,
		_w5294_
	);
	LUT2 #(
		.INIT('h8)
	) name4763 (
		\sa31_reg[4]/P0001 ,
		_w1266_,
		_w5295_
	);
	LUT2 #(
		.INIT('h1)
	) name4764 (
		_w1227_,
		_w5206_,
		_w5296_
	);
	LUT2 #(
		.INIT('h1)
	) name4765 (
		\sa31_reg[2]/P0001 ,
		_w5296_,
		_w5297_
	);
	LUT2 #(
		.INIT('h8)
	) name4766 (
		\sa31_reg[2]/P0001 ,
		_w1261_,
		_w5298_
	);
	LUT2 #(
		.INIT('h4)
	) name4767 (
		\sa31_reg[4]/P0001 ,
		_w5204_,
		_w5299_
	);
	LUT2 #(
		.INIT('h1)
	) name4768 (
		_w5231_,
		_w5299_,
		_w5300_
	);
	LUT2 #(
		.INIT('h4)
	) name4769 (
		_w5298_,
		_w5300_,
		_w5301_
	);
	LUT2 #(
		.INIT('h2)
	) name4770 (
		\sa31_reg[1]/P0001 ,
		_w5301_,
		_w5302_
	);
	LUT2 #(
		.INIT('h1)
	) name4771 (
		_w5295_,
		_w5297_,
		_w5303_
	);
	LUT2 #(
		.INIT('h4)
	) name4772 (
		_w5302_,
		_w5303_,
		_w5304_
	);
	LUT2 #(
		.INIT('h4)
	) name4773 (
		_w5294_,
		_w5304_,
		_w5305_
	);
	LUT2 #(
		.INIT('h4)
	) name4774 (
		_w5281_,
		_w5305_,
		_w5306_
	);
	LUT2 #(
		.INIT('h4)
	) name4775 (
		_w5237_,
		_w5306_,
		_w5307_
	);
	LUT2 #(
		.INIT('h2)
	) name4776 (
		\u0_w_reg[2][6]/P0001 ,
		_w5307_,
		_w5308_
	);
	LUT2 #(
		.INIT('h4)
	) name4777 (
		\u0_w_reg[2][6]/P0001 ,
		_w5307_,
		_w5309_
	);
	LUT2 #(
		.INIT('h1)
	) name4778 (
		_w5308_,
		_w5309_,
		_w5310_
	);
	LUT2 #(
		.INIT('h8)
	) name4779 (
		_w850_,
		_w5310_,
		_w5311_
	);
	LUT2 #(
		.INIT('h1)
	) name4780 (
		_w850_,
		_w5310_,
		_w5312_
	);
	LUT2 #(
		.INIT('h1)
	) name4781 (
		_w5311_,
		_w5312_,
		_w5313_
	);
	LUT2 #(
		.INIT('h4)
	) name4782 (
		_w5197_,
		_w5313_,
		_w5314_
	);
	LUT2 #(
		.INIT('h2)
	) name4783 (
		_w5197_,
		_w5313_,
		_w5315_
	);
	LUT2 #(
		.INIT('h1)
	) name4784 (
		\ld_r_reg/P0001 ,
		_w5314_,
		_w5316_
	);
	LUT2 #(
		.INIT('h4)
	) name4785 (
		_w5315_,
		_w5316_,
		_w5317_
	);
	LUT2 #(
		.INIT('h1)
	) name4786 (
		\text_in_r_reg[38]/P0001 ,
		\u0_w_reg[2][6]/P0001 ,
		_w5318_
	);
	LUT2 #(
		.INIT('h8)
	) name4787 (
		\text_in_r_reg[38]/P0001 ,
		\u0_w_reg[2][6]/P0001 ,
		_w5319_
	);
	LUT2 #(
		.INIT('h2)
	) name4788 (
		\ld_r_reg/P0001 ,
		_w5318_,
		_w5320_
	);
	LUT2 #(
		.INIT('h4)
	) name4789 (
		_w5319_,
		_w5320_,
		_w5321_
	);
	LUT2 #(
		.INIT('h1)
	) name4790 (
		_w5317_,
		_w5321_,
		_w5322_
	);
	LUT2 #(
		.INIT('h8)
	) name4791 (
		\sa02_reg[4]/P0001 ,
		_w982_,
		_w5323_
	);
	LUT2 #(
		.INIT('h1)
	) name4792 (
		_w1004_,
		_w5323_,
		_w5324_
	);
	LUT2 #(
		.INIT('h8)
	) name4793 (
		\sa02_reg[3]/P0001 ,
		_w1025_,
		_w5325_
	);
	LUT2 #(
		.INIT('h1)
	) name4794 (
		_w5155_,
		_w5325_,
		_w5326_
	);
	LUT2 #(
		.INIT('h8)
	) name4795 (
		_w5324_,
		_w5326_,
		_w5327_
	);
	LUT2 #(
		.INIT('h2)
	) name4796 (
		\sa02_reg[1]/P0001 ,
		_w5327_,
		_w5328_
	);
	LUT2 #(
		.INIT('h8)
	) name4797 (
		_w974_,
		_w1019_,
		_w5329_
	);
	LUT2 #(
		.INIT('h1)
	) name4798 (
		_w1022_,
		_w1031_,
		_w5330_
	);
	LUT2 #(
		.INIT('h4)
	) name4799 (
		_w5329_,
		_w5330_,
		_w5331_
	);
	LUT2 #(
		.INIT('h4)
	) name4800 (
		_w5328_,
		_w5331_,
		_w5332_
	);
	LUT2 #(
		.INIT('h2)
	) name4801 (
		\sa02_reg[2]/P0001 ,
		_w5332_,
		_w5333_
	);
	LUT2 #(
		.INIT('h8)
	) name4802 (
		_w984_,
		_w1090_,
		_w5334_
	);
	LUT2 #(
		.INIT('h4)
	) name4803 (
		\sa02_reg[2]/P0001 ,
		_w1025_,
		_w5335_
	);
	LUT2 #(
		.INIT('h1)
	) name4804 (
		_w1056_,
		_w5335_,
		_w5336_
	);
	LUT2 #(
		.INIT('h2)
	) name4805 (
		_w986_,
		_w5336_,
		_w5337_
	);
	LUT2 #(
		.INIT('h8)
	) name4806 (
		_w1011_,
		_w1039_,
		_w5338_
	);
	LUT2 #(
		.INIT('h8)
	) name4807 (
		_w1094_,
		_w5108_,
		_w5339_
	);
	LUT2 #(
		.INIT('h1)
	) name4808 (
		_w5338_,
		_w5339_,
		_w5340_
	);
	LUT2 #(
		.INIT('h2)
	) name4809 (
		\sa02_reg[1]/P0001 ,
		_w5340_,
		_w5341_
	);
	LUT2 #(
		.INIT('h8)
	) name4810 (
		\sa02_reg[2]/P0001 ,
		_w974_,
		_w5342_
	);
	LUT2 #(
		.INIT('h8)
	) name4811 (
		_w1003_,
		_w5342_,
		_w5343_
	);
	LUT2 #(
		.INIT('h2)
	) name4812 (
		\sa02_reg[2]/P0001 ,
		_w986_,
		_w5344_
	);
	LUT2 #(
		.INIT('h2)
	) name4813 (
		_w1025_,
		_w1035_,
		_w5345_
	);
	LUT2 #(
		.INIT('h4)
	) name4814 (
		_w5344_,
		_w5345_,
		_w5346_
	);
	LUT2 #(
		.INIT('h8)
	) name4815 (
		_w999_,
		_w1059_,
		_w5347_
	);
	LUT2 #(
		.INIT('h2)
	) name4816 (
		\sa02_reg[4]/P0001 ,
		_w999_,
		_w5348_
	);
	LUT2 #(
		.INIT('h1)
	) name4817 (
		\sa02_reg[2]/P0001 ,
		_w1020_,
		_w5349_
	);
	LUT2 #(
		.INIT('h8)
	) name4818 (
		_w5348_,
		_w5349_,
		_w5350_
	);
	LUT2 #(
		.INIT('h1)
	) name4819 (
		_w5343_,
		_w5347_,
		_w5351_
	);
	LUT2 #(
		.INIT('h4)
	) name4820 (
		_w5346_,
		_w5351_,
		_w5352_
	);
	LUT2 #(
		.INIT('h4)
	) name4821 (
		_w5350_,
		_w5352_,
		_w5353_
	);
	LUT2 #(
		.INIT('h1)
	) name4822 (
		\sa02_reg[1]/P0001 ,
		_w5353_,
		_w5354_
	);
	LUT2 #(
		.INIT('h2)
	) name4823 (
		\sa02_reg[0]/P0001 ,
		_w5334_,
		_w5355_
	);
	LUT2 #(
		.INIT('h4)
	) name4824 (
		_w5337_,
		_w5355_,
		_w5356_
	);
	LUT2 #(
		.INIT('h4)
	) name4825 (
		_w5341_,
		_w5356_,
		_w5357_
	);
	LUT2 #(
		.INIT('h4)
	) name4826 (
		_w5333_,
		_w5357_,
		_w5358_
	);
	LUT2 #(
		.INIT('h4)
	) name4827 (
		_w5354_,
		_w5358_,
		_w5359_
	);
	LUT2 #(
		.INIT('h1)
	) name4828 (
		_w5122_,
		_w5160_,
		_w5360_
	);
	LUT2 #(
		.INIT('h1)
	) name4829 (
		\sa02_reg[2]/P0001 ,
		_w5360_,
		_w5361_
	);
	LUT2 #(
		.INIT('h8)
	) name4830 (
		_w1037_,
		_w5168_,
		_w5362_
	);
	LUT2 #(
		.INIT('h8)
	) name4831 (
		_w1056_,
		_w5159_,
		_w5363_
	);
	LUT2 #(
		.INIT('h8)
	) name4832 (
		_w975_,
		_w1000_,
		_w5364_
	);
	LUT2 #(
		.INIT('h1)
	) name4833 (
		_w5363_,
		_w5364_,
		_w5365_
	);
	LUT2 #(
		.INIT('h2)
	) name4834 (
		_w984_,
		_w5365_,
		_w5366_
	);
	LUT2 #(
		.INIT('h2)
	) name4835 (
		\sa02_reg[5]/P0001 ,
		_w1023_,
		_w5367_
	);
	LUT2 #(
		.INIT('h4)
	) name4836 (
		_w1006_,
		_w5108_,
		_w5368_
	);
	LUT2 #(
		.INIT('h8)
	) name4837 (
		_w5367_,
		_w5368_,
		_w5369_
	);
	LUT2 #(
		.INIT('h1)
	) name4838 (
		_w979_,
		_w1039_,
		_w5370_
	);
	LUT2 #(
		.INIT('h2)
	) name4839 (
		_w5097_,
		_w5370_,
		_w5371_
	);
	LUT2 #(
		.INIT('h4)
	) name4840 (
		\sa02_reg[2]/P0001 ,
		_w5130_,
		_w5372_
	);
	LUT2 #(
		.INIT('h1)
	) name4841 (
		\sa02_reg[1]/P0001 ,
		_w5102_,
		_w5373_
	);
	LUT2 #(
		.INIT('h4)
	) name4842 (
		_w5372_,
		_w5373_,
		_w5374_
	);
	LUT2 #(
		.INIT('h4)
	) name4843 (
		_w5371_,
		_w5374_,
		_w5375_
	);
	LUT2 #(
		.INIT('h1)
	) name4844 (
		_w1130_,
		_w5159_,
		_w5376_
	);
	LUT2 #(
		.INIT('h2)
	) name4845 (
		_w1095_,
		_w5376_,
		_w5377_
	);
	LUT2 #(
		.INIT('h2)
	) name4846 (
		\sa02_reg[1]/P0001 ,
		_w1013_,
		_w5378_
	);
	LUT2 #(
		.INIT('h4)
	) name4847 (
		_w5156_,
		_w5378_,
		_w5379_
	);
	LUT2 #(
		.INIT('h1)
	) name4848 (
		_w5126_,
		_w5377_,
		_w5380_
	);
	LUT2 #(
		.INIT('h8)
	) name4849 (
		_w5379_,
		_w5380_,
		_w5381_
	);
	LUT2 #(
		.INIT('h1)
	) name4850 (
		_w5375_,
		_w5381_,
		_w5382_
	);
	LUT2 #(
		.INIT('h1)
	) name4851 (
		\sa02_reg[0]/P0001 ,
		_w5369_,
		_w5383_
	);
	LUT2 #(
		.INIT('h4)
	) name4852 (
		_w5362_,
		_w5383_,
		_w5384_
	);
	LUT2 #(
		.INIT('h4)
	) name4853 (
		_w5366_,
		_w5384_,
		_w5385_
	);
	LUT2 #(
		.INIT('h4)
	) name4854 (
		_w5361_,
		_w5385_,
		_w5386_
	);
	LUT2 #(
		.INIT('h4)
	) name4855 (
		_w5382_,
		_w5386_,
		_w5387_
	);
	LUT2 #(
		.INIT('h1)
	) name4856 (
		_w5359_,
		_w5387_,
		_w5388_
	);
	LUT2 #(
		.INIT('h1)
	) name4857 (
		_w1072_,
		_w5172_,
		_w5389_
	);
	LUT2 #(
		.INIT('h2)
	) name4858 (
		_w999_,
		_w5130_,
		_w5390_
	);
	LUT2 #(
		.INIT('h2)
	) name4859 (
		_w5389_,
		_w5390_,
		_w5391_
	);
	LUT2 #(
		.INIT('h2)
	) name4860 (
		_w1095_,
		_w5391_,
		_w5392_
	);
	LUT2 #(
		.INIT('h2)
	) name4861 (
		\sa02_reg[7]/NET0131 ,
		_w5324_,
		_w5393_
	);
	LUT2 #(
		.INIT('h4)
	) name4862 (
		\sa02_reg[6]/NET0131 ,
		_w1084_,
		_w5394_
	);
	LUT2 #(
		.INIT('h1)
	) name4863 (
		_w5393_,
		_w5394_,
		_w5395_
	);
	LUT2 #(
		.INIT('h1)
	) name4864 (
		\sa02_reg[3]/P0001 ,
		_w5395_,
		_w5396_
	);
	LUT2 #(
		.INIT('h1)
	) name4865 (
		_w1005_,
		_w1082_,
		_w5397_
	);
	LUT2 #(
		.INIT('h4)
	) name4866 (
		_w5396_,
		_w5397_,
		_w5398_
	);
	LUT2 #(
		.INIT('h2)
	) name4867 (
		\sa02_reg[2]/P0001 ,
		_w5398_,
		_w5399_
	);
	LUT2 #(
		.INIT('h1)
	) name4868 (
		_w5392_,
		_w5399_,
		_w5400_
	);
	LUT2 #(
		.INIT('h2)
	) name4869 (
		\sa02_reg[1]/P0001 ,
		_w5400_,
		_w5401_
	);
	LUT2 #(
		.INIT('h4)
	) name4870 (
		\sa02_reg[7]/NET0131 ,
		_w5171_,
		_w5402_
	);
	LUT2 #(
		.INIT('h4)
	) name4871 (
		\sa02_reg[5]/P0001 ,
		_w1091_,
		_w5403_
	);
	LUT2 #(
		.INIT('h1)
	) name4872 (
		_w5402_,
		_w5403_,
		_w5404_
	);
	LUT2 #(
		.INIT('h1)
	) name4873 (
		\sa02_reg[2]/P0001 ,
		_w5404_,
		_w5405_
	);
	LUT2 #(
		.INIT('h1)
	) name4874 (
		_w1037_,
		_w5140_,
		_w5406_
	);
	LUT2 #(
		.INIT('h4)
	) name4875 (
		_w5338_,
		_w5406_,
		_w5407_
	);
	LUT2 #(
		.INIT('h2)
	) name4876 (
		\sa02_reg[2]/P0001 ,
		_w5407_,
		_w5408_
	);
	LUT2 #(
		.INIT('h8)
	) name4877 (
		_w986_,
		_w993_,
		_w5409_
	);
	LUT2 #(
		.INIT('h8)
	) name4878 (
		_w1035_,
		_w5372_,
		_w5410_
	);
	LUT2 #(
		.INIT('h1)
	) name4879 (
		_w5369_,
		_w5409_,
		_w5411_
	);
	LUT2 #(
		.INIT('h4)
	) name4880 (
		_w5410_,
		_w5411_,
		_w5412_
	);
	LUT2 #(
		.INIT('h4)
	) name4881 (
		_w5408_,
		_w5412_,
		_w5413_
	);
	LUT2 #(
		.INIT('h1)
	) name4882 (
		\sa02_reg[1]/P0001 ,
		_w5413_,
		_w5414_
	);
	LUT2 #(
		.INIT('h1)
	) name4883 (
		_w5405_,
		_w5414_,
		_w5415_
	);
	LUT2 #(
		.INIT('h4)
	) name4884 (
		_w5388_,
		_w5415_,
		_w5416_
	);
	LUT2 #(
		.INIT('h4)
	) name4885 (
		_w5401_,
		_w5416_,
		_w5417_
	);
	LUT2 #(
		.INIT('h2)
	) name4886 (
		\sa13_reg[4]/P0001 ,
		_w532_,
		_w5418_
	);
	LUT2 #(
		.INIT('h4)
	) name4887 (
		_w855_,
		_w5418_,
		_w5419_
	);
	LUT2 #(
		.INIT('h1)
	) name4888 (
		_w861_,
		_w5419_,
		_w5420_
	);
	LUT2 #(
		.INIT('h1)
	) name4889 (
		\sa13_reg[2]/P0001 ,
		_w5420_,
		_w5421_
	);
	LUT2 #(
		.INIT('h4)
	) name4890 (
		\sa13_reg[7]/NET0131 ,
		_w620_,
		_w5422_
	);
	LUT2 #(
		.INIT('h8)
	) name4891 (
		_w532_,
		_w655_,
		_w5423_
	);
	LUT2 #(
		.INIT('h1)
	) name4892 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w5424_
	);
	LUT2 #(
		.INIT('h8)
	) name4893 (
		_w543_,
		_w5424_,
		_w5425_
	);
	LUT2 #(
		.INIT('h8)
	) name4894 (
		_w570_,
		_w653_,
		_w5426_
	);
	LUT2 #(
		.INIT('h8)
	) name4895 (
		\sa13_reg[2]/P0001 ,
		_w5426_,
		_w5427_
	);
	LUT2 #(
		.INIT('h1)
	) name4896 (
		_w5423_,
		_w5425_,
		_w5428_
	);
	LUT2 #(
		.INIT('h4)
	) name4897 (
		_w5422_,
		_w5428_,
		_w5429_
	);
	LUT2 #(
		.INIT('h4)
	) name4898 (
		_w5427_,
		_w5429_,
		_w5430_
	);
	LUT2 #(
		.INIT('h4)
	) name4899 (
		_w5421_,
		_w5430_,
		_w5431_
	);
	LUT2 #(
		.INIT('h1)
	) name4900 (
		\sa13_reg[1]/P0001 ,
		_w5431_,
		_w5432_
	);
	LUT2 #(
		.INIT('h4)
	) name4901 (
		\sa13_reg[2]/P0001 ,
		_w5422_,
		_w5433_
	);
	LUT2 #(
		.INIT('h4)
	) name4902 (
		\sa13_reg[3]/P0001 ,
		_w584_,
		_w5434_
	);
	LUT2 #(
		.INIT('h1)
	) name4903 (
		_w534_,
		_w858_,
		_w5435_
	);
	LUT2 #(
		.INIT('h4)
	) name4904 (
		_w5434_,
		_w5435_,
		_w5436_
	);
	LUT2 #(
		.INIT('h2)
	) name4905 (
		\sa13_reg[2]/P0001 ,
		_w5436_,
		_w5437_
	);
	LUT2 #(
		.INIT('h8)
	) name4906 (
		_w533_,
		_w900_,
		_w5438_
	);
	LUT2 #(
		.INIT('h8)
	) name4907 (
		_w623_,
		_w928_,
		_w5439_
	);
	LUT2 #(
		.INIT('h8)
	) name4908 (
		\sa13_reg[3]/P0001 ,
		_w913_,
		_w5440_
	);
	LUT2 #(
		.INIT('h1)
	) name4909 (
		_w563_,
		_w632_,
		_w5441_
	);
	LUT2 #(
		.INIT('h4)
	) name4910 (
		\sa13_reg[3]/P0001 ,
		_w556_,
		_w5442_
	);
	LUT2 #(
		.INIT('h1)
	) name4911 (
		_w544_,
		_w5442_,
		_w5443_
	);
	LUT2 #(
		.INIT('h8)
	) name4912 (
		_w5441_,
		_w5443_,
		_w5444_
	);
	LUT2 #(
		.INIT('h2)
	) name4913 (
		\sa13_reg[2]/P0001 ,
		_w5444_,
		_w5445_
	);
	LUT2 #(
		.INIT('h8)
	) name4914 (
		_w549_,
		_w565_,
		_w5446_
	);
	LUT2 #(
		.INIT('h1)
	) name4915 (
		_w5440_,
		_w5446_,
		_w5447_
	);
	LUT2 #(
		.INIT('h4)
	) name4916 (
		_w5445_,
		_w5447_,
		_w5448_
	);
	LUT2 #(
		.INIT('h2)
	) name4917 (
		\sa13_reg[1]/P0001 ,
		_w5448_,
		_w5449_
	);
	LUT2 #(
		.INIT('h2)
	) name4918 (
		\sa13_reg[0]/P0001 ,
		_w5438_,
		_w5450_
	);
	LUT2 #(
		.INIT('h4)
	) name4919 (
		_w5439_,
		_w5450_,
		_w5451_
	);
	LUT2 #(
		.INIT('h4)
	) name4920 (
		_w5433_,
		_w5451_,
		_w5452_
	);
	LUT2 #(
		.INIT('h4)
	) name4921 (
		_w5437_,
		_w5452_,
		_w5453_
	);
	LUT2 #(
		.INIT('h4)
	) name4922 (
		_w5432_,
		_w5453_,
		_w5454_
	);
	LUT2 #(
		.INIT('h4)
	) name4923 (
		_w5449_,
		_w5454_,
		_w5455_
	);
	LUT2 #(
		.INIT('h8)
	) name4924 (
		\sa13_reg[4]/P0001 ,
		_w570_,
		_w5456_
	);
	LUT2 #(
		.INIT('h8)
	) name4925 (
		_w623_,
		_w5456_,
		_w5457_
	);
	LUT2 #(
		.INIT('h4)
	) name4926 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w5458_
	);
	LUT2 #(
		.INIT('h4)
	) name4927 (
		\sa13_reg[2]/P0001 ,
		_w5458_,
		_w5459_
	);
	LUT2 #(
		.INIT('h1)
	) name4928 (
		_w561_,
		_w5459_,
		_w5460_
	);
	LUT2 #(
		.INIT('h1)
	) name4929 (
		_w887_,
		_w5457_,
		_w5461_
	);
	LUT2 #(
		.INIT('h8)
	) name4930 (
		_w5460_,
		_w5461_,
		_w5462_
	);
	LUT2 #(
		.INIT('h1)
	) name4931 (
		\sa13_reg[1]/P0001 ,
		_w5462_,
		_w5463_
	);
	LUT2 #(
		.INIT('h8)
	) name4932 (
		_w604_,
		_w623_,
		_w5464_
	);
	LUT2 #(
		.INIT('h4)
	) name4933 (
		\sa13_reg[6]/NET0131 ,
		_w5464_,
		_w5465_
	);
	LUT2 #(
		.INIT('h8)
	) name4934 (
		\sa13_reg[4]/P0001 ,
		_w557_,
		_w5466_
	);
	LUT2 #(
		.INIT('h1)
	) name4935 (
		_w907_,
		_w5466_,
		_w5467_
	);
	LUT2 #(
		.INIT('h2)
	) name4936 (
		_w623_,
		_w5467_,
		_w5468_
	);
	LUT2 #(
		.INIT('h1)
	) name4937 (
		_w540_,
		_w901_,
		_w5469_
	);
	LUT2 #(
		.INIT('h2)
	) name4938 (
		_w5424_,
		_w5469_,
		_w5470_
	);
	LUT2 #(
		.INIT('h1)
	) name4939 (
		_w609_,
		_w652_,
		_w5471_
	);
	LUT2 #(
		.INIT('h1)
	) name4940 (
		\sa13_reg[2]/P0001 ,
		_w5471_,
		_w5472_
	);
	LUT2 #(
		.INIT('h4)
	) name4941 (
		_w611_,
		_w621_,
		_w5473_
	);
	LUT2 #(
		.INIT('h1)
	) name4942 (
		_w648_,
		_w946_,
		_w5474_
	);
	LUT2 #(
		.INIT('h1)
	) name4943 (
		\sa13_reg[2]/P0001 ,
		_w5474_,
		_w5475_
	);
	LUT2 #(
		.INIT('h8)
	) name4944 (
		\sa13_reg[5]/P0001 ,
		_w864_,
		_w5476_
	);
	LUT2 #(
		.INIT('h1)
	) name4945 (
		_w5473_,
		_w5476_,
		_w5477_
	);
	LUT2 #(
		.INIT('h4)
	) name4946 (
		_w5475_,
		_w5477_,
		_w5478_
	);
	LUT2 #(
		.INIT('h2)
	) name4947 (
		\sa13_reg[1]/P0001 ,
		_w5478_,
		_w5479_
	);
	LUT2 #(
		.INIT('h1)
	) name4948 (
		\sa13_reg[0]/P0001 ,
		_w5465_,
		_w5480_
	);
	LUT2 #(
		.INIT('h4)
	) name4949 (
		_w5470_,
		_w5480_,
		_w5481_
	);
	LUT2 #(
		.INIT('h1)
	) name4950 (
		_w5468_,
		_w5472_,
		_w5482_
	);
	LUT2 #(
		.INIT('h8)
	) name4951 (
		_w5481_,
		_w5482_,
		_w5483_
	);
	LUT2 #(
		.INIT('h4)
	) name4952 (
		_w5463_,
		_w5483_,
		_w5484_
	);
	LUT2 #(
		.INIT('h4)
	) name4953 (
		_w5479_,
		_w5484_,
		_w5485_
	);
	LUT2 #(
		.INIT('h1)
	) name4954 (
		_w5455_,
		_w5485_,
		_w5486_
	);
	LUT2 #(
		.INIT('h1)
	) name4955 (
		_w888_,
		_w908_,
		_w5487_
	);
	LUT2 #(
		.INIT('h2)
	) name4956 (
		_w532_,
		_w5458_,
		_w5488_
	);
	LUT2 #(
		.INIT('h2)
	) name4957 (
		_w5487_,
		_w5488_,
		_w5489_
	);
	LUT2 #(
		.INIT('h2)
	) name4958 (
		_w581_,
		_w5489_,
		_w5490_
	);
	LUT2 #(
		.INIT('h2)
	) name4959 (
		\sa13_reg[7]/NET0131 ,
		_w5441_,
		_w5491_
	);
	LUT2 #(
		.INIT('h4)
	) name4960 (
		\sa13_reg[6]/NET0131 ,
		_w901_,
		_w5492_
	);
	LUT2 #(
		.INIT('h1)
	) name4961 (
		_w5491_,
		_w5492_,
		_w5493_
	);
	LUT2 #(
		.INIT('h1)
	) name4962 (
		\sa13_reg[3]/P0001 ,
		_w5493_,
		_w5494_
	);
	LUT2 #(
		.INIT('h1)
	) name4963 (
		_w571_,
		_w902_,
		_w5495_
	);
	LUT2 #(
		.INIT('h4)
	) name4964 (
		_w5494_,
		_w5495_,
		_w5496_
	);
	LUT2 #(
		.INIT('h2)
	) name4965 (
		\sa13_reg[2]/P0001 ,
		_w5496_,
		_w5497_
	);
	LUT2 #(
		.INIT('h1)
	) name4966 (
		_w5490_,
		_w5497_,
		_w5498_
	);
	LUT2 #(
		.INIT('h2)
	) name4967 (
		\sa13_reg[1]/P0001 ,
		_w5498_,
		_w5499_
	);
	LUT2 #(
		.INIT('h8)
	) name4968 (
		_w579_,
		_w946_,
		_w5500_
	);
	LUT2 #(
		.INIT('h1)
	) name4969 (
		_w863_,
		_w5500_,
		_w5501_
	);
	LUT2 #(
		.INIT('h1)
	) name4970 (
		\sa13_reg[2]/P0001 ,
		_w5501_,
		_w5502_
	);
	LUT2 #(
		.INIT('h8)
	) name4971 (
		_w550_,
		_w5459_,
		_w5503_
	);
	LUT2 #(
		.INIT('h8)
	) name4972 (
		_w533_,
		_w559_,
		_w5504_
	);
	LUT2 #(
		.INIT('h8)
	) name4973 (
		\sa13_reg[4]/P0001 ,
		_w535_,
		_w5505_
	);
	LUT2 #(
		.INIT('h4)
	) name4974 (
		\sa13_reg[3]/P0001 ,
		_w5505_,
		_w5506_
	);
	LUT2 #(
		.INIT('h1)
	) name4975 (
		_w854_,
		_w5440_,
		_w5507_
	);
	LUT2 #(
		.INIT('h4)
	) name4976 (
		_w5506_,
		_w5507_,
		_w5508_
	);
	LUT2 #(
		.INIT('h2)
	) name4977 (
		\sa13_reg[2]/P0001 ,
		_w5508_,
		_w5509_
	);
	LUT2 #(
		.INIT('h1)
	) name4978 (
		_w5503_,
		_w5504_,
		_w5510_
	);
	LUT2 #(
		.INIT('h4)
	) name4979 (
		_w5470_,
		_w5510_,
		_w5511_
	);
	LUT2 #(
		.INIT('h4)
	) name4980 (
		_w5509_,
		_w5511_,
		_w5512_
	);
	LUT2 #(
		.INIT('h1)
	) name4981 (
		\sa13_reg[1]/P0001 ,
		_w5512_,
		_w5513_
	);
	LUT2 #(
		.INIT('h1)
	) name4982 (
		_w5502_,
		_w5513_,
		_w5514_
	);
	LUT2 #(
		.INIT('h4)
	) name4983 (
		_w5486_,
		_w5514_,
		_w5515_
	);
	LUT2 #(
		.INIT('h4)
	) name4984 (
		_w5499_,
		_w5515_,
		_w5516_
	);
	LUT2 #(
		.INIT('h2)
	) name4985 (
		_w5417_,
		_w5516_,
		_w5517_
	);
	LUT2 #(
		.INIT('h4)
	) name4986 (
		_w5417_,
		_w5516_,
		_w5518_
	);
	LUT2 #(
		.INIT('h1)
	) name4987 (
		_w5517_,
		_w5518_,
		_w5519_
	);
	LUT2 #(
		.INIT('h1)
	) name4988 (
		_w5191_,
		_w5519_,
		_w5520_
	);
	LUT2 #(
		.INIT('h8)
	) name4989 (
		_w5191_,
		_w5519_,
		_w5521_
	);
	LUT2 #(
		.INIT('h1)
	) name4990 (
		_w5520_,
		_w5521_,
		_w5522_
	);
	LUT2 #(
		.INIT('h4)
	) name4991 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w5523_
	);
	LUT2 #(
		.INIT('h8)
	) name4992 (
		_w777_,
		_w5523_,
		_w5524_
	);
	LUT2 #(
		.INIT('h8)
	) name4993 (
		_w690_,
		_w745_,
		_w5525_
	);
	LUT2 #(
		.INIT('h2)
	) name4994 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w5526_
	);
	LUT2 #(
		.INIT('h4)
	) name4995 (
		\sa20_reg[3]/P0001 ,
		_w693_,
		_w5527_
	);
	LUT2 #(
		.INIT('h4)
	) name4996 (
		_w5526_,
		_w5527_,
		_w5528_
	);
	LUT2 #(
		.INIT('h4)
	) name4997 (
		\sa20_reg[4]/P0001 ,
		_w720_,
		_w5529_
	);
	LUT2 #(
		.INIT('h4)
	) name4998 (
		\sa20_reg[3]/P0001 ,
		_w5529_,
		_w5530_
	);
	LUT2 #(
		.INIT('h2)
	) name4999 (
		\sa20_reg[2]/P0001 ,
		_w5530_,
		_w5531_
	);
	LUT2 #(
		.INIT('h8)
	) name5000 (
		\sa20_reg[4]/P0001 ,
		_w701_,
		_w5532_
	);
	LUT2 #(
		.INIT('h1)
	) name5001 (
		\sa20_reg[2]/P0001 ,
		_w739_,
		_w5533_
	);
	LUT2 #(
		.INIT('h1)
	) name5002 (
		_w791_,
		_w5532_,
		_w5534_
	);
	LUT2 #(
		.INIT('h8)
	) name5003 (
		_w5533_,
		_w5534_,
		_w5535_
	);
	LUT2 #(
		.INIT('h1)
	) name5004 (
		_w5531_,
		_w5535_,
		_w5536_
	);
	LUT2 #(
		.INIT('h1)
	) name5005 (
		_w5524_,
		_w5525_,
		_w5537_
	);
	LUT2 #(
		.INIT('h4)
	) name5006 (
		_w5528_,
		_w5537_,
		_w5538_
	);
	LUT2 #(
		.INIT('h4)
	) name5007 (
		_w5536_,
		_w5538_,
		_w5539_
	);
	LUT2 #(
		.INIT('h1)
	) name5008 (
		\sa20_reg[1]/P0001 ,
		_w5539_,
		_w5540_
	);
	LUT2 #(
		.INIT('h8)
	) name5009 (
		_w735_,
		_w5526_,
		_w5541_
	);
	LUT2 #(
		.INIT('h8)
	) name5010 (
		\sa20_reg[3]/P0001 ,
		_w5541_,
		_w5542_
	);
	LUT2 #(
		.INIT('h8)
	) name5011 (
		\sa20_reg[4]/P0001 ,
		_w795_,
		_w5543_
	);
	LUT2 #(
		.INIT('h4)
	) name5012 (
		\sa20_reg[5]/P0001 ,
		_w705_,
		_w5544_
	);
	LUT2 #(
		.INIT('h8)
	) name5013 (
		_w747_,
		_w5544_,
		_w5545_
	);
	LUT2 #(
		.INIT('h1)
	) name5014 (
		_w5543_,
		_w5545_,
		_w5546_
	);
	LUT2 #(
		.INIT('h2)
	) name5015 (
		\sa20_reg[1]/P0001 ,
		_w5546_,
		_w5547_
	);
	LUT2 #(
		.INIT('h8)
	) name5016 (
		_w739_,
		_w747_,
		_w5548_
	);
	LUT2 #(
		.INIT('h8)
	) name5017 (
		_w691_,
		_w777_,
		_w5549_
	);
	LUT2 #(
		.INIT('h8)
	) name5018 (
		_w719_,
		_w736_,
		_w5550_
	);
	LUT2 #(
		.INIT('h1)
	) name5019 (
		_w719_,
		_w791_,
		_w5551_
	);
	LUT2 #(
		.INIT('h4)
	) name5020 (
		\sa20_reg[3]/P0001 ,
		_w723_,
		_w5552_
	);
	LUT2 #(
		.INIT('h1)
	) name5021 (
		_w699_,
		_w5552_,
		_w5553_
	);
	LUT2 #(
		.INIT('h8)
	) name5022 (
		_w5551_,
		_w5553_,
		_w5554_
	);
	LUT2 #(
		.INIT('h2)
	) name5023 (
		\sa20_reg[1]/P0001 ,
		_w5554_,
		_w5555_
	);
	LUT2 #(
		.INIT('h8)
	) name5024 (
		\sa20_reg[5]/P0001 ,
		_w739_,
		_w5556_
	);
	LUT2 #(
		.INIT('h1)
	) name5025 (
		_w692_,
		_w5550_,
		_w5557_
	);
	LUT2 #(
		.INIT('h4)
	) name5026 (
		_w5556_,
		_w5557_,
		_w5558_
	);
	LUT2 #(
		.INIT('h4)
	) name5027 (
		_w5555_,
		_w5558_,
		_w5559_
	);
	LUT2 #(
		.INIT('h2)
	) name5028 (
		\sa20_reg[2]/P0001 ,
		_w5559_,
		_w5560_
	);
	LUT2 #(
		.INIT('h1)
	) name5029 (
		_w5542_,
		_w5549_,
		_w5561_
	);
	LUT2 #(
		.INIT('h4)
	) name5030 (
		_w5548_,
		_w5561_,
		_w5562_
	);
	LUT2 #(
		.INIT('h4)
	) name5031 (
		_w5547_,
		_w5562_,
		_w5563_
	);
	LUT2 #(
		.INIT('h4)
	) name5032 (
		_w5540_,
		_w5563_,
		_w5564_
	);
	LUT2 #(
		.INIT('h4)
	) name5033 (
		_w5560_,
		_w5564_,
		_w5565_
	);
	LUT2 #(
		.INIT('h2)
	) name5034 (
		\sa20_reg[0]/P0001 ,
		_w5565_,
		_w5566_
	);
	LUT2 #(
		.INIT('h8)
	) name5035 (
		_w717_,
		_w719_,
		_w5567_
	);
	LUT2 #(
		.INIT('h1)
	) name5036 (
		_w827_,
		_w5567_,
		_w5568_
	);
	LUT2 #(
		.INIT('h2)
	) name5037 (
		_w690_,
		_w765_,
		_w5569_
	);
	LUT2 #(
		.INIT('h2)
	) name5038 (
		_w5568_,
		_w5569_,
		_w5570_
	);
	LUT2 #(
		.INIT('h2)
	) name5039 (
		_w763_,
		_w5570_,
		_w5571_
	);
	LUT2 #(
		.INIT('h2)
	) name5040 (
		\sa20_reg[7]/NET0131 ,
		_w5551_,
		_w5572_
	);
	LUT2 #(
		.INIT('h8)
	) name5041 (
		_w694_,
		_w723_,
		_w5573_
	);
	LUT2 #(
		.INIT('h1)
	) name5042 (
		_w5572_,
		_w5573_,
		_w5574_
	);
	LUT2 #(
		.INIT('h1)
	) name5043 (
		\sa20_reg[3]/P0001 ,
		_w5574_,
		_w5575_
	);
	LUT2 #(
		.INIT('h1)
	) name5044 (
		_w721_,
		_w778_,
		_w5576_
	);
	LUT2 #(
		.INIT('h4)
	) name5045 (
		_w5575_,
		_w5576_,
		_w5577_
	);
	LUT2 #(
		.INIT('h2)
	) name5046 (
		\sa20_reg[2]/P0001 ,
		_w5577_,
		_w5578_
	);
	LUT2 #(
		.INIT('h1)
	) name5047 (
		_w5571_,
		_w5578_,
		_w5579_
	);
	LUT2 #(
		.INIT('h2)
	) name5048 (
		\sa20_reg[1]/P0001 ,
		_w5579_,
		_w5580_
	);
	LUT2 #(
		.INIT('h8)
	) name5049 (
		\sa20_reg[2]/P0001 ,
		_w820_,
		_w5581_
	);
	LUT2 #(
		.INIT('h1)
	) name5050 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w5582_
	);
	LUT2 #(
		.INIT('h1)
	) name5051 (
		_w810_,
		_w5582_,
		_w5583_
	);
	LUT2 #(
		.INIT('h2)
	) name5052 (
		\sa20_reg[7]/NET0131 ,
		_w5583_,
		_w5584_
	);
	LUT2 #(
		.INIT('h8)
	) name5053 (
		\sa20_reg[4]/P0001 ,
		_w720_,
		_w5585_
	);
	LUT2 #(
		.INIT('h8)
	) name5054 (
		_w761_,
		_w5585_,
		_w5586_
	);
	LUT2 #(
		.INIT('h1)
	) name5055 (
		\sa20_reg[1]/P0001 ,
		_w5581_,
		_w5587_
	);
	LUT2 #(
		.INIT('h4)
	) name5056 (
		_w5586_,
		_w5587_,
		_w5588_
	);
	LUT2 #(
		.INIT('h4)
	) name5057 (
		_w5584_,
		_w5588_,
		_w5589_
	);
	LUT2 #(
		.INIT('h2)
	) name5058 (
		\sa20_reg[1]/P0001 ,
		_w834_,
		_w5590_
	);
	LUT2 #(
		.INIT('h8)
	) name5059 (
		_w693_,
		_w706_,
		_w5591_
	);
	LUT2 #(
		.INIT('h1)
	) name5060 (
		_w750_,
		_w5591_,
		_w5592_
	);
	LUT2 #(
		.INIT('h1)
	) name5061 (
		\sa20_reg[2]/P0001 ,
		_w5592_,
		_w5593_
	);
	LUT2 #(
		.INIT('h1)
	) name5062 (
		_w736_,
		_w819_,
		_w5594_
	);
	LUT2 #(
		.INIT('h2)
	) name5063 (
		_w767_,
		_w5594_,
		_w5595_
	);
	LUT2 #(
		.INIT('h2)
	) name5064 (
		_w5590_,
		_w5595_,
		_w5596_
	);
	LUT2 #(
		.INIT('h4)
	) name5065 (
		_w5593_,
		_w5596_,
		_w5597_
	);
	LUT2 #(
		.INIT('h1)
	) name5066 (
		_w5589_,
		_w5597_,
		_w5598_
	);
	LUT2 #(
		.INIT('h8)
	) name5067 (
		_w701_,
		_w736_,
		_w5599_
	);
	LUT2 #(
		.INIT('h8)
	) name5068 (
		_w777_,
		_w799_,
		_w5600_
	);
	LUT2 #(
		.INIT('h1)
	) name5069 (
		_w5599_,
		_w5600_,
		_w5601_
	);
	LUT2 #(
		.INIT('h1)
	) name5070 (
		_w779_,
		_w808_,
		_w5602_
	);
	LUT2 #(
		.INIT('h8)
	) name5071 (
		_w5601_,
		_w5602_,
		_w5603_
	);
	LUT2 #(
		.INIT('h1)
	) name5072 (
		\sa20_reg[2]/P0001 ,
		_w5603_,
		_w5604_
	);
	LUT2 #(
		.INIT('h8)
	) name5073 (
		_w701_,
		_w714_,
		_w5605_
	);
	LUT2 #(
		.INIT('h8)
	) name5074 (
		\sa20_reg[4]/P0001 ,
		_w724_,
		_w5606_
	);
	LUT2 #(
		.INIT('h1)
	) name5075 (
		_w710_,
		_w5605_,
		_w5607_
	);
	LUT2 #(
		.INIT('h4)
	) name5076 (
		_w5606_,
		_w5607_,
		_w5608_
	);
	LUT2 #(
		.INIT('h2)
	) name5077 (
		_w761_,
		_w5608_,
		_w5609_
	);
	LUT2 #(
		.INIT('h1)
	) name5078 (
		_w5604_,
		_w5609_,
		_w5610_
	);
	LUT2 #(
		.INIT('h4)
	) name5079 (
		_w5598_,
		_w5610_,
		_w5611_
	);
	LUT2 #(
		.INIT('h1)
	) name5080 (
		\sa20_reg[0]/P0001 ,
		_w5611_,
		_w5612_
	);
	LUT2 #(
		.INIT('h8)
	) name5081 (
		_w694_,
		_w5527_,
		_w5613_
	);
	LUT2 #(
		.INIT('h4)
	) name5082 (
		\sa20_reg[6]/NET0131 ,
		_w718_,
		_w5614_
	);
	LUT2 #(
		.INIT('h1)
	) name5083 (
		_w5613_,
		_w5614_,
		_w5615_
	);
	LUT2 #(
		.INIT('h1)
	) name5084 (
		\sa20_reg[2]/P0001 ,
		_w5615_,
		_w5616_
	);
	LUT2 #(
		.INIT('h8)
	) name5085 (
		_w691_,
		_w744_,
		_w5617_
	);
	LUT2 #(
		.INIT('h2)
	) name5086 (
		\sa20_reg[2]/P0001 ,
		_w5543_,
		_w5618_
	);
	LUT2 #(
		.INIT('h8)
	) name5087 (
		\sa20_reg[3]/P0001 ,
		_w708_,
		_w5619_
	);
	LUT2 #(
		.INIT('h4)
	) name5088 (
		\sa20_reg[7]/NET0131 ,
		_w5619_,
		_w5620_
	);
	LUT2 #(
		.INIT('h1)
	) name5089 (
		_w702_,
		_w5620_,
		_w5621_
	);
	LUT2 #(
		.INIT('h8)
	) name5090 (
		_w5618_,
		_w5621_,
		_w5622_
	);
	LUT2 #(
		.INIT('h1)
	) name5091 (
		\sa20_reg[2]/P0001 ,
		_w766_,
		_w5623_
	);
	LUT2 #(
		.INIT('h8)
	) name5092 (
		_w5601_,
		_w5623_,
		_w5624_
	);
	LUT2 #(
		.INIT('h1)
	) name5093 (
		_w5622_,
		_w5624_,
		_w5625_
	);
	LUT2 #(
		.INIT('h1)
	) name5094 (
		_w5617_,
		_w5625_,
		_w5626_
	);
	LUT2 #(
		.INIT('h1)
	) name5095 (
		\sa20_reg[1]/P0001 ,
		_w5626_,
		_w5627_
	);
	LUT2 #(
		.INIT('h1)
	) name5096 (
		_w5616_,
		_w5627_,
		_w5628_
	);
	LUT2 #(
		.INIT('h4)
	) name5097 (
		_w5612_,
		_w5628_,
		_w5629_
	);
	LUT2 #(
		.INIT('h4)
	) name5098 (
		_w5566_,
		_w5629_,
		_w5630_
	);
	LUT2 #(
		.INIT('h4)
	) name5099 (
		_w5580_,
		_w5630_,
		_w5631_
	);
	LUT2 #(
		.INIT('h2)
	) name5100 (
		\u0_w_reg[2][7]/P0001 ,
		_w5631_,
		_w5632_
	);
	LUT2 #(
		.INIT('h4)
	) name5101 (
		\u0_w_reg[2][7]/P0001 ,
		_w5631_,
		_w5633_
	);
	LUT2 #(
		.INIT('h1)
	) name5102 (
		_w5632_,
		_w5633_,
		_w5634_
	);
	LUT2 #(
		.INIT('h8)
	) name5103 (
		_w1300_,
		_w5634_,
		_w5635_
	);
	LUT2 #(
		.INIT('h1)
	) name5104 (
		_w1300_,
		_w5634_,
		_w5636_
	);
	LUT2 #(
		.INIT('h1)
	) name5105 (
		_w5635_,
		_w5636_,
		_w5637_
	);
	LUT2 #(
		.INIT('h1)
	) name5106 (
		_w5522_,
		_w5637_,
		_w5638_
	);
	LUT2 #(
		.INIT('h8)
	) name5107 (
		_w5522_,
		_w5637_,
		_w5639_
	);
	LUT2 #(
		.INIT('h1)
	) name5108 (
		\ld_r_reg/P0001 ,
		_w5638_,
		_w5640_
	);
	LUT2 #(
		.INIT('h4)
	) name5109 (
		_w5639_,
		_w5640_,
		_w5641_
	);
	LUT2 #(
		.INIT('h2)
	) name5110 (
		\text_in_r_reg[39]/P0001 ,
		\u0_w_reg[2][7]/P0001 ,
		_w5642_
	);
	LUT2 #(
		.INIT('h4)
	) name5111 (
		\text_in_r_reg[39]/P0001 ,
		\u0_w_reg[2][7]/P0001 ,
		_w5643_
	);
	LUT2 #(
		.INIT('h2)
	) name5112 (
		\ld_r_reg/P0001 ,
		_w5642_,
		_w5644_
	);
	LUT2 #(
		.INIT('h4)
	) name5113 (
		_w5643_,
		_w5644_,
		_w5645_
	);
	LUT2 #(
		.INIT('h1)
	) name5114 (
		_w5641_,
		_w5645_,
		_w5646_
	);
	LUT2 #(
		.INIT('h8)
	) name5115 (
		\sa13_reg[2]/P0001 ,
		_w588_,
		_w5647_
	);
	LUT2 #(
		.INIT('h8)
	) name5116 (
		\sa13_reg[5]/P0001 ,
		_w5459_,
		_w5648_
	);
	LUT2 #(
		.INIT('h8)
	) name5117 (
		_w611_,
		_w946_,
		_w5649_
	);
	LUT2 #(
		.INIT('h8)
	) name5118 (
		\sa13_reg[3]/P0001 ,
		_w583_,
		_w5650_
	);
	LUT2 #(
		.INIT('h4)
	) name5119 (
		\sa13_reg[4]/P0001 ,
		_w5650_,
		_w5651_
	);
	LUT2 #(
		.INIT('h1)
	) name5120 (
		\sa13_reg[1]/P0001 ,
		_w560_,
		_w5652_
	);
	LUT2 #(
		.INIT('h4)
	) name5121 (
		_w5647_,
		_w5652_,
		_w5653_
	);
	LUT2 #(
		.INIT('h1)
	) name5122 (
		_w5648_,
		_w5649_,
		_w5654_
	);
	LUT2 #(
		.INIT('h4)
	) name5123 (
		_w5651_,
		_w5654_,
		_w5655_
	);
	LUT2 #(
		.INIT('h8)
	) name5124 (
		_w5653_,
		_w5655_,
		_w5656_
	);
	LUT2 #(
		.INIT('h2)
	) name5125 (
		\sa13_reg[1]/P0001 ,
		_w681_,
		_w5657_
	);
	LUT2 #(
		.INIT('h8)
	) name5126 (
		\sa13_reg[7]/NET0131 ,
		_w632_,
		_w5658_
	);
	LUT2 #(
		.INIT('h1)
	) name5127 (
		_w865_,
		_w5658_,
		_w5659_
	);
	LUT2 #(
		.INIT('h1)
	) name5128 (
		\sa13_reg[2]/P0001 ,
		_w5659_,
		_w5660_
	);
	LUT2 #(
		.INIT('h8)
	) name5129 (
		_w549_,
		_w670_,
		_w5661_
	);
	LUT2 #(
		.INIT('h1)
	) name5130 (
		_w918_,
		_w5661_,
		_w5662_
	);
	LUT2 #(
		.INIT('h8)
	) name5131 (
		_w5657_,
		_w5662_,
		_w5663_
	);
	LUT2 #(
		.INIT('h4)
	) name5132 (
		_w5660_,
		_w5663_,
		_w5664_
	);
	LUT2 #(
		.INIT('h1)
	) name5133 (
		_w5656_,
		_w5664_,
		_w5665_
	);
	LUT2 #(
		.INIT('h1)
	) name5134 (
		_w616_,
		_w655_,
		_w5666_
	);
	LUT2 #(
		.INIT('h1)
	) name5135 (
		\sa13_reg[6]/NET0131 ,
		_w5666_,
		_w5667_
	);
	LUT2 #(
		.INIT('h2)
	) name5136 (
		\sa13_reg[2]/P0001 ,
		_w637_,
		_w5668_
	);
	LUT2 #(
		.INIT('h4)
	) name5137 (
		_w888_,
		_w5668_,
		_w5669_
	);
	LUT2 #(
		.INIT('h4)
	) name5138 (
		_w5667_,
		_w5669_,
		_w5670_
	);
	LUT2 #(
		.INIT('h8)
	) name5139 (
		_w550_,
		_w583_,
		_w5671_
	);
	LUT2 #(
		.INIT('h1)
	) name5140 (
		\sa13_reg[2]/P0001 ,
		_w5671_,
		_w5672_
	);
	LUT2 #(
		.INIT('h4)
	) name5141 (
		_w683_,
		_w5672_,
		_w5673_
	);
	LUT2 #(
		.INIT('h4)
	) name5142 (
		_w903_,
		_w5673_,
		_w5674_
	);
	LUT2 #(
		.INIT('h1)
	) name5143 (
		_w5670_,
		_w5674_,
		_w5675_
	);
	LUT2 #(
		.INIT('h1)
	) name5144 (
		_w5665_,
		_w5675_,
		_w5676_
	);
	LUT2 #(
		.INIT('h2)
	) name5145 (
		\sa13_reg[0]/P0001 ,
		_w5676_,
		_w5677_
	);
	LUT2 #(
		.INIT('h8)
	) name5146 (
		_w557_,
		_w653_,
		_w5678_
	);
	LUT2 #(
		.INIT('h8)
	) name5147 (
		_w547_,
		_w5458_,
		_w5679_
	);
	LUT2 #(
		.INIT('h4)
	) name5148 (
		\sa13_reg[3]/P0001 ,
		_w5679_,
		_w5680_
	);
	LUT2 #(
		.INIT('h2)
	) name5149 (
		\sa13_reg[5]/P0001 ,
		_w5443_,
		_w5681_
	);
	LUT2 #(
		.INIT('h8)
	) name5150 (
		_w547_,
		_w592_,
		_w5682_
	);
	LUT2 #(
		.INIT('h2)
	) name5151 (
		\sa13_reg[2]/P0001 ,
		_w5423_,
		_w5683_
	);
	LUT2 #(
		.INIT('h4)
	) name5152 (
		_w5680_,
		_w5683_,
		_w5684_
	);
	LUT2 #(
		.INIT('h4)
	) name5153 (
		_w5682_,
		_w5684_,
		_w5685_
	);
	LUT2 #(
		.INIT('h4)
	) name5154 (
		_w5681_,
		_w5685_,
		_w5686_
	);
	LUT2 #(
		.INIT('h8)
	) name5155 (
		\sa13_reg[5]/P0001 ,
		_w5651_,
		_w5687_
	);
	LUT2 #(
		.INIT('h1)
	) name5156 (
		\sa13_reg[2]/P0001 ,
		_w621_,
		_w5688_
	);
	LUT2 #(
		.INIT('h4)
	) name5157 (
		_w856_,
		_w5688_,
		_w5689_
	);
	LUT2 #(
		.INIT('h4)
	) name5158 (
		_w5687_,
		_w5689_,
		_w5690_
	);
	LUT2 #(
		.INIT('h1)
	) name5159 (
		_w5686_,
		_w5690_,
		_w5691_
	);
	LUT2 #(
		.INIT('h1)
	) name5160 (
		_w609_,
		_w5678_,
		_w5692_
	);
	LUT2 #(
		.INIT('h4)
	) name5161 (
		_w5691_,
		_w5692_,
		_w5693_
	);
	LUT2 #(
		.INIT('h1)
	) name5162 (
		\sa13_reg[1]/P0001 ,
		_w5693_,
		_w5694_
	);
	LUT2 #(
		.INIT('h4)
	) name5163 (
		\sa13_reg[2]/P0001 ,
		_w908_,
		_w5695_
	);
	LUT2 #(
		.INIT('h8)
	) name5164 (
		\sa13_reg[2]/P0001 ,
		_w5505_,
		_w5696_
	);
	LUT2 #(
		.INIT('h1)
	) name5165 (
		_w5695_,
		_w5696_,
		_w5697_
	);
	LUT2 #(
		.INIT('h2)
	) name5166 (
		\sa13_reg[3]/P0001 ,
		_w5697_,
		_w5698_
	);
	LUT2 #(
		.INIT('h8)
	) name5167 (
		\sa13_reg[7]/NET0131 ,
		_w668_,
		_w5699_
	);
	LUT2 #(
		.INIT('h1)
	) name5168 (
		_w634_,
		_w683_,
		_w5700_
	);
	LUT2 #(
		.INIT('h4)
	) name5169 (
		_w5699_,
		_w5700_,
		_w5701_
	);
	LUT2 #(
		.INIT('h1)
	) name5170 (
		\sa13_reg[2]/P0001 ,
		_w5701_,
		_w5702_
	);
	LUT2 #(
		.INIT('h8)
	) name5171 (
		_w567_,
		_w603_,
		_w5703_
	);
	LUT2 #(
		.INIT('h8)
	) name5172 (
		_w955_,
		_w5458_,
		_w5704_
	);
	LUT2 #(
		.INIT('h1)
	) name5173 (
		_w624_,
		_w5440_,
		_w5705_
	);
	LUT2 #(
		.INIT('h1)
	) name5174 (
		_w5703_,
		_w5704_,
		_w5706_
	);
	LUT2 #(
		.INIT('h8)
	) name5175 (
		_w5705_,
		_w5706_,
		_w5707_
	);
	LUT2 #(
		.INIT('h4)
	) name5176 (
		_w5702_,
		_w5707_,
		_w5708_
	);
	LUT2 #(
		.INIT('h2)
	) name5177 (
		\sa13_reg[1]/P0001 ,
		_w5708_,
		_w5709_
	);
	LUT2 #(
		.INIT('h1)
	) name5178 (
		_w914_,
		_w5492_,
		_w5710_
	);
	LUT2 #(
		.INIT('h1)
	) name5179 (
		\sa13_reg[3]/P0001 ,
		_w5710_,
		_w5711_
	);
	LUT2 #(
		.INIT('h8)
	) name5180 (
		_w653_,
		_w912_,
		_w5712_
	);
	LUT2 #(
		.INIT('h1)
	) name5181 (
		_w5500_,
		_w5712_,
		_w5713_
	);
	LUT2 #(
		.INIT('h2)
	) name5182 (
		\sa13_reg[2]/P0001 ,
		_w5713_,
		_w5714_
	);
	LUT2 #(
		.INIT('h8)
	) name5183 (
		\sa13_reg[3]/P0001 ,
		_w672_,
		_w5715_
	);
	LUT2 #(
		.INIT('h8)
	) name5184 (
		_w861_,
		_w5424_,
		_w5716_
	);
	LUT2 #(
		.INIT('h1)
	) name5185 (
		_w887_,
		_w5696_,
		_w5717_
	);
	LUT2 #(
		.INIT('h1)
	) name5186 (
		_w5715_,
		_w5716_,
		_w5718_
	);
	LUT2 #(
		.INIT('h8)
	) name5187 (
		_w5717_,
		_w5718_,
		_w5719_
	);
	LUT2 #(
		.INIT('h1)
	) name5188 (
		\sa13_reg[1]/P0001 ,
		_w5719_,
		_w5720_
	);
	LUT2 #(
		.INIT('h2)
	) name5189 (
		_w568_,
		_w655_,
		_w5721_
	);
	LUT2 #(
		.INIT('h1)
	) name5190 (
		_w5679_,
		_w5721_,
		_w5722_
	);
	LUT2 #(
		.INIT('h1)
	) name5191 (
		\sa13_reg[2]/P0001 ,
		_w5722_,
		_w5723_
	);
	LUT2 #(
		.INIT('h8)
	) name5192 (
		_w603_,
		_w5456_,
		_w5724_
	);
	LUT2 #(
		.INIT('h8)
	) name5193 (
		\sa13_reg[2]/P0001 ,
		_w861_,
		_w5725_
	);
	LUT2 #(
		.INIT('h1)
	) name5194 (
		_w545_,
		_w5724_,
		_w5726_
	);
	LUT2 #(
		.INIT('h4)
	) name5195 (
		_w5725_,
		_w5726_,
		_w5727_
	);
	LUT2 #(
		.INIT('h4)
	) name5196 (
		_w5723_,
		_w5727_,
		_w5728_
	);
	LUT2 #(
		.INIT('h2)
	) name5197 (
		\sa13_reg[1]/P0001 ,
		_w5728_,
		_w5729_
	);
	LUT2 #(
		.INIT('h1)
	) name5198 (
		_w5711_,
		_w5714_,
		_w5730_
	);
	LUT2 #(
		.INIT('h4)
	) name5199 (
		_w5720_,
		_w5730_,
		_w5731_
	);
	LUT2 #(
		.INIT('h4)
	) name5200 (
		_w5729_,
		_w5731_,
		_w5732_
	);
	LUT2 #(
		.INIT('h1)
	) name5201 (
		\sa13_reg[0]/P0001 ,
		_w5732_,
		_w5733_
	);
	LUT2 #(
		.INIT('h1)
	) name5202 (
		_w5698_,
		_w5709_,
		_w5734_
	);
	LUT2 #(
		.INIT('h4)
	) name5203 (
		_w5694_,
		_w5734_,
		_w5735_
	);
	LUT2 #(
		.INIT('h4)
	) name5204 (
		_w5733_,
		_w5735_,
		_w5736_
	);
	LUT2 #(
		.INIT('h4)
	) name5205 (
		_w5677_,
		_w5736_,
		_w5737_
	);
	LUT2 #(
		.INIT('h4)
	) name5206 (
		\sa02_reg[3]/P0001 ,
		_w1088_,
		_w5738_
	);
	LUT2 #(
		.INIT('h4)
	) name5207 (
		\sa02_reg[2]/P0001 ,
		_w5738_,
		_w5739_
	);
	LUT2 #(
		.INIT('h1)
	) name5208 (
		_w1116_,
		_w5739_,
		_w5740_
	);
	LUT2 #(
		.INIT('h1)
	) name5209 (
		\sa02_reg[1]/P0001 ,
		_w5740_,
		_w5741_
	);
	LUT2 #(
		.INIT('h1)
	) name5210 (
		_w5083_,
		_w5403_,
		_w5742_
	);
	LUT2 #(
		.INIT('h2)
	) name5211 (
		\sa02_reg[2]/P0001 ,
		_w5742_,
		_w5743_
	);
	LUT2 #(
		.INIT('h8)
	) name5212 (
		\sa02_reg[4]/P0001 ,
		_w975_,
		_w5744_
	);
	LUT2 #(
		.INIT('h1)
	) name5213 (
		_w980_,
		_w5744_,
		_w5745_
	);
	LUT2 #(
		.INIT('h2)
	) name5214 (
		_w5106_,
		_w5745_,
		_w5746_
	);
	LUT2 #(
		.INIT('h1)
	) name5215 (
		_w1077_,
		_w5394_,
		_w5747_
	);
	LUT2 #(
		.INIT('h1)
	) name5216 (
		\sa02_reg[3]/P0001 ,
		_w5747_,
		_w5748_
	);
	LUT2 #(
		.INIT('h2)
	) name5217 (
		_w1042_,
		_w1059_,
		_w5749_
	);
	LUT2 #(
		.INIT('h8)
	) name5218 (
		_w982_,
		_w5130_,
		_w5750_
	);
	LUT2 #(
		.INIT('h1)
	) name5219 (
		_w5749_,
		_w5750_,
		_w5751_
	);
	LUT2 #(
		.INIT('h1)
	) name5220 (
		\sa02_reg[2]/P0001 ,
		_w5751_,
		_w5752_
	);
	LUT2 #(
		.INIT('h8)
	) name5221 (
		\sa02_reg[2]/P0001 ,
		_w1056_,
		_w5753_
	);
	LUT2 #(
		.INIT('h8)
	) name5222 (
		\sa02_reg[6]/NET0131 ,
		_w5753_,
		_w5754_
	);
	LUT2 #(
		.INIT('h8)
	) name5223 (
		\sa02_reg[4]/P0001 ,
		_w1003_,
		_w5755_
	);
	LUT2 #(
		.INIT('h8)
	) name5224 (
		_w978_,
		_w5755_,
		_w5756_
	);
	LUT2 #(
		.INIT('h1)
	) name5225 (
		_w1123_,
		_w5754_,
		_w5757_
	);
	LUT2 #(
		.INIT('h4)
	) name5226 (
		_w5756_,
		_w5757_,
		_w5758_
	);
	LUT2 #(
		.INIT('h4)
	) name5227 (
		_w5752_,
		_w5758_,
		_w5759_
	);
	LUT2 #(
		.INIT('h2)
	) name5228 (
		\sa02_reg[1]/P0001 ,
		_w5759_,
		_w5760_
	);
	LUT2 #(
		.INIT('h1)
	) name5229 (
		_w5743_,
		_w5746_,
		_w5761_
	);
	LUT2 #(
		.INIT('h4)
	) name5230 (
		_w5748_,
		_w5761_,
		_w5762_
	);
	LUT2 #(
		.INIT('h4)
	) name5231 (
		_w5741_,
		_w5762_,
		_w5763_
	);
	LUT2 #(
		.INIT('h4)
	) name5232 (
		_w5760_,
		_w5763_,
		_w5764_
	);
	LUT2 #(
		.INIT('h1)
	) name5233 (
		\sa02_reg[0]/P0001 ,
		_w5764_,
		_w5765_
	);
	LUT2 #(
		.INIT('h8)
	) name5234 (
		_w1016_,
		_w5130_,
		_w5766_
	);
	LUT2 #(
		.INIT('h4)
	) name5235 (
		\sa02_reg[4]/P0001 ,
		_w1025_,
		_w5767_
	);
	LUT2 #(
		.INIT('h8)
	) name5236 (
		_w982_,
		_w1000_,
		_w5768_
	);
	LUT2 #(
		.INIT('h1)
	) name5237 (
		_w5767_,
		_w5768_,
		_w5769_
	);
	LUT2 #(
		.INIT('h1)
	) name5238 (
		\sa02_reg[2]/P0001 ,
		_w5769_,
		_w5770_
	);
	LUT2 #(
		.INIT('h2)
	) name5239 (
		\sa02_reg[1]/P0001 ,
		_w5766_,
		_w5771_
	);
	LUT2 #(
		.INIT('h4)
	) name5240 (
		_w1061_,
		_w5771_,
		_w5772_
	);
	LUT2 #(
		.INIT('h4)
	) name5241 (
		_w1110_,
		_w5772_,
		_w5773_
	);
	LUT2 #(
		.INIT('h4)
	) name5242 (
		_w5770_,
		_w5773_,
		_w5774_
	);
	LUT2 #(
		.INIT('h8)
	) name5243 (
		\sa02_reg[2]/P0001 ,
		_w1001_,
		_w5775_
	);
	LUT2 #(
		.INIT('h4)
	) name5244 (
		\sa02_reg[2]/P0001 ,
		_w1091_,
		_w5776_
	);
	LUT2 #(
		.INIT('h1)
	) name5245 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w5777_
	);
	LUT2 #(
		.INIT('h1)
	) name5246 (
		\sa02_reg[3]/P0001 ,
		_w5777_,
		_w5778_
	);
	LUT2 #(
		.INIT('h2)
	) name5247 (
		_w993_,
		_w5778_,
		_w5779_
	);
	LUT2 #(
		.INIT('h8)
	) name5248 (
		_w1068_,
		_w5130_,
		_w5780_
	);
	LUT2 #(
		.INIT('h1)
	) name5249 (
		\sa02_reg[1]/P0001 ,
		_w5780_,
		_w5781_
	);
	LUT2 #(
		.INIT('h4)
	) name5250 (
		_w5775_,
		_w5781_,
		_w5782_
	);
	LUT2 #(
		.INIT('h1)
	) name5251 (
		_w5776_,
		_w5779_,
		_w5783_
	);
	LUT2 #(
		.INIT('h8)
	) name5252 (
		_w5782_,
		_w5783_,
		_w5784_
	);
	LUT2 #(
		.INIT('h1)
	) name5253 (
		_w5774_,
		_w5784_,
		_w5785_
	);
	LUT2 #(
		.INIT('h4)
	) name5254 (
		\sa02_reg[7]/NET0131 ,
		_w986_,
		_w5786_
	);
	LUT2 #(
		.INIT('h8)
	) name5255 (
		_w1023_,
		_w1035_,
		_w5787_
	);
	LUT2 #(
		.INIT('h2)
	) name5256 (
		\sa02_reg[2]/P0001 ,
		_w1109_,
		_w5788_
	);
	LUT2 #(
		.INIT('h1)
	) name5257 (
		_w5172_,
		_w5786_,
		_w5789_
	);
	LUT2 #(
		.INIT('h4)
	) name5258 (
		_w5787_,
		_w5789_,
		_w5790_
	);
	LUT2 #(
		.INIT('h8)
	) name5259 (
		_w5788_,
		_w5790_,
		_w5791_
	);
	LUT2 #(
		.INIT('h8)
	) name5260 (
		_w1019_,
		_w1035_,
		_w5792_
	);
	LUT2 #(
		.INIT('h1)
	) name5261 (
		\sa02_reg[2]/P0001 ,
		_w1069_,
		_w5793_
	);
	LUT2 #(
		.INIT('h4)
	) name5262 (
		_w5792_,
		_w5793_,
		_w5794_
	);
	LUT2 #(
		.INIT('h4)
	) name5263 (
		_w5181_,
		_w5794_,
		_w5795_
	);
	LUT2 #(
		.INIT('h1)
	) name5264 (
		_w5791_,
		_w5795_,
		_w5796_
	);
	LUT2 #(
		.INIT('h1)
	) name5265 (
		_w5785_,
		_w5796_,
		_w5797_
	);
	LUT2 #(
		.INIT('h2)
	) name5266 (
		\sa02_reg[0]/P0001 ,
		_w5797_,
		_w5798_
	);
	LUT2 #(
		.INIT('h2)
	) name5267 (
		\sa02_reg[5]/P0001 ,
		_w5326_,
		_w5799_
	);
	LUT2 #(
		.INIT('h1)
	) name5268 (
		_w986_,
		_w1059_,
		_w5800_
	);
	LUT2 #(
		.INIT('h8)
	) name5269 (
		_w1094_,
		_w5800_,
		_w5801_
	);
	LUT2 #(
		.INIT('h2)
	) name5270 (
		\sa02_reg[2]/P0001 ,
		_w5347_,
		_w5802_
	);
	LUT2 #(
		.INIT('h4)
	) name5271 (
		_w5801_,
		_w5802_,
		_w5803_
	);
	LUT2 #(
		.INIT('h4)
	) name5272 (
		_w5799_,
		_w5803_,
		_w5804_
	);
	LUT2 #(
		.INIT('h8)
	) name5273 (
		_w1004_,
		_w1030_,
		_w5805_
	);
	LUT2 #(
		.INIT('h1)
	) name5274 (
		_w1012_,
		_w5805_,
		_w5806_
	);
	LUT2 #(
		.INIT('h8)
	) name5275 (
		_w1108_,
		_w5806_,
		_w5807_
	);
	LUT2 #(
		.INIT('h1)
	) name5276 (
		_w5804_,
		_w5807_,
		_w5808_
	);
	LUT2 #(
		.INIT('h4)
	) name5277 (
		\sa02_reg[3]/P0001 ,
		_w1084_,
		_w5809_
	);
	LUT2 #(
		.INIT('h4)
	) name5278 (
		\sa02_reg[6]/NET0131 ,
		_w5809_,
		_w5810_
	);
	LUT2 #(
		.INIT('h1)
	) name5279 (
		_w5122_,
		_w5810_,
		_w5811_
	);
	LUT2 #(
		.INIT('h4)
	) name5280 (
		_w5808_,
		_w5811_,
		_w5812_
	);
	LUT2 #(
		.INIT('h1)
	) name5281 (
		\sa02_reg[1]/P0001 ,
		_w5812_,
		_w5813_
	);
	LUT2 #(
		.INIT('h1)
	) name5282 (
		\sa02_reg[2]/P0001 ,
		_w1072_,
		_w5814_
	);
	LUT2 #(
		.INIT('h2)
	) name5283 (
		\sa02_reg[2]/P0001 ,
		_w5744_,
		_w5815_
	);
	LUT2 #(
		.INIT('h2)
	) name5284 (
		\sa02_reg[3]/P0001 ,
		_w5814_,
		_w5816_
	);
	LUT2 #(
		.INIT('h4)
	) name5285 (
		_w5815_,
		_w5816_,
		_w5817_
	);
	LUT2 #(
		.INIT('h8)
	) name5286 (
		_w1059_,
		_w1094_,
		_w5818_
	);
	LUT2 #(
		.INIT('h1)
	) name5287 (
		_w977_,
		_w5142_,
		_w5819_
	);
	LUT2 #(
		.INIT('h4)
	) name5288 (
		_w5181_,
		_w5819_,
		_w5820_
	);
	LUT2 #(
		.INIT('h1)
	) name5289 (
		\sa02_reg[2]/P0001 ,
		_w5820_,
		_w5821_
	);
	LUT2 #(
		.INIT('h1)
	) name5290 (
		_w1114_,
		_w5128_,
		_w5822_
	);
	LUT2 #(
		.INIT('h1)
	) name5291 (
		_w5338_,
		_w5818_,
		_w5823_
	);
	LUT2 #(
		.INIT('h8)
	) name5292 (
		_w5822_,
		_w5823_,
		_w5824_
	);
	LUT2 #(
		.INIT('h4)
	) name5293 (
		_w5821_,
		_w5824_,
		_w5825_
	);
	LUT2 #(
		.INIT('h2)
	) name5294 (
		\sa02_reg[1]/P0001 ,
		_w5825_,
		_w5826_
	);
	LUT2 #(
		.INIT('h1)
	) name5295 (
		_w5813_,
		_w5817_,
		_w5827_
	);
	LUT2 #(
		.INIT('h4)
	) name5296 (
		_w5826_,
		_w5827_,
		_w5828_
	);
	LUT2 #(
		.INIT('h4)
	) name5297 (
		_w5798_,
		_w5828_,
		_w5829_
	);
	LUT2 #(
		.INIT('h4)
	) name5298 (
		_w5765_,
		_w5829_,
		_w5830_
	);
	LUT2 #(
		.INIT('h2)
	) name5299 (
		_w5737_,
		_w5830_,
		_w5831_
	);
	LUT2 #(
		.INIT('h4)
	) name5300 (
		_w5737_,
		_w5830_,
		_w5832_
	);
	LUT2 #(
		.INIT('h1)
	) name5301 (
		_w5831_,
		_w5832_,
		_w5833_
	);
	LUT2 #(
		.INIT('h8)
	) name5302 (
		_w722_,
		_w831_,
		_w5834_
	);
	LUT2 #(
		.INIT('h8)
	) name5303 (
		_w691_,
		_w728_,
		_w5835_
	);
	LUT2 #(
		.INIT('h2)
	) name5304 (
		\sa20_reg[2]/P0001 ,
		_w5835_,
		_w5836_
	);
	LUT2 #(
		.INIT('h2)
	) name5305 (
		\sa20_reg[6]/NET0131 ,
		_w706_,
		_w5837_
	);
	LUT2 #(
		.INIT('h2)
	) name5306 (
		_w709_,
		_w5837_,
		_w5838_
	);
	LUT2 #(
		.INIT('h8)
	) name5307 (
		_w716_,
		_w744_,
		_w5839_
	);
	LUT2 #(
		.INIT('h1)
	) name5308 (
		_w5838_,
		_w5839_,
		_w5840_
	);
	LUT2 #(
		.INIT('h8)
	) name5309 (
		_w5836_,
		_w5840_,
		_w5841_
	);
	LUT2 #(
		.INIT('h1)
	) name5310 (
		_w5834_,
		_w5841_,
		_w5842_
	);
	LUT2 #(
		.INIT('h8)
	) name5311 (
		_w705_,
		_w763_,
		_w5843_
	);
	LUT2 #(
		.INIT('h8)
	) name5312 (
		_w693_,
		_w799_,
		_w5844_
	);
	LUT2 #(
		.INIT('h1)
	) name5313 (
		\sa20_reg[2]/P0001 ,
		_w692_,
		_w5845_
	);
	LUT2 #(
		.INIT('h4)
	) name5314 (
		_w5844_,
		_w5845_,
		_w5846_
	);
	LUT2 #(
		.INIT('h2)
	) name5315 (
		\sa20_reg[2]/P0001 ,
		_w833_,
		_w5847_
	);
	LUT2 #(
		.INIT('h4)
	) name5316 (
		_w5556_,
		_w5847_,
		_w5848_
	);
	LUT2 #(
		.INIT('h1)
	) name5317 (
		_w5846_,
		_w5848_,
		_w5849_
	);
	LUT2 #(
		.INIT('h2)
	) name5318 (
		\sa20_reg[1]/P0001 ,
		_w737_,
		_w5850_
	);
	LUT2 #(
		.INIT('h1)
	) name5319 (
		_w740_,
		_w5839_,
		_w5851_
	);
	LUT2 #(
		.INIT('h4)
	) name5320 (
		_w5843_,
		_w5851_,
		_w5852_
	);
	LUT2 #(
		.INIT('h4)
	) name5321 (
		_w5613_,
		_w5850_,
		_w5853_
	);
	LUT2 #(
		.INIT('h4)
	) name5322 (
		_w5620_,
		_w5853_,
		_w5854_
	);
	LUT2 #(
		.INIT('h8)
	) name5323 (
		_w5852_,
		_w5854_,
		_w5855_
	);
	LUT2 #(
		.INIT('h4)
	) name5324 (
		_w5849_,
		_w5855_,
		_w5856_
	);
	LUT2 #(
		.INIT('h8)
	) name5325 (
		_w736_,
		_w791_,
		_w5857_
	);
	LUT2 #(
		.INIT('h8)
	) name5326 (
		\sa20_reg[6]/NET0131 ,
		_w744_,
		_w5858_
	);
	LUT2 #(
		.INIT('h8)
	) name5327 (
		_w799_,
		_w5858_,
		_w5859_
	);
	LUT2 #(
		.INIT('h8)
	) name5328 (
		_w5526_,
		_w5619_,
		_w5860_
	);
	LUT2 #(
		.INIT('h1)
	) name5329 (
		\sa20_reg[1]/P0001 ,
		_w821_,
		_w5861_
	);
	LUT2 #(
		.INIT('h1)
	) name5330 (
		_w5857_,
		_w5859_,
		_w5862_
	);
	LUT2 #(
		.INIT('h4)
	) name5331 (
		_w5860_,
		_w5862_,
		_w5863_
	);
	LUT2 #(
		.INIT('h8)
	) name5332 (
		_w5861_,
		_w5863_,
		_w5864_
	);
	LUT2 #(
		.INIT('h1)
	) name5333 (
		_w5856_,
		_w5864_,
		_w5865_
	);
	LUT2 #(
		.INIT('h1)
	) name5334 (
		\sa20_reg[0]/P0001 ,
		_w710_,
		_w5866_
	);
	LUT2 #(
		.INIT('h4)
	) name5335 (
		_w5842_,
		_w5866_,
		_w5867_
	);
	LUT2 #(
		.INIT('h4)
	) name5336 (
		_w5865_,
		_w5867_,
		_w5868_
	);
	LUT2 #(
		.INIT('h4)
	) name5337 (
		_w714_,
		_w748_,
		_w5869_
	);
	LUT2 #(
		.INIT('h1)
	) name5338 (
		_w810_,
		_w5869_,
		_w5870_
	);
	LUT2 #(
		.INIT('h2)
	) name5339 (
		\sa20_reg[1]/P0001 ,
		_w5870_,
		_w5871_
	);
	LUT2 #(
		.INIT('h8)
	) name5340 (
		_w693_,
		_w745_,
		_w5872_
	);
	LUT2 #(
		.INIT('h1)
	) name5341 (
		_w778_,
		_w5872_,
		_w5873_
	);
	LUT2 #(
		.INIT('h4)
	) name5342 (
		\sa20_reg[4]/P0001 ,
		_w777_,
		_w5874_
	);
	LUT2 #(
		.INIT('h1)
	) name5343 (
		\sa20_reg[2]/P0001 ,
		_w5874_,
		_w5875_
	);
	LUT2 #(
		.INIT('h8)
	) name5344 (
		_w5873_,
		_w5875_,
		_w5876_
	);
	LUT2 #(
		.INIT('h4)
	) name5345 (
		_w5871_,
		_w5876_,
		_w5877_
	);
	LUT2 #(
		.INIT('h8)
	) name5346 (
		_w728_,
		_w799_,
		_w5878_
	);
	LUT2 #(
		.INIT('h2)
	) name5347 (
		\sa20_reg[2]/P0001 ,
		_w703_,
		_w5879_
	);
	LUT2 #(
		.INIT('h4)
	) name5348 (
		_w5878_,
		_w5879_,
		_w5880_
	);
	LUT2 #(
		.INIT('h1)
	) name5349 (
		_w5877_,
		_w5880_,
		_w5881_
	);
	LUT2 #(
		.INIT('h8)
	) name5350 (
		_w763_,
		_w5544_,
		_w5882_
	);
	LUT2 #(
		.INIT('h4)
	) name5351 (
		\sa20_reg[4]/P0001 ,
		_w735_,
		_w5883_
	);
	LUT2 #(
		.INIT('h8)
	) name5352 (
		_w716_,
		_w723_,
		_w5884_
	);
	LUT2 #(
		.INIT('h1)
	) name5353 (
		_w5883_,
		_w5884_,
		_w5885_
	);
	LUT2 #(
		.INIT('h2)
	) name5354 (
		\sa20_reg[2]/P0001 ,
		_w5885_,
		_w5886_
	);
	LUT2 #(
		.INIT('h1)
	) name5355 (
		\sa20_reg[1]/P0001 ,
		_w778_,
		_w5887_
	);
	LUT2 #(
		.INIT('h4)
	) name5356 (
		_w5524_,
		_w5887_,
		_w5888_
	);
	LUT2 #(
		.INIT('h1)
	) name5357 (
		_w703_,
		_w5882_,
		_w5889_
	);
	LUT2 #(
		.INIT('h8)
	) name5358 (
		_w5888_,
		_w5889_,
		_w5890_
	);
	LUT2 #(
		.INIT('h4)
	) name5359 (
		_w5886_,
		_w5890_,
		_w5891_
	);
	LUT2 #(
		.INIT('h4)
	) name5360 (
		\sa20_reg[3]/P0001 ,
		_w715_,
		_w5892_
	);
	LUT2 #(
		.INIT('h1)
	) name5361 (
		_w752_,
		_w5892_,
		_w5893_
	);
	LUT2 #(
		.INIT('h8)
	) name5362 (
		_w691_,
		_w820_,
		_w5894_
	);
	LUT2 #(
		.INIT('h8)
	) name5363 (
		_w705_,
		_w745_,
		_w5895_
	);
	LUT2 #(
		.INIT('h2)
	) name5364 (
		\sa20_reg[1]/P0001 ,
		_w5895_,
		_w5896_
	);
	LUT2 #(
		.INIT('h4)
	) name5365 (
		_w5894_,
		_w5896_,
		_w5897_
	);
	LUT2 #(
		.INIT('h8)
	) name5366 (
		_w5893_,
		_w5897_,
		_w5898_
	);
	LUT2 #(
		.INIT('h1)
	) name5367 (
		_w5891_,
		_w5898_,
		_w5899_
	);
	LUT2 #(
		.INIT('h8)
	) name5368 (
		_w5523_,
		_w5585_,
		_w5900_
	);
	LUT2 #(
		.INIT('h8)
	) name5369 (
		_w694_,
		_w699_,
		_w5901_
	);
	LUT2 #(
		.INIT('h2)
	) name5370 (
		\sa20_reg[0]/P0001 ,
		_w5900_,
		_w5902_
	);
	LUT2 #(
		.INIT('h4)
	) name5371 (
		_w5901_,
		_w5902_,
		_w5903_
	);
	LUT2 #(
		.INIT('h4)
	) name5372 (
		_w5881_,
		_w5903_,
		_w5904_
	);
	LUT2 #(
		.INIT('h4)
	) name5373 (
		_w5899_,
		_w5904_,
		_w5905_
	);
	LUT2 #(
		.INIT('h1)
	) name5374 (
		_w5868_,
		_w5905_,
		_w5906_
	);
	LUT2 #(
		.INIT('h8)
	) name5375 (
		_w714_,
		_w735_,
		_w5907_
	);
	LUT2 #(
		.INIT('h8)
	) name5376 (
		_w694_,
		_w736_,
		_w5908_
	);
	LUT2 #(
		.INIT('h1)
	) name5377 (
		_w5907_,
		_w5908_,
		_w5909_
	);
	LUT2 #(
		.INIT('h4)
	) name5378 (
		_w779_,
		_w5909_,
		_w5910_
	);
	LUT2 #(
		.INIT('h1)
	) name5379 (
		\sa20_reg[1]/P0001 ,
		_w5910_,
		_w5911_
	);
	LUT2 #(
		.INIT('h1)
	) name5380 (
		_w737_,
		_w817_,
		_w5912_
	);
	LUT2 #(
		.INIT('h4)
	) name5381 (
		_w5911_,
		_w5912_,
		_w5913_
	);
	LUT2 #(
		.INIT('h1)
	) name5382 (
		\sa20_reg[2]/P0001 ,
		_w5913_,
		_w5914_
	);
	LUT2 #(
		.INIT('h8)
	) name5383 (
		\sa20_reg[3]/P0001 ,
		_w710_,
		_w5915_
	);
	LUT2 #(
		.INIT('h2)
	) name5384 (
		\sa20_reg[2]/P0001 ,
		_w790_,
		_w5916_
	);
	LUT2 #(
		.INIT('h1)
	) name5385 (
		_w831_,
		_w5916_,
		_w5917_
	);
	LUT2 #(
		.INIT('h2)
	) name5386 (
		\sa20_reg[1]/P0001 ,
		_w5915_,
		_w5918_
	);
	LUT2 #(
		.INIT('h4)
	) name5387 (
		_w5917_,
		_w5918_,
		_w5919_
	);
	LUT2 #(
		.INIT('h1)
	) name5388 (
		_w728_,
		_w5544_,
		_w5920_
	);
	LUT2 #(
		.INIT('h4)
	) name5389 (
		_w5858_,
		_w5920_,
		_w5921_
	);
	LUT2 #(
		.INIT('h2)
	) name5390 (
		_w691_,
		_w5921_,
		_w5922_
	);
	LUT2 #(
		.INIT('h1)
	) name5391 (
		_w751_,
		_w5922_,
		_w5923_
	);
	LUT2 #(
		.INIT('h2)
	) name5392 (
		\sa20_reg[2]/P0001 ,
		_w5923_,
		_w5924_
	);
	LUT2 #(
		.INIT('h1)
	) name5393 (
		\sa20_reg[1]/P0001 ,
		_w809_,
		_w5925_
	);
	LUT2 #(
		.INIT('h4)
	) name5394 (
		_w5924_,
		_w5925_,
		_w5926_
	);
	LUT2 #(
		.INIT('h1)
	) name5395 (
		_w5919_,
		_w5926_,
		_w5927_
	);
	LUT2 #(
		.INIT('h8)
	) name5396 (
		_w761_,
		_w5606_,
		_w5928_
	);
	LUT2 #(
		.INIT('h1)
	) name5397 (
		_w5914_,
		_w5928_,
		_w5929_
	);
	LUT2 #(
		.INIT('h4)
	) name5398 (
		_w5927_,
		_w5929_,
		_w5930_
	);
	LUT2 #(
		.INIT('h4)
	) name5399 (
		_w5906_,
		_w5930_,
		_w5931_
	);
	LUT2 #(
		.INIT('h2)
	) name5400 (
		_w973_,
		_w5931_,
		_w5932_
	);
	LUT2 #(
		.INIT('h4)
	) name5401 (
		_w973_,
		_w5931_,
		_w5933_
	);
	LUT2 #(
		.INIT('h1)
	) name5402 (
		_w5932_,
		_w5933_,
		_w5934_
	);
	LUT2 #(
		.INIT('h2)
	) name5403 (
		\u0_w_reg[2][29]/P0001 ,
		_w5307_,
		_w5935_
	);
	LUT2 #(
		.INIT('h4)
	) name5404 (
		\u0_w_reg[2][29]/P0001 ,
		_w5307_,
		_w5936_
	);
	LUT2 #(
		.INIT('h1)
	) name5405 (
		_w5935_,
		_w5936_,
		_w5937_
	);
	LUT2 #(
		.INIT('h8)
	) name5406 (
		_w5934_,
		_w5937_,
		_w5938_
	);
	LUT2 #(
		.INIT('h1)
	) name5407 (
		_w5934_,
		_w5937_,
		_w5939_
	);
	LUT2 #(
		.INIT('h1)
	) name5408 (
		_w5938_,
		_w5939_,
		_w5940_
	);
	LUT2 #(
		.INIT('h4)
	) name5409 (
		_w5833_,
		_w5940_,
		_w5941_
	);
	LUT2 #(
		.INIT('h2)
	) name5410 (
		_w5833_,
		_w5940_,
		_w5942_
	);
	LUT2 #(
		.INIT('h1)
	) name5411 (
		\ld_r_reg/P0001 ,
		_w5941_,
		_w5943_
	);
	LUT2 #(
		.INIT('h4)
	) name5412 (
		_w5942_,
		_w5943_,
		_w5944_
	);
	LUT2 #(
		.INIT('h2)
	) name5413 (
		\text_in_r_reg[61]/P0001 ,
		\u0_w_reg[2][29]/P0001 ,
		_w5945_
	);
	LUT2 #(
		.INIT('h4)
	) name5414 (
		\text_in_r_reg[61]/P0001 ,
		\u0_w_reg[2][29]/P0001 ,
		_w5946_
	);
	LUT2 #(
		.INIT('h2)
	) name5415 (
		\ld_r_reg/P0001 ,
		_w5945_,
		_w5947_
	);
	LUT2 #(
		.INIT('h4)
	) name5416 (
		_w5946_,
		_w5947_,
		_w5948_
	);
	LUT2 #(
		.INIT('h1)
	) name5417 (
		_w5944_,
		_w5948_,
		_w5949_
	);
	LUT2 #(
		.INIT('h1)
	) name5418 (
		_w5191_,
		_w5934_,
		_w5950_
	);
	LUT2 #(
		.INIT('h8)
	) name5419 (
		_w5191_,
		_w5934_,
		_w5951_
	);
	LUT2 #(
		.INIT('h1)
	) name5420 (
		_w5950_,
		_w5951_,
		_w5952_
	);
	LUT2 #(
		.INIT('h2)
	) name5421 (
		\u0_w_reg[2][22]/P0001 ,
		_w1300_,
		_w5953_
	);
	LUT2 #(
		.INIT('h4)
	) name5422 (
		\u0_w_reg[2][22]/P0001 ,
		_w1300_,
		_w5954_
	);
	LUT2 #(
		.INIT('h1)
	) name5423 (
		_w5953_,
		_w5954_,
		_w5955_
	);
	LUT2 #(
		.INIT('h8)
	) name5424 (
		_w850_,
		_w5955_,
		_w5956_
	);
	LUT2 #(
		.INIT('h1)
	) name5425 (
		_w850_,
		_w5955_,
		_w5957_
	);
	LUT2 #(
		.INIT('h1)
	) name5426 (
		_w5956_,
		_w5957_,
		_w5958_
	);
	LUT2 #(
		.INIT('h1)
	) name5427 (
		_w5952_,
		_w5958_,
		_w5959_
	);
	LUT2 #(
		.INIT('h8)
	) name5428 (
		_w5952_,
		_w5958_,
		_w5960_
	);
	LUT2 #(
		.INIT('h1)
	) name5429 (
		\ld_r_reg/P0001 ,
		_w5959_,
		_w5961_
	);
	LUT2 #(
		.INIT('h4)
	) name5430 (
		_w5960_,
		_w5961_,
		_w5962_
	);
	LUT2 #(
		.INIT('h2)
	) name5431 (
		\text_in_r_reg[54]/P0001 ,
		\u0_w_reg[2][22]/P0001 ,
		_w5963_
	);
	LUT2 #(
		.INIT('h4)
	) name5432 (
		\text_in_r_reg[54]/P0001 ,
		\u0_w_reg[2][22]/P0001 ,
		_w5964_
	);
	LUT2 #(
		.INIT('h2)
	) name5433 (
		\ld_r_reg/P0001 ,
		_w5963_,
		_w5965_
	);
	LUT2 #(
		.INIT('h4)
	) name5434 (
		_w5964_,
		_w5965_,
		_w5966_
	);
	LUT2 #(
		.INIT('h1)
	) name5435 (
		_w5962_,
		_w5966_,
		_w5967_
	);
	LUT2 #(
		.INIT('h8)
	) name5436 (
		_w724_,
		_w799_,
		_w5968_
	);
	LUT2 #(
		.INIT('h1)
	) name5437 (
		_w5541_,
		_w5900_,
		_w5969_
	);
	LUT2 #(
		.INIT('h1)
	) name5438 (
		\sa20_reg[3]/P0001 ,
		_w5969_,
		_w5970_
	);
	LUT2 #(
		.INIT('h8)
	) name5439 (
		_w716_,
		_w5581_,
		_w5971_
	);
	LUT2 #(
		.INIT('h8)
	) name5440 (
		\sa20_reg[2]/P0001 ,
		_w5532_,
		_w5972_
	);
	LUT2 #(
		.INIT('h8)
	) name5441 (
		\sa20_reg[5]/P0001 ,
		_w5527_,
		_w5973_
	);
	LUT2 #(
		.INIT('h4)
	) name5442 (
		\sa20_reg[2]/P0001 ,
		_w5973_,
		_w5974_
	);
	LUT2 #(
		.INIT('h1)
	) name5443 (
		_w829_,
		_w5581_,
		_w5975_
	);
	LUT2 #(
		.INIT('h4)
	) name5444 (
		_w5972_,
		_w5975_,
		_w5976_
	);
	LUT2 #(
		.INIT('h4)
	) name5445 (
		_w5974_,
		_w5976_,
		_w5977_
	);
	LUT2 #(
		.INIT('h1)
	) name5446 (
		\sa20_reg[1]/P0001 ,
		_w5977_,
		_w5978_
	);
	LUT2 #(
		.INIT('h8)
	) name5447 (
		\sa20_reg[5]/P0001 ,
		_w705_,
		_w5979_
	);
	LUT2 #(
		.INIT('h4)
	) name5448 (
		_w745_,
		_w5979_,
		_w5980_
	);
	LUT2 #(
		.INIT('h8)
	) name5449 (
		_w708_,
		_w765_,
		_w5981_
	);
	LUT2 #(
		.INIT('h1)
	) name5450 (
		_w5980_,
		_w5981_,
		_w5982_
	);
	LUT2 #(
		.INIT('h1)
	) name5451 (
		\sa20_reg[2]/P0001 ,
		_w5982_,
		_w5983_
	);
	LUT2 #(
		.INIT('h2)
	) name5452 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w5984_
	);
	LUT2 #(
		.INIT('h8)
	) name5453 (
		_w701_,
		_w5984_,
		_w5985_
	);
	LUT2 #(
		.INIT('h8)
	) name5454 (
		_w819_,
		_w5585_,
		_w5986_
	);
	LUT2 #(
		.INIT('h1)
	) name5455 (
		_w700_,
		_w5985_,
		_w5987_
	);
	LUT2 #(
		.INIT('h4)
	) name5456 (
		_w5986_,
		_w5987_,
		_w5988_
	);
	LUT2 #(
		.INIT('h4)
	) name5457 (
		_w5983_,
		_w5988_,
		_w5989_
	);
	LUT2 #(
		.INIT('h2)
	) name5458 (
		\sa20_reg[1]/P0001 ,
		_w5989_,
		_w5990_
	);
	LUT2 #(
		.INIT('h1)
	) name5459 (
		_w5968_,
		_w5971_,
		_w5991_
	);
	LUT2 #(
		.INIT('h4)
	) name5460 (
		_w5970_,
		_w5991_,
		_w5992_
	);
	LUT2 #(
		.INIT('h4)
	) name5461 (
		_w5978_,
		_w5992_,
		_w5993_
	);
	LUT2 #(
		.INIT('h4)
	) name5462 (
		_w5990_,
		_w5993_,
		_w5994_
	);
	LUT2 #(
		.INIT('h1)
	) name5463 (
		\sa20_reg[0]/P0001 ,
		_w5994_,
		_w5995_
	);
	LUT2 #(
		.INIT('h2)
	) name5464 (
		\sa20_reg[1]/P0001 ,
		_w817_,
		_w5996_
	);
	LUT2 #(
		.INIT('h4)
	) name5465 (
		\sa20_reg[4]/P0001 ,
		_w693_,
		_w5997_
	);
	LUT2 #(
		.INIT('h8)
	) name5466 (
		_w708_,
		_w714_,
		_w5998_
	);
	LUT2 #(
		.INIT('h1)
	) name5467 (
		_w5997_,
		_w5998_,
		_w5999_
	);
	LUT2 #(
		.INIT('h1)
	) name5468 (
		\sa20_reg[2]/P0001 ,
		_w5999_,
		_w6000_
	);
	LUT2 #(
		.INIT('h8)
	) name5469 (
		_w705_,
		_w5526_,
		_w6001_
	);
	LUT2 #(
		.INIT('h1)
	) name5470 (
		_w5894_,
		_w6001_,
		_w6002_
	);
	LUT2 #(
		.INIT('h8)
	) name5471 (
		_w5996_,
		_w6002_,
		_w6003_
	);
	LUT2 #(
		.INIT('h4)
	) name5472 (
		_w6000_,
		_w6003_,
		_w6004_
	);
	LUT2 #(
		.INIT('h8)
	) name5473 (
		_w745_,
		_w826_,
		_w6005_
	);
	LUT2 #(
		.INIT('h1)
	) name5474 (
		\sa20_reg[1]/P0001 ,
		_w6005_,
		_w6006_
	);
	LUT2 #(
		.INIT('h8)
	) name5475 (
		_w763_,
		_w807_,
		_w6007_
	);
	LUT2 #(
		.INIT('h8)
	) name5476 (
		\sa20_reg[2]/P0001 ,
		_w715_,
		_w6008_
	);
	LUT2 #(
		.INIT('h1)
	) name5477 (
		\sa20_reg[3]/P0001 ,
		_w5582_,
		_w6009_
	);
	LUT2 #(
		.INIT('h2)
	) name5478 (
		_w744_,
		_w6009_,
		_w6010_
	);
	LUT2 #(
		.INIT('h2)
	) name5479 (
		_w6006_,
		_w6007_,
		_w6011_
	);
	LUT2 #(
		.INIT('h1)
	) name5480 (
		_w6008_,
		_w6010_,
		_w6012_
	);
	LUT2 #(
		.INIT('h8)
	) name5481 (
		_w6011_,
		_w6012_,
		_w6013_
	);
	LUT2 #(
		.INIT('h1)
	) name5482 (
		_w6004_,
		_w6013_,
		_w6014_
	);
	LUT2 #(
		.INIT('h2)
	) name5483 (
		_w796_,
		_w5872_,
		_w6015_
	);
	LUT2 #(
		.INIT('h4)
	) name5484 (
		_w824_,
		_w6015_,
		_w6016_
	);
	LUT2 #(
		.INIT('h1)
	) name5485 (
		_w707_,
		_w789_,
		_w6017_
	);
	LUT2 #(
		.INIT('h4)
	) name5486 (
		_w816_,
		_w6017_,
		_w6018_
	);
	LUT2 #(
		.INIT('h8)
	) name5487 (
		_w828_,
		_w6018_,
		_w6019_
	);
	LUT2 #(
		.INIT('h1)
	) name5488 (
		_w6016_,
		_w6019_,
		_w6020_
	);
	LUT2 #(
		.INIT('h1)
	) name5489 (
		_w6014_,
		_w6020_,
		_w6021_
	);
	LUT2 #(
		.INIT('h2)
	) name5490 (
		\sa20_reg[0]/P0001 ,
		_w6021_,
		_w6022_
	);
	LUT2 #(
		.INIT('h8)
	) name5491 (
		_w782_,
		_w5523_,
		_w6023_
	);
	LUT2 #(
		.INIT('h1)
	) name5492 (
		_w5972_,
		_w6023_,
		_w6024_
	);
	LUT2 #(
		.INIT('h2)
	) name5493 (
		\sa20_reg[3]/P0001 ,
		_w6024_,
		_w6025_
	);
	LUT2 #(
		.INIT('h1)
	) name5494 (
		_w792_,
		_w824_,
		_w6026_
	);
	LUT2 #(
		.INIT('h4)
	) name5495 (
		_w5859_,
		_w6026_,
		_w6027_
	);
	LUT2 #(
		.INIT('h1)
	) name5496 (
		\sa20_reg[2]/P0001 ,
		_w6027_,
		_w6028_
	);
	LUT2 #(
		.INIT('h4)
	) name5497 (
		\sa20_reg[5]/P0001 ,
		_w5895_,
		_w6029_
	);
	LUT2 #(
		.INIT('h8)
	) name5498 (
		_w739_,
		_w819_,
		_w6030_
	);
	LUT2 #(
		.INIT('h1)
	) name5499 (
		_w762_,
		_w5543_,
		_w6031_
	);
	LUT2 #(
		.INIT('h1)
	) name5500 (
		_w6029_,
		_w6030_,
		_w6032_
	);
	LUT2 #(
		.INIT('h8)
	) name5501 (
		_w6031_,
		_w6032_,
		_w6033_
	);
	LUT2 #(
		.INIT('h4)
	) name5502 (
		_w6028_,
		_w6033_,
		_w6034_
	);
	LUT2 #(
		.INIT('h2)
	) name5503 (
		\sa20_reg[1]/P0001 ,
		_w6034_,
		_w6035_
	);
	LUT2 #(
		.INIT('h8)
	) name5504 (
		_w714_,
		_w5619_,
		_w6036_
	);
	LUT2 #(
		.INIT('h8)
	) name5505 (
		\sa20_reg[7]/NET0131 ,
		_w800_,
		_w6037_
	);
	LUT2 #(
		.INIT('h2)
	) name5506 (
		\sa20_reg[2]/P0001 ,
		_w778_,
		_w6038_
	);
	LUT2 #(
		.INIT('h4)
	) name5507 (
		_w5525_,
		_w6038_,
		_w6039_
	);
	LUT2 #(
		.INIT('h1)
	) name5508 (
		_w725_,
		_w6036_,
		_w6040_
	);
	LUT2 #(
		.INIT('h4)
	) name5509 (
		_w6037_,
		_w6040_,
		_w6041_
	);
	LUT2 #(
		.INIT('h8)
	) name5510 (
		_w6039_,
		_w6041_,
		_w6042_
	);
	LUT2 #(
		.INIT('h8)
	) name5511 (
		_w810_,
		_w826_,
		_w6043_
	);
	LUT2 #(
		.INIT('h1)
	) name5512 (
		\sa20_reg[3]/P0001 ,
		_w709_,
		_w6044_
	);
	LUT2 #(
		.INIT('h8)
	) name5513 (
		_w735_,
		_w6044_,
		_w6045_
	);
	LUT2 #(
		.INIT('h1)
	) name5514 (
		\sa20_reg[2]/P0001 ,
		_w779_,
		_w6046_
	);
	LUT2 #(
		.INIT('h1)
	) name5515 (
		_w6043_,
		_w6045_,
		_w6047_
	);
	LUT2 #(
		.INIT('h8)
	) name5516 (
		_w6046_,
		_w6047_,
		_w6048_
	);
	LUT2 #(
		.INIT('h1)
	) name5517 (
		_w6042_,
		_w6048_,
		_w6049_
	);
	LUT2 #(
		.INIT('h1)
	) name5518 (
		_w5968_,
		_w6049_,
		_w6050_
	);
	LUT2 #(
		.INIT('h1)
	) name5519 (
		\sa20_reg[1]/P0001 ,
		_w6050_,
		_w6051_
	);
	LUT2 #(
		.INIT('h1)
	) name5520 (
		_w6025_,
		_w6035_,
		_w6052_
	);
	LUT2 #(
		.INIT('h4)
	) name5521 (
		_w6022_,
		_w6052_,
		_w6053_
	);
	LUT2 #(
		.INIT('h4)
	) name5522 (
		_w6051_,
		_w6053_,
		_w6054_
	);
	LUT2 #(
		.INIT('h4)
	) name5523 (
		_w5995_,
		_w6054_,
		_w6055_
	);
	LUT2 #(
		.INIT('h2)
	) name5524 (
		_w5737_,
		_w6055_,
		_w6056_
	);
	LUT2 #(
		.INIT('h4)
	) name5525 (
		_w5737_,
		_w6055_,
		_w6057_
	);
	LUT2 #(
		.INIT('h1)
	) name5526 (
		_w6056_,
		_w6057_,
		_w6058_
	);
	LUT2 #(
		.INIT('h1)
	) name5527 (
		_w1142_,
		_w6058_,
		_w6059_
	);
	LUT2 #(
		.INIT('h8)
	) name5528 (
		_w1142_,
		_w6058_,
		_w6060_
	);
	LUT2 #(
		.INIT('h1)
	) name5529 (
		_w6059_,
		_w6060_,
		_w6061_
	);
	LUT2 #(
		.INIT('h2)
	) name5530 (
		\u0_w_reg[2][21]/P0001 ,
		_w5307_,
		_w6062_
	);
	LUT2 #(
		.INIT('h4)
	) name5531 (
		\u0_w_reg[2][21]/P0001 ,
		_w5307_,
		_w6063_
	);
	LUT2 #(
		.INIT('h1)
	) name5532 (
		_w6062_,
		_w6063_,
		_w6064_
	);
	LUT2 #(
		.INIT('h8)
	) name5533 (
		_w5931_,
		_w6064_,
		_w6065_
	);
	LUT2 #(
		.INIT('h1)
	) name5534 (
		_w5931_,
		_w6064_,
		_w6066_
	);
	LUT2 #(
		.INIT('h1)
	) name5535 (
		_w6065_,
		_w6066_,
		_w6067_
	);
	LUT2 #(
		.INIT('h1)
	) name5536 (
		_w6061_,
		_w6067_,
		_w6068_
	);
	LUT2 #(
		.INIT('h8)
	) name5537 (
		_w6061_,
		_w6067_,
		_w6069_
	);
	LUT2 #(
		.INIT('h1)
	) name5538 (
		\ld_r_reg/P0001 ,
		_w6068_,
		_w6070_
	);
	LUT2 #(
		.INIT('h4)
	) name5539 (
		_w6069_,
		_w6070_,
		_w6071_
	);
	LUT2 #(
		.INIT('h2)
	) name5540 (
		\text_in_r_reg[53]/P0001 ,
		\u0_w_reg[2][21]/P0001 ,
		_w6072_
	);
	LUT2 #(
		.INIT('h4)
	) name5541 (
		\text_in_r_reg[53]/P0001 ,
		\u0_w_reg[2][21]/P0001 ,
		_w6073_
	);
	LUT2 #(
		.INIT('h2)
	) name5542 (
		\ld_r_reg/P0001 ,
		_w6072_,
		_w6074_
	);
	LUT2 #(
		.INIT('h4)
	) name5543 (
		_w6073_,
		_w6074_,
		_w6075_
	);
	LUT2 #(
		.INIT('h1)
	) name5544 (
		_w6071_,
		_w6075_,
		_w6076_
	);
	LUT2 #(
		.INIT('h1)
	) name5545 (
		_w1145_,
		_w6055_,
		_w6077_
	);
	LUT2 #(
		.INIT('h8)
	) name5546 (
		_w1145_,
		_w6055_,
		_w6078_
	);
	LUT2 #(
		.INIT('h1)
	) name5547 (
		_w6077_,
		_w6078_,
		_w6079_
	);
	LUT2 #(
		.INIT('h4)
	) name5548 (
		\sa31_reg[6]/NET0131 ,
		_w1181_,
		_w6080_
	);
	LUT2 #(
		.INIT('h4)
	) name5549 (
		\sa31_reg[3]/P0001 ,
		_w5241_,
		_w6081_
	);
	LUT2 #(
		.INIT('h1)
	) name5550 (
		_w6080_,
		_w6081_,
		_w6082_
	);
	LUT2 #(
		.INIT('h2)
	) name5551 (
		\sa31_reg[2]/P0001 ,
		_w6082_,
		_w6083_
	);
	LUT2 #(
		.INIT('h4)
	) name5552 (
		\sa31_reg[6]/NET0131 ,
		_w5268_,
		_w6084_
	);
	LUT2 #(
		.INIT('h1)
	) name5553 (
		_w5262_,
		_w6084_,
		_w6085_
	);
	LUT2 #(
		.INIT('h1)
	) name5554 (
		\sa31_reg[3]/P0001 ,
		_w6085_,
		_w6086_
	);
	LUT2 #(
		.INIT('h8)
	) name5555 (
		\sa31_reg[2]/P0001 ,
		_w1194_,
		_w6087_
	);
	LUT2 #(
		.INIT('h2)
	) name5556 (
		_w1147_,
		_w1225_,
		_w6088_
	);
	LUT2 #(
		.INIT('h4)
	) name5557 (
		\sa31_reg[4]/P0001 ,
		_w5239_,
		_w6089_
	);
	LUT2 #(
		.INIT('h1)
	) name5558 (
		_w6088_,
		_w6089_,
		_w6090_
	);
	LUT2 #(
		.INIT('h1)
	) name5559 (
		\sa31_reg[2]/P0001 ,
		_w6090_,
		_w6091_
	);
	LUT2 #(
		.INIT('h8)
	) name5560 (
		\sa31_reg[4]/P0001 ,
		_w1182_,
		_w6092_
	);
	LUT2 #(
		.INIT('h8)
	) name5561 (
		_w1279_,
		_w6092_,
		_w6093_
	);
	LUT2 #(
		.INIT('h2)
	) name5562 (
		\sa31_reg[1]/P0001 ,
		_w1200_,
		_w6094_
	);
	LUT2 #(
		.INIT('h1)
	) name5563 (
		_w6087_,
		_w6093_,
		_w6095_
	);
	LUT2 #(
		.INIT('h8)
	) name5564 (
		_w6094_,
		_w6095_,
		_w6096_
	);
	LUT2 #(
		.INIT('h4)
	) name5565 (
		_w6091_,
		_w6096_,
		_w6097_
	);
	LUT2 #(
		.INIT('h8)
	) name5566 (
		\sa31_reg[2]/P0001 ,
		_w1219_,
		_w6098_
	);
	LUT2 #(
		.INIT('h1)
	) name5567 (
		\sa31_reg[1]/P0001 ,
		_w6098_,
		_w6099_
	);
	LUT2 #(
		.INIT('h8)
	) name5568 (
		_w1162_,
		_w1193_,
		_w6100_
	);
	LUT2 #(
		.INIT('h1)
	) name5569 (
		_w1226_,
		_w6100_,
		_w6101_
	);
	LUT2 #(
		.INIT('h1)
	) name5570 (
		\sa31_reg[7]/P0001 ,
		_w6101_,
		_w6102_
	);
	LUT2 #(
		.INIT('h8)
	) name5571 (
		\sa31_reg[2]/P0001 ,
		_w1277_,
		_w6103_
	);
	LUT2 #(
		.INIT('h2)
	) name5572 (
		_w6099_,
		_w6103_,
		_w6104_
	);
	LUT2 #(
		.INIT('h4)
	) name5573 (
		_w6102_,
		_w6104_,
		_w6105_
	);
	LUT2 #(
		.INIT('h1)
	) name5574 (
		_w6097_,
		_w6105_,
		_w6106_
	);
	LUT2 #(
		.INIT('h1)
	) name5575 (
		_w6083_,
		_w6086_,
		_w6107_
	);
	LUT2 #(
		.INIT('h4)
	) name5576 (
		_w6106_,
		_w6107_,
		_w6108_
	);
	LUT2 #(
		.INIT('h1)
	) name5577 (
		\sa31_reg[0]/P0002 ,
		_w6108_,
		_w6109_
	);
	LUT2 #(
		.INIT('h8)
	) name5578 (
		_w1163_,
		_w1180_,
		_w6110_
	);
	LUT2 #(
		.INIT('h4)
	) name5579 (
		\sa31_reg[2]/P0001 ,
		_w6110_,
		_w6111_
	);
	LUT2 #(
		.INIT('h1)
	) name5580 (
		_w6103_,
		_w6111_,
		_w6112_
	);
	LUT2 #(
		.INIT('h2)
	) name5581 (
		\sa31_reg[3]/P0001 ,
		_w6112_,
		_w6113_
	);
	LUT2 #(
		.INIT('h2)
	) name5582 (
		\sa31_reg[2]/P0001 ,
		_w1207_,
		_w6114_
	);
	LUT2 #(
		.INIT('h8)
	) name5583 (
		_w1163_,
		_w1166_,
		_w6115_
	);
	LUT2 #(
		.INIT('h1)
	) name5584 (
		_w1226_,
		_w5252_,
		_w6116_
	);
	LUT2 #(
		.INIT('h4)
	) name5585 (
		_w6115_,
		_w6116_,
		_w6117_
	);
	LUT2 #(
		.INIT('h8)
	) name5586 (
		_w6114_,
		_w6117_,
		_w6118_
	);
	LUT2 #(
		.INIT('h8)
	) name5587 (
		_w1182_,
		_w5269_,
		_w6119_
	);
	LUT2 #(
		.INIT('h1)
	) name5588 (
		\sa31_reg[2]/P0001 ,
		_w5271_,
		_w6120_
	);
	LUT2 #(
		.INIT('h4)
	) name5589 (
		_w6119_,
		_w6120_,
		_w6121_
	);
	LUT2 #(
		.INIT('h4)
	) name5590 (
		_w1231_,
		_w6121_,
		_w6122_
	);
	LUT2 #(
		.INIT('h1)
	) name5591 (
		_w6118_,
		_w6122_,
		_w6123_
	);
	LUT2 #(
		.INIT('h4)
	) name5592 (
		\sa31_reg[6]/NET0131 ,
		_w6092_,
		_w6124_
	);
	LUT2 #(
		.INIT('h1)
	) name5593 (
		_w5199_,
		_w6124_,
		_w6125_
	);
	LUT2 #(
		.INIT('h1)
	) name5594 (
		\sa31_reg[2]/P0001 ,
		_w6125_,
		_w6126_
	);
	LUT2 #(
		.INIT('h8)
	) name5595 (
		_w1146_,
		_w1244_,
		_w6127_
	);
	LUT2 #(
		.INIT('h2)
	) name5596 (
		\sa31_reg[1]/P0001 ,
		_w6127_,
		_w6128_
	);
	LUT2 #(
		.INIT('h4)
	) name5597 (
		_w1227_,
		_w6128_,
		_w6129_
	);
	LUT2 #(
		.INIT('h4)
	) name5598 (
		_w5253_,
		_w6129_,
		_w6130_
	);
	LUT2 #(
		.INIT('h4)
	) name5599 (
		_w6126_,
		_w6130_,
		_w6131_
	);
	LUT2 #(
		.INIT('h4)
	) name5600 (
		\sa31_reg[2]/P0001 ,
		_w5242_,
		_w6132_
	);
	LUT2 #(
		.INIT('h1)
	) name5601 (
		\sa31_reg[1]/P0001 ,
		_w6132_,
		_w6133_
	);
	LUT2 #(
		.INIT('h8)
	) name5602 (
		_w1225_,
		_w1256_,
		_w6134_
	);
	LUT2 #(
		.INIT('h8)
	) name5603 (
		\sa31_reg[2]/P0001 ,
		_w1179_,
		_w6135_
	);
	LUT2 #(
		.INIT('h1)
	) name5604 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w6136_
	);
	LUT2 #(
		.INIT('h1)
	) name5605 (
		\sa31_reg[3]/P0001 ,
		_w6136_,
		_w6137_
	);
	LUT2 #(
		.INIT('h2)
	) name5606 (
		_w1166_,
		_w6137_,
		_w6138_
	);
	LUT2 #(
		.INIT('h1)
	) name5607 (
		_w6134_,
		_w6135_,
		_w6139_
	);
	LUT2 #(
		.INIT('h4)
	) name5608 (
		_w6138_,
		_w6139_,
		_w6140_
	);
	LUT2 #(
		.INIT('h8)
	) name5609 (
		_w6133_,
		_w6140_,
		_w6141_
	);
	LUT2 #(
		.INIT('h1)
	) name5610 (
		_w6131_,
		_w6141_,
		_w6142_
	);
	LUT2 #(
		.INIT('h1)
	) name5611 (
		_w6123_,
		_w6142_,
		_w6143_
	);
	LUT2 #(
		.INIT('h2)
	) name5612 (
		\sa31_reg[0]/P0002 ,
		_w6143_,
		_w6144_
	);
	LUT2 #(
		.INIT('h8)
	) name5613 (
		_w1225_,
		_w5239_,
		_w6145_
	);
	LUT2 #(
		.INIT('h8)
	) name5614 (
		_w1149_,
		_w1279_,
		_w6146_
	);
	LUT2 #(
		.INIT('h8)
	) name5615 (
		\sa31_reg[4]/P0001 ,
		_w6146_,
		_w6147_
	);
	LUT2 #(
		.INIT('h8)
	) name5616 (
		\sa31_reg[7]/P0001 ,
		_w1247_,
		_w6148_
	);
	LUT2 #(
		.INIT('h1)
	) name5617 (
		_w1231_,
		_w1258_,
		_w6149_
	);
	LUT2 #(
		.INIT('h4)
	) name5618 (
		_w6148_,
		_w6149_,
		_w6150_
	);
	LUT2 #(
		.INIT('h1)
	) name5619 (
		\sa31_reg[2]/P0001 ,
		_w6150_,
		_w6151_
	);
	LUT2 #(
		.INIT('h8)
	) name5620 (
		_w1159_,
		_w1256_,
		_w6152_
	);
	LUT2 #(
		.INIT('h4)
	) name5621 (
		\sa31_reg[5]/P0001 ,
		_w6152_,
		_w6153_
	);
	LUT2 #(
		.INIT('h2)
	) name5622 (
		\sa31_reg[1]/P0001 ,
		_w1266_,
		_w6154_
	);
	LUT2 #(
		.INIT('h1)
	) name5623 (
		_w6145_,
		_w6147_,
		_w6155_
	);
	LUT2 #(
		.INIT('h4)
	) name5624 (
		_w6153_,
		_w6155_,
		_w6156_
	);
	LUT2 #(
		.INIT('h8)
	) name5625 (
		_w6154_,
		_w6156_,
		_w6157_
	);
	LUT2 #(
		.INIT('h4)
	) name5626 (
		_w6151_,
		_w6157_,
		_w6158_
	);
	LUT2 #(
		.INIT('h8)
	) name5627 (
		_w1178_,
		_w1230_,
		_w6159_
	);
	LUT2 #(
		.INIT('h8)
	) name5628 (
		_w1256_,
		_w5263_,
		_w6160_
	);
	LUT2 #(
		.INIT('h1)
	) name5629 (
		\sa31_reg[2]/P0001 ,
		_w6160_,
		_w6161_
	);
	LUT2 #(
		.INIT('h4)
	) name5630 (
		\sa31_reg[5]/P0001 ,
		_w1260_,
		_w6162_
	);
	LUT2 #(
		.INIT('h1)
	) name5631 (
		_w5206_,
		_w6162_,
		_w6163_
	);
	LUT2 #(
		.INIT('h8)
	) name5632 (
		_w6161_,
		_w6163_,
		_w6164_
	);
	LUT2 #(
		.INIT('h1)
	) name5633 (
		_w1196_,
		_w1225_,
		_w6165_
	);
	LUT2 #(
		.INIT('h8)
	) name5634 (
		_w5239_,
		_w6165_,
		_w6166_
	);
	LUT2 #(
		.INIT('h4)
	) name5635 (
		\sa31_reg[6]/NET0131 ,
		_w5263_,
		_w6167_
	);
	LUT2 #(
		.INIT('h4)
	) name5636 (
		\sa31_reg[3]/P0001 ,
		_w1187_,
		_w6168_
	);
	LUT2 #(
		.INIT('h2)
	) name5637 (
		\sa31_reg[2]/P0001 ,
		_w5270_,
		_w6169_
	);
	LUT2 #(
		.INIT('h4)
	) name5638 (
		_w6166_,
		_w6169_,
		_w6170_
	);
	LUT2 #(
		.INIT('h1)
	) name5639 (
		_w6167_,
		_w6168_,
		_w6171_
	);
	LUT2 #(
		.INIT('h8)
	) name5640 (
		_w6170_,
		_w6171_,
		_w6172_
	);
	LUT2 #(
		.INIT('h1)
	) name5641 (
		_w6164_,
		_w6172_,
		_w6173_
	);
	LUT2 #(
		.INIT('h1)
	) name5642 (
		\sa31_reg[1]/P0001 ,
		_w1278_,
		_w6174_
	);
	LUT2 #(
		.INIT('h4)
	) name5643 (
		_w6159_,
		_w6174_,
		_w6175_
	);
	LUT2 #(
		.INIT('h4)
	) name5644 (
		_w6173_,
		_w6175_,
		_w6176_
	);
	LUT2 #(
		.INIT('h1)
	) name5645 (
		_w6158_,
		_w6176_,
		_w6177_
	);
	LUT2 #(
		.INIT('h1)
	) name5646 (
		_w6113_,
		_w6177_,
		_w6178_
	);
	LUT2 #(
		.INIT('h4)
	) name5647 (
		_w6109_,
		_w6178_,
		_w6179_
	);
	LUT2 #(
		.INIT('h4)
	) name5648 (
		_w6144_,
		_w6179_,
		_w6180_
	);
	LUT2 #(
		.INIT('h2)
	) name5649 (
		\u0_w_reg[2][13]/P0001 ,
		_w6180_,
		_w6181_
	);
	LUT2 #(
		.INIT('h4)
	) name5650 (
		\u0_w_reg[2][13]/P0001 ,
		_w6180_,
		_w6182_
	);
	LUT2 #(
		.INIT('h1)
	) name5651 (
		_w6181_,
		_w6182_,
		_w6183_
	);
	LUT2 #(
		.INIT('h8)
	) name5652 (
		_w5307_,
		_w6183_,
		_w6184_
	);
	LUT2 #(
		.INIT('h1)
	) name5653 (
		_w5307_,
		_w6183_,
		_w6185_
	);
	LUT2 #(
		.INIT('h1)
	) name5654 (
		_w6184_,
		_w6185_,
		_w6186_
	);
	LUT2 #(
		.INIT('h1)
	) name5655 (
		_w6079_,
		_w6186_,
		_w6187_
	);
	LUT2 #(
		.INIT('h8)
	) name5656 (
		_w6079_,
		_w6186_,
		_w6188_
	);
	LUT2 #(
		.INIT('h1)
	) name5657 (
		\ld_r_reg/P0001 ,
		_w6187_,
		_w6189_
	);
	LUT2 #(
		.INIT('h4)
	) name5658 (
		_w6188_,
		_w6189_,
		_w6190_
	);
	LUT2 #(
		.INIT('h1)
	) name5659 (
		\text_in_r_reg[45]/P0001 ,
		\u0_w_reg[2][13]/P0001 ,
		_w6191_
	);
	LUT2 #(
		.INIT('h8)
	) name5660 (
		\text_in_r_reg[45]/P0001 ,
		\u0_w_reg[2][13]/P0001 ,
		_w6192_
	);
	LUT2 #(
		.INIT('h2)
	) name5661 (
		\ld_r_reg/P0001 ,
		_w6191_,
		_w6193_
	);
	LUT2 #(
		.INIT('h4)
	) name5662 (
		_w6192_,
		_w6193_,
		_w6194_
	);
	LUT2 #(
		.INIT('h1)
	) name5663 (
		_w6190_,
		_w6194_,
		_w6195_
	);
	LUT2 #(
		.INIT('h1)
	) name5664 (
		_w5194_,
		_w5931_,
		_w6196_
	);
	LUT2 #(
		.INIT('h8)
	) name5665 (
		_w5194_,
		_w5931_,
		_w6197_
	);
	LUT2 #(
		.INIT('h1)
	) name5666 (
		_w6196_,
		_w6197_,
		_w6198_
	);
	LUT2 #(
		.INIT('h2)
	) name5667 (
		\u0_w_reg[2][14]/P0001 ,
		_w1300_,
		_w6199_
	);
	LUT2 #(
		.INIT('h4)
	) name5668 (
		\u0_w_reg[2][14]/P0001 ,
		_w1300_,
		_w6200_
	);
	LUT2 #(
		.INIT('h1)
	) name5669 (
		_w6199_,
		_w6200_,
		_w6201_
	);
	LUT2 #(
		.INIT('h8)
	) name5670 (
		_w5307_,
		_w6201_,
		_w6202_
	);
	LUT2 #(
		.INIT('h1)
	) name5671 (
		_w5307_,
		_w6201_,
		_w6203_
	);
	LUT2 #(
		.INIT('h1)
	) name5672 (
		_w6202_,
		_w6203_,
		_w6204_
	);
	LUT2 #(
		.INIT('h1)
	) name5673 (
		_w6198_,
		_w6204_,
		_w6205_
	);
	LUT2 #(
		.INIT('h8)
	) name5674 (
		_w6198_,
		_w6204_,
		_w6206_
	);
	LUT2 #(
		.INIT('h1)
	) name5675 (
		\ld_r_reg/P0001 ,
		_w6205_,
		_w6207_
	);
	LUT2 #(
		.INIT('h4)
	) name5676 (
		_w6206_,
		_w6207_,
		_w6208_
	);
	LUT2 #(
		.INIT('h2)
	) name5677 (
		\text_in_r_reg[46]/P0001 ,
		\u0_w_reg[2][14]/P0001 ,
		_w6209_
	);
	LUT2 #(
		.INIT('h4)
	) name5678 (
		\text_in_r_reg[46]/P0001 ,
		\u0_w_reg[2][14]/P0001 ,
		_w6210_
	);
	LUT2 #(
		.INIT('h2)
	) name5679 (
		\ld_r_reg/P0001 ,
		_w6209_,
		_w6211_
	);
	LUT2 #(
		.INIT('h4)
	) name5680 (
		_w6210_,
		_w6211_,
		_w6212_
	);
	LUT2 #(
		.INIT('h1)
	) name5681 (
		_w6208_,
		_w6212_,
		_w6213_
	);
	LUT2 #(
		.INIT('h1)
	) name5682 (
		_w541_,
		_w605_,
		_w6214_
	);
	LUT2 #(
		.INIT('h2)
	) name5683 (
		\sa13_reg[2]/P0001 ,
		_w6214_,
		_w6215_
	);
	LUT2 #(
		.INIT('h8)
	) name5684 (
		\sa13_reg[6]/NET0131 ,
		_w550_,
		_w6216_
	);
	LUT2 #(
		.INIT('h8)
	) name5685 (
		\sa13_reg[4]/P0001 ,
		_w6216_,
		_w6217_
	);
	LUT2 #(
		.INIT('h1)
	) name5686 (
		_w610_,
		_w617_,
		_w6218_
	);
	LUT2 #(
		.INIT('h4)
	) name5687 (
		_w6217_,
		_w6218_,
		_w6219_
	);
	LUT2 #(
		.INIT('h1)
	) name5688 (
		\sa13_reg[2]/P0001 ,
		_w6219_,
		_w6220_
	);
	LUT2 #(
		.INIT('h4)
	) name5689 (
		_w854_,
		_w904_,
		_w6221_
	);
	LUT2 #(
		.INIT('h4)
	) name5690 (
		_w6215_,
		_w6221_,
		_w6222_
	);
	LUT2 #(
		.INIT('h4)
	) name5691 (
		_w6220_,
		_w6222_,
		_w6223_
	);
	LUT2 #(
		.INIT('h2)
	) name5692 (
		\sa13_reg[1]/P0001 ,
		_w6223_,
		_w6224_
	);
	LUT2 #(
		.INIT('h1)
	) name5693 (
		_w536_,
		_w650_,
		_w6225_
	);
	LUT2 #(
		.INIT('h2)
	) name5694 (
		_w603_,
		_w6225_,
		_w6226_
	);
	LUT2 #(
		.INIT('h1)
	) name5695 (
		_w921_,
		_w5687_,
		_w6227_
	);
	LUT2 #(
		.INIT('h1)
	) name5696 (
		\sa13_reg[2]/P0001 ,
		_w6227_,
		_w6228_
	);
	LUT2 #(
		.INIT('h1)
	) name5697 (
		\sa13_reg[2]/P0001 ,
		_w572_,
		_w6229_
	);
	LUT2 #(
		.INIT('h4)
	) name5698 (
		_w665_,
		_w6229_,
		_w6230_
	);
	LUT2 #(
		.INIT('h2)
	) name5699 (
		\sa13_reg[2]/P0001 ,
		_w5671_,
		_w6231_
	);
	LUT2 #(
		.INIT('h4)
	) name5700 (
		_w862_,
		_w6231_,
		_w6232_
	);
	LUT2 #(
		.INIT('h1)
	) name5701 (
		_w6230_,
		_w6232_,
		_w6233_
	);
	LUT2 #(
		.INIT('h1)
	) name5702 (
		_w649_,
		_w5687_,
		_w6234_
	);
	LUT2 #(
		.INIT('h4)
	) name5703 (
		_w6233_,
		_w6234_,
		_w6235_
	);
	LUT2 #(
		.INIT('h1)
	) name5704 (
		\sa13_reg[1]/P0001 ,
		_w6235_,
		_w6236_
	);
	LUT2 #(
		.INIT('h1)
	) name5705 (
		_w654_,
		_w953_,
		_w6237_
	);
	LUT2 #(
		.INIT('h4)
	) name5706 (
		_w6226_,
		_w6237_,
		_w6238_
	);
	LUT2 #(
		.INIT('h4)
	) name5707 (
		_w6228_,
		_w6238_,
		_w6239_
	);
	LUT2 #(
		.INIT('h4)
	) name5708 (
		_w6224_,
		_w6239_,
		_w6240_
	);
	LUT2 #(
		.INIT('h4)
	) name5709 (
		_w6236_,
		_w6240_,
		_w6241_
	);
	LUT2 #(
		.INIT('h1)
	) name5710 (
		\sa13_reg[0]/P0001 ,
		_w6241_,
		_w6242_
	);
	LUT2 #(
		.INIT('h8)
	) name5711 (
		_w540_,
		_w555_,
		_w6243_
	);
	LUT2 #(
		.INIT('h1)
	) name5712 (
		_w571_,
		_w6243_,
		_w6244_
	);
	LUT2 #(
		.INIT('h8)
	) name5713 (
		\sa13_reg[4]/P0001 ,
		_w912_,
		_w6245_
	);
	LUT2 #(
		.INIT('h4)
	) name5714 (
		\sa13_reg[5]/P0001 ,
		_w5458_,
		_w6246_
	);
	LUT2 #(
		.INIT('h1)
	) name5715 (
		_w5650_,
		_w6245_,
		_w6247_
	);
	LUT2 #(
		.INIT('h4)
	) name5716 (
		_w6246_,
		_w6247_,
		_w6248_
	);
	LUT2 #(
		.INIT('h2)
	) name5717 (
		\sa13_reg[2]/P0001 ,
		_w6248_,
		_w6249_
	);
	LUT2 #(
		.INIT('h2)
	) name5718 (
		_w6244_,
		_w6249_,
		_w6250_
	);
	LUT2 #(
		.INIT('h2)
	) name5719 (
		\sa13_reg[1]/P0001 ,
		_w6250_,
		_w6251_
	);
	LUT2 #(
		.INIT('h4)
	) name5720 (
		\sa13_reg[3]/P0001 ,
		_w5458_,
		_w6252_
	);
	LUT2 #(
		.INIT('h8)
	) name5721 (
		_w532_,
		_w6252_,
		_w6253_
	);
	LUT2 #(
		.INIT('h1)
	) name5722 (
		_w608_,
		_w928_,
		_w6254_
	);
	LUT2 #(
		.INIT('h1)
	) name5723 (
		\sa13_reg[7]/NET0131 ,
		_w6254_,
		_w6255_
	);
	LUT2 #(
		.INIT('h4)
	) name5724 (
		_w670_,
		_w864_,
		_w6256_
	);
	LUT2 #(
		.INIT('h1)
	) name5725 (
		_w6253_,
		_w6256_,
		_w6257_
	);
	LUT2 #(
		.INIT('h4)
	) name5726 (
		_w6255_,
		_w6257_,
		_w6258_
	);
	LUT2 #(
		.INIT('h1)
	) name5727 (
		\sa13_reg[1]/P0001 ,
		_w6258_,
		_w6259_
	);
	LUT2 #(
		.INIT('h1)
	) name5728 (
		_w862_,
		_w908_,
		_w6260_
	);
	LUT2 #(
		.INIT('h1)
	) name5729 (
		_w5466_,
		_w5476_,
		_w6261_
	);
	LUT2 #(
		.INIT('h8)
	) name5730 (
		_w6260_,
		_w6261_,
		_w6262_
	);
	LUT2 #(
		.INIT('h1)
	) name5731 (
		\sa13_reg[2]/P0001 ,
		_w6262_,
		_w6263_
	);
	LUT2 #(
		.INIT('h8)
	) name5732 (
		\sa13_reg[2]/P0001 ,
		_w855_,
		_w6264_
	);
	LUT2 #(
		.INIT('h1)
	) name5733 (
		_w913_,
		_w5466_,
		_w6265_
	);
	LUT2 #(
		.INIT('h4)
	) name5734 (
		_w6264_,
		_w6265_,
		_w6266_
	);
	LUT2 #(
		.INIT('h1)
	) name5735 (
		\sa13_reg[3]/P0001 ,
		_w6266_,
		_w6267_
	);
	LUT2 #(
		.INIT('h1)
	) name5736 (
		_w6259_,
		_w6263_,
		_w6268_
	);
	LUT2 #(
		.INIT('h4)
	) name5737 (
		_w6267_,
		_w6268_,
		_w6269_
	);
	LUT2 #(
		.INIT('h4)
	) name5738 (
		_w6251_,
		_w6269_,
		_w6270_
	);
	LUT2 #(
		.INIT('h2)
	) name5739 (
		\sa13_reg[0]/P0001 ,
		_w6270_,
		_w6271_
	);
	LUT2 #(
		.INIT('h4)
	) name5740 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[2]/P0001 ,
		_w6272_
	);
	LUT2 #(
		.INIT('h4)
	) name5741 (
		\sa13_reg[5]/P0001 ,
		_w617_,
		_w6273_
	);
	LUT2 #(
		.INIT('h1)
	) name5742 (
		_w654_,
		_w6273_,
		_w6274_
	);
	LUT2 #(
		.INIT('h4)
	) name5743 (
		_w542_,
		_w6274_,
		_w6275_
	);
	LUT2 #(
		.INIT('h2)
	) name5744 (
		_w6272_,
		_w6275_,
		_w6276_
	);
	LUT2 #(
		.INIT('h4)
	) name5745 (
		_w587_,
		_w920_,
		_w6277_
	);
	LUT2 #(
		.INIT('h1)
	) name5746 (
		_w537_,
		_w548_,
		_w6278_
	);
	LUT2 #(
		.INIT('h4)
	) name5747 (
		_w6277_,
		_w6278_,
		_w6279_
	);
	LUT2 #(
		.INIT('h2)
	) name5748 (
		_w680_,
		_w6279_,
		_w6280_
	);
	LUT2 #(
		.INIT('h8)
	) name5749 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w6281_
	);
	LUT2 #(
		.INIT('h8)
	) name5750 (
		_w551_,
		_w6281_,
		_w6282_
	);
	LUT2 #(
		.INIT('h8)
	) name5751 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w6283_
	);
	LUT2 #(
		.INIT('h8)
	) name5752 (
		_w547_,
		_w611_,
		_w6284_
	);
	LUT2 #(
		.INIT('h8)
	) name5753 (
		_w6283_,
		_w6284_,
		_w6285_
	);
	LUT2 #(
		.INIT('h8)
	) name5754 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[2]/P0001 ,
		_w6286_
	);
	LUT2 #(
		.INIT('h1)
	) name5755 (
		_w571_,
		_w5505_,
		_w6287_
	);
	LUT2 #(
		.INIT('h2)
	) name5756 (
		\sa13_reg[3]/P0001 ,
		_w6287_,
		_w6288_
	);
	LUT2 #(
		.INIT('h1)
	) name5757 (
		_w622_,
		_w6288_,
		_w6289_
	);
	LUT2 #(
		.INIT('h2)
	) name5758 (
		_w6286_,
		_w6289_,
		_w6290_
	);
	LUT2 #(
		.INIT('h1)
	) name5759 (
		_w561_,
		_w648_,
		_w6291_
	);
	LUT2 #(
		.INIT('h4)
	) name5760 (
		_w918_,
		_w6291_,
		_w6292_
	);
	LUT2 #(
		.INIT('h1)
	) name5761 (
		\sa13_reg[2]/P0001 ,
		_w6292_,
		_w6293_
	);
	LUT2 #(
		.INIT('h1)
	) name5762 (
		_w558_,
		_w5682_,
		_w6294_
	);
	LUT2 #(
		.INIT('h4)
	) name5763 (
		_w6293_,
		_w6294_,
		_w6295_
	);
	LUT2 #(
		.INIT('h1)
	) name5764 (
		\sa13_reg[1]/P0001 ,
		_w6295_,
		_w6296_
	);
	LUT2 #(
		.INIT('h1)
	) name5765 (
		_w6282_,
		_w6285_,
		_w6297_
	);
	LUT2 #(
		.INIT('h4)
	) name5766 (
		_w5465_,
		_w6297_,
		_w6298_
	);
	LUT2 #(
		.INIT('h4)
	) name5767 (
		_w6280_,
		_w6298_,
		_w6299_
	);
	LUT2 #(
		.INIT('h4)
	) name5768 (
		_w6276_,
		_w6299_,
		_w6300_
	);
	LUT2 #(
		.INIT('h4)
	) name5769 (
		_w6290_,
		_w6300_,
		_w6301_
	);
	LUT2 #(
		.INIT('h4)
	) name5770 (
		_w6296_,
		_w6301_,
		_w6302_
	);
	LUT2 #(
		.INIT('h4)
	) name5771 (
		_w6271_,
		_w6302_,
		_w6303_
	);
	LUT2 #(
		.INIT('h4)
	) name5772 (
		_w6242_,
		_w6303_,
		_w6304_
	);
	LUT2 #(
		.INIT('h8)
	) name5773 (
		_w1035_,
		_w5082_,
		_w6305_
	);
	LUT2 #(
		.INIT('h1)
	) name5774 (
		_w5084_,
		_w5163_,
		_w6306_
	);
	LUT2 #(
		.INIT('h1)
	) name5775 (
		\sa02_reg[2]/P0001 ,
		_w6306_,
		_w6307_
	);
	LUT2 #(
		.INIT('h1)
	) name5776 (
		\sa02_reg[1]/P0001 ,
		_w5805_,
		_w6308_
	);
	LUT2 #(
		.INIT('h4)
	) name5777 (
		_w6305_,
		_w6308_,
		_w6309_
	);
	LUT2 #(
		.INIT('h4)
	) name5778 (
		_w6307_,
		_w6309_,
		_w6310_
	);
	LUT2 #(
		.INIT('h8)
	) name5779 (
		_w1011_,
		_w1038_,
		_w6311_
	);
	LUT2 #(
		.INIT('h4)
	) name5780 (
		\sa02_reg[3]/P0001 ,
		_w1023_,
		_w6312_
	);
	LUT2 #(
		.INIT('h1)
	) name5781 (
		_w983_,
		_w6311_,
		_w6313_
	);
	LUT2 #(
		.INIT('h4)
	) name5782 (
		_w6312_,
		_w6313_,
		_w6314_
	);
	LUT2 #(
		.INIT('h1)
	) name5783 (
		\sa02_reg[2]/P0001 ,
		_w6314_,
		_w6315_
	);
	LUT2 #(
		.INIT('h2)
	) name5784 (
		\sa02_reg[1]/P0001 ,
		_w1037_,
		_w6316_
	);
	LUT2 #(
		.INIT('h8)
	) name5785 (
		_w1083_,
		_w6316_,
		_w6317_
	);
	LUT2 #(
		.INIT('h4)
	) name5786 (
		_w6315_,
		_w6317_,
		_w6318_
	);
	LUT2 #(
		.INIT('h1)
	) name5787 (
		_w6310_,
		_w6318_,
		_w6319_
	);
	LUT2 #(
		.INIT('h8)
	) name5788 (
		\sa02_reg[2]/P0001 ,
		_w1058_,
		_w6320_
	);
	LUT2 #(
		.INIT('h1)
	) name5789 (
		_w5738_,
		_w5792_,
		_w6321_
	);
	LUT2 #(
		.INIT('h2)
	) name5790 (
		_w5106_,
		_w6321_,
		_w6322_
	);
	LUT2 #(
		.INIT('h1)
	) name5791 (
		_w1063_,
		_w5805_,
		_w6323_
	);
	LUT2 #(
		.INIT('h1)
	) name5792 (
		\sa02_reg[2]/P0001 ,
		_w6323_,
		_w6324_
	);
	LUT2 #(
		.INIT('h4)
	) name5793 (
		\sa02_reg[3]/P0001 ,
		_w976_,
		_w6325_
	);
	LUT2 #(
		.INIT('h1)
	) name5794 (
		_w994_,
		_w6325_,
		_w6326_
	);
	LUT2 #(
		.INIT('h2)
	) name5795 (
		_w5154_,
		_w6326_,
		_w6327_
	);
	LUT2 #(
		.INIT('h1)
	) name5796 (
		_w980_,
		_w1015_,
		_w6328_
	);
	LUT2 #(
		.INIT('h2)
	) name5797 (
		_w978_,
		_w6328_,
		_w6329_
	);
	LUT2 #(
		.INIT('h1)
	) name5798 (
		_w1121_,
		_w6320_,
		_w6330_
	);
	LUT2 #(
		.INIT('h4)
	) name5799 (
		_w6329_,
		_w6330_,
		_w6331_
	);
	LUT2 #(
		.INIT('h1)
	) name5800 (
		_w6322_,
		_w6324_,
		_w6332_
	);
	LUT2 #(
		.INIT('h4)
	) name5801 (
		_w6327_,
		_w6332_,
		_w6333_
	);
	LUT2 #(
		.INIT('h8)
	) name5802 (
		_w6331_,
		_w6333_,
		_w6334_
	);
	LUT2 #(
		.INIT('h4)
	) name5803 (
		_w6319_,
		_w6334_,
		_w6335_
	);
	LUT2 #(
		.INIT('h1)
	) name5804 (
		\sa02_reg[0]/P0001 ,
		_w6335_,
		_w6336_
	);
	LUT2 #(
		.INIT('h8)
	) name5805 (
		_w976_,
		_w1038_,
		_w6337_
	);
	LUT2 #(
		.INIT('h1)
	) name5806 (
		_w1005_,
		_w6337_,
		_w6338_
	);
	LUT2 #(
		.INIT('h1)
	) name5807 (
		\sa02_reg[5]/P0001 ,
		_w1015_,
		_w6339_
	);
	LUT2 #(
		.INIT('h4)
	) name5808 (
		_w5159_,
		_w6339_,
		_w6340_
	);
	LUT2 #(
		.INIT('h8)
	) name5809 (
		\sa02_reg[7]/NET0131 ,
		_w1068_,
		_w6341_
	);
	LUT2 #(
		.INIT('h1)
	) name5810 (
		_w6340_,
		_w6341_,
		_w6342_
	);
	LUT2 #(
		.INIT('h2)
	) name5811 (
		\sa02_reg[2]/P0001 ,
		_w6342_,
		_w6343_
	);
	LUT2 #(
		.INIT('h2)
	) name5812 (
		_w6338_,
		_w6343_,
		_w6344_
	);
	LUT2 #(
		.INIT('h2)
	) name5813 (
		\sa02_reg[1]/P0001 ,
		_w6344_,
		_w6345_
	);
	LUT2 #(
		.INIT('h2)
	) name5814 (
		_w1020_,
		_w5777_,
		_w6346_
	);
	LUT2 #(
		.INIT('h1)
	) name5815 (
		_w5363_,
		_w6346_,
		_w6347_
	);
	LUT2 #(
		.INIT('h1)
	) name5816 (
		\sa02_reg[3]/P0001 ,
		_w6347_,
		_w6348_
	);
	LUT2 #(
		.INIT('h1)
	) name5817 (
		_w1072_,
		_w5363_,
		_w6349_
	);
	LUT2 #(
		.INIT('h4)
	) name5818 (
		_w5156_,
		_w6349_,
		_w6350_
	);
	LUT2 #(
		.INIT('h4)
	) name5819 (
		_w5738_,
		_w6350_,
		_w6351_
	);
	LUT2 #(
		.INIT('h1)
	) name5820 (
		\sa02_reg[2]/P0001 ,
		_w6351_,
		_w6352_
	);
	LUT2 #(
		.INIT('h8)
	) name5821 (
		_w999_,
		_w1122_,
		_w6353_
	);
	LUT2 #(
		.INIT('h2)
	) name5822 (
		_w1024_,
		_w5168_,
		_w6354_
	);
	LUT2 #(
		.INIT('h1)
	) name5823 (
		_w1057_,
		_w1072_,
		_w6355_
	);
	LUT2 #(
		.INIT('h4)
	) name5824 (
		_w6353_,
		_w6355_,
		_w6356_
	);
	LUT2 #(
		.INIT('h4)
	) name5825 (
		_w6354_,
		_w6356_,
		_w6357_
	);
	LUT2 #(
		.INIT('h1)
	) name5826 (
		\sa02_reg[1]/P0001 ,
		_w6357_,
		_w6358_
	);
	LUT2 #(
		.INIT('h1)
	) name5827 (
		_w6348_,
		_w6352_,
		_w6359_
	);
	LUT2 #(
		.INIT('h4)
	) name5828 (
		_w6358_,
		_w6359_,
		_w6360_
	);
	LUT2 #(
		.INIT('h4)
	) name5829 (
		_w6345_,
		_w6360_,
		_w6361_
	);
	LUT2 #(
		.INIT('h2)
	) name5830 (
		\sa02_reg[0]/P0001 ,
		_w6361_,
		_w6362_
	);
	LUT2 #(
		.INIT('h1)
	) name5831 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		_w6363_
	);
	LUT2 #(
		.INIT('h8)
	) name5832 (
		_w1025_,
		_w1035_,
		_w6364_
	);
	LUT2 #(
		.INIT('h1)
	) name5833 (
		_w5102_,
		_w6364_,
		_w6365_
	);
	LUT2 #(
		.INIT('h4)
	) name5834 (
		_w1061_,
		_w6365_,
		_w6366_
	);
	LUT2 #(
		.INIT('h2)
	) name5835 (
		_w6363_,
		_w6366_,
		_w6367_
	);
	LUT2 #(
		.INIT('h4)
	) name5836 (
		_w1000_,
		_w1062_,
		_w6368_
	);
	LUT2 #(
		.INIT('h1)
	) name5837 (
		_w5081_,
		_w5099_,
		_w6369_
	);
	LUT2 #(
		.INIT('h4)
	) name5838 (
		_w1037_,
		_w6369_,
		_w6370_
	);
	LUT2 #(
		.INIT('h4)
	) name5839 (
		_w6368_,
		_w6370_,
		_w6371_
	);
	LUT2 #(
		.INIT('h2)
	) name5840 (
		_w5179_,
		_w6371_,
		_w6372_
	);
	LUT2 #(
		.INIT('h2)
	) name5841 (
		_w1020_,
		_w5800_,
		_w6373_
	);
	LUT2 #(
		.INIT('h8)
	) name5842 (
		\sa02_reg[3]/P0001 ,
		_w5744_,
		_w6374_
	);
	LUT2 #(
		.INIT('h1)
	) name5843 (
		_w6373_,
		_w6374_,
		_w6375_
	);
	LUT2 #(
		.INIT('h2)
	) name5844 (
		\sa02_reg[1]/P0001 ,
		_w6375_,
		_w6376_
	);
	LUT2 #(
		.INIT('h8)
	) name5845 (
		_w1038_,
		_w1094_,
		_w6377_
	);
	LUT2 #(
		.INIT('h1)
	) name5846 (
		_w1117_,
		_w6377_,
		_w6378_
	);
	LUT2 #(
		.INIT('h4)
	) name5847 (
		_w6376_,
		_w6378_,
		_w6379_
	);
	LUT2 #(
		.INIT('h2)
	) name5848 (
		\sa02_reg[2]/P0001 ,
		_w6379_,
		_w6380_
	);
	LUT2 #(
		.INIT('h4)
	) name5849 (
		\sa02_reg[3]/P0001 ,
		_w1094_,
		_w6381_
	);
	LUT2 #(
		.INIT('h1)
	) name5850 (
		_w1071_,
		_w1121_,
		_w6382_
	);
	LUT2 #(
		.INIT('h4)
	) name5851 (
		_w6381_,
		_w6382_,
		_w6383_
	);
	LUT2 #(
		.INIT('h2)
	) name5852 (
		\sa02_reg[2]/P0001 ,
		_w6383_,
		_w6384_
	);
	LUT2 #(
		.INIT('h1)
	) name5853 (
		_w1058_,
		_w6377_,
		_w6385_
	);
	LUT2 #(
		.INIT('h4)
	) name5854 (
		_w6384_,
		_w6385_,
		_w6386_
	);
	LUT2 #(
		.INIT('h1)
	) name5855 (
		\sa02_reg[1]/P0001 ,
		_w6386_,
		_w6387_
	);
	LUT2 #(
		.INIT('h1)
	) name5856 (
		_w6367_,
		_w6372_,
		_w6388_
	);
	LUT2 #(
		.INIT('h4)
	) name5857 (
		_w6380_,
		_w6388_,
		_w6389_
	);
	LUT2 #(
		.INIT('h4)
	) name5858 (
		_w6387_,
		_w6389_,
		_w6390_
	);
	LUT2 #(
		.INIT('h4)
	) name5859 (
		_w6336_,
		_w6390_,
		_w6391_
	);
	LUT2 #(
		.INIT('h4)
	) name5860 (
		_w6362_,
		_w6391_,
		_w6392_
	);
	LUT2 #(
		.INIT('h1)
	) name5861 (
		_w6304_,
		_w6392_,
		_w6393_
	);
	LUT2 #(
		.INIT('h8)
	) name5862 (
		_w6304_,
		_w6392_,
		_w6394_
	);
	LUT2 #(
		.INIT('h1)
	) name5863 (
		_w6393_,
		_w6394_,
		_w6395_
	);
	LUT2 #(
		.INIT('h8)
	) name5864 (
		_w1003_,
		_w5108_,
		_w6396_
	);
	LUT2 #(
		.INIT('h8)
	) name5865 (
		_w5159_,
		_w6396_,
		_w6397_
	);
	LUT2 #(
		.INIT('h2)
	) name5866 (
		_w1059_,
		_w5367_,
		_w6398_
	);
	LUT2 #(
		.INIT('h4)
	) name5867 (
		\sa02_reg[5]/P0001 ,
		_w5155_,
		_w6399_
	);
	LUT2 #(
		.INIT('h1)
	) name5868 (
		_w1031_,
		_w1076_,
		_w6400_
	);
	LUT2 #(
		.INIT('h4)
	) name5869 (
		_w6399_,
		_w6400_,
		_w6401_
	);
	LUT2 #(
		.INIT('h2)
	) name5870 (
		\sa02_reg[2]/P0001 ,
		_w6401_,
		_w6402_
	);
	LUT2 #(
		.INIT('h1)
	) name5871 (
		_w5809_,
		_w6397_,
		_w6403_
	);
	LUT2 #(
		.INIT('h4)
	) name5872 (
		_w6398_,
		_w6403_,
		_w6404_
	);
	LUT2 #(
		.INIT('h4)
	) name5873 (
		_w6402_,
		_w6404_,
		_w6405_
	);
	LUT2 #(
		.INIT('h2)
	) name5874 (
		\sa02_reg[0]/P0001 ,
		_w6405_,
		_w6406_
	);
	LUT2 #(
		.INIT('h1)
	) name5875 (
		_w975_,
		_w1094_,
		_w6407_
	);
	LUT2 #(
		.INIT('h2)
	) name5876 (
		_w974_,
		_w6407_,
		_w6408_
	);
	LUT2 #(
		.INIT('h2)
	) name5877 (
		_w1107_,
		_w6408_,
		_w6409_
	);
	LUT2 #(
		.INIT('h1)
	) name5878 (
		_w1130_,
		_w5082_,
		_w6410_
	);
	LUT2 #(
		.INIT('h4)
	) name5879 (
		_w5394_,
		_w6410_,
		_w6411_
	);
	LUT2 #(
		.INIT('h1)
	) name5880 (
		\sa02_reg[3]/P0001 ,
		_w6411_,
		_w6412_
	);
	LUT2 #(
		.INIT('h1)
	) name5881 (
		\sa02_reg[2]/P0001 ,
		_w1070_,
		_w6413_
	);
	LUT2 #(
		.INIT('h4)
	) name5882 (
		_w6412_,
		_w6413_,
		_w6414_
	);
	LUT2 #(
		.INIT('h1)
	) name5883 (
		_w6409_,
		_w6414_,
		_w6415_
	);
	LUT2 #(
		.INIT('h1)
	) name5884 (
		_w6406_,
		_w6415_,
		_w6416_
	);
	LUT2 #(
		.INIT('h1)
	) name5885 (
		\sa02_reg[1]/P0001 ,
		_w6416_,
		_w6417_
	);
	LUT2 #(
		.INIT('h8)
	) name5886 (
		\sa02_reg[6]/NET0131 ,
		_w1030_,
		_w6418_
	);
	LUT2 #(
		.INIT('h1)
	) name5887 (
		_w1063_,
		_w6418_,
		_w6419_
	);
	LUT2 #(
		.INIT('h4)
	) name5888 (
		_w5148_,
		_w6419_,
		_w6420_
	);
	LUT2 #(
		.INIT('h1)
	) name5889 (
		\sa02_reg[2]/P0001 ,
		_w6420_,
		_w6421_
	);
	LUT2 #(
		.INIT('h8)
	) name5890 (
		\sa02_reg[4]/P0001 ,
		_w6341_,
		_w6422_
	);
	LUT2 #(
		.INIT('h2)
	) name5891 (
		_w979_,
		_w1038_,
		_w6423_
	);
	LUT2 #(
		.INIT('h8)
	) name5892 (
		_w1068_,
		_w5753_,
		_w6424_
	);
	LUT2 #(
		.INIT('h1)
	) name5893 (
		_w6396_,
		_w6423_,
		_w6425_
	);
	LUT2 #(
		.INIT('h4)
	) name5894 (
		_w6422_,
		_w6425_,
		_w6426_
	);
	LUT2 #(
		.INIT('h4)
	) name5895 (
		_w6424_,
		_w6426_,
		_w6427_
	);
	LUT2 #(
		.INIT('h2)
	) name5896 (
		\sa02_reg[1]/P0001 ,
		_w6427_,
		_w6428_
	);
	LUT2 #(
		.INIT('h1)
	) name5897 (
		\sa02_reg[3]/P0001 ,
		_w5389_,
		_w6429_
	);
	LUT2 #(
		.INIT('h1)
	) name5898 (
		_w5776_,
		_w6429_,
		_w6430_
	);
	LUT2 #(
		.INIT('h1)
	) name5899 (
		\sa02_reg[1]/P0001 ,
		_w6430_,
		_w6431_
	);
	LUT2 #(
		.INIT('h1)
	) name5900 (
		_w1011_,
		_w5091_,
		_w6432_
	);
	LUT2 #(
		.INIT('h2)
	) name5901 (
		_w1059_,
		_w6432_,
		_w6433_
	);
	LUT2 #(
		.INIT('h4)
	) name5902 (
		\sa02_reg[1]/P0001 ,
		_w993_,
		_w6434_
	);
	LUT2 #(
		.INIT('h4)
	) name5903 (
		_w1068_,
		_w6434_,
		_w6435_
	);
	LUT2 #(
		.INIT('h1)
	) name5904 (
		_w6433_,
		_w6435_,
		_w6436_
	);
	LUT2 #(
		.INIT('h2)
	) name5905 (
		\sa02_reg[2]/P0001 ,
		_w6436_,
		_w6437_
	);
	LUT2 #(
		.INIT('h1)
	) name5906 (
		_w6421_,
		_w6428_,
		_w6438_
	);
	LUT2 #(
		.INIT('h1)
	) name5907 (
		_w6431_,
		_w6437_,
		_w6439_
	);
	LUT2 #(
		.INIT('h8)
	) name5908 (
		_w6438_,
		_w6439_,
		_w6440_
	);
	LUT2 #(
		.INIT('h1)
	) name5909 (
		\sa02_reg[0]/P0001 ,
		_w6440_,
		_w6441_
	);
	LUT2 #(
		.INIT('h8)
	) name5910 (
		\sa02_reg[6]/NET0131 ,
		_w5132_,
		_w6442_
	);
	LUT2 #(
		.INIT('h8)
	) name5911 (
		_w5168_,
		_w5738_,
		_w6443_
	);
	LUT2 #(
		.INIT('h8)
	) name5912 (
		_w994_,
		_w5108_,
		_w6444_
	);
	LUT2 #(
		.INIT('h1)
	) name5913 (
		_w1110_,
		_w5098_,
		_w6445_
	);
	LUT2 #(
		.INIT('h1)
	) name5914 (
		_w5181_,
		_w6444_,
		_w6446_
	);
	LUT2 #(
		.INIT('h8)
	) name5915 (
		_w6445_,
		_w6446_,
		_w6447_
	);
	LUT2 #(
		.INIT('h4)
	) name5916 (
		_w1014_,
		_w6447_,
		_w6448_
	);
	LUT2 #(
		.INIT('h2)
	) name5917 (
		\sa02_reg[1]/P0001 ,
		_w6448_,
		_w6449_
	);
	LUT2 #(
		.INIT('h1)
	) name5918 (
		_w1063_,
		_w5750_,
		_w6450_
	);
	LUT2 #(
		.INIT('h8)
	) name5919 (
		_w5103_,
		_w6450_,
		_w6451_
	);
	LUT2 #(
		.INIT('h2)
	) name5920 (
		\sa02_reg[2]/P0001 ,
		_w6451_,
		_w6452_
	);
	LUT2 #(
		.INIT('h8)
	) name5921 (
		\sa02_reg[5]/P0001 ,
		_w5786_,
		_w6453_
	);
	LUT2 #(
		.INIT('h1)
	) name5922 (
		_w5364_,
		_w6453_,
		_w6454_
	);
	LUT2 #(
		.INIT('h1)
	) name5923 (
		\sa02_reg[2]/P0001 ,
		_w6454_,
		_w6455_
	);
	LUT2 #(
		.INIT('h1)
	) name5924 (
		_w1011_,
		_w1015_,
		_w6456_
	);
	LUT2 #(
		.INIT('h2)
	) name5925 (
		_w1095_,
		_w6456_,
		_w6457_
	);
	LUT2 #(
		.INIT('h1)
	) name5926 (
		_w975_,
		_w980_,
		_w6458_
	);
	LUT2 #(
		.INIT('h1)
	) name5927 (
		\sa02_reg[2]/P0001 ,
		_w6458_,
		_w6459_
	);
	LUT2 #(
		.INIT('h1)
	) name5928 (
		_w5163_,
		_w6459_,
		_w6460_
	);
	LUT2 #(
		.INIT('h2)
	) name5929 (
		\sa02_reg[1]/P0001 ,
		_w6460_,
		_w6461_
	);
	LUT2 #(
		.INIT('h1)
	) name5930 (
		_w5738_,
		_w5818_,
		_w6462_
	);
	LUT2 #(
		.INIT('h4)
	) name5931 (
		_w6457_,
		_w6462_,
		_w6463_
	);
	LUT2 #(
		.INIT('h4)
	) name5932 (
		_w6455_,
		_w6463_,
		_w6464_
	);
	LUT2 #(
		.INIT('h4)
	) name5933 (
		_w6452_,
		_w6464_,
		_w6465_
	);
	LUT2 #(
		.INIT('h4)
	) name5934 (
		_w6461_,
		_w6465_,
		_w6466_
	);
	LUT2 #(
		.INIT('h2)
	) name5935 (
		\sa02_reg[0]/P0001 ,
		_w6466_,
		_w6467_
	);
	LUT2 #(
		.INIT('h1)
	) name5936 (
		_w6442_,
		_w6443_,
		_w6468_
	);
	LUT2 #(
		.INIT('h4)
	) name5937 (
		_w6449_,
		_w6468_,
		_w6469_
	);
	LUT2 #(
		.INIT('h4)
	) name5938 (
		_w6417_,
		_w6469_,
		_w6470_
	);
	LUT2 #(
		.INIT('h1)
	) name5939 (
		_w6441_,
		_w6467_,
		_w6471_
	);
	LUT2 #(
		.INIT('h8)
	) name5940 (
		_w6470_,
		_w6471_,
		_w6472_
	);
	LUT2 #(
		.INIT('h1)
	) name5941 (
		_w5417_,
		_w6472_,
		_w6473_
	);
	LUT2 #(
		.INIT('h8)
	) name5942 (
		_w5417_,
		_w6472_,
		_w6474_
	);
	LUT2 #(
		.INIT('h1)
	) name5943 (
		_w6473_,
		_w6474_,
		_w6475_
	);
	LUT2 #(
		.INIT('h2)
	) name5944 (
		_w6395_,
		_w6475_,
		_w6476_
	);
	LUT2 #(
		.INIT('h4)
	) name5945 (
		_w6395_,
		_w6475_,
		_w6477_
	);
	LUT2 #(
		.INIT('h1)
	) name5946 (
		_w6476_,
		_w6477_,
		_w6478_
	);
	LUT2 #(
		.INIT('h1)
	) name5947 (
		_w1193_,
		_w1219_,
		_w6479_
	);
	LUT2 #(
		.INIT('h1)
	) name5948 (
		\sa31_reg[2]/P0001 ,
		_w6479_,
		_w6480_
	);
	LUT2 #(
		.INIT('h1)
	) name5949 (
		_w1239_,
		_w6480_,
		_w6481_
	);
	LUT2 #(
		.INIT('h2)
	) name5950 (
		\sa31_reg[1]/P0001 ,
		_w6481_,
		_w6482_
	);
	LUT2 #(
		.INIT('h8)
	) name5951 (
		\sa31_reg[3]/P0001 ,
		_w1151_,
		_w6483_
	);
	LUT2 #(
		.INIT('h4)
	) name5952 (
		\sa31_reg[4]/P0001 ,
		_w1276_,
		_w6484_
	);
	LUT2 #(
		.INIT('h1)
	) name5953 (
		_w6483_,
		_w6484_,
		_w6485_
	);
	LUT2 #(
		.INIT('h1)
	) name5954 (
		\sa31_reg[2]/P0001 ,
		_w6485_,
		_w6486_
	);
	LUT2 #(
		.INIT('h8)
	) name5955 (
		_w1158_,
		_w1196_,
		_w6487_
	);
	LUT2 #(
		.INIT('h8)
	) name5956 (
		\sa31_reg[7]/P0001 ,
		_w1277_,
		_w6488_
	);
	LUT2 #(
		.INIT('h1)
	) name5957 (
		_w6487_,
		_w6488_,
		_w6489_
	);
	LUT2 #(
		.INIT('h1)
	) name5958 (
		\sa31_reg[2]/P0001 ,
		_w6489_,
		_w6490_
	);
	LUT2 #(
		.INIT('h4)
	) name5959 (
		\sa31_reg[3]/P0001 ,
		_w1194_,
		_w6491_
	);
	LUT2 #(
		.INIT('h1)
	) name5960 (
		_w1168_,
		_w6089_,
		_w6492_
	);
	LUT2 #(
		.INIT('h8)
	) name5961 (
		_w5251_,
		_w6492_,
		_w6493_
	);
	LUT2 #(
		.INIT('h2)
	) name5962 (
		\sa31_reg[2]/P0001 ,
		_w6493_,
		_w6494_
	);
	LUT2 #(
		.INIT('h8)
	) name5963 (
		_w1162_,
		_w5239_,
		_w6495_
	);
	LUT2 #(
		.INIT('h8)
	) name5964 (
		\sa31_reg[4]/P0001 ,
		_w6495_,
		_w6496_
	);
	LUT2 #(
		.INIT('h2)
	) name5965 (
		\sa31_reg[5]/P0001 ,
		_w1146_,
		_w6497_
	);
	LUT2 #(
		.INIT('h2)
	) name5966 (
		_w1225_,
		_w6497_,
		_w6498_
	);
	LUT2 #(
		.INIT('h8)
	) name5967 (
		_w1152_,
		_w1158_,
		_w6499_
	);
	LUT2 #(
		.INIT('h1)
	) name5968 (
		_w1220_,
		_w5261_,
		_w6500_
	);
	LUT2 #(
		.INIT('h4)
	) name5969 (
		_w5209_,
		_w6500_,
		_w6501_
	);
	LUT2 #(
		.INIT('h2)
	) name5970 (
		\sa31_reg[2]/P0001 ,
		_w6501_,
		_w6502_
	);
	LUT2 #(
		.INIT('h1)
	) name5971 (
		_w6498_,
		_w6499_,
		_w6503_
	);
	LUT2 #(
		.INIT('h4)
	) name5972 (
		_w6496_,
		_w6503_,
		_w6504_
	);
	LUT2 #(
		.INIT('h4)
	) name5973 (
		_w6502_,
		_w6504_,
		_w6505_
	);
	LUT2 #(
		.INIT('h1)
	) name5974 (
		\sa31_reg[1]/P0001 ,
		_w6505_,
		_w6506_
	);
	LUT2 #(
		.INIT('h1)
	) name5975 (
		_w6145_,
		_w6491_,
		_w6507_
	);
	LUT2 #(
		.INIT('h4)
	) name5976 (
		_w6486_,
		_w6507_,
		_w6508_
	);
	LUT2 #(
		.INIT('h4)
	) name5977 (
		_w6490_,
		_w6508_,
		_w6509_
	);
	LUT2 #(
		.INIT('h4)
	) name5978 (
		_w6482_,
		_w6509_,
		_w6510_
	);
	LUT2 #(
		.INIT('h4)
	) name5979 (
		_w6494_,
		_w6510_,
		_w6511_
	);
	LUT2 #(
		.INIT('h4)
	) name5980 (
		_w6506_,
		_w6511_,
		_w6512_
	);
	LUT2 #(
		.INIT('h2)
	) name5981 (
		\sa31_reg[0]/P0002 ,
		_w6512_,
		_w6513_
	);
	LUT2 #(
		.INIT('h4)
	) name5982 (
		\sa31_reg[1]/P0001 ,
		\sa31_reg[2]/P0001 ,
		_w6514_
	);
	LUT2 #(
		.INIT('h2)
	) name5983 (
		_w1166_,
		_w5269_,
		_w6515_
	);
	LUT2 #(
		.INIT('h8)
	) name5984 (
		_w6514_,
		_w6515_,
		_w6516_
	);
	LUT2 #(
		.INIT('h1)
	) name5985 (
		_w6110_,
		_w6115_,
		_w6517_
	);
	LUT2 #(
		.INIT('h1)
	) name5986 (
		\sa31_reg[3]/P0001 ,
		_w6517_,
		_w6518_
	);
	LUT2 #(
		.INIT('h2)
	) name5987 (
		_w6133_,
		_w6518_,
		_w6519_
	);
	LUT2 #(
		.INIT('h8)
	) name5988 (
		_w1194_,
		_w1265_,
		_w6520_
	);
	LUT2 #(
		.INIT('h4)
	) name5989 (
		_w1159_,
		_w1186_,
		_w6521_
	);
	LUT2 #(
		.INIT('h8)
	) name5990 (
		_w1162_,
		_w1182_,
		_w6522_
	);
	LUT2 #(
		.INIT('h2)
	) name5991 (
		\sa31_reg[1]/P0001 ,
		_w6152_,
		_w6523_
	);
	LUT2 #(
		.INIT('h1)
	) name5992 (
		_w6521_,
		_w6522_,
		_w6524_
	);
	LUT2 #(
		.INIT('h8)
	) name5993 (
		_w6523_,
		_w6524_,
		_w6525_
	);
	LUT2 #(
		.INIT('h4)
	) name5994 (
		_w6520_,
		_w6525_,
		_w6526_
	);
	LUT2 #(
		.INIT('h1)
	) name5995 (
		_w6519_,
		_w6526_,
		_w6527_
	);
	LUT2 #(
		.INIT('h8)
	) name5996 (
		_w1166_,
		_w5269_,
		_w6528_
	);
	LUT2 #(
		.INIT('h1)
	) name5997 (
		_w5250_,
		_w6528_,
		_w6529_
	);
	LUT2 #(
		.INIT('h4)
	) name5998 (
		\sa31_reg[4]/P0001 ,
		_w1229_,
		_w6530_
	);
	LUT2 #(
		.INIT('h4)
	) name5999 (
		\sa31_reg[3]/P0001 ,
		_w6530_,
		_w6531_
	);
	LUT2 #(
		.INIT('h2)
	) name6000 (
		_w6529_,
		_w6531_,
		_w6532_
	);
	LUT2 #(
		.INIT('h1)
	) name6001 (
		\sa31_reg[2]/P0001 ,
		_w6532_,
		_w6533_
	);
	LUT2 #(
		.INIT('h1)
	) name6002 (
		_w1151_,
		_w1187_,
		_w6534_
	);
	LUT2 #(
		.INIT('h2)
	) name6003 (
		_w1248_,
		_w6534_,
		_w6535_
	);
	LUT2 #(
		.INIT('h1)
	) name6004 (
		_w6516_,
		_w6535_,
		_w6536_
	);
	LUT2 #(
		.INIT('h4)
	) name6005 (
		_w6527_,
		_w6536_,
		_w6537_
	);
	LUT2 #(
		.INIT('h4)
	) name6006 (
		_w6533_,
		_w6537_,
		_w6538_
	);
	LUT2 #(
		.INIT('h1)
	) name6007 (
		\sa31_reg[0]/P0002 ,
		_w6538_,
		_w6539_
	);
	LUT2 #(
		.INIT('h8)
	) name6008 (
		\sa31_reg[7]/P0001 ,
		_w6531_,
		_w6540_
	);
	LUT2 #(
		.INIT('h1)
	) name6009 (
		_w1247_,
		_w6540_,
		_w6541_
	);
	LUT2 #(
		.INIT('h2)
	) name6010 (
		\sa31_reg[2]/P0001 ,
		_w6541_,
		_w6542_
	);
	LUT2 #(
		.INIT('h8)
	) name6011 (
		_w1152_,
		_w1178_,
		_w6543_
	);
	LUT2 #(
		.INIT('h1)
	) name6012 (
		_w1260_,
		_w6543_,
		_w6544_
	);
	LUT2 #(
		.INIT('h1)
	) name6013 (
		\sa31_reg[7]/P0001 ,
		_w6544_,
		_w6545_
	);
	LUT2 #(
		.INIT('h4)
	) name6014 (
		\sa31_reg[3]/P0001 ,
		_w1173_,
		_w6546_
	);
	LUT2 #(
		.INIT('h1)
	) name6015 (
		_w5264_,
		_w6546_,
		_w6547_
	);
	LUT2 #(
		.INIT('h4)
	) name6016 (
		_w6545_,
		_w6547_,
		_w6548_
	);
	LUT2 #(
		.INIT('h1)
	) name6017 (
		\sa31_reg[2]/P0001 ,
		_w6548_,
		_w6549_
	);
	LUT2 #(
		.INIT('h1)
	) name6018 (
		_w5295_,
		_w6542_,
		_w6550_
	);
	LUT2 #(
		.INIT('h4)
	) name6019 (
		_w6549_,
		_w6550_,
		_w6551_
	);
	LUT2 #(
		.INIT('h1)
	) name6020 (
		\sa31_reg[1]/P0001 ,
		_w6551_,
		_w6552_
	);
	LUT2 #(
		.INIT('h8)
	) name6021 (
		\sa31_reg[2]/P0001 ,
		_w6162_,
		_w6553_
	);
	LUT2 #(
		.INIT('h1)
	) name6022 (
		_w6167_,
		_w6553_,
		_w6554_
	);
	LUT2 #(
		.INIT('h1)
	) name6023 (
		\sa31_reg[7]/P0001 ,
		_w6554_,
		_w6555_
	);
	LUT2 #(
		.INIT('h8)
	) name6024 (
		_w1166_,
		_w1196_,
		_w6556_
	);
	LUT2 #(
		.INIT('h1)
	) name6025 (
		\sa31_reg[2]/P0001 ,
		_w6556_,
		_w6557_
	);
	LUT2 #(
		.INIT('h1)
	) name6026 (
		_w6114_,
		_w6557_,
		_w6558_
	);
	LUT2 #(
		.INIT('h1)
	) name6027 (
		_w1231_,
		_w6558_,
		_w6559_
	);
	LUT2 #(
		.INIT('h4)
	) name6028 (
		_w6555_,
		_w6559_,
		_w6560_
	);
	LUT2 #(
		.INIT('h2)
	) name6029 (
		\sa31_reg[1]/P0001 ,
		_w6560_,
		_w6561_
	);
	LUT2 #(
		.INIT('h8)
	) name6030 (
		\sa31_reg[6]/NET0131 ,
		_w1222_,
		_w6562_
	);
	LUT2 #(
		.INIT('h8)
	) name6031 (
		_w1152_,
		_w6087_,
		_w6563_
	);
	LUT2 #(
		.INIT('h1)
	) name6032 (
		_w6562_,
		_w6563_,
		_w6564_
	);
	LUT2 #(
		.INIT('h4)
	) name6033 (
		_w6561_,
		_w6564_,
		_w6565_
	);
	LUT2 #(
		.INIT('h4)
	) name6034 (
		_w6539_,
		_w6565_,
		_w6566_
	);
	LUT2 #(
		.INIT('h4)
	) name6035 (
		_w6552_,
		_w6566_,
		_w6567_
	);
	LUT2 #(
		.INIT('h4)
	) name6036 (
		_w6513_,
		_w6567_,
		_w6568_
	);
	LUT2 #(
		.INIT('h4)
	) name6037 (
		\sa31_reg[3]/P0001 ,
		_w1149_,
		_w6569_
	);
	LUT2 #(
		.INIT('h4)
	) name6038 (
		_w1244_,
		_w6569_,
		_w6570_
	);
	LUT2 #(
		.INIT('h4)
	) name6039 (
		\sa31_reg[4]/P0001 ,
		_w1182_,
		_w6571_
	);
	LUT2 #(
		.INIT('h8)
	) name6040 (
		_w1279_,
		_w6571_,
		_w6572_
	);
	LUT2 #(
		.INIT('h2)
	) name6041 (
		\sa31_reg[4]/P0001 ,
		_w1178_,
		_w6573_
	);
	LUT2 #(
		.INIT('h4)
	) name6042 (
		_w5205_,
		_w6573_,
		_w6574_
	);
	LUT2 #(
		.INIT('h1)
	) name6043 (
		_w1194_,
		_w6574_,
		_w6575_
	);
	LUT2 #(
		.INIT('h1)
	) name6044 (
		\sa31_reg[2]/P0001 ,
		_w6575_,
		_w6576_
	);
	LUT2 #(
		.INIT('h1)
	) name6045 (
		_w6167_,
		_w6570_,
		_w6577_
	);
	LUT2 #(
		.INIT('h4)
	) name6046 (
		_w6572_,
		_w6577_,
		_w6578_
	);
	LUT2 #(
		.INIT('h4)
	) name6047 (
		_w6576_,
		_w6578_,
		_w6579_
	);
	LUT2 #(
		.INIT('h2)
	) name6048 (
		\sa31_reg[0]/P0002 ,
		_w6579_,
		_w6580_
	);
	LUT2 #(
		.INIT('h4)
	) name6049 (
		\sa31_reg[3]/P0001 ,
		_w1201_,
		_w6581_
	);
	LUT2 #(
		.INIT('h1)
	) name6050 (
		_w6499_,
		_w6581_,
		_w6582_
	);
	LUT2 #(
		.INIT('h1)
	) name6051 (
		\sa31_reg[2]/P0001 ,
		_w6582_,
		_w6583_
	);
	LUT2 #(
		.INIT('h8)
	) name6052 (
		_w5238_,
		_w6571_,
		_w6584_
	);
	LUT2 #(
		.INIT('h1)
	) name6053 (
		_w6556_,
		_w6584_,
		_w6585_
	);
	LUT2 #(
		.INIT('h4)
	) name6054 (
		_w6583_,
		_w6585_,
		_w6586_
	);
	LUT2 #(
		.INIT('h4)
	) name6055 (
		_w6580_,
		_w6586_,
		_w6587_
	);
	LUT2 #(
		.INIT('h1)
	) name6056 (
		\sa31_reg[1]/P0001 ,
		_w6587_,
		_w6588_
	);
	LUT2 #(
		.INIT('h4)
	) name6057 (
		\sa31_reg[4]/P0001 ,
		_w1256_,
		_w6589_
	);
	LUT2 #(
		.INIT('h1)
	) name6058 (
		_w5198_,
		_w6589_,
		_w6590_
	);
	LUT2 #(
		.INIT('h1)
	) name6059 (
		\sa31_reg[3]/P0001 ,
		_w6590_,
		_w6591_
	);
	LUT2 #(
		.INIT('h1)
	) name6060 (
		_w5209_,
		_w6591_,
		_w6592_
	);
	LUT2 #(
		.INIT('h2)
	) name6061 (
		\sa31_reg[2]/P0001 ,
		_w6592_,
		_w6593_
	);
	LUT2 #(
		.INIT('h1)
	) name6062 (
		_w6153_,
		_w6495_,
		_w6594_
	);
	LUT2 #(
		.INIT('h2)
	) name6063 (
		\sa31_reg[1]/P0001 ,
		_w6594_,
		_w6595_
	);
	LUT2 #(
		.INIT('h2)
	) name6064 (
		\sa31_reg[4]/P0001 ,
		_w1276_,
		_w6596_
	);
	LUT2 #(
		.INIT('h2)
	) name6065 (
		\sa31_reg[6]/NET0131 ,
		_w6596_,
		_w6597_
	);
	LUT2 #(
		.INIT('h8)
	) name6066 (
		\sa31_reg[4]/P0001 ,
		_w1229_,
		_w6598_
	);
	LUT2 #(
		.INIT('h4)
	) name6067 (
		\sa31_reg[3]/P0001 ,
		_w1186_,
		_w6599_
	);
	LUT2 #(
		.INIT('h1)
	) name6068 (
		_w6598_,
		_w6599_,
		_w6600_
	);
	LUT2 #(
		.INIT('h4)
	) name6069 (
		_w6597_,
		_w6600_,
		_w6601_
	);
	LUT2 #(
		.INIT('h2)
	) name6070 (
		_w1232_,
		_w6601_,
		_w6602_
	);
	LUT2 #(
		.INIT('h8)
	) name6071 (
		_w1151_,
		_w1248_,
		_w6603_
	);
	LUT2 #(
		.INIT('h8)
	) name6072 (
		_w1150_,
		_w1162_,
		_w6604_
	);
	LUT2 #(
		.INIT('h1)
	) name6073 (
		_w6487_,
		_w6603_,
		_w6605_
	);
	LUT2 #(
		.INIT('h4)
	) name6074 (
		_w6604_,
		_w6605_,
		_w6606_
	);
	LUT2 #(
		.INIT('h4)
	) name6075 (
		_w6595_,
		_w6606_,
		_w6607_
	);
	LUT2 #(
		.INIT('h4)
	) name6076 (
		_w6602_,
		_w6607_,
		_w6608_
	);
	LUT2 #(
		.INIT('h4)
	) name6077 (
		_w6593_,
		_w6608_,
		_w6609_
	);
	LUT2 #(
		.INIT('h2)
	) name6078 (
		\sa31_reg[0]/P0002 ,
		_w6609_,
		_w6610_
	);
	LUT2 #(
		.INIT('h1)
	) name6079 (
		_w6084_,
		_w6589_,
		_w6611_
	);
	LUT2 #(
		.INIT('h4)
	) name6080 (
		_w6124_,
		_w6611_,
		_w6612_
	);
	LUT2 #(
		.INIT('h1)
	) name6081 (
		\sa31_reg[3]/P0001 ,
		_w6612_,
		_w6613_
	);
	LUT2 #(
		.INIT('h1)
	) name6082 (
		_w1183_,
		_w5270_,
		_w6614_
	);
	LUT2 #(
		.INIT('h4)
	) name6083 (
		_w6613_,
		_w6614_,
		_w6615_
	);
	LUT2 #(
		.INIT('h2)
	) name6084 (
		_w1232_,
		_w6615_,
		_w6616_
	);
	LUT2 #(
		.INIT('h1)
	) name6085 (
		_w5207_,
		_w6080_,
		_w6617_
	);
	LUT2 #(
		.INIT('h1)
	) name6086 (
		\sa31_reg[2]/P0001 ,
		_w6617_,
		_w6618_
	);
	LUT2 #(
		.INIT('h1)
	) name6087 (
		_w1187_,
		_w5198_,
		_w6619_
	);
	LUT2 #(
		.INIT('h8)
	) name6088 (
		_w6517_,
		_w6619_,
		_w6620_
	);
	LUT2 #(
		.INIT('h8)
	) name6089 (
		\sa31_reg[1]/P0001 ,
		_w5238_,
		_w6621_
	);
	LUT2 #(
		.INIT('h4)
	) name6090 (
		_w6620_,
		_w6621_,
		_w6622_
	);
	LUT2 #(
		.INIT('h8)
	) name6091 (
		\sa31_reg[5]/P0001 ,
		_w1260_,
		_w6623_
	);
	LUT2 #(
		.INIT('h1)
	) name6092 (
		_w5204_,
		_w6153_,
		_w6624_
	);
	LUT2 #(
		.INIT('h4)
	) name6093 (
		_w6623_,
		_w6624_,
		_w6625_
	);
	LUT2 #(
		.INIT('h2)
	) name6094 (
		_w6514_,
		_w6625_,
		_w6626_
	);
	LUT2 #(
		.INIT('h8)
	) name6095 (
		\sa31_reg[4]/P0001 ,
		_w1187_,
		_w6627_
	);
	LUT2 #(
		.INIT('h1)
	) name6096 (
		_w6488_,
		_w6627_,
		_w6628_
	);
	LUT2 #(
		.INIT('h2)
	) name6097 (
		\sa31_reg[3]/P0001 ,
		_w6628_,
		_w6629_
	);
	LUT2 #(
		.INIT('h2)
	) name6098 (
		\sa31_reg[2]/P0001 ,
		_w6629_,
		_w6630_
	);
	LUT2 #(
		.INIT('h1)
	) name6099 (
		\sa31_reg[2]/P0001 ,
		_w1278_,
		_w6631_
	);
	LUT2 #(
		.INIT('h4)
	) name6100 (
		_w1233_,
		_w6582_,
		_w6632_
	);
	LUT2 #(
		.INIT('h8)
	) name6101 (
		_w6631_,
		_w6632_,
		_w6633_
	);
	LUT2 #(
		.INIT('h1)
	) name6102 (
		_w6630_,
		_w6633_,
		_w6634_
	);
	LUT2 #(
		.INIT('h2)
	) name6103 (
		\sa31_reg[1]/P0001 ,
		_w1240_,
		_w6635_
	);
	LUT2 #(
		.INIT('h8)
	) name6104 (
		\sa31_reg[7]/P0001 ,
		_w6162_,
		_w6636_
	);
	LUT2 #(
		.INIT('h1)
	) name6105 (
		_w1160_,
		_w1217_,
		_w6637_
	);
	LUT2 #(
		.INIT('h1)
	) name6106 (
		\sa31_reg[2]/P0001 ,
		_w6637_,
		_w6638_
	);
	LUT2 #(
		.INIT('h4)
	) name6107 (
		_w6553_,
		_w6635_,
		_w6639_
	);
	LUT2 #(
		.INIT('h1)
	) name6108 (
		_w6636_,
		_w6638_,
		_w6640_
	);
	LUT2 #(
		.INIT('h8)
	) name6109 (
		_w6639_,
		_w6640_,
		_w6641_
	);
	LUT2 #(
		.INIT('h1)
	) name6110 (
		_w5263_,
		_w6136_,
		_w6642_
	);
	LUT2 #(
		.INIT('h2)
	) name6111 (
		\sa31_reg[7]/P0001 ,
		_w6642_,
		_w6643_
	);
	LUT2 #(
		.INIT('h8)
	) name6112 (
		_w1265_,
		_w6092_,
		_w6644_
	);
	LUT2 #(
		.INIT('h2)
	) name6113 (
		_w6099_,
		_w6644_,
		_w6645_
	);
	LUT2 #(
		.INIT('h4)
	) name6114 (
		_w6643_,
		_w6645_,
		_w6646_
	);
	LUT2 #(
		.INIT('h1)
	) name6115 (
		_w6641_,
		_w6646_,
		_w6647_
	);
	LUT2 #(
		.INIT('h8)
	) name6116 (
		_w1225_,
		_w6098_,
		_w6648_
	);
	LUT2 #(
		.INIT('h1)
	) name6117 (
		_w6634_,
		_w6648_,
		_w6649_
	);
	LUT2 #(
		.INIT('h4)
	) name6118 (
		_w6647_,
		_w6649_,
		_w6650_
	);
	LUT2 #(
		.INIT('h1)
	) name6119 (
		\sa31_reg[0]/P0002 ,
		_w6650_,
		_w6651_
	);
	LUT2 #(
		.INIT('h1)
	) name6120 (
		_w6618_,
		_w6622_,
		_w6652_
	);
	LUT2 #(
		.INIT('h4)
	) name6121 (
		_w6626_,
		_w6652_,
		_w6653_
	);
	LUT2 #(
		.INIT('h4)
	) name6122 (
		_w6616_,
		_w6653_,
		_w6654_
	);
	LUT2 #(
		.INIT('h4)
	) name6123 (
		_w6588_,
		_w6654_,
		_w6655_
	);
	LUT2 #(
		.INIT('h4)
	) name6124 (
		_w6610_,
		_w6655_,
		_w6656_
	);
	LUT2 #(
		.INIT('h4)
	) name6125 (
		_w6651_,
		_w6656_,
		_w6657_
	);
	LUT2 #(
		.INIT('h2)
	) name6126 (
		_w6568_,
		_w6657_,
		_w6658_
	);
	LUT2 #(
		.INIT('h4)
	) name6127 (
		_w6568_,
		_w6657_,
		_w6659_
	);
	LUT2 #(
		.INIT('h1)
	) name6128 (
		_w6658_,
		_w6659_,
		_w6660_
	);
	LUT2 #(
		.INIT('h1)
	) name6129 (
		_w781_,
		_w5599_,
		_w6661_
	);
	LUT2 #(
		.INIT('h2)
	) name6130 (
		\sa20_reg[2]/P0001 ,
		_w6661_,
		_w6662_
	);
	LUT2 #(
		.INIT('h2)
	) name6131 (
		\sa20_reg[4]/P0001 ,
		_w698_,
		_w6663_
	);
	LUT2 #(
		.INIT('h2)
	) name6132 (
		_w748_,
		_w6663_,
		_w6664_
	);
	LUT2 #(
		.INIT('h1)
	) name6133 (
		_w769_,
		_w6664_,
		_w6665_
	);
	LUT2 #(
		.INIT('h1)
	) name6134 (
		\sa20_reg[2]/P0001 ,
		_w6665_,
		_w6666_
	);
	LUT2 #(
		.INIT('h4)
	) name6135 (
		_w5620_,
		_w5873_,
		_w6667_
	);
	LUT2 #(
		.INIT('h4)
	) name6136 (
		_w6662_,
		_w6667_,
		_w6668_
	);
	LUT2 #(
		.INIT('h4)
	) name6137 (
		_w6666_,
		_w6668_,
		_w6669_
	);
	LUT2 #(
		.INIT('h2)
	) name6138 (
		\sa20_reg[1]/P0001 ,
		_w6669_,
		_w6670_
	);
	LUT2 #(
		.INIT('h1)
	) name6139 (
		_w795_,
		_w5973_,
		_w6671_
	);
	LUT2 #(
		.INIT('h2)
	) name6140 (
		\sa20_reg[2]/P0001 ,
		_w6671_,
		_w6672_
	);
	LUT2 #(
		.INIT('h1)
	) name6141 (
		_w738_,
		_w832_,
		_w6673_
	);
	LUT2 #(
		.INIT('h1)
	) name6142 (
		\sa20_reg[2]/P0001 ,
		_w6673_,
		_w6674_
	);
	LUT2 #(
		.INIT('h1)
	) name6143 (
		_w822_,
		_w6043_,
		_w6675_
	);
	LUT2 #(
		.INIT('h4)
	) name6144 (
		_w6672_,
		_w6675_,
		_w6676_
	);
	LUT2 #(
		.INIT('h4)
	) name6145 (
		_w6674_,
		_w6676_,
		_w6677_
	);
	LUT2 #(
		.INIT('h1)
	) name6146 (
		\sa20_reg[1]/P0001 ,
		_w6677_,
		_w6678_
	);
	LUT2 #(
		.INIT('h1)
	) name6147 (
		_w5892_,
		_w6043_,
		_w6679_
	);
	LUT2 #(
		.INIT('h1)
	) name6148 (
		\sa20_reg[2]/P0001 ,
		_w6679_,
		_w6680_
	);
	LUT2 #(
		.INIT('h1)
	) name6149 (
		_w709_,
		_w820_,
		_w6681_
	);
	LUT2 #(
		.INIT('h2)
	) name6150 (
		_w819_,
		_w6681_,
		_w6682_
	);
	LUT2 #(
		.INIT('h1)
	) name6151 (
		_w809_,
		_w5928_,
		_w6683_
	);
	LUT2 #(
		.INIT('h4)
	) name6152 (
		_w6682_,
		_w6683_,
		_w6684_
	);
	LUT2 #(
		.INIT('h4)
	) name6153 (
		_w6680_,
		_w6684_,
		_w6685_
	);
	LUT2 #(
		.INIT('h4)
	) name6154 (
		_w6670_,
		_w6685_,
		_w6686_
	);
	LUT2 #(
		.INIT('h4)
	) name6155 (
		_w6678_,
		_w6686_,
		_w6687_
	);
	LUT2 #(
		.INIT('h1)
	) name6156 (
		\sa20_reg[0]/P0001 ,
		_w6687_,
		_w6688_
	);
	LUT2 #(
		.INIT('h8)
	) name6157 (
		_w716_,
		_w5858_,
		_w6689_
	);
	LUT2 #(
		.INIT('h1)
	) name6158 (
		_w721_,
		_w6689_,
		_w6690_
	);
	LUT2 #(
		.INIT('h8)
	) name6159 (
		\sa20_reg[7]/NET0131 ,
		_w698_,
		_w6691_
	);
	LUT2 #(
		.INIT('h1)
	) name6160 (
		_w767_,
		_w5529_,
		_w6692_
	);
	LUT2 #(
		.INIT('h4)
	) name6161 (
		_w6691_,
		_w6692_,
		_w6693_
	);
	LUT2 #(
		.INIT('h2)
	) name6162 (
		\sa20_reg[2]/P0001 ,
		_w6693_,
		_w6694_
	);
	LUT2 #(
		.INIT('h2)
	) name6163 (
		_w6690_,
		_w6694_,
		_w6695_
	);
	LUT2 #(
		.INIT('h2)
	) name6164 (
		\sa20_reg[1]/P0001 ,
		_w6695_,
		_w6696_
	);
	LUT2 #(
		.INIT('h2)
	) name6165 (
		_w716_,
		_w826_,
		_w6697_
	);
	LUT2 #(
		.INIT('h4)
	) name6166 (
		_w717_,
		_w6697_,
		_w6698_
	);
	LUT2 #(
		.INIT('h4)
	) name6167 (
		\sa20_reg[6]/NET0131 ,
		_w5908_,
		_w6699_
	);
	LUT2 #(
		.INIT('h1)
	) name6168 (
		_w5567_,
		_w5843_,
		_w6700_
	);
	LUT2 #(
		.INIT('h4)
	) name6169 (
		_w6698_,
		_w6700_,
		_w6701_
	);
	LUT2 #(
		.INIT('h4)
	) name6170 (
		_w6699_,
		_w6701_,
		_w6702_
	);
	LUT2 #(
		.INIT('h1)
	) name6171 (
		\sa20_reg[1]/P0001 ,
		_w6702_,
		_w6703_
	);
	LUT2 #(
		.INIT('h2)
	) name6172 (
		_w737_,
		_w5582_,
		_w6704_
	);
	LUT2 #(
		.INIT('h8)
	) name6173 (
		\sa20_reg[4]/P0001 ,
		_w725_,
		_w6705_
	);
	LUT2 #(
		.INIT('h1)
	) name6174 (
		_w834_,
		_w5567_,
		_w6706_
	);
	LUT2 #(
		.INIT('h1)
	) name6175 (
		_w5606_,
		_w5973_,
		_w6707_
	);
	LUT2 #(
		.INIT('h8)
	) name6176 (
		_w6706_,
		_w6707_,
		_w6708_
	);
	LUT2 #(
		.INIT('h1)
	) name6177 (
		\sa20_reg[2]/P0001 ,
		_w6708_,
		_w6709_
	);
	LUT2 #(
		.INIT('h1)
	) name6178 (
		_w6704_,
		_w6705_,
		_w6710_
	);
	LUT2 #(
		.INIT('h4)
	) name6179 (
		_w6703_,
		_w6710_,
		_w6711_
	);
	LUT2 #(
		.INIT('h4)
	) name6180 (
		_w6709_,
		_w6711_,
		_w6712_
	);
	LUT2 #(
		.INIT('h4)
	) name6181 (
		_w6696_,
		_w6712_,
		_w6713_
	);
	LUT2 #(
		.INIT('h2)
	) name6182 (
		\sa20_reg[0]/P0001 ,
		_w6713_,
		_w6714_
	);
	LUT2 #(
		.INIT('h4)
	) name6183 (
		\sa20_reg[3]/P0001 ,
		_w690_,
		_w6715_
	);
	LUT2 #(
		.INIT('h1)
	) name6184 (
		_w710_,
		_w6715_,
		_w6716_
	);
	LUT2 #(
		.INIT('h4)
	) name6185 (
		_w5620_,
		_w6716_,
		_w6717_
	);
	LUT2 #(
		.INIT('h1)
	) name6186 (
		_w714_,
		_w6717_,
		_w6718_
	);
	LUT2 #(
		.INIT('h1)
	) name6187 (
		_w695_,
		_w6718_,
		_w6719_
	);
	LUT2 #(
		.INIT('h2)
	) name6188 (
		_w815_,
		_w6719_,
		_w6720_
	);
	LUT2 #(
		.INIT('h1)
	) name6189 (
		_w721_,
		_w5532_,
		_w6721_
	);
	LUT2 #(
		.INIT('h2)
	) name6190 (
		\sa20_reg[3]/P0001 ,
		_w6721_,
		_w6722_
	);
	LUT2 #(
		.INIT('h1)
	) name6191 (
		_w768_,
		_w6722_,
		_w6723_
	);
	LUT2 #(
		.INIT('h2)
	) name6192 (
		_w806_,
		_w6723_,
		_w6724_
	);
	LUT2 #(
		.INIT('h1)
	) name6193 (
		_w710_,
		_w5998_,
		_w6725_
	);
	LUT2 #(
		.INIT('h2)
	) name6194 (
		_w761_,
		_w6725_,
		_w6726_
	);
	LUT2 #(
		.INIT('h4)
	) name6195 (
		\sa20_reg[1]/P0001 ,
		\sa20_reg[2]/P0001 ,
		_w6727_
	);
	LUT2 #(
		.INIT('h8)
	) name6196 (
		_w708_,
		_w736_,
		_w6728_
	);
	LUT2 #(
		.INIT('h1)
	) name6197 (
		_w809_,
		_w6728_,
		_w6729_
	);
	LUT2 #(
		.INIT('h4)
	) name6198 (
		_w703_,
		_w6729_,
		_w6730_
	);
	LUT2 #(
		.INIT('h2)
	) name6199 (
		_w6727_,
		_w6730_,
		_w6731_
	);
	LUT2 #(
		.INIT('h1)
	) name6200 (
		_w746_,
		_w5591_,
		_w6732_
	);
	LUT2 #(
		.INIT('h4)
	) name6201 (
		_w5894_,
		_w6732_,
		_w6733_
	);
	LUT2 #(
		.INIT('h1)
	) name6202 (
		\sa20_reg[2]/P0001 ,
		_w6733_,
		_w6734_
	);
	LUT2 #(
		.INIT('h1)
	) name6203 (
		_w752_,
		_w6036_,
		_w6735_
	);
	LUT2 #(
		.INIT('h4)
	) name6204 (
		_w6734_,
		_w6735_,
		_w6736_
	);
	LUT2 #(
		.INIT('h1)
	) name6205 (
		\sa20_reg[1]/P0001 ,
		_w6736_,
		_w6737_
	);
	LUT2 #(
		.INIT('h1)
	) name6206 (
		_w6726_,
		_w6731_,
		_w6738_
	);
	LUT2 #(
		.INIT('h4)
	) name6207 (
		_w6724_,
		_w6738_,
		_w6739_
	);
	LUT2 #(
		.INIT('h4)
	) name6208 (
		_w6720_,
		_w6739_,
		_w6740_
	);
	LUT2 #(
		.INIT('h4)
	) name6209 (
		_w6737_,
		_w6740_,
		_w6741_
	);
	LUT2 #(
		.INIT('h4)
	) name6210 (
		_w6688_,
		_w6741_,
		_w6742_
	);
	LUT2 #(
		.INIT('h4)
	) name6211 (
		_w6714_,
		_w6742_,
		_w6743_
	);
	LUT2 #(
		.INIT('h2)
	) name6212 (
		\u0_w_reg[2][1]/P0001 ,
		_w6743_,
		_w6744_
	);
	LUT2 #(
		.INIT('h4)
	) name6213 (
		\u0_w_reg[2][1]/P0001 ,
		_w6743_,
		_w6745_
	);
	LUT2 #(
		.INIT('h1)
	) name6214 (
		_w6744_,
		_w6745_,
		_w6746_
	);
	LUT2 #(
		.INIT('h8)
	) name6215 (
		_w6660_,
		_w6746_,
		_w6747_
	);
	LUT2 #(
		.INIT('h1)
	) name6216 (
		_w6660_,
		_w6746_,
		_w6748_
	);
	LUT2 #(
		.INIT('h1)
	) name6217 (
		_w6747_,
		_w6748_,
		_w6749_
	);
	LUT2 #(
		.INIT('h1)
	) name6218 (
		_w6478_,
		_w6749_,
		_w6750_
	);
	LUT2 #(
		.INIT('h8)
	) name6219 (
		_w6478_,
		_w6749_,
		_w6751_
	);
	LUT2 #(
		.INIT('h1)
	) name6220 (
		\ld_r_reg/P0001 ,
		_w6750_,
		_w6752_
	);
	LUT2 #(
		.INIT('h4)
	) name6221 (
		_w6751_,
		_w6752_,
		_w6753_
	);
	LUT2 #(
		.INIT('h1)
	) name6222 (
		\text_in_r_reg[33]/P0001 ,
		\u0_w_reg[2][1]/P0001 ,
		_w6754_
	);
	LUT2 #(
		.INIT('h8)
	) name6223 (
		\text_in_r_reg[33]/P0001 ,
		\u0_w_reg[2][1]/P0001 ,
		_w6755_
	);
	LUT2 #(
		.INIT('h2)
	) name6224 (
		\ld_r_reg/P0001 ,
		_w6754_,
		_w6756_
	);
	LUT2 #(
		.INIT('h4)
	) name6225 (
		_w6755_,
		_w6756_,
		_w6757_
	);
	LUT2 #(
		.INIT('h1)
	) name6226 (
		_w6753_,
		_w6757_,
		_w6758_
	);
	LUT2 #(
		.INIT('h8)
	) name6227 (
		\sa31_reg[4]/P0001 ,
		_w6483_,
		_w6759_
	);
	LUT2 #(
		.INIT('h1)
	) name6228 (
		_w1269_,
		_w6530_,
		_w6760_
	);
	LUT2 #(
		.INIT('h4)
	) name6229 (
		_w6759_,
		_w6760_,
		_w6761_
	);
	LUT2 #(
		.INIT('h1)
	) name6230 (
		\sa31_reg[2]/P0001 ,
		_w6761_,
		_w6762_
	);
	LUT2 #(
		.INIT('h1)
	) name6231 (
		_w1280_,
		_w6581_,
		_w6763_
	);
	LUT2 #(
		.INIT('h2)
	) name6232 (
		\sa31_reg[2]/P0001 ,
		_w6763_,
		_w6764_
	);
	LUT2 #(
		.INIT('h2)
	) name6233 (
		\sa31_reg[1]/P0001 ,
		_w5204_,
		_w6765_
	);
	LUT2 #(
		.INIT('h8)
	) name6234 (
		_w5272_,
		_w6765_,
		_w6766_
	);
	LUT2 #(
		.INIT('h4)
	) name6235 (
		_w6762_,
		_w6766_,
		_w6767_
	);
	LUT2 #(
		.INIT('h4)
	) name6236 (
		_w6764_,
		_w6767_,
		_w6768_
	);
	LUT2 #(
		.INIT('h8)
	) name6237 (
		\sa31_reg[6]/NET0131 ,
		_w1181_,
		_w6769_
	);
	LUT2 #(
		.INIT('h1)
	) name6238 (
		_w6119_,
		_w6491_,
		_w6770_
	);
	LUT2 #(
		.INIT('h2)
	) name6239 (
		\sa31_reg[2]/P0001 ,
		_w6770_,
		_w6771_
	);
	LUT2 #(
		.INIT('h1)
	) name6240 (
		_w1154_,
		_w1239_,
		_w6772_
	);
	LUT2 #(
		.INIT('h1)
	) name6241 (
		\sa31_reg[2]/P0001 ,
		_w6772_,
		_w6773_
	);
	LUT2 #(
		.INIT('h1)
	) name6242 (
		\sa31_reg[1]/P0001 ,
		_w6160_,
		_w6774_
	);
	LUT2 #(
		.INIT('h4)
	) name6243 (
		_w6769_,
		_w6774_,
		_w6775_
	);
	LUT2 #(
		.INIT('h4)
	) name6244 (
		_w6771_,
		_w6775_,
		_w6776_
	);
	LUT2 #(
		.INIT('h4)
	) name6245 (
		_w6773_,
		_w6776_,
		_w6777_
	);
	LUT2 #(
		.INIT('h1)
	) name6246 (
		_w6768_,
		_w6777_,
		_w6778_
	);
	LUT2 #(
		.INIT('h4)
	) name6247 (
		_w5250_,
		_w6161_,
		_w6779_
	);
	LUT2 #(
		.INIT('h2)
	) name6248 (
		\sa31_reg[2]/P0001 ,
		_w1230_,
		_w6780_
	);
	LUT2 #(
		.INIT('h4)
	) name6249 (
		_w1220_,
		_w6780_,
		_w6781_
	);
	LUT2 #(
		.INIT('h1)
	) name6250 (
		_w6779_,
		_w6781_,
		_w6782_
	);
	LUT2 #(
		.INIT('h1)
	) name6251 (
		_w1234_,
		_w5295_,
		_w6783_
	);
	LUT2 #(
		.INIT('h4)
	) name6252 (
		_w6782_,
		_w6783_,
		_w6784_
	);
	LUT2 #(
		.INIT('h4)
	) name6253 (
		_w6778_,
		_w6784_,
		_w6785_
	);
	LUT2 #(
		.INIT('h1)
	) name6254 (
		\sa31_reg[0]/P0002 ,
		_w6785_,
		_w6786_
	);
	LUT2 #(
		.INIT('h8)
	) name6255 (
		\sa31_reg[3]/P0001 ,
		_w6488_,
		_w6787_
	);
	LUT2 #(
		.INIT('h1)
	) name6256 (
		_w1183_,
		_w6787_,
		_w6788_
	);
	LUT2 #(
		.INIT('h8)
	) name6257 (
		\sa31_reg[4]/P0001 ,
		_w1151_,
		_w6789_
	);
	LUT2 #(
		.INIT('h8)
	) name6258 (
		\sa31_reg[7]/P0001 ,
		_w5269_,
		_w6790_
	);
	LUT2 #(
		.INIT('h1)
	) name6259 (
		_w6571_,
		_w6789_,
		_w6791_
	);
	LUT2 #(
		.INIT('h4)
	) name6260 (
		_w6790_,
		_w6791_,
		_w6792_
	);
	LUT2 #(
		.INIT('h2)
	) name6261 (
		\sa31_reg[2]/P0001 ,
		_w6792_,
		_w6793_
	);
	LUT2 #(
		.INIT('h2)
	) name6262 (
		_w6788_,
		_w6793_,
		_w6794_
	);
	LUT2 #(
		.INIT('h2)
	) name6263 (
		\sa31_reg[1]/P0001 ,
		_w6794_,
		_w6795_
	);
	LUT2 #(
		.INIT('h2)
	) name6264 (
		_w5205_,
		_w6136_,
		_w6796_
	);
	LUT2 #(
		.INIT('h1)
	) name6265 (
		_w6627_,
		_w6796_,
		_w6797_
	);
	LUT2 #(
		.INIT('h1)
	) name6266 (
		\sa31_reg[3]/P0001 ,
		_w6797_,
		_w6798_
	);
	LUT2 #(
		.INIT('h1)
	) name6267 (
		_w1240_,
		_w6110_,
		_w6799_
	);
	LUT2 #(
		.INIT('h1)
	) name6268 (
		_w6491_,
		_w6627_,
		_w6800_
	);
	LUT2 #(
		.INIT('h8)
	) name6269 (
		_w6799_,
		_w6800_,
		_w6801_
	);
	LUT2 #(
		.INIT('h1)
	) name6270 (
		\sa31_reg[2]/P0001 ,
		_w6801_,
		_w6802_
	);
	LUT2 #(
		.INIT('h2)
	) name6271 (
		_w1159_,
		_w1180_,
		_w6803_
	);
	LUT2 #(
		.INIT('h4)
	) name6272 (
		_w1256_,
		_w6803_,
		_w6804_
	);
	LUT2 #(
		.INIT('h8)
	) name6273 (
		_w1153_,
		_w1178_,
		_w6805_
	);
	LUT2 #(
		.INIT('h8)
	) name6274 (
		_w1146_,
		_w5238_,
		_w6806_
	);
	LUT2 #(
		.INIT('h1)
	) name6275 (
		_w6110_,
		_w6806_,
		_w6807_
	);
	LUT2 #(
		.INIT('h4)
	) name6276 (
		_w6804_,
		_w6807_,
		_w6808_
	);
	LUT2 #(
		.INIT('h4)
	) name6277 (
		_w6805_,
		_w6808_,
		_w6809_
	);
	LUT2 #(
		.INIT('h1)
	) name6278 (
		\sa31_reg[1]/P0001 ,
		_w6809_,
		_w6810_
	);
	LUT2 #(
		.INIT('h1)
	) name6279 (
		_w6798_,
		_w6802_,
		_w6811_
	);
	LUT2 #(
		.INIT('h4)
	) name6280 (
		_w6810_,
		_w6811_,
		_w6812_
	);
	LUT2 #(
		.INIT('h4)
	) name6281 (
		_w6795_,
		_w6812_,
		_w6813_
	);
	LUT2 #(
		.INIT('h2)
	) name6282 (
		\sa31_reg[0]/P0002 ,
		_w6813_,
		_w6814_
	);
	LUT2 #(
		.INIT('h4)
	) name6283 (
		\sa31_reg[5]/P0001 ,
		_w1269_,
		_w6815_
	);
	LUT2 #(
		.INIT('h1)
	) name6284 (
		_w1202_,
		_w1234_,
		_w6816_
	);
	LUT2 #(
		.INIT('h4)
	) name6285 (
		_w6815_,
		_w6816_,
		_w6817_
	);
	LUT2 #(
		.INIT('h2)
	) name6286 (
		_w6514_,
		_w6817_,
		_w6818_
	);
	LUT2 #(
		.INIT('h1)
	) name6287 (
		_w5204_,
		_w6543_,
		_w6819_
	);
	LUT2 #(
		.INIT('h4)
	) name6288 (
		_w1195_,
		_w6819_,
		_w6820_
	);
	LUT2 #(
		.INIT('h1)
	) name6289 (
		_w1205_,
		_w6168_,
		_w6821_
	);
	LUT2 #(
		.INIT('h8)
	) name6290 (
		_w6820_,
		_w6821_,
		_w6822_
	);
	LUT2 #(
		.INIT('h2)
	) name6291 (
		_w1224_,
		_w6822_,
		_w6823_
	);
	LUT2 #(
		.INIT('h4)
	) name6292 (
		\sa31_reg[6]/NET0131 ,
		_w6644_,
		_w6824_
	);
	LUT2 #(
		.INIT('h1)
	) name6293 (
		_w1183_,
		_w1277_,
		_w6825_
	);
	LUT2 #(
		.INIT('h2)
	) name6294 (
		\sa31_reg[3]/P0001 ,
		_w6825_,
		_w6826_
	);
	LUT2 #(
		.INIT('h1)
	) name6295 (
		_w6636_,
		_w6826_,
		_w6827_
	);
	LUT2 #(
		.INIT('h2)
	) name6296 (
		_w1232_,
		_w6827_,
		_w6828_
	);
	LUT2 #(
		.INIT('h1)
	) name6297 (
		_w1168_,
		_w1217_,
		_w6829_
	);
	LUT2 #(
		.INIT('h4)
	) name6298 (
		_w5253_,
		_w6829_,
		_w6830_
	);
	LUT2 #(
		.INIT('h1)
	) name6299 (
		\sa31_reg[2]/P0001 ,
		_w6830_,
		_w6831_
	);
	LUT2 #(
		.INIT('h8)
	) name6300 (
		_w1160_,
		_w1182_,
		_w6832_
	);
	LUT2 #(
		.INIT('h1)
	) name6301 (
		_w1161_,
		_w6832_,
		_w6833_
	);
	LUT2 #(
		.INIT('h4)
	) name6302 (
		_w6831_,
		_w6833_,
		_w6834_
	);
	LUT2 #(
		.INIT('h1)
	) name6303 (
		\sa31_reg[1]/P0001 ,
		_w6834_,
		_w6835_
	);
	LUT2 #(
		.INIT('h1)
	) name6304 (
		_w6648_,
		_w6824_,
		_w6836_
	);
	LUT2 #(
		.INIT('h4)
	) name6305 (
		_w6818_,
		_w6836_,
		_w6837_
	);
	LUT2 #(
		.INIT('h1)
	) name6306 (
		_w6823_,
		_w6828_,
		_w6838_
	);
	LUT2 #(
		.INIT('h8)
	) name6307 (
		_w6837_,
		_w6838_,
		_w6839_
	);
	LUT2 #(
		.INIT('h4)
	) name6308 (
		_w6835_,
		_w6839_,
		_w6840_
	);
	LUT2 #(
		.INIT('h4)
	) name6309 (
		_w6786_,
		_w6840_,
		_w6841_
	);
	LUT2 #(
		.INIT('h4)
	) name6310 (
		_w6814_,
		_w6841_,
		_w6842_
	);
	LUT2 #(
		.INIT('h2)
	) name6311 (
		\u0_w_reg[2][9]/P0001 ,
		_w6842_,
		_w6843_
	);
	LUT2 #(
		.INIT('h4)
	) name6312 (
		\u0_w_reg[2][9]/P0001 ,
		_w6842_,
		_w6844_
	);
	LUT2 #(
		.INIT('h1)
	) name6313 (
		_w6843_,
		_w6844_,
		_w6845_
	);
	LUT2 #(
		.INIT('h8)
	) name6314 (
		_w6660_,
		_w6845_,
		_w6846_
	);
	LUT2 #(
		.INIT('h1)
	) name6315 (
		_w6660_,
		_w6845_,
		_w6847_
	);
	LUT2 #(
		.INIT('h1)
	) name6316 (
		_w6846_,
		_w6847_,
		_w6848_
	);
	LUT2 #(
		.INIT('h4)
	) name6317 (
		\sa20_reg[4]/P0001 ,
		_w706_,
		_w6849_
	);
	LUT2 #(
		.INIT('h4)
	) name6318 (
		\sa20_reg[2]/P0001 ,
		_w5857_,
		_w6850_
	);
	LUT2 #(
		.INIT('h4)
	) name6319 (
		\sa20_reg[3]/P0001 ,
		_w820_,
		_w6851_
	);
	LUT2 #(
		.INIT('h1)
	) name6320 (
		_w5556_,
		_w5907_,
		_w6852_
	);
	LUT2 #(
		.INIT('h4)
	) name6321 (
		_w6851_,
		_w6852_,
		_w6853_
	);
	LUT2 #(
		.INIT('h2)
	) name6322 (
		\sa20_reg[2]/P0001 ,
		_w6853_,
		_w6854_
	);
	LUT2 #(
		.INIT('h1)
	) name6323 (
		_w5600_,
		_w5895_,
		_w6855_
	);
	LUT2 #(
		.INIT('h4)
	) name6324 (
		_w6849_,
		_w6855_,
		_w6856_
	);
	LUT2 #(
		.INIT('h4)
	) name6325 (
		_w6850_,
		_w6856_,
		_w6857_
	);
	LUT2 #(
		.INIT('h4)
	) name6326 (
		_w6854_,
		_w6857_,
		_w6858_
	);
	LUT2 #(
		.INIT('h1)
	) name6327 (
		\sa20_reg[1]/P0001 ,
		_w6858_,
		_w6859_
	);
	LUT2 #(
		.INIT('h1)
	) name6328 (
		_w746_,
		_w5981_,
		_w6860_
	);
	LUT2 #(
		.INIT('h8)
	) name6329 (
		_w5893_,
		_w6860_,
		_w6861_
	);
	LUT2 #(
		.INIT('h2)
	) name6330 (
		\sa20_reg[2]/P0001 ,
		_w6861_,
		_w6862_
	);
	LUT2 #(
		.INIT('h1)
	) name6331 (
		_w5549_,
		_w5605_,
		_w6863_
	);
	LUT2 #(
		.INIT('h1)
	) name6332 (
		\sa20_reg[2]/P0001 ,
		_w6863_,
		_w6864_
	);
	LUT2 #(
		.INIT('h1)
	) name6333 (
		_w709_,
		_w735_,
		_w6865_
	);
	LUT2 #(
		.INIT('h2)
	) name6334 (
		_w763_,
		_w6865_,
		_w6866_
	);
	LUT2 #(
		.INIT('h1)
	) name6335 (
		\sa20_reg[2]/P0001 ,
		_w690_,
		_w6867_
	);
	LUT2 #(
		.INIT('h1)
	) name6336 (
		\sa20_reg[5]/P0001 ,
		_w723_,
		_w6868_
	);
	LUT2 #(
		.INIT('h2)
	) name6337 (
		_w6867_,
		_w6868_,
		_w6869_
	);
	LUT2 #(
		.INIT('h1)
	) name6338 (
		_w832_,
		_w6869_,
		_w6870_
	);
	LUT2 #(
		.INIT('h2)
	) name6339 (
		\sa20_reg[1]/P0001 ,
		_w6870_,
		_w6871_
	);
	LUT2 #(
		.INIT('h1)
	) name6340 (
		_w5973_,
		_w6029_,
		_w6872_
	);
	LUT2 #(
		.INIT('h4)
	) name6341 (
		_w6866_,
		_w6872_,
		_w6873_
	);
	LUT2 #(
		.INIT('h4)
	) name6342 (
		_w6864_,
		_w6873_,
		_w6874_
	);
	LUT2 #(
		.INIT('h4)
	) name6343 (
		_w6871_,
		_w6874_,
		_w6875_
	);
	LUT2 #(
		.INIT('h4)
	) name6344 (
		_w6862_,
		_w6875_,
		_w6876_
	);
	LUT2 #(
		.INIT('h4)
	) name6345 (
		_w6859_,
		_w6876_,
		_w6877_
	);
	LUT2 #(
		.INIT('h2)
	) name6346 (
		\sa20_reg[0]/P0001 ,
		_w6877_,
		_w6878_
	);
	LUT2 #(
		.INIT('h8)
	) name6347 (
		\sa20_reg[6]/NET0131 ,
		_w833_,
		_w6879_
	);
	LUT2 #(
		.INIT('h1)
	) name6348 (
		_w5892_,
		_w6879_,
		_w6880_
	);
	LUT2 #(
		.INIT('h4)
	) name6349 (
		_w800_,
		_w6880_,
		_w6881_
	);
	LUT2 #(
		.INIT('h1)
	) name6350 (
		\sa20_reg[2]/P0001 ,
		_w6881_,
		_w6882_
	);
	LUT2 #(
		.INIT('h1)
	) name6351 (
		_w724_,
		_w735_,
		_w6883_
	);
	LUT2 #(
		.INIT('h8)
	) name6352 (
		\sa20_reg[2]/P0001 ,
		_w745_,
		_w6884_
	);
	LUT2 #(
		.INIT('h4)
	) name6353 (
		_w6883_,
		_w6884_,
		_w6885_
	);
	LUT2 #(
		.INIT('h4)
	) name6354 (
		_w698_,
		_w744_,
		_w6886_
	);
	LUT2 #(
		.INIT('h8)
	) name6355 (
		_w6727_,
		_w6886_,
		_w6887_
	);
	LUT2 #(
		.INIT('h1)
	) name6356 (
		\sa20_reg[3]/P0001 ,
		_w5568_,
		_w6888_
	);
	LUT2 #(
		.INIT('h1)
	) name6357 (
		_w6007_,
		_w6888_,
		_w6889_
	);
	LUT2 #(
		.INIT('h1)
	) name6358 (
		\sa20_reg[1]/P0001 ,
		_w6889_,
		_w6890_
	);
	LUT2 #(
		.INIT('h8)
	) name6359 (
		_w720_,
		_w747_,
		_w6891_
	);
	LUT2 #(
		.INIT('h1)
	) name6360 (
		_w716_,
		_w723_,
		_w6892_
	);
	LUT2 #(
		.INIT('h1)
	) name6361 (
		_w6697_,
		_w6892_,
		_w6893_
	);
	LUT2 #(
		.INIT('h8)
	) name6362 (
		\sa20_reg[2]/P0001 ,
		_w698_,
		_w6894_
	);
	LUT2 #(
		.INIT('h8)
	) name6363 (
		_w777_,
		_w6894_,
		_w6895_
	);
	LUT2 #(
		.INIT('h1)
	) name6364 (
		_w6891_,
		_w6893_,
		_w6896_
	);
	LUT2 #(
		.INIT('h4)
	) name6365 (
		_w6895_,
		_w6896_,
		_w6897_
	);
	LUT2 #(
		.INIT('h2)
	) name6366 (
		\sa20_reg[1]/P0001 ,
		_w6897_,
		_w6898_
	);
	LUT2 #(
		.INIT('h1)
	) name6367 (
		_w6885_,
		_w6887_,
		_w6899_
	);
	LUT2 #(
		.INIT('h4)
	) name6368 (
		_w6882_,
		_w6899_,
		_w6900_
	);
	LUT2 #(
		.INIT('h1)
	) name6369 (
		_w6890_,
		_w6898_,
		_w6901_
	);
	LUT2 #(
		.INIT('h8)
	) name6370 (
		_w6900_,
		_w6901_,
		_w6902_
	);
	LUT2 #(
		.INIT('h1)
	) name6371 (
		\sa20_reg[0]/P0001 ,
		_w6902_,
		_w6903_
	);
	LUT2 #(
		.INIT('h8)
	) name6372 (
		_w729_,
		_w5523_,
		_w6904_
	);
	LUT2 #(
		.INIT('h8)
	) name6373 (
		_w5526_,
		_w5973_,
		_w6905_
	);
	LUT2 #(
		.INIT('h8)
	) name6374 (
		\sa20_reg[2]/P0001 ,
		_w799_,
		_w6906_
	);
	LUT2 #(
		.INIT('h1)
	) name6375 (
		_w701_,
		_w5544_,
		_w6907_
	);
	LUT2 #(
		.INIT('h2)
	) name6376 (
		_w6906_,
		_w6907_,
		_w6908_
	);
	LUT2 #(
		.INIT('h8)
	) name6377 (
		_w695_,
		_w763_,
		_w6909_
	);
	LUT2 #(
		.INIT('h4)
	) name6378 (
		_w694_,
		_w5527_,
		_w6910_
	);
	LUT2 #(
		.INIT('h1)
	) name6379 (
		_w5968_,
		_w6910_,
		_w6911_
	);
	LUT2 #(
		.INIT('h1)
	) name6380 (
		\sa20_reg[2]/P0001 ,
		_w6911_,
		_w6912_
	);
	LUT2 #(
		.INIT('h1)
	) name6381 (
		\sa20_reg[1]/P0001 ,
		_w6909_,
		_w6913_
	);
	LUT2 #(
		.INIT('h4)
	) name6382 (
		_w5928_,
		_w6913_,
		_w6914_
	);
	LUT2 #(
		.INIT('h4)
	) name6383 (
		_w6908_,
		_w6914_,
		_w6915_
	);
	LUT2 #(
		.INIT('h4)
	) name6384 (
		_w6912_,
		_w6915_,
		_w6916_
	);
	LUT2 #(
		.INIT('h8)
	) name6385 (
		\sa20_reg[2]/P0001 ,
		_w707_,
		_w6917_
	);
	LUT2 #(
		.INIT('h1)
	) name6386 (
		\sa20_reg[2]/P0001 ,
		_w5617_,
		_w6918_
	);
	LUT2 #(
		.INIT('h1)
	) name6387 (
		_w5836_,
		_w6918_,
		_w6919_
	);
	LUT2 #(
		.INIT('h1)
	) name6388 (
		_w824_,
		_w6917_,
		_w6920_
	);
	LUT2 #(
		.INIT('h8)
	) name6389 (
		_w5996_,
		_w6920_,
		_w6921_
	);
	LUT2 #(
		.INIT('h4)
	) name6390 (
		_w6919_,
		_w6921_,
		_w6922_
	);
	LUT2 #(
		.INIT('h1)
	) name6391 (
		_w6916_,
		_w6922_,
		_w6923_
	);
	LUT2 #(
		.INIT('h1)
	) name6392 (
		_w6904_,
		_w6905_,
		_w6924_
	);
	LUT2 #(
		.INIT('h4)
	) name6393 (
		_w6923_,
		_w6924_,
		_w6925_
	);
	LUT2 #(
		.INIT('h4)
	) name6394 (
		_w6903_,
		_w6925_,
		_w6926_
	);
	LUT2 #(
		.INIT('h4)
	) name6395 (
		_w6878_,
		_w6926_,
		_w6927_
	);
	LUT2 #(
		.INIT('h2)
	) name6396 (
		_w5631_,
		_w6927_,
		_w6928_
	);
	LUT2 #(
		.INIT('h4)
	) name6397 (
		_w5631_,
		_w6927_,
		_w6929_
	);
	LUT2 #(
		.INIT('h1)
	) name6398 (
		_w6928_,
		_w6929_,
		_w6930_
	);
	LUT2 #(
		.INIT('h8)
	) name6399 (
		_w6395_,
		_w6930_,
		_w6931_
	);
	LUT2 #(
		.INIT('h1)
	) name6400 (
		_w6395_,
		_w6930_,
		_w6932_
	);
	LUT2 #(
		.INIT('h1)
	) name6401 (
		_w6931_,
		_w6932_,
		_w6933_
	);
	LUT2 #(
		.INIT('h1)
	) name6402 (
		_w6848_,
		_w6933_,
		_w6934_
	);
	LUT2 #(
		.INIT('h8)
	) name6403 (
		_w6848_,
		_w6933_,
		_w6935_
	);
	LUT2 #(
		.INIT('h1)
	) name6404 (
		\ld_r_reg/P0001 ,
		_w6934_,
		_w6936_
	);
	LUT2 #(
		.INIT('h4)
	) name6405 (
		_w6935_,
		_w6936_,
		_w6937_
	);
	LUT2 #(
		.INIT('h1)
	) name6406 (
		\text_in_r_reg[41]/P0001 ,
		\u0_w_reg[2][9]/P0001 ,
		_w6938_
	);
	LUT2 #(
		.INIT('h8)
	) name6407 (
		\text_in_r_reg[41]/P0001 ,
		\u0_w_reg[2][9]/P0001 ,
		_w6939_
	);
	LUT2 #(
		.INIT('h2)
	) name6408 (
		\ld_r_reg/P0001 ,
		_w6938_,
		_w6940_
	);
	LUT2 #(
		.INIT('h4)
	) name6409 (
		_w6939_,
		_w6940_,
		_w6941_
	);
	LUT2 #(
		.INIT('h1)
	) name6410 (
		_w6937_,
		_w6941_,
		_w6942_
	);
	LUT2 #(
		.INIT('h1)
	) name6411 (
		_w1145_,
		_w5830_,
		_w6943_
	);
	LUT2 #(
		.INIT('h8)
	) name6412 (
		_w1145_,
		_w5830_,
		_w6944_
	);
	LUT2 #(
		.INIT('h1)
	) name6413 (
		_w6943_,
		_w6944_,
		_w6945_
	);
	LUT2 #(
		.INIT('h2)
	) name6414 (
		\u0_w_reg[2][5]/P0001 ,
		_w6180_,
		_w6946_
	);
	LUT2 #(
		.INIT('h4)
	) name6415 (
		\u0_w_reg[2][5]/P0001 ,
		_w6180_,
		_w6947_
	);
	LUT2 #(
		.INIT('h1)
	) name6416 (
		_w6946_,
		_w6947_,
		_w6948_
	);
	LUT2 #(
		.INIT('h8)
	) name6417 (
		_w5931_,
		_w6948_,
		_w6949_
	);
	LUT2 #(
		.INIT('h1)
	) name6418 (
		_w5931_,
		_w6948_,
		_w6950_
	);
	LUT2 #(
		.INIT('h1)
	) name6419 (
		_w6949_,
		_w6950_,
		_w6951_
	);
	LUT2 #(
		.INIT('h1)
	) name6420 (
		_w6945_,
		_w6951_,
		_w6952_
	);
	LUT2 #(
		.INIT('h8)
	) name6421 (
		_w6945_,
		_w6951_,
		_w6953_
	);
	LUT2 #(
		.INIT('h1)
	) name6422 (
		\ld_r_reg/P0001 ,
		_w6952_,
		_w6954_
	);
	LUT2 #(
		.INIT('h4)
	) name6423 (
		_w6953_,
		_w6954_,
		_w6955_
	);
	LUT2 #(
		.INIT('h1)
	) name6424 (
		\text_in_r_reg[37]/P0001 ,
		\u0_w_reg[2][5]/P0001 ,
		_w6956_
	);
	LUT2 #(
		.INIT('h8)
	) name6425 (
		\text_in_r_reg[37]/P0001 ,
		\u0_w_reg[2][5]/P0001 ,
		_w6957_
	);
	LUT2 #(
		.INIT('h2)
	) name6426 (
		\ld_r_reg/P0001 ,
		_w6956_,
		_w6958_
	);
	LUT2 #(
		.INIT('h4)
	) name6427 (
		_w6957_,
		_w6958_,
		_w6959_
	);
	LUT2 #(
		.INIT('h1)
	) name6428 (
		_w6955_,
		_w6959_,
		_w6960_
	);
	LUT2 #(
		.INIT('h2)
	) name6429 (
		\u0_w_reg[2][28]/P0001 ,
		_w6180_,
		_w6961_
	);
	LUT2 #(
		.INIT('h4)
	) name6430 (
		\u0_w_reg[2][28]/P0001 ,
		_w6180_,
		_w6962_
	);
	LUT2 #(
		.INIT('h1)
	) name6431 (
		_w6961_,
		_w6962_,
		_w6963_
	);
	LUT2 #(
		.INIT('h8)
	) name6432 (
		_w6058_,
		_w6963_,
		_w6964_
	);
	LUT2 #(
		.INIT('h1)
	) name6433 (
		_w6058_,
		_w6963_,
		_w6965_
	);
	LUT2 #(
		.INIT('h1)
	) name6434 (
		_w6964_,
		_w6965_,
		_w6966_
	);
	LUT2 #(
		.INIT('h4)
	) name6435 (
		\sa02_reg[2]/P0001 ,
		_w1043_,
		_w6967_
	);
	LUT2 #(
		.INIT('h1)
	) name6436 (
		_w996_,
		_w5141_,
		_w6968_
	);
	LUT2 #(
		.INIT('h2)
	) name6437 (
		\sa02_reg[2]/P0001 ,
		_w6968_,
		_w6969_
	);
	LUT2 #(
		.INIT('h1)
	) name6438 (
		_w977_,
		_w5787_,
		_w6970_
	);
	LUT2 #(
		.INIT('h4)
	) name6439 (
		_w6337_,
		_w6970_,
		_w6971_
	);
	LUT2 #(
		.INIT('h4)
	) name6440 (
		_w6967_,
		_w6971_,
		_w6972_
	);
	LUT2 #(
		.INIT('h4)
	) name6441 (
		_w6969_,
		_w6972_,
		_w6973_
	);
	LUT2 #(
		.INIT('h2)
	) name6442 (
		\sa02_reg[1]/P0001 ,
		_w6973_,
		_w6974_
	);
	LUT2 #(
		.INIT('h2)
	) name6443 (
		_w1006_,
		_w1017_,
		_w6975_
	);
	LUT2 #(
		.INIT('h8)
	) name6444 (
		_w974_,
		_w1003_,
		_w6976_
	);
	LUT2 #(
		.INIT('h8)
	) name6445 (
		\sa02_reg[7]/NET0131 ,
		_w978_,
		_w6977_
	);
	LUT2 #(
		.INIT('h4)
	) name6446 (
		_w982_,
		_w6977_,
		_w6978_
	);
	LUT2 #(
		.INIT('h1)
	) name6447 (
		_w5182_,
		_w6976_,
		_w6979_
	);
	LUT2 #(
		.INIT('h1)
	) name6448 (
		_w6975_,
		_w6978_,
		_w6980_
	);
	LUT2 #(
		.INIT('h8)
	) name6449 (
		_w6979_,
		_w6980_,
		_w6981_
	);
	LUT2 #(
		.INIT('h1)
	) name6450 (
		\sa02_reg[1]/P0001 ,
		_w6981_,
		_w6982_
	);
	LUT2 #(
		.INIT('h1)
	) name6451 (
		\sa02_reg[2]/P0001 ,
		_w5080_,
		_w6983_
	);
	LUT2 #(
		.INIT('h8)
	) name6452 (
		_w984_,
		_w996_,
		_w6984_
	);
	LUT2 #(
		.INIT('h1)
	) name6453 (
		_w1073_,
		_w5173_,
		_w6985_
	);
	LUT2 #(
		.INIT('h4)
	) name6454 (
		_w6984_,
		_w6985_,
		_w6986_
	);
	LUT2 #(
		.INIT('h4)
	) name6455 (
		_w6983_,
		_w6986_,
		_w6987_
	);
	LUT2 #(
		.INIT('h4)
	) name6456 (
		_w6982_,
		_w6987_,
		_w6988_
	);
	LUT2 #(
		.INIT('h4)
	) name6457 (
		_w6974_,
		_w6988_,
		_w6989_
	);
	LUT2 #(
		.INIT('h1)
	) name6458 (
		\sa02_reg[0]/P0001 ,
		_w6989_,
		_w6990_
	);
	LUT2 #(
		.INIT('h1)
	) name6459 (
		_w1021_,
		_w6364_,
		_w6991_
	);
	LUT2 #(
		.INIT('h1)
	) name6460 (
		\sa02_reg[2]/P0001 ,
		_w6991_,
		_w6992_
	);
	LUT2 #(
		.INIT('h4)
	) name6461 (
		_w5159_,
		_w5753_,
		_w6993_
	);
	LUT2 #(
		.INIT('h1)
	) name6462 (
		_w1121_,
		_w5171_,
		_w6994_
	);
	LUT2 #(
		.INIT('h4)
	) name6463 (
		_w5098_,
		_w6994_,
		_w6995_
	);
	LUT2 #(
		.INIT('h1)
	) name6464 (
		_w6377_,
		_w6993_,
		_w6996_
	);
	LUT2 #(
		.INIT('h8)
	) name6465 (
		_w6995_,
		_w6996_,
		_w6997_
	);
	LUT2 #(
		.INIT('h4)
	) name6466 (
		_w6992_,
		_w6997_,
		_w6998_
	);
	LUT2 #(
		.INIT('h1)
	) name6467 (
		\sa02_reg[1]/P0001 ,
		_w6998_,
		_w6999_
	);
	LUT2 #(
		.INIT('h1)
	) name6468 (
		_w1042_,
		_w1062_,
		_w7000_
	);
	LUT2 #(
		.INIT('h4)
	) name6469 (
		_w5755_,
		_w7000_,
		_w7001_
	);
	LUT2 #(
		.INIT('h2)
	) name6470 (
		\sa02_reg[2]/P0001 ,
		_w7001_,
		_w7002_
	);
	LUT2 #(
		.INIT('h2)
	) name6471 (
		_w994_,
		_w1068_,
		_w7003_
	);
	LUT2 #(
		.INIT('h8)
	) name6472 (
		_w1025_,
		_w5108_,
		_w7004_
	);
	LUT2 #(
		.INIT('h1)
	) name6473 (
		_w5792_,
		_w7004_,
		_w7005_
	);
	LUT2 #(
		.INIT('h4)
	) name6474 (
		_w5119_,
		_w7005_,
		_w7006_
	);
	LUT2 #(
		.INIT('h4)
	) name6475 (
		_w7003_,
		_w7006_,
		_w7007_
	);
	LUT2 #(
		.INIT('h4)
	) name6476 (
		_w7002_,
		_w7007_,
		_w7008_
	);
	LUT2 #(
		.INIT('h2)
	) name6477 (
		\sa02_reg[1]/P0001 ,
		_w7008_,
		_w7009_
	);
	LUT2 #(
		.INIT('h2)
	) name6478 (
		_w6419_,
		_w6976_,
		_w7010_
	);
	LUT2 #(
		.INIT('h1)
	) name6479 (
		\sa02_reg[2]/P0001 ,
		_w7010_,
		_w7011_
	);
	LUT2 #(
		.INIT('h4)
	) name6480 (
		_w1024_,
		_w1131_,
		_w7012_
	);
	LUT2 #(
		.INIT('h2)
	) name6481 (
		_w1128_,
		_w7012_,
		_w7013_
	);
	LUT2 #(
		.INIT('h1)
	) name6482 (
		_w1070_,
		_w7013_,
		_w7014_
	);
	LUT2 #(
		.INIT('h4)
	) name6483 (
		_w7011_,
		_w7014_,
		_w7015_
	);
	LUT2 #(
		.INIT('h4)
	) name6484 (
		_w6999_,
		_w7015_,
		_w7016_
	);
	LUT2 #(
		.INIT('h4)
	) name6485 (
		_w7009_,
		_w7016_,
		_w7017_
	);
	LUT2 #(
		.INIT('h2)
	) name6486 (
		\sa02_reg[0]/P0001 ,
		_w7017_,
		_w7018_
	);
	LUT2 #(
		.INIT('h4)
	) name6487 (
		\sa02_reg[2]/P0001 ,
		_w5818_,
		_w7019_
	);
	LUT2 #(
		.INIT('h1)
	) name6488 (
		_w5323_,
		_w5767_,
		_w7020_
	);
	LUT2 #(
		.INIT('h4)
	) name6489 (
		_w1043_,
		_w7020_,
		_w7021_
	);
	LUT2 #(
		.INIT('h2)
	) name6490 (
		_w5108_,
		_w7021_,
		_w7022_
	);
	LUT2 #(
		.INIT('h1)
	) name6491 (
		_w5775_,
		_w7019_,
		_w7023_
	);
	LUT2 #(
		.INIT('h4)
	) name6492 (
		_w7022_,
		_w7023_,
		_w7024_
	);
	LUT2 #(
		.INIT('h2)
	) name6493 (
		\sa02_reg[1]/P0001 ,
		_w7024_,
		_w7025_
	);
	LUT2 #(
		.INIT('h1)
	) name6494 (
		_w1061_,
		_w1073_,
		_w7026_
	);
	LUT2 #(
		.INIT('h2)
	) name6495 (
		_w5106_,
		_w7026_,
		_w7027_
	);
	LUT2 #(
		.INIT('h8)
	) name6496 (
		\sa02_reg[6]/NET0131 ,
		_w1078_,
		_w7028_
	);
	LUT2 #(
		.INIT('h1)
	) name6497 (
		_w5792_,
		_w7028_,
		_w7029_
	);
	LUT2 #(
		.INIT('h2)
	) name6498 (
		_w5154_,
		_w7029_,
		_w7030_
	);
	LUT2 #(
		.INIT('h8)
	) name6499 (
		_w5780_,
		_w6363_,
		_w7031_
	);
	LUT2 #(
		.INIT('h1)
	) name6500 (
		_w1005_,
		_w5768_,
		_w7032_
	);
	LUT2 #(
		.INIT('h2)
	) name6501 (
		_w984_,
		_w7032_,
		_w7033_
	);
	LUT2 #(
		.INIT('h1)
	) name6502 (
		_w6305_,
		_w7031_,
		_w7034_
	);
	LUT2 #(
		.INIT('h4)
	) name6503 (
		_w7033_,
		_w7034_,
		_w7035_
	);
	LUT2 #(
		.INIT('h4)
	) name6504 (
		_w7027_,
		_w7035_,
		_w7036_
	);
	LUT2 #(
		.INIT('h4)
	) name6505 (
		_w7030_,
		_w7036_,
		_w7037_
	);
	LUT2 #(
		.INIT('h4)
	) name6506 (
		_w7025_,
		_w7037_,
		_w7038_
	);
	LUT2 #(
		.INIT('h4)
	) name6507 (
		_w6990_,
		_w7038_,
		_w7039_
	);
	LUT2 #(
		.INIT('h4)
	) name6508 (
		_w7018_,
		_w7039_,
		_w7040_
	);
	LUT2 #(
		.INIT('h8)
	) name6509 (
		_w532_,
		_w5459_,
		_w7041_
	);
	LUT2 #(
		.INIT('h1)
	) name6510 (
		_w604_,
		_w638_,
		_w7042_
	);
	LUT2 #(
		.INIT('h2)
	) name6511 (
		\sa13_reg[2]/P0001 ,
		_w7042_,
		_w7043_
	);
	LUT2 #(
		.INIT('h1)
	) name6512 (
		_w551_,
		_w5699_,
		_w7044_
	);
	LUT2 #(
		.INIT('h1)
	) name6513 (
		_w6243_,
		_w7041_,
		_w7045_
	);
	LUT2 #(
		.INIT('h8)
	) name6514 (
		_w7044_,
		_w7045_,
		_w7046_
	);
	LUT2 #(
		.INIT('h4)
	) name6515 (
		_w7043_,
		_w7046_,
		_w7047_
	);
	LUT2 #(
		.INIT('h2)
	) name6516 (
		\sa13_reg[1]/P0001 ,
		_w7047_,
		_w7048_
	);
	LUT2 #(
		.INIT('h1)
	) name6517 (
		\sa13_reg[2]/P0001 ,
		_w546_,
		_w7049_
	);
	LUT2 #(
		.INIT('h8)
	) name6518 (
		_w591_,
		_w653_,
		_w7050_
	);
	LUT2 #(
		.INIT('h2)
	) name6519 (
		\sa13_reg[7]/NET0131 ,
		_w547_,
		_w7051_
	);
	LUT2 #(
		.INIT('h8)
	) name6520 (
		_w603_,
		_w7051_,
		_w7052_
	);
	LUT2 #(
		.INIT('h8)
	) name6521 (
		_w556_,
		_w6281_,
		_w7053_
	);
	LUT2 #(
		.INIT('h1)
	) name6522 (
		_w5426_,
		_w7053_,
		_w7054_
	);
	LUT2 #(
		.INIT('h4)
	) name6523 (
		_w652_,
		_w7054_,
		_w7055_
	);
	LUT2 #(
		.INIT('h1)
	) name6524 (
		_w679_,
		_w7052_,
		_w7056_
	);
	LUT2 #(
		.INIT('h8)
	) name6525 (
		_w7055_,
		_w7056_,
		_w7057_
	);
	LUT2 #(
		.INIT('h1)
	) name6526 (
		\sa13_reg[1]/P0001 ,
		_w7057_,
		_w7058_
	);
	LUT2 #(
		.INIT('h1)
	) name6527 (
		_w671_,
		_w5464_,
		_w7059_
	);
	LUT2 #(
		.INIT('h4)
	) name6528 (
		_w7050_,
		_w7059_,
		_w7060_
	);
	LUT2 #(
		.INIT('h4)
	) name6529 (
		_w7049_,
		_w7060_,
		_w7061_
	);
	LUT2 #(
		.INIT('h4)
	) name6530 (
		_w7058_,
		_w7061_,
		_w7062_
	);
	LUT2 #(
		.INIT('h4)
	) name6531 (
		_w7048_,
		_w7062_,
		_w7063_
	);
	LUT2 #(
		.INIT('h1)
	) name6532 (
		\sa13_reg[0]/P0001 ,
		_w7063_,
		_w7064_
	);
	LUT2 #(
		.INIT('h4)
	) name6533 (
		_w901_,
		_w926_,
		_w7065_
	);
	LUT2 #(
		.INIT('h2)
	) name6534 (
		\sa13_reg[2]/P0001 ,
		_w7065_,
		_w7066_
	);
	LUT2 #(
		.INIT('h1)
	) name6535 (
		_w648_,
		_w856_,
		_w7067_
	);
	LUT2 #(
		.INIT('h1)
	) name6536 (
		\sa13_reg[2]/P0001 ,
		_w7067_,
		_w7068_
	);
	LUT2 #(
		.INIT('h1)
	) name6537 (
		_w654_,
		_w668_,
		_w7069_
	);
	LUT2 #(
		.INIT('h4)
	) name6538 (
		_w5682_,
		_w7069_,
		_w7070_
	);
	LUT2 #(
		.INIT('h4)
	) name6539 (
		_w7066_,
		_w7070_,
		_w7071_
	);
	LUT2 #(
		.INIT('h4)
	) name6540 (
		_w7068_,
		_w7071_,
		_w7072_
	);
	LUT2 #(
		.INIT('h1)
	) name6541 (
		\sa13_reg[1]/P0001 ,
		_w7072_,
		_w7073_
	);
	LUT2 #(
		.INIT('h1)
	) name6542 (
		_w568_,
		_w920_,
		_w7074_
	);
	LUT2 #(
		.INIT('h4)
	) name6543 (
		_w5456_,
		_w7074_,
		_w7075_
	);
	LUT2 #(
		.INIT('h2)
	) name6544 (
		\sa13_reg[2]/P0001 ,
		_w7075_,
		_w7076_
	);
	LUT2 #(
		.INIT('h1)
	) name6545 (
		_w588_,
		_w5425_,
		_w7077_
	);
	LUT2 #(
		.INIT('h1)
	) name6546 (
		_w5504_,
		_w5671_,
		_w7078_
	);
	LUT2 #(
		.INIT('h4)
	) name6547 (
		_w6284_,
		_w7078_,
		_w7079_
	);
	LUT2 #(
		.INIT('h8)
	) name6548 (
		_w7077_,
		_w7079_,
		_w7080_
	);
	LUT2 #(
		.INIT('h4)
	) name6549 (
		_w7076_,
		_w7080_,
		_w7081_
	);
	LUT2 #(
		.INIT('h2)
	) name6550 (
		\sa13_reg[1]/P0001 ,
		_w7081_,
		_w7082_
	);
	LUT2 #(
		.INIT('h8)
	) name6551 (
		\sa13_reg[3]/P0001 ,
		_w540_,
		_w7083_
	);
	LUT2 #(
		.INIT('h1)
	) name6552 (
		_w921_,
		_w7083_,
		_w7084_
	);
	LUT2 #(
		.INIT('h4)
	) name6553 (
		_w5426_,
		_w7084_,
		_w7085_
	);
	LUT2 #(
		.INIT('h1)
	) name6554 (
		\sa13_reg[2]/P0001 ,
		_w7085_,
		_w7086_
	);
	LUT2 #(
		.INIT('h1)
	) name6555 (
		_w864_,
		_w944_,
		_w7087_
	);
	LUT2 #(
		.INIT('h2)
	) name6556 (
		_w6281_,
		_w7087_,
		_w7088_
	);
	LUT2 #(
		.INIT('h1)
	) name6557 (
		_w911_,
		_w7088_,
		_w7089_
	);
	LUT2 #(
		.INIT('h4)
	) name6558 (
		_w7086_,
		_w7089_,
		_w7090_
	);
	LUT2 #(
		.INIT('h4)
	) name6559 (
		_w7082_,
		_w7090_,
		_w7091_
	);
	LUT2 #(
		.INIT('h4)
	) name6560 (
		_w7073_,
		_w7091_,
		_w7092_
	);
	LUT2 #(
		.INIT('h2)
	) name6561 (
		\sa13_reg[0]/P0001 ,
		_w7092_,
		_w7093_
	);
	LUT2 #(
		.INIT('h8)
	) name6562 (
		_w571_,
		_w623_,
		_w7094_
	);
	LUT2 #(
		.INIT('h1)
	) name6563 (
		_w632_,
		_w865_,
		_w7095_
	);
	LUT2 #(
		.INIT('h4)
	) name6564 (
		_w569_,
		_w7095_,
		_w7096_
	);
	LUT2 #(
		.INIT('h2)
	) name6565 (
		_w5424_,
		_w7096_,
		_w7097_
	);
	LUT2 #(
		.INIT('h8)
	) name6566 (
		_w955_,
		_w5459_,
		_w7098_
	);
	LUT2 #(
		.INIT('h1)
	) name6567 (
		_w5647_,
		_w7098_,
		_w7099_
	);
	LUT2 #(
		.INIT('h4)
	) name6568 (
		_w7097_,
		_w7099_,
		_w7100_
	);
	LUT2 #(
		.INIT('h2)
	) name6569 (
		\sa13_reg[1]/P0001 ,
		_w7100_,
		_w7101_
	);
	LUT2 #(
		.INIT('h1)
	) name6570 (
		_w918_,
		_w7050_,
		_w7102_
	);
	LUT2 #(
		.INIT('h2)
	) name6571 (
		_w6272_,
		_w7102_,
		_w7103_
	);
	LUT2 #(
		.INIT('h8)
	) name6572 (
		\sa13_reg[6]/NET0131 ,
		_w656_,
		_w7104_
	);
	LUT2 #(
		.INIT('h1)
	) name6573 (
		_w5671_,
		_w7104_,
		_w7105_
	);
	LUT2 #(
		.INIT('h2)
	) name6574 (
		_w6286_,
		_w7105_,
		_w7106_
	);
	LUT2 #(
		.INIT('h8)
	) name6575 (
		_w962_,
		_w5651_,
		_w7107_
	);
	LUT2 #(
		.INIT('h1)
	) name6576 (
		_w649_,
		_w6282_,
		_w7108_
	);
	LUT2 #(
		.INIT('h4)
	) name6577 (
		_w7094_,
		_w7108_,
		_w7109_
	);
	LUT2 #(
		.INIT('h4)
	) name6578 (
		_w7107_,
		_w7109_,
		_w7110_
	);
	LUT2 #(
		.INIT('h4)
	) name6579 (
		_w7106_,
		_w7110_,
		_w7111_
	);
	LUT2 #(
		.INIT('h4)
	) name6580 (
		_w7103_,
		_w7111_,
		_w7112_
	);
	LUT2 #(
		.INIT('h4)
	) name6581 (
		_w7101_,
		_w7112_,
		_w7113_
	);
	LUT2 #(
		.INIT('h4)
	) name6582 (
		_w7064_,
		_w7113_,
		_w7114_
	);
	LUT2 #(
		.INIT('h4)
	) name6583 (
		_w7093_,
		_w7114_,
		_w7115_
	);
	LUT2 #(
		.INIT('h2)
	) name6584 (
		_w7040_,
		_w7115_,
		_w7116_
	);
	LUT2 #(
		.INIT('h4)
	) name6585 (
		_w7040_,
		_w7115_,
		_w7117_
	);
	LUT2 #(
		.INIT('h1)
	) name6586 (
		_w7116_,
		_w7117_,
		_w7118_
	);
	LUT2 #(
		.INIT('h4)
	) name6587 (
		_w5519_,
		_w7118_,
		_w7119_
	);
	LUT2 #(
		.INIT('h2)
	) name6588 (
		_w5519_,
		_w7118_,
		_w7120_
	);
	LUT2 #(
		.INIT('h1)
	) name6589 (
		_w7119_,
		_w7120_,
		_w7121_
	);
	LUT2 #(
		.INIT('h2)
	) name6590 (
		_w6966_,
		_w7121_,
		_w7122_
	);
	LUT2 #(
		.INIT('h4)
	) name6591 (
		_w6966_,
		_w7121_,
		_w7123_
	);
	LUT2 #(
		.INIT('h1)
	) name6592 (
		\ld_r_reg/P0001 ,
		_w7122_,
		_w7124_
	);
	LUT2 #(
		.INIT('h4)
	) name6593 (
		_w7123_,
		_w7124_,
		_w7125_
	);
	LUT2 #(
		.INIT('h2)
	) name6594 (
		\text_in_r_reg[60]/P0001 ,
		\u0_w_reg[2][28]/P0001 ,
		_w7126_
	);
	LUT2 #(
		.INIT('h4)
	) name6595 (
		\text_in_r_reg[60]/P0001 ,
		\u0_w_reg[2][28]/P0001 ,
		_w7127_
	);
	LUT2 #(
		.INIT('h2)
	) name6596 (
		\ld_r_reg/P0001 ,
		_w7126_,
		_w7128_
	);
	LUT2 #(
		.INIT('h4)
	) name6597 (
		_w7127_,
		_w7128_,
		_w7129_
	);
	LUT2 #(
		.INIT('h1)
	) name6598 (
		_w7125_,
		_w7129_,
		_w7130_
	);
	LUT2 #(
		.INIT('h4)
	) name6599 (
		_w5530_,
		_w6880_,
		_w7131_
	);
	LUT2 #(
		.INIT('h1)
	) name6600 (
		\sa20_reg[2]/P0001 ,
		_w7131_,
		_w7132_
	);
	LUT2 #(
		.INIT('h1)
	) name6601 (
		_w820_,
		_w5527_,
		_w7133_
	);
	LUT2 #(
		.INIT('h1)
	) name6602 (
		\sa20_reg[2]/P0001 ,
		_w7133_,
		_w7134_
	);
	LUT2 #(
		.INIT('h1)
	) name6603 (
		_w715_,
		_w795_,
		_w7135_
	);
	LUT2 #(
		.INIT('h4)
	) name6604 (
		_w5617_,
		_w7135_,
		_w7136_
	);
	LUT2 #(
		.INIT('h4)
	) name6605 (
		_w7134_,
		_w7136_,
		_w7137_
	);
	LUT2 #(
		.INIT('h2)
	) name6606 (
		\sa20_reg[1]/P0001 ,
		_w7137_,
		_w7138_
	);
	LUT2 #(
		.INIT('h1)
	) name6607 (
		_w737_,
		_w5591_,
		_w7139_
	);
	LUT2 #(
		.INIT('h1)
	) name6608 (
		\sa20_reg[2]/P0001 ,
		_w7139_,
		_w7140_
	);
	LUT2 #(
		.INIT('h1)
	) name6609 (
		_w694_,
		_w701_,
		_w7141_
	);
	LUT2 #(
		.INIT('h2)
	) name6610 (
		_w5984_,
		_w7141_,
		_w7142_
	);
	LUT2 #(
		.INIT('h1)
	) name6611 (
		_w809_,
		_w838_,
		_w7143_
	);
	LUT2 #(
		.INIT('h4)
	) name6612 (
		_w6036_,
		_w7143_,
		_w7144_
	);
	LUT2 #(
		.INIT('h1)
	) name6613 (
		_w6917_,
		_w7142_,
		_w7145_
	);
	LUT2 #(
		.INIT('h8)
	) name6614 (
		_w7144_,
		_w7145_,
		_w7146_
	);
	LUT2 #(
		.INIT('h4)
	) name6615 (
		_w7140_,
		_w7146_,
		_w7147_
	);
	LUT2 #(
		.INIT('h1)
	) name6616 (
		\sa20_reg[1]/P0001 ,
		_w7147_,
		_w7148_
	);
	LUT2 #(
		.INIT('h8)
	) name6617 (
		\sa20_reg[3]/P0001 ,
		_w705_,
		_w7149_
	);
	LUT2 #(
		.INIT('h2)
	) name6618 (
		_w5920_,
		_w7149_,
		_w7150_
	);
	LUT2 #(
		.INIT('h2)
	) name6619 (
		\sa20_reg[4]/P0001 ,
		_w7150_,
		_w7151_
	);
	LUT2 #(
		.INIT('h1)
	) name6620 (
		_w5585_,
		_w5979_,
		_w7152_
	);
	LUT2 #(
		.INIT('h4)
	) name6621 (
		_w6715_,
		_w7152_,
		_w7153_
	);
	LUT2 #(
		.INIT('h2)
	) name6622 (
		\sa20_reg[1]/P0001 ,
		_w7153_,
		_w7154_
	);
	LUT2 #(
		.INIT('h1)
	) name6623 (
		_w7151_,
		_w7154_,
		_w7155_
	);
	LUT2 #(
		.INIT('h2)
	) name6624 (
		\sa20_reg[2]/P0001 ,
		_w7155_,
		_w7156_
	);
	LUT2 #(
		.INIT('h1)
	) name6625 (
		_w5901_,
		_w7132_,
		_w7157_
	);
	LUT2 #(
		.INIT('h4)
	) name6626 (
		_w7138_,
		_w7157_,
		_w7158_
	);
	LUT2 #(
		.INIT('h1)
	) name6627 (
		_w7148_,
		_w7156_,
		_w7159_
	);
	LUT2 #(
		.INIT('h8)
	) name6628 (
		_w7158_,
		_w7159_,
		_w7160_
	);
	LUT2 #(
		.INIT('h2)
	) name6629 (
		\sa20_reg[0]/P0001 ,
		_w7160_,
		_w7161_
	);
	LUT2 #(
		.INIT('h1)
	) name6630 (
		_w782_,
		_w790_,
		_w7162_
	);
	LUT2 #(
		.INIT('h2)
	) name6631 (
		\sa20_reg[2]/P0001 ,
		_w7162_,
		_w7163_
	);
	LUT2 #(
		.INIT('h4)
	) name6632 (
		\sa20_reg[2]/P0001 ,
		_w740_,
		_w7164_
	);
	LUT2 #(
		.INIT('h1)
	) name6633 (
		_w707_,
		_w5859_,
		_w7165_
	);
	LUT2 #(
		.INIT('h1)
	) name6634 (
		_w6689_,
		_w7164_,
		_w7166_
	);
	LUT2 #(
		.INIT('h8)
	) name6635 (
		_w7165_,
		_w7166_,
		_w7167_
	);
	LUT2 #(
		.INIT('h4)
	) name6636 (
		_w7163_,
		_w7167_,
		_w7168_
	);
	LUT2 #(
		.INIT('h2)
	) name6637 (
		\sa20_reg[1]/P0001 ,
		_w7168_,
		_w7169_
	);
	LUT2 #(
		.INIT('h4)
	) name6638 (
		\sa20_reg[2]/P0001 ,
		_w704_,
		_w7170_
	);
	LUT2 #(
		.INIT('h4)
	) name6639 (
		\sa20_reg[7]/NET0131 ,
		_w6849_,
		_w7171_
	);
	LUT2 #(
		.INIT('h2)
	) name6640 (
		_w828_,
		_w7171_,
		_w7172_
	);
	LUT2 #(
		.INIT('h1)
	) name6641 (
		_w7170_,
		_w7172_,
		_w7173_
	);
	LUT2 #(
		.INIT('h4)
	) name6642 (
		_w708_,
		_w736_,
		_w7174_
	);
	LUT2 #(
		.INIT('h1)
	) name6643 (
		_w807_,
		_w7174_,
		_w7175_
	);
	LUT2 #(
		.INIT('h2)
	) name6644 (
		\sa20_reg[2]/P0001 ,
		_w7175_,
		_w7176_
	);
	LUT2 #(
		.INIT('h1)
	) name6645 (
		_w808_,
		_w825_,
		_w7177_
	);
	LUT2 #(
		.INIT('h4)
	) name6646 (
		_w5530_,
		_w7177_,
		_w7178_
	);
	LUT2 #(
		.INIT('h4)
	) name6647 (
		_w7176_,
		_w7178_,
		_w7179_
	);
	LUT2 #(
		.INIT('h1)
	) name6648 (
		\sa20_reg[1]/P0001 ,
		_w7179_,
		_w7180_
	);
	LUT2 #(
		.INIT('h1)
	) name6649 (
		_w5878_,
		_w7173_,
		_w7181_
	);
	LUT2 #(
		.INIT('h4)
	) name6650 (
		_w7169_,
		_w7181_,
		_w7182_
	);
	LUT2 #(
		.INIT('h4)
	) name6651 (
		_w7180_,
		_w7182_,
		_w7183_
	);
	LUT2 #(
		.INIT('h1)
	) name6652 (
		\sa20_reg[0]/P0001 ,
		_w7183_,
		_w7184_
	);
	LUT2 #(
		.INIT('h8)
	) name6653 (
		_w763_,
		_w5981_,
		_w7185_
	);
	LUT2 #(
		.INIT('h1)
	) name6654 (
		_w694_,
		_w720_,
		_w7186_
	);
	LUT2 #(
		.INIT('h2)
	) name6655 (
		_w6894_,
		_w7186_,
		_w7187_
	);
	LUT2 #(
		.INIT('h1)
	) name6656 (
		_w740_,
		_w791_,
		_w7188_
	);
	LUT2 #(
		.INIT('h4)
	) name6657 (
		_w5997_,
		_w7188_,
		_w7189_
	);
	LUT2 #(
		.INIT('h2)
	) name6658 (
		_w747_,
		_w7189_,
		_w7190_
	);
	LUT2 #(
		.INIT('h1)
	) name6659 (
		_w6008_,
		_w7185_,
		_w7191_
	);
	LUT2 #(
		.INIT('h4)
	) name6660 (
		_w7187_,
		_w7191_,
		_w7192_
	);
	LUT2 #(
		.INIT('h4)
	) name6661 (
		_w7190_,
		_w7192_,
		_w7193_
	);
	LUT2 #(
		.INIT('h2)
	) name6662 (
		\sa20_reg[1]/P0001 ,
		_w7193_,
		_w7194_
	);
	LUT2 #(
		.INIT('h1)
	) name6663 (
		_w721_,
		_w5998_,
		_w7195_
	);
	LUT2 #(
		.INIT('h2)
	) name6664 (
		_w761_,
		_w7195_,
		_w7196_
	);
	LUT2 #(
		.INIT('h1)
	) name6665 (
		\sa20_reg[2]/P0001 ,
		_w6005_,
		_w7197_
	);
	LUT2 #(
		.INIT('h2)
	) name6666 (
		\sa20_reg[2]/P0001 ,
		_w5878_,
		_w7198_
	);
	LUT2 #(
		.INIT('h4)
	) name6667 (
		_w5894_,
		_w7198_,
		_w7199_
	);
	LUT2 #(
		.INIT('h1)
	) name6668 (
		\sa20_reg[1]/P0001 ,
		_w7197_,
		_w7200_
	);
	LUT2 #(
		.INIT('h4)
	) name6669 (
		_w7199_,
		_w7200_,
		_w7201_
	);
	LUT2 #(
		.INIT('h1)
	) name6670 (
		_w822_,
		_w7196_,
		_w7202_
	);
	LUT2 #(
		.INIT('h4)
	) name6671 (
		_w7201_,
		_w7202_,
		_w7203_
	);
	LUT2 #(
		.INIT('h4)
	) name6672 (
		_w7194_,
		_w7203_,
		_w7204_
	);
	LUT2 #(
		.INIT('h4)
	) name6673 (
		_w7161_,
		_w7204_,
		_w7205_
	);
	LUT2 #(
		.INIT('h4)
	) name6674 (
		_w7184_,
		_w7205_,
		_w7206_
	);
	LUT2 #(
		.INIT('h2)
	) name6675 (
		_w7115_,
		_w7206_,
		_w7207_
	);
	LUT2 #(
		.INIT('h4)
	) name6676 (
		_w7115_,
		_w7206_,
		_w7208_
	);
	LUT2 #(
		.INIT('h1)
	) name6677 (
		_w7207_,
		_w7208_,
		_w7209_
	);
	LUT2 #(
		.INIT('h2)
	) name6678 (
		_w5516_,
		_w5830_,
		_w7210_
	);
	LUT2 #(
		.INIT('h4)
	) name6679 (
		_w5516_,
		_w5830_,
		_w7211_
	);
	LUT2 #(
		.INIT('h1)
	) name6680 (
		_w7210_,
		_w7211_,
		_w7212_
	);
	LUT2 #(
		.INIT('h8)
	) name6681 (
		_w7209_,
		_w7212_,
		_w7213_
	);
	LUT2 #(
		.INIT('h1)
	) name6682 (
		_w7209_,
		_w7212_,
		_w7214_
	);
	LUT2 #(
		.INIT('h1)
	) name6683 (
		_w7213_,
		_w7214_,
		_w7215_
	);
	LUT2 #(
		.INIT('h1)
	) name6684 (
		_w5631_,
		_w6055_,
		_w7216_
	);
	LUT2 #(
		.INIT('h8)
	) name6685 (
		_w5631_,
		_w6055_,
		_w7217_
	);
	LUT2 #(
		.INIT('h1)
	) name6686 (
		_w7216_,
		_w7217_,
		_w7218_
	);
	LUT2 #(
		.INIT('h2)
	) name6687 (
		\u0_w_reg[2][20]/P0001 ,
		_w6180_,
		_w7219_
	);
	LUT2 #(
		.INIT('h4)
	) name6688 (
		\u0_w_reg[2][20]/P0001 ,
		_w6180_,
		_w7220_
	);
	LUT2 #(
		.INIT('h1)
	) name6689 (
		_w7219_,
		_w7220_,
		_w7221_
	);
	LUT2 #(
		.INIT('h8)
	) name6690 (
		_w7218_,
		_w7221_,
		_w7222_
	);
	LUT2 #(
		.INIT('h1)
	) name6691 (
		_w7218_,
		_w7221_,
		_w7223_
	);
	LUT2 #(
		.INIT('h1)
	) name6692 (
		_w7222_,
		_w7223_,
		_w7224_
	);
	LUT2 #(
		.INIT('h2)
	) name6693 (
		_w7215_,
		_w7224_,
		_w7225_
	);
	LUT2 #(
		.INIT('h4)
	) name6694 (
		_w7215_,
		_w7224_,
		_w7226_
	);
	LUT2 #(
		.INIT('h1)
	) name6695 (
		\ld_r_reg/P0001 ,
		_w7225_,
		_w7227_
	);
	LUT2 #(
		.INIT('h4)
	) name6696 (
		_w7226_,
		_w7227_,
		_w7228_
	);
	LUT2 #(
		.INIT('h2)
	) name6697 (
		\text_in_r_reg[52]/P0001 ,
		\u0_w_reg[2][20]/P0001 ,
		_w7229_
	);
	LUT2 #(
		.INIT('h4)
	) name6698 (
		\text_in_r_reg[52]/P0001 ,
		\u0_w_reg[2][20]/P0001 ,
		_w7230_
	);
	LUT2 #(
		.INIT('h2)
	) name6699 (
		\ld_r_reg/P0001 ,
		_w7229_,
		_w7231_
	);
	LUT2 #(
		.INIT('h4)
	) name6700 (
		_w7230_,
		_w7231_,
		_w7232_
	);
	LUT2 #(
		.INIT('h1)
	) name6701 (
		_w7228_,
		_w7232_,
		_w7233_
	);
	LUT2 #(
		.INIT('h1)
	) name6702 (
		_w6180_,
		_w6657_,
		_w7234_
	);
	LUT2 #(
		.INIT('h8)
	) name6703 (
		_w6180_,
		_w6657_,
		_w7235_
	);
	LUT2 #(
		.INIT('h1)
	) name6704 (
		_w7234_,
		_w7235_,
		_w7236_
	);
	LUT2 #(
		.INIT('h1)
	) name6705 (
		_w1217_,
		_w5206_,
		_w7237_
	);
	LUT2 #(
		.INIT('h1)
	) name6706 (
		\sa31_reg[2]/P0001 ,
		_w7237_,
		_w7238_
	);
	LUT2 #(
		.INIT('h1)
	) name6707 (
		_w1194_,
		_w5268_,
		_w7239_
	);
	LUT2 #(
		.INIT('h4)
	) name6708 (
		_w1207_,
		_w7239_,
		_w7240_
	);
	LUT2 #(
		.INIT('h2)
	) name6709 (
		\sa31_reg[2]/P0001 ,
		_w7240_,
		_w7241_
	);
	LUT2 #(
		.INIT('h1)
	) name6710 (
		_w1234_,
		_w1247_,
		_w7242_
	);
	LUT2 #(
		.INIT('h4)
	) name6711 (
		_w6832_,
		_w7242_,
		_w7243_
	);
	LUT2 #(
		.INIT('h4)
	) name6712 (
		_w7238_,
		_w7243_,
		_w7244_
	);
	LUT2 #(
		.INIT('h4)
	) name6713 (
		_w7241_,
		_w7244_,
		_w7245_
	);
	LUT2 #(
		.INIT('h1)
	) name6714 (
		\sa31_reg[1]/P0001 ,
		_w7245_,
		_w7246_
	);
	LUT2 #(
		.INIT('h8)
	) name6715 (
		\sa31_reg[4]/P0001 ,
		_w6515_,
		_w7247_
	);
	LUT2 #(
		.INIT('h2)
	) name6716 (
		_w1178_,
		_w1276_,
		_w7248_
	);
	LUT2 #(
		.INIT('h1)
	) name6717 (
		_w6092_,
		_w7248_,
		_w7249_
	);
	LUT2 #(
		.INIT('h2)
	) name6718 (
		\sa31_reg[2]/P0001 ,
		_w7249_,
		_w7250_
	);
	LUT2 #(
		.INIT('h1)
	) name6719 (
		_w1219_,
		_w6569_,
		_w7251_
	);
	LUT2 #(
		.INIT('h1)
	) name6720 (
		\sa31_reg[2]/P0001 ,
		_w7251_,
		_w7252_
	);
	LUT2 #(
		.INIT('h1)
	) name6721 (
		_w6119_,
		_w7247_,
		_w7253_
	);
	LUT2 #(
		.INIT('h4)
	) name6722 (
		_w7250_,
		_w7253_,
		_w7254_
	);
	LUT2 #(
		.INIT('h4)
	) name6723 (
		_w7252_,
		_w7254_,
		_w7255_
	);
	LUT2 #(
		.INIT('h2)
	) name6724 (
		\sa31_reg[1]/P0001 ,
		_w7255_,
		_w7256_
	);
	LUT2 #(
		.INIT('h8)
	) name6725 (
		_w1152_,
		_w1182_,
		_w7257_
	);
	LUT2 #(
		.INIT('h2)
	) name6726 (
		_w6529_,
		_w7257_,
		_w7258_
	);
	LUT2 #(
		.INIT('h1)
	) name6727 (
		\sa31_reg[2]/P0001 ,
		_w7258_,
		_w7259_
	);
	LUT2 #(
		.INIT('h4)
	) name6728 (
		_w1206_,
		_w5287_,
		_w7260_
	);
	LUT2 #(
		.INIT('h2)
	) name6729 (
		_w1215_,
		_w7260_,
		_w7261_
	);
	LUT2 #(
		.INIT('h1)
	) name6730 (
		_w5264_,
		_w7261_,
		_w7262_
	);
	LUT2 #(
		.INIT('h4)
	) name6731 (
		_w7259_,
		_w7262_,
		_w7263_
	);
	LUT2 #(
		.INIT('h4)
	) name6732 (
		_w7256_,
		_w7263_,
		_w7264_
	);
	LUT2 #(
		.INIT('h4)
	) name6733 (
		_w7246_,
		_w7264_,
		_w7265_
	);
	LUT2 #(
		.INIT('h2)
	) name6734 (
		\sa31_reg[0]/P0002 ,
		_w7265_,
		_w7266_
	);
	LUT2 #(
		.INIT('h8)
	) name6735 (
		_w1147_,
		_w6136_,
		_w7267_
	);
	LUT2 #(
		.INIT('h1)
	) name6736 (
		_w1204_,
		_w1261_,
		_w7268_
	);
	LUT2 #(
		.INIT('h2)
	) name6737 (
		\sa31_reg[2]/P0001 ,
		_w7268_,
		_w7269_
	);
	LUT2 #(
		.INIT('h1)
	) name6738 (
		_w1207_,
		_w6148_,
		_w7270_
	);
	LUT2 #(
		.INIT('h4)
	) name6739 (
		_w7267_,
		_w7270_,
		_w7271_
	);
	LUT2 #(
		.INIT('h4)
	) name6740 (
		_w6787_,
		_w7271_,
		_w7272_
	);
	LUT2 #(
		.INIT('h4)
	) name6741 (
		_w7269_,
		_w7272_,
		_w7273_
	);
	LUT2 #(
		.INIT('h2)
	) name6742 (
		\sa31_reg[1]/P0001 ,
		_w7273_,
		_w7274_
	);
	LUT2 #(
		.INIT('h8)
	) name6743 (
		_w1186_,
		_w1215_,
		_w7275_
	);
	LUT2 #(
		.INIT('h2)
	) name6744 (
		\sa31_reg[7]/P0001 ,
		_w1229_,
		_w7276_
	);
	LUT2 #(
		.INIT('h8)
	) name6745 (
		_w1279_,
		_w7276_,
		_w7277_
	);
	LUT2 #(
		.INIT('h1)
	) name6746 (
		_w7257_,
		_w7275_,
		_w7278_
	);
	LUT2 #(
		.INIT('h4)
	) name6747 (
		_w1233_,
		_w7278_,
		_w7279_
	);
	LUT2 #(
		.INIT('h4)
	) name6748 (
		_w7277_,
		_w7279_,
		_w7280_
	);
	LUT2 #(
		.INIT('h4)
	) name6749 (
		_w1223_,
		_w7280_,
		_w7281_
	);
	LUT2 #(
		.INIT('h1)
	) name6750 (
		\sa31_reg[1]/P0001 ,
		_w7281_,
		_w7282_
	);
	LUT2 #(
		.INIT('h1)
	) name6751 (
		\sa31_reg[2]/P0001 ,
		_w1203_,
		_w7283_
	);
	LUT2 #(
		.INIT('h8)
	) name6752 (
		_w1204_,
		_w1265_,
		_w7284_
	);
	LUT2 #(
		.INIT('h1)
	) name6753 (
		_w1245_,
		_w5258_,
		_w7285_
	);
	LUT2 #(
		.INIT('h4)
	) name6754 (
		_w7284_,
		_w7285_,
		_w7286_
	);
	LUT2 #(
		.INIT('h4)
	) name6755 (
		_w7283_,
		_w7286_,
		_w7287_
	);
	LUT2 #(
		.INIT('h4)
	) name6756 (
		_w7282_,
		_w7287_,
		_w7288_
	);
	LUT2 #(
		.INIT('h4)
	) name6757 (
		_w7274_,
		_w7288_,
		_w7289_
	);
	LUT2 #(
		.INIT('h1)
	) name6758 (
		\sa31_reg[0]/P0002 ,
		_w7289_,
		_w7290_
	);
	LUT2 #(
		.INIT('h1)
	) name6759 (
		_w5199_,
		_w6598_,
		_w7291_
	);
	LUT2 #(
		.INIT('h4)
	) name6760 (
		_w1148_,
		_w7291_,
		_w7292_
	);
	LUT2 #(
		.INIT('h2)
	) name6761 (
		_w1162_,
		_w7292_,
		_w7293_
	);
	LUT2 #(
		.INIT('h8)
	) name6762 (
		\sa31_reg[6]/NET0131 ,
		_w5263_,
		_w7294_
	);
	LUT2 #(
		.INIT('h1)
	) name6763 (
		_w6119_,
		_w7294_,
		_w7295_
	);
	LUT2 #(
		.INIT('h2)
	) name6764 (
		\sa31_reg[2]/P0001 ,
		_w7295_,
		_w7296_
	);
	LUT2 #(
		.INIT('h4)
	) name6765 (
		\sa31_reg[6]/NET0131 ,
		_w6584_,
		_w7297_
	);
	LUT2 #(
		.INIT('h1)
	) name6766 (
		_w6135_,
		_w7297_,
		_w7298_
	);
	LUT2 #(
		.INIT('h4)
	) name6767 (
		_w7293_,
		_w7298_,
		_w7299_
	);
	LUT2 #(
		.INIT('h4)
	) name6768 (
		_w7296_,
		_w7299_,
		_w7300_
	);
	LUT2 #(
		.INIT('h2)
	) name6769 (
		\sa31_reg[1]/P0001 ,
		_w7300_,
		_w7301_
	);
	LUT2 #(
		.INIT('h1)
	) name6770 (
		_w1233_,
		_w6110_,
		_w7302_
	);
	LUT2 #(
		.INIT('h2)
	) name6771 (
		_w1279_,
		_w7302_,
		_w7303_
	);
	LUT2 #(
		.INIT('h8)
	) name6772 (
		_w6136_,
		_w6790_,
		_w7304_
	);
	LUT2 #(
		.INIT('h1)
	) name6773 (
		_w7303_,
		_w7304_,
		_w7305_
	);
	LUT2 #(
		.INIT('h1)
	) name6774 (
		\sa31_reg[1]/P0001 ,
		_w7305_,
		_w7306_
	);
	LUT2 #(
		.INIT('h1)
	) name6775 (
		_w1183_,
		_w6124_,
		_w7307_
	);
	LUT2 #(
		.INIT('h2)
	) name6776 (
		_w1265_,
		_w7307_,
		_w7308_
	);
	LUT2 #(
		.INIT('h1)
	) name6777 (
		_w6769_,
		_w7308_,
		_w7309_
	);
	LUT2 #(
		.INIT('h4)
	) name6778 (
		_w7306_,
		_w7309_,
		_w7310_
	);
	LUT2 #(
		.INIT('h4)
	) name6779 (
		_w7301_,
		_w7310_,
		_w7311_
	);
	LUT2 #(
		.INIT('h4)
	) name6780 (
		_w7266_,
		_w7311_,
		_w7312_
	);
	LUT2 #(
		.INIT('h4)
	) name6781 (
		_w7290_,
		_w7312_,
		_w7313_
	);
	LUT2 #(
		.INIT('h2)
	) name6782 (
		\u0_w_reg[2][12]/P0001 ,
		_w7313_,
		_w7314_
	);
	LUT2 #(
		.INIT('h4)
	) name6783 (
		\u0_w_reg[2][12]/P0001 ,
		_w7313_,
		_w7315_
	);
	LUT2 #(
		.INIT('h1)
	) name6784 (
		_w7314_,
		_w7315_,
		_w7316_
	);
	LUT2 #(
		.INIT('h8)
	) name6785 (
		_w7236_,
		_w7316_,
		_w7317_
	);
	LUT2 #(
		.INIT('h1)
	) name6786 (
		_w7236_,
		_w7316_,
		_w7318_
	);
	LUT2 #(
		.INIT('h1)
	) name6787 (
		_w7317_,
		_w7318_,
		_w7319_
	);
	LUT2 #(
		.INIT('h2)
	) name6788 (
		_w5631_,
		_w7206_,
		_w7320_
	);
	LUT2 #(
		.INIT('h4)
	) name6789 (
		_w5631_,
		_w7206_,
		_w7321_
	);
	LUT2 #(
		.INIT('h1)
	) name6790 (
		_w7320_,
		_w7321_,
		_w7322_
	);
	LUT2 #(
		.INIT('h4)
	) name6791 (
		_w5833_,
		_w7322_,
		_w7323_
	);
	LUT2 #(
		.INIT('h2)
	) name6792 (
		_w5833_,
		_w7322_,
		_w7324_
	);
	LUT2 #(
		.INIT('h1)
	) name6793 (
		_w7323_,
		_w7324_,
		_w7325_
	);
	LUT2 #(
		.INIT('h1)
	) name6794 (
		_w7319_,
		_w7325_,
		_w7326_
	);
	LUT2 #(
		.INIT('h8)
	) name6795 (
		_w7319_,
		_w7325_,
		_w7327_
	);
	LUT2 #(
		.INIT('h1)
	) name6796 (
		\ld_r_reg/P0001 ,
		_w7326_,
		_w7328_
	);
	LUT2 #(
		.INIT('h4)
	) name6797 (
		_w7327_,
		_w7328_,
		_w7329_
	);
	LUT2 #(
		.INIT('h2)
	) name6798 (
		\text_in_r_reg[44]/P0001 ,
		\u0_w_reg[2][12]/P0001 ,
		_w7330_
	);
	LUT2 #(
		.INIT('h4)
	) name6799 (
		\text_in_r_reg[44]/P0001 ,
		\u0_w_reg[2][12]/P0001 ,
		_w7331_
	);
	LUT2 #(
		.INIT('h2)
	) name6800 (
		\ld_r_reg/P0001 ,
		_w7330_,
		_w7332_
	);
	LUT2 #(
		.INIT('h4)
	) name6801 (
		_w7331_,
		_w7332_,
		_w7333_
	);
	LUT2 #(
		.INIT('h1)
	) name6802 (
		_w7329_,
		_w7333_,
		_w7334_
	);
	LUT2 #(
		.INIT('h2)
	) name6803 (
		\sa13_reg[5]/P0001 ,
		_w549_,
		_w7335_
	);
	LUT2 #(
		.INIT('h2)
	) name6804 (
		_w655_,
		_w7335_,
		_w7336_
	);
	LUT2 #(
		.INIT('h8)
	) name6805 (
		\sa13_reg[4]/P0001 ,
		_w5446_,
		_w7337_
	);
	LUT2 #(
		.INIT('h8)
	) name6806 (
		_w653_,
		_w900_,
		_w7338_
	);
	LUT2 #(
		.INIT('h1)
	) name6807 (
		_w651_,
		_w913_,
		_w7339_
	);
	LUT2 #(
		.INIT('h4)
	) name6808 (
		_w858_,
		_w7339_,
		_w7340_
	);
	LUT2 #(
		.INIT('h2)
	) name6809 (
		\sa13_reg[2]/P0001 ,
		_w7340_,
		_w7341_
	);
	LUT2 #(
		.INIT('h1)
	) name6810 (
		_w7336_,
		_w7338_,
		_w7342_
	);
	LUT2 #(
		.INIT('h4)
	) name6811 (
		_w7337_,
		_w7342_,
		_w7343_
	);
	LUT2 #(
		.INIT('h4)
	) name6812 (
		_w7341_,
		_w7343_,
		_w7344_
	);
	LUT2 #(
		.INIT('h1)
	) name6813 (
		\sa13_reg[1]/P0001 ,
		_w7344_,
		_w7345_
	);
	LUT2 #(
		.INIT('h1)
	) name6814 (
		_w921_,
		_w5679_,
		_w7346_
	);
	LUT2 #(
		.INIT('h8)
	) name6815 (
		_w562_,
		_w7346_,
		_w7347_
	);
	LUT2 #(
		.INIT('h2)
	) name6816 (
		\sa13_reg[2]/P0001 ,
		_w7347_,
		_w7348_
	);
	LUT2 #(
		.INIT('h1)
	) name6817 (
		_w907_,
		_w5438_,
		_w7349_
	);
	LUT2 #(
		.INIT('h1)
	) name6818 (
		\sa13_reg[2]/P0001 ,
		_w7349_,
		_w7350_
	);
	LUT2 #(
		.INIT('h1)
	) name6819 (
		_w536_,
		_w912_,
		_w7351_
	);
	LUT2 #(
		.INIT('h2)
	) name6820 (
		_w581_,
		_w7351_,
		_w7352_
	);
	LUT2 #(
		.INIT('h1)
	) name6821 (
		_w535_,
		_w650_,
		_w7353_
	);
	LUT2 #(
		.INIT('h1)
	) name6822 (
		\sa13_reg[2]/P0001 ,
		_w7353_,
		_w7354_
	);
	LUT2 #(
		.INIT('h1)
	) name6823 (
		_w665_,
		_w7354_,
		_w7355_
	);
	LUT2 #(
		.INIT('h2)
	) name6824 (
		\sa13_reg[1]/P0001 ,
		_w7355_,
		_w7356_
	);
	LUT2 #(
		.INIT('h1)
	) name6825 (
		_w862_,
		_w5704_,
		_w7357_
	);
	LUT2 #(
		.INIT('h4)
	) name6826 (
		_w7352_,
		_w7357_,
		_w7358_
	);
	LUT2 #(
		.INIT('h4)
	) name6827 (
		_w7350_,
		_w7358_,
		_w7359_
	);
	LUT2 #(
		.INIT('h4)
	) name6828 (
		_w7348_,
		_w7359_,
		_w7360_
	);
	LUT2 #(
		.INIT('h4)
	) name6829 (
		_w7356_,
		_w7360_,
		_w7361_
	);
	LUT2 #(
		.INIT('h4)
	) name6830 (
		_w7345_,
		_w7361_,
		_w7362_
	);
	LUT2 #(
		.INIT('h2)
	) name6831 (
		\sa13_reg[0]/P0001 ,
		_w7362_,
		_w7363_
	);
	LUT2 #(
		.INIT('h4)
	) name6832 (
		_w642_,
		_w7084_,
		_w7364_
	);
	LUT2 #(
		.INIT('h1)
	) name6833 (
		\sa13_reg[2]/P0001 ,
		_w7364_,
		_w7365_
	);
	LUT2 #(
		.INIT('h1)
	) name6834 (
		_w557_,
		_w912_,
		_w7366_
	);
	LUT2 #(
		.INIT('h2)
	) name6835 (
		_w883_,
		_w7366_,
		_w7367_
	);
	LUT2 #(
		.INIT('h1)
	) name6836 (
		_w568_,
		_w963_,
		_w7368_
	);
	LUT2 #(
		.INIT('h2)
	) name6837 (
		_w6272_,
		_w7368_,
		_w7369_
	);
	LUT2 #(
		.INIT('h1)
	) name6838 (
		_w555_,
		_w556_,
		_w7370_
	);
	LUT2 #(
		.INIT('h1)
	) name6839 (
		_w635_,
		_w7370_,
		_w7371_
	);
	LUT2 #(
		.INIT('h8)
	) name6840 (
		_w623_,
		_w861_,
		_w7372_
	);
	LUT2 #(
		.INIT('h8)
	) name6841 (
		_w570_,
		_w5424_,
		_w7373_
	);
	LUT2 #(
		.INIT('h2)
	) name6842 (
		\sa13_reg[1]/P0001 ,
		_w5442_,
		_w7374_
	);
	LUT2 #(
		.INIT('h4)
	) name6843 (
		_w7373_,
		_w7374_,
		_w7375_
	);
	LUT2 #(
		.INIT('h1)
	) name6844 (
		_w7371_,
		_w7372_,
		_w7376_
	);
	LUT2 #(
		.INIT('h8)
	) name6845 (
		_w7375_,
		_w7376_,
		_w7377_
	);
	LUT2 #(
		.INIT('h1)
	) name6846 (
		\sa13_reg[3]/P0001 ,
		_w5487_,
		_w7378_
	);
	LUT2 #(
		.INIT('h1)
	) name6847 (
		\sa13_reg[1]/P0001 ,
		_w5649_,
		_w7379_
	);
	LUT2 #(
		.INIT('h4)
	) name6848 (
		_w7378_,
		_w7379_,
		_w7380_
	);
	LUT2 #(
		.INIT('h1)
	) name6849 (
		_w7377_,
		_w7380_,
		_w7381_
	);
	LUT2 #(
		.INIT('h1)
	) name6850 (
		_w7367_,
		_w7369_,
		_w7382_
	);
	LUT2 #(
		.INIT('h4)
	) name6851 (
		_w7365_,
		_w7382_,
		_w7383_
	);
	LUT2 #(
		.INIT('h4)
	) name6852 (
		_w7381_,
		_w7383_,
		_w7384_
	);
	LUT2 #(
		.INIT('h1)
	) name6853 (
		\sa13_reg[0]/P0001 ,
		_w7384_,
		_w7385_
	);
	LUT2 #(
		.INIT('h1)
	) name6854 (
		_w668_,
		_w5680_,
		_w7386_
	);
	LUT2 #(
		.INIT('h2)
	) name6855 (
		_w6272_,
		_w7386_,
		_w7387_
	);
	LUT2 #(
		.INIT('h8)
	) name6856 (
		_w603_,
		_w901_,
		_w7388_
	);
	LUT2 #(
		.INIT('h1)
	) name6857 (
		_w625_,
		_w7388_,
		_w7389_
	);
	LUT2 #(
		.INIT('h2)
	) name6858 (
		\sa13_reg[6]/NET0131 ,
		_w7389_,
		_w7390_
	);
	LUT2 #(
		.INIT('h4)
	) name6859 (
		\sa13_reg[2]/P0001 ,
		_w5504_,
		_w7391_
	);
	LUT2 #(
		.INIT('h8)
	) name6860 (
		\sa13_reg[4]/P0001 ,
		_w877_,
		_w7392_
	);
	LUT2 #(
		.INIT('h1)
	) name6861 (
		_w551_,
		_w7392_,
		_w7393_
	);
	LUT2 #(
		.INIT('h2)
	) name6862 (
		\sa13_reg[2]/P0001 ,
		_w7393_,
		_w7394_
	);
	LUT2 #(
		.INIT('h1)
	) name6863 (
		_w683_,
		_w7391_,
		_w7395_
	);
	LUT2 #(
		.INIT('h8)
	) name6864 (
		_w5657_,
		_w7395_,
		_w7396_
	);
	LUT2 #(
		.INIT('h4)
	) name6865 (
		_w7394_,
		_w7396_,
		_w7397_
	);
	LUT2 #(
		.INIT('h1)
	) name6866 (
		_w877_,
		_w911_,
		_w7398_
	);
	LUT2 #(
		.INIT('h1)
	) name6867 (
		_w5422_,
		_w5678_,
		_w7399_
	);
	LUT2 #(
		.INIT('h8)
	) name6868 (
		_w7398_,
		_w7399_,
		_w7400_
	);
	LUT2 #(
		.INIT('h1)
	) name6869 (
		\sa13_reg[2]/P0001 ,
		_w7400_,
		_w7401_
	);
	LUT2 #(
		.INIT('h1)
	) name6870 (
		\sa13_reg[1]/P0001 ,
		_w953_,
		_w7402_
	);
	LUT2 #(
		.INIT('h4)
	) name6871 (
		_w7401_,
		_w7402_,
		_w7403_
	);
	LUT2 #(
		.INIT('h1)
	) name6872 (
		_w7397_,
		_w7403_,
		_w7404_
	);
	LUT2 #(
		.INIT('h1)
	) name6873 (
		_w7387_,
		_w7390_,
		_w7405_
	);
	LUT2 #(
		.INIT('h4)
	) name6874 (
		_w7404_,
		_w7405_,
		_w7406_
	);
	LUT2 #(
		.INIT('h4)
	) name6875 (
		_w7385_,
		_w7406_,
		_w7407_
	);
	LUT2 #(
		.INIT('h4)
	) name6876 (
		_w7363_,
		_w7407_,
		_w7408_
	);
	LUT2 #(
		.INIT('h2)
	) name6877 (
		_w5516_,
		_w7408_,
		_w7409_
	);
	LUT2 #(
		.INIT('h4)
	) name6878 (
		_w5516_,
		_w7408_,
		_w7410_
	);
	LUT2 #(
		.INIT('h1)
	) name6879 (
		_w7409_,
		_w7410_,
		_w7411_
	);
	LUT2 #(
		.INIT('h2)
	) name6880 (
		_w6392_,
		_w6927_,
		_w7412_
	);
	LUT2 #(
		.INIT('h4)
	) name6881 (
		_w6392_,
		_w6927_,
		_w7413_
	);
	LUT2 #(
		.INIT('h1)
	) name6882 (
		_w7412_,
		_w7413_,
		_w7414_
	);
	LUT2 #(
		.INIT('h8)
	) name6883 (
		_w7411_,
		_w7414_,
		_w7415_
	);
	LUT2 #(
		.INIT('h1)
	) name6884 (
		_w7411_,
		_w7414_,
		_w7416_
	);
	LUT2 #(
		.INIT('h1)
	) name6885 (
		_w7415_,
		_w7416_,
		_w7417_
	);
	LUT2 #(
		.INIT('h1)
	) name6886 (
		\u0_w_reg[2][17]/P0001 ,
		_w6842_,
		_w7418_
	);
	LUT2 #(
		.INIT('h8)
	) name6887 (
		\u0_w_reg[2][17]/P0001 ,
		_w6842_,
		_w7419_
	);
	LUT2 #(
		.INIT('h1)
	) name6888 (
		_w7418_,
		_w7419_,
		_w7420_
	);
	LUT2 #(
		.INIT('h2)
	) name6889 (
		_w5631_,
		_w6743_,
		_w7421_
	);
	LUT2 #(
		.INIT('h4)
	) name6890 (
		_w5631_,
		_w6743_,
		_w7422_
	);
	LUT2 #(
		.INIT('h1)
	) name6891 (
		_w7421_,
		_w7422_,
		_w7423_
	);
	LUT2 #(
		.INIT('h8)
	) name6892 (
		_w7420_,
		_w7423_,
		_w7424_
	);
	LUT2 #(
		.INIT('h1)
	) name6893 (
		_w7420_,
		_w7423_,
		_w7425_
	);
	LUT2 #(
		.INIT('h1)
	) name6894 (
		_w7424_,
		_w7425_,
		_w7426_
	);
	LUT2 #(
		.INIT('h1)
	) name6895 (
		_w7417_,
		_w7426_,
		_w7427_
	);
	LUT2 #(
		.INIT('h8)
	) name6896 (
		_w7417_,
		_w7426_,
		_w7428_
	);
	LUT2 #(
		.INIT('h1)
	) name6897 (
		\ld_r_reg/P0001 ,
		_w7427_,
		_w7429_
	);
	LUT2 #(
		.INIT('h4)
	) name6898 (
		_w7428_,
		_w7429_,
		_w7430_
	);
	LUT2 #(
		.INIT('h1)
	) name6899 (
		\text_in_r_reg[49]/P0001 ,
		\u0_w_reg[2][17]/P0001 ,
		_w7431_
	);
	LUT2 #(
		.INIT('h8)
	) name6900 (
		\text_in_r_reg[49]/P0001 ,
		\u0_w_reg[2][17]/P0001 ,
		_w7432_
	);
	LUT2 #(
		.INIT('h2)
	) name6901 (
		\ld_r_reg/P0001 ,
		_w7431_,
		_w7433_
	);
	LUT2 #(
		.INIT('h4)
	) name6902 (
		_w7432_,
		_w7433_,
		_w7434_
	);
	LUT2 #(
		.INIT('h1)
	) name6903 (
		_w7430_,
		_w7434_,
		_w7435_
	);
	LUT2 #(
		.INIT('h1)
	) name6904 (
		_w654_,
		_w913_,
		_w7436_
	);
	LUT2 #(
		.INIT('h1)
	) name6905 (
		\sa13_reg[2]/P0001 ,
		_w7436_,
		_w7437_
	);
	LUT2 #(
		.INIT('h8)
	) name6906 (
		_w543_,
		_w603_,
		_w7438_
	);
	LUT2 #(
		.INIT('h1)
	) name6907 (
		_w5661_,
		_w7338_,
		_w7439_
	);
	LUT2 #(
		.INIT('h4)
	) name6908 (
		_w7438_,
		_w7439_,
		_w7440_
	);
	LUT2 #(
		.INIT('h1)
	) name6909 (
		_w589_,
		_w5651_,
		_w7441_
	);
	LUT2 #(
		.INIT('h4)
	) name6910 (
		_w5725_,
		_w7441_,
		_w7442_
	);
	LUT2 #(
		.INIT('h4)
	) name6911 (
		_w7437_,
		_w7440_,
		_w7443_
	);
	LUT2 #(
		.INIT('h8)
	) name6912 (
		_w7442_,
		_w7443_,
		_w7444_
	);
	LUT2 #(
		.INIT('h1)
	) name6913 (
		\sa13_reg[1]/P0001 ,
		_w7444_,
		_w7445_
	);
	LUT2 #(
		.INIT('h8)
	) name6914 (
		\sa13_reg[1]/P0001 ,
		_w672_,
		_w7446_
	);
	LUT2 #(
		.INIT('h1)
	) name6915 (
		_w540_,
		_w665_,
		_w7447_
	);
	LUT2 #(
		.INIT('h4)
	) name6916 (
		_w5466_,
		_w7447_,
		_w7448_
	);
	LUT2 #(
		.INIT('h2)
	) name6917 (
		\sa13_reg[3]/P0001 ,
		_w7448_,
		_w7449_
	);
	LUT2 #(
		.INIT('h1)
	) name6918 (
		_w862_,
		_w7446_,
		_w7450_
	);
	LUT2 #(
		.INIT('h4)
	) name6919 (
		_w7449_,
		_w7450_,
		_w7451_
	);
	LUT2 #(
		.INIT('h2)
	) name6920 (
		\sa13_reg[2]/P0001 ,
		_w7451_,
		_w7452_
	);
	LUT2 #(
		.INIT('h1)
	) name6921 (
		_w620_,
		_w632_,
		_w7453_
	);
	LUT2 #(
		.INIT('h4)
	) name6922 (
		_w911_,
		_w7453_,
		_w7454_
	);
	LUT2 #(
		.INIT('h2)
	) name6923 (
		_w680_,
		_w7454_,
		_w7455_
	);
	LUT2 #(
		.INIT('h1)
	) name6924 (
		_w5678_,
		_w5680_,
		_w7456_
	);
	LUT2 #(
		.INIT('h4)
	) name6925 (
		_w7455_,
		_w7456_,
		_w7457_
	);
	LUT2 #(
		.INIT('h4)
	) name6926 (
		_w7445_,
		_w7457_,
		_w7458_
	);
	LUT2 #(
		.INIT('h4)
	) name6927 (
		_w7452_,
		_w7458_,
		_w7459_
	);
	LUT2 #(
		.INIT('h2)
	) name6928 (
		\sa13_reg[0]/P0001 ,
		_w7459_,
		_w7460_
	);
	LUT2 #(
		.INIT('h1)
	) name6929 (
		_w609_,
		_w669_,
		_w7461_
	);
	LUT2 #(
		.INIT('h4)
	) name6930 (
		_w5492_,
		_w7461_,
		_w7462_
	);
	LUT2 #(
		.INIT('h8)
	) name6931 (
		_w590_,
		_w7462_,
		_w7463_
	);
	LUT2 #(
		.INIT('h2)
	) name6932 (
		\sa13_reg[2]/P0001 ,
		_w955_,
		_w7464_
	);
	LUT2 #(
		.INIT('h4)
	) name6933 (
		_w5504_,
		_w7464_,
		_w7465_
	);
	LUT2 #(
		.INIT('h4)
	) name6934 (
		_w5687_,
		_w7465_,
		_w7466_
	);
	LUT2 #(
		.INIT('h1)
	) name6935 (
		_w7463_,
		_w7466_,
		_w7467_
	);
	LUT2 #(
		.INIT('h1)
	) name6936 (
		_w533_,
		_w536_,
		_w7468_
	);
	LUT2 #(
		.INIT('h8)
	) name6937 (
		_w547_,
		_w7468_,
		_w7469_
	);
	LUT2 #(
		.INIT('h1)
	) name6938 (
		_w7467_,
		_w7469_,
		_w7470_
	);
	LUT2 #(
		.INIT('h1)
	) name6939 (
		\sa13_reg[1]/P0001 ,
		_w7470_,
		_w7471_
	);
	LUT2 #(
		.INIT('h4)
	) name6940 (
		\sa13_reg[6]/NET0131 ,
		_w884_,
		_w7472_
	);
	LUT2 #(
		.INIT('h2)
	) name6941 (
		_w6244_,
		_w7472_,
		_w7473_
	);
	LUT2 #(
		.INIT('h1)
	) name6942 (
		\sa13_reg[2]/P0001 ,
		_w7473_,
		_w7474_
	);
	LUT2 #(
		.INIT('h1)
	) name6943 (
		_w856_,
		_w7474_,
		_w7475_
	);
	LUT2 #(
		.INIT('h2)
	) name6944 (
		\sa13_reg[1]/P0001 ,
		_w7475_,
		_w7476_
	);
	LUT2 #(
		.INIT('h8)
	) name6945 (
		\sa13_reg[2]/P0001 ,
		_w6283_,
		_w7477_
	);
	LUT2 #(
		.INIT('h8)
	) name6946 (
		_w908_,
		_w7477_,
		_w7478_
	);
	LUT2 #(
		.INIT('h1)
	) name6947 (
		_w557_,
		_w570_,
		_w7479_
	);
	LUT2 #(
		.INIT('h2)
	) name6948 (
		_w653_,
		_w7479_,
		_w7480_
	);
	LUT2 #(
		.INIT('h1)
	) name6949 (
		_w913_,
		_w6252_,
		_w7481_
	);
	LUT2 #(
		.INIT('h2)
	) name6950 (
		\sa13_reg[1]/P0001 ,
		_w7481_,
		_w7482_
	);
	LUT2 #(
		.INIT('h1)
	) name6951 (
		_w7480_,
		_w7482_,
		_w7483_
	);
	LUT2 #(
		.INIT('h2)
	) name6952 (
		\sa13_reg[2]/P0001 ,
		_w7483_,
		_w7484_
	);
	LUT2 #(
		.INIT('h2)
	) name6953 (
		\sa13_reg[2]/P0001 ,
		_w5442_,
		_w7485_
	);
	LUT2 #(
		.INIT('h4)
	) name6954 (
		_w903_,
		_w7485_,
		_w7486_
	);
	LUT2 #(
		.INIT('h1)
	) name6955 (
		\sa13_reg[2]/P0001 ,
		_w604_,
		_w7487_
	);
	LUT2 #(
		.INIT('h1)
	) name6956 (
		_w5650_,
		_w6216_,
		_w7488_
	);
	LUT2 #(
		.INIT('h8)
	) name6957 (
		_w7487_,
		_w7488_,
		_w7489_
	);
	LUT2 #(
		.INIT('h1)
	) name6958 (
		_w7486_,
		_w7489_,
		_w7490_
	);
	LUT2 #(
		.INIT('h1)
	) name6959 (
		_w5476_,
		_w7490_,
		_w7491_
	);
	LUT2 #(
		.INIT('h2)
	) name6960 (
		\sa13_reg[1]/P0001 ,
		_w7491_,
		_w7492_
	);
	LUT2 #(
		.INIT('h4)
	) name6961 (
		\sa13_reg[1]/P0001 ,
		_w900_,
		_w7493_
	);
	LUT2 #(
		.INIT('h1)
	) name6962 (
		_w5492_,
		_w7493_,
		_w7494_
	);
	LUT2 #(
		.INIT('h2)
	) name6963 (
		_w581_,
		_w7494_,
		_w7495_
	);
	LUT2 #(
		.INIT('h8)
	) name6964 (
		_w5671_,
		_w6281_,
		_w7496_
	);
	LUT2 #(
		.INIT('h4)
	) name6965 (
		\sa13_reg[1]/P0001 ,
		_w5504_,
		_w7497_
	);
	LUT2 #(
		.INIT('h1)
	) name6966 (
		_w588_,
		_w7496_,
		_w7498_
	);
	LUT2 #(
		.INIT('h4)
	) name6967 (
		_w7497_,
		_w7498_,
		_w7499_
	);
	LUT2 #(
		.INIT('h4)
	) name6968 (
		_w7495_,
		_w7499_,
		_w7500_
	);
	LUT2 #(
		.INIT('h4)
	) name6969 (
		_w7492_,
		_w7500_,
		_w7501_
	);
	LUT2 #(
		.INIT('h1)
	) name6970 (
		\sa13_reg[0]/P0001 ,
		_w7501_,
		_w7502_
	);
	LUT2 #(
		.INIT('h1)
	) name6971 (
		_w7098_,
		_w7478_,
		_w7503_
	);
	LUT2 #(
		.INIT('h4)
	) name6972 (
		_w7484_,
		_w7503_,
		_w7504_
	);
	LUT2 #(
		.INIT('h4)
	) name6973 (
		_w7476_,
		_w7504_,
		_w7505_
	);
	LUT2 #(
		.INIT('h4)
	) name6974 (
		_w7471_,
		_w7505_,
		_w7506_
	);
	LUT2 #(
		.INIT('h4)
	) name6975 (
		_w7502_,
		_w7506_,
		_w7507_
	);
	LUT2 #(
		.INIT('h4)
	) name6976 (
		_w7460_,
		_w7507_,
		_w7508_
	);
	LUT2 #(
		.INIT('h4)
	) name6977 (
		_w1068_,
		_w5348_,
		_w7509_
	);
	LUT2 #(
		.INIT('h1)
	) name6978 (
		_w1070_,
		_w7509_,
		_w7510_
	);
	LUT2 #(
		.INIT('h1)
	) name6979 (
		\sa02_reg[2]/P0001 ,
		_w7510_,
		_w7511_
	);
	LUT2 #(
		.INIT('h1)
	) name6980 (
		_w5169_,
		_w7511_,
		_w7512_
	);
	LUT2 #(
		.INIT('h2)
	) name6981 (
		\sa02_reg[1]/P0001 ,
		_w7512_,
		_w7513_
	);
	LUT2 #(
		.INIT('h1)
	) name6982 (
		_w976_,
		_w5363_,
		_w7514_
	);
	LUT2 #(
		.INIT('h4)
	) name6983 (
		_w5163_,
		_w7514_,
		_w7515_
	);
	LUT2 #(
		.INIT('h2)
	) name6984 (
		_w984_,
		_w7515_,
		_w7516_
	);
	LUT2 #(
		.INIT('h1)
	) name6985 (
		_w5394_,
		_w5750_,
		_w7517_
	);
	LUT2 #(
		.INIT('h4)
	) name6986 (
		_w5754_,
		_w7517_,
		_w7518_
	);
	LUT2 #(
		.INIT('h1)
	) name6987 (
		\sa02_reg[3]/P0001 ,
		_w7518_,
		_w7519_
	);
	LUT2 #(
		.INIT('h1)
	) name6988 (
		_w1076_,
		_w1121_,
		_w7520_
	);
	LUT2 #(
		.INIT('h1)
	) name6989 (
		\sa02_reg[2]/P0001 ,
		_w7520_,
		_w7521_
	);
	LUT2 #(
		.INIT('h1)
	) name6990 (
		_w1113_,
		_w5766_,
		_w7522_
	);
	LUT2 #(
		.INIT('h4)
	) name6991 (
		_w5780_,
		_w7522_,
		_w7523_
	);
	LUT2 #(
		.INIT('h1)
	) name6992 (
		_w5092_,
		_w5754_,
		_w7524_
	);
	LUT2 #(
		.INIT('h4)
	) name6993 (
		_w5809_,
		_w7524_,
		_w7525_
	);
	LUT2 #(
		.INIT('h4)
	) name6994 (
		_w7521_,
		_w7523_,
		_w7526_
	);
	LUT2 #(
		.INIT('h8)
	) name6995 (
		_w7525_,
		_w7526_,
		_w7527_
	);
	LUT2 #(
		.INIT('h1)
	) name6996 (
		\sa02_reg[1]/P0001 ,
		_w7527_,
		_w7528_
	);
	LUT2 #(
		.INIT('h1)
	) name6997 (
		_w7516_,
		_w7519_,
		_w7529_
	);
	LUT2 #(
		.INIT('h4)
	) name6998 (
		_w7513_,
		_w7529_,
		_w7530_
	);
	LUT2 #(
		.INIT('h4)
	) name6999 (
		_w7528_,
		_w7530_,
		_w7531_
	);
	LUT2 #(
		.INIT('h2)
	) name7000 (
		\sa02_reg[0]/P0001 ,
		_w7531_,
		_w7532_
	);
	LUT2 #(
		.INIT('h1)
	) name7001 (
		_w1069_,
		_w5155_,
		_w7533_
	);
	LUT2 #(
		.INIT('h2)
	) name7002 (
		\sa02_reg[2]/P0001 ,
		_w7533_,
		_w7534_
	);
	LUT2 #(
		.INIT('h1)
	) name7003 (
		_w1015_,
		_w1068_,
		_w7535_
	);
	LUT2 #(
		.INIT('h1)
	) name7004 (
		\sa02_reg[2]/P0001 ,
		_w1056_,
		_w7536_
	);
	LUT2 #(
		.INIT('h4)
	) name7005 (
		_w7535_,
		_w7536_,
		_w7537_
	);
	LUT2 #(
		.INIT('h1)
	) name7006 (
		_w5156_,
		_w7537_,
		_w7538_
	);
	LUT2 #(
		.INIT('h4)
	) name7007 (
		_w7534_,
		_w7538_,
		_w7539_
	);
	LUT2 #(
		.INIT('h2)
	) name7008 (
		\sa02_reg[1]/P0001 ,
		_w7539_,
		_w7540_
	);
	LUT2 #(
		.INIT('h8)
	) name7009 (
		_w986_,
		_w6434_,
		_w7541_
	);
	LUT2 #(
		.INIT('h4)
	) name7010 (
		\sa02_reg[1]/P0001 ,
		_w5127_,
		_w7542_
	);
	LUT2 #(
		.INIT('h1)
	) name7011 (
		_w1110_,
		_w7542_,
		_w7543_
	);
	LUT2 #(
		.INIT('h1)
	) name7012 (
		\sa02_reg[2]/P0001 ,
		_w7543_,
		_w7544_
	);
	LUT2 #(
		.INIT('h8)
	) name7013 (
		\sa02_reg[2]/P0001 ,
		_w5338_,
		_w7545_
	);
	LUT2 #(
		.INIT('h1)
	) name7014 (
		_w1001_,
		_w7541_,
		_w7546_
	);
	LUT2 #(
		.INIT('h4)
	) name7015 (
		_w7545_,
		_w7546_,
		_w7547_
	);
	LUT2 #(
		.INIT('h4)
	) name7016 (
		_w7544_,
		_w7547_,
		_w7548_
	);
	LUT2 #(
		.INIT('h4)
	) name7017 (
		_w7540_,
		_w7548_,
		_w7549_
	);
	LUT2 #(
		.INIT('h1)
	) name7018 (
		\sa02_reg[0]/P0001 ,
		_w7549_,
		_w7550_
	);
	LUT2 #(
		.INIT('h1)
	) name7019 (
		_w1076_,
		_w1122_,
		_w7551_
	);
	LUT2 #(
		.INIT('h2)
	) name7020 (
		_w5154_,
		_w7551_,
		_w7552_
	);
	LUT2 #(
		.INIT('h8)
	) name7021 (
		\sa02_reg[1]/P0001 ,
		_w984_,
		_w7553_
	);
	LUT2 #(
		.INIT('h8)
	) name7022 (
		_w1072_,
		_w7553_,
		_w7554_
	);
	LUT2 #(
		.INIT('h1)
	) name7023 (
		_w1003_,
		_w5091_,
		_w7555_
	);
	LUT2 #(
		.INIT('h2)
	) name7024 (
		_w5342_,
		_w7555_,
		_w7556_
	);
	LUT2 #(
		.INIT('h1)
	) name7025 (
		\sa02_reg[6]/NET0131 ,
		_w986_,
		_w7557_
	);
	LUT2 #(
		.INIT('h8)
	) name7026 (
		_w6339_,
		_w7557_,
		_w7558_
	);
	LUT2 #(
		.INIT('h1)
	) name7027 (
		\sa02_reg[2]/P0001 ,
		_w5167_,
		_w7559_
	);
	LUT2 #(
		.INIT('h4)
	) name7028 (
		_w5092_,
		_w7559_,
		_w7560_
	);
	LUT2 #(
		.INIT('h1)
	) name7029 (
		_w5122_,
		_w5394_,
		_w7561_
	);
	LUT2 #(
		.INIT('h8)
	) name7030 (
		_w7560_,
		_w7561_,
		_w7562_
	);
	LUT2 #(
		.INIT('h2)
	) name7031 (
		\sa02_reg[2]/P0001 ,
		_w1036_,
		_w7563_
	);
	LUT2 #(
		.INIT('h4)
	) name7032 (
		_w5409_,
		_w7563_,
		_w7564_
	);
	LUT2 #(
		.INIT('h4)
	) name7033 (
		_w5805_,
		_w7564_,
		_w7565_
	);
	LUT2 #(
		.INIT('h1)
	) name7034 (
		_w7562_,
		_w7565_,
		_w7566_
	);
	LUT2 #(
		.INIT('h1)
	) name7035 (
		\sa02_reg[1]/P0001 ,
		_w7558_,
		_w7567_
	);
	LUT2 #(
		.INIT('h4)
	) name7036 (
		_w7566_,
		_w7567_,
		_w7568_
	);
	LUT2 #(
		.INIT('h8)
	) name7037 (
		\sa02_reg[4]/P0001 ,
		_w6312_,
		_w7569_
	);
	LUT2 #(
		.INIT('h2)
	) name7038 (
		_w6338_,
		_w7569_,
		_w7570_
	);
	LUT2 #(
		.INIT('h1)
	) name7039 (
		\sa02_reg[2]/P0001 ,
		_w7570_,
		_w7571_
	);
	LUT2 #(
		.INIT('h2)
	) name7040 (
		\sa02_reg[1]/P0001 ,
		_w1021_,
		_w7572_
	);
	LUT2 #(
		.INIT('h4)
	) name7041 (
		_w7571_,
		_w7572_,
		_w7573_
	);
	LUT2 #(
		.INIT('h1)
	) name7042 (
		_w7568_,
		_w7573_,
		_w7574_
	);
	LUT2 #(
		.INIT('h1)
	) name7043 (
		_w7019_,
		_w7554_,
		_w7575_
	);
	LUT2 #(
		.INIT('h1)
	) name7044 (
		_w7552_,
		_w7556_,
		_w7576_
	);
	LUT2 #(
		.INIT('h8)
	) name7045 (
		_w7575_,
		_w7576_,
		_w7577_
	);
	LUT2 #(
		.INIT('h4)
	) name7046 (
		_w7550_,
		_w7577_,
		_w7578_
	);
	LUT2 #(
		.INIT('h4)
	) name7047 (
		_w7574_,
		_w7578_,
		_w7579_
	);
	LUT2 #(
		.INIT('h4)
	) name7048 (
		_w7532_,
		_w7579_,
		_w7580_
	);
	LUT2 #(
		.INIT('h2)
	) name7049 (
		_w7508_,
		_w7580_,
		_w7581_
	);
	LUT2 #(
		.INIT('h4)
	) name7050 (
		_w7508_,
		_w7580_,
		_w7582_
	);
	LUT2 #(
		.INIT('h1)
	) name7051 (
		_w7581_,
		_w7582_,
		_w7583_
	);
	LUT2 #(
		.INIT('h1)
	) name7052 (
		_w6392_,
		_w7583_,
		_w7584_
	);
	LUT2 #(
		.INIT('h8)
	) name7053 (
		_w6392_,
		_w7583_,
		_w7585_
	);
	LUT2 #(
		.INIT('h1)
	) name7054 (
		_w7584_,
		_w7585_,
		_w7586_
	);
	LUT2 #(
		.INIT('h8)
	) name7055 (
		\sa20_reg[4]/P0001 ,
		_w769_,
		_w7587_
	);
	LUT2 #(
		.INIT('h2)
	) name7056 (
		_w6690_,
		_w7587_,
		_w7588_
	);
	LUT2 #(
		.INIT('h1)
	) name7057 (
		\sa20_reg[2]/P0001 ,
		_w7588_,
		_w7589_
	);
	LUT2 #(
		.INIT('h1)
	) name7058 (
		_w737_,
		_w7589_,
		_w7590_
	);
	LUT2 #(
		.INIT('h2)
	) name7059 (
		\sa20_reg[1]/P0001 ,
		_w7590_,
		_w7591_
	);
	LUT2 #(
		.INIT('h1)
	) name7060 (
		\sa20_reg[2]/P0001 ,
		_w839_,
		_w7592_
	);
	LUT2 #(
		.INIT('h4)
	) name7061 (
		_w5573_,
		_w7592_,
		_w7593_
	);
	LUT2 #(
		.INIT('h1)
	) name7062 (
		_w725_,
		_w779_,
		_w7594_
	);
	LUT2 #(
		.INIT('h8)
	) name7063 (
		_w7593_,
		_w7594_,
		_w7595_
	);
	LUT2 #(
		.INIT('h2)
	) name7064 (
		\sa20_reg[2]/P0001 ,
		_w5617_,
		_w7596_
	);
	LUT2 #(
		.INIT('h4)
	) name7065 (
		_w5619_,
		_w7596_,
		_w7597_
	);
	LUT2 #(
		.INIT('h4)
	) name7066 (
		_w6043_,
		_w7597_,
		_w7598_
	);
	LUT2 #(
		.INIT('h1)
	) name7067 (
		_w7595_,
		_w7598_,
		_w7599_
	);
	LUT2 #(
		.INIT('h4)
	) name7068 (
		_w691_,
		_w708_,
		_w7600_
	);
	LUT2 #(
		.INIT('h4)
	) name7069 (
		_w709_,
		_w7600_,
		_w7601_
	);
	LUT2 #(
		.INIT('h1)
	) name7070 (
		_w7599_,
		_w7601_,
		_w7602_
	);
	LUT2 #(
		.INIT('h1)
	) name7071 (
		\sa20_reg[1]/P0001 ,
		_w7602_,
		_w7603_
	);
	LUT2 #(
		.INIT('h1)
	) name7072 (
		_w736_,
		_w5591_,
		_w7604_
	);
	LUT2 #(
		.INIT('h1)
	) name7073 (
		\sa20_reg[4]/P0001 ,
		_w7604_,
		_w7605_
	);
	LUT2 #(
		.INIT('h1)
	) name7074 (
		_w5907_,
		_w7605_,
		_w7606_
	);
	LUT2 #(
		.INIT('h2)
	) name7075 (
		_w806_,
		_w7606_,
		_w7607_
	);
	LUT2 #(
		.INIT('h1)
	) name7076 (
		_w720_,
		_w724_,
		_w7608_
	);
	LUT2 #(
		.INIT('h2)
	) name7077 (
		_w6906_,
		_w7608_,
		_w7609_
	);
	LUT2 #(
		.INIT('h1)
	) name7078 (
		_w832_,
		_w5858_,
		_w7610_
	);
	LUT2 #(
		.INIT('h4)
	) name7079 (
		_w5606_,
		_w7610_,
		_w7611_
	);
	LUT2 #(
		.INIT('h2)
	) name7080 (
		_w761_,
		_w7611_,
		_w7612_
	);
	LUT2 #(
		.INIT('h1)
	) name7081 (
		_w809_,
		_w5907_,
		_w7613_
	);
	LUT2 #(
		.INIT('h1)
	) name7082 (
		\sa20_reg[2]/P0001 ,
		_w7613_,
		_w7614_
	);
	LUT2 #(
		.INIT('h8)
	) name7083 (
		_w693_,
		_w819_,
		_w7615_
	);
	LUT2 #(
		.INIT('h1)
	) name7084 (
		_w5600_,
		_w5985_,
		_w7616_
	);
	LUT2 #(
		.INIT('h1)
	) name7085 (
		_w6001_,
		_w7615_,
		_w7617_
	);
	LUT2 #(
		.INIT('h8)
	) name7086 (
		_w7616_,
		_w7617_,
		_w7618_
	);
	LUT2 #(
		.INIT('h4)
	) name7087 (
		_w725_,
		_w6006_,
		_w7619_
	);
	LUT2 #(
		.INIT('h8)
	) name7088 (
		_w7618_,
		_w7619_,
		_w7620_
	);
	LUT2 #(
		.INIT('h4)
	) name7089 (
		_w7614_,
		_w7620_,
		_w7621_
	);
	LUT2 #(
		.INIT('h8)
	) name7090 (
		_w723_,
		_w5526_,
		_w7622_
	);
	LUT2 #(
		.INIT('h8)
	) name7091 (
		_w6663_,
		_w6867_,
		_w7623_
	);
	LUT2 #(
		.INIT('h2)
	) name7092 (
		\sa20_reg[1]/P0001 ,
		_w7622_,
		_w7624_
	);
	LUT2 #(
		.INIT('h4)
	) name7093 (
		_w6909_,
		_w7624_,
		_w7625_
	);
	LUT2 #(
		.INIT('h4)
	) name7094 (
		_w7623_,
		_w7625_,
		_w7626_
	);
	LUT2 #(
		.INIT('h1)
	) name7095 (
		_w7621_,
		_w7626_,
		_w7627_
	);
	LUT2 #(
		.INIT('h1)
	) name7096 (
		_w809_,
		_w7615_,
		_w7628_
	);
	LUT2 #(
		.INIT('h2)
	) name7097 (
		\sa20_reg[5]/P0001 ,
		_w7628_,
		_w7629_
	);
	LUT2 #(
		.INIT('h2)
	) name7098 (
		\sa20_reg[0]/P0001 ,
		_w6037_,
		_w7630_
	);
	LUT2 #(
		.INIT('h4)
	) name7099 (
		_w7629_,
		_w7630_,
		_w7631_
	);
	LUT2 #(
		.INIT('h4)
	) name7100 (
		_w7612_,
		_w7631_,
		_w7632_
	);
	LUT2 #(
		.INIT('h4)
	) name7101 (
		_w7627_,
		_w7632_,
		_w7633_
	);
	LUT2 #(
		.INIT('h1)
	) name7102 (
		_w698_,
		_w709_,
		_w7634_
	);
	LUT2 #(
		.INIT('h2)
	) name7103 (
		\sa20_reg[1]/P0001 ,
		_w777_,
		_w7635_
	);
	LUT2 #(
		.INIT('h1)
	) name7104 (
		\sa20_reg[2]/P0001 ,
		_w7635_,
		_w7636_
	);
	LUT2 #(
		.INIT('h1)
	) name7105 (
		_w7634_,
		_w7636_,
		_w7637_
	);
	LUT2 #(
		.INIT('h1)
	) name7106 (
		_w817_,
		_w7637_,
		_w7638_
	);
	LUT2 #(
		.INIT('h1)
	) name7107 (
		_w5618_,
		_w7638_,
		_w7639_
	);
	LUT2 #(
		.INIT('h1)
	) name7108 (
		_w5552_,
		_w5872_,
		_w7640_
	);
	LUT2 #(
		.INIT('h2)
	) name7109 (
		\sa20_reg[2]/P0001 ,
		_w7640_,
		_w7641_
	);
	LUT2 #(
		.INIT('h2)
	) name7110 (
		_w5590_,
		_w7641_,
		_w7642_
	);
	LUT2 #(
		.INIT('h8)
	) name7111 (
		_w763_,
		_w777_,
		_w7643_
	);
	LUT2 #(
		.INIT('h1)
	) name7112 (
		\sa20_reg[1]/P0001 ,
		_w5617_,
		_w7644_
	);
	LUT2 #(
		.INIT('h4)
	) name7113 (
		_w7643_,
		_w7644_,
		_w7645_
	);
	LUT2 #(
		.INIT('h1)
	) name7114 (
		_w7642_,
		_w7645_,
		_w7646_
	);
	LUT2 #(
		.INIT('h1)
	) name7115 (
		\sa20_reg[0]/P0001 ,
		_w715_,
		_w7647_
	);
	LUT2 #(
		.INIT('h4)
	) name7116 (
		_w7639_,
		_w7647_,
		_w7648_
	);
	LUT2 #(
		.INIT('h4)
	) name7117 (
		_w7646_,
		_w7648_,
		_w7649_
	);
	LUT2 #(
		.INIT('h1)
	) name7118 (
		_w7633_,
		_w7649_,
		_w7650_
	);
	LUT2 #(
		.INIT('h1)
	) name7119 (
		_w7185_,
		_w7609_,
		_w7651_
	);
	LUT2 #(
		.INIT('h4)
	) name7120 (
		_w7607_,
		_w7651_,
		_w7652_
	);
	LUT2 #(
		.INIT('h4)
	) name7121 (
		_w7591_,
		_w7652_,
		_w7653_
	);
	LUT2 #(
		.INIT('h4)
	) name7122 (
		_w7603_,
		_w7653_,
		_w7654_
	);
	LUT2 #(
		.INIT('h4)
	) name7123 (
		_w7650_,
		_w7654_,
		_w7655_
	);
	LUT2 #(
		.INIT('h2)
	) name7124 (
		\u0_w_reg[2][2]/P0001 ,
		_w7655_,
		_w7656_
	);
	LUT2 #(
		.INIT('h4)
	) name7125 (
		\u0_w_reg[2][2]/P0001 ,
		_w7655_,
		_w7657_
	);
	LUT2 #(
		.INIT('h1)
	) name7126 (
		_w7656_,
		_w7657_,
		_w7658_
	);
	LUT2 #(
		.INIT('h8)
	) name7127 (
		_w6842_,
		_w7658_,
		_w7659_
	);
	LUT2 #(
		.INIT('h1)
	) name7128 (
		_w6842_,
		_w7658_,
		_w7660_
	);
	LUT2 #(
		.INIT('h1)
	) name7129 (
		_w7659_,
		_w7660_,
		_w7661_
	);
	LUT2 #(
		.INIT('h4)
	) name7130 (
		_w7586_,
		_w7661_,
		_w7662_
	);
	LUT2 #(
		.INIT('h2)
	) name7131 (
		_w7586_,
		_w7661_,
		_w7663_
	);
	LUT2 #(
		.INIT('h1)
	) name7132 (
		\ld_r_reg/P0001 ,
		_w7662_,
		_w7664_
	);
	LUT2 #(
		.INIT('h4)
	) name7133 (
		_w7663_,
		_w7664_,
		_w7665_
	);
	LUT2 #(
		.INIT('h1)
	) name7134 (
		\text_in_r_reg[34]/P0001 ,
		\u0_w_reg[2][2]/P0001 ,
		_w7666_
	);
	LUT2 #(
		.INIT('h8)
	) name7135 (
		\text_in_r_reg[34]/P0001 ,
		\u0_w_reg[2][2]/P0001 ,
		_w7667_
	);
	LUT2 #(
		.INIT('h2)
	) name7136 (
		\ld_r_reg/P0001 ,
		_w7666_,
		_w7668_
	);
	LUT2 #(
		.INIT('h4)
	) name7137 (
		_w7667_,
		_w7668_,
		_w7669_
	);
	LUT2 #(
		.INIT('h1)
	) name7138 (
		_w7665_,
		_w7669_,
		_w7670_
	);
	LUT2 #(
		.INIT('h4)
	) name7139 (
		_w6304_,
		_w6743_,
		_w7671_
	);
	LUT2 #(
		.INIT('h2)
	) name7140 (
		_w6304_,
		_w6743_,
		_w7672_
	);
	LUT2 #(
		.INIT('h1)
	) name7141 (
		_w7671_,
		_w7672_,
		_w7673_
	);
	LUT2 #(
		.INIT('h2)
	) name7142 (
		\u0_w_reg[2][25]/P0001 ,
		_w6842_,
		_w7674_
	);
	LUT2 #(
		.INIT('h4)
	) name7143 (
		\u0_w_reg[2][25]/P0001 ,
		_w6842_,
		_w7675_
	);
	LUT2 #(
		.INIT('h1)
	) name7144 (
		_w7674_,
		_w7675_,
		_w7676_
	);
	LUT2 #(
		.INIT('h8)
	) name7145 (
		_w7673_,
		_w7676_,
		_w7677_
	);
	LUT2 #(
		.INIT('h1)
	) name7146 (
		_w7673_,
		_w7676_,
		_w7678_
	);
	LUT2 #(
		.INIT('h1)
	) name7147 (
		_w7677_,
		_w7678_,
		_w7679_
	);
	LUT2 #(
		.INIT('h8)
	) name7148 (
		_w6475_,
		_w7411_,
		_w7680_
	);
	LUT2 #(
		.INIT('h1)
	) name7149 (
		_w6475_,
		_w7411_,
		_w7681_
	);
	LUT2 #(
		.INIT('h1)
	) name7150 (
		_w7680_,
		_w7681_,
		_w7682_
	);
	LUT2 #(
		.INIT('h1)
	) name7151 (
		_w7679_,
		_w7682_,
		_w7683_
	);
	LUT2 #(
		.INIT('h8)
	) name7152 (
		_w7679_,
		_w7682_,
		_w7684_
	);
	LUT2 #(
		.INIT('h1)
	) name7153 (
		\ld_r_reg/P0001 ,
		_w7683_,
		_w7685_
	);
	LUT2 #(
		.INIT('h4)
	) name7154 (
		_w7684_,
		_w7685_,
		_w7686_
	);
	LUT2 #(
		.INIT('h1)
	) name7155 (
		\text_in_r_reg[57]/P0001 ,
		\u0_w_reg[2][25]/P0001 ,
		_w7687_
	);
	LUT2 #(
		.INIT('h8)
	) name7156 (
		\text_in_r_reg[57]/P0001 ,
		\u0_w_reg[2][25]/P0001 ,
		_w7688_
	);
	LUT2 #(
		.INIT('h2)
	) name7157 (
		\ld_r_reg/P0001 ,
		_w7687_,
		_w7689_
	);
	LUT2 #(
		.INIT('h4)
	) name7158 (
		_w7688_,
		_w7689_,
		_w7690_
	);
	LUT2 #(
		.INIT('h1)
	) name7159 (
		_w7686_,
		_w7690_,
		_w7691_
	);
	LUT2 #(
		.INIT('h1)
	) name7160 (
		_w850_,
		_w5519_,
		_w7692_
	);
	LUT2 #(
		.INIT('h8)
	) name7161 (
		_w850_,
		_w5519_,
		_w7693_
	);
	LUT2 #(
		.INIT('h1)
	) name7162 (
		_w7692_,
		_w7693_,
		_w7694_
	);
	LUT2 #(
		.INIT('h2)
	) name7163 (
		\u0_w_reg[2][15]/P0001 ,
		_w6657_,
		_w7695_
	);
	LUT2 #(
		.INIT('h4)
	) name7164 (
		\u0_w_reg[2][15]/P0001 ,
		_w6657_,
		_w7696_
	);
	LUT2 #(
		.INIT('h1)
	) name7165 (
		_w7695_,
		_w7696_,
		_w7697_
	);
	LUT2 #(
		.INIT('h8)
	) name7166 (
		_w1300_,
		_w7697_,
		_w7698_
	);
	LUT2 #(
		.INIT('h1)
	) name7167 (
		_w1300_,
		_w7697_,
		_w7699_
	);
	LUT2 #(
		.INIT('h1)
	) name7168 (
		_w7698_,
		_w7699_,
		_w7700_
	);
	LUT2 #(
		.INIT('h1)
	) name7169 (
		_w7694_,
		_w7700_,
		_w7701_
	);
	LUT2 #(
		.INIT('h8)
	) name7170 (
		_w7694_,
		_w7700_,
		_w7702_
	);
	LUT2 #(
		.INIT('h1)
	) name7171 (
		\ld_r_reg/P0001 ,
		_w7701_,
		_w7703_
	);
	LUT2 #(
		.INIT('h4)
	) name7172 (
		_w7702_,
		_w7703_,
		_w7704_
	);
	LUT2 #(
		.INIT('h2)
	) name7173 (
		\text_in_r_reg[47]/P0001 ,
		\u0_w_reg[2][15]/P0001 ,
		_w7705_
	);
	LUT2 #(
		.INIT('h4)
	) name7174 (
		\text_in_r_reg[47]/P0001 ,
		\u0_w_reg[2][15]/P0001 ,
		_w7706_
	);
	LUT2 #(
		.INIT('h2)
	) name7175 (
		\ld_r_reg/P0001 ,
		_w7705_,
		_w7707_
	);
	LUT2 #(
		.INIT('h4)
	) name7176 (
		_w7706_,
		_w7707_,
		_w7708_
	);
	LUT2 #(
		.INIT('h1)
	) name7177 (
		_w7704_,
		_w7708_,
		_w7709_
	);
	LUT2 #(
		.INIT('h2)
	) name7178 (
		_w5417_,
		_w7040_,
		_w7710_
	);
	LUT2 #(
		.INIT('h4)
	) name7179 (
		_w5417_,
		_w7040_,
		_w7711_
	);
	LUT2 #(
		.INIT('h1)
	) name7180 (
		_w7710_,
		_w7711_,
		_w7712_
	);
	LUT2 #(
		.INIT('h8)
	) name7181 (
		_w5833_,
		_w7712_,
		_w7713_
	);
	LUT2 #(
		.INIT('h1)
	) name7182 (
		_w5833_,
		_w7712_,
		_w7714_
	);
	LUT2 #(
		.INIT('h1)
	) name7183 (
		_w7713_,
		_w7714_,
		_w7715_
	);
	LUT2 #(
		.INIT('h1)
	) name7184 (
		_w6055_,
		_w6657_,
		_w7716_
	);
	LUT2 #(
		.INIT('h8)
	) name7185 (
		_w6055_,
		_w6657_,
		_w7717_
	);
	LUT2 #(
		.INIT('h1)
	) name7186 (
		_w7716_,
		_w7717_,
		_w7718_
	);
	LUT2 #(
		.INIT('h2)
	) name7187 (
		\u0_w_reg[2][4]/P0001 ,
		_w7313_,
		_w7719_
	);
	LUT2 #(
		.INIT('h4)
	) name7188 (
		\u0_w_reg[2][4]/P0001 ,
		_w7313_,
		_w7720_
	);
	LUT2 #(
		.INIT('h1)
	) name7189 (
		_w7719_,
		_w7720_,
		_w7721_
	);
	LUT2 #(
		.INIT('h8)
	) name7190 (
		_w7718_,
		_w7721_,
		_w7722_
	);
	LUT2 #(
		.INIT('h1)
	) name7191 (
		_w7718_,
		_w7721_,
		_w7723_
	);
	LUT2 #(
		.INIT('h1)
	) name7192 (
		_w7722_,
		_w7723_,
		_w7724_
	);
	LUT2 #(
		.INIT('h2)
	) name7193 (
		_w7715_,
		_w7724_,
		_w7725_
	);
	LUT2 #(
		.INIT('h4)
	) name7194 (
		_w7715_,
		_w7724_,
		_w7726_
	);
	LUT2 #(
		.INIT('h1)
	) name7195 (
		\ld_r_reg/P0001 ,
		_w7725_,
		_w7727_
	);
	LUT2 #(
		.INIT('h4)
	) name7196 (
		_w7726_,
		_w7727_,
		_w7728_
	);
	LUT2 #(
		.INIT('h2)
	) name7197 (
		\text_in_r_reg[36]/P0001 ,
		\u0_w_reg[2][4]/P0001 ,
		_w7729_
	);
	LUT2 #(
		.INIT('h4)
	) name7198 (
		\text_in_r_reg[36]/P0001 ,
		\u0_w_reg[2][4]/P0001 ,
		_w7730_
	);
	LUT2 #(
		.INIT('h2)
	) name7199 (
		\ld_r_reg/P0001 ,
		_w7729_,
		_w7731_
	);
	LUT2 #(
		.INIT('h4)
	) name7200 (
		_w7730_,
		_w7731_,
		_w7732_
	);
	LUT2 #(
		.INIT('h1)
	) name7201 (
		_w7728_,
		_w7732_,
		_w7733_
	);
	LUT2 #(
		.INIT('h2)
	) name7202 (
		\u0_w_reg[2][27]/P0001 ,
		_w7313_,
		_w7734_
	);
	LUT2 #(
		.INIT('h4)
	) name7203 (
		\u0_w_reg[2][27]/P0001 ,
		_w7313_,
		_w7735_
	);
	LUT2 #(
		.INIT('h1)
	) name7204 (
		_w7734_,
		_w7735_,
		_w7736_
	);
	LUT2 #(
		.INIT('h8)
	) name7205 (
		_w7209_,
		_w7736_,
		_w7737_
	);
	LUT2 #(
		.INIT('h1)
	) name7206 (
		_w7209_,
		_w7736_,
		_w7738_
	);
	LUT2 #(
		.INIT('h1)
	) name7207 (
		_w7737_,
		_w7738_,
		_w7739_
	);
	LUT2 #(
		.INIT('h4)
	) name7208 (
		_w5519_,
		_w7583_,
		_w7740_
	);
	LUT2 #(
		.INIT('h2)
	) name7209 (
		_w5519_,
		_w7583_,
		_w7741_
	);
	LUT2 #(
		.INIT('h1)
	) name7210 (
		_w7740_,
		_w7741_,
		_w7742_
	);
	LUT2 #(
		.INIT('h2)
	) name7211 (
		_w7739_,
		_w7742_,
		_w7743_
	);
	LUT2 #(
		.INIT('h4)
	) name7212 (
		_w7739_,
		_w7742_,
		_w7744_
	);
	LUT2 #(
		.INIT('h1)
	) name7213 (
		\ld_r_reg/P0001 ,
		_w7743_,
		_w7745_
	);
	LUT2 #(
		.INIT('h4)
	) name7214 (
		_w7744_,
		_w7745_,
		_w7746_
	);
	LUT2 #(
		.INIT('h2)
	) name7215 (
		\text_in_r_reg[59]/P0001 ,
		\u0_w_reg[2][27]/P0001 ,
		_w7747_
	);
	LUT2 #(
		.INIT('h4)
	) name7216 (
		\text_in_r_reg[59]/P0001 ,
		\u0_w_reg[2][27]/P0001 ,
		_w7748_
	);
	LUT2 #(
		.INIT('h2)
	) name7217 (
		\ld_r_reg/P0001 ,
		_w7747_,
		_w7749_
	);
	LUT2 #(
		.INIT('h4)
	) name7218 (
		_w7748_,
		_w7749_,
		_w7750_
	);
	LUT2 #(
		.INIT('h1)
	) name7219 (
		_w7746_,
		_w7750_,
		_w7751_
	);
	LUT2 #(
		.INIT('h2)
	) name7220 (
		\u0_w_reg[2][19]/P0001 ,
		_w7313_,
		_w7752_
	);
	LUT2 #(
		.INIT('h4)
	) name7221 (
		\u0_w_reg[2][19]/P0001 ,
		_w7313_,
		_w7753_
	);
	LUT2 #(
		.INIT('h1)
	) name7222 (
		_w7752_,
		_w7753_,
		_w7754_
	);
	LUT2 #(
		.INIT('h8)
	) name7223 (
		_w7322_,
		_w7754_,
		_w7755_
	);
	LUT2 #(
		.INIT('h1)
	) name7224 (
		_w7322_,
		_w7754_,
		_w7756_
	);
	LUT2 #(
		.INIT('h1)
	) name7225 (
		_w7755_,
		_w7756_,
		_w7757_
	);
	LUT2 #(
		.INIT('h2)
	) name7226 (
		_w7508_,
		_w7655_,
		_w7758_
	);
	LUT2 #(
		.INIT('h4)
	) name7227 (
		_w7508_,
		_w7655_,
		_w7759_
	);
	LUT2 #(
		.INIT('h1)
	) name7228 (
		_w7758_,
		_w7759_,
		_w7760_
	);
	LUT2 #(
		.INIT('h2)
	) name7229 (
		_w5516_,
		_w7040_,
		_w7761_
	);
	LUT2 #(
		.INIT('h4)
	) name7230 (
		_w5516_,
		_w7040_,
		_w7762_
	);
	LUT2 #(
		.INIT('h1)
	) name7231 (
		_w7761_,
		_w7762_,
		_w7763_
	);
	LUT2 #(
		.INIT('h8)
	) name7232 (
		_w7760_,
		_w7763_,
		_w7764_
	);
	LUT2 #(
		.INIT('h1)
	) name7233 (
		_w7760_,
		_w7763_,
		_w7765_
	);
	LUT2 #(
		.INIT('h1)
	) name7234 (
		_w7764_,
		_w7765_,
		_w7766_
	);
	LUT2 #(
		.INIT('h1)
	) name7235 (
		_w7757_,
		_w7766_,
		_w7767_
	);
	LUT2 #(
		.INIT('h8)
	) name7236 (
		_w7757_,
		_w7766_,
		_w7768_
	);
	LUT2 #(
		.INIT('h1)
	) name7237 (
		\ld_r_reg/P0001 ,
		_w7767_,
		_w7769_
	);
	LUT2 #(
		.INIT('h4)
	) name7238 (
		_w7768_,
		_w7769_,
		_w7770_
	);
	LUT2 #(
		.INIT('h2)
	) name7239 (
		\text_in_r_reg[51]/P0001 ,
		\u0_w_reg[2][19]/P0001 ,
		_w7771_
	);
	LUT2 #(
		.INIT('h4)
	) name7240 (
		\text_in_r_reg[51]/P0001 ,
		\u0_w_reg[2][19]/P0001 ,
		_w7772_
	);
	LUT2 #(
		.INIT('h2)
	) name7241 (
		\ld_r_reg/P0001 ,
		_w7771_,
		_w7773_
	);
	LUT2 #(
		.INIT('h4)
	) name7242 (
		_w7772_,
		_w7773_,
		_w7774_
	);
	LUT2 #(
		.INIT('h1)
	) name7243 (
		_w7770_,
		_w7774_,
		_w7775_
	);
	LUT2 #(
		.INIT('h2)
	) name7244 (
		_w5631_,
		_w7655_,
		_w7776_
	);
	LUT2 #(
		.INIT('h4)
	) name7245 (
		_w5631_,
		_w7655_,
		_w7777_
	);
	LUT2 #(
		.INIT('h1)
	) name7246 (
		_w7776_,
		_w7777_,
		_w7778_
	);
	LUT2 #(
		.INIT('h8)
	) name7247 (
		_w7118_,
		_w7778_,
		_w7779_
	);
	LUT2 #(
		.INIT('h1)
	) name7248 (
		_w7118_,
		_w7778_,
		_w7780_
	);
	LUT2 #(
		.INIT('h1)
	) name7249 (
		_w7779_,
		_w7780_,
		_w7781_
	);
	LUT2 #(
		.INIT('h1)
	) name7250 (
		_w1182_,
		_w1187_,
		_w7782_
	);
	LUT2 #(
		.INIT('h4)
	) name7251 (
		\sa31_reg[3]/P0001 ,
		_w1244_,
		_w7783_
	);
	LUT2 #(
		.INIT('h4)
	) name7252 (
		_w7782_,
		_w7783_,
		_w7784_
	);
	LUT2 #(
		.INIT('h4)
	) name7253 (
		\sa31_reg[5]/P0001 ,
		_w1160_,
		_w7785_
	);
	LUT2 #(
		.INIT('h1)
	) name7254 (
		_w1246_,
		_w6084_,
		_w7786_
	);
	LUT2 #(
		.INIT('h4)
	) name7255 (
		_w6168_,
		_w7786_,
		_w7787_
	);
	LUT2 #(
		.INIT('h8)
	) name7256 (
		_w6631_,
		_w7787_,
		_w7788_
	);
	LUT2 #(
		.INIT('h4)
	) name7257 (
		\sa31_reg[6]/NET0131 ,
		_w1216_,
		_w7789_
	);
	LUT2 #(
		.INIT('h2)
	) name7258 (
		\sa31_reg[2]/P0001 ,
		_w6556_,
		_w7790_
	);
	LUT2 #(
		.INIT('h4)
	) name7259 (
		_w7789_,
		_w7790_,
		_w7791_
	);
	LUT2 #(
		.INIT('h4)
	) name7260 (
		_w6160_,
		_w7791_,
		_w7792_
	);
	LUT2 #(
		.INIT('h1)
	) name7261 (
		_w7788_,
		_w7792_,
		_w7793_
	);
	LUT2 #(
		.INIT('h1)
	) name7262 (
		\sa31_reg[1]/P0001 ,
		_w6089_,
		_w7794_
	);
	LUT2 #(
		.INIT('h4)
	) name7263 (
		_w7785_,
		_w7794_,
		_w7795_
	);
	LUT2 #(
		.INIT('h4)
	) name7264 (
		_w7793_,
		_w7795_,
		_w7796_
	);
	LUT2 #(
		.INIT('h8)
	) name7265 (
		\sa31_reg[4]/P0001 ,
		_w1269_,
		_w7797_
	);
	LUT2 #(
		.INIT('h1)
	) name7266 (
		\sa31_reg[2]/P0001 ,
		_w7797_,
		_w7798_
	);
	LUT2 #(
		.INIT('h8)
	) name7267 (
		_w6788_,
		_w7798_,
		_w7799_
	);
	LUT2 #(
		.INIT('h8)
	) name7268 (
		_w1276_,
		_w5241_,
		_w7800_
	);
	LUT2 #(
		.INIT('h2)
	) name7269 (
		\sa31_reg[2]/P0001 ,
		_w1153_,
		_w7801_
	);
	LUT2 #(
		.INIT('h4)
	) name7270 (
		_w5261_,
		_w7801_,
		_w7802_
	);
	LUT2 #(
		.INIT('h4)
	) name7271 (
		_w7800_,
		_w7802_,
		_w7803_
	);
	LUT2 #(
		.INIT('h1)
	) name7272 (
		_w7799_,
		_w7803_,
		_w7804_
	);
	LUT2 #(
		.INIT('h2)
	) name7273 (
		\sa31_reg[1]/P0001 ,
		_w5206_,
		_w7805_
	);
	LUT2 #(
		.INIT('h4)
	) name7274 (
		_w7804_,
		_w7805_,
		_w7806_
	);
	LUT2 #(
		.INIT('h1)
	) name7275 (
		_w7796_,
		_w7806_,
		_w7807_
	);
	LUT2 #(
		.INIT('h1)
	) name7276 (
		_w1201_,
		_w1239_,
		_w7808_
	);
	LUT2 #(
		.INIT('h4)
	) name7277 (
		_w6627_,
		_w7808_,
		_w7809_
	);
	LUT2 #(
		.INIT('h2)
	) name7278 (
		_w1265_,
		_w7809_,
		_w7810_
	);
	LUT2 #(
		.INIT('h8)
	) name7279 (
		_w6136_,
		_w6599_,
		_w7811_
	);
	LUT2 #(
		.INIT('h1)
	) name7280 (
		\sa31_reg[1]/P0001 ,
		_w6127_,
		_w7812_
	);
	LUT2 #(
		.INIT('h1)
	) name7281 (
		_w6134_,
		_w6146_,
		_w7813_
	);
	LUT2 #(
		.INIT('h4)
	) name7282 (
		_w6499_,
		_w7813_,
		_w7814_
	);
	LUT2 #(
		.INIT('h4)
	) name7283 (
		_w5262_,
		_w7812_,
		_w7815_
	);
	LUT2 #(
		.INIT('h1)
	) name7284 (
		_w6087_,
		_w6168_,
		_w7816_
	);
	LUT2 #(
		.INIT('h4)
	) name7285 (
		_w7811_,
		_w7816_,
		_w7817_
	);
	LUT2 #(
		.INIT('h8)
	) name7286 (
		_w7814_,
		_w7815_,
		_w7818_
	);
	LUT2 #(
		.INIT('h8)
	) name7287 (
		_w7817_,
		_w7818_,
		_w7819_
	);
	LUT2 #(
		.INIT('h8)
	) name7288 (
		\sa31_reg[2]/P0001 ,
		_w5220_,
		_w7820_
	);
	LUT2 #(
		.INIT('h4)
	) name7289 (
		_w5269_,
		_w6573_,
		_w7821_
	);
	LUT2 #(
		.INIT('h1)
	) name7290 (
		_w5264_,
		_w7821_,
		_w7822_
	);
	LUT2 #(
		.INIT('h1)
	) name7291 (
		\sa31_reg[2]/P0001 ,
		_w7822_,
		_w7823_
	);
	LUT2 #(
		.INIT('h2)
	) name7292 (
		\sa31_reg[1]/P0001 ,
		_w7820_,
		_w7824_
	);
	LUT2 #(
		.INIT('h4)
	) name7293 (
		_w7823_,
		_w7824_,
		_w7825_
	);
	LUT2 #(
		.INIT('h1)
	) name7294 (
		_w7819_,
		_w7825_,
		_w7826_
	);
	LUT2 #(
		.INIT('h8)
	) name7295 (
		_w1194_,
		_w1279_,
		_w7827_
	);
	LUT2 #(
		.INIT('h2)
	) name7296 (
		\sa31_reg[0]/P0002 ,
		_w6159_,
		_w7828_
	);
	LUT2 #(
		.INIT('h4)
	) name7297 (
		_w7827_,
		_w7828_,
		_w7829_
	);
	LUT2 #(
		.INIT('h4)
	) name7298 (
		_w6540_,
		_w7829_,
		_w7830_
	);
	LUT2 #(
		.INIT('h4)
	) name7299 (
		_w7810_,
		_w7830_,
		_w7831_
	);
	LUT2 #(
		.INIT('h4)
	) name7300 (
		_w7826_,
		_w7831_,
		_w7832_
	);
	LUT2 #(
		.INIT('h2)
	) name7301 (
		\sa31_reg[2]/P0001 ,
		_w5271_,
		_w7833_
	);
	LUT2 #(
		.INIT('h4)
	) name7302 (
		_w6599_,
		_w7833_,
		_w7834_
	);
	LUT2 #(
		.INIT('h4)
	) name7303 (
		_w1158_,
		_w5269_,
		_w7835_
	);
	LUT2 #(
		.INIT('h1)
	) name7304 (
		\sa31_reg[2]/P0001 ,
		_w1204_,
		_w7836_
	);
	LUT2 #(
		.INIT('h4)
	) name7305 (
		_w7835_,
		_w7836_,
		_w7837_
	);
	LUT2 #(
		.INIT('h1)
	) name7306 (
		_w7834_,
		_w7837_,
		_w7838_
	);
	LUT2 #(
		.INIT('h2)
	) name7307 (
		_w6635_,
		_w7838_,
		_w7839_
	);
	LUT2 #(
		.INIT('h8)
	) name7308 (
		_w1158_,
		_w5238_,
		_w7840_
	);
	LUT2 #(
		.INIT('h1)
	) name7309 (
		\sa31_reg[1]/P0001 ,
		_w6556_,
		_w7841_
	);
	LUT2 #(
		.INIT('h4)
	) name7310 (
		_w7840_,
		_w7841_,
		_w7842_
	);
	LUT2 #(
		.INIT('h1)
	) name7311 (
		_w7839_,
		_w7842_,
		_w7843_
	);
	LUT2 #(
		.INIT('h8)
	) name7312 (
		\sa31_reg[2]/P0001 ,
		_w6153_,
		_w7844_
	);
	LUT2 #(
		.INIT('h4)
	) name7313 (
		\sa31_reg[2]/P0001 ,
		_w1227_,
		_w7845_
	);
	LUT2 #(
		.INIT('h1)
	) name7314 (
		\sa31_reg[0]/P0002 ,
		_w1179_,
		_w7846_
	);
	LUT2 #(
		.INIT('h4)
	) name7315 (
		_w7844_,
		_w7846_,
		_w7847_
	);
	LUT2 #(
		.INIT('h4)
	) name7316 (
		_w7845_,
		_w7847_,
		_w7848_
	);
	LUT2 #(
		.INIT('h4)
	) name7317 (
		_w7843_,
		_w7848_,
		_w7849_
	);
	LUT2 #(
		.INIT('h1)
	) name7318 (
		_w7832_,
		_w7849_,
		_w7850_
	);
	LUT2 #(
		.INIT('h1)
	) name7319 (
		_w7297_,
		_w7784_,
		_w7851_
	);
	LUT2 #(
		.INIT('h4)
	) name7320 (
		_w7807_,
		_w7851_,
		_w7852_
	);
	LUT2 #(
		.INIT('h4)
	) name7321 (
		_w7850_,
		_w7852_,
		_w7853_
	);
	LUT2 #(
		.INIT('h2)
	) name7322 (
		_w6657_,
		_w7853_,
		_w7854_
	);
	LUT2 #(
		.INIT('h4)
	) name7323 (
		_w6657_,
		_w7853_,
		_w7855_
	);
	LUT2 #(
		.INIT('h1)
	) name7324 (
		_w7854_,
		_w7855_,
		_w7856_
	);
	LUT2 #(
		.INIT('h2)
	) name7325 (
		\u0_w_reg[2][11]/P0001 ,
		_w7313_,
		_w7857_
	);
	LUT2 #(
		.INIT('h4)
	) name7326 (
		\u0_w_reg[2][11]/P0001 ,
		_w7313_,
		_w7858_
	);
	LUT2 #(
		.INIT('h1)
	) name7327 (
		_w7857_,
		_w7858_,
		_w7859_
	);
	LUT2 #(
		.INIT('h8)
	) name7328 (
		_w7856_,
		_w7859_,
		_w7860_
	);
	LUT2 #(
		.INIT('h1)
	) name7329 (
		_w7856_,
		_w7859_,
		_w7861_
	);
	LUT2 #(
		.INIT('h1)
	) name7330 (
		_w7860_,
		_w7861_,
		_w7862_
	);
	LUT2 #(
		.INIT('h1)
	) name7331 (
		_w7781_,
		_w7862_,
		_w7863_
	);
	LUT2 #(
		.INIT('h8)
	) name7332 (
		_w7781_,
		_w7862_,
		_w7864_
	);
	LUT2 #(
		.INIT('h1)
	) name7333 (
		\ld_r_reg/P0001 ,
		_w7863_,
		_w7865_
	);
	LUT2 #(
		.INIT('h4)
	) name7334 (
		_w7864_,
		_w7865_,
		_w7866_
	);
	LUT2 #(
		.INIT('h2)
	) name7335 (
		\text_in_r_reg[43]/P0001 ,
		\u0_w_reg[2][11]/P0001 ,
		_w7867_
	);
	LUT2 #(
		.INIT('h4)
	) name7336 (
		\text_in_r_reg[43]/P0001 ,
		\u0_w_reg[2][11]/P0001 ,
		_w7868_
	);
	LUT2 #(
		.INIT('h2)
	) name7337 (
		\ld_r_reg/P0001 ,
		_w7867_,
		_w7869_
	);
	LUT2 #(
		.INIT('h4)
	) name7338 (
		_w7868_,
		_w7869_,
		_w7870_
	);
	LUT2 #(
		.INIT('h1)
	) name7339 (
		_w7866_,
		_w7870_,
		_w7871_
	);
	LUT2 #(
		.INIT('h2)
	) name7340 (
		\u0_w_reg[2][26]/P0001 ,
		_w7853_,
		_w7872_
	);
	LUT2 #(
		.INIT('h4)
	) name7341 (
		\u0_w_reg[2][26]/P0001 ,
		_w7853_,
		_w7873_
	);
	LUT2 #(
		.INIT('h1)
	) name7342 (
		_w7872_,
		_w7873_,
		_w7874_
	);
	LUT2 #(
		.INIT('h8)
	) name7343 (
		_w7760_,
		_w7874_,
		_w7875_
	);
	LUT2 #(
		.INIT('h1)
	) name7344 (
		_w7760_,
		_w7874_,
		_w7876_
	);
	LUT2 #(
		.INIT('h1)
	) name7345 (
		_w7875_,
		_w7876_,
		_w7877_
	);
	LUT2 #(
		.INIT('h4)
	) name7346 (
		_w6395_,
		_w7877_,
		_w7878_
	);
	LUT2 #(
		.INIT('h2)
	) name7347 (
		_w6395_,
		_w7877_,
		_w7879_
	);
	LUT2 #(
		.INIT('h1)
	) name7348 (
		\ld_r_reg/P0001 ,
		_w7878_,
		_w7880_
	);
	LUT2 #(
		.INIT('h4)
	) name7349 (
		_w7879_,
		_w7880_,
		_w7881_
	);
	LUT2 #(
		.INIT('h1)
	) name7350 (
		\text_in_r_reg[58]/P0001 ,
		\u0_w_reg[2][26]/P0001 ,
		_w7882_
	);
	LUT2 #(
		.INIT('h8)
	) name7351 (
		\text_in_r_reg[58]/P0001 ,
		\u0_w_reg[2][26]/P0001 ,
		_w7883_
	);
	LUT2 #(
		.INIT('h2)
	) name7352 (
		\ld_r_reg/P0001 ,
		_w7882_,
		_w7884_
	);
	LUT2 #(
		.INIT('h4)
	) name7353 (
		_w7883_,
		_w7884_,
		_w7885_
	);
	LUT2 #(
		.INIT('h1)
	) name7354 (
		_w7881_,
		_w7885_,
		_w7886_
	);
	LUT2 #(
		.INIT('h2)
	) name7355 (
		_w5417_,
		_w7580_,
		_w7887_
	);
	LUT2 #(
		.INIT('h4)
	) name7356 (
		_w5417_,
		_w7580_,
		_w7888_
	);
	LUT2 #(
		.INIT('h1)
	) name7357 (
		_w7887_,
		_w7888_,
		_w7889_
	);
	LUT2 #(
		.INIT('h8)
	) name7358 (
		_w7118_,
		_w7889_,
		_w7890_
	);
	LUT2 #(
		.INIT('h1)
	) name7359 (
		_w7118_,
		_w7889_,
		_w7891_
	);
	LUT2 #(
		.INIT('h1)
	) name7360 (
		_w7890_,
		_w7891_,
		_w7892_
	);
	LUT2 #(
		.INIT('h2)
	) name7361 (
		\u0_w_reg[2][3]/P0001 ,
		_w7206_,
		_w7893_
	);
	LUT2 #(
		.INIT('h4)
	) name7362 (
		\u0_w_reg[2][3]/P0001 ,
		_w7206_,
		_w7894_
	);
	LUT2 #(
		.INIT('h1)
	) name7363 (
		_w7893_,
		_w7894_,
		_w7895_
	);
	LUT2 #(
		.INIT('h8)
	) name7364 (
		_w7856_,
		_w7895_,
		_w7896_
	);
	LUT2 #(
		.INIT('h1)
	) name7365 (
		_w7856_,
		_w7895_,
		_w7897_
	);
	LUT2 #(
		.INIT('h1)
	) name7366 (
		_w7896_,
		_w7897_,
		_w7898_
	);
	LUT2 #(
		.INIT('h1)
	) name7367 (
		_w7892_,
		_w7898_,
		_w7899_
	);
	LUT2 #(
		.INIT('h8)
	) name7368 (
		_w7892_,
		_w7898_,
		_w7900_
	);
	LUT2 #(
		.INIT('h1)
	) name7369 (
		\ld_r_reg/P0001 ,
		_w7899_,
		_w7901_
	);
	LUT2 #(
		.INIT('h4)
	) name7370 (
		_w7900_,
		_w7901_,
		_w7902_
	);
	LUT2 #(
		.INIT('h2)
	) name7371 (
		\text_in_r_reg[35]/P0001 ,
		\u0_w_reg[2][3]/P0001 ,
		_w7903_
	);
	LUT2 #(
		.INIT('h4)
	) name7372 (
		\text_in_r_reg[35]/P0001 ,
		\u0_w_reg[2][3]/P0001 ,
		_w7904_
	);
	LUT2 #(
		.INIT('h2)
	) name7373 (
		\ld_r_reg/P0001 ,
		_w7903_,
		_w7905_
	);
	LUT2 #(
		.INIT('h4)
	) name7374 (
		_w7904_,
		_w7905_,
		_w7906_
	);
	LUT2 #(
		.INIT('h1)
	) name7375 (
		_w7902_,
		_w7906_,
		_w7907_
	);
	LUT2 #(
		.INIT('h2)
	) name7376 (
		\u0_w_reg[2][31]/P0001 ,
		_w5516_,
		_w7908_
	);
	LUT2 #(
		.INIT('h4)
	) name7377 (
		\u0_w_reg[2][31]/P0001 ,
		_w5516_,
		_w7909_
	);
	LUT2 #(
		.INIT('h1)
	) name7378 (
		_w7908_,
		_w7909_,
		_w7910_
	);
	LUT2 #(
		.INIT('h2)
	) name7379 (
		_w5631_,
		_w6657_,
		_w7911_
	);
	LUT2 #(
		.INIT('h4)
	) name7380 (
		_w5631_,
		_w6657_,
		_w7912_
	);
	LUT2 #(
		.INIT('h1)
	) name7381 (
		_w7911_,
		_w7912_,
		_w7913_
	);
	LUT2 #(
		.INIT('h8)
	) name7382 (
		_w5194_,
		_w7913_,
		_w7914_
	);
	LUT2 #(
		.INIT('h1)
	) name7383 (
		_w5194_,
		_w7913_,
		_w7915_
	);
	LUT2 #(
		.INIT('h1)
	) name7384 (
		_w7914_,
		_w7915_,
		_w7916_
	);
	LUT2 #(
		.INIT('h4)
	) name7385 (
		_w7910_,
		_w7916_,
		_w7917_
	);
	LUT2 #(
		.INIT('h2)
	) name7386 (
		_w7910_,
		_w7916_,
		_w7918_
	);
	LUT2 #(
		.INIT('h1)
	) name7387 (
		\ld_r_reg/P0001 ,
		_w7917_,
		_w7919_
	);
	LUT2 #(
		.INIT('h4)
	) name7388 (
		_w7918_,
		_w7919_,
		_w7920_
	);
	LUT2 #(
		.INIT('h2)
	) name7389 (
		\text_in_r_reg[63]/P0001 ,
		\u0_w_reg[2][31]/P0001 ,
		_w7921_
	);
	LUT2 #(
		.INIT('h4)
	) name7390 (
		\text_in_r_reg[63]/P0001 ,
		\u0_w_reg[2][31]/P0001 ,
		_w7922_
	);
	LUT2 #(
		.INIT('h2)
	) name7391 (
		\ld_r_reg/P0001 ,
		_w7921_,
		_w7923_
	);
	LUT2 #(
		.INIT('h4)
	) name7392 (
		_w7922_,
		_w7923_,
		_w7924_
	);
	LUT2 #(
		.INIT('h1)
	) name7393 (
		_w7920_,
		_w7924_,
		_w7925_
	);
	LUT2 #(
		.INIT('h1)
	) name7394 (
		\u0_w_reg[2][24]/P0001 ,
		_w6568_,
		_w7926_
	);
	LUT2 #(
		.INIT('h8)
	) name7395 (
		\u0_w_reg[2][24]/P0001 ,
		_w6568_,
		_w7927_
	);
	LUT2 #(
		.INIT('h1)
	) name7396 (
		_w7926_,
		_w7927_,
		_w7928_
	);
	LUT2 #(
		.INIT('h2)
	) name7397 (
		_w6927_,
		_w7408_,
		_w7929_
	);
	LUT2 #(
		.INIT('h4)
	) name7398 (
		_w6927_,
		_w7408_,
		_w7930_
	);
	LUT2 #(
		.INIT('h1)
	) name7399 (
		_w7929_,
		_w7930_,
		_w7931_
	);
	LUT2 #(
		.INIT('h4)
	) name7400 (
		_w5519_,
		_w7931_,
		_w7932_
	);
	LUT2 #(
		.INIT('h2)
	) name7401 (
		_w5519_,
		_w7931_,
		_w7933_
	);
	LUT2 #(
		.INIT('h1)
	) name7402 (
		_w7932_,
		_w7933_,
		_w7934_
	);
	LUT2 #(
		.INIT('h1)
	) name7403 (
		_w7928_,
		_w7934_,
		_w7935_
	);
	LUT2 #(
		.INIT('h8)
	) name7404 (
		_w7928_,
		_w7934_,
		_w7936_
	);
	LUT2 #(
		.INIT('h1)
	) name7405 (
		\ld_r_reg/P0001 ,
		_w7935_,
		_w7937_
	);
	LUT2 #(
		.INIT('h4)
	) name7406 (
		_w7936_,
		_w7937_,
		_w7938_
	);
	LUT2 #(
		.INIT('h1)
	) name7407 (
		\text_in_r_reg[56]/P0001 ,
		\u0_w_reg[2][24]/P0001 ,
		_w7939_
	);
	LUT2 #(
		.INIT('h8)
	) name7408 (
		\text_in_r_reg[56]/P0001 ,
		\u0_w_reg[2][24]/P0001 ,
		_w7940_
	);
	LUT2 #(
		.INIT('h2)
	) name7409 (
		\ld_r_reg/P0001 ,
		_w7939_,
		_w7941_
	);
	LUT2 #(
		.INIT('h4)
	) name7410 (
		_w7940_,
		_w7941_,
		_w7942_
	);
	LUT2 #(
		.INIT('h1)
	) name7411 (
		_w7938_,
		_w7942_,
		_w7943_
	);
	LUT2 #(
		.INIT('h1)
	) name7412 (
		\u0_w_reg[2][16]/P0001 ,
		_w6568_,
		_w7944_
	);
	LUT2 #(
		.INIT('h8)
	) name7413 (
		\u0_w_reg[2][16]/P0001 ,
		_w6568_,
		_w7945_
	);
	LUT2 #(
		.INIT('h1)
	) name7414 (
		_w7944_,
		_w7945_,
		_w7946_
	);
	LUT2 #(
		.INIT('h2)
	) name7415 (
		_w5516_,
		_w6472_,
		_w7947_
	);
	LUT2 #(
		.INIT('h4)
	) name7416 (
		_w5516_,
		_w6472_,
		_w7948_
	);
	LUT2 #(
		.INIT('h1)
	) name7417 (
		_w7947_,
		_w7948_,
		_w7949_
	);
	LUT2 #(
		.INIT('h8)
	) name7418 (
		_w6930_,
		_w7949_,
		_w7950_
	);
	LUT2 #(
		.INIT('h1)
	) name7419 (
		_w6930_,
		_w7949_,
		_w7951_
	);
	LUT2 #(
		.INIT('h1)
	) name7420 (
		_w7950_,
		_w7951_,
		_w7952_
	);
	LUT2 #(
		.INIT('h4)
	) name7421 (
		_w7946_,
		_w7952_,
		_w7953_
	);
	LUT2 #(
		.INIT('h2)
	) name7422 (
		_w7946_,
		_w7952_,
		_w7954_
	);
	LUT2 #(
		.INIT('h1)
	) name7423 (
		\ld_r_reg/P0001 ,
		_w7953_,
		_w7955_
	);
	LUT2 #(
		.INIT('h4)
	) name7424 (
		_w7954_,
		_w7955_,
		_w7956_
	);
	LUT2 #(
		.INIT('h1)
	) name7425 (
		\text_in_r_reg[48]/P0001 ,
		\u0_w_reg[2][16]/P0001 ,
		_w7957_
	);
	LUT2 #(
		.INIT('h8)
	) name7426 (
		\text_in_r_reg[48]/P0001 ,
		\u0_w_reg[2][16]/P0001 ,
		_w7958_
	);
	LUT2 #(
		.INIT('h2)
	) name7427 (
		\ld_r_reg/P0001 ,
		_w7957_,
		_w7959_
	);
	LUT2 #(
		.INIT('h4)
	) name7428 (
		_w7958_,
		_w7959_,
		_w7960_
	);
	LUT2 #(
		.INIT('h1)
	) name7429 (
		_w7956_,
		_w7960_,
		_w7961_
	);
	LUT2 #(
		.INIT('h1)
	) name7430 (
		_w7580_,
		_w7673_,
		_w7962_
	);
	LUT2 #(
		.INIT('h8)
	) name7431 (
		_w7580_,
		_w7673_,
		_w7963_
	);
	LUT2 #(
		.INIT('h1)
	) name7432 (
		_w7962_,
		_w7963_,
		_w7964_
	);
	LUT2 #(
		.INIT('h2)
	) name7433 (
		\u0_w_reg[2][18]/P0001 ,
		_w7853_,
		_w7965_
	);
	LUT2 #(
		.INIT('h4)
	) name7434 (
		\u0_w_reg[2][18]/P0001 ,
		_w7853_,
		_w7966_
	);
	LUT2 #(
		.INIT('h1)
	) name7435 (
		_w7965_,
		_w7966_,
		_w7967_
	);
	LUT2 #(
		.INIT('h8)
	) name7436 (
		_w7655_,
		_w7967_,
		_w7968_
	);
	LUT2 #(
		.INIT('h1)
	) name7437 (
		_w7655_,
		_w7967_,
		_w7969_
	);
	LUT2 #(
		.INIT('h1)
	) name7438 (
		_w7968_,
		_w7969_,
		_w7970_
	);
	LUT2 #(
		.INIT('h1)
	) name7439 (
		_w7964_,
		_w7970_,
		_w7971_
	);
	LUT2 #(
		.INIT('h8)
	) name7440 (
		_w7964_,
		_w7970_,
		_w7972_
	);
	LUT2 #(
		.INIT('h1)
	) name7441 (
		\ld_r_reg/P0001 ,
		_w7971_,
		_w7973_
	);
	LUT2 #(
		.INIT('h4)
	) name7442 (
		_w7972_,
		_w7973_,
		_w7974_
	);
	LUT2 #(
		.INIT('h2)
	) name7443 (
		\text_in_r_reg[50]/P0001 ,
		\u0_w_reg[2][18]/P0001 ,
		_w7975_
	);
	LUT2 #(
		.INIT('h4)
	) name7444 (
		\text_in_r_reg[50]/P0001 ,
		\u0_w_reg[2][18]/P0001 ,
		_w7976_
	);
	LUT2 #(
		.INIT('h2)
	) name7445 (
		\ld_r_reg/P0001 ,
		_w7975_,
		_w7977_
	);
	LUT2 #(
		.INIT('h4)
	) name7446 (
		_w7976_,
		_w7977_,
		_w7978_
	);
	LUT2 #(
		.INIT('h1)
	) name7447 (
		_w7974_,
		_w7978_,
		_w7979_
	);
	LUT2 #(
		.INIT('h1)
	) name7448 (
		_w853_,
		_w5417_,
		_w7980_
	);
	LUT2 #(
		.INIT('h8)
	) name7449 (
		_w853_,
		_w5417_,
		_w7981_
	);
	LUT2 #(
		.INIT('h1)
	) name7450 (
		_w7980_,
		_w7981_,
		_w7982_
	);
	LUT2 #(
		.INIT('h1)
	) name7451 (
		\u0_w_reg[2][23]/P0001 ,
		_w7913_,
		_w7983_
	);
	LUT2 #(
		.INIT('h8)
	) name7452 (
		\u0_w_reg[2][23]/P0001 ,
		_w7913_,
		_w7984_
	);
	LUT2 #(
		.INIT('h1)
	) name7453 (
		_w7983_,
		_w7984_,
		_w7985_
	);
	LUT2 #(
		.INIT('h1)
	) name7454 (
		_w7982_,
		_w7985_,
		_w7986_
	);
	LUT2 #(
		.INIT('h8)
	) name7455 (
		_w7982_,
		_w7985_,
		_w7987_
	);
	LUT2 #(
		.INIT('h1)
	) name7456 (
		\ld_r_reg/P0001 ,
		_w7986_,
		_w7988_
	);
	LUT2 #(
		.INIT('h4)
	) name7457 (
		_w7987_,
		_w7988_,
		_w7989_
	);
	LUT2 #(
		.INIT('h2)
	) name7458 (
		\text_in_r_reg[55]/P0001 ,
		\u0_w_reg[2][23]/P0001 ,
		_w7990_
	);
	LUT2 #(
		.INIT('h4)
	) name7459 (
		\text_in_r_reg[55]/P0001 ,
		\u0_w_reg[2][23]/P0001 ,
		_w7991_
	);
	LUT2 #(
		.INIT('h2)
	) name7460 (
		\ld_r_reg/P0001 ,
		_w7990_,
		_w7992_
	);
	LUT2 #(
		.INIT('h4)
	) name7461 (
		_w7991_,
		_w7992_,
		_w7993_
	);
	LUT2 #(
		.INIT('h1)
	) name7462 (
		_w7989_,
		_w7993_,
		_w7994_
	);
	LUT2 #(
		.INIT('h1)
	) name7463 (
		\u0_w_reg[2][8]/P0001 ,
		_w6568_,
		_w7995_
	);
	LUT2 #(
		.INIT('h8)
	) name7464 (
		\u0_w_reg[2][8]/P0001 ,
		_w6568_,
		_w7996_
	);
	LUT2 #(
		.INIT('h1)
	) name7465 (
		_w7995_,
		_w7996_,
		_w7997_
	);
	LUT2 #(
		.INIT('h2)
	) name7466 (
		_w6472_,
		_w7408_,
		_w7998_
	);
	LUT2 #(
		.INIT('h4)
	) name7467 (
		_w6472_,
		_w7408_,
		_w7999_
	);
	LUT2 #(
		.INIT('h1)
	) name7468 (
		_w7998_,
		_w7999_,
		_w8000_
	);
	LUT2 #(
		.INIT('h8)
	) name7469 (
		_w7913_,
		_w8000_,
		_w8001_
	);
	LUT2 #(
		.INIT('h1)
	) name7470 (
		_w7913_,
		_w8000_,
		_w8002_
	);
	LUT2 #(
		.INIT('h1)
	) name7471 (
		_w8001_,
		_w8002_,
		_w8003_
	);
	LUT2 #(
		.INIT('h1)
	) name7472 (
		_w7997_,
		_w8003_,
		_w8004_
	);
	LUT2 #(
		.INIT('h8)
	) name7473 (
		_w7997_,
		_w8003_,
		_w8005_
	);
	LUT2 #(
		.INIT('h1)
	) name7474 (
		\ld_r_reg/P0001 ,
		_w8004_,
		_w8006_
	);
	LUT2 #(
		.INIT('h4)
	) name7475 (
		_w8005_,
		_w8006_,
		_w8007_
	);
	LUT2 #(
		.INIT('h2)
	) name7476 (
		\text_in_r_reg[40]/P0001 ,
		\u0_w_reg[2][8]/P0001 ,
		_w8008_
	);
	LUT2 #(
		.INIT('h4)
	) name7477 (
		\text_in_r_reg[40]/P0001 ,
		\u0_w_reg[2][8]/P0001 ,
		_w8009_
	);
	LUT2 #(
		.INIT('h2)
	) name7478 (
		\ld_r_reg/P0001 ,
		_w8008_,
		_w8010_
	);
	LUT2 #(
		.INIT('h4)
	) name7479 (
		_w8009_,
		_w8010_,
		_w8011_
	);
	LUT2 #(
		.INIT('h1)
	) name7480 (
		_w8007_,
		_w8011_,
		_w8012_
	);
	LUT2 #(
		.INIT('h1)
	) name7481 (
		_w6743_,
		_w7583_,
		_w8013_
	);
	LUT2 #(
		.INIT('h8)
	) name7482 (
		_w6743_,
		_w7583_,
		_w8014_
	);
	LUT2 #(
		.INIT('h1)
	) name7483 (
		_w8013_,
		_w8014_,
		_w8015_
	);
	LUT2 #(
		.INIT('h2)
	) name7484 (
		\u0_w_reg[2][10]/P0001 ,
		_w7853_,
		_w8016_
	);
	LUT2 #(
		.INIT('h4)
	) name7485 (
		\u0_w_reg[2][10]/P0001 ,
		_w7853_,
		_w8017_
	);
	LUT2 #(
		.INIT('h1)
	) name7486 (
		_w8016_,
		_w8017_,
		_w8018_
	);
	LUT2 #(
		.INIT('h8)
	) name7487 (
		_w6842_,
		_w8018_,
		_w8019_
	);
	LUT2 #(
		.INIT('h1)
	) name7488 (
		_w6842_,
		_w8018_,
		_w8020_
	);
	LUT2 #(
		.INIT('h1)
	) name7489 (
		_w8019_,
		_w8020_,
		_w8021_
	);
	LUT2 #(
		.INIT('h1)
	) name7490 (
		_w8015_,
		_w8021_,
		_w8022_
	);
	LUT2 #(
		.INIT('h8)
	) name7491 (
		_w8015_,
		_w8021_,
		_w8023_
	);
	LUT2 #(
		.INIT('h1)
	) name7492 (
		\ld_r_reg/P0001 ,
		_w8022_,
		_w8024_
	);
	LUT2 #(
		.INIT('h4)
	) name7493 (
		_w8023_,
		_w8024_,
		_w8025_
	);
	LUT2 #(
		.INIT('h2)
	) name7494 (
		\text_in_r_reg[42]/P0001 ,
		\u0_w_reg[2][10]/P0001 ,
		_w8026_
	);
	LUT2 #(
		.INIT('h4)
	) name7495 (
		\text_in_r_reg[42]/P0001 ,
		\u0_w_reg[2][10]/P0001 ,
		_w8027_
	);
	LUT2 #(
		.INIT('h2)
	) name7496 (
		\ld_r_reg/P0001 ,
		_w8026_,
		_w8028_
	);
	LUT2 #(
		.INIT('h4)
	) name7497 (
		_w8027_,
		_w8028_,
		_w8029_
	);
	LUT2 #(
		.INIT('h1)
	) name7498 (
		_w8025_,
		_w8029_,
		_w8030_
	);
	LUT2 #(
		.INIT('h1)
	) name7499 (
		\u0_w_reg[2][5]/P0001 ,
		_w5307_,
		_w8031_
	);
	LUT2 #(
		.INIT('h8)
	) name7500 (
		\u0_w_reg[2][5]/P0001 ,
		_w5307_,
		_w8032_
	);
	LUT2 #(
		.INIT('h1)
	) name7501 (
		_w8031_,
		_w8032_,
		_w8033_
	);
	LUT2 #(
		.INIT('h1)
	) name7502 (
		\u0_w_reg[2][6]/P0001 ,
		_w1300_,
		_w8034_
	);
	LUT2 #(
		.INIT('h8)
	) name7503 (
		\u0_w_reg[2][6]/P0001 ,
		_w1300_,
		_w8035_
	);
	LUT2 #(
		.INIT('h1)
	) name7504 (
		_w8034_,
		_w8035_,
		_w8036_
	);
	LUT2 #(
		.INIT('h1)
	) name7505 (
		\u0_w_reg[2][4]/P0001 ,
		_w6180_,
		_w8037_
	);
	LUT2 #(
		.INIT('h8)
	) name7506 (
		\u0_w_reg[2][4]/P0001 ,
		_w6180_,
		_w8038_
	);
	LUT2 #(
		.INIT('h1)
	) name7507 (
		_w8037_,
		_w8038_,
		_w8039_
	);
	LUT2 #(
		.INIT('h1)
	) name7508 (
		\u0_w_reg[2][0]/P0001 ,
		_w6568_,
		_w8040_
	);
	LUT2 #(
		.INIT('h8)
	) name7509 (
		\u0_w_reg[2][0]/P0001 ,
		_w6568_,
		_w8041_
	);
	LUT2 #(
		.INIT('h1)
	) name7510 (
		_w8040_,
		_w8041_,
		_w8042_
	);
	LUT2 #(
		.INIT('h1)
	) name7511 (
		\u0_w_reg[2][3]/P0001 ,
		_w7313_,
		_w8043_
	);
	LUT2 #(
		.INIT('h8)
	) name7512 (
		\u0_w_reg[2][3]/P0001 ,
		_w7313_,
		_w8044_
	);
	LUT2 #(
		.INIT('h1)
	) name7513 (
		_w8043_,
		_w8044_,
		_w8045_
	);
	LUT2 #(
		.INIT('h1)
	) name7514 (
		\u0_w_reg[2][1]/P0001 ,
		_w6842_,
		_w8046_
	);
	LUT2 #(
		.INIT('h8)
	) name7515 (
		\u0_w_reg[2][1]/P0001 ,
		_w6842_,
		_w8047_
	);
	LUT2 #(
		.INIT('h1)
	) name7516 (
		_w8046_,
		_w8047_,
		_w8048_
	);
	LUT2 #(
		.INIT('h1)
	) name7517 (
		\u0_w_reg[2][2]/P0001 ,
		_w7853_,
		_w8049_
	);
	LUT2 #(
		.INIT('h8)
	) name7518 (
		\u0_w_reg[2][2]/P0001 ,
		_w7853_,
		_w8050_
	);
	LUT2 #(
		.INIT('h1)
	) name7519 (
		_w8049_,
		_w8050_,
		_w8051_
	);
	LUT2 #(
		.INIT('h1)
	) name7520 (
		\u0_w_reg[2][7]/P0001 ,
		_w6657_,
		_w8052_
	);
	LUT2 #(
		.INIT('h8)
	) name7521 (
		\u0_w_reg[2][7]/P0001 ,
		_w6657_,
		_w8053_
	);
	LUT2 #(
		.INIT('h1)
	) name7522 (
		_w8052_,
		_w8053_,
		_w8054_
	);
	LUT2 #(
		.INIT('h1)
	) name7523 (
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w8055_
	);
	LUT2 #(
		.INIT('h8)
	) name7524 (
		\sa12_reg[5]/P0001 ,
		_w8055_,
		_w8056_
	);
	LUT2 #(
		.INIT('h8)
	) name7525 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		_w8057_
	);
	LUT2 #(
		.INIT('h8)
	) name7526 (
		_w8056_,
		_w8057_,
		_w8058_
	);
	LUT2 #(
		.INIT('h2)
	) name7527 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		_w8059_
	);
	LUT2 #(
		.INIT('h2)
	) name7528 (
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w8060_
	);
	LUT2 #(
		.INIT('h8)
	) name7529 (
		\sa12_reg[4]/P0001 ,
		_w8060_,
		_w8061_
	);
	LUT2 #(
		.INIT('h8)
	) name7530 (
		_w8059_,
		_w8061_,
		_w8062_
	);
	LUT2 #(
		.INIT('h1)
	) name7531 (
		_w8058_,
		_w8062_,
		_w8063_
	);
	LUT2 #(
		.INIT('h2)
	) name7532 (
		\sa12_reg[1]/P0001 ,
		_w8063_,
		_w8064_
	);
	LUT2 #(
		.INIT('h8)
	) name7533 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w8065_
	);
	LUT2 #(
		.INIT('h8)
	) name7534 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w8066_
	);
	LUT2 #(
		.INIT('h8)
	) name7535 (
		_w8065_,
		_w8066_,
		_w8067_
	);
	LUT2 #(
		.INIT('h4)
	) name7536 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w8068_
	);
	LUT2 #(
		.INIT('h1)
	) name7537 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w8069_
	);
	LUT2 #(
		.INIT('h8)
	) name7538 (
		_w8068_,
		_w8069_,
		_w8070_
	);
	LUT2 #(
		.INIT('h4)
	) name7539 (
		\sa12_reg[2]/P0001 ,
		_w8070_,
		_w8071_
	);
	LUT2 #(
		.INIT('h1)
	) name7540 (
		_w8067_,
		_w8071_,
		_w8072_
	);
	LUT2 #(
		.INIT('h2)
	) name7541 (
		\sa12_reg[3]/P0001 ,
		_w8072_,
		_w8073_
	);
	LUT2 #(
		.INIT('h2)
	) name7542 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w8074_
	);
	LUT2 #(
		.INIT('h8)
	) name7543 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w8075_
	);
	LUT2 #(
		.INIT('h8)
	) name7544 (
		_w8074_,
		_w8075_,
		_w8076_
	);
	LUT2 #(
		.INIT('h2)
	) name7545 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w8077_
	);
	LUT2 #(
		.INIT('h2)
	) name7546 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w8078_
	);
	LUT2 #(
		.INIT('h8)
	) name7547 (
		_w8077_,
		_w8078_,
		_w8079_
	);
	LUT2 #(
		.INIT('h8)
	) name7548 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w8080_
	);
	LUT2 #(
		.INIT('h8)
	) name7549 (
		\sa12_reg[3]/P0001 ,
		_w8080_,
		_w8081_
	);
	LUT2 #(
		.INIT('h1)
	) name7550 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w8082_
	);
	LUT2 #(
		.INIT('h8)
	) name7551 (
		_w8081_,
		_w8082_,
		_w8083_
	);
	LUT2 #(
		.INIT('h4)
	) name7552 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w8084_
	);
	LUT2 #(
		.INIT('h4)
	) name7553 (
		\sa12_reg[4]/P0001 ,
		_w8084_,
		_w8085_
	);
	LUT2 #(
		.INIT('h8)
	) name7554 (
		_w8082_,
		_w8085_,
		_w8086_
	);
	LUT2 #(
		.INIT('h4)
	) name7555 (
		\sa12_reg[3]/P0001 ,
		_w8056_,
		_w8087_
	);
	LUT2 #(
		.INIT('h2)
	) name7556 (
		\sa12_reg[2]/P0001 ,
		_w8076_,
		_w8088_
	);
	LUT2 #(
		.INIT('h4)
	) name7557 (
		_w8079_,
		_w8088_,
		_w8089_
	);
	LUT2 #(
		.INIT('h1)
	) name7558 (
		_w8083_,
		_w8086_,
		_w8090_
	);
	LUT2 #(
		.INIT('h4)
	) name7559 (
		_w8087_,
		_w8090_,
		_w8091_
	);
	LUT2 #(
		.INIT('h8)
	) name7560 (
		_w8089_,
		_w8091_,
		_w8092_
	);
	LUT2 #(
		.INIT('h4)
	) name7561 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w8093_
	);
	LUT2 #(
		.INIT('h4)
	) name7562 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w8094_
	);
	LUT2 #(
		.INIT('h8)
	) name7563 (
		_w8093_,
		_w8094_,
		_w8095_
	);
	LUT2 #(
		.INIT('h8)
	) name7564 (
		_w8084_,
		_w8093_,
		_w8096_
	);
	LUT2 #(
		.INIT('h8)
	) name7565 (
		_w8065_,
		_w8078_,
		_w8097_
	);
	LUT2 #(
		.INIT('h8)
	) name7566 (
		\sa12_reg[7]/NET0131 ,
		_w8097_,
		_w8098_
	);
	LUT2 #(
		.INIT('h1)
	) name7567 (
		\sa12_reg[2]/P0001 ,
		_w8095_,
		_w8099_
	);
	LUT2 #(
		.INIT('h4)
	) name7568 (
		_w8096_,
		_w8099_,
		_w8100_
	);
	LUT2 #(
		.INIT('h4)
	) name7569 (
		_w8098_,
		_w8100_,
		_w8101_
	);
	LUT2 #(
		.INIT('h1)
	) name7570 (
		_w8092_,
		_w8101_,
		_w8102_
	);
	LUT2 #(
		.INIT('h8)
	) name7571 (
		\sa12_reg[4]/P0001 ,
		_w8076_,
		_w8103_
	);
	LUT2 #(
		.INIT('h1)
	) name7572 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w8104_
	);
	LUT2 #(
		.INIT('h8)
	) name7573 (
		_w8056_,
		_w8104_,
		_w8105_
	);
	LUT2 #(
		.INIT('h1)
	) name7574 (
		\sa12_reg[1]/P0001 ,
		_w8103_,
		_w8106_
	);
	LUT2 #(
		.INIT('h4)
	) name7575 (
		_w8105_,
		_w8106_,
		_w8107_
	);
	LUT2 #(
		.INIT('h4)
	) name7576 (
		_w8102_,
		_w8107_,
		_w8108_
	);
	LUT2 #(
		.INIT('h8)
	) name7577 (
		_w8081_,
		_w8093_,
		_w8109_
	);
	LUT2 #(
		.INIT('h2)
	) name7578 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		_w8110_
	);
	LUT2 #(
		.INIT('h4)
	) name7579 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w8111_
	);
	LUT2 #(
		.INIT('h8)
	) name7580 (
		_w8110_,
		_w8111_,
		_w8112_
	);
	LUT2 #(
		.INIT('h4)
	) name7581 (
		\sa12_reg[6]/NET0131 ,
		_w8112_,
		_w8113_
	);
	LUT2 #(
		.INIT('h8)
	) name7582 (
		_w8065_,
		_w8084_,
		_w8114_
	);
	LUT2 #(
		.INIT('h4)
	) name7583 (
		\sa12_reg[4]/P0001 ,
		_w8114_,
		_w8115_
	);
	LUT2 #(
		.INIT('h4)
	) name7584 (
		_w8055_,
		_w8110_,
		_w8116_
	);
	LUT2 #(
		.INIT('h8)
	) name7585 (
		_w8082_,
		_w8104_,
		_w8117_
	);
	LUT2 #(
		.INIT('h4)
	) name7586 (
		\sa12_reg[7]/NET0131 ,
		_w8117_,
		_w8118_
	);
	LUT2 #(
		.INIT('h1)
	) name7587 (
		_w8115_,
		_w8116_,
		_w8119_
	);
	LUT2 #(
		.INIT('h4)
	) name7588 (
		_w8118_,
		_w8119_,
		_w8120_
	);
	LUT2 #(
		.INIT('h1)
	) name7589 (
		\sa12_reg[2]/P0001 ,
		_w8120_,
		_w8121_
	);
	LUT2 #(
		.INIT('h2)
	) name7590 (
		\sa12_reg[1]/P0001 ,
		_w8109_,
		_w8122_
	);
	LUT2 #(
		.INIT('h4)
	) name7591 (
		_w8113_,
		_w8122_,
		_w8123_
	);
	LUT2 #(
		.INIT('h4)
	) name7592 (
		_w8121_,
		_w8123_,
		_w8124_
	);
	LUT2 #(
		.INIT('h1)
	) name7593 (
		_w8108_,
		_w8124_,
		_w8125_
	);
	LUT2 #(
		.INIT('h4)
	) name7594 (
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w8126_
	);
	LUT2 #(
		.INIT('h8)
	) name7595 (
		_w8110_,
		_w8126_,
		_w8127_
	);
	LUT2 #(
		.INIT('h2)
	) name7596 (
		\sa12_reg[2]/P0001 ,
		_w8127_,
		_w8128_
	);
	LUT2 #(
		.INIT('h4)
	) name7597 (
		\sa12_reg[6]/NET0131 ,
		_w8078_,
		_w8129_
	);
	LUT2 #(
		.INIT('h8)
	) name7598 (
		\sa12_reg[7]/NET0131 ,
		_w8065_,
		_w8130_
	);
	LUT2 #(
		.INIT('h1)
	) name7599 (
		_w8094_,
		_w8130_,
		_w8131_
	);
	LUT2 #(
		.INIT('h1)
	) name7600 (
		_w8080_,
		_w8131_,
		_w8132_
	);
	LUT2 #(
		.INIT('h2)
	) name7601 (
		_w8128_,
		_w8129_,
		_w8133_
	);
	LUT2 #(
		.INIT('h4)
	) name7602 (
		_w8132_,
		_w8133_,
		_w8134_
	);
	LUT2 #(
		.INIT('h4)
	) name7603 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w8135_
	);
	LUT2 #(
		.INIT('h8)
	) name7604 (
		_w8075_,
		_w8135_,
		_w8136_
	);
	LUT2 #(
		.INIT('h1)
	) name7605 (
		\sa12_reg[2]/P0001 ,
		_w8136_,
		_w8137_
	);
	LUT2 #(
		.INIT('h8)
	) name7606 (
		_w8060_,
		_w8078_,
		_w8138_
	);
	LUT2 #(
		.INIT('h1)
	) name7607 (
		_w8118_,
		_w8138_,
		_w8139_
	);
	LUT2 #(
		.INIT('h8)
	) name7608 (
		_w8137_,
		_w8139_,
		_w8140_
	);
	LUT2 #(
		.INIT('h1)
	) name7609 (
		_w8134_,
		_w8140_,
		_w8141_
	);
	LUT2 #(
		.INIT('h4)
	) name7610 (
		\sa12_reg[7]/NET0131 ,
		_w8082_,
		_w8142_
	);
	LUT2 #(
		.INIT('h8)
	) name7611 (
		_w8094_,
		_w8142_,
		_w8143_
	);
	LUT2 #(
		.INIT('h2)
	) name7612 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w8144_
	);
	LUT2 #(
		.INIT('h8)
	) name7613 (
		_w8126_,
		_w8144_,
		_w8145_
	);
	LUT2 #(
		.INIT('h4)
	) name7614 (
		\sa12_reg[4]/P0001 ,
		_w8060_,
		_w8146_
	);
	LUT2 #(
		.INIT('h8)
	) name7615 (
		_w8080_,
		_w8082_,
		_w8147_
	);
	LUT2 #(
		.INIT('h1)
	) name7616 (
		_w8146_,
		_w8147_,
		_w8148_
	);
	LUT2 #(
		.INIT('h1)
	) name7617 (
		\sa12_reg[2]/P0001 ,
		_w8148_,
		_w8149_
	);
	LUT2 #(
		.INIT('h8)
	) name7618 (
		_w8074_,
		_w8129_,
		_w8150_
	);
	LUT2 #(
		.INIT('h2)
	) name7619 (
		\sa12_reg[1]/P0001 ,
		_w8145_,
		_w8151_
	);
	LUT2 #(
		.INIT('h4)
	) name7620 (
		_w8143_,
		_w8151_,
		_w8152_
	);
	LUT2 #(
		.INIT('h4)
	) name7621 (
		_w8150_,
		_w8152_,
		_w8153_
	);
	LUT2 #(
		.INIT('h4)
	) name7622 (
		_w8149_,
		_w8153_,
		_w8154_
	);
	LUT2 #(
		.INIT('h4)
	) name7623 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		_w8155_
	);
	LUT2 #(
		.INIT('h8)
	) name7624 (
		\sa12_reg[4]/P0001 ,
		_w8055_,
		_w8156_
	);
	LUT2 #(
		.INIT('h8)
	) name7625 (
		_w8155_,
		_w8156_,
		_w8157_
	);
	LUT2 #(
		.INIT('h1)
	) name7626 (
		\sa12_reg[1]/P0001 ,
		_w8157_,
		_w8158_
	);
	LUT2 #(
		.INIT('h8)
	) name7627 (
		\sa12_reg[7]/NET0131 ,
		_w8075_,
		_w8159_
	);
	LUT2 #(
		.INIT('h4)
	) name7628 (
		\sa12_reg[4]/P0001 ,
		_w8159_,
		_w8160_
	);
	LUT2 #(
		.INIT('h8)
	) name7629 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w8161_
	);
	LUT2 #(
		.INIT('h1)
	) name7630 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w8162_
	);
	LUT2 #(
		.INIT('h1)
	) name7631 (
		\sa12_reg[3]/P0001 ,
		_w8162_,
		_w8163_
	);
	LUT2 #(
		.INIT('h2)
	) name7632 (
		_w8161_,
		_w8163_,
		_w8164_
	);
	LUT2 #(
		.INIT('h8)
	) name7633 (
		\sa12_reg[4]/P0001 ,
		_w8161_,
		_w8165_
	);
	LUT2 #(
		.INIT('h4)
	) name7634 (
		\sa12_reg[6]/NET0131 ,
		_w8165_,
		_w8166_
	);
	LUT2 #(
		.INIT('h8)
	) name7635 (
		\sa12_reg[2]/P0001 ,
		_w8166_,
		_w8167_
	);
	LUT2 #(
		.INIT('h1)
	) name7636 (
		_w8160_,
		_w8164_,
		_w8168_
	);
	LUT2 #(
		.INIT('h8)
	) name7637 (
		_w8158_,
		_w8168_,
		_w8169_
	);
	LUT2 #(
		.INIT('h4)
	) name7638 (
		_w8167_,
		_w8169_,
		_w8170_
	);
	LUT2 #(
		.INIT('h1)
	) name7639 (
		_w8154_,
		_w8170_,
		_w8171_
	);
	LUT2 #(
		.INIT('h2)
	) name7640 (
		\sa12_reg[0]/P0001 ,
		_w8141_,
		_w8172_
	);
	LUT2 #(
		.INIT('h4)
	) name7641 (
		_w8171_,
		_w8172_,
		_w8173_
	);
	LUT2 #(
		.INIT('h8)
	) name7642 (
		\sa12_reg[5]/P0001 ,
		_w8060_,
		_w8174_
	);
	LUT2 #(
		.INIT('h4)
	) name7643 (
		\sa12_reg[3]/P0001 ,
		_w8174_,
		_w8175_
	);
	LUT2 #(
		.INIT('h4)
	) name7644 (
		\sa12_reg[1]/P0001 ,
		_w8175_,
		_w8176_
	);
	LUT2 #(
		.INIT('h8)
	) name7645 (
		\sa12_reg[7]/NET0131 ,
		_w8095_,
		_w8177_
	);
	LUT2 #(
		.INIT('h1)
	) name7646 (
		_w8176_,
		_w8177_,
		_w8178_
	);
	LUT2 #(
		.INIT('h1)
	) name7647 (
		\sa12_reg[2]/P0001 ,
		_w8178_,
		_w8179_
	);
	LUT2 #(
		.INIT('h8)
	) name7648 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w8180_
	);
	LUT2 #(
		.INIT('h8)
	) name7649 (
		_w8060_,
		_w8180_,
		_w8181_
	);
	LUT2 #(
		.INIT('h8)
	) name7650 (
		\sa12_reg[4]/P0001 ,
		_w8135_,
		_w8182_
	);
	LUT2 #(
		.INIT('h8)
	) name7651 (
		_w8059_,
		_w8182_,
		_w8183_
	);
	LUT2 #(
		.INIT('h8)
	) name7652 (
		_w8082_,
		_w8111_,
		_w8184_
	);
	LUT2 #(
		.INIT('h8)
	) name7653 (
		\sa12_reg[5]/P0001 ,
		_w8126_,
		_w8185_
	);
	LUT2 #(
		.INIT('h4)
	) name7654 (
		_w8078_,
		_w8185_,
		_w8186_
	);
	LUT2 #(
		.INIT('h1)
	) name7655 (
		_w8184_,
		_w8186_,
		_w8187_
	);
	LUT2 #(
		.INIT('h1)
	) name7656 (
		\sa12_reg[2]/P0001 ,
		_w8187_,
		_w8188_
	);
	LUT2 #(
		.INIT('h8)
	) name7657 (
		\sa12_reg[2]/P0001 ,
		_w8174_,
		_w8189_
	);
	LUT2 #(
		.INIT('h2)
	) name7658 (
		\sa12_reg[1]/P0001 ,
		_w8181_,
		_w8190_
	);
	LUT2 #(
		.INIT('h4)
	) name7659 (
		_w8183_,
		_w8190_,
		_w8191_
	);
	LUT2 #(
		.INIT('h4)
	) name7660 (
		_w8189_,
		_w8191_,
		_w8192_
	);
	LUT2 #(
		.INIT('h4)
	) name7661 (
		_w8188_,
		_w8192_,
		_w8193_
	);
	LUT2 #(
		.INIT('h8)
	) name7662 (
		\sa12_reg[2]/P0001 ,
		_w8142_,
		_w8194_
	);
	LUT2 #(
		.INIT('h4)
	) name7663 (
		\sa12_reg[7]/NET0131 ,
		_w8129_,
		_w8195_
	);
	LUT2 #(
		.INIT('h1)
	) name7664 (
		\sa12_reg[1]/P0001 ,
		_w8067_,
		_w8196_
	);
	LUT2 #(
		.INIT('h4)
	) name7665 (
		_w8194_,
		_w8196_,
		_w8197_
	);
	LUT2 #(
		.INIT('h4)
	) name7666 (
		_w8195_,
		_w8197_,
		_w8198_
	);
	LUT2 #(
		.INIT('h1)
	) name7667 (
		_w8193_,
		_w8198_,
		_w8199_
	);
	LUT2 #(
		.INIT('h8)
	) name7668 (
		_w8069_,
		_w8180_,
		_w8200_
	);
	LUT2 #(
		.INIT('h4)
	) name7669 (
		\sa12_reg[6]/NET0131 ,
		_w8200_,
		_w8201_
	);
	LUT2 #(
		.INIT('h4)
	) name7670 (
		\sa12_reg[4]/P0001 ,
		_w8093_,
		_w8202_
	);
	LUT2 #(
		.INIT('h4)
	) name7671 (
		\sa12_reg[3]/P0001 ,
		_w8202_,
		_w8203_
	);
	LUT2 #(
		.INIT('h1)
	) name7672 (
		_w8201_,
		_w8203_,
		_w8204_
	);
	LUT2 #(
		.INIT('h2)
	) name7673 (
		\sa12_reg[2]/P0001 ,
		_w8204_,
		_w8205_
	);
	LUT2 #(
		.INIT('h1)
	) name7674 (
		\sa12_reg[0]/P0001 ,
		_w8105_,
		_w8206_
	);
	LUT2 #(
		.INIT('h4)
	) name7675 (
		_w8205_,
		_w8206_,
		_w8207_
	);
	LUT2 #(
		.INIT('h4)
	) name7676 (
		_w8179_,
		_w8207_,
		_w8208_
	);
	LUT2 #(
		.INIT('h4)
	) name7677 (
		_w8199_,
		_w8208_,
		_w8209_
	);
	LUT2 #(
		.INIT('h1)
	) name7678 (
		_w8173_,
		_w8209_,
		_w8210_
	);
	LUT2 #(
		.INIT('h1)
	) name7679 (
		_w8064_,
		_w8073_,
		_w8211_
	);
	LUT2 #(
		.INIT('h4)
	) name7680 (
		_w8125_,
		_w8211_,
		_w8212_
	);
	LUT2 #(
		.INIT('h4)
	) name7681 (
		_w8210_,
		_w8212_,
		_w8213_
	);
	LUT2 #(
		.INIT('h4)
	) name7682 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w8214_
	);
	LUT2 #(
		.INIT('h1)
	) name7683 (
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w8215_
	);
	LUT2 #(
		.INIT('h4)
	) name7684 (
		\sa01_reg[5]/P0001 ,
		_w8215_,
		_w8216_
	);
	LUT2 #(
		.INIT('h8)
	) name7685 (
		_w8214_,
		_w8216_,
		_w8217_
	);
	LUT2 #(
		.INIT('h2)
	) name7686 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w8218_
	);
	LUT2 #(
		.INIT('h8)
	) name7687 (
		\sa01_reg[5]/P0001 ,
		_w8215_,
		_w8219_
	);
	LUT2 #(
		.INIT('h8)
	) name7688 (
		_w8218_,
		_w8219_,
		_w8220_
	);
	LUT2 #(
		.INIT('h4)
	) name7689 (
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w8221_
	);
	LUT2 #(
		.INIT('h2)
	) name7690 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w8222_
	);
	LUT2 #(
		.INIT('h8)
	) name7691 (
		_w8221_,
		_w8222_,
		_w8223_
	);
	LUT2 #(
		.INIT('h8)
	) name7692 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w8224_
	);
	LUT2 #(
		.INIT('h4)
	) name7693 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w8225_
	);
	LUT2 #(
		.INIT('h1)
	) name7694 (
		_w8224_,
		_w8225_,
		_w8226_
	);
	LUT2 #(
		.INIT('h1)
	) name7695 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w8227_
	);
	LUT2 #(
		.INIT('h2)
	) name7696 (
		\sa01_reg[7]/NET0131 ,
		_w8227_,
		_w8228_
	);
	LUT2 #(
		.INIT('h1)
	) name7697 (
		\sa01_reg[2]/P0001 ,
		_w8226_,
		_w8229_
	);
	LUT2 #(
		.INIT('h4)
	) name7698 (
		_w8228_,
		_w8229_,
		_w8230_
	);
	LUT2 #(
		.INIT('h2)
	) name7699 (
		\sa01_reg[1]/P0001 ,
		_w8223_,
		_w8231_
	);
	LUT2 #(
		.INIT('h4)
	) name7700 (
		_w8217_,
		_w8231_,
		_w8232_
	);
	LUT2 #(
		.INIT('h4)
	) name7701 (
		_w8220_,
		_w8232_,
		_w8233_
	);
	LUT2 #(
		.INIT('h4)
	) name7702 (
		_w8230_,
		_w8233_,
		_w8234_
	);
	LUT2 #(
		.INIT('h8)
	) name7703 (
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w8235_
	);
	LUT2 #(
		.INIT('h8)
	) name7704 (
		_w8218_,
		_w8235_,
		_w8236_
	);
	LUT2 #(
		.INIT('h1)
	) name7705 (
		\sa01_reg[1]/P0001 ,
		_w8236_,
		_w8237_
	);
	LUT2 #(
		.INIT('h8)
	) name7706 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w8238_
	);
	LUT2 #(
		.INIT('h4)
	) name7707 (
		\sa01_reg[6]/NET0131 ,
		_w8238_,
		_w8239_
	);
	LUT2 #(
		.INIT('h1)
	) name7708 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w8240_
	);
	LUT2 #(
		.INIT('h8)
	) name7709 (
		_w8239_,
		_w8240_,
		_w8241_
	);
	LUT2 #(
		.INIT('h2)
	) name7710 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w8242_
	);
	LUT2 #(
		.INIT('h8)
	) name7711 (
		_w8224_,
		_w8242_,
		_w8243_
	);
	LUT2 #(
		.INIT('h8)
	) name7712 (
		\sa01_reg[2]/P0001 ,
		_w8243_,
		_w8244_
	);
	LUT2 #(
		.INIT('h8)
	) name7713 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w8245_
	);
	LUT2 #(
		.INIT('h1)
	) name7714 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w8246_
	);
	LUT2 #(
		.INIT('h1)
	) name7715 (
		\sa01_reg[3]/P0001 ,
		_w8246_,
		_w8247_
	);
	LUT2 #(
		.INIT('h2)
	) name7716 (
		_w8245_,
		_w8247_,
		_w8248_
	);
	LUT2 #(
		.INIT('h2)
	) name7717 (
		_w8237_,
		_w8241_,
		_w8249_
	);
	LUT2 #(
		.INIT('h1)
	) name7718 (
		_w8244_,
		_w8248_,
		_w8250_
	);
	LUT2 #(
		.INIT('h8)
	) name7719 (
		_w8249_,
		_w8250_,
		_w8251_
	);
	LUT2 #(
		.INIT('h1)
	) name7720 (
		_w8234_,
		_w8251_,
		_w8252_
	);
	LUT2 #(
		.INIT('h2)
	) name7721 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w8253_
	);
	LUT2 #(
		.INIT('h4)
	) name7722 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w8254_
	);
	LUT2 #(
		.INIT('h8)
	) name7723 (
		_w8253_,
		_w8254_,
		_w8255_
	);
	LUT2 #(
		.INIT('h4)
	) name7724 (
		\sa01_reg[4]/P0001 ,
		_w8253_,
		_w8256_
	);
	LUT2 #(
		.INIT('h8)
	) name7725 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w8257_
	);
	LUT2 #(
		.INIT('h8)
	) name7726 (
		\sa01_reg[7]/NET0131 ,
		_w8257_,
		_w8258_
	);
	LUT2 #(
		.INIT('h1)
	) name7727 (
		_w8214_,
		_w8256_,
		_w8259_
	);
	LUT2 #(
		.INIT('h4)
	) name7728 (
		_w8258_,
		_w8259_,
		_w8260_
	);
	LUT2 #(
		.INIT('h1)
	) name7729 (
		_w8224_,
		_w8260_,
		_w8261_
	);
	LUT2 #(
		.INIT('h2)
	) name7730 (
		\sa01_reg[2]/P0001 ,
		_w8255_,
		_w8262_
	);
	LUT2 #(
		.INIT('h4)
	) name7731 (
		_w8261_,
		_w8262_,
		_w8263_
	);
	LUT2 #(
		.INIT('h8)
	) name7732 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w8264_
	);
	LUT2 #(
		.INIT('h1)
	) name7733 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w8265_
	);
	LUT2 #(
		.INIT('h8)
	) name7734 (
		_w8264_,
		_w8265_,
		_w8266_
	);
	LUT2 #(
		.INIT('h1)
	) name7735 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w8267_
	);
	LUT2 #(
		.INIT('h8)
	) name7736 (
		_w8216_,
		_w8267_,
		_w8268_
	);
	LUT2 #(
		.INIT('h8)
	) name7737 (
		_w8254_,
		_w8264_,
		_w8269_
	);
	LUT2 #(
		.INIT('h1)
	) name7738 (
		\sa01_reg[2]/P0001 ,
		_w8266_,
		_w8270_
	);
	LUT2 #(
		.INIT('h4)
	) name7739 (
		_w8269_,
		_w8270_,
		_w8271_
	);
	LUT2 #(
		.INIT('h4)
	) name7740 (
		_w8268_,
		_w8271_,
		_w8272_
	);
	LUT2 #(
		.INIT('h1)
	) name7741 (
		_w8263_,
		_w8272_,
		_w8273_
	);
	LUT2 #(
		.INIT('h1)
	) name7742 (
		_w8252_,
		_w8273_,
		_w8274_
	);
	LUT2 #(
		.INIT('h2)
	) name7743 (
		\sa01_reg[0]/P0001 ,
		_w8274_,
		_w8275_
	);
	LUT2 #(
		.INIT('h2)
	) name7744 (
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w8276_
	);
	LUT2 #(
		.INIT('h8)
	) name7745 (
		\sa01_reg[5]/P0001 ,
		_w8276_,
		_w8277_
	);
	LUT2 #(
		.INIT('h8)
	) name7746 (
		\sa01_reg[2]/P0001 ,
		_w8277_,
		_w8278_
	);
	LUT2 #(
		.INIT('h8)
	) name7747 (
		\sa01_reg[5]/P0001 ,
		_w8221_,
		_w8279_
	);
	LUT2 #(
		.INIT('h4)
	) name7748 (
		_w8218_,
		_w8279_,
		_w8280_
	);
	LUT2 #(
		.INIT('h4)
	) name7749 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w8281_
	);
	LUT2 #(
		.INIT('h4)
	) name7750 (
		\sa01_reg[5]/P0001 ,
		_w8281_,
		_w8282_
	);
	LUT2 #(
		.INIT('h4)
	) name7751 (
		\sa01_reg[6]/NET0131 ,
		_w8282_,
		_w8283_
	);
	LUT2 #(
		.INIT('h1)
	) name7752 (
		_w8280_,
		_w8283_,
		_w8284_
	);
	LUT2 #(
		.INIT('h1)
	) name7753 (
		\sa01_reg[2]/P0001 ,
		_w8284_,
		_w8285_
	);
	LUT2 #(
		.INIT('h8)
	) name7754 (
		_w8238_,
		_w8276_,
		_w8286_
	);
	LUT2 #(
		.INIT('h8)
	) name7755 (
		\sa01_reg[2]/P0001 ,
		_w8214_,
		_w8287_
	);
	LUT2 #(
		.INIT('h8)
	) name7756 (
		_w8254_,
		_w8287_,
		_w8288_
	);
	LUT2 #(
		.INIT('h2)
	) name7757 (
		\sa01_reg[1]/P0001 ,
		_w8286_,
		_w8289_
	);
	LUT2 #(
		.INIT('h4)
	) name7758 (
		_w8278_,
		_w8289_,
		_w8290_
	);
	LUT2 #(
		.INIT('h4)
	) name7759 (
		_w8288_,
		_w8290_,
		_w8291_
	);
	LUT2 #(
		.INIT('h4)
	) name7760 (
		_w8285_,
		_w8291_,
		_w8292_
	);
	LUT2 #(
		.INIT('h4)
	) name7761 (
		\sa01_reg[3]/P0001 ,
		_w8277_,
		_w8293_
	);
	LUT2 #(
		.INIT('h4)
	) name7762 (
		\sa01_reg[2]/P0001 ,
		_w8293_,
		_w8294_
	);
	LUT2 #(
		.INIT('h8)
	) name7763 (
		\sa01_reg[4]/P0001 ,
		_w8257_,
		_w8295_
	);
	LUT2 #(
		.INIT('h1)
	) name7764 (
		_w8216_,
		_w8295_,
		_w8296_
	);
	LUT2 #(
		.INIT('h2)
	) name7765 (
		\sa01_reg[2]/P0001 ,
		_w8296_,
		_w8297_
	);
	LUT2 #(
		.INIT('h8)
	) name7766 (
		_w8215_,
		_w8218_,
		_w8298_
	);
	LUT2 #(
		.INIT('h1)
	) name7767 (
		\sa01_reg[1]/P0001 ,
		_w8298_,
		_w8299_
	);
	LUT2 #(
		.INIT('h4)
	) name7768 (
		_w8294_,
		_w8299_,
		_w8300_
	);
	LUT2 #(
		.INIT('h4)
	) name7769 (
		_w8297_,
		_w8300_,
		_w8301_
	);
	LUT2 #(
		.INIT('h1)
	) name7770 (
		_w8292_,
		_w8301_,
		_w8302_
	);
	LUT2 #(
		.INIT('h2)
	) name7771 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[5]/P0001 ,
		_w8303_
	);
	LUT2 #(
		.INIT('h8)
	) name7772 (
		\sa01_reg[6]/NET0131 ,
		_w8267_,
		_w8304_
	);
	LUT2 #(
		.INIT('h8)
	) name7773 (
		_w8215_,
		_w8238_,
		_w8305_
	);
	LUT2 #(
		.INIT('h1)
	) name7774 (
		_w8304_,
		_w8305_,
		_w8306_
	);
	LUT2 #(
		.INIT('h2)
	) name7775 (
		_w8303_,
		_w8306_,
		_w8307_
	);
	LUT2 #(
		.INIT('h4)
	) name7776 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		_w8308_
	);
	LUT2 #(
		.INIT('h8)
	) name7777 (
		_w8215_,
		_w8308_,
		_w8309_
	);
	LUT2 #(
		.INIT('h4)
	) name7778 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w8310_
	);
	LUT2 #(
		.INIT('h4)
	) name7779 (
		\sa01_reg[2]/P0001 ,
		_w8224_,
		_w8311_
	);
	LUT2 #(
		.INIT('h8)
	) name7780 (
		_w8310_,
		_w8311_,
		_w8312_
	);
	LUT2 #(
		.INIT('h1)
	) name7781 (
		_w8309_,
		_w8312_,
		_w8313_
	);
	LUT2 #(
		.INIT('h1)
	) name7782 (
		\sa01_reg[3]/P0001 ,
		_w8313_,
		_w8314_
	);
	LUT2 #(
		.INIT('h1)
	) name7783 (
		_w8307_,
		_w8314_,
		_w8315_
	);
	LUT2 #(
		.INIT('h4)
	) name7784 (
		_w8302_,
		_w8315_,
		_w8316_
	);
	LUT2 #(
		.INIT('h1)
	) name7785 (
		\sa01_reg[0]/P0001 ,
		_w8316_,
		_w8317_
	);
	LUT2 #(
		.INIT('h2)
	) name7786 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		_w8318_
	);
	LUT2 #(
		.INIT('h4)
	) name7787 (
		_w8215_,
		_w8318_,
		_w8319_
	);
	LUT2 #(
		.INIT('h8)
	) name7788 (
		\sa01_reg[7]/NET0131 ,
		_w8267_,
		_w8320_
	);
	LUT2 #(
		.INIT('h8)
	) name7789 (
		\sa01_reg[5]/P0001 ,
		_w8320_,
		_w8321_
	);
	LUT2 #(
		.INIT('h8)
	) name7790 (
		\sa01_reg[6]/NET0131 ,
		_w8321_,
		_w8322_
	);
	LUT2 #(
		.INIT('h1)
	) name7791 (
		_w8268_,
		_w8319_,
		_w8323_
	);
	LUT2 #(
		.INIT('h4)
	) name7792 (
		_w8322_,
		_w8323_,
		_w8324_
	);
	LUT2 #(
		.INIT('h1)
	) name7793 (
		\sa01_reg[2]/P0001 ,
		_w8324_,
		_w8325_
	);
	LUT2 #(
		.INIT('h4)
	) name7794 (
		\sa01_reg[3]/P0001 ,
		_w8276_,
		_w8326_
	);
	LUT2 #(
		.INIT('h8)
	) name7795 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w8327_
	);
	LUT2 #(
		.INIT('h8)
	) name7796 (
		_w8326_,
		_w8327_,
		_w8328_
	);
	LUT2 #(
		.INIT('h8)
	) name7797 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		_w8329_
	);
	LUT2 #(
		.INIT('h8)
	) name7798 (
		_w8219_,
		_w8329_,
		_w8330_
	);
	LUT2 #(
		.INIT('h4)
	) name7799 (
		\sa01_reg[5]/P0001 ,
		_w8224_,
		_w8331_
	);
	LUT2 #(
		.INIT('h8)
	) name7800 (
		_w8264_,
		_w8331_,
		_w8332_
	);
	LUT2 #(
		.INIT('h8)
	) name7801 (
		_w8254_,
		_w8256_,
		_w8333_
	);
	LUT2 #(
		.INIT('h2)
	) name7802 (
		\sa01_reg[1]/P0001 ,
		_w8328_,
		_w8334_
	);
	LUT2 #(
		.INIT('h1)
	) name7803 (
		_w8330_,
		_w8332_,
		_w8335_
	);
	LUT2 #(
		.INIT('h4)
	) name7804 (
		_w8333_,
		_w8335_,
		_w8336_
	);
	LUT2 #(
		.INIT('h8)
	) name7805 (
		_w8334_,
		_w8336_,
		_w8337_
	);
	LUT2 #(
		.INIT('h4)
	) name7806 (
		_w8325_,
		_w8337_,
		_w8338_
	);
	LUT2 #(
		.INIT('h4)
	) name7807 (
		\sa01_reg[3]/P0001 ,
		_w8215_,
		_w8339_
	);
	LUT2 #(
		.INIT('h8)
	) name7808 (
		\sa01_reg[5]/P0001 ,
		_w8339_,
		_w8340_
	);
	LUT2 #(
		.INIT('h8)
	) name7809 (
		_w8253_,
		_w8308_,
		_w8341_
	);
	LUT2 #(
		.INIT('h2)
	) name7810 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w8342_
	);
	LUT2 #(
		.INIT('h8)
	) name7811 (
		_w8264_,
		_w8342_,
		_w8343_
	);
	LUT2 #(
		.INIT('h4)
	) name7812 (
		\sa01_reg[5]/P0001 ,
		_w8221_,
		_w8344_
	);
	LUT2 #(
		.INIT('h1)
	) name7813 (
		_w8214_,
		_w8218_,
		_w8345_
	);
	LUT2 #(
		.INIT('h8)
	) name7814 (
		_w8344_,
		_w8345_,
		_w8346_
	);
	LUT2 #(
		.INIT('h2)
	) name7815 (
		\sa01_reg[2]/P0001 ,
		_w8341_,
		_w8347_
	);
	LUT2 #(
		.INIT('h4)
	) name7816 (
		_w8343_,
		_w8347_,
		_w8348_
	);
	LUT2 #(
		.INIT('h1)
	) name7817 (
		_w8340_,
		_w8346_,
		_w8349_
	);
	LUT2 #(
		.INIT('h8)
	) name7818 (
		_w8348_,
		_w8349_,
		_w8350_
	);
	LUT2 #(
		.INIT('h1)
	) name7819 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		_w8351_
	);
	LUT2 #(
		.INIT('h8)
	) name7820 (
		_w8235_,
		_w8351_,
		_w8352_
	);
	LUT2 #(
		.INIT('h1)
	) name7821 (
		\sa01_reg[2]/P0001 ,
		_w8352_,
		_w8353_
	);
	LUT2 #(
		.INIT('h8)
	) name7822 (
		\sa01_reg[3]/P0001 ,
		_w8308_,
		_w8354_
	);
	LUT2 #(
		.INIT('h8)
	) name7823 (
		_w8235_,
		_w8354_,
		_w8355_
	);
	LUT2 #(
		.INIT('h8)
	) name7824 (
		_w8214_,
		_w8310_,
		_w8356_
	);
	LUT2 #(
		.INIT('h2)
	) name7825 (
		_w8353_,
		_w8356_,
		_w8357_
	);
	LUT2 #(
		.INIT('h4)
	) name7826 (
		_w8355_,
		_w8357_,
		_w8358_
	);
	LUT2 #(
		.INIT('h1)
	) name7827 (
		_w8350_,
		_w8358_,
		_w8359_
	);
	LUT2 #(
		.INIT('h8)
	) name7828 (
		_w8238_,
		_w8342_,
		_w8360_
	);
	LUT2 #(
		.INIT('h8)
	) name7829 (
		\sa01_reg[6]/NET0131 ,
		_w8360_,
		_w8361_
	);
	LUT2 #(
		.INIT('h8)
	) name7830 (
		_w8215_,
		_w8267_,
		_w8362_
	);
	LUT2 #(
		.INIT('h8)
	) name7831 (
		\sa01_reg[5]/P0001 ,
		_w8362_,
		_w8363_
	);
	LUT2 #(
		.INIT('h1)
	) name7832 (
		\sa01_reg[1]/P0001 ,
		_w8361_,
		_w8364_
	);
	LUT2 #(
		.INIT('h4)
	) name7833 (
		_w8363_,
		_w8364_,
		_w8365_
	);
	LUT2 #(
		.INIT('h4)
	) name7834 (
		_w8359_,
		_w8365_,
		_w8366_
	);
	LUT2 #(
		.INIT('h1)
	) name7835 (
		_w8338_,
		_w8366_,
		_w8367_
	);
	LUT2 #(
		.INIT('h1)
	) name7836 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w8368_
	);
	LUT2 #(
		.INIT('h8)
	) name7837 (
		_w8225_,
		_w8368_,
		_w8369_
	);
	LUT2 #(
		.INIT('h1)
	) name7838 (
		\sa01_reg[2]/P0001 ,
		_w8369_,
		_w8370_
	);
	LUT2 #(
		.INIT('h2)
	) name7839 (
		\sa01_reg[2]/P0001 ,
		_w8295_,
		_w8371_
	);
	LUT2 #(
		.INIT('h2)
	) name7840 (
		\sa01_reg[3]/P0001 ,
		_w8370_,
		_w8372_
	);
	LUT2 #(
		.INIT('h4)
	) name7841 (
		_w8371_,
		_w8372_,
		_w8373_
	);
	LUT2 #(
		.INIT('h1)
	) name7842 (
		_w8367_,
		_w8373_,
		_w8374_
	);
	LUT2 #(
		.INIT('h4)
	) name7843 (
		_w8275_,
		_w8374_,
		_w8375_
	);
	LUT2 #(
		.INIT('h4)
	) name7844 (
		_w8317_,
		_w8375_,
		_w8376_
	);
	LUT2 #(
		.INIT('h2)
	) name7845 (
		_w8213_,
		_w8376_,
		_w8377_
	);
	LUT2 #(
		.INIT('h4)
	) name7846 (
		_w8213_,
		_w8376_,
		_w8378_
	);
	LUT2 #(
		.INIT('h1)
	) name7847 (
		_w8377_,
		_w8378_,
		_w8379_
	);
	LUT2 #(
		.INIT('h8)
	) name7848 (
		_w8077_,
		_w8094_,
		_w8380_
	);
	LUT2 #(
		.INIT('h8)
	) name7849 (
		\sa12_reg[3]/P0001 ,
		_w8126_,
		_w8381_
	);
	LUT2 #(
		.INIT('h4)
	) name7850 (
		\sa12_reg[3]/P0001 ,
		_w8146_,
		_w8382_
	);
	LUT2 #(
		.INIT('h1)
	) name7851 (
		_w8380_,
		_w8381_,
		_w8383_
	);
	LUT2 #(
		.INIT('h4)
	) name7852 (
		_w8382_,
		_w8383_,
		_w8384_
	);
	LUT2 #(
		.INIT('h1)
	) name7853 (
		\sa12_reg[2]/P0001 ,
		_w8384_,
		_w8385_
	);
	LUT2 #(
		.INIT('h8)
	) name7854 (
		_w8161_,
		_w8180_,
		_w8386_
	);
	LUT2 #(
		.INIT('h8)
	) name7855 (
		_w8055_,
		_w8110_,
		_w8387_
	);
	LUT2 #(
		.INIT('h8)
	) name7856 (
		_w8077_,
		_w8111_,
		_w8388_
	);
	LUT2 #(
		.INIT('h8)
	) name7857 (
		\sa12_reg[3]/P0001 ,
		_w8161_,
		_w8389_
	);
	LUT2 #(
		.INIT('h8)
	) name7858 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w8390_
	);
	LUT2 #(
		.INIT('h8)
	) name7859 (
		_w8074_,
		_w8390_,
		_w8391_
	);
	LUT2 #(
		.INIT('h1)
	) name7860 (
		_w8389_,
		_w8391_,
		_w8392_
	);
	LUT2 #(
		.INIT('h2)
	) name7861 (
		\sa12_reg[2]/P0001 ,
		_w8392_,
		_w8393_
	);
	LUT2 #(
		.INIT('h8)
	) name7862 (
		_w8065_,
		_w8104_,
		_w8394_
	);
	LUT2 #(
		.INIT('h4)
	) name7863 (
		\sa12_reg[7]/NET0131 ,
		_w8394_,
		_w8395_
	);
	LUT2 #(
		.INIT('h1)
	) name7864 (
		_w8096_,
		_w8386_,
		_w8396_
	);
	LUT2 #(
		.INIT('h1)
	) name7865 (
		_w8387_,
		_w8388_,
		_w8397_
	);
	LUT2 #(
		.INIT('h8)
	) name7866 (
		_w8396_,
		_w8397_,
		_w8398_
	);
	LUT2 #(
		.INIT('h4)
	) name7867 (
		_w8395_,
		_w8398_,
		_w8399_
	);
	LUT2 #(
		.INIT('h4)
	) name7868 (
		_w8393_,
		_w8399_,
		_w8400_
	);
	LUT2 #(
		.INIT('h4)
	) name7869 (
		_w8385_,
		_w8400_,
		_w8401_
	);
	LUT2 #(
		.INIT('h2)
	) name7870 (
		\sa12_reg[1]/P0001 ,
		_w8401_,
		_w8402_
	);
	LUT2 #(
		.INIT('h8)
	) name7871 (
		\sa12_reg[2]/P0001 ,
		_w8129_,
		_w8403_
	);
	LUT2 #(
		.INIT('h4)
	) name7872 (
		\sa12_reg[6]/NET0131 ,
		_w8084_,
		_w8404_
	);
	LUT2 #(
		.INIT('h8)
	) name7873 (
		\sa12_reg[4]/P0001 ,
		_w8404_,
		_w8405_
	);
	LUT2 #(
		.INIT('h1)
	) name7874 (
		_w8403_,
		_w8405_,
		_w8406_
	);
	LUT2 #(
		.INIT('h1)
	) name7875 (
		\sa12_reg[5]/P0001 ,
		_w8406_,
		_w8407_
	);
	LUT2 #(
		.INIT('h4)
	) name7876 (
		\sa12_reg[3]/P0001 ,
		_w8194_,
		_w8408_
	);
	LUT2 #(
		.INIT('h1)
	) name7877 (
		_w8115_,
		_w8408_,
		_w8409_
	);
	LUT2 #(
		.INIT('h4)
	) name7878 (
		_w8407_,
		_w8409_,
		_w8410_
	);
	LUT2 #(
		.INIT('h1)
	) name7879 (
		\sa12_reg[1]/P0001 ,
		_w8410_,
		_w8411_
	);
	LUT2 #(
		.INIT('h4)
	) name7880 (
		\sa12_reg[5]/P0001 ,
		_w8060_,
		_w8412_
	);
	LUT2 #(
		.INIT('h4)
	) name7881 (
		\sa12_reg[3]/P0001 ,
		_w8412_,
		_w8413_
	);
	LUT2 #(
		.INIT('h4)
	) name7882 (
		\sa12_reg[4]/P0001 ,
		_w8069_,
		_w8414_
	);
	LUT2 #(
		.INIT('h1)
	) name7883 (
		_w8413_,
		_w8414_,
		_w8415_
	);
	LUT2 #(
		.INIT('h1)
	) name7884 (
		_w8104_,
		_w8415_,
		_w8416_
	);
	LUT2 #(
		.INIT('h4)
	) name7885 (
		\sa12_reg[4]/P0001 ,
		_w8055_,
		_w8417_
	);
	LUT2 #(
		.INIT('h1)
	) name7886 (
		_w8386_,
		_w8417_,
		_w8418_
	);
	LUT2 #(
		.INIT('h4)
	) name7887 (
		_w8416_,
		_w8418_,
		_w8419_
	);
	LUT2 #(
		.INIT('h2)
	) name7888 (
		\sa12_reg[2]/P0001 ,
		_w8419_,
		_w8420_
	);
	LUT2 #(
		.INIT('h4)
	) name7889 (
		\sa12_reg[2]/P0001 ,
		_w8166_,
		_w8421_
	);
	LUT2 #(
		.INIT('h8)
	) name7890 (
		_w8068_,
		_w8135_,
		_w8422_
	);
	LUT2 #(
		.INIT('h1)
	) name7891 (
		_w8200_,
		_w8422_,
		_w8423_
	);
	LUT2 #(
		.INIT('h1)
	) name7892 (
		\sa12_reg[2]/P0001 ,
		_w8423_,
		_w8424_
	);
	LUT2 #(
		.INIT('h4)
	) name7893 (
		\sa12_reg[4]/P0001 ,
		_w8142_,
		_w8425_
	);
	LUT2 #(
		.INIT('h1)
	) name7894 (
		_w8421_,
		_w8425_,
		_w8426_
	);
	LUT2 #(
		.INIT('h4)
	) name7895 (
		_w8424_,
		_w8426_,
		_w8427_
	);
	LUT2 #(
		.INIT('h4)
	) name7896 (
		_w8411_,
		_w8427_,
		_w8428_
	);
	LUT2 #(
		.INIT('h4)
	) name7897 (
		_w8420_,
		_w8428_,
		_w8429_
	);
	LUT2 #(
		.INIT('h4)
	) name7898 (
		_w8402_,
		_w8429_,
		_w8430_
	);
	LUT2 #(
		.INIT('h1)
	) name7899 (
		\sa12_reg[0]/P0001 ,
		_w8430_,
		_w8431_
	);
	LUT2 #(
		.INIT('h8)
	) name7900 (
		_w8065_,
		_w8080_,
		_w8432_
	);
	LUT2 #(
		.INIT('h4)
	) name7901 (
		\sa12_reg[3]/P0001 ,
		_w8432_,
		_w8433_
	);
	LUT2 #(
		.INIT('h8)
	) name7902 (
		_w8055_,
		_w8180_,
		_w8434_
	);
	LUT2 #(
		.INIT('h2)
	) name7903 (
		\sa12_reg[2]/P0001 ,
		_w8202_,
		_w8435_
	);
	LUT2 #(
		.INIT('h4)
	) name7904 (
		_w8434_,
		_w8435_,
		_w8436_
	);
	LUT2 #(
		.INIT('h1)
	) name7905 (
		\sa12_reg[2]/P0001 ,
		_w8127_,
		_w8437_
	);
	LUT2 #(
		.INIT('h4)
	) name7906 (
		_w8174_,
		_w8437_,
		_w8438_
	);
	LUT2 #(
		.INIT('h1)
	) name7907 (
		_w8436_,
		_w8438_,
		_w8439_
	);
	LUT2 #(
		.INIT('h1)
	) name7908 (
		_w8076_,
		_w8433_,
		_w8440_
	);
	LUT2 #(
		.INIT('h4)
	) name7909 (
		_w8439_,
		_w8440_,
		_w8441_
	);
	LUT2 #(
		.INIT('h1)
	) name7910 (
		\sa12_reg[1]/P0001 ,
		_w8441_,
		_w8442_
	);
	LUT2 #(
		.INIT('h4)
	) name7911 (
		\sa12_reg[4]/P0001 ,
		_w8074_,
		_w8443_
	);
	LUT2 #(
		.INIT('h1)
	) name7912 (
		_w8076_,
		_w8138_,
		_w8444_
	);
	LUT2 #(
		.INIT('h4)
	) name7913 (
		_w8443_,
		_w8444_,
		_w8445_
	);
	LUT2 #(
		.INIT('h1)
	) name7914 (
		\sa12_reg[2]/P0001 ,
		_w8445_,
		_w8446_
	);
	LUT2 #(
		.INIT('h8)
	) name7915 (
		\sa12_reg[2]/P0001 ,
		_w8104_,
		_w8447_
	);
	LUT2 #(
		.INIT('h8)
	) name7916 (
		_w8412_,
		_w8447_,
		_w8448_
	);
	LUT2 #(
		.INIT('h4)
	) name7917 (
		\sa12_reg[7]/NET0131 ,
		_w8097_,
		_w8449_
	);
	LUT2 #(
		.INIT('h8)
	) name7918 (
		\sa12_reg[2]/P0001 ,
		_w8094_,
		_w8450_
	);
	LUT2 #(
		.INIT('h8)
	) name7919 (
		_w8130_,
		_w8450_,
		_w8451_
	);
	LUT2 #(
		.INIT('h8)
	) name7920 (
		_w8080_,
		_w8093_,
		_w8452_
	);
	LUT2 #(
		.INIT('h4)
	) name7921 (
		\sa12_reg[2]/P0001 ,
		_w8452_,
		_w8453_
	);
	LUT2 #(
		.INIT('h2)
	) name7922 (
		\sa12_reg[5]/P0001 ,
		_w8078_,
		_w8454_
	);
	LUT2 #(
		.INIT('h2)
	) name7923 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[2]/P0001 ,
		_w8455_
	);
	LUT2 #(
		.INIT('h4)
	) name7924 (
		_w8080_,
		_w8455_,
		_w8456_
	);
	LUT2 #(
		.INIT('h4)
	) name7925 (
		_w8202_,
		_w8456_,
		_w8457_
	);
	LUT2 #(
		.INIT('h4)
	) name7926 (
		_w8454_,
		_w8457_,
		_w8458_
	);
	LUT2 #(
		.INIT('h4)
	) name7927 (
		\sa12_reg[6]/NET0131 ,
		_w8180_,
		_w8459_
	);
	LUT2 #(
		.INIT('h8)
	) name7928 (
		_w8074_,
		_w8459_,
		_w8460_
	);
	LUT2 #(
		.INIT('h8)
	) name7929 (
		\sa12_reg[7]/NET0131 ,
		_w8380_,
		_w8461_
	);
	LUT2 #(
		.INIT('h1)
	) name7930 (
		_w8460_,
		_w8461_,
		_w8462_
	);
	LUT2 #(
		.INIT('h8)
	) name7931 (
		_w8078_,
		_w8126_,
		_w8463_
	);
	LUT2 #(
		.INIT('h1)
	) name7932 (
		_w8143_,
		_w8463_,
		_w8464_
	);
	LUT2 #(
		.INIT('h8)
	) name7933 (
		_w8462_,
		_w8464_,
		_w8465_
	);
	LUT2 #(
		.INIT('h2)
	) name7934 (
		\sa12_reg[1]/P0001 ,
		_w8465_,
		_w8466_
	);
	LUT2 #(
		.INIT('h1)
	) name7935 (
		_w8448_,
		_w8449_,
		_w8467_
	);
	LUT2 #(
		.INIT('h1)
	) name7936 (
		_w8451_,
		_w8453_,
		_w8468_
	);
	LUT2 #(
		.INIT('h8)
	) name7937 (
		_w8467_,
		_w8468_,
		_w8469_
	);
	LUT2 #(
		.INIT('h4)
	) name7938 (
		_w8458_,
		_w8469_,
		_w8470_
	);
	LUT2 #(
		.INIT('h4)
	) name7939 (
		_w8446_,
		_w8470_,
		_w8471_
	);
	LUT2 #(
		.INIT('h4)
	) name7940 (
		_w8466_,
		_w8471_,
		_w8472_
	);
	LUT2 #(
		.INIT('h4)
	) name7941 (
		_w8442_,
		_w8472_,
		_w8473_
	);
	LUT2 #(
		.INIT('h2)
	) name7942 (
		\sa12_reg[0]/P0001 ,
		_w8473_,
		_w8474_
	);
	LUT2 #(
		.INIT('h1)
	) name7943 (
		_w8085_,
		_w8181_,
		_w8475_
	);
	LUT2 #(
		.INIT('h2)
	) name7944 (
		\sa12_reg[5]/P0001 ,
		_w8475_,
		_w8476_
	);
	LUT2 #(
		.INIT('h1)
	) name7945 (
		_w8452_,
		_w8476_,
		_w8477_
	);
	LUT2 #(
		.INIT('h1)
	) name7946 (
		\sa12_reg[2]/P0001 ,
		_w8477_,
		_w8478_
	);
	LUT2 #(
		.INIT('h8)
	) name7947 (
		\sa12_reg[2]/P0001 ,
		_w8180_,
		_w8479_
	);
	LUT2 #(
		.INIT('h8)
	) name7948 (
		_w8077_,
		_w8479_,
		_w8480_
	);
	LUT2 #(
		.INIT('h4)
	) name7949 (
		\sa12_reg[5]/P0001 ,
		_w8126_,
		_w8481_
	);
	LUT2 #(
		.INIT('h1)
	) name7950 (
		_w8412_,
		_w8481_,
		_w8482_
	);
	LUT2 #(
		.INIT('h4)
	) name7951 (
		_w8130_,
		_w8482_,
		_w8483_
	);
	LUT2 #(
		.INIT('h2)
	) name7952 (
		_w8450_,
		_w8483_,
		_w8484_
	);
	LUT2 #(
		.INIT('h8)
	) name7953 (
		_w8055_,
		_w8104_,
		_w8485_
	);
	LUT2 #(
		.INIT('h1)
	) name7954 (
		_w8480_,
		_w8485_,
		_w8486_
	);
	LUT2 #(
		.INIT('h4)
	) name7955 (
		_w8484_,
		_w8486_,
		_w8487_
	);
	LUT2 #(
		.INIT('h4)
	) name7956 (
		_w8478_,
		_w8487_,
		_w8488_
	);
	LUT2 #(
		.INIT('h1)
	) name7957 (
		\sa12_reg[1]/P0001 ,
		_w8488_,
		_w8489_
	);
	LUT2 #(
		.INIT('h8)
	) name7958 (
		\sa12_reg[5]/P0001 ,
		_w8156_,
		_w8490_
	);
	LUT2 #(
		.INIT('h8)
	) name7959 (
		_w8057_,
		_w8490_,
		_w8491_
	);
	LUT2 #(
		.INIT('h1)
	) name7960 (
		_w8096_,
		_w8150_,
		_w8492_
	);
	LUT2 #(
		.INIT('h1)
	) name7961 (
		\sa12_reg[2]/P0001 ,
		_w8492_,
		_w8493_
	);
	LUT2 #(
		.INIT('h8)
	) name7962 (
		_w8074_,
		_w8094_,
		_w8494_
	);
	LUT2 #(
		.INIT('h8)
	) name7963 (
		\sa12_reg[6]/NET0131 ,
		_w8494_,
		_w8495_
	);
	LUT2 #(
		.INIT('h8)
	) name7964 (
		\sa12_reg[2]/P0001 ,
		_w8495_,
		_w8496_
	);
	LUT2 #(
		.INIT('h4)
	) name7965 (
		\sa12_reg[6]/NET0131 ,
		_w8110_,
		_w8497_
	);
	LUT2 #(
		.INIT('h1)
	) name7966 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w8498_
	);
	LUT2 #(
		.INIT('h8)
	) name7967 (
		_w8497_,
		_w8498_,
		_w8499_
	);
	LUT2 #(
		.INIT('h1)
	) name7968 (
		_w8421_,
		_w8499_,
		_w8500_
	);
	LUT2 #(
		.INIT('h4)
	) name7969 (
		_w8496_,
		_w8500_,
		_w8501_
	);
	LUT2 #(
		.INIT('h2)
	) name7970 (
		\sa12_reg[1]/P0001 ,
		_w8501_,
		_w8502_
	);
	LUT2 #(
		.INIT('h1)
	) name7971 (
		_w8491_,
		_w8493_,
		_w8503_
	);
	LUT2 #(
		.INIT('h4)
	) name7972 (
		_w8502_,
		_w8503_,
		_w8504_
	);
	LUT2 #(
		.INIT('h4)
	) name7973 (
		_w8489_,
		_w8504_,
		_w8505_
	);
	LUT2 #(
		.INIT('h4)
	) name7974 (
		_w8474_,
		_w8505_,
		_w8506_
	);
	LUT2 #(
		.INIT('h4)
	) name7975 (
		_w8431_,
		_w8506_,
		_w8507_
	);
	LUT2 #(
		.INIT('h2)
	) name7976 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w8508_
	);
	LUT2 #(
		.INIT('h4)
	) name7977 (
		\sa23_reg[3]/P0001 ,
		_w8508_,
		_w8509_
	);
	LUT2 #(
		.INIT('h8)
	) name7978 (
		\sa23_reg[4]/P0001 ,
		_w8509_,
		_w8510_
	);
	LUT2 #(
		.INIT('h4)
	) name7979 (
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w8511_
	);
	LUT2 #(
		.INIT('h8)
	) name7980 (
		\sa23_reg[3]/P0001 ,
		_w8511_,
		_w8512_
	);
	LUT2 #(
		.INIT('h2)
	) name7981 (
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w8513_
	);
	LUT2 #(
		.INIT('h4)
	) name7982 (
		\sa23_reg[4]/P0001 ,
		_w8513_,
		_w8514_
	);
	LUT2 #(
		.INIT('h4)
	) name7983 (
		\sa23_reg[3]/P0001 ,
		_w8514_,
		_w8515_
	);
	LUT2 #(
		.INIT('h1)
	) name7984 (
		_w8510_,
		_w8512_,
		_w8516_
	);
	LUT2 #(
		.INIT('h4)
	) name7985 (
		_w8515_,
		_w8516_,
		_w8517_
	);
	LUT2 #(
		.INIT('h1)
	) name7986 (
		\sa23_reg[2]/P0001 ,
		_w8517_,
		_w8518_
	);
	LUT2 #(
		.INIT('h4)
	) name7987 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w8519_
	);
	LUT2 #(
		.INIT('h8)
	) name7988 (
		_w8508_,
		_w8519_,
		_w8520_
	);
	LUT2 #(
		.INIT('h8)
	) name7989 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w8521_
	);
	LUT2 #(
		.INIT('h1)
	) name7990 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w8522_
	);
	LUT2 #(
		.INIT('h4)
	) name7991 (
		\sa23_reg[7]/NET0131 ,
		_w8522_,
		_w8523_
	);
	LUT2 #(
		.INIT('h8)
	) name7992 (
		_w8521_,
		_w8523_,
		_w8524_
	);
	LUT2 #(
		.INIT('h4)
	) name7993 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w8525_
	);
	LUT2 #(
		.INIT('h4)
	) name7994 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w8526_
	);
	LUT2 #(
		.INIT('h8)
	) name7995 (
		_w8525_,
		_w8526_,
		_w8527_
	);
	LUT2 #(
		.INIT('h1)
	) name7996 (
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w8528_
	);
	LUT2 #(
		.INIT('h2)
	) name7997 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		_w8529_
	);
	LUT2 #(
		.INIT('h8)
	) name7998 (
		_w8528_,
		_w8529_,
		_w8530_
	);
	LUT2 #(
		.INIT('h8)
	) name7999 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w8531_
	);
	LUT2 #(
		.INIT('h8)
	) name8000 (
		\sa23_reg[3]/P0001 ,
		_w8531_,
		_w8532_
	);
	LUT2 #(
		.INIT('h8)
	) name8001 (
		\sa23_reg[4]/P0001 ,
		_w8521_,
		_w8533_
	);
	LUT2 #(
		.INIT('h4)
	) name8002 (
		\sa23_reg[7]/NET0131 ,
		_w8533_,
		_w8534_
	);
	LUT2 #(
		.INIT('h1)
	) name8003 (
		_w8532_,
		_w8534_,
		_w8535_
	);
	LUT2 #(
		.INIT('h2)
	) name8004 (
		\sa23_reg[2]/P0001 ,
		_w8535_,
		_w8536_
	);
	LUT2 #(
		.INIT('h8)
	) name8005 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w8537_
	);
	LUT2 #(
		.INIT('h8)
	) name8006 (
		_w8531_,
		_w8537_,
		_w8538_
	);
	LUT2 #(
		.INIT('h1)
	) name8007 (
		_w8520_,
		_w8527_,
		_w8539_
	);
	LUT2 #(
		.INIT('h1)
	) name8008 (
		_w8530_,
		_w8538_,
		_w8540_
	);
	LUT2 #(
		.INIT('h8)
	) name8009 (
		_w8539_,
		_w8540_,
		_w8541_
	);
	LUT2 #(
		.INIT('h4)
	) name8010 (
		_w8524_,
		_w8541_,
		_w8542_
	);
	LUT2 #(
		.INIT('h4)
	) name8011 (
		_w8536_,
		_w8542_,
		_w8543_
	);
	LUT2 #(
		.INIT('h4)
	) name8012 (
		_w8518_,
		_w8543_,
		_w8544_
	);
	LUT2 #(
		.INIT('h2)
	) name8013 (
		\sa23_reg[1]/P0001 ,
		_w8544_,
		_w8545_
	);
	LUT2 #(
		.INIT('h8)
	) name8014 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		_w8546_
	);
	LUT2 #(
		.INIT('h1)
	) name8015 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w8547_
	);
	LUT2 #(
		.INIT('h4)
	) name8016 (
		\sa23_reg[4]/P0001 ,
		_w8547_,
		_w8548_
	);
	LUT2 #(
		.INIT('h8)
	) name8017 (
		_w8546_,
		_w8548_,
		_w8549_
	);
	LUT2 #(
		.INIT('h4)
	) name8018 (
		\sa23_reg[6]/NET0131 ,
		_w8526_,
		_w8550_
	);
	LUT2 #(
		.INIT('h8)
	) name8019 (
		\sa23_reg[4]/P0001 ,
		_w8550_,
		_w8551_
	);
	LUT2 #(
		.INIT('h4)
	) name8020 (
		\sa23_reg[3]/P0001 ,
		_w8528_,
		_w8552_
	);
	LUT2 #(
		.INIT('h8)
	) name8021 (
		\sa23_reg[2]/P0001 ,
		_w8552_,
		_w8553_
	);
	LUT2 #(
		.INIT('h1)
	) name8022 (
		_w8551_,
		_w8553_,
		_w8554_
	);
	LUT2 #(
		.INIT('h1)
	) name8023 (
		\sa23_reg[5]/P0001 ,
		_w8554_,
		_w8555_
	);
	LUT2 #(
		.INIT('h4)
	) name8024 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w8556_
	);
	LUT2 #(
		.INIT('h8)
	) name8025 (
		_w8531_,
		_w8556_,
		_w8557_
	);
	LUT2 #(
		.INIT('h4)
	) name8026 (
		\sa23_reg[3]/P0001 ,
		_w8557_,
		_w8558_
	);
	LUT2 #(
		.INIT('h1)
	) name8027 (
		_w8549_,
		_w8558_,
		_w8559_
	);
	LUT2 #(
		.INIT('h4)
	) name8028 (
		_w8555_,
		_w8559_,
		_w8560_
	);
	LUT2 #(
		.INIT('h1)
	) name8029 (
		\sa23_reg[1]/P0001 ,
		_w8560_,
		_w8561_
	);
	LUT2 #(
		.INIT('h4)
	) name8030 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w8562_
	);
	LUT2 #(
		.INIT('h8)
	) name8031 (
		_w8556_,
		_w8562_,
		_w8563_
	);
	LUT2 #(
		.INIT('h1)
	) name8032 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w8564_
	);
	LUT2 #(
		.INIT('h8)
	) name8033 (
		_w8537_,
		_w8564_,
		_w8565_
	);
	LUT2 #(
		.INIT('h1)
	) name8034 (
		_w8563_,
		_w8565_,
		_w8566_
	);
	LUT2 #(
		.INIT('h1)
	) name8035 (
		\sa23_reg[2]/P0001 ,
		_w8566_,
		_w8567_
	);
	LUT2 #(
		.INIT('h4)
	) name8036 (
		\sa23_reg[7]/NET0131 ,
		_w8548_,
		_w8568_
	);
	LUT2 #(
		.INIT('h8)
	) name8037 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w8569_
	);
	LUT2 #(
		.INIT('h8)
	) name8038 (
		_w8508_,
		_w8569_,
		_w8570_
	);
	LUT2 #(
		.INIT('h4)
	) name8039 (
		\sa23_reg[2]/P0001 ,
		_w8570_,
		_w8571_
	);
	LUT2 #(
		.INIT('h2)
	) name8040 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w8572_
	);
	LUT2 #(
		.INIT('h4)
	) name8041 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w8573_
	);
	LUT2 #(
		.INIT('h8)
	) name8042 (
		\sa23_reg[6]/NET0131 ,
		_w8573_,
		_w8574_
	);
	LUT2 #(
		.INIT('h1)
	) name8043 (
		_w8572_,
		_w8574_,
		_w8575_
	);
	LUT2 #(
		.INIT('h2)
	) name8044 (
		_w8564_,
		_w8575_,
		_w8576_
	);
	LUT2 #(
		.INIT('h1)
	) name8045 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w8577_
	);
	LUT2 #(
		.INIT('h4)
	) name8046 (
		\sa23_reg[6]/NET0131 ,
		_w8577_,
		_w8578_
	);
	LUT2 #(
		.INIT('h1)
	) name8047 (
		_w8538_,
		_w8578_,
		_w8579_
	);
	LUT2 #(
		.INIT('h4)
	) name8048 (
		_w8576_,
		_w8579_,
		_w8580_
	);
	LUT2 #(
		.INIT('h2)
	) name8049 (
		\sa23_reg[2]/P0001 ,
		_w8580_,
		_w8581_
	);
	LUT2 #(
		.INIT('h1)
	) name8050 (
		_w8568_,
		_w8571_,
		_w8582_
	);
	LUT2 #(
		.INIT('h4)
	) name8051 (
		_w8567_,
		_w8582_,
		_w8583_
	);
	LUT2 #(
		.INIT('h4)
	) name8052 (
		_w8581_,
		_w8583_,
		_w8584_
	);
	LUT2 #(
		.INIT('h4)
	) name8053 (
		_w8561_,
		_w8584_,
		_w8585_
	);
	LUT2 #(
		.INIT('h4)
	) name8054 (
		_w8545_,
		_w8585_,
		_w8586_
	);
	LUT2 #(
		.INIT('h1)
	) name8055 (
		\sa23_reg[0]/P0001 ,
		_w8586_,
		_w8587_
	);
	LUT2 #(
		.INIT('h8)
	) name8056 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w8588_
	);
	LUT2 #(
		.INIT('h2)
	) name8057 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w8589_
	);
	LUT2 #(
		.INIT('h8)
	) name8058 (
		_w8588_,
		_w8589_,
		_w8590_
	);
	LUT2 #(
		.INIT('h8)
	) name8059 (
		_w8513_,
		_w8572_,
		_w8591_
	);
	LUT2 #(
		.INIT('h1)
	) name8060 (
		_w8590_,
		_w8591_,
		_w8592_
	);
	LUT2 #(
		.INIT('h8)
	) name8061 (
		\sa23_reg[5]/P0001 ,
		_w8572_,
		_w8593_
	);
	LUT2 #(
		.INIT('h1)
	) name8062 (
		\sa23_reg[5]/P0001 ,
		_w8556_,
		_w8594_
	);
	LUT2 #(
		.INIT('h4)
	) name8063 (
		_w8569_,
		_w8594_,
		_w8595_
	);
	LUT2 #(
		.INIT('h1)
	) name8064 (
		_w8593_,
		_w8595_,
		_w8596_
	);
	LUT2 #(
		.INIT('h2)
	) name8065 (
		\sa23_reg[1]/P0001 ,
		_w8596_,
		_w8597_
	);
	LUT2 #(
		.INIT('h4)
	) name8066 (
		\sa23_reg[4]/P0001 ,
		_w8589_,
		_w8598_
	);
	LUT2 #(
		.INIT('h2)
	) name8067 (
		_w8592_,
		_w8598_,
		_w8599_
	);
	LUT2 #(
		.INIT('h4)
	) name8068 (
		_w8597_,
		_w8599_,
		_w8600_
	);
	LUT2 #(
		.INIT('h2)
	) name8069 (
		\sa23_reg[0]/P0001 ,
		_w8600_,
		_w8601_
	);
	LUT2 #(
		.INIT('h8)
	) name8070 (
		_w8525_,
		_w8569_,
		_w8602_
	);
	LUT2 #(
		.INIT('h4)
	) name8071 (
		\sa23_reg[3]/P0001 ,
		_w8519_,
		_w8603_
	);
	LUT2 #(
		.INIT('h8)
	) name8072 (
		_w8513_,
		_w8537_,
		_w8604_
	);
	LUT2 #(
		.INIT('h1)
	) name8073 (
		_w8603_,
		_w8604_,
		_w8605_
	);
	LUT2 #(
		.INIT('h2)
	) name8074 (
		\sa23_reg[5]/P0001 ,
		_w8605_,
		_w8606_
	);
	LUT2 #(
		.INIT('h1)
	) name8075 (
		_w8602_,
		_w8606_,
		_w8607_
	);
	LUT2 #(
		.INIT('h1)
	) name8076 (
		\sa23_reg[1]/P0001 ,
		_w8607_,
		_w8608_
	);
	LUT2 #(
		.INIT('h8)
	) name8077 (
		_w8528_,
		_w8593_,
		_w8609_
	);
	LUT2 #(
		.INIT('h1)
	) name8078 (
		_w8527_,
		_w8609_,
		_w8610_
	);
	LUT2 #(
		.INIT('h4)
	) name8079 (
		_w8608_,
		_w8610_,
		_w8611_
	);
	LUT2 #(
		.INIT('h4)
	) name8080 (
		_w8601_,
		_w8611_,
		_w8612_
	);
	LUT2 #(
		.INIT('h1)
	) name8081 (
		\sa23_reg[2]/P0001 ,
		_w8612_,
		_w8613_
	);
	LUT2 #(
		.INIT('h8)
	) name8082 (
		\sa23_reg[5]/P0001 ,
		_w8513_,
		_w8614_
	);
	LUT2 #(
		.INIT('h8)
	) name8083 (
		_w8511_,
		_w8529_,
		_w8615_
	);
	LUT2 #(
		.INIT('h1)
	) name8084 (
		_w8614_,
		_w8615_,
		_w8616_
	);
	LUT2 #(
		.INIT('h1)
	) name8085 (
		\sa23_reg[2]/P0001 ,
		_w8616_,
		_w8617_
	);
	LUT2 #(
		.INIT('h8)
	) name8086 (
		\sa23_reg[3]/P0001 ,
		_w8589_,
		_w8618_
	);
	LUT2 #(
		.INIT('h8)
	) name8087 (
		_w8531_,
		_w8573_,
		_w8619_
	);
	LUT2 #(
		.INIT('h1)
	) name8088 (
		_w8618_,
		_w8619_,
		_w8620_
	);
	LUT2 #(
		.INIT('h2)
	) name8089 (
		\sa23_reg[6]/NET0131 ,
		_w8620_,
		_w8621_
	);
	LUT2 #(
		.INIT('h4)
	) name8090 (
		\sa23_reg[4]/P0001 ,
		_w8525_,
		_w8622_
	);
	LUT2 #(
		.INIT('h2)
	) name8091 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w8623_
	);
	LUT2 #(
		.INIT('h2)
	) name8092 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w8624_
	);
	LUT2 #(
		.INIT('h8)
	) name8093 (
		_w8623_,
		_w8624_,
		_w8625_
	);
	LUT2 #(
		.INIT('h1)
	) name8094 (
		_w8622_,
		_w8625_,
		_w8626_
	);
	LUT2 #(
		.INIT('h2)
	) name8095 (
		\sa23_reg[2]/P0001 ,
		_w8626_,
		_w8627_
	);
	LUT2 #(
		.INIT('h1)
	) name8096 (
		_w8617_,
		_w8621_,
		_w8628_
	);
	LUT2 #(
		.INIT('h4)
	) name8097 (
		_w8627_,
		_w8628_,
		_w8629_
	);
	LUT2 #(
		.INIT('h1)
	) name8098 (
		\sa23_reg[1]/P0001 ,
		_w8629_,
		_w8630_
	);
	LUT2 #(
		.INIT('h8)
	) name8099 (
		\sa23_reg[5]/P0001 ,
		_w8528_,
		_w8631_
	);
	LUT2 #(
		.INIT('h8)
	) name8100 (
		_w8537_,
		_w8631_,
		_w8632_
	);
	LUT2 #(
		.INIT('h8)
	) name8101 (
		_w8509_,
		_w8569_,
		_w8633_
	);
	LUT2 #(
		.INIT('h1)
	) name8102 (
		_w8632_,
		_w8633_,
		_w8634_
	);
	LUT2 #(
		.INIT('h4)
	) name8103 (
		\sa23_reg[7]/NET0131 ,
		_w8573_,
		_w8635_
	);
	LUT2 #(
		.INIT('h8)
	) name8104 (
		_w8547_,
		_w8635_,
		_w8636_
	);
	LUT2 #(
		.INIT('h4)
	) name8105 (
		\sa23_reg[4]/P0001 ,
		_w8512_,
		_w8637_
	);
	LUT2 #(
		.INIT('h1)
	) name8106 (
		_w8636_,
		_w8637_,
		_w8638_
	);
	LUT2 #(
		.INIT('h8)
	) name8107 (
		_w8634_,
		_w8638_,
		_w8639_
	);
	LUT2 #(
		.INIT('h2)
	) name8108 (
		\sa23_reg[1]/P0001 ,
		_w8639_,
		_w8640_
	);
	LUT2 #(
		.INIT('h8)
	) name8109 (
		_w8531_,
		_w8574_,
		_w8641_
	);
	LUT2 #(
		.INIT('h4)
	) name8110 (
		\sa23_reg[3]/P0001 ,
		_w8525_,
		_w8642_
	);
	LUT2 #(
		.INIT('h8)
	) name8111 (
		_w8577_,
		_w8642_,
		_w8643_
	);
	LUT2 #(
		.INIT('h1)
	) name8112 (
		_w8641_,
		_w8643_,
		_w8644_
	);
	LUT2 #(
		.INIT('h2)
	) name8113 (
		\sa23_reg[2]/P0001 ,
		_w8644_,
		_w8645_
	);
	LUT2 #(
		.INIT('h4)
	) name8114 (
		\sa23_reg[2]/P0001 ,
		_w8602_,
		_w8646_
	);
	LUT2 #(
		.INIT('h8)
	) name8115 (
		_w8572_,
		_w8614_,
		_w8647_
	);
	LUT2 #(
		.INIT('h1)
	) name8116 (
		_w8646_,
		_w8647_,
		_w8648_
	);
	LUT2 #(
		.INIT('h4)
	) name8117 (
		_w8645_,
		_w8648_,
		_w8649_
	);
	LUT2 #(
		.INIT('h4)
	) name8118 (
		_w8640_,
		_w8649_,
		_w8650_
	);
	LUT2 #(
		.INIT('h4)
	) name8119 (
		_w8630_,
		_w8650_,
		_w8651_
	);
	LUT2 #(
		.INIT('h2)
	) name8120 (
		\sa23_reg[0]/P0001 ,
		_w8651_,
		_w8652_
	);
	LUT2 #(
		.INIT('h8)
	) name8121 (
		\sa23_reg[6]/NET0131 ,
		_w8531_,
		_w8653_
	);
	LUT2 #(
		.INIT('h4)
	) name8122 (
		\sa23_reg[5]/P0001 ,
		_w8511_,
		_w8654_
	);
	LUT2 #(
		.INIT('h4)
	) name8123 (
		\sa23_reg[5]/P0001 ,
		_w8513_,
		_w8655_
	);
	LUT2 #(
		.INIT('h1)
	) name8124 (
		_w8654_,
		_w8655_,
		_w8656_
	);
	LUT2 #(
		.INIT('h4)
	) name8125 (
		_w8653_,
		_w8656_,
		_w8657_
	);
	LUT2 #(
		.INIT('h8)
	) name8126 (
		\sa23_reg[2]/P0001 ,
		_w8573_,
		_w8658_
	);
	LUT2 #(
		.INIT('h4)
	) name8127 (
		_w8657_,
		_w8658_,
		_w8659_
	);
	LUT2 #(
		.INIT('h2)
	) name8128 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w8660_
	);
	LUT2 #(
		.INIT('h8)
	) name8129 (
		\sa23_reg[5]/P0001 ,
		_w8537_,
		_w8661_
	);
	LUT2 #(
		.INIT('h8)
	) name8130 (
		_w8660_,
		_w8661_,
		_w8662_
	);
	LUT2 #(
		.INIT('h8)
	) name8131 (
		_w8522_,
		_w8528_,
		_w8663_
	);
	LUT2 #(
		.INIT('h1)
	) name8132 (
		_w8662_,
		_w8663_,
		_w8664_
	);
	LUT2 #(
		.INIT('h4)
	) name8133 (
		_w8659_,
		_w8664_,
		_w8665_
	);
	LUT2 #(
		.INIT('h1)
	) name8134 (
		\sa23_reg[1]/P0001 ,
		_w8665_,
		_w8666_
	);
	LUT2 #(
		.INIT('h8)
	) name8135 (
		_w8508_,
		_w8623_,
		_w8667_
	);
	LUT2 #(
		.INIT('h8)
	) name8136 (
		_w8546_,
		_w8667_,
		_w8668_
	);
	LUT2 #(
		.INIT('h8)
	) name8137 (
		_w8614_,
		_w8658_,
		_w8669_
	);
	LUT2 #(
		.INIT('h8)
	) name8138 (
		_w8529_,
		_w8578_,
		_w8670_
	);
	LUT2 #(
		.INIT('h1)
	) name8139 (
		_w8571_,
		_w8669_,
		_w8671_
	);
	LUT2 #(
		.INIT('h4)
	) name8140 (
		_w8670_,
		_w8671_,
		_w8672_
	);
	LUT2 #(
		.INIT('h2)
	) name8141 (
		\sa23_reg[1]/P0001 ,
		_w8672_,
		_w8673_
	);
	LUT2 #(
		.INIT('h1)
	) name8142 (
		_w8668_,
		_w8673_,
		_w8674_
	);
	LUT2 #(
		.INIT('h4)
	) name8143 (
		_w8666_,
		_w8674_,
		_w8675_
	);
	LUT2 #(
		.INIT('h4)
	) name8144 (
		_w8613_,
		_w8675_,
		_w8676_
	);
	LUT2 #(
		.INIT('h4)
	) name8145 (
		_w8652_,
		_w8676_,
		_w8677_
	);
	LUT2 #(
		.INIT('h4)
	) name8146 (
		_w8587_,
		_w8677_,
		_w8678_
	);
	LUT2 #(
		.INIT('h2)
	) name8147 (
		_w8507_,
		_w8678_,
		_w8679_
	);
	LUT2 #(
		.INIT('h4)
	) name8148 (
		_w8507_,
		_w8678_,
		_w8680_
	);
	LUT2 #(
		.INIT('h1)
	) name8149 (
		_w8679_,
		_w8680_,
		_w8681_
	);
	LUT2 #(
		.INIT('h4)
	) name8150 (
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w8682_
	);
	LUT2 #(
		.INIT('h8)
	) name8151 (
		\sa30_reg[3]/P0001 ,
		_w8682_,
		_w8683_
	);
	LUT2 #(
		.INIT('h2)
	) name8152 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w8684_
	);
	LUT2 #(
		.INIT('h8)
	) name8153 (
		\sa30_reg[4]/P0001 ,
		_w8684_,
		_w8685_
	);
	LUT2 #(
		.INIT('h2)
	) name8154 (
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w8686_
	);
	LUT2 #(
		.INIT('h4)
	) name8155 (
		\sa30_reg[4]/P0001 ,
		_w8686_,
		_w8687_
	);
	LUT2 #(
		.INIT('h1)
	) name8156 (
		_w8685_,
		_w8687_,
		_w8688_
	);
	LUT2 #(
		.INIT('h1)
	) name8157 (
		\sa30_reg[3]/P0001 ,
		_w8688_,
		_w8689_
	);
	LUT2 #(
		.INIT('h1)
	) name8158 (
		_w8683_,
		_w8689_,
		_w8690_
	);
	LUT2 #(
		.INIT('h1)
	) name8159 (
		\sa30_reg[2]/P0001 ,
		_w8690_,
		_w8691_
	);
	LUT2 #(
		.INIT('h8)
	) name8160 (
		\sa30_reg[7]/P0001 ,
		_w8684_,
		_w8692_
	);
	LUT2 #(
		.INIT('h4)
	) name8161 (
		\sa30_reg[4]/P0001 ,
		_w8692_,
		_w8693_
	);
	LUT2 #(
		.INIT('h8)
	) name8162 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w8694_
	);
	LUT2 #(
		.INIT('h8)
	) name8163 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w8695_
	);
	LUT2 #(
		.INIT('h8)
	) name8164 (
		_w8694_,
		_w8695_,
		_w8696_
	);
	LUT2 #(
		.INIT('h8)
	) name8165 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w8697_
	);
	LUT2 #(
		.INIT('h1)
	) name8166 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w8698_
	);
	LUT2 #(
		.INIT('h8)
	) name8167 (
		_w8697_,
		_w8698_,
		_w8699_
	);
	LUT2 #(
		.INIT('h4)
	) name8168 (
		\sa30_reg[7]/P0001 ,
		_w8699_,
		_w8700_
	);
	LUT2 #(
		.INIT('h1)
	) name8169 (
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w8701_
	);
	LUT2 #(
		.INIT('h2)
	) name8170 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		_w8702_
	);
	LUT2 #(
		.INIT('h8)
	) name8171 (
		_w8701_,
		_w8702_,
		_w8703_
	);
	LUT2 #(
		.INIT('h8)
	) name8172 (
		\sa30_reg[3]/P0001 ,
		_w8694_,
		_w8704_
	);
	LUT2 #(
		.INIT('h4)
	) name8173 (
		\sa30_reg[7]/P0001 ,
		_w8697_,
		_w8705_
	);
	LUT2 #(
		.INIT('h8)
	) name8174 (
		\sa30_reg[4]/P0001 ,
		_w8705_,
		_w8706_
	);
	LUT2 #(
		.INIT('h1)
	) name8175 (
		_w8704_,
		_w8706_,
		_w8707_
	);
	LUT2 #(
		.INIT('h2)
	) name8176 (
		\sa30_reg[2]/P0001 ,
		_w8707_,
		_w8708_
	);
	LUT2 #(
		.INIT('h8)
	) name8177 (
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w8709_
	);
	LUT2 #(
		.INIT('h4)
	) name8178 (
		\sa30_reg[5]/P0001 ,
		_w8709_,
		_w8710_
	);
	LUT2 #(
		.INIT('h4)
	) name8179 (
		\sa30_reg[3]/P0001 ,
		_w8710_,
		_w8711_
	);
	LUT2 #(
		.INIT('h1)
	) name8180 (
		_w8696_,
		_w8703_,
		_w8712_
	);
	LUT2 #(
		.INIT('h4)
	) name8181 (
		_w8693_,
		_w8712_,
		_w8713_
	);
	LUT2 #(
		.INIT('h1)
	) name8182 (
		_w8700_,
		_w8711_,
		_w8714_
	);
	LUT2 #(
		.INIT('h8)
	) name8183 (
		_w8713_,
		_w8714_,
		_w8715_
	);
	LUT2 #(
		.INIT('h4)
	) name8184 (
		_w8708_,
		_w8715_,
		_w8716_
	);
	LUT2 #(
		.INIT('h4)
	) name8185 (
		_w8691_,
		_w8716_,
		_w8717_
	);
	LUT2 #(
		.INIT('h2)
	) name8186 (
		\sa30_reg[1]/P0001 ,
		_w8717_,
		_w8718_
	);
	LUT2 #(
		.INIT('h8)
	) name8187 (
		\sa30_reg[7]/P0001 ,
		_w8698_,
		_w8719_
	);
	LUT2 #(
		.INIT('h8)
	) name8188 (
		_w8697_,
		_w8719_,
		_w8720_
	);
	LUT2 #(
		.INIT('h4)
	) name8189 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w8721_
	);
	LUT2 #(
		.INIT('h8)
	) name8190 (
		_w8682_,
		_w8721_,
		_w8722_
	);
	LUT2 #(
		.INIT('h1)
	) name8191 (
		\sa30_reg[2]/P0001 ,
		_w8722_,
		_w8723_
	);
	LUT2 #(
		.INIT('h4)
	) name8192 (
		\sa30_reg[3]/P0001 ,
		_w8701_,
		_w8724_
	);
	LUT2 #(
		.INIT('h2)
	) name8193 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w8725_
	);
	LUT2 #(
		.INIT('h4)
	) name8194 (
		\sa30_reg[6]/NET0131 ,
		_w8725_,
		_w8726_
	);
	LUT2 #(
		.INIT('h1)
	) name8195 (
		_w8722_,
		_w8724_,
		_w8727_
	);
	LUT2 #(
		.INIT('h4)
	) name8196 (
		_w8726_,
		_w8727_,
		_w8728_
	);
	LUT2 #(
		.INIT('h1)
	) name8197 (
		\sa30_reg[5]/P0001 ,
		_w8723_,
		_w8729_
	);
	LUT2 #(
		.INIT('h4)
	) name8198 (
		_w8728_,
		_w8729_,
		_w8730_
	);
	LUT2 #(
		.INIT('h1)
	) name8199 (
		_w8720_,
		_w8730_,
		_w8731_
	);
	LUT2 #(
		.INIT('h1)
	) name8200 (
		\sa30_reg[1]/P0001 ,
		_w8731_,
		_w8732_
	);
	LUT2 #(
		.INIT('h4)
	) name8201 (
		\sa30_reg[4]/P0001 ,
		_w8701_,
		_w8733_
	);
	LUT2 #(
		.INIT('h1)
	) name8202 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w8734_
	);
	LUT2 #(
		.INIT('h8)
	) name8203 (
		\sa30_reg[6]/NET0131 ,
		_w8721_,
		_w8735_
	);
	LUT2 #(
		.INIT('h1)
	) name8204 (
		_w8725_,
		_w8735_,
		_w8736_
	);
	LUT2 #(
		.INIT('h2)
	) name8205 (
		_w8734_,
		_w8736_,
		_w8737_
	);
	LUT2 #(
		.INIT('h1)
	) name8206 (
		_w8696_,
		_w8733_,
		_w8738_
	);
	LUT2 #(
		.INIT('h4)
	) name8207 (
		_w8737_,
		_w8738_,
		_w8739_
	);
	LUT2 #(
		.INIT('h2)
	) name8208 (
		\sa30_reg[2]/P0001 ,
		_w8739_,
		_w8740_
	);
	LUT2 #(
		.INIT('h4)
	) name8209 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w8741_
	);
	LUT2 #(
		.INIT('h8)
	) name8210 (
		_w8692_,
		_w8741_,
		_w8742_
	);
	LUT2 #(
		.INIT('h4)
	) name8211 (
		\sa30_reg[4]/P0001 ,
		_w8709_,
		_w8743_
	);
	LUT2 #(
		.INIT('h4)
	) name8212 (
		\sa30_reg[5]/P0001 ,
		_w8743_,
		_w8744_
	);
	LUT2 #(
		.INIT('h8)
	) name8213 (
		_w8695_,
		_w8734_,
		_w8745_
	);
	LUT2 #(
		.INIT('h1)
	) name8214 (
		_w8744_,
		_w8745_,
		_w8746_
	);
	LUT2 #(
		.INIT('h1)
	) name8215 (
		\sa30_reg[2]/P0001 ,
		_w8746_,
		_w8747_
	);
	LUT2 #(
		.INIT('h4)
	) name8216 (
		\sa30_reg[4]/P0001 ,
		_w8734_,
		_w8748_
	);
	LUT2 #(
		.INIT('h4)
	) name8217 (
		\sa30_reg[6]/NET0131 ,
		_w8748_,
		_w8749_
	);
	LUT2 #(
		.INIT('h1)
	) name8218 (
		_w8742_,
		_w8749_,
		_w8750_
	);
	LUT2 #(
		.INIT('h4)
	) name8219 (
		_w8747_,
		_w8750_,
		_w8751_
	);
	LUT2 #(
		.INIT('h4)
	) name8220 (
		_w8740_,
		_w8751_,
		_w8752_
	);
	LUT2 #(
		.INIT('h4)
	) name8221 (
		_w8732_,
		_w8752_,
		_w8753_
	);
	LUT2 #(
		.INIT('h4)
	) name8222 (
		_w8718_,
		_w8753_,
		_w8754_
	);
	LUT2 #(
		.INIT('h1)
	) name8223 (
		\sa30_reg[0]/P0002 ,
		_w8754_,
		_w8755_
	);
	LUT2 #(
		.INIT('h2)
	) name8224 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w8756_
	);
	LUT2 #(
		.INIT('h4)
	) name8225 (
		\sa30_reg[4]/P0001 ,
		_w8756_,
		_w8757_
	);
	LUT2 #(
		.INIT('h8)
	) name8226 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w8758_
	);
	LUT2 #(
		.INIT('h8)
	) name8227 (
		_w8756_,
		_w8758_,
		_w8759_
	);
	LUT2 #(
		.INIT('h8)
	) name8228 (
		_w8686_,
		_w8725_,
		_w8760_
	);
	LUT2 #(
		.INIT('h1)
	) name8229 (
		_w8759_,
		_w8760_,
		_w8761_
	);
	LUT2 #(
		.INIT('h4)
	) name8230 (
		_w8757_,
		_w8761_,
		_w8762_
	);
	LUT2 #(
		.INIT('h1)
	) name8231 (
		\sa30_reg[2]/P0001 ,
		_w8762_,
		_w8763_
	);
	LUT2 #(
		.INIT('h8)
	) name8232 (
		_w8705_,
		_w8725_,
		_w8764_
	);
	LUT2 #(
		.INIT('h8)
	) name8233 (
		_w8710_,
		_w8741_,
		_w8765_
	);
	LUT2 #(
		.INIT('h4)
	) name8234 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w8766_
	);
	LUT2 #(
		.INIT('h8)
	) name8235 (
		_w8734_,
		_w8766_,
		_w8767_
	);
	LUT2 #(
		.INIT('h4)
	) name8236 (
		\sa30_reg[3]/P0001 ,
		_w8767_,
		_w8768_
	);
	LUT2 #(
		.INIT('h8)
	) name8237 (
		_w8694_,
		_w8735_,
		_w8769_
	);
	LUT2 #(
		.INIT('h1)
	) name8238 (
		_w8768_,
		_w8769_,
		_w8770_
	);
	LUT2 #(
		.INIT('h2)
	) name8239 (
		\sa30_reg[2]/P0001 ,
		_w8770_,
		_w8771_
	);
	LUT2 #(
		.INIT('h2)
	) name8240 (
		\sa30_reg[1]/P0001 ,
		\sa30_reg[2]/P0001 ,
		_w8772_
	);
	LUT2 #(
		.INIT('h8)
	) name8241 (
		\sa30_reg[5]/P0001 ,
		_w8725_,
		_w8773_
	);
	LUT2 #(
		.INIT('h8)
	) name8242 (
		\sa30_reg[4]/P0001 ,
		_w8734_,
		_w8774_
	);
	LUT2 #(
		.INIT('h1)
	) name8243 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w8775_
	);
	LUT2 #(
		.INIT('h4)
	) name8244 (
		\sa30_reg[4]/P0001 ,
		_w8775_,
		_w8776_
	);
	LUT2 #(
		.INIT('h1)
	) name8245 (
		_w8773_,
		_w8774_,
		_w8777_
	);
	LUT2 #(
		.INIT('h4)
	) name8246 (
		_w8776_,
		_w8777_,
		_w8778_
	);
	LUT2 #(
		.INIT('h2)
	) name8247 (
		_w8772_,
		_w8778_,
		_w8779_
	);
	LUT2 #(
		.INIT('h8)
	) name8248 (
		_w8695_,
		_w8756_,
		_w8780_
	);
	LUT2 #(
		.INIT('h4)
	) name8249 (
		\sa30_reg[6]/NET0131 ,
		_w8780_,
		_w8781_
	);
	LUT2 #(
		.INIT('h4)
	) name8250 (
		\sa30_reg[4]/P0001 ,
		_w8683_,
		_w8782_
	);
	LUT2 #(
		.INIT('h4)
	) name8251 (
		\sa30_reg[7]/P0001 ,
		_w8721_,
		_w8783_
	);
	LUT2 #(
		.INIT('h8)
	) name8252 (
		_w8775_,
		_w8783_,
		_w8784_
	);
	LUT2 #(
		.INIT('h8)
	) name8253 (
		_w8694_,
		_w8721_,
		_w8785_
	);
	LUT2 #(
		.INIT('h4)
	) name8254 (
		\sa30_reg[6]/NET0131 ,
		_w8785_,
		_w8786_
	);
	LUT2 #(
		.INIT('h1)
	) name8255 (
		_w8781_,
		_w8782_,
		_w8787_
	);
	LUT2 #(
		.INIT('h1)
	) name8256 (
		_w8784_,
		_w8786_,
		_w8788_
	);
	LUT2 #(
		.INIT('h8)
	) name8257 (
		_w8787_,
		_w8788_,
		_w8789_
	);
	LUT2 #(
		.INIT('h2)
	) name8258 (
		\sa30_reg[1]/P0001 ,
		_w8789_,
		_w8790_
	);
	LUT2 #(
		.INIT('h8)
	) name8259 (
		_w8695_,
		_w8701_,
		_w8791_
	);
	LUT2 #(
		.INIT('h4)
	) name8260 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w8792_
	);
	LUT2 #(
		.INIT('h4)
	) name8261 (
		\sa30_reg[4]/P0001 ,
		_w8792_,
		_w8793_
	);
	LUT2 #(
		.INIT('h1)
	) name8262 (
		_w8791_,
		_w8793_,
		_w8794_
	);
	LUT2 #(
		.INIT('h2)
	) name8263 (
		\sa30_reg[2]/P0001 ,
		_w8794_,
		_w8795_
	);
	LUT2 #(
		.INIT('h8)
	) name8264 (
		_w8682_,
		_w8702_,
		_w8796_
	);
	LUT2 #(
		.INIT('h1)
	) name8265 (
		_w8705_,
		_w8796_,
		_w8797_
	);
	LUT2 #(
		.INIT('h1)
	) name8266 (
		\sa30_reg[2]/P0001 ,
		_w8797_,
		_w8798_
	);
	LUT2 #(
		.INIT('h1)
	) name8267 (
		_w8759_,
		_w8769_,
		_w8799_
	);
	LUT2 #(
		.INIT('h4)
	) name8268 (
		_w8795_,
		_w8799_,
		_w8800_
	);
	LUT2 #(
		.INIT('h4)
	) name8269 (
		_w8798_,
		_w8800_,
		_w8801_
	);
	LUT2 #(
		.INIT('h1)
	) name8270 (
		\sa30_reg[1]/P0001 ,
		_w8801_,
		_w8802_
	);
	LUT2 #(
		.INIT('h1)
	) name8271 (
		_w8764_,
		_w8765_,
		_w8803_
	);
	LUT2 #(
		.INIT('h4)
	) name8272 (
		_w8763_,
		_w8803_,
		_w8804_
	);
	LUT2 #(
		.INIT('h1)
	) name8273 (
		_w8771_,
		_w8779_,
		_w8805_
	);
	LUT2 #(
		.INIT('h8)
	) name8274 (
		_w8804_,
		_w8805_,
		_w8806_
	);
	LUT2 #(
		.INIT('h4)
	) name8275 (
		_w8790_,
		_w8806_,
		_w8807_
	);
	LUT2 #(
		.INIT('h4)
	) name8276 (
		_w8802_,
		_w8807_,
		_w8808_
	);
	LUT2 #(
		.INIT('h2)
	) name8277 (
		\sa30_reg[0]/P0002 ,
		_w8808_,
		_w8809_
	);
	LUT2 #(
		.INIT('h8)
	) name8278 (
		_w8698_,
		_w8701_,
		_w8810_
	);
	LUT2 #(
		.INIT('h8)
	) name8279 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w8811_
	);
	LUT2 #(
		.INIT('h2)
	) name8280 (
		\sa30_reg[3]/P0001 ,
		_w8684_,
		_w8812_
	);
	LUT2 #(
		.INIT('h4)
	) name8281 (
		\sa30_reg[5]/P0001 ,
		_w8682_,
		_w8813_
	);
	LUT2 #(
		.INIT('h4)
	) name8282 (
		\sa30_reg[5]/P0001 ,
		_w8686_,
		_w8814_
	);
	LUT2 #(
		.INIT('h1)
	) name8283 (
		_w8813_,
		_w8814_,
		_w8815_
	);
	LUT2 #(
		.INIT('h8)
	) name8284 (
		\sa30_reg[6]/NET0131 ,
		_w8694_,
		_w8816_
	);
	LUT2 #(
		.INIT('h1)
	) name8285 (
		\sa30_reg[3]/P0001 ,
		_w8816_,
		_w8817_
	);
	LUT2 #(
		.INIT('h8)
	) name8286 (
		_w8815_,
		_w8817_,
		_w8818_
	);
	LUT2 #(
		.INIT('h2)
	) name8287 (
		_w8811_,
		_w8812_,
		_w8819_
	);
	LUT2 #(
		.INIT('h4)
	) name8288 (
		_w8818_,
		_w8819_,
		_w8820_
	);
	LUT2 #(
		.INIT('h8)
	) name8289 (
		_w8695_,
		_w8697_,
		_w8821_
	);
	LUT2 #(
		.INIT('h4)
	) name8290 (
		\sa30_reg[7]/P0001 ,
		_w8821_,
		_w8822_
	);
	LUT2 #(
		.INIT('h8)
	) name8291 (
		\sa30_reg[4]/P0001 ,
		_w8710_,
		_w8823_
	);
	LUT2 #(
		.INIT('h8)
	) name8292 (
		_w8694_,
		_w8698_,
		_w8824_
	);
	LUT2 #(
		.INIT('h1)
	) name8293 (
		_w8822_,
		_w8824_,
		_w8825_
	);
	LUT2 #(
		.INIT('h4)
	) name8294 (
		_w8823_,
		_w8825_,
		_w8826_
	);
	LUT2 #(
		.INIT('h1)
	) name8295 (
		\sa30_reg[2]/P0001 ,
		_w8826_,
		_w8827_
	);
	LUT2 #(
		.INIT('h1)
	) name8296 (
		_w8810_,
		_w8820_,
		_w8828_
	);
	LUT2 #(
		.INIT('h4)
	) name8297 (
		_w8827_,
		_w8828_,
		_w8829_
	);
	LUT2 #(
		.INIT('h1)
	) name8298 (
		\sa30_reg[1]/P0001 ,
		_w8829_,
		_w8830_
	);
	LUT2 #(
		.INIT('h8)
	) name8299 (
		_w8726_,
		_w8756_,
		_w8831_
	);
	LUT2 #(
		.INIT('h4)
	) name8300 (
		\sa30_reg[2]/P0001 ,
		_w8831_,
		_w8832_
	);
	LUT2 #(
		.INIT('h1)
	) name8301 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		_w8833_
	);
	LUT2 #(
		.INIT('h8)
	) name8302 (
		_w8710_,
		_w8833_,
		_w8834_
	);
	LUT2 #(
		.INIT('h4)
	) name8303 (
		\sa30_reg[3]/P0001 ,
		_w8686_,
		_w8835_
	);
	LUT2 #(
		.INIT('h8)
	) name8304 (
		_w8811_,
		_w8835_,
		_w8836_
	);
	LUT2 #(
		.INIT('h8)
	) name8305 (
		\sa30_reg[5]/P0001 ,
		_w8836_,
		_w8837_
	);
	LUT2 #(
		.INIT('h4)
	) name8306 (
		\sa30_reg[7]/P0001 ,
		_w8725_,
		_w8838_
	);
	LUT2 #(
		.INIT('h4)
	) name8307 (
		\sa30_reg[5]/P0001 ,
		_w8838_,
		_w8839_
	);
	LUT2 #(
		.INIT('h4)
	) name8308 (
		\sa30_reg[6]/NET0131 ,
		_w8839_,
		_w8840_
	);
	LUT2 #(
		.INIT('h1)
	) name8309 (
		_w8742_,
		_w8837_,
		_w8841_
	);
	LUT2 #(
		.INIT('h4)
	) name8310 (
		_w8840_,
		_w8841_,
		_w8842_
	);
	LUT2 #(
		.INIT('h2)
	) name8311 (
		\sa30_reg[1]/P0001 ,
		_w8842_,
		_w8843_
	);
	LUT2 #(
		.INIT('h8)
	) name8312 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		_w8844_
	);
	LUT2 #(
		.INIT('h8)
	) name8313 (
		\sa30_reg[5]/P0001 ,
		_w8701_,
		_w8845_
	);
	LUT2 #(
		.INIT('h8)
	) name8314 (
		_w8844_,
		_w8845_,
		_w8846_
	);
	LUT2 #(
		.INIT('h8)
	) name8315 (
		\sa30_reg[4]/P0001 ,
		_w8846_,
		_w8847_
	);
	LUT2 #(
		.INIT('h1)
	) name8316 (
		_w8832_,
		_w8834_,
		_w8848_
	);
	LUT2 #(
		.INIT('h4)
	) name8317 (
		_w8847_,
		_w8848_,
		_w8849_
	);
	LUT2 #(
		.INIT('h4)
	) name8318 (
		_w8843_,
		_w8849_,
		_w8850_
	);
	LUT2 #(
		.INIT('h4)
	) name8319 (
		_w8830_,
		_w8850_,
		_w8851_
	);
	LUT2 #(
		.INIT('h4)
	) name8320 (
		_w8755_,
		_w8851_,
		_w8852_
	);
	LUT2 #(
		.INIT('h4)
	) name8321 (
		_w8809_,
		_w8852_,
		_w8853_
	);
	LUT2 #(
		.INIT('h2)
	) name8322 (
		\u0_w_reg[1][29]/P0002 ,
		_w8853_,
		_w8854_
	);
	LUT2 #(
		.INIT('h4)
	) name8323 (
		\u0_w_reg[1][29]/P0002 ,
		_w8853_,
		_w8855_
	);
	LUT2 #(
		.INIT('h1)
	) name8324 (
		_w8854_,
		_w8855_,
		_w8856_
	);
	LUT2 #(
		.INIT('h8)
	) name8325 (
		_w8681_,
		_w8856_,
		_w8857_
	);
	LUT2 #(
		.INIT('h1)
	) name8326 (
		_w8681_,
		_w8856_,
		_w8858_
	);
	LUT2 #(
		.INIT('h1)
	) name8327 (
		_w8857_,
		_w8858_,
		_w8859_
	);
	LUT2 #(
		.INIT('h4)
	) name8328 (
		_w8379_,
		_w8859_,
		_w8860_
	);
	LUT2 #(
		.INIT('h2)
	) name8329 (
		_w8379_,
		_w8859_,
		_w8861_
	);
	LUT2 #(
		.INIT('h1)
	) name8330 (
		\ld_r_reg/P0001 ,
		_w8860_,
		_w8862_
	);
	LUT2 #(
		.INIT('h4)
	) name8331 (
		_w8861_,
		_w8862_,
		_w8863_
	);
	LUT2 #(
		.INIT('h2)
	) name8332 (
		\text_in_r_reg[93]/P0001 ,
		\u0_w_reg[1][29]/P0002 ,
		_w8864_
	);
	LUT2 #(
		.INIT('h4)
	) name8333 (
		\text_in_r_reg[93]/P0001 ,
		\u0_w_reg[1][29]/P0002 ,
		_w8865_
	);
	LUT2 #(
		.INIT('h2)
	) name8334 (
		\ld_r_reg/P0001 ,
		_w8864_,
		_w8866_
	);
	LUT2 #(
		.INIT('h4)
	) name8335 (
		_w8865_,
		_w8866_,
		_w8867_
	);
	LUT2 #(
		.INIT('h1)
	) name8336 (
		_w8863_,
		_w8867_,
		_w8868_
	);
	LUT2 #(
		.INIT('h8)
	) name8337 (
		_w8694_,
		_w8725_,
		_w8869_
	);
	LUT2 #(
		.INIT('h1)
	) name8338 (
		_w8781_,
		_w8869_,
		_w8870_
	);
	LUT2 #(
		.INIT('h4)
	) name8339 (
		\sa30_reg[5]/P0001 ,
		_w8833_,
		_w8871_
	);
	LUT2 #(
		.INIT('h4)
	) name8340 (
		_w8766_,
		_w8871_,
		_w8872_
	);
	LUT2 #(
		.INIT('h8)
	) name8341 (
		\sa30_reg[4]/P0001 ,
		_w8686_,
		_w8873_
	);
	LUT2 #(
		.INIT('h4)
	) name8342 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w8874_
	);
	LUT2 #(
		.INIT('h8)
	) name8343 (
		_w8698_,
		_w8874_,
		_w8875_
	);
	LUT2 #(
		.INIT('h8)
	) name8344 (
		\sa30_reg[6]/NET0131 ,
		_w8875_,
		_w8876_
	);
	LUT2 #(
		.INIT('h1)
	) name8345 (
		_w8693_,
		_w8873_,
		_w8877_
	);
	LUT2 #(
		.INIT('h4)
	) name8346 (
		_w8876_,
		_w8877_,
		_w8878_
	);
	LUT2 #(
		.INIT('h2)
	) name8347 (
		\sa30_reg[2]/P0001 ,
		_w8878_,
		_w8879_
	);
	LUT2 #(
		.INIT('h2)
	) name8348 (
		_w8870_,
		_w8872_,
		_w8880_
	);
	LUT2 #(
		.INIT('h4)
	) name8349 (
		_w8879_,
		_w8880_,
		_w8881_
	);
	LUT2 #(
		.INIT('h2)
	) name8350 (
		\sa30_reg[1]/P0001 ,
		_w8881_,
		_w8882_
	);
	LUT2 #(
		.INIT('h8)
	) name8351 (
		_w8756_,
		_w8766_,
		_w8883_
	);
	LUT2 #(
		.INIT('h4)
	) name8352 (
		\sa30_reg[3]/P0001 ,
		_w8684_,
		_w8884_
	);
	LUT2 #(
		.INIT('h8)
	) name8353 (
		\sa30_reg[4]/P0001 ,
		_w8884_,
		_w8885_
	);
	LUT2 #(
		.INIT('h1)
	) name8354 (
		_w8883_,
		_w8885_,
		_w8886_
	);
	LUT2 #(
		.INIT('h1)
	) name8355 (
		\sa30_reg[2]/P0001 ,
		_w8886_,
		_w8887_
	);
	LUT2 #(
		.INIT('h8)
	) name8356 (
		\sa30_reg[3]/P0001 ,
		_w8686_,
		_w8888_
	);
	LUT2 #(
		.INIT('h8)
	) name8357 (
		\sa30_reg[4]/P0001 ,
		_w8888_,
		_w8889_
	);
	LUT2 #(
		.INIT('h1)
	) name8358 (
		_w8769_,
		_w8889_,
		_w8890_
	);
	LUT2 #(
		.INIT('h1)
	) name8359 (
		_w8749_,
		_w8796_,
		_w8891_
	);
	LUT2 #(
		.INIT('h8)
	) name8360 (
		_w8890_,
		_w8891_,
		_w8892_
	);
	LUT2 #(
		.INIT('h2)
	) name8361 (
		\sa30_reg[2]/P0001 ,
		_w8892_,
		_w8893_
	);
	LUT2 #(
		.INIT('h4)
	) name8362 (
		\sa30_reg[3]/P0001 ,
		_w8845_,
		_w8894_
	);
	LUT2 #(
		.INIT('h4)
	) name8363 (
		\sa30_reg[2]/P0001 ,
		_w8894_,
		_w8895_
	);
	LUT2 #(
		.INIT('h8)
	) name8364 (
		\sa30_reg[7]/P0001 ,
		_w8695_,
		_w8896_
	);
	LUT2 #(
		.INIT('h1)
	) name8365 (
		_w8814_,
		_w8896_,
		_w8897_
	);
	LUT2 #(
		.INIT('h2)
	) name8366 (
		\sa30_reg[2]/P0001 ,
		_w8897_,
		_w8898_
	);
	LUT2 #(
		.INIT('h8)
	) name8367 (
		\sa30_reg[7]/P0001 ,
		_w8685_,
		_w8899_
	);
	LUT2 #(
		.INIT('h1)
	) name8368 (
		_w8895_,
		_w8899_,
		_w8900_
	);
	LUT2 #(
		.INIT('h4)
	) name8369 (
		_w8898_,
		_w8900_,
		_w8901_
	);
	LUT2 #(
		.INIT('h4)
	) name8370 (
		_w8747_,
		_w8901_,
		_w8902_
	);
	LUT2 #(
		.INIT('h1)
	) name8371 (
		\sa30_reg[1]/P0001 ,
		_w8902_,
		_w8903_
	);
	LUT2 #(
		.INIT('h1)
	) name8372 (
		_w8887_,
		_w8893_,
		_w8904_
	);
	LUT2 #(
		.INIT('h4)
	) name8373 (
		_w8882_,
		_w8904_,
		_w8905_
	);
	LUT2 #(
		.INIT('h4)
	) name8374 (
		_w8903_,
		_w8905_,
		_w8906_
	);
	LUT2 #(
		.INIT('h2)
	) name8375 (
		\sa30_reg[0]/P0002 ,
		_w8906_,
		_w8907_
	);
	LUT2 #(
		.INIT('h2)
	) name8376 (
		\sa30_reg[4]/P0001 ,
		_w8709_,
		_w8908_
	);
	LUT2 #(
		.INIT('h4)
	) name8377 (
		_w8701_,
		_w8702_,
		_w8909_
	);
	LUT2 #(
		.INIT('h4)
	) name8378 (
		_w8908_,
		_w8909_,
		_w8910_
	);
	LUT2 #(
		.INIT('h1)
	) name8379 (
		_w8705_,
		_w8775_,
		_w8911_
	);
	LUT2 #(
		.INIT('h2)
	) name8380 (
		_w8721_,
		_w8911_,
		_w8912_
	);
	LUT2 #(
		.INIT('h1)
	) name8381 (
		\sa30_reg[2]/P0001 ,
		_w8910_,
		_w8913_
	);
	LUT2 #(
		.INIT('h4)
	) name8382 (
		_w8912_,
		_w8913_,
		_w8914_
	);
	LUT2 #(
		.INIT('h8)
	) name8383 (
		_w8710_,
		_w8721_,
		_w8915_
	);
	LUT2 #(
		.INIT('h8)
	) name8384 (
		_w8698_,
		_w8775_,
		_w8916_
	);
	LUT2 #(
		.INIT('h2)
	) name8385 (
		\sa30_reg[2]/P0001 ,
		_w8916_,
		_w8917_
	);
	LUT2 #(
		.INIT('h4)
	) name8386 (
		_w8915_,
		_w8917_,
		_w8918_
	);
	LUT2 #(
		.INIT('h1)
	) name8387 (
		_w8914_,
		_w8918_,
		_w8919_
	);
	LUT2 #(
		.INIT('h8)
	) name8388 (
		_w8682_,
		_w8698_,
		_w8920_
	);
	LUT2 #(
		.INIT('h4)
	) name8389 (
		\sa30_reg[2]/P0001 ,
		_w8896_,
		_w8921_
	);
	LUT2 #(
		.INIT('h8)
	) name8390 (
		_w8725_,
		_w8874_,
		_w8922_
	);
	LUT2 #(
		.INIT('h1)
	) name8391 (
		\sa30_reg[1]/P0001 ,
		_w8883_,
		_w8923_
	);
	LUT2 #(
		.INIT('h1)
	) name8392 (
		_w8920_,
		_w8922_,
		_w8924_
	);
	LUT2 #(
		.INIT('h8)
	) name8393 (
		_w8923_,
		_w8924_,
		_w8925_
	);
	LUT2 #(
		.INIT('h1)
	) name8394 (
		_w8846_,
		_w8915_,
		_w8926_
	);
	LUT2 #(
		.INIT('h4)
	) name8395 (
		_w8921_,
		_w8926_,
		_w8927_
	);
	LUT2 #(
		.INIT('h8)
	) name8396 (
		_w8925_,
		_w8927_,
		_w8928_
	);
	LUT2 #(
		.INIT('h2)
	) name8397 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		_w8929_
	);
	LUT2 #(
		.INIT('h8)
	) name8398 (
		\sa30_reg[4]/P0001 ,
		_w8694_,
		_w8930_
	);
	LUT2 #(
		.INIT('h1)
	) name8399 (
		_w8748_,
		_w8930_,
		_w8931_
	);
	LUT2 #(
		.INIT('h2)
	) name8400 (
		_w8929_,
		_w8931_,
		_w8932_
	);
	LUT2 #(
		.INIT('h4)
	) name8401 (
		\sa30_reg[2]/P0001 ,
		_w8749_,
		_w8933_
	);
	LUT2 #(
		.INIT('h2)
	) name8402 (
		\sa30_reg[1]/P0001 ,
		_w8822_,
		_w8934_
	);
	LUT2 #(
		.INIT('h4)
	) name8403 (
		_w8932_,
		_w8934_,
		_w8935_
	);
	LUT2 #(
		.INIT('h4)
	) name8404 (
		_w8933_,
		_w8935_,
		_w8936_
	);
	LUT2 #(
		.INIT('h1)
	) name8405 (
		_w8928_,
		_w8936_,
		_w8937_
	);
	LUT2 #(
		.INIT('h1)
	) name8406 (
		_w8919_,
		_w8937_,
		_w8938_
	);
	LUT2 #(
		.INIT('h1)
	) name8407 (
		\sa30_reg[0]/P0002 ,
		_w8938_,
		_w8939_
	);
	LUT2 #(
		.INIT('h4)
	) name8408 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		_w8940_
	);
	LUT2 #(
		.INIT('h8)
	) name8409 (
		_w8899_,
		_w8940_,
		_w8941_
	);
	LUT2 #(
		.INIT('h8)
	) name8410 (
		_w8772_,
		_w8831_,
		_w8942_
	);
	LUT2 #(
		.INIT('h4)
	) name8411 (
		\sa30_reg[7]/P0001 ,
		_w8698_,
		_w8943_
	);
	LUT2 #(
		.INIT('h1)
	) name8412 (
		_w8774_,
		_w8869_,
		_w8944_
	);
	LUT2 #(
		.INIT('h4)
	) name8413 (
		_w8943_,
		_w8944_,
		_w8945_
	);
	LUT2 #(
		.INIT('h8)
	) name8414 (
		\sa30_reg[1]/P0001 ,
		\sa30_reg[2]/P0001 ,
		_w8946_
	);
	LUT2 #(
		.INIT('h4)
	) name8415 (
		\sa30_reg[6]/NET0131 ,
		_w8946_,
		_w8947_
	);
	LUT2 #(
		.INIT('h4)
	) name8416 (
		_w8945_,
		_w8947_,
		_w8948_
	);
	LUT2 #(
		.INIT('h8)
	) name8417 (
		_w8775_,
		_w8943_,
		_w8949_
	);
	LUT2 #(
		.INIT('h4)
	) name8418 (
		\sa30_reg[5]/P0001 ,
		_w8701_,
		_w8950_
	);
	LUT2 #(
		.INIT('h4)
	) name8419 (
		\sa30_reg[3]/P0001 ,
		_w8950_,
		_w8951_
	);
	LUT2 #(
		.INIT('h8)
	) name8420 (
		_w8694_,
		_w8766_,
		_w8952_
	);
	LUT2 #(
		.INIT('h4)
	) name8421 (
		\sa30_reg[7]/P0001 ,
		_w8726_,
		_w8953_
	);
	LUT2 #(
		.INIT('h1)
	) name8422 (
		_w8952_,
		_w8953_,
		_w8954_
	);
	LUT2 #(
		.INIT('h1)
	) name8423 (
		\sa30_reg[1]/P0001 ,
		_w8954_,
		_w8955_
	);
	LUT2 #(
		.INIT('h8)
	) name8424 (
		_w8695_,
		_w8814_,
		_w8956_
	);
	LUT2 #(
		.INIT('h1)
	) name8425 (
		_w8951_,
		_w8956_,
		_w8957_
	);
	LUT2 #(
		.INIT('h4)
	) name8426 (
		_w8955_,
		_w8957_,
		_w8958_
	);
	LUT2 #(
		.INIT('h2)
	) name8427 (
		\sa30_reg[2]/P0001 ,
		_w8958_,
		_w8959_
	);
	LUT2 #(
		.INIT('h2)
	) name8428 (
		_w8692_,
		_w8698_,
		_w8960_
	);
	LUT2 #(
		.INIT('h4)
	) name8429 (
		\sa30_reg[5]/P0001 ,
		_w8873_,
		_w8961_
	);
	LUT2 #(
		.INIT('h1)
	) name8430 (
		_w8960_,
		_w8961_,
		_w8962_
	);
	LUT2 #(
		.INIT('h1)
	) name8431 (
		\sa30_reg[2]/P0001 ,
		_w8962_,
		_w8963_
	);
	LUT2 #(
		.INIT('h8)
	) name8432 (
		_w8682_,
		_w8695_,
		_w8964_
	);
	LUT2 #(
		.INIT('h1)
	) name8433 (
		_w8699_,
		_w8964_,
		_w8965_
	);
	LUT2 #(
		.INIT('h4)
	) name8434 (
		_w8963_,
		_w8965_,
		_w8966_
	);
	LUT2 #(
		.INIT('h1)
	) name8435 (
		\sa30_reg[1]/P0001 ,
		_w8966_,
		_w8967_
	);
	LUT2 #(
		.INIT('h1)
	) name8436 (
		_w8941_,
		_w8949_,
		_w8968_
	);
	LUT2 #(
		.INIT('h4)
	) name8437 (
		_w8942_,
		_w8968_,
		_w8969_
	);
	LUT2 #(
		.INIT('h4)
	) name8438 (
		_w8948_,
		_w8969_,
		_w8970_
	);
	LUT2 #(
		.INIT('h4)
	) name8439 (
		_w8959_,
		_w8970_,
		_w8971_
	);
	LUT2 #(
		.INIT('h4)
	) name8440 (
		_w8967_,
		_w8971_,
		_w8972_
	);
	LUT2 #(
		.INIT('h4)
	) name8441 (
		_w8939_,
		_w8972_,
		_w8973_
	);
	LUT2 #(
		.INIT('h4)
	) name8442 (
		_w8907_,
		_w8973_,
		_w8974_
	);
	LUT2 #(
		.INIT('h2)
	) name8443 (
		\u0_w_reg[1][30]/P0001 ,
		_w8974_,
		_w8975_
	);
	LUT2 #(
		.INIT('h4)
	) name8444 (
		\u0_w_reg[1][30]/P0001 ,
		_w8974_,
		_w8976_
	);
	LUT2 #(
		.INIT('h1)
	) name8445 (
		_w8975_,
		_w8976_,
		_w8977_
	);
	LUT2 #(
		.INIT('h1)
	) name8446 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		_w8978_
	);
	LUT2 #(
		.INIT('h1)
	) name8447 (
		\sa12_reg[5]/P0001 ,
		_w8068_,
		_w8979_
	);
	LUT2 #(
		.INIT('h8)
	) name8448 (
		_w8978_,
		_w8979_,
		_w8980_
	);
	LUT2 #(
		.INIT('h8)
	) name8449 (
		_w8084_,
		_w8202_,
		_w8981_
	);
	LUT2 #(
		.INIT('h1)
	) name8450 (
		_w8061_,
		_w8388_,
		_w8982_
	);
	LUT2 #(
		.INIT('h4)
	) name8451 (
		_w8981_,
		_w8982_,
		_w8983_
	);
	LUT2 #(
		.INIT('h2)
	) name8452 (
		\sa12_reg[2]/P0001 ,
		_w8983_,
		_w8984_
	);
	LUT2 #(
		.INIT('h8)
	) name8453 (
		_w8078_,
		_w8161_,
		_w8985_
	);
	LUT2 #(
		.INIT('h1)
	) name8454 (
		_w8460_,
		_w8985_,
		_w8986_
	);
	LUT2 #(
		.INIT('h4)
	) name8455 (
		_w8980_,
		_w8986_,
		_w8987_
	);
	LUT2 #(
		.INIT('h4)
	) name8456 (
		_w8984_,
		_w8987_,
		_w8988_
	);
	LUT2 #(
		.INIT('h2)
	) name8457 (
		\sa12_reg[1]/P0001 ,
		_w8988_,
		_w8989_
	);
	LUT2 #(
		.INIT('h8)
	) name8458 (
		_w8065_,
		_w8498_,
		_w8990_
	);
	LUT2 #(
		.INIT('h1)
	) name8459 (
		_w8380_,
		_w8990_,
		_w8991_
	);
	LUT2 #(
		.INIT('h1)
	) name8460 (
		\sa12_reg[2]/P0001 ,
		_w8991_,
		_w8992_
	);
	LUT2 #(
		.INIT('h1)
	) name8461 (
		_w8181_,
		_w8433_,
		_w8993_
	);
	LUT2 #(
		.INIT('h1)
	) name8462 (
		_w8127_,
		_w8425_,
		_w8994_
	);
	LUT2 #(
		.INIT('h8)
	) name8463 (
		_w8993_,
		_w8994_,
		_w8995_
	);
	LUT2 #(
		.INIT('h2)
	) name8464 (
		\sa12_reg[2]/P0001 ,
		_w8995_,
		_w8996_
	);
	LUT2 #(
		.INIT('h1)
	) name8465 (
		\sa12_reg[2]/P0001 ,
		_w8087_,
		_w8997_
	);
	LUT2 #(
		.INIT('h2)
	) name8466 (
		\sa12_reg[2]/P0001 ,
		_w8081_,
		_w8998_
	);
	LUT2 #(
		.INIT('h4)
	) name8467 (
		_w8412_,
		_w8998_,
		_w8999_
	);
	LUT2 #(
		.INIT('h1)
	) name8468 (
		_w8997_,
		_w8999_,
		_w9000_
	);
	LUT2 #(
		.INIT('h1)
	) name8469 (
		_w8166_,
		_w8424_,
		_w9001_
	);
	LUT2 #(
		.INIT('h4)
	) name8470 (
		_w9000_,
		_w9001_,
		_w9002_
	);
	LUT2 #(
		.INIT('h1)
	) name8471 (
		\sa12_reg[1]/P0001 ,
		_w9002_,
		_w9003_
	);
	LUT2 #(
		.INIT('h1)
	) name8472 (
		_w8992_,
		_w8996_,
		_w9004_
	);
	LUT2 #(
		.INIT('h4)
	) name8473 (
		_w8989_,
		_w9004_,
		_w9005_
	);
	LUT2 #(
		.INIT('h4)
	) name8474 (
		_w9003_,
		_w9005_,
		_w9006_
	);
	LUT2 #(
		.INIT('h2)
	) name8475 (
		\sa12_reg[0]/P0001 ,
		_w9006_,
		_w9007_
	);
	LUT2 #(
		.INIT('h1)
	) name8476 (
		_w8165_,
		_w8414_,
		_w9008_
	);
	LUT2 #(
		.INIT('h2)
	) name8477 (
		_w8059_,
		_w9008_,
		_w9009_
	);
	LUT2 #(
		.INIT('h8)
	) name8478 (
		_w8142_,
		_w8162_,
		_w9010_
	);
	LUT2 #(
		.INIT('h2)
	) name8479 (
		\sa12_reg[1]/P0001 ,
		_w8103_,
		_w9011_
	);
	LUT2 #(
		.INIT('h4)
	) name8480 (
		_w9010_,
		_w9011_,
		_w9012_
	);
	LUT2 #(
		.INIT('h4)
	) name8481 (
		_w9009_,
		_w9012_,
		_w9013_
	);
	LUT2 #(
		.INIT('h8)
	) name8482 (
		_w8080_,
		_w8155_,
		_w9014_
	);
	LUT2 #(
		.INIT('h4)
	) name8483 (
		\sa12_reg[6]/NET0131 ,
		_w8085_,
		_w9015_
	);
	LUT2 #(
		.INIT('h1)
	) name8484 (
		\sa12_reg[1]/P0001 ,
		_w8112_,
		_w9016_
	);
	LUT2 #(
		.INIT('h1)
	) name8485 (
		_w8990_,
		_w9014_,
		_w9017_
	);
	LUT2 #(
		.INIT('h8)
	) name8486 (
		_w9016_,
		_w9017_,
		_w9018_
	);
	LUT2 #(
		.INIT('h1)
	) name8487 (
		_w8058_,
		_w8177_,
		_w9019_
	);
	LUT2 #(
		.INIT('h4)
	) name8488 (
		_w9015_,
		_w9019_,
		_w9020_
	);
	LUT2 #(
		.INIT('h8)
	) name8489 (
		_w9018_,
		_w9020_,
		_w9021_
	);
	LUT2 #(
		.INIT('h1)
	) name8490 (
		_w9013_,
		_w9021_,
		_w9022_
	);
	LUT2 #(
		.INIT('h2)
	) name8491 (
		\sa12_reg[2]/P0001 ,
		_w8117_,
		_w9023_
	);
	LUT2 #(
		.INIT('h4)
	) name8492 (
		_w8177_,
		_w9023_,
		_w9024_
	);
	LUT2 #(
		.INIT('h8)
	) name8493 (
		\sa12_reg[4]/P0001 ,
		_w8082_,
		_w9025_
	);
	LUT2 #(
		.INIT('h1)
	) name8494 (
		_w8116_,
		_w9025_,
		_w9026_
	);
	LUT2 #(
		.INIT('h1)
	) name8495 (
		_w8180_,
		_w9026_,
		_w9027_
	);
	LUT2 #(
		.INIT('h2)
	) name8496 (
		_w8137_,
		_w8495_,
		_w9028_
	);
	LUT2 #(
		.INIT('h4)
	) name8497 (
		_w9027_,
		_w9028_,
		_w9029_
	);
	LUT2 #(
		.INIT('h1)
	) name8498 (
		_w9024_,
		_w9029_,
		_w9030_
	);
	LUT2 #(
		.INIT('h1)
	) name8499 (
		_w9022_,
		_w9030_,
		_w9031_
	);
	LUT2 #(
		.INIT('h1)
	) name8500 (
		\sa12_reg[0]/P0001 ,
		_w9031_,
		_w9032_
	);
	LUT2 #(
		.INIT('h8)
	) name8501 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[2]/P0001 ,
		_w9033_
	);
	LUT2 #(
		.INIT('h8)
	) name8502 (
		\sa12_reg[4]/P0001 ,
		_w8142_,
		_w9034_
	);
	LUT2 #(
		.INIT('h8)
	) name8503 (
		\sa12_reg[5]/P0001 ,
		_w8381_,
		_w9035_
	);
	LUT2 #(
		.INIT('h4)
	) name8504 (
		\sa12_reg[4]/P0001 ,
		_w9035_,
		_w9036_
	);
	LUT2 #(
		.INIT('h1)
	) name8505 (
		_w8485_,
		_w9034_,
		_w9037_
	);
	LUT2 #(
		.INIT('h4)
	) name8506 (
		_w9036_,
		_w9037_,
		_w9038_
	);
	LUT2 #(
		.INIT('h2)
	) name8507 (
		_w9033_,
		_w9038_,
		_w9039_
	);
	LUT2 #(
		.INIT('h8)
	) name8508 (
		_w8150_,
		_w8455_,
		_w9040_
	);
	LUT2 #(
		.INIT('h8)
	) name8509 (
		_w8155_,
		_w8166_,
		_w9041_
	);
	LUT2 #(
		.INIT('h8)
	) name8510 (
		_w8069_,
		_w8075_,
		_w9042_
	);
	LUT2 #(
		.INIT('h8)
	) name8511 (
		_w8066_,
		_w9042_,
		_w9043_
	);
	LUT2 #(
		.INIT('h8)
	) name8512 (
		_w8068_,
		_w8161_,
		_w9044_
	);
	LUT2 #(
		.INIT('h1)
	) name8513 (
		_w8195_,
		_w9044_,
		_w9045_
	);
	LUT2 #(
		.INIT('h2)
	) name8514 (
		\sa12_reg[2]/P0001 ,
		_w9045_,
		_w9046_
	);
	LUT2 #(
		.INIT('h8)
	) name8515 (
		_w8126_,
		_w8180_,
		_w9047_
	);
	LUT2 #(
		.INIT('h4)
	) name8516 (
		_w8104_,
		_w8185_,
		_w9048_
	);
	LUT2 #(
		.INIT('h8)
	) name8517 (
		_w8069_,
		_w8390_,
		_w9049_
	);
	LUT2 #(
		.INIT('h1)
	) name8518 (
		_w9048_,
		_w9049_,
		_w9050_
	);
	LUT2 #(
		.INIT('h1)
	) name8519 (
		\sa12_reg[2]/P0001 ,
		_w9050_,
		_w9051_
	);
	LUT2 #(
		.INIT('h1)
	) name8520 (
		_w8394_,
		_w9047_,
		_w9052_
	);
	LUT2 #(
		.INIT('h4)
	) name8521 (
		_w9046_,
		_w9052_,
		_w9053_
	);
	LUT2 #(
		.INIT('h4)
	) name8522 (
		_w9051_,
		_w9053_,
		_w9054_
	);
	LUT2 #(
		.INIT('h1)
	) name8523 (
		\sa12_reg[1]/P0001 ,
		_w9054_,
		_w9055_
	);
	LUT2 #(
		.INIT('h1)
	) name8524 (
		_w8118_,
		_w9043_,
		_w9056_
	);
	LUT2 #(
		.INIT('h4)
	) name8525 (
		_w8408_,
		_w9056_,
		_w9057_
	);
	LUT2 #(
		.INIT('h1)
	) name8526 (
		_w9040_,
		_w9041_,
		_w9058_
	);
	LUT2 #(
		.INIT('h8)
	) name8527 (
		_w9057_,
		_w9058_,
		_w9059_
	);
	LUT2 #(
		.INIT('h4)
	) name8528 (
		_w9039_,
		_w9059_,
		_w9060_
	);
	LUT2 #(
		.INIT('h4)
	) name8529 (
		_w9055_,
		_w9060_,
		_w9061_
	);
	LUT2 #(
		.INIT('h4)
	) name8530 (
		_w9032_,
		_w9061_,
		_w9062_
	);
	LUT2 #(
		.INIT('h4)
	) name8531 (
		_w9007_,
		_w9062_,
		_w9063_
	);
	LUT2 #(
		.INIT('h4)
	) name8532 (
		\sa23_reg[3]/P0001 ,
		_w8631_,
		_w9064_
	);
	LUT2 #(
		.INIT('h4)
	) name8533 (
		\sa23_reg[2]/P0001 ,
		_w9064_,
		_w9065_
	);
	LUT2 #(
		.INIT('h8)
	) name8534 (
		\sa23_reg[3]/P0001 ,
		_w8569_,
		_w9066_
	);
	LUT2 #(
		.INIT('h1)
	) name8535 (
		_w8655_,
		_w9066_,
		_w9067_
	);
	LUT2 #(
		.INIT('h2)
	) name8536 (
		\sa23_reg[2]/P0001 ,
		_w9067_,
		_w9068_
	);
	LUT2 #(
		.INIT('h1)
	) name8537 (
		_w8567_,
		_w8570_,
		_w9069_
	);
	LUT2 #(
		.INIT('h1)
	) name8538 (
		_w9065_,
		_w9068_,
		_w9070_
	);
	LUT2 #(
		.INIT('h8)
	) name8539 (
		_w9069_,
		_w9070_,
		_w9071_
	);
	LUT2 #(
		.INIT('h1)
	) name8540 (
		\sa23_reg[1]/P0001 ,
		_w9071_,
		_w9072_
	);
	LUT2 #(
		.INIT('h8)
	) name8541 (
		\sa23_reg[4]/P0001 ,
		_w8513_,
		_w9073_
	);
	LUT2 #(
		.INIT('h8)
	) name8542 (
		_w8525_,
		_w8603_,
		_w9074_
	);
	LUT2 #(
		.INIT('h1)
	) name8543 (
		_w8520_,
		_w9073_,
		_w9075_
	);
	LUT2 #(
		.INIT('h4)
	) name8544 (
		_w9074_,
		_w9075_,
		_w9076_
	);
	LUT2 #(
		.INIT('h2)
	) name8545 (
		\sa23_reg[2]/P0001 ,
		_w9076_,
		_w9077_
	);
	LUT2 #(
		.INIT('h8)
	) name8546 (
		_w8531_,
		_w8572_,
		_w9078_
	);
	LUT2 #(
		.INIT('h1)
	) name8547 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		_w9079_
	);
	LUT2 #(
		.INIT('h8)
	) name8548 (
		_w8594_,
		_w9079_,
		_w9080_
	);
	LUT2 #(
		.INIT('h1)
	) name8549 (
		_w8632_,
		_w9078_,
		_w9081_
	);
	LUT2 #(
		.INIT('h4)
	) name8550 (
		_w9080_,
		_w9081_,
		_w9082_
	);
	LUT2 #(
		.INIT('h4)
	) name8551 (
		_w9077_,
		_w9082_,
		_w9083_
	);
	LUT2 #(
		.INIT('h2)
	) name8552 (
		\sa23_reg[1]/P0001 ,
		_w9083_,
		_w9084_
	);
	LUT2 #(
		.INIT('h8)
	) name8553 (
		_w8521_,
		_w8577_,
		_w9085_
	);
	LUT2 #(
		.INIT('h1)
	) name8554 (
		_w8510_,
		_w9085_,
		_w9086_
	);
	LUT2 #(
		.INIT('h1)
	) name8555 (
		\sa23_reg[2]/P0001 ,
		_w9086_,
		_w9087_
	);
	LUT2 #(
		.INIT('h1)
	) name8556 (
		_w8604_,
		_w8641_,
		_w9088_
	);
	LUT2 #(
		.INIT('h1)
	) name8557 (
		_w8568_,
		_w8615_,
		_w9089_
	);
	LUT2 #(
		.INIT('h8)
	) name8558 (
		_w9088_,
		_w9089_,
		_w9090_
	);
	LUT2 #(
		.INIT('h2)
	) name8559 (
		\sa23_reg[2]/P0001 ,
		_w9090_,
		_w9091_
	);
	LUT2 #(
		.INIT('h1)
	) name8560 (
		_w9087_,
		_w9091_,
		_w9092_
	);
	LUT2 #(
		.INIT('h4)
	) name8561 (
		_w9072_,
		_w9092_,
		_w9093_
	);
	LUT2 #(
		.INIT('h4)
	) name8562 (
		_w9084_,
		_w9093_,
		_w9094_
	);
	LUT2 #(
		.INIT('h2)
	) name8563 (
		\sa23_reg[0]/P0001 ,
		_w9094_,
		_w9095_
	);
	LUT2 #(
		.INIT('h8)
	) name8564 (
		\sa23_reg[7]/NET0131 ,
		_w8588_,
		_w9096_
	);
	LUT2 #(
		.INIT('h4)
	) name8565 (
		\sa23_reg[5]/P0001 ,
		_w9096_,
		_w9097_
	);
	LUT2 #(
		.INIT('h1)
	) name8566 (
		\sa23_reg[2]/P0001 ,
		_w9097_,
		_w9098_
	);
	LUT2 #(
		.INIT('h8)
	) name8567 (
		\sa23_reg[4]/P0001 ,
		_w8547_,
		_w9099_
	);
	LUT2 #(
		.INIT('h4)
	) name8568 (
		_w8528_,
		_w8529_,
		_w9100_
	);
	LUT2 #(
		.INIT('h8)
	) name8569 (
		_w8574_,
		_w8589_,
		_w9101_
	);
	LUT2 #(
		.INIT('h1)
	) name8570 (
		_w9099_,
		_w9100_,
		_w9102_
	);
	LUT2 #(
		.INIT('h4)
	) name8571 (
		_w9101_,
		_w9102_,
		_w9103_
	);
	LUT2 #(
		.INIT('h1)
	) name8572 (
		_w8537_,
		_w9103_,
		_w9104_
	);
	LUT2 #(
		.INIT('h2)
	) name8573 (
		_w9098_,
		_w9104_,
		_w9105_
	);
	LUT2 #(
		.INIT('h8)
	) name8574 (
		_w8522_,
		_w8547_,
		_w9106_
	);
	LUT2 #(
		.INIT('h4)
	) name8575 (
		\sa23_reg[3]/P0001 ,
		_w8602_,
		_w9107_
	);
	LUT2 #(
		.INIT('h2)
	) name8576 (
		\sa23_reg[2]/P0001 ,
		_w9106_,
		_w9108_
	);
	LUT2 #(
		.INIT('h4)
	) name8577 (
		_w9107_,
		_w9108_,
		_w9109_
	);
	LUT2 #(
		.INIT('h1)
	) name8578 (
		_w9105_,
		_w9109_,
		_w9110_
	);
	LUT2 #(
		.INIT('h4)
	) name8579 (
		\sa23_reg[2]/P0001 ,
		_w8568_,
		_w9111_
	);
	LUT2 #(
		.INIT('h2)
	) name8580 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		_w9112_
	);
	LUT2 #(
		.INIT('h8)
	) name8581 (
		\sa23_reg[4]/P0001 ,
		_w8531_,
		_w9113_
	);
	LUT2 #(
		.INIT('h4)
	) name8582 (
		\sa23_reg[4]/P0001 ,
		_w8564_,
		_w9114_
	);
	LUT2 #(
		.INIT('h1)
	) name8583 (
		_w9113_,
		_w9114_,
		_w9115_
	);
	LUT2 #(
		.INIT('h2)
	) name8584 (
		_w9112_,
		_w9115_,
		_w9116_
	);
	LUT2 #(
		.INIT('h8)
	) name8585 (
		_w8537_,
		_w8614_,
		_w9117_
	);
	LUT2 #(
		.INIT('h1)
	) name8586 (
		_w9111_,
		_w9117_,
		_w9118_
	);
	LUT2 #(
		.INIT('h4)
	) name8587 (
		_w9116_,
		_w9118_,
		_w9119_
	);
	LUT2 #(
		.INIT('h2)
	) name8588 (
		\sa23_reg[1]/P0001 ,
		_w9119_,
		_w9120_
	);
	LUT2 #(
		.INIT('h1)
	) name8589 (
		_w9110_,
		_w9120_,
		_w9121_
	);
	LUT2 #(
		.INIT('h1)
	) name8590 (
		\sa23_reg[0]/P0001 ,
		_w9121_,
		_w9122_
	);
	LUT2 #(
		.INIT('h1)
	) name8591 (
		_w8523_,
		_w9078_,
		_w9123_
	);
	LUT2 #(
		.INIT('h1)
	) name8592 (
		\sa23_reg[6]/NET0131 ,
		_w9123_,
		_w9124_
	);
	LUT2 #(
		.INIT('h4)
	) name8593 (
		\sa23_reg[7]/NET0131 ,
		_w9099_,
		_w9125_
	);
	LUT2 #(
		.INIT('h1)
	) name8594 (
		_w9124_,
		_w9125_,
		_w9126_
	);
	LUT2 #(
		.INIT('h2)
	) name8595 (
		\sa23_reg[1]/P0001 ,
		_w9126_,
		_w9127_
	);
	LUT2 #(
		.INIT('h4)
	) name8596 (
		\sa23_reg[5]/P0001 ,
		_w8552_,
		_w9128_
	);
	LUT2 #(
		.INIT('h8)
	) name8597 (
		_w8525_,
		_w8537_,
		_w9129_
	);
	LUT2 #(
		.INIT('h4)
	) name8598 (
		\sa23_reg[7]/NET0131 ,
		_w9129_,
		_w9130_
	);
	LUT2 #(
		.INIT('h1)
	) name8599 (
		_w9128_,
		_w9130_,
		_w9131_
	);
	LUT2 #(
		.INIT('h4)
	) name8600 (
		_w9127_,
		_w9131_,
		_w9132_
	);
	LUT2 #(
		.INIT('h2)
	) name8601 (
		\sa23_reg[2]/P0001 ,
		_w9132_,
		_w9133_
	);
	LUT2 #(
		.INIT('h8)
	) name8602 (
		\sa23_reg[3]/P0001 ,
		_w8571_,
		_w9134_
	);
	LUT2 #(
		.INIT('h4)
	) name8603 (
		\sa23_reg[2]/P0001 ,
		_w8609_,
		_w9135_
	);
	LUT2 #(
		.INIT('h8)
	) name8604 (
		\sa23_reg[1]/P0001 ,
		_w9135_,
		_w9136_
	);
	LUT2 #(
		.INIT('h8)
	) name8605 (
		_w8523_,
		_w8547_,
		_w9137_
	);
	LUT2 #(
		.INIT('h8)
	) name8606 (
		_w8511_,
		_w8522_,
		_w9138_
	);
	LUT2 #(
		.INIT('h8)
	) name8607 (
		_w8519_,
		_w8529_,
		_w9139_
	);
	LUT2 #(
		.INIT('h4)
	) name8608 (
		\sa23_reg[2]/P0001 ,
		_w9066_,
		_w9140_
	);
	LUT2 #(
		.INIT('h8)
	) name8609 (
		_w8618_,
		_w8660_,
		_w9141_
	);
	LUT2 #(
		.INIT('h1)
	) name8610 (
		_w9085_,
		_w9138_,
		_w9142_
	);
	LUT2 #(
		.INIT('h4)
	) name8611 (
		_w9139_,
		_w9142_,
		_w9143_
	);
	LUT2 #(
		.INIT('h1)
	) name8612 (
		_w9107_,
		_w9140_,
		_w9144_
	);
	LUT2 #(
		.INIT('h4)
	) name8613 (
		_w9141_,
		_w9144_,
		_w9145_
	);
	LUT2 #(
		.INIT('h8)
	) name8614 (
		_w9143_,
		_w9145_,
		_w9146_
	);
	LUT2 #(
		.INIT('h1)
	) name8615 (
		\sa23_reg[0]/P0001 ,
		_w9146_,
		_w9147_
	);
	LUT2 #(
		.INIT('h2)
	) name8616 (
		\sa23_reg[2]/P0001 ,
		_w8557_,
		_w9148_
	);
	LUT2 #(
		.INIT('h8)
	) name8617 (
		_w8577_,
		_w8624_,
		_w9149_
	);
	LUT2 #(
		.INIT('h2)
	) name8618 (
		_w9148_,
		_w9149_,
		_w9150_
	);
	LUT2 #(
		.INIT('h8)
	) name8619 (
		\sa23_reg[4]/P0001 ,
		_w8525_,
		_w9151_
	);
	LUT2 #(
		.INIT('h4)
	) name8620 (
		\sa23_reg[7]/NET0131 ,
		_w9151_,
		_w9152_
	);
	LUT2 #(
		.INIT('h1)
	) name8621 (
		\sa23_reg[2]/P0001 ,
		_w9152_,
		_w9153_
	);
	LUT2 #(
		.INIT('h4)
	) name8622 (
		\sa23_reg[6]/NET0131 ,
		_w8532_,
		_w9154_
	);
	LUT2 #(
		.INIT('h1)
	) name8623 (
		_w8570_,
		_w9154_,
		_w9155_
	);
	LUT2 #(
		.INIT('h8)
	) name8624 (
		_w9153_,
		_w9155_,
		_w9156_
	);
	LUT2 #(
		.INIT('h1)
	) name8625 (
		_w9150_,
		_w9156_,
		_w9157_
	);
	LUT2 #(
		.INIT('h8)
	) name8626 (
		_w8521_,
		_w8522_,
		_w9158_
	);
	LUT2 #(
		.INIT('h8)
	) name8627 (
		_w8569_,
		_w8624_,
		_w9159_
	);
	LUT2 #(
		.INIT('h1)
	) name8628 (
		_w9158_,
		_w9159_,
		_w9160_
	);
	LUT2 #(
		.INIT('h4)
	) name8629 (
		_w9157_,
		_w9160_,
		_w9161_
	);
	LUT2 #(
		.INIT('h4)
	) name8630 (
		_w9147_,
		_w9161_,
		_w9162_
	);
	LUT2 #(
		.INIT('h1)
	) name8631 (
		\sa23_reg[1]/P0001 ,
		_w9162_,
		_w9163_
	);
	LUT2 #(
		.INIT('h1)
	) name8632 (
		_w9134_,
		_w9137_,
		_w9164_
	);
	LUT2 #(
		.INIT('h4)
	) name8633 (
		_w9136_,
		_w9164_,
		_w9165_
	);
	LUT2 #(
		.INIT('h4)
	) name8634 (
		_w9133_,
		_w9165_,
		_w9166_
	);
	LUT2 #(
		.INIT('h4)
	) name8635 (
		_w9122_,
		_w9166_,
		_w9167_
	);
	LUT2 #(
		.INIT('h4)
	) name8636 (
		_w9163_,
		_w9167_,
		_w9168_
	);
	LUT2 #(
		.INIT('h4)
	) name8637 (
		_w9095_,
		_w9168_,
		_w9169_
	);
	LUT2 #(
		.INIT('h2)
	) name8638 (
		_w9063_,
		_w9169_,
		_w9170_
	);
	LUT2 #(
		.INIT('h4)
	) name8639 (
		_w9063_,
		_w9169_,
		_w9171_
	);
	LUT2 #(
		.INIT('h1)
	) name8640 (
		_w9170_,
		_w9171_,
		_w9172_
	);
	LUT2 #(
		.INIT('h8)
	) name8641 (
		\sa01_reg[3]/P0001 ,
		_w8245_,
		_w9173_
	);
	LUT2 #(
		.INIT('h8)
	) name8642 (
		\sa01_reg[4]/P0001 ,
		_w9173_,
		_w9174_
	);
	LUT2 #(
		.INIT('h8)
	) name8643 (
		\sa01_reg[4]/P0001 ,
		_w8276_,
		_w9175_
	);
	LUT2 #(
		.INIT('h8)
	) name8644 (
		\sa01_reg[5]/P0001 ,
		_w9175_,
		_w9176_
	);
	LUT2 #(
		.INIT('h1)
	) name8645 (
		_w9173_,
		_w9176_,
		_w9177_
	);
	LUT2 #(
		.INIT('h2)
	) name8646 (
		\sa01_reg[2]/P0001 ,
		_w9177_,
		_w9178_
	);
	LUT2 #(
		.INIT('h8)
	) name8647 (
		_w8253_,
		_w8368_,
		_w9179_
	);
	LUT2 #(
		.INIT('h8)
	) name8648 (
		_w8221_,
		_w8308_,
		_w9180_
	);
	LUT2 #(
		.INIT('h8)
	) name8649 (
		_w8267_,
		_w8277_,
		_w9181_
	);
	LUT2 #(
		.INIT('h4)
	) name8650 (
		\sa01_reg[7]/NET0131 ,
		_w8304_,
		_w9182_
	);
	LUT2 #(
		.INIT('h8)
	) name8651 (
		\sa01_reg[3]/P0001 ,
		_w8221_,
		_w9183_
	);
	LUT2 #(
		.INIT('h4)
	) name8652 (
		\sa01_reg[3]/P0001 ,
		_w8242_,
		_w9184_
	);
	LUT2 #(
		.INIT('h8)
	) name8653 (
		\sa01_reg[4]/P0001 ,
		_w9184_,
		_w9185_
	);
	LUT2 #(
		.INIT('h1)
	) name8654 (
		_w9182_,
		_w9183_,
		_w9186_
	);
	LUT2 #(
		.INIT('h4)
	) name8655 (
		_w9185_,
		_w9186_,
		_w9187_
	);
	LUT2 #(
		.INIT('h1)
	) name8656 (
		\sa01_reg[2]/P0001 ,
		_w9187_,
		_w9188_
	);
	LUT2 #(
		.INIT('h1)
	) name8657 (
		_w8352_,
		_w9179_,
		_w9189_
	);
	LUT2 #(
		.INIT('h4)
	) name8658 (
		_w9180_,
		_w9189_,
		_w9190_
	);
	LUT2 #(
		.INIT('h1)
	) name8659 (
		_w9174_,
		_w9181_,
		_w9191_
	);
	LUT2 #(
		.INIT('h8)
	) name8660 (
		_w9190_,
		_w9191_,
		_w9192_
	);
	LUT2 #(
		.INIT('h4)
	) name8661 (
		_w9178_,
		_w9192_,
		_w9193_
	);
	LUT2 #(
		.INIT('h4)
	) name8662 (
		_w9188_,
		_w9193_,
		_w9194_
	);
	LUT2 #(
		.INIT('h2)
	) name8663 (
		\sa01_reg[1]/P0001 ,
		_w9194_,
		_w9195_
	);
	LUT2 #(
		.INIT('h8)
	) name8664 (
		_w8214_,
		_w8221_,
		_w9196_
	);
	LUT2 #(
		.INIT('h2)
	) name8665 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		_w9197_
	);
	LUT2 #(
		.INIT('h8)
	) name8666 (
		_w8215_,
		_w9197_,
		_w9198_
	);
	LUT2 #(
		.INIT('h1)
	) name8667 (
		_w9196_,
		_w9198_,
		_w9199_
	);
	LUT2 #(
		.INIT('h1)
	) name8668 (
		\sa01_reg[5]/P0001 ,
		_w9199_,
		_w9200_
	);
	LUT2 #(
		.INIT('h4)
	) name8669 (
		\sa01_reg[4]/P0001 ,
		_w8227_,
		_w9201_
	);
	LUT2 #(
		.INIT('h8)
	) name8670 (
		_w8329_,
		_w9201_,
		_w9202_
	);
	LUT2 #(
		.INIT('h1)
	) name8671 (
		_w8322_,
		_w9202_,
		_w9203_
	);
	LUT2 #(
		.INIT('h4)
	) name8672 (
		_w9200_,
		_w9203_,
		_w9204_
	);
	LUT2 #(
		.INIT('h1)
	) name8673 (
		\sa01_reg[1]/P0001 ,
		_w9204_,
		_w9205_
	);
	LUT2 #(
		.INIT('h4)
	) name8674 (
		\sa01_reg[5]/P0001 ,
		_w8276_,
		_w9206_
	);
	LUT2 #(
		.INIT('h8)
	) name8675 (
		_w8287_,
		_w9206_,
		_w9207_
	);
	LUT2 #(
		.INIT('h8)
	) name8676 (
		_w8215_,
		_w8222_,
		_w9208_
	);
	LUT2 #(
		.INIT('h4)
	) name8677 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w9209_
	);
	LUT2 #(
		.INIT('h8)
	) name8678 (
		_w8279_,
		_w9209_,
		_w9210_
	);
	LUT2 #(
		.INIT('h8)
	) name8679 (
		_w8238_,
		_w8368_,
		_w9211_
	);
	LUT2 #(
		.INIT('h8)
	) name8680 (
		_w8225_,
		_w8254_,
		_w9212_
	);
	LUT2 #(
		.INIT('h1)
	) name8681 (
		_w9211_,
		_w9212_,
		_w9213_
	);
	LUT2 #(
		.INIT('h1)
	) name8682 (
		\sa01_reg[2]/P0001 ,
		_w9213_,
		_w9214_
	);
	LUT2 #(
		.INIT('h8)
	) name8683 (
		\sa01_reg[4]/P0001 ,
		_w8245_,
		_w9215_
	);
	LUT2 #(
		.INIT('h4)
	) name8684 (
		\sa01_reg[4]/P0001 ,
		_w8368_,
		_w9216_
	);
	LUT2 #(
		.INIT('h1)
	) name8685 (
		_w9215_,
		_w9216_,
		_w9217_
	);
	LUT2 #(
		.INIT('h2)
	) name8686 (
		_w8329_,
		_w9217_,
		_w9218_
	);
	LUT2 #(
		.INIT('h8)
	) name8687 (
		_w8227_,
		_w8265_,
		_w9219_
	);
	LUT2 #(
		.INIT('h1)
	) name8688 (
		_w9208_,
		_w9219_,
		_w9220_
	);
	LUT2 #(
		.INIT('h4)
	) name8689 (
		_w9207_,
		_w9220_,
		_w9221_
	);
	LUT2 #(
		.INIT('h4)
	) name8690 (
		_w9210_,
		_w9221_,
		_w9222_
	);
	LUT2 #(
		.INIT('h1)
	) name8691 (
		_w9214_,
		_w9218_,
		_w9223_
	);
	LUT2 #(
		.INIT('h8)
	) name8692 (
		_w9222_,
		_w9223_,
		_w9224_
	);
	LUT2 #(
		.INIT('h4)
	) name8693 (
		_w9205_,
		_w9224_,
		_w9225_
	);
	LUT2 #(
		.INIT('h4)
	) name8694 (
		_w9195_,
		_w9225_,
		_w9226_
	);
	LUT2 #(
		.INIT('h1)
	) name8695 (
		\sa01_reg[0]/P0001 ,
		_w9226_,
		_w9227_
	);
	LUT2 #(
		.INIT('h4)
	) name8696 (
		\sa01_reg[5]/P0001 ,
		_w8226_,
		_w9228_
	);
	LUT2 #(
		.INIT('h1)
	) name8697 (
		_w8354_,
		_w9228_,
		_w9229_
	);
	LUT2 #(
		.INIT('h2)
	) name8698 (
		\sa01_reg[1]/P0001 ,
		_w9229_,
		_w9230_
	);
	LUT2 #(
		.INIT('h4)
	) name8699 (
		\sa01_reg[4]/P0001 ,
		_w8342_,
		_w9231_
	);
	LUT2 #(
		.INIT('h1)
	) name8700 (
		_w8266_,
		_w8343_,
		_w9232_
	);
	LUT2 #(
		.INIT('h4)
	) name8701 (
		_w9231_,
		_w9232_,
		_w9233_
	);
	LUT2 #(
		.INIT('h4)
	) name8702 (
		_w9230_,
		_w9233_,
		_w9234_
	);
	LUT2 #(
		.INIT('h1)
	) name8703 (
		\sa01_reg[2]/P0001 ,
		_w9234_,
		_w9235_
	);
	LUT2 #(
		.INIT('h4)
	) name8704 (
		\sa01_reg[6]/NET0131 ,
		_w8360_,
		_w9236_
	);
	LUT2 #(
		.INIT('h8)
	) name8705 (
		_w8214_,
		_w8279_,
		_w9237_
	);
	LUT2 #(
		.INIT('h8)
	) name8706 (
		\sa01_reg[7]/NET0131 ,
		_w8256_,
		_w9238_
	);
	LUT2 #(
		.INIT('h1)
	) name8707 (
		_w8217_,
		_w9236_,
		_w9239_
	);
	LUT2 #(
		.INIT('h1)
	) name8708 (
		_w9237_,
		_w9238_,
		_w9240_
	);
	LUT2 #(
		.INIT('h8)
	) name8709 (
		_w9239_,
		_w9240_,
		_w9241_
	);
	LUT2 #(
		.INIT('h2)
	) name8710 (
		\sa01_reg[1]/P0001 ,
		_w9241_,
		_w9242_
	);
	LUT2 #(
		.INIT('h8)
	) name8711 (
		_w8214_,
		_w8258_,
		_w9243_
	);
	LUT2 #(
		.INIT('h1)
	) name8712 (
		\sa01_reg[2]/P0001 ,
		_w8277_,
		_w9244_
	);
	LUT2 #(
		.INIT('h4)
	) name8713 (
		_w8255_,
		_w9244_,
		_w9245_
	);
	LUT2 #(
		.INIT('h4)
	) name8714 (
		\sa01_reg[5]/P0001 ,
		_w8225_,
		_w9246_
	);
	LUT2 #(
		.INIT('h2)
	) name8715 (
		\sa01_reg[2]/P0001 ,
		_w8305_,
		_w9247_
	);
	LUT2 #(
		.INIT('h4)
	) name8716 (
		_w9246_,
		_w9247_,
		_w9248_
	);
	LUT2 #(
		.INIT('h1)
	) name8717 (
		_w9245_,
		_w9248_,
		_w9249_
	);
	LUT2 #(
		.INIT('h1)
	) name8718 (
		_w8343_,
		_w9243_,
		_w9250_
	);
	LUT2 #(
		.INIT('h4)
	) name8719 (
		_w9249_,
		_w9250_,
		_w9251_
	);
	LUT2 #(
		.INIT('h1)
	) name8720 (
		\sa01_reg[1]/P0001 ,
		_w9251_,
		_w9252_
	);
	LUT2 #(
		.INIT('h8)
	) name8721 (
		_w8304_,
		_w8368_,
		_w9253_
	);
	LUT2 #(
		.INIT('h1)
	) name8722 (
		_w9243_,
		_w9253_,
		_w9254_
	);
	LUT2 #(
		.INIT('h2)
	) name8723 (
		\sa01_reg[2]/P0001 ,
		_w9254_,
		_w9255_
	);
	LUT2 #(
		.INIT('h8)
	) name8724 (
		_w8276_,
		_w8354_,
		_w9256_
	);
	LUT2 #(
		.INIT('h1)
	) name8725 (
		_w8312_,
		_w9256_,
		_w9257_
	);
	LUT2 #(
		.INIT('h4)
	) name8726 (
		_w9255_,
		_w9257_,
		_w9258_
	);
	LUT2 #(
		.INIT('h4)
	) name8727 (
		_w9242_,
		_w9258_,
		_w9259_
	);
	LUT2 #(
		.INIT('h4)
	) name8728 (
		_w9235_,
		_w9259_,
		_w9260_
	);
	LUT2 #(
		.INIT('h4)
	) name8729 (
		_w9252_,
		_w9260_,
		_w9261_
	);
	LUT2 #(
		.INIT('h2)
	) name8730 (
		\sa01_reg[0]/P0001 ,
		_w9261_,
		_w9262_
	);
	LUT2 #(
		.INIT('h1)
	) name8731 (
		_w8344_,
		_w9206_,
		_w9263_
	);
	LUT2 #(
		.INIT('h4)
	) name8732 (
		_w8258_,
		_w9263_,
		_w9264_
	);
	LUT2 #(
		.INIT('h2)
	) name8733 (
		_w8287_,
		_w9264_,
		_w9265_
	);
	LUT2 #(
		.INIT('h8)
	) name8734 (
		\sa01_reg[5]/P0001 ,
		_w8253_,
		_w9266_
	);
	LUT2 #(
		.INIT('h8)
	) name8735 (
		_w8327_,
		_w9266_,
		_w9267_
	);
	LUT2 #(
		.INIT('h8)
	) name8736 (
		\sa01_reg[6]/NET0131 ,
		_w8331_,
		_w9268_
	);
	LUT2 #(
		.INIT('h1)
	) name8737 (
		_w8321_,
		_w8361_,
		_w9269_
	);
	LUT2 #(
		.INIT('h4)
	) name8738 (
		_w9268_,
		_w9269_,
		_w9270_
	);
	LUT2 #(
		.INIT('h1)
	) name8739 (
		\sa01_reg[2]/P0001 ,
		_w9270_,
		_w9271_
	);
	LUT2 #(
		.INIT('h1)
	) name8740 (
		_w8362_,
		_w9267_,
		_w9272_
	);
	LUT2 #(
		.INIT('h4)
	) name8741 (
		_w9265_,
		_w9272_,
		_w9273_
	);
	LUT2 #(
		.INIT('h4)
	) name8742 (
		_w9271_,
		_w9273_,
		_w9274_
	);
	LUT2 #(
		.INIT('h1)
	) name8743 (
		\sa01_reg[1]/P0001 ,
		_w9274_,
		_w9275_
	);
	LUT2 #(
		.INIT('h8)
	) name8744 (
		\sa01_reg[4]/P0001 ,
		_w8219_,
		_w9276_
	);
	LUT2 #(
		.INIT('h8)
	) name8745 (
		_w8329_,
		_w9276_,
		_w9277_
	);
	LUT2 #(
		.INIT('h1)
	) name8746 (
		_w8220_,
		_w8352_,
		_w9278_
	);
	LUT2 #(
		.INIT('h1)
	) name8747 (
		\sa01_reg[2]/P0001 ,
		_w9278_,
		_w9279_
	);
	LUT2 #(
		.INIT('h8)
	) name8748 (
		_w8277_,
		_w8287_,
		_w9280_
	);
	LUT2 #(
		.INIT('h8)
	) name8749 (
		_w8253_,
		_w9216_,
		_w9281_
	);
	LUT2 #(
		.INIT('h1)
	) name8750 (
		_w9210_,
		_w9280_,
		_w9282_
	);
	LUT2 #(
		.INIT('h4)
	) name8751 (
		_w9281_,
		_w9282_,
		_w9283_
	);
	LUT2 #(
		.INIT('h2)
	) name8752 (
		\sa01_reg[1]/P0001 ,
		_w9283_,
		_w9284_
	);
	LUT2 #(
		.INIT('h1)
	) name8753 (
		_w9277_,
		_w9279_,
		_w9285_
	);
	LUT2 #(
		.INIT('h4)
	) name8754 (
		_w9284_,
		_w9285_,
		_w9286_
	);
	LUT2 #(
		.INIT('h4)
	) name8755 (
		_w9275_,
		_w9286_,
		_w9287_
	);
	LUT2 #(
		.INIT('h4)
	) name8756 (
		_w9227_,
		_w9287_,
		_w9288_
	);
	LUT2 #(
		.INIT('h4)
	) name8757 (
		_w9262_,
		_w9288_,
		_w9289_
	);
	LUT2 #(
		.INIT('h2)
	) name8758 (
		_w8507_,
		_w9289_,
		_w9290_
	);
	LUT2 #(
		.INIT('h4)
	) name8759 (
		_w8507_,
		_w9289_,
		_w9291_
	);
	LUT2 #(
		.INIT('h1)
	) name8760 (
		_w9290_,
		_w9291_,
		_w9292_
	);
	LUT2 #(
		.INIT('h8)
	) name8761 (
		_w9172_,
		_w9292_,
		_w9293_
	);
	LUT2 #(
		.INIT('h1)
	) name8762 (
		_w9172_,
		_w9292_,
		_w9294_
	);
	LUT2 #(
		.INIT('h1)
	) name8763 (
		_w9293_,
		_w9294_,
		_w9295_
	);
	LUT2 #(
		.INIT('h4)
	) name8764 (
		_w8977_,
		_w9295_,
		_w9296_
	);
	LUT2 #(
		.INIT('h2)
	) name8765 (
		_w8977_,
		_w9295_,
		_w9297_
	);
	LUT2 #(
		.INIT('h1)
	) name8766 (
		\ld_r_reg/P0001 ,
		_w9296_,
		_w9298_
	);
	LUT2 #(
		.INIT('h4)
	) name8767 (
		_w9297_,
		_w9298_,
		_w9299_
	);
	LUT2 #(
		.INIT('h2)
	) name8768 (
		\text_in_r_reg[94]/P0001 ,
		\u0_w_reg[1][30]/P0001 ,
		_w9300_
	);
	LUT2 #(
		.INIT('h4)
	) name8769 (
		\text_in_r_reg[94]/P0001 ,
		\u0_w_reg[1][30]/P0001 ,
		_w9301_
	);
	LUT2 #(
		.INIT('h2)
	) name8770 (
		\ld_r_reg/P0001 ,
		_w9300_,
		_w9302_
	);
	LUT2 #(
		.INIT('h4)
	) name8771 (
		_w9301_,
		_w9302_,
		_w9303_
	);
	LUT2 #(
		.INIT('h1)
	) name8772 (
		_w9299_,
		_w9303_,
		_w9304_
	);
	LUT2 #(
		.INIT('h8)
	) name8773 (
		_w8240_,
		_w9184_,
		_w9305_
	);
	LUT2 #(
		.INIT('h1)
	) name8774 (
		_w8243_,
		_w9305_,
		_w9306_
	);
	LUT2 #(
		.INIT('h4)
	) name8775 (
		_w9214_,
		_w9306_,
		_w9307_
	);
	LUT2 #(
		.INIT('h1)
	) name8776 (
		\sa01_reg[1]/P0001 ,
		_w9307_,
		_w9308_
	);
	LUT2 #(
		.INIT('h8)
	) name8777 (
		_w8276_,
		_w8308_,
		_w9309_
	);
	LUT2 #(
		.INIT('h2)
	) name8778 (
		\sa01_reg[1]/P0001 ,
		_w8225_,
		_w9310_
	);
	LUT2 #(
		.INIT('h8)
	) name8779 (
		_w8351_,
		_w9310_,
		_w9311_
	);
	LUT2 #(
		.INIT('h1)
	) name8780 (
		_w9185_,
		_w9309_,
		_w9312_
	);
	LUT2 #(
		.INIT('h4)
	) name8781 (
		_w9311_,
		_w9312_,
		_w9313_
	);
	LUT2 #(
		.INIT('h1)
	) name8782 (
		\sa01_reg[2]/P0001 ,
		_w9313_,
		_w9314_
	);
	LUT2 #(
		.INIT('h8)
	) name8783 (
		_w8218_,
		_w8245_,
		_w9315_
	);
	LUT2 #(
		.INIT('h1)
	) name8784 (
		_w9236_,
		_w9315_,
		_w9316_
	);
	LUT2 #(
		.INIT('h2)
	) name8785 (
		\sa01_reg[1]/P0001 ,
		_w9316_,
		_w9317_
	);
	LUT2 #(
		.INIT('h4)
	) name8786 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[2]/P0001 ,
		_w9318_
	);
	LUT2 #(
		.INIT('h8)
	) name8787 (
		\sa01_reg[3]/P0001 ,
		_w8224_,
		_w9319_
	);
	LUT2 #(
		.INIT('h1)
	) name8788 (
		_w9206_,
		_w9319_,
		_w9320_
	);
	LUT2 #(
		.INIT('h2)
	) name8789 (
		_w9318_,
		_w9320_,
		_w9321_
	);
	LUT2 #(
		.INIT('h8)
	) name8790 (
		_w8329_,
		_w8344_,
		_w9322_
	);
	LUT2 #(
		.INIT('h1)
	) name8791 (
		_w8286_,
		_w9243_,
		_w9323_
	);
	LUT2 #(
		.INIT('h8)
	) name8792 (
		_w8254_,
		_w8304_,
		_w9324_
	);
	LUT2 #(
		.INIT('h1)
	) name8793 (
		_w9175_,
		_w9180_,
		_w9325_
	);
	LUT2 #(
		.INIT('h4)
	) name8794 (
		_w9324_,
		_w9325_,
		_w9326_
	);
	LUT2 #(
		.INIT('h2)
	) name8795 (
		\sa01_reg[1]/P0001 ,
		_w9326_,
		_w9327_
	);
	LUT2 #(
		.INIT('h4)
	) name8796 (
		_w9219_,
		_w9323_,
		_w9328_
	);
	LUT2 #(
		.INIT('h4)
	) name8797 (
		_w9327_,
		_w9328_,
		_w9329_
	);
	LUT2 #(
		.INIT('h2)
	) name8798 (
		\sa01_reg[2]/P0001 ,
		_w9329_,
		_w9330_
	);
	LUT2 #(
		.INIT('h1)
	) name8799 (
		_w9321_,
		_w9322_,
		_w9331_
	);
	LUT2 #(
		.INIT('h4)
	) name8800 (
		_w9317_,
		_w9331_,
		_w9332_
	);
	LUT2 #(
		.INIT('h4)
	) name8801 (
		_w9308_,
		_w9332_,
		_w9333_
	);
	LUT2 #(
		.INIT('h4)
	) name8802 (
		_w9314_,
		_w9333_,
		_w9334_
	);
	LUT2 #(
		.INIT('h4)
	) name8803 (
		_w9330_,
		_w9334_,
		_w9335_
	);
	LUT2 #(
		.INIT('h2)
	) name8804 (
		\sa01_reg[0]/P0001 ,
		_w9335_,
		_w9336_
	);
	LUT2 #(
		.INIT('h8)
	) name8805 (
		_w8221_,
		_w8267_,
		_w9337_
	);
	LUT2 #(
		.INIT('h8)
	) name8806 (
		\sa01_reg[7]/NET0131 ,
		_w8356_,
		_w9338_
	);
	LUT2 #(
		.INIT('h1)
	) name8807 (
		_w8282_,
		_w8311_,
		_w9339_
	);
	LUT2 #(
		.INIT('h2)
	) name8808 (
		\sa01_reg[3]/P0001 ,
		_w9339_,
		_w9340_
	);
	LUT2 #(
		.INIT('h1)
	) name8809 (
		\sa01_reg[1]/P0001 ,
		_w9309_,
		_w9341_
	);
	LUT2 #(
		.INIT('h4)
	) name8810 (
		_w9337_,
		_w9341_,
		_w9342_
	);
	LUT2 #(
		.INIT('h1)
	) name8811 (
		_w8330_,
		_w9338_,
		_w9343_
	);
	LUT2 #(
		.INIT('h8)
	) name8812 (
		_w9342_,
		_w9343_,
		_w9344_
	);
	LUT2 #(
		.INIT('h4)
	) name8813 (
		_w9340_,
		_w9344_,
		_w9345_
	);
	LUT2 #(
		.INIT('h2)
	) name8814 (
		_w9197_,
		_w9217_,
		_w9346_
	);
	LUT2 #(
		.INIT('h4)
	) name8815 (
		\sa01_reg[2]/P0001 ,
		_w9219_,
		_w9347_
	);
	LUT2 #(
		.INIT('h2)
	) name8816 (
		\sa01_reg[1]/P0001 ,
		_w8361_,
		_w9348_
	);
	LUT2 #(
		.INIT('h4)
	) name8817 (
		_w9347_,
		_w9348_,
		_w9349_
	);
	LUT2 #(
		.INIT('h4)
	) name8818 (
		_w9346_,
		_w9349_,
		_w9350_
	);
	LUT2 #(
		.INIT('h1)
	) name8819 (
		_w9345_,
		_w9350_,
		_w9351_
	);
	LUT2 #(
		.INIT('h8)
	) name8820 (
		\sa01_reg[4]/P0001 ,
		_w8227_,
		_w9352_
	);
	LUT2 #(
		.INIT('h4)
	) name8821 (
		\sa01_reg[3]/P0001 ,
		_w9352_,
		_w9353_
	);
	LUT2 #(
		.INIT('h2)
	) name8822 (
		\sa01_reg[4]/P0001 ,
		_w8235_,
		_w9354_
	);
	LUT2 #(
		.INIT('h2)
	) name8823 (
		_w8319_,
		_w9354_,
		_w9355_
	);
	LUT2 #(
		.INIT('h8)
	) name8824 (
		_w8214_,
		_w8342_,
		_w9356_
	);
	LUT2 #(
		.INIT('h8)
	) name8825 (
		\sa01_reg[6]/NET0131 ,
		_w9356_,
		_w9357_
	);
	LUT2 #(
		.INIT('h1)
	) name8826 (
		\sa01_reg[2]/P0001 ,
		_w9353_,
		_w9358_
	);
	LUT2 #(
		.INIT('h1)
	) name8827 (
		_w9355_,
		_w9357_,
		_w9359_
	);
	LUT2 #(
		.INIT('h8)
	) name8828 (
		_w9358_,
		_w9359_,
		_w9360_
	);
	LUT2 #(
		.INIT('h4)
	) name8829 (
		\sa01_reg[3]/P0001 ,
		_w9201_,
		_w9361_
	);
	LUT2 #(
		.INIT('h2)
	) name8830 (
		\sa01_reg[2]/P0001 ,
		_w9338_,
		_w9362_
	);
	LUT2 #(
		.INIT('h4)
	) name8831 (
		_w9361_,
		_w9362_,
		_w9363_
	);
	LUT2 #(
		.INIT('h1)
	) name8832 (
		_w9360_,
		_w9363_,
		_w9364_
	);
	LUT2 #(
		.INIT('h1)
	) name8833 (
		_w9351_,
		_w9364_,
		_w9365_
	);
	LUT2 #(
		.INIT('h1)
	) name8834 (
		\sa01_reg[0]/P0001 ,
		_w9365_,
		_w9366_
	);
	LUT2 #(
		.INIT('h8)
	) name8835 (
		\sa01_reg[3]/P0001 ,
		_w9208_,
		_w9367_
	);
	LUT2 #(
		.INIT('h4)
	) name8836 (
		\sa01_reg[5]/P0001 ,
		_w9175_,
		_w9368_
	);
	LUT2 #(
		.INIT('h4)
	) name8837 (
		\sa01_reg[6]/NET0131 ,
		_w9173_,
		_w9369_
	);
	LUT2 #(
		.INIT('h1)
	) name8838 (
		_w8243_,
		_w9368_,
		_w9370_
	);
	LUT2 #(
		.INIT('h4)
	) name8839 (
		_w9369_,
		_w9370_,
		_w9371_
	);
	LUT2 #(
		.INIT('h1)
	) name8840 (
		\sa01_reg[2]/P0001 ,
		_w9371_,
		_w9372_
	);
	LUT2 #(
		.INIT('h8)
	) name8841 (
		_w8235_,
		_w8308_,
		_w9373_
	);
	LUT2 #(
		.INIT('h8)
	) name8842 (
		\sa01_reg[2]/P0001 ,
		_w9373_,
		_w9374_
	);
	LUT2 #(
		.INIT('h8)
	) name8843 (
		_w8224_,
		_w8253_,
		_w9375_
	);
	LUT2 #(
		.INIT('h8)
	) name8844 (
		_w8257_,
		_w8267_,
		_w9376_
	);
	LUT2 #(
		.INIT('h1)
	) name8845 (
		_w9375_,
		_w9376_,
		_w9377_
	);
	LUT2 #(
		.INIT('h4)
	) name8846 (
		_w9367_,
		_w9377_,
		_w9378_
	);
	LUT2 #(
		.INIT('h4)
	) name8847 (
		_w9374_,
		_w9378_,
		_w9379_
	);
	LUT2 #(
		.INIT('h4)
	) name8848 (
		_w9372_,
		_w9379_,
		_w9380_
	);
	LUT2 #(
		.INIT('h1)
	) name8849 (
		\sa01_reg[1]/P0001 ,
		_w9380_,
		_w9381_
	);
	LUT2 #(
		.INIT('h2)
	) name8850 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[2]/P0001 ,
		_w9382_
	);
	LUT2 #(
		.INIT('h8)
	) name8851 (
		_w8220_,
		_w9382_,
		_w9383_
	);
	LUT2 #(
		.INIT('h1)
	) name8852 (
		_w8286_,
		_w8339_,
		_w9384_
	);
	LUT2 #(
		.INIT('h2)
	) name8853 (
		_w8303_,
		_w9384_,
		_w9385_
	);
	LUT2 #(
		.INIT('h4)
	) name8854 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		_w9386_
	);
	LUT2 #(
		.INIT('h8)
	) name8855 (
		_w8243_,
		_w9386_,
		_w9387_
	);
	LUT2 #(
		.INIT('h8)
	) name8856 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[2]/P0001 ,
		_w9388_
	);
	LUT2 #(
		.INIT('h8)
	) name8857 (
		\sa01_reg[4]/P0001 ,
		_w8216_,
		_w9389_
	);
	LUT2 #(
		.INIT('h4)
	) name8858 (
		\sa01_reg[4]/P0001 ,
		_w9369_,
		_w9390_
	);
	LUT2 #(
		.INIT('h1)
	) name8859 (
		_w8362_,
		_w9389_,
		_w9391_
	);
	LUT2 #(
		.INIT('h4)
	) name8860 (
		_w9390_,
		_w9391_,
		_w9392_
	);
	LUT2 #(
		.INIT('h2)
	) name8861 (
		_w9388_,
		_w9392_,
		_w9393_
	);
	LUT2 #(
		.INIT('h1)
	) name8862 (
		_w8268_,
		_w9387_,
		_w9394_
	);
	LUT2 #(
		.INIT('h4)
	) name8863 (
		_w9383_,
		_w9394_,
		_w9395_
	);
	LUT2 #(
		.INIT('h4)
	) name8864 (
		_w9385_,
		_w9395_,
		_w9396_
	);
	LUT2 #(
		.INIT('h4)
	) name8865 (
		_w9393_,
		_w9396_,
		_w9397_
	);
	LUT2 #(
		.INIT('h4)
	) name8866 (
		_w9381_,
		_w9397_,
		_w9398_
	);
	LUT2 #(
		.INIT('h4)
	) name8867 (
		_w9366_,
		_w9398_,
		_w9399_
	);
	LUT2 #(
		.INIT('h4)
	) name8868 (
		_w9336_,
		_w9399_,
		_w9400_
	);
	LUT2 #(
		.INIT('h1)
	) name8869 (
		_w8681_,
		_w9400_,
		_w9401_
	);
	LUT2 #(
		.INIT('h8)
	) name8870 (
		_w8681_,
		_w9400_,
		_w9402_
	);
	LUT2 #(
		.INIT('h1)
	) name8871 (
		_w9401_,
		_w9402_,
		_w9403_
	);
	LUT2 #(
		.INIT('h2)
	) name8872 (
		\u0_w_reg[1][22]/P0001 ,
		_w8974_,
		_w9404_
	);
	LUT2 #(
		.INIT('h4)
	) name8873 (
		\u0_w_reg[1][22]/P0001 ,
		_w8974_,
		_w9405_
	);
	LUT2 #(
		.INIT('h1)
	) name8874 (
		_w9404_,
		_w9405_,
		_w9406_
	);
	LUT2 #(
		.INIT('h8)
	) name8875 (
		_w9169_,
		_w9406_,
		_w9407_
	);
	LUT2 #(
		.INIT('h1)
	) name8876 (
		_w9169_,
		_w9406_,
		_w9408_
	);
	LUT2 #(
		.INIT('h1)
	) name8877 (
		_w9407_,
		_w9408_,
		_w9409_
	);
	LUT2 #(
		.INIT('h1)
	) name8878 (
		_w9403_,
		_w9409_,
		_w9410_
	);
	LUT2 #(
		.INIT('h8)
	) name8879 (
		_w9403_,
		_w9409_,
		_w9411_
	);
	LUT2 #(
		.INIT('h1)
	) name8880 (
		\ld_r_reg/P0001 ,
		_w9410_,
		_w9412_
	);
	LUT2 #(
		.INIT('h4)
	) name8881 (
		_w9411_,
		_w9412_,
		_w9413_
	);
	LUT2 #(
		.INIT('h2)
	) name8882 (
		\text_in_r_reg[86]/P0001 ,
		\u0_w_reg[1][22]/P0001 ,
		_w9414_
	);
	LUT2 #(
		.INIT('h4)
	) name8883 (
		\text_in_r_reg[86]/P0001 ,
		\u0_w_reg[1][22]/P0001 ,
		_w9415_
	);
	LUT2 #(
		.INIT('h2)
	) name8884 (
		\ld_r_reg/P0001 ,
		_w9414_,
		_w9416_
	);
	LUT2 #(
		.INIT('h4)
	) name8885 (
		_w9415_,
		_w9416_,
		_w9417_
	);
	LUT2 #(
		.INIT('h1)
	) name8886 (
		_w9413_,
		_w9417_,
		_w9418_
	);
	LUT2 #(
		.INIT('h8)
	) name8887 (
		_w8519_,
		_w8660_,
		_w9419_
	);
	LUT2 #(
		.INIT('h8)
	) name8888 (
		_w8547_,
		_w8569_,
		_w9420_
	);
	LUT2 #(
		.INIT('h1)
	) name8889 (
		_w8514_,
		_w9420_,
		_w9421_
	);
	LUT2 #(
		.INIT('h1)
	) name8890 (
		\sa23_reg[2]/P0001 ,
		_w9421_,
		_w9422_
	);
	LUT2 #(
		.INIT('h2)
	) name8891 (
		\sa23_reg[1]/P0001 ,
		_w9419_,
		_w9423_
	);
	LUT2 #(
		.INIT('h4)
	) name8892 (
		_w8609_,
		_w9423_,
		_w9424_
	);
	LUT2 #(
		.INIT('h4)
	) name8893 (
		_w8636_,
		_w9424_,
		_w9425_
	);
	LUT2 #(
		.INIT('h4)
	) name8894 (
		_w9422_,
		_w9425_,
		_w9426_
	);
	LUT2 #(
		.INIT('h1)
	) name8895 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w9427_
	);
	LUT2 #(
		.INIT('h1)
	) name8896 (
		\sa23_reg[3]/P0001 ,
		_w9427_,
		_w9428_
	);
	LUT2 #(
		.INIT('h2)
	) name8897 (
		_w8531_,
		_w9428_,
		_w9429_
	);
	LUT2 #(
		.INIT('h8)
	) name8898 (
		_w8519_,
		_w8588_,
		_w9430_
	);
	LUT2 #(
		.INIT('h4)
	) name8899 (
		\sa23_reg[2]/P0001 ,
		_w8625_,
		_w9431_
	);
	LUT2 #(
		.INIT('h1)
	) name8900 (
		\sa23_reg[1]/P0001 ,
		_w9431_,
		_w9432_
	);
	LUT2 #(
		.INIT('h8)
	) name8901 (
		\sa23_reg[2]/P0001 ,
		_w8570_,
		_w9433_
	);
	LUT2 #(
		.INIT('h1)
	) name8902 (
		_w9429_,
		_w9430_,
		_w9434_
	);
	LUT2 #(
		.INIT('h4)
	) name8903 (
		_w9433_,
		_w9434_,
		_w9435_
	);
	LUT2 #(
		.INIT('h8)
	) name8904 (
		_w9432_,
		_w9435_,
		_w9436_
	);
	LUT2 #(
		.INIT('h1)
	) name8905 (
		_w9426_,
		_w9436_,
		_w9437_
	);
	LUT2 #(
		.INIT('h2)
	) name8906 (
		\sa23_reg[2]/P0001 ,
		_w8615_,
		_w9438_
	);
	LUT2 #(
		.INIT('h1)
	) name8907 (
		_w8624_,
		_w8653_,
		_w9439_
	);
	LUT2 #(
		.INIT('h1)
	) name8908 (
		\sa23_reg[4]/P0001 ,
		_w9439_,
		_w9440_
	);
	LUT2 #(
		.INIT('h4)
	) name8909 (
		_w8635_,
		_w9438_,
		_w9441_
	);
	LUT2 #(
		.INIT('h4)
	) name8910 (
		_w9440_,
		_w9441_,
		_w9442_
	);
	LUT2 #(
		.INIT('h1)
	) name8911 (
		_w8591_,
		_w9137_,
		_w9443_
	);
	LUT2 #(
		.INIT('h8)
	) name8912 (
		_w9098_,
		_w9443_,
		_w9444_
	);
	LUT2 #(
		.INIT('h1)
	) name8913 (
		_w9442_,
		_w9444_,
		_w9445_
	);
	LUT2 #(
		.INIT('h1)
	) name8914 (
		_w9437_,
		_w9445_,
		_w9446_
	);
	LUT2 #(
		.INIT('h2)
	) name8915 (
		\sa23_reg[0]/P0001 ,
		_w9446_,
		_w9447_
	);
	LUT2 #(
		.INIT('h1)
	) name8916 (
		_w8558_,
		_w9100_,
		_w9448_
	);
	LUT2 #(
		.INIT('h4)
	) name8917 (
		_w9137_,
		_w9448_,
		_w9449_
	);
	LUT2 #(
		.INIT('h1)
	) name8918 (
		\sa23_reg[2]/P0001 ,
		_w9449_,
		_w9450_
	);
	LUT2 #(
		.INIT('h8)
	) name8919 (
		_w8513_,
		_w9112_,
		_w9451_
	);
	LUT2 #(
		.INIT('h8)
	) name8920 (
		\sa23_reg[4]/P0001 ,
		_w9451_,
		_w9452_
	);
	LUT2 #(
		.INIT('h4)
	) name8921 (
		\sa23_reg[5]/P0001 ,
		_w8519_,
		_w9453_
	);
	LUT2 #(
		.INIT('h8)
	) name8922 (
		_w8624_,
		_w9453_,
		_w9454_
	);
	LUT2 #(
		.INIT('h8)
	) name8923 (
		\sa23_reg[7]/NET0131 ,
		_w9129_,
		_w9455_
	);
	LUT2 #(
		.INIT('h1)
	) name8924 (
		_w9141_,
		_w9452_,
		_w9456_
	);
	LUT2 #(
		.INIT('h1)
	) name8925 (
		_w9454_,
		_w9455_,
		_w9457_
	);
	LUT2 #(
		.INIT('h8)
	) name8926 (
		_w9456_,
		_w9457_,
		_w9458_
	);
	LUT2 #(
		.INIT('h4)
	) name8927 (
		_w9450_,
		_w9458_,
		_w9459_
	);
	LUT2 #(
		.INIT('h2)
	) name8928 (
		\sa23_reg[1]/P0001 ,
		_w9459_,
		_w9460_
	);
	LUT2 #(
		.INIT('h8)
	) name8929 (
		_w8533_,
		_w8546_,
		_w9461_
	);
	LUT2 #(
		.INIT('h8)
	) name8930 (
		_w8514_,
		_w8529_,
		_w9462_
	);
	LUT2 #(
		.INIT('h4)
	) name8931 (
		\sa23_reg[2]/P0001 ,
		_w9462_,
		_w9463_
	);
	LUT2 #(
		.INIT('h8)
	) name8932 (
		_w8508_,
		_w8523_,
		_w9464_
	);
	LUT2 #(
		.INIT('h2)
	) name8933 (
		\sa23_reg[2]/P0001 ,
		_w8590_,
		_w9465_
	);
	LUT2 #(
		.INIT('h8)
	) name8934 (
		_w8508_,
		_w8572_,
		_w9466_
	);
	LUT2 #(
		.INIT('h8)
	) name8935 (
		_w8547_,
		_w9066_,
		_w9467_
	);
	LUT2 #(
		.INIT('h4)
	) name8936 (
		\sa23_reg[5]/P0001 ,
		_w8603_,
		_w9468_
	);
	LUT2 #(
		.INIT('h4)
	) name8937 (
		\sa23_reg[6]/NET0131 ,
		_w9468_,
		_w9469_
	);
	LUT2 #(
		.INIT('h1)
	) name8938 (
		_w9064_,
		_w9466_,
		_w9470_
	);
	LUT2 #(
		.INIT('h2)
	) name8939 (
		_w9465_,
		_w9467_,
		_w9471_
	);
	LUT2 #(
		.INIT('h8)
	) name8940 (
		_w9470_,
		_w9471_,
		_w9472_
	);
	LUT2 #(
		.INIT('h4)
	) name8941 (
		_w9469_,
		_w9472_,
		_w9473_
	);
	LUT2 #(
		.INIT('h1)
	) name8942 (
		\sa23_reg[2]/P0001 ,
		_w9117_,
		_w9474_
	);
	LUT2 #(
		.INIT('h4)
	) name8943 (
		_w8577_,
		_w8642_,
		_w9475_
	);
	LUT2 #(
		.INIT('h8)
	) name8944 (
		\sa23_reg[6]/NET0131 ,
		_w9078_,
		_w9476_
	);
	LUT2 #(
		.INIT('h1)
	) name8945 (
		_w9475_,
		_w9476_,
		_w9477_
	);
	LUT2 #(
		.INIT('h8)
	) name8946 (
		_w9474_,
		_w9477_,
		_w9478_
	);
	LUT2 #(
		.INIT('h1)
	) name8947 (
		_w9473_,
		_w9478_,
		_w9479_
	);
	LUT2 #(
		.INIT('h1)
	) name8948 (
		_w9464_,
		_w9479_,
		_w9480_
	);
	LUT2 #(
		.INIT('h1)
	) name8949 (
		\sa23_reg[1]/P0001 ,
		_w9480_,
		_w9481_
	);
	LUT2 #(
		.INIT('h8)
	) name8950 (
		_w8508_,
		_w8577_,
		_w9482_
	);
	LUT2 #(
		.INIT('h1)
	) name8951 (
		_w8646_,
		_w9482_,
		_w9483_
	);
	LUT2 #(
		.INIT('h1)
	) name8952 (
		\sa23_reg[3]/P0001 ,
		_w9483_,
		_w9484_
	);
	LUT2 #(
		.INIT('h4)
	) name8953 (
		\sa23_reg[5]/P0001 ,
		_w8625_,
		_w9485_
	);
	LUT2 #(
		.INIT('h4)
	) name8954 (
		\sa23_reg[4]/P0001 ,
		_w8642_,
		_w9486_
	);
	LUT2 #(
		.INIT('h1)
	) name8955 (
		_w9485_,
		_w9486_,
		_w9487_
	);
	LUT2 #(
		.INIT('h2)
	) name8956 (
		\sa23_reg[2]/P0001 ,
		_w9487_,
		_w9488_
	);
	LUT2 #(
		.INIT('h4)
	) name8957 (
		\sa23_reg[5]/P0001 ,
		_w8528_,
		_w9489_
	);
	LUT2 #(
		.INIT('h1)
	) name8958 (
		_w8533_,
		_w9489_,
		_w9490_
	);
	LUT2 #(
		.INIT('h2)
	) name8959 (
		\sa23_reg[2]/P0001 ,
		_w9490_,
		_w9491_
	);
	LUT2 #(
		.INIT('h4)
	) name8960 (
		\sa23_reg[3]/P0001 ,
		_w8614_,
		_w9492_
	);
	LUT2 #(
		.INIT('h4)
	) name8961 (
		\sa23_reg[2]/P0001 ,
		_w9492_,
		_w9493_
	);
	LUT2 #(
		.INIT('h1)
	) name8962 (
		_w9149_,
		_w9491_,
		_w9494_
	);
	LUT2 #(
		.INIT('h4)
	) name8963 (
		_w9493_,
		_w9494_,
		_w9495_
	);
	LUT2 #(
		.INIT('h1)
	) name8964 (
		\sa23_reg[1]/P0001 ,
		_w9495_,
		_w9496_
	);
	LUT2 #(
		.INIT('h2)
	) name8965 (
		\sa23_reg[2]/P0001 ,
		_w8614_,
		_w9497_
	);
	LUT2 #(
		.INIT('h8)
	) name8966 (
		_w8519_,
		_w8547_,
		_w9498_
	);
	LUT2 #(
		.INIT('h8)
	) name8967 (
		\sa23_reg[5]/P0001 ,
		_w8511_,
		_w9499_
	);
	LUT2 #(
		.INIT('h4)
	) name8968 (
		_w8572_,
		_w9499_,
		_w9500_
	);
	LUT2 #(
		.INIT('h1)
	) name8969 (
		\sa23_reg[2]/P0001 ,
		_w9498_,
		_w9501_
	);
	LUT2 #(
		.INIT('h4)
	) name8970 (
		_w9500_,
		_w9501_,
		_w9502_
	);
	LUT2 #(
		.INIT('h1)
	) name8971 (
		_w9497_,
		_w9502_,
		_w9503_
	);
	LUT2 #(
		.INIT('h8)
	) name8972 (
		_w8562_,
		_w8658_,
		_w9504_
	);
	LUT2 #(
		.INIT('h1)
	) name8973 (
		_w8604_,
		_w9504_,
		_w9505_
	);
	LUT2 #(
		.INIT('h4)
	) name8974 (
		_w9503_,
		_w9505_,
		_w9506_
	);
	LUT2 #(
		.INIT('h2)
	) name8975 (
		\sa23_reg[1]/P0001 ,
		_w9506_,
		_w9507_
	);
	LUT2 #(
		.INIT('h1)
	) name8976 (
		_w9484_,
		_w9488_,
		_w9508_
	);
	LUT2 #(
		.INIT('h4)
	) name8977 (
		_w9496_,
		_w9508_,
		_w9509_
	);
	LUT2 #(
		.INIT('h4)
	) name8978 (
		_w9507_,
		_w9509_,
		_w9510_
	);
	LUT2 #(
		.INIT('h1)
	) name8979 (
		\sa23_reg[0]/P0001 ,
		_w9510_,
		_w9511_
	);
	LUT2 #(
		.INIT('h1)
	) name8980 (
		_w9461_,
		_w9463_,
		_w9512_
	);
	LUT2 #(
		.INIT('h4)
	) name8981 (
		_w9460_,
		_w9512_,
		_w9513_
	);
	LUT2 #(
		.INIT('h4)
	) name8982 (
		_w9447_,
		_w9513_,
		_w9514_
	);
	LUT2 #(
		.INIT('h4)
	) name8983 (
		_w9481_,
		_w9514_,
		_w9515_
	);
	LUT2 #(
		.INIT('h4)
	) name8984 (
		_w9511_,
		_w9515_,
		_w9516_
	);
	LUT2 #(
		.INIT('h2)
	) name8985 (
		_w8213_,
		_w9516_,
		_w9517_
	);
	LUT2 #(
		.INIT('h4)
	) name8986 (
		_w8213_,
		_w9516_,
		_w9518_
	);
	LUT2 #(
		.INIT('h1)
	) name8987 (
		_w9517_,
		_w9518_,
		_w9519_
	);
	LUT2 #(
		.INIT('h1)
	) name8988 (
		_w9289_,
		_w9519_,
		_w9520_
	);
	LUT2 #(
		.INIT('h8)
	) name8989 (
		_w9289_,
		_w9519_,
		_w9521_
	);
	LUT2 #(
		.INIT('h1)
	) name8990 (
		_w9520_,
		_w9521_,
		_w9522_
	);
	LUT2 #(
		.INIT('h2)
	) name8991 (
		\u0_w_reg[1][21]/P0001 ,
		_w8853_,
		_w9523_
	);
	LUT2 #(
		.INIT('h4)
	) name8992 (
		\u0_w_reg[1][21]/P0001 ,
		_w8853_,
		_w9524_
	);
	LUT2 #(
		.INIT('h1)
	) name8993 (
		_w9523_,
		_w9524_,
		_w9525_
	);
	LUT2 #(
		.INIT('h8)
	) name8994 (
		_w8678_,
		_w9525_,
		_w9526_
	);
	LUT2 #(
		.INIT('h1)
	) name8995 (
		_w8678_,
		_w9525_,
		_w9527_
	);
	LUT2 #(
		.INIT('h1)
	) name8996 (
		_w9526_,
		_w9527_,
		_w9528_
	);
	LUT2 #(
		.INIT('h1)
	) name8997 (
		_w9522_,
		_w9528_,
		_w9529_
	);
	LUT2 #(
		.INIT('h8)
	) name8998 (
		_w9522_,
		_w9528_,
		_w9530_
	);
	LUT2 #(
		.INIT('h1)
	) name8999 (
		\ld_r_reg/P0001 ,
		_w9529_,
		_w9531_
	);
	LUT2 #(
		.INIT('h4)
	) name9000 (
		_w9530_,
		_w9531_,
		_w9532_
	);
	LUT2 #(
		.INIT('h2)
	) name9001 (
		\text_in_r_reg[85]/P0001 ,
		\u0_w_reg[1][21]/P0001 ,
		_w9533_
	);
	LUT2 #(
		.INIT('h4)
	) name9002 (
		\text_in_r_reg[85]/P0001 ,
		\u0_w_reg[1][21]/P0001 ,
		_w9534_
	);
	LUT2 #(
		.INIT('h2)
	) name9003 (
		\ld_r_reg/P0001 ,
		_w9533_,
		_w9535_
	);
	LUT2 #(
		.INIT('h4)
	) name9004 (
		_w9534_,
		_w9535_,
		_w9536_
	);
	LUT2 #(
		.INIT('h1)
	) name9005 (
		_w9532_,
		_w9536_,
		_w9537_
	);
	LUT2 #(
		.INIT('h1)
	) name9006 (
		_w9292_,
		_w9516_,
		_w9538_
	);
	LUT2 #(
		.INIT('h8)
	) name9007 (
		_w9292_,
		_w9516_,
		_w9539_
	);
	LUT2 #(
		.INIT('h1)
	) name9008 (
		_w9538_,
		_w9539_,
		_w9540_
	);
	LUT2 #(
		.INIT('h4)
	) name9009 (
		\sa30_reg[3]/P0001 ,
		_w8765_,
		_w9541_
	);
	LUT2 #(
		.INIT('h2)
	) name9010 (
		_w8692_,
		_w8725_,
		_w9542_
	);
	LUT2 #(
		.INIT('h4)
	) name9011 (
		\sa30_reg[4]/P0001 ,
		_w8813_,
		_w9543_
	);
	LUT2 #(
		.INIT('h1)
	) name9012 (
		_w9542_,
		_w9543_,
		_w9544_
	);
	LUT2 #(
		.INIT('h1)
	) name9013 (
		\sa30_reg[2]/P0001 ,
		_w9544_,
		_w9545_
	);
	LUT2 #(
		.INIT('h8)
	) name9014 (
		\sa30_reg[2]/P0001 ,
		_w8705_,
		_w9546_
	);
	LUT2 #(
		.INIT('h8)
	) name9015 (
		\sa30_reg[4]/P0001 ,
		_w8874_,
		_w9547_
	);
	LUT2 #(
		.INIT('h8)
	) name9016 (
		_w8929_,
		_w9547_,
		_w9548_
	);
	LUT2 #(
		.INIT('h1)
	) name9017 (
		_w8889_,
		_w9546_,
		_w9549_
	);
	LUT2 #(
		.INIT('h4)
	) name9018 (
		_w9548_,
		_w9549_,
		_w9550_
	);
	LUT2 #(
		.INIT('h4)
	) name9019 (
		_w9545_,
		_w9550_,
		_w9551_
	);
	LUT2 #(
		.INIT('h2)
	) name9020 (
		\sa30_reg[1]/P0001 ,
		_w9551_,
		_w9552_
	);
	LUT2 #(
		.INIT('h8)
	) name9021 (
		\sa30_reg[2]/P0001 ,
		_w8950_,
		_w9553_
	);
	LUT2 #(
		.INIT('h4)
	) name9022 (
		\sa30_reg[7]/P0001 ,
		_w8833_,
		_w9554_
	);
	LUT2 #(
		.INIT('h1)
	) name9023 (
		_w8811_,
		_w9554_,
		_w9555_
	);
	LUT2 #(
		.INIT('h2)
	) name9024 (
		_w8697_,
		_w9555_,
		_w9556_
	);
	LUT2 #(
		.INIT('h1)
	) name9025 (
		_w8953_,
		_w9553_,
		_w9557_
	);
	LUT2 #(
		.INIT('h4)
	) name9026 (
		_w9556_,
		_w9557_,
		_w9558_
	);
	LUT2 #(
		.INIT('h1)
	) name9027 (
		\sa30_reg[1]/P0001 ,
		_w9558_,
		_w9559_
	);
	LUT2 #(
		.INIT('h4)
	) name9028 (
		\sa30_reg[6]/NET0131 ,
		_w8695_,
		_w9560_
	);
	LUT2 #(
		.INIT('h8)
	) name9029 (
		_w8734_,
		_w9560_,
		_w9561_
	);
	LUT2 #(
		.INIT('h8)
	) name9030 (
		_w8698_,
		_w8792_,
		_w9562_
	);
	LUT2 #(
		.INIT('h1)
	) name9031 (
		_w9561_,
		_w9562_,
		_w9563_
	);
	LUT2 #(
		.INIT('h2)
	) name9032 (
		\sa30_reg[2]/P0001 ,
		_w9563_,
		_w9564_
	);
	LUT2 #(
		.INIT('h8)
	) name9033 (
		_w8684_,
		_w8698_,
		_w9565_
	);
	LUT2 #(
		.INIT('h4)
	) name9034 (
		\sa30_reg[7]/P0001 ,
		_w9565_,
		_w9566_
	);
	LUT2 #(
		.INIT('h1)
	) name9035 (
		_w9541_,
		_w9566_,
		_w9567_
	);
	LUT2 #(
		.INIT('h4)
	) name9036 (
		_w9564_,
		_w9567_,
		_w9568_
	);
	LUT2 #(
		.INIT('h4)
	) name9037 (
		_w9559_,
		_w9568_,
		_w9569_
	);
	LUT2 #(
		.INIT('h4)
	) name9038 (
		_w9552_,
		_w9569_,
		_w9570_
	);
	LUT2 #(
		.INIT('h1)
	) name9039 (
		\sa30_reg[0]/P0002 ,
		_w9570_,
		_w9571_
	);
	LUT2 #(
		.INIT('h8)
	) name9040 (
		\sa30_reg[4]/P0001 ,
		_w8813_,
		_w9572_
	);
	LUT2 #(
		.INIT('h1)
	) name9041 (
		_w8687_,
		_w9572_,
		_w9573_
	);
	LUT2 #(
		.INIT('h1)
	) name9042 (
		\sa30_reg[2]/P0001 ,
		_w9573_,
		_w9574_
	);
	LUT2 #(
		.INIT('h2)
	) name9043 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w9575_
	);
	LUT2 #(
		.INIT('h8)
	) name9044 (
		_w8682_,
		_w9575_,
		_w9576_
	);
	LUT2 #(
		.INIT('h2)
	) name9045 (
		\sa30_reg[1]/P0001 ,
		_w9576_,
		_w9577_
	);
	LUT2 #(
		.INIT('h4)
	) name9046 (
		_w8784_,
		_w9577_,
		_w9578_
	);
	LUT2 #(
		.INIT('h4)
	) name9047 (
		_w8831_,
		_w9578_,
		_w9579_
	);
	LUT2 #(
		.INIT('h4)
	) name9048 (
		_w9574_,
		_w9579_,
		_w9580_
	);
	LUT2 #(
		.INIT('h4)
	) name9049 (
		\sa30_reg[2]/P0001 ,
		_w8791_,
		_w9581_
	);
	LUT2 #(
		.INIT('h1)
	) name9050 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w9582_
	);
	LUT2 #(
		.INIT('h1)
	) name9051 (
		\sa30_reg[3]/P0001 ,
		_w9582_,
		_w9583_
	);
	LUT2 #(
		.INIT('h2)
	) name9052 (
		_w8694_,
		_w9583_,
		_w9584_
	);
	LUT2 #(
		.INIT('h8)
	) name9053 (
		_w8692_,
		_w8811_,
		_w9585_
	);
	LUT2 #(
		.INIT('h8)
	) name9054 (
		\sa30_reg[3]/P0001 ,
		_w8743_,
		_w9586_
	);
	LUT2 #(
		.INIT('h1)
	) name9055 (
		\sa30_reg[1]/P0001 ,
		_w9586_,
		_w9587_
	);
	LUT2 #(
		.INIT('h1)
	) name9056 (
		_w9581_,
		_w9584_,
		_w9588_
	);
	LUT2 #(
		.INIT('h4)
	) name9057 (
		_w9585_,
		_w9588_,
		_w9589_
	);
	LUT2 #(
		.INIT('h8)
	) name9058 (
		_w9587_,
		_w9589_,
		_w9590_
	);
	LUT2 #(
		.INIT('h1)
	) name9059 (
		_w9580_,
		_w9590_,
		_w9591_
	);
	LUT2 #(
		.INIT('h2)
	) name9060 (
		\sa30_reg[2]/P0001 ,
		_w8796_,
		_w9592_
	);
	LUT2 #(
		.INIT('h1)
	) name9061 (
		_w8726_,
		_w8783_,
		_w9593_
	);
	LUT2 #(
		.INIT('h4)
	) name9062 (
		_w8952_,
		_w9593_,
		_w9594_
	);
	LUT2 #(
		.INIT('h8)
	) name9063 (
		_w9592_,
		_w9594_,
		_w9595_
	);
	LUT2 #(
		.INIT('h8)
	) name9064 (
		_w8758_,
		_w8874_,
		_w9596_
	);
	LUT2 #(
		.INIT('h1)
	) name9065 (
		\sa30_reg[2]/P0001 ,
		_w8760_,
		_w9597_
	);
	LUT2 #(
		.INIT('h4)
	) name9066 (
		_w9596_,
		_w9597_,
		_w9598_
	);
	LUT2 #(
		.INIT('h4)
	) name9067 (
		_w8949_,
		_w9598_,
		_w9599_
	);
	LUT2 #(
		.INIT('h1)
	) name9068 (
		_w9595_,
		_w9599_,
		_w9600_
	);
	LUT2 #(
		.INIT('h1)
	) name9069 (
		_w9591_,
		_w9600_,
		_w9601_
	);
	LUT2 #(
		.INIT('h2)
	) name9070 (
		\sa30_reg[0]/P0002 ,
		_w9601_,
		_w9602_
	);
	LUT2 #(
		.INIT('h8)
	) name9071 (
		_w8695_,
		_w8709_,
		_w9603_
	);
	LUT2 #(
		.INIT('h4)
	) name9072 (
		\sa30_reg[5]/P0001 ,
		_w9603_,
		_w9604_
	);
	LUT2 #(
		.INIT('h1)
	) name9073 (
		_w8720_,
		_w8909_,
		_w9605_
	);
	LUT2 #(
		.INIT('h4)
	) name9074 (
		_w8949_,
		_w9605_,
		_w9606_
	);
	LUT2 #(
		.INIT('h1)
	) name9075 (
		\sa30_reg[2]/P0001 ,
		_w9606_,
		_w9607_
	);
	LUT2 #(
		.INIT('h4)
	) name9076 (
		\sa30_reg[6]/NET0131 ,
		_w8922_,
		_w9608_
	);
	LUT2 #(
		.INIT('h2)
	) name9077 (
		\sa30_reg[1]/P0001 ,
		_w8836_,
		_w9609_
	);
	LUT2 #(
		.INIT('h1)
	) name9078 (
		_w8846_,
		_w9604_,
		_w9610_
	);
	LUT2 #(
		.INIT('h4)
	) name9079 (
		_w9608_,
		_w9610_,
		_w9611_
	);
	LUT2 #(
		.INIT('h8)
	) name9080 (
		_w9609_,
		_w9611_,
		_w9612_
	);
	LUT2 #(
		.INIT('h4)
	) name9081 (
		_w9607_,
		_w9612_,
		_w9613_
	);
	LUT2 #(
		.INIT('h8)
	) name9082 (
		\sa30_reg[4]/P0001 ,
		_w8792_,
		_w9614_
	);
	LUT2 #(
		.INIT('h1)
	) name9083 (
		_w8710_,
		_w9614_,
		_w9615_
	);
	LUT2 #(
		.INIT('h1)
	) name9084 (
		\sa30_reg[3]/P0001 ,
		_w9615_,
		_w9616_
	);
	LUT2 #(
		.INIT('h8)
	) name9085 (
		_w8709_,
		_w8773_,
		_w9617_
	);
	LUT2 #(
		.INIT('h1)
	) name9086 (
		\sa30_reg[2]/P0001 ,
		_w9617_,
		_w9618_
	);
	LUT2 #(
		.INIT('h4)
	) name9087 (
		_w9616_,
		_w9618_,
		_w9619_
	);
	LUT2 #(
		.INIT('h8)
	) name9088 (
		_w8684_,
		_w8725_,
		_w9620_
	);
	LUT2 #(
		.INIT('h1)
	) name9089 (
		_w8721_,
		_w8725_,
		_w9621_
	);
	LUT2 #(
		.INIT('h8)
	) name9090 (
		_w8813_,
		_w9621_,
		_w9622_
	);
	LUT2 #(
		.INIT('h2)
	) name9091 (
		\sa30_reg[2]/P0001 ,
		_w8759_,
		_w9623_
	);
	LUT2 #(
		.INIT('h4)
	) name9092 (
		_w9620_,
		_w9623_,
		_w9624_
	);
	LUT2 #(
		.INIT('h1)
	) name9093 (
		_w8894_,
		_w9622_,
		_w9625_
	);
	LUT2 #(
		.INIT('h8)
	) name9094 (
		_w9624_,
		_w9625_,
		_w9626_
	);
	LUT2 #(
		.INIT('h1)
	) name9095 (
		_w9619_,
		_w9626_,
		_w9627_
	);
	LUT2 #(
		.INIT('h1)
	) name9096 (
		\sa30_reg[1]/P0001 ,
		_w8822_,
		_w9628_
	);
	LUT2 #(
		.INIT('h4)
	) name9097 (
		_w9566_,
		_w9628_,
		_w9629_
	);
	LUT2 #(
		.INIT('h4)
	) name9098 (
		_w9627_,
		_w9629_,
		_w9630_
	);
	LUT2 #(
		.INIT('h1)
	) name9099 (
		_w9613_,
		_w9630_,
		_w9631_
	);
	LUT2 #(
		.INIT('h8)
	) name9100 (
		_w8734_,
		_w8758_,
		_w9632_
	);
	LUT2 #(
		.INIT('h1)
	) name9101 (
		\sa30_reg[2]/P0001 ,
		_w9632_,
		_w9633_
	);
	LUT2 #(
		.INIT('h2)
	) name9102 (
		\sa30_reg[2]/P0001 ,
		_w8821_,
		_w9634_
	);
	LUT2 #(
		.INIT('h1)
	) name9103 (
		_w8741_,
		_w9633_,
		_w9635_
	);
	LUT2 #(
		.INIT('h4)
	) name9104 (
		_w9634_,
		_w9635_,
		_w9636_
	);
	LUT2 #(
		.INIT('h1)
	) name9105 (
		_w9631_,
		_w9636_,
		_w9637_
	);
	LUT2 #(
		.INIT('h4)
	) name9106 (
		_w9571_,
		_w9637_,
		_w9638_
	);
	LUT2 #(
		.INIT('h4)
	) name9107 (
		_w9602_,
		_w9638_,
		_w9639_
	);
	LUT2 #(
		.INIT('h2)
	) name9108 (
		\u0_w_reg[1][13]/P0001 ,
		_w9639_,
		_w9640_
	);
	LUT2 #(
		.INIT('h4)
	) name9109 (
		\u0_w_reg[1][13]/P0001 ,
		_w9639_,
		_w9641_
	);
	LUT2 #(
		.INIT('h1)
	) name9110 (
		_w9640_,
		_w9641_,
		_w9642_
	);
	LUT2 #(
		.INIT('h8)
	) name9111 (
		_w8853_,
		_w9642_,
		_w9643_
	);
	LUT2 #(
		.INIT('h1)
	) name9112 (
		_w8853_,
		_w9642_,
		_w9644_
	);
	LUT2 #(
		.INIT('h1)
	) name9113 (
		_w9643_,
		_w9644_,
		_w9645_
	);
	LUT2 #(
		.INIT('h4)
	) name9114 (
		_w9540_,
		_w9645_,
		_w9646_
	);
	LUT2 #(
		.INIT('h2)
	) name9115 (
		_w9540_,
		_w9645_,
		_w9647_
	);
	LUT2 #(
		.INIT('h1)
	) name9116 (
		\ld_r_reg/P0001 ,
		_w9646_,
		_w9648_
	);
	LUT2 #(
		.INIT('h4)
	) name9117 (
		_w9647_,
		_w9648_,
		_w9649_
	);
	LUT2 #(
		.INIT('h1)
	) name9118 (
		\text_in_r_reg[77]/P0001 ,
		\u0_w_reg[1][13]/P0001 ,
		_w9650_
	);
	LUT2 #(
		.INIT('h8)
	) name9119 (
		\text_in_r_reg[77]/P0001 ,
		\u0_w_reg[1][13]/P0001 ,
		_w9651_
	);
	LUT2 #(
		.INIT('h2)
	) name9120 (
		\ld_r_reg/P0001 ,
		_w9650_,
		_w9652_
	);
	LUT2 #(
		.INIT('h4)
	) name9121 (
		_w9651_,
		_w9652_,
		_w9653_
	);
	LUT2 #(
		.INIT('h1)
	) name9122 (
		_w9649_,
		_w9653_,
		_w9654_
	);
	LUT2 #(
		.INIT('h2)
	) name9123 (
		_w9063_,
		_w9400_,
		_w9655_
	);
	LUT2 #(
		.INIT('h4)
	) name9124 (
		_w9063_,
		_w9400_,
		_w9656_
	);
	LUT2 #(
		.INIT('h1)
	) name9125 (
		_w9655_,
		_w9656_,
		_w9657_
	);
	LUT2 #(
		.INIT('h1)
	) name9126 (
		_w8678_,
		_w9657_,
		_w9658_
	);
	LUT2 #(
		.INIT('h8)
	) name9127 (
		_w8678_,
		_w9657_,
		_w9659_
	);
	LUT2 #(
		.INIT('h1)
	) name9128 (
		_w9658_,
		_w9659_,
		_w9660_
	);
	LUT2 #(
		.INIT('h2)
	) name9129 (
		\u0_w_reg[1][14]/P0001 ,
		_w8974_,
		_w9661_
	);
	LUT2 #(
		.INIT('h4)
	) name9130 (
		\u0_w_reg[1][14]/P0001 ,
		_w8974_,
		_w9662_
	);
	LUT2 #(
		.INIT('h1)
	) name9131 (
		_w9661_,
		_w9662_,
		_w9663_
	);
	LUT2 #(
		.INIT('h8)
	) name9132 (
		_w8853_,
		_w9663_,
		_w9664_
	);
	LUT2 #(
		.INIT('h1)
	) name9133 (
		_w8853_,
		_w9663_,
		_w9665_
	);
	LUT2 #(
		.INIT('h1)
	) name9134 (
		_w9664_,
		_w9665_,
		_w9666_
	);
	LUT2 #(
		.INIT('h1)
	) name9135 (
		_w9660_,
		_w9666_,
		_w9667_
	);
	LUT2 #(
		.INIT('h8)
	) name9136 (
		_w9660_,
		_w9666_,
		_w9668_
	);
	LUT2 #(
		.INIT('h1)
	) name9137 (
		\ld_r_reg/P0001 ,
		_w9667_,
		_w9669_
	);
	LUT2 #(
		.INIT('h4)
	) name9138 (
		_w9668_,
		_w9669_,
		_w9670_
	);
	LUT2 #(
		.INIT('h2)
	) name9139 (
		\text_in_r_reg[78]/P0001 ,
		\u0_w_reg[1][14]/P0001 ,
		_w9671_
	);
	LUT2 #(
		.INIT('h4)
	) name9140 (
		\text_in_r_reg[78]/P0001 ,
		\u0_w_reg[1][14]/P0001 ,
		_w9672_
	);
	LUT2 #(
		.INIT('h2)
	) name9141 (
		\ld_r_reg/P0001 ,
		_w9671_,
		_w9673_
	);
	LUT2 #(
		.INIT('h4)
	) name9142 (
		_w9672_,
		_w9673_,
		_w9674_
	);
	LUT2 #(
		.INIT('h1)
	) name9143 (
		_w9670_,
		_w9674_,
		_w9675_
	);
	LUT2 #(
		.INIT('h1)
	) name9144 (
		_w9289_,
		_w9657_,
		_w9676_
	);
	LUT2 #(
		.INIT('h8)
	) name9145 (
		_w9289_,
		_w9657_,
		_w9677_
	);
	LUT2 #(
		.INIT('h1)
	) name9146 (
		_w9676_,
		_w9677_,
		_w9678_
	);
	LUT2 #(
		.INIT('h2)
	) name9147 (
		\u0_w_reg[1][6]/P0001 ,
		_w9169_,
		_w9679_
	);
	LUT2 #(
		.INIT('h4)
	) name9148 (
		\u0_w_reg[1][6]/P0001 ,
		_w9169_,
		_w9680_
	);
	LUT2 #(
		.INIT('h1)
	) name9149 (
		_w9679_,
		_w9680_,
		_w9681_
	);
	LUT2 #(
		.INIT('h8)
	) name9150 (
		_w8853_,
		_w9681_,
		_w9682_
	);
	LUT2 #(
		.INIT('h1)
	) name9151 (
		_w8853_,
		_w9681_,
		_w9683_
	);
	LUT2 #(
		.INIT('h1)
	) name9152 (
		_w9682_,
		_w9683_,
		_w9684_
	);
	LUT2 #(
		.INIT('h4)
	) name9153 (
		_w9678_,
		_w9684_,
		_w9685_
	);
	LUT2 #(
		.INIT('h2)
	) name9154 (
		_w9678_,
		_w9684_,
		_w9686_
	);
	LUT2 #(
		.INIT('h1)
	) name9155 (
		\ld_r_reg/P0001 ,
		_w9685_,
		_w9687_
	);
	LUT2 #(
		.INIT('h4)
	) name9156 (
		_w9686_,
		_w9687_,
		_w9688_
	);
	LUT2 #(
		.INIT('h1)
	) name9157 (
		\text_in_r_reg[70]/P0001 ,
		\u0_w_reg[1][6]/P0001 ,
		_w9689_
	);
	LUT2 #(
		.INIT('h8)
	) name9158 (
		\text_in_r_reg[70]/P0001 ,
		\u0_w_reg[1][6]/P0001 ,
		_w9690_
	);
	LUT2 #(
		.INIT('h2)
	) name9159 (
		\ld_r_reg/P0001 ,
		_w9689_,
		_w9691_
	);
	LUT2 #(
		.INIT('h4)
	) name9160 (
		_w9690_,
		_w9691_,
		_w9692_
	);
	LUT2 #(
		.INIT('h1)
	) name9161 (
		_w9688_,
		_w9692_,
		_w9693_
	);
	LUT2 #(
		.INIT('h1)
	) name9162 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		_w9694_
	);
	LUT2 #(
		.INIT('h8)
	) name9163 (
		_w8344_,
		_w9694_,
		_w9695_
	);
	LUT2 #(
		.INIT('h1)
	) name9164 (
		_w8332_,
		_w9695_,
		_w9696_
	);
	LUT2 #(
		.INIT('h2)
	) name9165 (
		\sa01_reg[1]/P0001 ,
		_w9696_,
		_w9697_
	);
	LUT2 #(
		.INIT('h8)
	) name9166 (
		\sa01_reg[2]/P0001 ,
		_w8218_,
		_w9698_
	);
	LUT2 #(
		.INIT('h8)
	) name9167 (
		_w8310_,
		_w9698_,
		_w9699_
	);
	LUT2 #(
		.INIT('h8)
	) name9168 (
		_w8326_,
		_w9209_,
		_w9700_
	);
	LUT2 #(
		.INIT('h1)
	) name9169 (
		_w8225_,
		_w9352_,
		_w9701_
	);
	LUT2 #(
		.INIT('h4)
	) name9170 (
		\sa01_reg[7]/NET0131 ,
		_w8264_,
		_w9702_
	);
	LUT2 #(
		.INIT('h1)
	) name9171 (
		_w8339_,
		_w9702_,
		_w9703_
	);
	LUT2 #(
		.INIT('h8)
	) name9172 (
		_w9701_,
		_w9703_,
		_w9704_
	);
	LUT2 #(
		.INIT('h2)
	) name9173 (
		_w9388_,
		_w9704_,
		_w9705_
	);
	LUT2 #(
		.INIT('h8)
	) name9174 (
		\sa01_reg[7]/NET0131 ,
		_w8304_,
		_w9706_
	);
	LUT2 #(
		.INIT('h1)
	) name9175 (
		_w9176_,
		_w9185_,
		_w9707_
	);
	LUT2 #(
		.INIT('h4)
	) name9176 (
		_w9706_,
		_w9707_,
		_w9708_
	);
	LUT2 #(
		.INIT('h2)
	) name9177 (
		\sa01_reg[2]/P0001 ,
		_w9708_,
		_w9709_
	);
	LUT2 #(
		.INIT('h8)
	) name9178 (
		_w8281_,
		_w8351_,
		_w9710_
	);
	LUT2 #(
		.INIT('h2)
	) name9179 (
		\sa01_reg[2]/P0001 ,
		_w9710_,
		_w9711_
	);
	LUT2 #(
		.INIT('h1)
	) name9180 (
		_w9244_,
		_w9711_,
		_w9712_
	);
	LUT2 #(
		.INIT('h4)
	) name9181 (
		_w8222_,
		_w8326_,
		_w9713_
	);
	LUT2 #(
		.INIT('h1)
	) name9182 (
		_w8295_,
		_w9175_,
		_w9714_
	);
	LUT2 #(
		.INIT('h4)
	) name9183 (
		_w9352_,
		_w9714_,
		_w9715_
	);
	LUT2 #(
		.INIT('h1)
	) name9184 (
		\sa01_reg[2]/P0001 ,
		_w9715_,
		_w9716_
	);
	LUT2 #(
		.INIT('h1)
	) name9185 (
		_w8341_,
		_w9713_,
		_w9717_
	);
	LUT2 #(
		.INIT('h4)
	) name9186 (
		_w9712_,
		_w9717_,
		_w9718_
	);
	LUT2 #(
		.INIT('h4)
	) name9187 (
		_w9716_,
		_w9718_,
		_w9719_
	);
	LUT2 #(
		.INIT('h1)
	) name9188 (
		\sa01_reg[1]/P0001 ,
		_w9719_,
		_w9720_
	);
	LUT2 #(
		.INIT('h1)
	) name9189 (
		_w9356_,
		_w9699_,
		_w9721_
	);
	LUT2 #(
		.INIT('h4)
	) name9190 (
		_w9700_,
		_w9721_,
		_w9722_
	);
	LUT2 #(
		.INIT('h4)
	) name9191 (
		_w9697_,
		_w9722_,
		_w9723_
	);
	LUT2 #(
		.INIT('h4)
	) name9192 (
		_w9705_,
		_w9723_,
		_w9724_
	);
	LUT2 #(
		.INIT('h4)
	) name9193 (
		_w9709_,
		_w9724_,
		_w9725_
	);
	LUT2 #(
		.INIT('h4)
	) name9194 (
		_w9720_,
		_w9725_,
		_w9726_
	);
	LUT2 #(
		.INIT('h2)
	) name9195 (
		\sa01_reg[0]/P0001 ,
		_w9726_,
		_w9727_
	);
	LUT2 #(
		.INIT('h1)
	) name9196 (
		_w8369_,
		_w9373_,
		_w9728_
	);
	LUT2 #(
		.INIT('h2)
	) name9197 (
		_w8242_,
		_w8281_,
		_w9729_
	);
	LUT2 #(
		.INIT('h2)
	) name9198 (
		_w9728_,
		_w9729_,
		_w9730_
	);
	LUT2 #(
		.INIT('h2)
	) name9199 (
		_w9386_,
		_w9730_,
		_w9731_
	);
	LUT2 #(
		.INIT('h2)
	) name9200 (
		\sa01_reg[7]/NET0131 ,
		_w9701_,
		_w9732_
	);
	LUT2 #(
		.INIT('h1)
	) name9201 (
		_w8309_,
		_w9732_,
		_w9733_
	);
	LUT2 #(
		.INIT('h1)
	) name9202 (
		\sa01_reg[3]/P0001 ,
		_w9733_,
		_w9734_
	);
	LUT2 #(
		.INIT('h1)
	) name9203 (
		_w8343_,
		_w9212_,
		_w9735_
	);
	LUT2 #(
		.INIT('h4)
	) name9204 (
		_w9734_,
		_w9735_,
		_w9736_
	);
	LUT2 #(
		.INIT('h2)
	) name9205 (
		\sa01_reg[2]/P0001 ,
		_w9736_,
		_w9737_
	);
	LUT2 #(
		.INIT('h1)
	) name9206 (
		_w9731_,
		_w9737_,
		_w9738_
	);
	LUT2 #(
		.INIT('h2)
	) name9207 (
		\sa01_reg[1]/P0001 ,
		_w9738_,
		_w9739_
	);
	LUT2 #(
		.INIT('h4)
	) name9208 (
		_w8240_,
		_w8356_,
		_w9740_
	);
	LUT2 #(
		.INIT('h8)
	) name9209 (
		_w8276_,
		_w8318_,
		_w9741_
	);
	LUT2 #(
		.INIT('h1)
	) name9210 (
		_w8239_,
		_w9741_,
		_w9742_
	);
	LUT2 #(
		.INIT('h1)
	) name9211 (
		\sa01_reg[2]/P0001 ,
		_w9742_,
		_w9743_
	);
	LUT2 #(
		.INIT('h2)
	) name9212 (
		\sa01_reg[1]/P0001 ,
		_w9369_,
		_w9744_
	);
	LUT2 #(
		.INIT('h4)
	) name9213 (
		_w9740_,
		_w9744_,
		_w9745_
	);
	LUT2 #(
		.INIT('h4)
	) name9214 (
		_w9743_,
		_w9745_,
		_w9746_
	);
	LUT2 #(
		.INIT('h1)
	) name9215 (
		_w8215_,
		_w9319_,
		_w9747_
	);
	LUT2 #(
		.INIT('h2)
	) name9216 (
		_w8303_,
		_w9747_,
		_w9748_
	);
	LUT2 #(
		.INIT('h4)
	) name9217 (
		\sa01_reg[2]/P0001 ,
		_w8281_,
		_w9749_
	);
	LUT2 #(
		.INIT('h1)
	) name9218 (
		\sa01_reg[1]/P0001 ,
		_w9315_,
		_w9750_
	);
	LUT2 #(
		.INIT('h4)
	) name9219 (
		_w9749_,
		_w9750_,
		_w9751_
	);
	LUT2 #(
		.INIT('h4)
	) name9220 (
		_w9748_,
		_w9751_,
		_w9752_
	);
	LUT2 #(
		.INIT('h1)
	) name9221 (
		_w9746_,
		_w9752_,
		_w9753_
	);
	LUT2 #(
		.INIT('h8)
	) name9222 (
		_w8224_,
		_w8257_,
		_w9754_
	);
	LUT2 #(
		.INIT('h1)
	) name9223 (
		_w9276_,
		_w9754_,
		_w9755_
	);
	LUT2 #(
		.INIT('h2)
	) name9224 (
		_w8329_,
		_w9755_,
		_w9756_
	);
	LUT2 #(
		.INIT('h8)
	) name9225 (
		_w8329_,
		_w9219_,
		_w9757_
	);
	LUT2 #(
		.INIT('h1)
	) name9226 (
		_w8361_,
		_w9389_,
		_w9758_
	);
	LUT2 #(
		.INIT('h1)
	) name9227 (
		\sa01_reg[2]/P0001 ,
		_w9758_,
		_w9759_
	);
	LUT2 #(
		.INIT('h1)
	) name9228 (
		_w8258_,
		_w9231_,
		_w9760_
	);
	LUT2 #(
		.INIT('h2)
	) name9229 (
		_w9694_,
		_w9760_,
		_w9761_
	);
	LUT2 #(
		.INIT('h1)
	) name9230 (
		_w9757_,
		_w9761_,
		_w9762_
	);
	LUT2 #(
		.INIT('h4)
	) name9231 (
		_w9756_,
		_w9762_,
		_w9763_
	);
	LUT2 #(
		.INIT('h4)
	) name9232 (
		_w9759_,
		_w9763_,
		_w9764_
	);
	LUT2 #(
		.INIT('h4)
	) name9233 (
		_w9753_,
		_w9764_,
		_w9765_
	);
	LUT2 #(
		.INIT('h1)
	) name9234 (
		\sa01_reg[0]/P0001 ,
		_w9765_,
		_w9766_
	);
	LUT2 #(
		.INIT('h4)
	) name9235 (
		\sa01_reg[5]/P0001 ,
		_w8305_,
		_w9767_
	);
	LUT2 #(
		.INIT('h1)
	) name9236 (
		_w9181_,
		_w9767_,
		_w9768_
	);
	LUT2 #(
		.INIT('h1)
	) name9237 (
		\sa01_reg[2]/P0001 ,
		_w9768_,
		_w9769_
	);
	LUT2 #(
		.INIT('h4)
	) name9238 (
		\sa01_reg[3]/P0001 ,
		_w8295_,
		_w9770_
	);
	LUT2 #(
		.INIT('h1)
	) name9239 (
		_w8332_,
		_w9179_,
		_w9771_
	);
	LUT2 #(
		.INIT('h4)
	) name9240 (
		_w9770_,
		_w9771_,
		_w9772_
	);
	LUT2 #(
		.INIT('h2)
	) name9241 (
		\sa01_reg[2]/P0001 ,
		_w9772_,
		_w9773_
	);
	LUT2 #(
		.INIT('h8)
	) name9242 (
		_w8214_,
		_w8245_,
		_w9774_
	);
	LUT2 #(
		.INIT('h8)
	) name9243 (
		_w8282_,
		_w9386_,
		_w9775_
	);
	LUT2 #(
		.INIT('h1)
	) name9244 (
		_w9774_,
		_w9775_,
		_w9776_
	);
	LUT2 #(
		.INIT('h4)
	) name9245 (
		_w9761_,
		_w9776_,
		_w9777_
	);
	LUT2 #(
		.INIT('h4)
	) name9246 (
		_w9773_,
		_w9777_,
		_w9778_
	);
	LUT2 #(
		.INIT('h1)
	) name9247 (
		\sa01_reg[1]/P0001 ,
		_w9778_,
		_w9779_
	);
	LUT2 #(
		.INIT('h1)
	) name9248 (
		_w9769_,
		_w9779_,
		_w9780_
	);
	LUT2 #(
		.INIT('h4)
	) name9249 (
		_w9766_,
		_w9780_,
		_w9781_
	);
	LUT2 #(
		.INIT('h4)
	) name9250 (
		_w9727_,
		_w9781_,
		_w9782_
	);
	LUT2 #(
		.INIT('h4)
	) name9251 (
		_w9739_,
		_w9782_,
		_w9783_
	);
	LUT2 #(
		.INIT('h1)
	) name9252 (
		_w8070_,
		_w9044_,
		_w9784_
	);
	LUT2 #(
		.INIT('h2)
	) name9253 (
		_w8077_,
		_w8111_,
		_w9785_
	);
	LUT2 #(
		.INIT('h2)
	) name9254 (
		_w9784_,
		_w9785_,
		_w9786_
	);
	LUT2 #(
		.INIT('h2)
	) name9255 (
		_w8155_,
		_w9786_,
		_w9787_
	);
	LUT2 #(
		.INIT('h1)
	) name9256 (
		_w8068_,
		_w9025_,
		_w9788_
	);
	LUT2 #(
		.INIT('h2)
	) name9257 (
		\sa12_reg[7]/NET0131 ,
		_w9788_,
		_w9789_
	);
	LUT2 #(
		.INIT('h8)
	) name9258 (
		_w8077_,
		_w8498_,
		_w9790_
	);
	LUT2 #(
		.INIT('h1)
	) name9259 (
		_w9789_,
		_w9790_,
		_w9791_
	);
	LUT2 #(
		.INIT('h1)
	) name9260 (
		\sa12_reg[3]/P0001 ,
		_w9791_,
		_w9792_
	);
	LUT2 #(
		.INIT('h1)
	) name9261 (
		_w8076_,
		_w8422_,
		_w9793_
	);
	LUT2 #(
		.INIT('h4)
	) name9262 (
		_w9792_,
		_w9793_,
		_w9794_
	);
	LUT2 #(
		.INIT('h2)
	) name9263 (
		\sa12_reg[2]/P0001 ,
		_w9794_,
		_w9795_
	);
	LUT2 #(
		.INIT('h1)
	) name9264 (
		_w9787_,
		_w9795_,
		_w9796_
	);
	LUT2 #(
		.INIT('h2)
	) name9265 (
		\sa12_reg[1]/P0001 ,
		_w9796_,
		_w9797_
	);
	LUT2 #(
		.INIT('h4)
	) name9266 (
		_w8135_,
		_w8390_,
		_w9798_
	);
	LUT2 #(
		.INIT('h1)
	) name9267 (
		_w9025_,
		_w9798_,
		_w9799_
	);
	LUT2 #(
		.INIT('h1)
	) name9268 (
		\sa12_reg[2]/P0001 ,
		_w9799_,
		_w9800_
	);
	LUT2 #(
		.INIT('h8)
	) name9269 (
		_w8104_,
		_w8135_,
		_w9801_
	);
	LUT2 #(
		.INIT('h8)
	) name9270 (
		\sa12_reg[2]/P0001 ,
		_w9801_,
		_w9802_
	);
	LUT2 #(
		.INIT('h2)
	) name9271 (
		\sa12_reg[2]/P0001 ,
		_w8094_,
		_w9803_
	);
	LUT2 #(
		.INIT('h2)
	) name9272 (
		_w8060_,
		_w8110_,
		_w9804_
	);
	LUT2 #(
		.INIT('h4)
	) name9273 (
		_w9803_,
		_w9804_,
		_w9805_
	);
	LUT2 #(
		.INIT('h1)
	) name9274 (
		_w8079_,
		_w9802_,
		_w9806_
	);
	LUT2 #(
		.INIT('h4)
	) name9275 (
		_w9805_,
		_w9806_,
		_w9807_
	);
	LUT2 #(
		.INIT('h4)
	) name9276 (
		_w9800_,
		_w9807_,
		_w9808_
	);
	LUT2 #(
		.INIT('h1)
	) name9277 (
		\sa12_reg[1]/P0001 ,
		_w9808_,
		_w9809_
	);
	LUT2 #(
		.INIT('h8)
	) name9278 (
		_w8061_,
		_w8978_,
		_w9810_
	);
	LUT2 #(
		.INIT('h1)
	) name9279 (
		_w8084_,
		_w8110_,
		_w9811_
	);
	LUT2 #(
		.INIT('h2)
	) name9280 (
		_w8068_,
		_w9811_,
		_w9812_
	);
	LUT2 #(
		.INIT('h1)
	) name9281 (
		_w8380_,
		_w8391_,
		_w9813_
	);
	LUT2 #(
		.INIT('h4)
	) name9282 (
		_w9812_,
		_w9813_,
		_w9814_
	);
	LUT2 #(
		.INIT('h2)
	) name9283 (
		\sa12_reg[2]/P0001 ,
		_w9814_,
		_w9815_
	);
	LUT2 #(
		.INIT('h8)
	) name9284 (
		\sa12_reg[3]/P0001 ,
		_w8060_,
		_w9816_
	);
	LUT2 #(
		.INIT('h4)
	) name9285 (
		\sa12_reg[3]/P0001 ,
		_w8055_,
		_w9817_
	);
	LUT2 #(
		.INIT('h1)
	) name9286 (
		_w9816_,
		_w9817_,
		_w9818_
	);
	LUT2 #(
		.INIT('h8)
	) name9287 (
		_w9788_,
		_w9818_,
		_w9819_
	);
	LUT2 #(
		.INIT('h2)
	) name9288 (
		\sa12_reg[2]/P0001 ,
		_w9819_,
		_w9820_
	);
	LUT2 #(
		.INIT('h8)
	) name9289 (
		_w8135_,
		_w8978_,
		_w9821_
	);
	LUT2 #(
		.INIT('h4)
	) name9290 (
		\sa12_reg[6]/NET0131 ,
		_w9821_,
		_w9822_
	);
	LUT2 #(
		.INIT('h1)
	) name9291 (
		_w8109_,
		_w9822_,
		_w9823_
	);
	LUT2 #(
		.INIT('h4)
	) name9292 (
		_w9820_,
		_w9823_,
		_w9824_
	);
	LUT2 #(
		.INIT('h2)
	) name9293 (
		\sa12_reg[1]/P0001 ,
		_w9824_,
		_w9825_
	);
	LUT2 #(
		.INIT('h1)
	) name9294 (
		_w8494_,
		_w9810_,
		_w9826_
	);
	LUT2 #(
		.INIT('h4)
	) name9295 (
		_w9815_,
		_w9826_,
		_w9827_
	);
	LUT2 #(
		.INIT('h4)
	) name9296 (
		_w9809_,
		_w9827_,
		_w9828_
	);
	LUT2 #(
		.INIT('h4)
	) name9297 (
		_w9825_,
		_w9828_,
		_w9829_
	);
	LUT2 #(
		.INIT('h2)
	) name9298 (
		\sa12_reg[0]/P0001 ,
		_w9829_,
		_w9830_
	);
	LUT2 #(
		.INIT('h1)
	) name9299 (
		_w8432_,
		_w8490_,
		_w9831_
	);
	LUT2 #(
		.INIT('h2)
	) name9300 (
		_w8057_,
		_w9831_,
		_w9832_
	);
	LUT2 #(
		.INIT('h1)
	) name9301 (
		_w8103_,
		_w9034_,
		_w9833_
	);
	LUT2 #(
		.INIT('h1)
	) name9302 (
		\sa12_reg[2]/P0001 ,
		_w9833_,
		_w9834_
	);
	LUT2 #(
		.INIT('h1)
	) name9303 (
		_w8130_,
		_w8443_,
		_w9835_
	);
	LUT2 #(
		.INIT('h2)
	) name9304 (
		_w8978_,
		_w9835_,
		_w9836_
	);
	LUT2 #(
		.INIT('h8)
	) name9305 (
		_w8055_,
		_w8144_,
		_w9837_
	);
	LUT2 #(
		.INIT('h8)
	) name9306 (
		_w8110_,
		_w9837_,
		_w9838_
	);
	LUT2 #(
		.INIT('h1)
	) name9307 (
		_w8459_,
		_w9042_,
		_w9839_
	);
	LUT2 #(
		.INIT('h1)
	) name9308 (
		\sa12_reg[2]/P0001 ,
		_w9839_,
		_w9840_
	);
	LUT2 #(
		.INIT('h1)
	) name9309 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w9841_
	);
	LUT2 #(
		.INIT('h2)
	) name9310 (
		_w8095_,
		_w9841_,
		_w9842_
	);
	LUT2 #(
		.INIT('h1)
	) name9311 (
		_w9035_,
		_w9842_,
		_w9843_
	);
	LUT2 #(
		.INIT('h4)
	) name9312 (
		_w9840_,
		_w9843_,
		_w9844_
	);
	LUT2 #(
		.INIT('h2)
	) name9313 (
		\sa12_reg[1]/P0001 ,
		_w9844_,
		_w9845_
	);
	LUT2 #(
		.INIT('h4)
	) name9314 (
		\sa12_reg[2]/P0001 ,
		_w8111_,
		_w9846_
	);
	LUT2 #(
		.INIT('h8)
	) name9315 (
		_w8135_,
		_w8479_,
		_w9847_
	);
	LUT2 #(
		.INIT('h1)
	) name9316 (
		_w8985_,
		_w9846_,
		_w9848_
	);
	LUT2 #(
		.INIT('h4)
	) name9317 (
		_w8194_,
		_w9848_,
		_w9849_
	);
	LUT2 #(
		.INIT('h4)
	) name9318 (
		_w9847_,
		_w9849_,
		_w9850_
	);
	LUT2 #(
		.INIT('h1)
	) name9319 (
		\sa12_reg[1]/P0001 ,
		_w9850_,
		_w9851_
	);
	LUT2 #(
		.INIT('h1)
	) name9320 (
		_w9836_,
		_w9838_,
		_w9852_
	);
	LUT2 #(
		.INIT('h4)
	) name9321 (
		_w9832_,
		_w9852_,
		_w9853_
	);
	LUT2 #(
		.INIT('h4)
	) name9322 (
		_w9834_,
		_w9853_,
		_w9854_
	);
	LUT2 #(
		.INIT('h1)
	) name9323 (
		_w9845_,
		_w9851_,
		_w9855_
	);
	LUT2 #(
		.INIT('h8)
	) name9324 (
		_w9854_,
		_w9855_,
		_w9856_
	);
	LUT2 #(
		.INIT('h1)
	) name9325 (
		\sa12_reg[0]/P0001 ,
		_w9856_,
		_w9857_
	);
	LUT2 #(
		.INIT('h1)
	) name9326 (
		_w8201_,
		_w8395_,
		_w9858_
	);
	LUT2 #(
		.INIT('h1)
	) name9327 (
		\sa12_reg[2]/P0001 ,
		_w9858_,
		_w9859_
	);
	LUT2 #(
		.INIT('h8)
	) name9328 (
		\sa12_reg[4]/P0001 ,
		_w8065_,
		_w9860_
	);
	LUT2 #(
		.INIT('h4)
	) name9329 (
		\sa12_reg[3]/P0001 ,
		_w9860_,
		_w9861_
	);
	LUT2 #(
		.INIT('h1)
	) name9330 (
		_w8109_,
		_w8387_,
		_w9862_
	);
	LUT2 #(
		.INIT('h4)
	) name9331 (
		_w9861_,
		_w9862_,
		_w9863_
	);
	LUT2 #(
		.INIT('h2)
	) name9332 (
		\sa12_reg[2]/P0001 ,
		_w9863_,
		_w9864_
	);
	LUT2 #(
		.INIT('h8)
	) name9333 (
		_w8094_,
		_w8161_,
		_w9865_
	);
	LUT2 #(
		.INIT('h8)
	) name9334 (
		_w8110_,
		_w9846_,
		_w9866_
	);
	LUT2 #(
		.INIT('h1)
	) name9335 (
		_w9865_,
		_w9866_,
		_w9867_
	);
	LUT2 #(
		.INIT('h4)
	) name9336 (
		_w9836_,
		_w9867_,
		_w9868_
	);
	LUT2 #(
		.INIT('h4)
	) name9337 (
		_w9864_,
		_w9868_,
		_w9869_
	);
	LUT2 #(
		.INIT('h1)
	) name9338 (
		\sa12_reg[1]/P0001 ,
		_w9869_,
		_w9870_
	);
	LUT2 #(
		.INIT('h1)
	) name9339 (
		_w9859_,
		_w9870_,
		_w9871_
	);
	LUT2 #(
		.INIT('h4)
	) name9340 (
		_w9857_,
		_w9871_,
		_w9872_
	);
	LUT2 #(
		.INIT('h4)
	) name9341 (
		_w9797_,
		_w9872_,
		_w9873_
	);
	LUT2 #(
		.INIT('h4)
	) name9342 (
		_w9830_,
		_w9873_,
		_w9874_
	);
	LUT2 #(
		.INIT('h1)
	) name9343 (
		_w9783_,
		_w9874_,
		_w9875_
	);
	LUT2 #(
		.INIT('h8)
	) name9344 (
		_w9783_,
		_w9874_,
		_w9876_
	);
	LUT2 #(
		.INIT('h1)
	) name9345 (
		_w9875_,
		_w9876_,
		_w9877_
	);
	LUT2 #(
		.INIT('h1)
	) name9346 (
		_w9400_,
		_w9877_,
		_w9878_
	);
	LUT2 #(
		.INIT('h8)
	) name9347 (
		_w9400_,
		_w9877_,
		_w9879_
	);
	LUT2 #(
		.INIT('h1)
	) name9348 (
		_w9878_,
		_w9879_,
		_w9880_
	);
	LUT2 #(
		.INIT('h8)
	) name9349 (
		\sa23_reg[3]/P0001 ,
		_w8513_,
		_w9881_
	);
	LUT2 #(
		.INIT('h1)
	) name9350 (
		_w8552_,
		_w8556_,
		_w9882_
	);
	LUT2 #(
		.INIT('h1)
	) name9351 (
		_w9099_,
		_w9881_,
		_w9883_
	);
	LUT2 #(
		.INIT('h8)
	) name9352 (
		_w9882_,
		_w9883_,
		_w9884_
	);
	LUT2 #(
		.INIT('h2)
	) name9353 (
		\sa23_reg[1]/P0001 ,
		_w9884_,
		_w9885_
	);
	LUT2 #(
		.INIT('h8)
	) name9354 (
		\sa23_reg[7]/NET0131 ,
		_w8556_,
		_w9886_
	);
	LUT2 #(
		.INIT('h4)
	) name9355 (
		\sa23_reg[3]/P0001 ,
		_w9886_,
		_w9887_
	);
	LUT2 #(
		.INIT('h1)
	) name9356 (
		_w8510_,
		_w8534_,
		_w9888_
	);
	LUT2 #(
		.INIT('h4)
	) name9357 (
		_w9887_,
		_w9888_,
		_w9889_
	);
	LUT2 #(
		.INIT('h4)
	) name9358 (
		_w9885_,
		_w9889_,
		_w9890_
	);
	LUT2 #(
		.INIT('h2)
	) name9359 (
		\sa23_reg[2]/P0001 ,
		_w9890_,
		_w9891_
	);
	LUT2 #(
		.INIT('h8)
	) name9360 (
		_w9073_,
		_w9079_,
		_w9892_
	);
	LUT2 #(
		.INIT('h4)
	) name9361 (
		\sa23_reg[5]/P0001 ,
		_w8550_,
		_w9893_
	);
	LUT2 #(
		.INIT('h4)
	) name9362 (
		\sa23_reg[2]/P0001 ,
		_w9893_,
		_w9894_
	);
	LUT2 #(
		.INIT('h1)
	) name9363 (
		_w9455_,
		_w9894_,
		_w9895_
	);
	LUT2 #(
		.INIT('h2)
	) name9364 (
		\sa23_reg[1]/P0001 ,
		_w9895_,
		_w9896_
	);
	LUT2 #(
		.INIT('h8)
	) name9365 (
		\sa23_reg[2]/P0001 ,
		_w8572_,
		_w9897_
	);
	LUT2 #(
		.INIT('h8)
	) name9366 (
		_w8525_,
		_w9897_,
		_w9898_
	);
	LUT2 #(
		.INIT('h8)
	) name9367 (
		\sa23_reg[5]/P0001 ,
		_w8635_,
		_w9899_
	);
	LUT2 #(
		.INIT('h2)
	) name9368 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w9900_
	);
	LUT2 #(
		.INIT('h2)
	) name9369 (
		_w8513_,
		_w9900_,
		_w9901_
	);
	LUT2 #(
		.INIT('h8)
	) name9370 (
		\sa23_reg[2]/P0001 ,
		_w9453_,
		_w9902_
	);
	LUT2 #(
		.INIT('h1)
	) name9371 (
		_w9901_,
		_w9902_,
		_w9903_
	);
	LUT2 #(
		.INIT('h1)
	) name9372 (
		\sa23_reg[3]/P0001 ,
		_w9903_,
		_w9904_
	);
	LUT2 #(
		.INIT('h4)
	) name9373 (
		_w8519_,
		_w8521_,
		_w9905_
	);
	LUT2 #(
		.INIT('h1)
	) name9374 (
		_w9073_,
		_w9099_,
		_w9906_
	);
	LUT2 #(
		.INIT('h4)
	) name9375 (
		_w9905_,
		_w9906_,
		_w9907_
	);
	LUT2 #(
		.INIT('h1)
	) name9376 (
		\sa23_reg[2]/P0001 ,
		_w9907_,
		_w9908_
	);
	LUT2 #(
		.INIT('h1)
	) name9377 (
		_w9466_,
		_w9904_,
		_w9909_
	);
	LUT2 #(
		.INIT('h4)
	) name9378 (
		_w9908_,
		_w9909_,
		_w9910_
	);
	LUT2 #(
		.INIT('h1)
	) name9379 (
		\sa23_reg[1]/P0001 ,
		_w9910_,
		_w9911_
	);
	LUT2 #(
		.INIT('h1)
	) name9380 (
		_w9892_,
		_w9898_,
		_w9912_
	);
	LUT2 #(
		.INIT('h4)
	) name9381 (
		_w9899_,
		_w9912_,
		_w9913_
	);
	LUT2 #(
		.INIT('h4)
	) name9382 (
		_w9896_,
		_w9913_,
		_w9914_
	);
	LUT2 #(
		.INIT('h4)
	) name9383 (
		_w9891_,
		_w9914_,
		_w9915_
	);
	LUT2 #(
		.INIT('h4)
	) name9384 (
		_w9911_,
		_w9915_,
		_w9916_
	);
	LUT2 #(
		.INIT('h2)
	) name9385 (
		\sa23_reg[0]/P0001 ,
		_w9916_,
		_w9917_
	);
	LUT2 #(
		.INIT('h8)
	) name9386 (
		_w8564_,
		_w8660_,
		_w9918_
	);
	LUT2 #(
		.INIT('h8)
	) name9387 (
		_w8572_,
		_w9918_,
		_w9919_
	);
	LUT2 #(
		.INIT('h8)
	) name9388 (
		\sa23_reg[4]/P0001 ,
		_w8562_,
		_w9920_
	);
	LUT2 #(
		.INIT('h8)
	) name9389 (
		_w8546_,
		_w9920_,
		_w9921_
	);
	LUT2 #(
		.INIT('h8)
	) name9390 (
		\sa23_reg[7]/NET0131 ,
		_w9427_,
		_w9922_
	);
	LUT2 #(
		.INIT('h1)
	) name9391 (
		\sa23_reg[1]/P0001 ,
		_w9078_,
		_w9923_
	);
	LUT2 #(
		.INIT('h1)
	) name9392 (
		_w9918_,
		_w9922_,
		_w9924_
	);
	LUT2 #(
		.INIT('h8)
	) name9393 (
		_w9923_,
		_w9924_,
		_w9925_
	);
	LUT2 #(
		.INIT('h4)
	) name9394 (
		_w9921_,
		_w9925_,
		_w9926_
	);
	LUT2 #(
		.INIT('h8)
	) name9395 (
		_w8513_,
		_w8529_,
		_w9927_
	);
	LUT2 #(
		.INIT('h4)
	) name9396 (
		\sa23_reg[6]/NET0131 ,
		_w8537_,
		_w9928_
	);
	LUT2 #(
		.INIT('h1)
	) name9397 (
		_w9927_,
		_w9928_,
		_w9929_
	);
	LUT2 #(
		.INIT('h1)
	) name9398 (
		\sa23_reg[2]/P0001 ,
		_w9929_,
		_w9930_
	);
	LUT2 #(
		.INIT('h8)
	) name9399 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w9931_
	);
	LUT2 #(
		.INIT('h1)
	) name9400 (
		_w8569_,
		_w9931_,
		_w9932_
	);
	LUT2 #(
		.INIT('h2)
	) name9401 (
		_w8642_,
		_w9932_,
		_w9933_
	);
	LUT2 #(
		.INIT('h2)
	) name9402 (
		\sa23_reg[1]/P0001 ,
		_w9154_,
		_w9934_
	);
	LUT2 #(
		.INIT('h4)
	) name9403 (
		_w9933_,
		_w9934_,
		_w9935_
	);
	LUT2 #(
		.INIT('h4)
	) name9404 (
		_w9930_,
		_w9935_,
		_w9936_
	);
	LUT2 #(
		.INIT('h1)
	) name9405 (
		_w9926_,
		_w9936_,
		_w9937_
	);
	LUT2 #(
		.INIT('h8)
	) name9406 (
		_w8521_,
		_w8569_,
		_w9938_
	);
	LUT2 #(
		.INIT('h1)
	) name9407 (
		_w8667_,
		_w9938_,
		_w9939_
	);
	LUT2 #(
		.INIT('h2)
	) name9408 (
		\sa23_reg[3]/P0001 ,
		_w9939_,
		_w9940_
	);
	LUT2 #(
		.INIT('h2)
	) name9409 (
		\sa23_reg[2]/P0001 ,
		_w9940_,
		_w9941_
	);
	LUT2 #(
		.INIT('h8)
	) name9410 (
		_w8521_,
		_w8526_,
		_w9942_
	);
	LUT2 #(
		.INIT('h8)
	) name9411 (
		_w8522_,
		_w8589_,
		_w9943_
	);
	LUT2 #(
		.INIT('h1)
	) name9412 (
		_w9942_,
		_w9943_,
		_w9944_
	);
	LUT2 #(
		.INIT('h4)
	) name9413 (
		_w9125_,
		_w9944_,
		_w9945_
	);
	LUT2 #(
		.INIT('h8)
	) name9414 (
		_w9474_,
		_w9945_,
		_w9946_
	);
	LUT2 #(
		.INIT('h1)
	) name9415 (
		_w9941_,
		_w9946_,
		_w9947_
	);
	LUT2 #(
		.INIT('h1)
	) name9416 (
		_w9919_,
		_w9947_,
		_w9948_
	);
	LUT2 #(
		.INIT('h4)
	) name9417 (
		_w9937_,
		_w9948_,
		_w9949_
	);
	LUT2 #(
		.INIT('h1)
	) name9418 (
		\sa23_reg[0]/P0001 ,
		_w9949_,
		_w9950_
	);
	LUT2 #(
		.INIT('h1)
	) name9419 (
		_w8524_,
		_w9485_,
		_w9951_
	);
	LUT2 #(
		.INIT('h1)
	) name9420 (
		\sa23_reg[2]/P0001 ,
		_w9951_,
		_w9952_
	);
	LUT2 #(
		.INIT('h2)
	) name9421 (
		\sa23_reg[2]/P0001 ,
		_w8619_,
		_w9953_
	);
	LUT2 #(
		.INIT('h1)
	) name9422 (
		\sa23_reg[1]/P0001 ,
		_w9953_,
		_w9954_
	);
	LUT2 #(
		.INIT('h1)
	) name9423 (
		_w8619_,
		_w9139_,
		_w9955_
	);
	LUT2 #(
		.INIT('h8)
	) name9424 (
		_w9944_,
		_w9955_,
		_w9956_
	);
	LUT2 #(
		.INIT('h2)
	) name9425 (
		_w9954_,
		_w9956_,
		_w9957_
	);
	LUT2 #(
		.INIT('h4)
	) name9426 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[2]/P0001 ,
		_w9958_
	);
	LUT2 #(
		.INIT('h8)
	) name9427 (
		\sa23_reg[5]/P0001 ,
		_w8574_,
		_w9959_
	);
	LUT2 #(
		.INIT('h1)
	) name9428 (
		_w8530_,
		_w9455_,
		_w9960_
	);
	LUT2 #(
		.INIT('h4)
	) name9429 (
		_w9959_,
		_w9960_,
		_w9961_
	);
	LUT2 #(
		.INIT('h2)
	) name9430 (
		_w9958_,
		_w9961_,
		_w9962_
	);
	LUT2 #(
		.INIT('h2)
	) name9431 (
		_w8508_,
		_w8519_,
		_w9963_
	);
	LUT2 #(
		.INIT('h8)
	) name9432 (
		_w8525_,
		_w8577_,
		_w9964_
	);
	LUT2 #(
		.INIT('h1)
	) name9433 (
		_w8557_,
		_w9964_,
		_w9965_
	);
	LUT2 #(
		.INIT('h4)
	) name9434 (
		_w9963_,
		_w9965_,
		_w9966_
	);
	LUT2 #(
		.INIT('h2)
	) name9435 (
		\sa23_reg[3]/P0001 ,
		_w9966_,
		_w9967_
	);
	LUT2 #(
		.INIT('h1)
	) name9436 (
		\sa23_reg[2]/P0001 ,
		_w9967_,
		_w9968_
	);
	LUT2 #(
		.INIT('h1)
	) name9437 (
		_w9420_,
		_w9482_,
		_w9969_
	);
	LUT2 #(
		.INIT('h4)
	) name9438 (
		_w9886_,
		_w9969_,
		_w9970_
	);
	LUT2 #(
		.INIT('h1)
	) name9439 (
		\sa23_reg[3]/P0001 ,
		_w9970_,
		_w9971_
	);
	LUT2 #(
		.INIT('h4)
	) name9440 (
		_w8563_,
		_w9465_,
		_w9972_
	);
	LUT2 #(
		.INIT('h4)
	) name9441 (
		_w9971_,
		_w9972_,
		_w9973_
	);
	LUT2 #(
		.INIT('h2)
	) name9442 (
		\sa23_reg[1]/P0001 ,
		_w9968_,
		_w9974_
	);
	LUT2 #(
		.INIT('h4)
	) name9443 (
		_w9973_,
		_w9974_,
		_w9975_
	);
	LUT2 #(
		.INIT('h1)
	) name9444 (
		_w9952_,
		_w9957_,
		_w9976_
	);
	LUT2 #(
		.INIT('h4)
	) name9445 (
		_w9962_,
		_w9976_,
		_w9977_
	);
	LUT2 #(
		.INIT('h4)
	) name9446 (
		_w9975_,
		_w9977_,
		_w9978_
	);
	LUT2 #(
		.INIT('h4)
	) name9447 (
		_w9950_,
		_w9978_,
		_w9979_
	);
	LUT2 #(
		.INIT('h4)
	) name9448 (
		_w9917_,
		_w9979_,
		_w9980_
	);
	LUT2 #(
		.INIT('h2)
	) name9449 (
		\u0_w_reg[1][7]/P0001 ,
		_w9980_,
		_w9981_
	);
	LUT2 #(
		.INIT('h4)
	) name9450 (
		\u0_w_reg[1][7]/P0001 ,
		_w9980_,
		_w9982_
	);
	LUT2 #(
		.INIT('h1)
	) name9451 (
		_w9981_,
		_w9982_,
		_w9983_
	);
	LUT2 #(
		.INIT('h8)
	) name9452 (
		_w8974_,
		_w9983_,
		_w9984_
	);
	LUT2 #(
		.INIT('h1)
	) name9453 (
		_w8974_,
		_w9983_,
		_w9985_
	);
	LUT2 #(
		.INIT('h1)
	) name9454 (
		_w9984_,
		_w9985_,
		_w9986_
	);
	LUT2 #(
		.INIT('h4)
	) name9455 (
		_w9880_,
		_w9986_,
		_w9987_
	);
	LUT2 #(
		.INIT('h2)
	) name9456 (
		_w9880_,
		_w9986_,
		_w9988_
	);
	LUT2 #(
		.INIT('h1)
	) name9457 (
		\ld_r_reg/P0001 ,
		_w9987_,
		_w9989_
	);
	LUT2 #(
		.INIT('h4)
	) name9458 (
		_w9988_,
		_w9989_,
		_w9990_
	);
	LUT2 #(
		.INIT('h2)
	) name9459 (
		\text_in_r_reg[71]/P0001 ,
		\u0_w_reg[1][7]/P0001 ,
		_w9991_
	);
	LUT2 #(
		.INIT('h4)
	) name9460 (
		\text_in_r_reg[71]/P0001 ,
		\u0_w_reg[1][7]/P0001 ,
		_w9992_
	);
	LUT2 #(
		.INIT('h2)
	) name9461 (
		\ld_r_reg/P0001 ,
		_w9991_,
		_w9993_
	);
	LUT2 #(
		.INIT('h4)
	) name9462 (
		_w9992_,
		_w9993_,
		_w9994_
	);
	LUT2 #(
		.INIT('h1)
	) name9463 (
		_w9990_,
		_w9994_,
		_w9995_
	);
	LUT2 #(
		.INIT('h8)
	) name9464 (
		_w8075_,
		_w8165_,
		_w9996_
	);
	LUT2 #(
		.INIT('h1)
	) name9465 (
		_w8422_,
		_w9996_,
		_w9997_
	);
	LUT2 #(
		.INIT('h1)
	) name9466 (
		_w8111_,
		_w8390_,
		_w9998_
	);
	LUT2 #(
		.INIT('h1)
	) name9467 (
		\sa12_reg[5]/P0001 ,
		_w9998_,
		_w9999_
	);
	LUT2 #(
		.INIT('h1)
	) name9468 (
		_w8159_,
		_w9999_,
		_w10000_
	);
	LUT2 #(
		.INIT('h2)
	) name9469 (
		\sa12_reg[2]/P0001 ,
		_w10000_,
		_w10001_
	);
	LUT2 #(
		.INIT('h2)
	) name9470 (
		_w9997_,
		_w10001_,
		_w10002_
	);
	LUT2 #(
		.INIT('h2)
	) name9471 (
		\sa12_reg[1]/P0001 ,
		_w10002_,
		_w10003_
	);
	LUT2 #(
		.INIT('h8)
	) name9472 (
		\sa12_reg[5]/P0001 ,
		_w9015_,
		_w10004_
	);
	LUT2 #(
		.INIT('h8)
	) name9473 (
		_w8074_,
		_w8180_,
		_w10005_
	);
	LUT2 #(
		.INIT('h4)
	) name9474 (
		_w8144_,
		_w8381_,
		_w10006_
	);
	LUT2 #(
		.INIT('h1)
	) name9475 (
		_w8070_,
		_w10005_,
		_w10007_
	);
	LUT2 #(
		.INIT('h4)
	) name9476 (
		_w10006_,
		_w10007_,
		_w10008_
	);
	LUT2 #(
		.INIT('h4)
	) name9477 (
		_w10004_,
		_w10008_,
		_w10009_
	);
	LUT2 #(
		.INIT('h1)
	) name9478 (
		\sa12_reg[1]/P0001 ,
		_w10009_,
		_w10010_
	);
	LUT2 #(
		.INIT('h2)
	) name9479 (
		_w8096_,
		_w8162_,
		_w10011_
	);
	LUT2 #(
		.INIT('h8)
	) name9480 (
		\sa12_reg[4]/P0001 ,
		_w8087_,
		_w10012_
	);
	LUT2 #(
		.INIT('h1)
	) name9481 (
		_w8070_,
		_w8175_,
		_w10013_
	);
	LUT2 #(
		.INIT('h1)
	) name9482 (
		_w8490_,
		_w9035_,
		_w10014_
	);
	LUT2 #(
		.INIT('h8)
	) name9483 (
		_w10013_,
		_w10014_,
		_w10015_
	);
	LUT2 #(
		.INIT('h1)
	) name9484 (
		\sa12_reg[2]/P0001 ,
		_w10015_,
		_w10016_
	);
	LUT2 #(
		.INIT('h1)
	) name9485 (
		_w10011_,
		_w10012_,
		_w10017_
	);
	LUT2 #(
		.INIT('h4)
	) name9486 (
		_w10010_,
		_w10017_,
		_w10018_
	);
	LUT2 #(
		.INIT('h4)
	) name9487 (
		_w10016_,
		_w10018_,
		_w10019_
	);
	LUT2 #(
		.INIT('h4)
	) name9488 (
		_w10003_,
		_w10019_,
		_w10020_
	);
	LUT2 #(
		.INIT('h2)
	) name9489 (
		\sa12_reg[0]/P0001 ,
		_w10020_,
		_w10021_
	);
	LUT2 #(
		.INIT('h1)
	) name9490 (
		_w8981_,
		_w9049_,
		_w10022_
	);
	LUT2 #(
		.INIT('h1)
	) name9491 (
		\sa12_reg[2]/P0001 ,
		_w10022_,
		_w10023_
	);
	LUT2 #(
		.INIT('h8)
	) name9492 (
		\sa12_reg[4]/P0001 ,
		_w9042_,
		_w10024_
	);
	LUT2 #(
		.INIT('h1)
	) name9493 (
		_w8136_,
		_w8175_,
		_w10025_
	);
	LUT2 #(
		.INIT('h2)
	) name9494 (
		\sa12_reg[2]/P0001 ,
		_w10025_,
		_w10026_
	);
	LUT2 #(
		.INIT('h1)
	) name9495 (
		_w8098_,
		_w10024_,
		_w10027_
	);
	LUT2 #(
		.INIT('h4)
	) name9496 (
		_w10023_,
		_w10027_,
		_w10028_
	);
	LUT2 #(
		.INIT('h4)
	) name9497 (
		_w10026_,
		_w10028_,
		_w10029_
	);
	LUT2 #(
		.INIT('h1)
	) name9498 (
		\sa12_reg[1]/P0001 ,
		_w10029_,
		_w10030_
	);
	LUT2 #(
		.INIT('h2)
	) name9499 (
		\sa12_reg[4]/P0001 ,
		_w8075_,
		_w10031_
	);
	LUT2 #(
		.INIT('h2)
	) name9500 (
		_w8979_,
		_w10031_,
		_w10032_
	);
	LUT2 #(
		.INIT('h1)
	) name9501 (
		_w8404_,
		_w10032_,
		_w10033_
	);
	LUT2 #(
		.INIT('h1)
	) name9502 (
		\sa12_reg[2]/P0001 ,
		_w10033_,
		_w10034_
	);
	LUT2 #(
		.INIT('h1)
	) name9503 (
		_w8114_,
		_w8165_,
		_w10035_
	);
	LUT2 #(
		.INIT('h2)
	) name9504 (
		\sa12_reg[2]/P0001 ,
		_w10035_,
		_w10036_
	);
	LUT2 #(
		.INIT('h4)
	) name9505 (
		_w8387_,
		_w8444_,
		_w10037_
	);
	LUT2 #(
		.INIT('h4)
	) name9506 (
		_w10036_,
		_w10037_,
		_w10038_
	);
	LUT2 #(
		.INIT('h4)
	) name9507 (
		_w10034_,
		_w10038_,
		_w10039_
	);
	LUT2 #(
		.INIT('h2)
	) name9508 (
		\sa12_reg[1]/P0001 ,
		_w10039_,
		_w10040_
	);
	LUT2 #(
		.INIT('h1)
	) name9509 (
		_w8142_,
		_w8498_,
		_w10041_
	);
	LUT2 #(
		.INIT('h2)
	) name9510 (
		_w8059_,
		_w10041_,
		_w10042_
	);
	LUT2 #(
		.INIT('h1)
	) name9511 (
		_w8098_,
		_w8461_,
		_w10043_
	);
	LUT2 #(
		.INIT('h1)
	) name9512 (
		\sa12_reg[2]/P0001 ,
		_w10043_,
		_w10044_
	);
	LUT2 #(
		.INIT('h1)
	) name9513 (
		_w8485_,
		_w8491_,
		_w10045_
	);
	LUT2 #(
		.INIT('h4)
	) name9514 (
		_w10042_,
		_w10045_,
		_w10046_
	);
	LUT2 #(
		.INIT('h4)
	) name9515 (
		_w10044_,
		_w10046_,
		_w10047_
	);
	LUT2 #(
		.INIT('h4)
	) name9516 (
		_w10040_,
		_w10047_,
		_w10048_
	);
	LUT2 #(
		.INIT('h4)
	) name9517 (
		_w10030_,
		_w10048_,
		_w10049_
	);
	LUT2 #(
		.INIT('h1)
	) name9518 (
		\sa12_reg[0]/P0001 ,
		_w10049_,
		_w10050_
	);
	LUT2 #(
		.INIT('h1)
	) name9519 (
		_w8422_,
		_w9860_,
		_w10051_
	);
	LUT2 #(
		.INIT('h2)
	) name9520 (
		\sa12_reg[3]/P0001 ,
		_w10051_,
		_w10052_
	);
	LUT2 #(
		.INIT('h1)
	) name9521 (
		_w8177_,
		_w10052_,
		_w10053_
	);
	LUT2 #(
		.INIT('h2)
	) name9522 (
		_w9033_,
		_w10053_,
		_w10054_
	);
	LUT2 #(
		.INIT('h4)
	) name9523 (
		\sa12_reg[3]/P0001 ,
		_w8077_,
		_w10055_
	);
	LUT2 #(
		.INIT('h1)
	) name9524 (
		_w8425_,
		_w10055_,
		_w10056_
	);
	LUT2 #(
		.INIT('h1)
	) name9525 (
		_w8080_,
		_w10056_,
		_w10057_
	);
	LUT2 #(
		.INIT('h1)
	) name9526 (
		_w8990_,
		_w10057_,
		_w10058_
	);
	LUT2 #(
		.INIT('h2)
	) name9527 (
		_w8455_,
		_w10058_,
		_w10059_
	);
	LUT2 #(
		.INIT('h1)
	) name9528 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[2]/P0001 ,
		_w10060_
	);
	LUT2 #(
		.INIT('h1)
	) name9529 (
		_w8066_,
		_w10060_,
		_w10061_
	);
	LUT2 #(
		.INIT('h8)
	) name9530 (
		_w8387_,
		_w10061_,
		_w10062_
	);
	LUT2 #(
		.INIT('h8)
	) name9531 (
		\sa12_reg[2]/P0001 ,
		_w8083_,
		_w10063_
	);
	LUT2 #(
		.INIT('h4)
	) name9532 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[2]/P0001 ,
		_w10064_
	);
	LUT2 #(
		.INIT('h1)
	) name9533 (
		_w8417_,
		_w8432_,
		_w10065_
	);
	LUT2 #(
		.INIT('h4)
	) name9534 (
		_w8481_,
		_w10065_,
		_w10066_
	);
	LUT2 #(
		.INIT('h4)
	) name9535 (
		\sa12_reg[3]/P0001 ,
		_w10064_,
		_w10067_
	);
	LUT2 #(
		.INIT('h4)
	) name9536 (
		_w10066_,
		_w10067_,
		_w10068_
	);
	LUT2 #(
		.INIT('h1)
	) name9537 (
		_w8985_,
		_w9042_,
		_w10069_
	);
	LUT2 #(
		.INIT('h4)
	) name9538 (
		_w8143_,
		_w10069_,
		_w10070_
	);
	LUT2 #(
		.INIT('h1)
	) name9539 (
		\sa12_reg[2]/P0001 ,
		_w10070_,
		_w10071_
	);
	LUT2 #(
		.INIT('h1)
	) name9540 (
		_w8083_,
		_w8460_,
		_w10072_
	);
	LUT2 #(
		.INIT('h4)
	) name9541 (
		_w10071_,
		_w10072_,
		_w10073_
	);
	LUT2 #(
		.INIT('h1)
	) name9542 (
		\sa12_reg[1]/P0001 ,
		_w10073_,
		_w10074_
	);
	LUT2 #(
		.INIT('h1)
	) name9543 (
		_w10062_,
		_w10063_,
		_w10075_
	);
	LUT2 #(
		.INIT('h4)
	) name9544 (
		_w10068_,
		_w10075_,
		_w10076_
	);
	LUT2 #(
		.INIT('h4)
	) name9545 (
		_w10054_,
		_w10076_,
		_w10077_
	);
	LUT2 #(
		.INIT('h4)
	) name9546 (
		_w10059_,
		_w10077_,
		_w10078_
	);
	LUT2 #(
		.INIT('h4)
	) name9547 (
		_w10074_,
		_w10078_,
		_w10079_
	);
	LUT2 #(
		.INIT('h4)
	) name9548 (
		_w10021_,
		_w10079_,
		_w10080_
	);
	LUT2 #(
		.INIT('h4)
	) name9549 (
		_w10050_,
		_w10080_,
		_w10081_
	);
	LUT2 #(
		.INIT('h4)
	) name9550 (
		_w8246_,
		_w8352_,
		_w10082_
	);
	LUT2 #(
		.INIT('h8)
	) name9551 (
		_w8238_,
		_w8258_,
		_w10083_
	);
	LUT2 #(
		.INIT('h1)
	) name9552 (
		_w9212_,
		_w10083_,
		_w10084_
	);
	LUT2 #(
		.INIT('h8)
	) name9553 (
		\sa01_reg[3]/P0001 ,
		_w8235_,
		_w10085_
	);
	LUT2 #(
		.INIT('h8)
	) name9554 (
		\sa01_reg[4]/P0001 ,
		_w8310_,
		_w10086_
	);
	LUT2 #(
		.INIT('h1)
	) name9555 (
		_w8282_,
		_w10085_,
		_w10087_
	);
	LUT2 #(
		.INIT('h4)
	) name9556 (
		_w10086_,
		_w10087_,
		_w10088_
	);
	LUT2 #(
		.INIT('h2)
	) name9557 (
		\sa01_reg[2]/P0001 ,
		_w10088_,
		_w10089_
	);
	LUT2 #(
		.INIT('h2)
	) name9558 (
		_w10084_,
		_w10089_,
		_w10090_
	);
	LUT2 #(
		.INIT('h2)
	) name9559 (
		\sa01_reg[1]/P0001 ,
		_w10090_,
		_w10091_
	);
	LUT2 #(
		.INIT('h4)
	) name9560 (
		\sa01_reg[3]/P0001 ,
		_w9276_,
		_w10092_
	);
	LUT2 #(
		.INIT('h2)
	) name9561 (
		\sa01_reg[2]/P0001 ,
		_w10092_,
		_w10093_
	);
	LUT2 #(
		.INIT('h1)
	) name9562 (
		_w8293_,
		_w8369_,
		_w10094_
	);
	LUT2 #(
		.INIT('h1)
	) name9563 (
		_w9276_,
		_w9369_,
		_w10095_
	);
	LUT2 #(
		.INIT('h8)
	) name9564 (
		_w10094_,
		_w10095_,
		_w10096_
	);
	LUT2 #(
		.INIT('h1)
	) name9565 (
		_w10093_,
		_w10096_,
		_w10097_
	);
	LUT2 #(
		.INIT('h4)
	) name9566 (
		_w8222_,
		_w9183_,
		_w10098_
	);
	LUT2 #(
		.INIT('h4)
	) name9567 (
		\sa01_reg[6]/NET0131 ,
		_w8321_,
		_w10099_
	);
	LUT2 #(
		.INIT('h1)
	) name9568 (
		_w8360_,
		_w8369_,
		_w10100_
	);
	LUT2 #(
		.INIT('h4)
	) name9569 (
		_w10098_,
		_w10100_,
		_w10101_
	);
	LUT2 #(
		.INIT('h4)
	) name9570 (
		_w10099_,
		_w10101_,
		_w10102_
	);
	LUT2 #(
		.INIT('h1)
	) name9571 (
		\sa01_reg[1]/P0001 ,
		_w10102_,
		_w10103_
	);
	LUT2 #(
		.INIT('h1)
	) name9572 (
		_w10082_,
		_w10097_,
		_w10104_
	);
	LUT2 #(
		.INIT('h4)
	) name9573 (
		_w10103_,
		_w10104_,
		_w10105_
	);
	LUT2 #(
		.INIT('h4)
	) name9574 (
		_w10091_,
		_w10105_,
		_w10106_
	);
	LUT2 #(
		.INIT('h2)
	) name9575 (
		\sa01_reg[0]/P0001 ,
		_w10106_,
		_w10107_
	);
	LUT2 #(
		.INIT('h4)
	) name9576 (
		\sa01_reg[3]/P0001 ,
		_w8221_,
		_w10108_
	);
	LUT2 #(
		.INIT('h8)
	) name9577 (
		\sa01_reg[3]/P0001 ,
		_w10086_,
		_w10109_
	);
	LUT2 #(
		.INIT('h1)
	) name9578 (
		_w9201_,
		_w10108_,
		_w10110_
	);
	LUT2 #(
		.INIT('h4)
	) name9579 (
		_w10109_,
		_w10110_,
		_w10111_
	);
	LUT2 #(
		.INIT('h1)
	) name9580 (
		\sa01_reg[2]/P0001 ,
		_w10111_,
		_w10112_
	);
	LUT2 #(
		.INIT('h2)
	) name9581 (
		\sa01_reg[1]/P0001 ,
		_w9179_,
		_w10113_
	);
	LUT2 #(
		.INIT('h8)
	) name9582 (
		_w9232_,
		_w10113_,
		_w10114_
	);
	LUT2 #(
		.INIT('h4)
	) name9583 (
		_w10112_,
		_w10114_,
		_w10115_
	);
	LUT2 #(
		.INIT('h8)
	) name9584 (
		_w8238_,
		_w9206_,
		_w10116_
	);
	LUT2 #(
		.INIT('h1)
	) name9585 (
		_w9324_,
		_w9368_,
		_w10117_
	);
	LUT2 #(
		.INIT('h1)
	) name9586 (
		\sa01_reg[2]/P0001 ,
		_w10117_,
		_w10118_
	);
	LUT2 #(
		.INIT('h1)
	) name9587 (
		\sa01_reg[1]/P0001 ,
		_w8355_,
		_w10119_
	);
	LUT2 #(
		.INIT('h4)
	) name9588 (
		_w10116_,
		_w10119_,
		_w10120_
	);
	LUT2 #(
		.INIT('h4)
	) name9589 (
		_w10118_,
		_w10120_,
		_w10121_
	);
	LUT2 #(
		.INIT('h1)
	) name9590 (
		_w10115_,
		_w10121_,
		_w10122_
	);
	LUT2 #(
		.INIT('h4)
	) name9591 (
		\sa01_reg[3]/P0001 ,
		_w8258_,
		_w10123_
	);
	LUT2 #(
		.INIT('h1)
	) name9592 (
		_w9215_,
		_w10123_,
		_w10124_
	);
	LUT2 #(
		.INIT('h2)
	) name9593 (
		_w9388_,
		_w10124_,
		_w10125_
	);
	LUT2 #(
		.INIT('h1)
	) name9594 (
		_w8355_,
		_w9237_,
		_w10126_
	);
	LUT2 #(
		.INIT('h1)
	) name9595 (
		\sa01_reg[2]/P0001 ,
		_w10126_,
		_w10127_
	);
	LUT2 #(
		.INIT('h1)
	) name9596 (
		_w8269_,
		_w8293_,
		_w10128_
	);
	LUT2 #(
		.INIT('h2)
	) name9597 (
		_w9318_,
		_w10128_,
		_w10129_
	);
	LUT2 #(
		.INIT('h1)
	) name9598 (
		_w8216_,
		_w8265_,
		_w10130_
	);
	LUT2 #(
		.INIT('h2)
	) name9599 (
		_w9197_,
		_w10130_,
		_w10131_
	);
	LUT2 #(
		.INIT('h1)
	) name9600 (
		_w8362_,
		_w9277_,
		_w10132_
	);
	LUT2 #(
		.INIT('h4)
	) name9601 (
		_w10131_,
		_w10132_,
		_w10133_
	);
	LUT2 #(
		.INIT('h1)
	) name9602 (
		_w10125_,
		_w10127_,
		_w10134_
	);
	LUT2 #(
		.INIT('h4)
	) name9603 (
		_w10129_,
		_w10134_,
		_w10135_
	);
	LUT2 #(
		.INIT('h8)
	) name9604 (
		_w10133_,
		_w10135_,
		_w10136_
	);
	LUT2 #(
		.INIT('h4)
	) name9605 (
		_w10122_,
		_w10136_,
		_w10137_
	);
	LUT2 #(
		.INIT('h1)
	) name9606 (
		\sa01_reg[0]/P0001 ,
		_w10137_,
		_w10138_
	);
	LUT2 #(
		.INIT('h1)
	) name9607 (
		_w9184_,
		_w9219_,
		_w10139_
	);
	LUT2 #(
		.INIT('h1)
	) name9608 (
		_w8224_,
		_w10139_,
		_w10140_
	);
	LUT2 #(
		.INIT('h1)
	) name9609 (
		_w9179_,
		_w9309_,
		_w10141_
	);
	LUT2 #(
		.INIT('h4)
	) name9610 (
		_w10140_,
		_w10141_,
		_w10142_
	);
	LUT2 #(
		.INIT('h2)
	) name9611 (
		_w9382_,
		_w10142_,
		_w10143_
	);
	LUT2 #(
		.INIT('h8)
	) name9612 (
		_w8303_,
		_w9375_,
		_w10144_
	);
	LUT2 #(
		.INIT('h1)
	) name9613 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[2]/P0001 ,
		_w10145_
	);
	LUT2 #(
		.INIT('h1)
	) name9614 (
		_w9315_,
		_w9741_,
		_w10146_
	);
	LUT2 #(
		.INIT('h4)
	) name9615 (
		_w8217_,
		_w10146_,
		_w10147_
	);
	LUT2 #(
		.INIT('h2)
	) name9616 (
		_w10145_,
		_w10147_,
		_w10148_
	);
	LUT2 #(
		.INIT('h1)
	) name9617 (
		_w8295_,
		_w9212_,
		_w10149_
	);
	LUT2 #(
		.INIT('h2)
	) name9618 (
		\sa01_reg[3]/P0001 ,
		_w10149_,
		_w10150_
	);
	LUT2 #(
		.INIT('h1)
	) name9619 (
		_w9338_,
		_w10150_,
		_w10151_
	);
	LUT2 #(
		.INIT('h2)
	) name9620 (
		_w9388_,
		_w10151_,
		_w10152_
	);
	LUT2 #(
		.INIT('h8)
	) name9621 (
		_w8221_,
		_w8351_,
		_w10153_
	);
	LUT2 #(
		.INIT('h1)
	) name9622 (
		_w8362_,
		_w10153_,
		_w10154_
	);
	LUT2 #(
		.INIT('h4)
	) name9623 (
		_w9243_,
		_w10154_,
		_w10155_
	);
	LUT2 #(
		.INIT('h2)
	) name9624 (
		\sa01_reg[2]/P0001 ,
		_w10155_,
		_w10156_
	);
	LUT2 #(
		.INIT('h8)
	) name9625 (
		_w8239_,
		_w8254_,
		_w10157_
	);
	LUT2 #(
		.INIT('h1)
	) name9626 (
		_w9236_,
		_w10157_,
		_w10158_
	);
	LUT2 #(
		.INIT('h4)
	) name9627 (
		_w10156_,
		_w10158_,
		_w10159_
	);
	LUT2 #(
		.INIT('h1)
	) name9628 (
		\sa01_reg[1]/P0001 ,
		_w10159_,
		_w10160_
	);
	LUT2 #(
		.INIT('h1)
	) name9629 (
		_w9757_,
		_w10144_,
		_w10161_
	);
	LUT2 #(
		.INIT('h4)
	) name9630 (
		_w10148_,
		_w10161_,
		_w10162_
	);
	LUT2 #(
		.INIT('h4)
	) name9631 (
		_w10143_,
		_w10162_,
		_w10163_
	);
	LUT2 #(
		.INIT('h4)
	) name9632 (
		_w10152_,
		_w10163_,
		_w10164_
	);
	LUT2 #(
		.INIT('h4)
	) name9633 (
		_w10160_,
		_w10164_,
		_w10165_
	);
	LUT2 #(
		.INIT('h4)
	) name9634 (
		_w10107_,
		_w10165_,
		_w10166_
	);
	LUT2 #(
		.INIT('h4)
	) name9635 (
		_w10138_,
		_w10166_,
		_w10167_
	);
	LUT2 #(
		.INIT('h1)
	) name9636 (
		_w10081_,
		_w10167_,
		_w10168_
	);
	LUT2 #(
		.INIT('h8)
	) name9637 (
		_w10081_,
		_w10167_,
		_w10169_
	);
	LUT2 #(
		.INIT('h1)
	) name9638 (
		_w10168_,
		_w10169_,
		_w10170_
	);
	LUT2 #(
		.INIT('h1)
	) name9639 (
		_w8216_,
		_w8257_,
		_w10171_
	);
	LUT2 #(
		.INIT('h1)
	) name9640 (
		\sa01_reg[2]/P0001 ,
		_w10171_,
		_w10172_
	);
	LUT2 #(
		.INIT('h1)
	) name9641 (
		_w9368_,
		_w10172_,
		_w10173_
	);
	LUT2 #(
		.INIT('h2)
	) name9642 (
		\sa01_reg[1]/P0001 ,
		_w10173_,
		_w10174_
	);
	LUT2 #(
		.INIT('h1)
	) name9643 (
		_w8265_,
		_w8310_,
		_w10175_
	);
	LUT2 #(
		.INIT('h2)
	) name9644 (
		_w9386_,
		_w10175_,
		_w10176_
	);
	LUT2 #(
		.INIT('h1)
	) name9645 (
		_w9356_,
		_w9754_,
		_w10177_
	);
	LUT2 #(
		.INIT('h1)
	) name9646 (
		\sa01_reg[2]/P0001 ,
		_w10177_,
		_w10178_
	);
	LUT2 #(
		.INIT('h1)
	) name9647 (
		_w8283_,
		_w9237_,
		_w10179_
	);
	LUT2 #(
		.INIT('h8)
	) name9648 (
		_w9316_,
		_w10179_,
		_w10180_
	);
	LUT2 #(
		.INIT('h2)
	) name9649 (
		\sa01_reg[2]/P0001 ,
		_w10180_,
		_w10181_
	);
	LUT2 #(
		.INIT('h8)
	) name9650 (
		_w9209_,
		_w10153_,
		_w10182_
	);
	LUT2 #(
		.INIT('h2)
	) name9651 (
		\sa01_reg[5]/P0001 ,
		_w8221_,
		_w10183_
	);
	LUT2 #(
		.INIT('h2)
	) name9652 (
		_w8218_,
		_w10183_,
		_w10184_
	);
	LUT2 #(
		.INIT('h8)
	) name9653 (
		_w8267_,
		_w8342_,
		_w10185_
	);
	LUT2 #(
		.INIT('h8)
	) name9654 (
		_w8215_,
		_w8351_,
		_w10186_
	);
	LUT2 #(
		.INIT('h1)
	) name9655 (
		_w9176_,
		_w10186_,
		_w10187_
	);
	LUT2 #(
		.INIT('h4)
	) name9656 (
		_w9268_,
		_w10187_,
		_w10188_
	);
	LUT2 #(
		.INIT('h2)
	) name9657 (
		\sa01_reg[2]/P0001 ,
		_w10188_,
		_w10189_
	);
	LUT2 #(
		.INIT('h1)
	) name9658 (
		_w10182_,
		_w10185_,
		_w10190_
	);
	LUT2 #(
		.INIT('h4)
	) name9659 (
		_w10184_,
		_w10190_,
		_w10191_
	);
	LUT2 #(
		.INIT('h4)
	) name9660 (
		_w10189_,
		_w10191_,
		_w10192_
	);
	LUT2 #(
		.INIT('h1)
	) name9661 (
		\sa01_reg[1]/P0001 ,
		_w10192_,
		_w10193_
	);
	LUT2 #(
		.INIT('h1)
	) name9662 (
		_w8293_,
		_w8333_,
		_w10194_
	);
	LUT2 #(
		.INIT('h4)
	) name9663 (
		_w10176_,
		_w10194_,
		_w10195_
	);
	LUT2 #(
		.INIT('h4)
	) name9664 (
		_w10178_,
		_w10195_,
		_w10196_
	);
	LUT2 #(
		.INIT('h4)
	) name9665 (
		_w10174_,
		_w10196_,
		_w10197_
	);
	LUT2 #(
		.INIT('h4)
	) name9666 (
		_w10181_,
		_w10197_,
		_w10198_
	);
	LUT2 #(
		.INIT('h4)
	) name9667 (
		_w10193_,
		_w10198_,
		_w10199_
	);
	LUT2 #(
		.INIT('h2)
	) name9668 (
		\sa01_reg[0]/P0001 ,
		_w10199_,
		_w10200_
	);
	LUT2 #(
		.INIT('h8)
	) name9669 (
		_w8222_,
		_w8293_,
		_w10201_
	);
	LUT2 #(
		.INIT('h8)
	) name9670 (
		\sa01_reg[6]/NET0131 ,
		_w9173_,
		_w10202_
	);
	LUT2 #(
		.INIT('h1)
	) name9671 (
		_w9237_,
		_w10202_,
		_w10203_
	);
	LUT2 #(
		.INIT('h4)
	) name9672 (
		_w9361_,
		_w10203_,
		_w10204_
	);
	LUT2 #(
		.INIT('h1)
	) name9673 (
		\sa01_reg[2]/P0001 ,
		_w10204_,
		_w10205_
	);
	LUT2 #(
		.INIT('h1)
	) name9674 (
		_w8219_,
		_w8310_,
		_w10206_
	);
	LUT2 #(
		.INIT('h2)
	) name9675 (
		_w9698_,
		_w10206_,
		_w10207_
	);
	LUT2 #(
		.INIT('h2)
	) name9676 (
		_w8245_,
		_w8264_,
		_w10208_
	);
	LUT2 #(
		.INIT('h8)
	) name9677 (
		_w9318_,
		_w10208_,
		_w10209_
	);
	LUT2 #(
		.INIT('h1)
	) name9678 (
		\sa01_reg[3]/P0001 ,
		_w9728_,
		_w10210_
	);
	LUT2 #(
		.INIT('h1)
	) name9679 (
		_w8241_,
		_w10210_,
		_w10211_
	);
	LUT2 #(
		.INIT('h1)
	) name9680 (
		\sa01_reg[1]/P0001 ,
		_w10211_,
		_w10212_
	);
	LUT2 #(
		.INIT('h8)
	) name9681 (
		_w8254_,
		_w9694_,
		_w10213_
	);
	LUT2 #(
		.INIT('h2)
	) name9682 (
		_w8215_,
		_w8238_,
		_w10214_
	);
	LUT2 #(
		.INIT('h8)
	) name9683 (
		_w8235_,
		_w8238_,
		_w10215_
	);
	LUT2 #(
		.INIT('h8)
	) name9684 (
		_w8277_,
		_w8329_,
		_w10216_
	);
	LUT2 #(
		.INIT('h1)
	) name9685 (
		_w10213_,
		_w10214_,
		_w10217_
	);
	LUT2 #(
		.INIT('h4)
	) name9686 (
		_w10215_,
		_w10217_,
		_w10218_
	);
	LUT2 #(
		.INIT('h4)
	) name9687 (
		_w10216_,
		_w10218_,
		_w10219_
	);
	LUT2 #(
		.INIT('h2)
	) name9688 (
		\sa01_reg[1]/P0001 ,
		_w10219_,
		_w10220_
	);
	LUT2 #(
		.INIT('h1)
	) name9689 (
		_w10207_,
		_w10209_,
		_w10221_
	);
	LUT2 #(
		.INIT('h4)
	) name9690 (
		_w10205_,
		_w10221_,
		_w10222_
	);
	LUT2 #(
		.INIT('h1)
	) name9691 (
		_w10212_,
		_w10220_,
		_w10223_
	);
	LUT2 #(
		.INIT('h8)
	) name9692 (
		_w10222_,
		_w10223_,
		_w10224_
	);
	LUT2 #(
		.INIT('h1)
	) name9693 (
		\sa01_reg[0]/P0001 ,
		_w10224_,
		_w10225_
	);
	LUT2 #(
		.INIT('h4)
	) name9694 (
		_w8308_,
		_w8326_,
		_w10226_
	);
	LUT2 #(
		.INIT('h1)
	) name9695 (
		_w8363_,
		_w10226_,
		_w10227_
	);
	LUT2 #(
		.INIT('h1)
	) name9696 (
		\sa01_reg[2]/P0001 ,
		_w10227_,
		_w10228_
	);
	LUT2 #(
		.INIT('h4)
	) name9697 (
		\sa01_reg[2]/P0001 ,
		_w9256_,
		_w10229_
	);
	LUT2 #(
		.INIT('h8)
	) name9698 (
		\sa01_reg[2]/P0001 ,
		_w8267_,
		_w10230_
	);
	LUT2 #(
		.INIT('h1)
	) name9699 (
		_w8257_,
		_w8344_,
		_w10231_
	);
	LUT2 #(
		.INIT('h2)
	) name9700 (
		_w10230_,
		_w10231_,
		_w10232_
	);
	LUT2 #(
		.INIT('h1)
	) name9701 (
		_w9277_,
		_w10229_,
		_w10233_
	);
	LUT2 #(
		.INIT('h4)
	) name9702 (
		_w10232_,
		_w10233_,
		_w10234_
	);
	LUT2 #(
		.INIT('h4)
	) name9703 (
		_w10228_,
		_w10234_,
		_w10235_
	);
	LUT2 #(
		.INIT('h1)
	) name9704 (
		\sa01_reg[1]/P0001 ,
		_w10235_,
		_w10236_
	);
	LUT2 #(
		.INIT('h8)
	) name9705 (
		\sa01_reg[1]/P0001 ,
		_w9774_,
		_w10237_
	);
	LUT2 #(
		.INIT('h1)
	) name9706 (
		_w10215_,
		_w10237_,
		_w10238_
	);
	LUT2 #(
		.INIT('h1)
	) name9707 (
		\sa01_reg[2]/P0001 ,
		_w10238_,
		_w10239_
	);
	LUT2 #(
		.INIT('h1)
	) name9708 (
		_w8220_,
		_w8268_,
		_w10240_
	);
	LUT2 #(
		.INIT('h1)
	) name9709 (
		_w9207_,
		_w9322_,
		_w10241_
	);
	LUT2 #(
		.INIT('h8)
	) name9710 (
		_w10240_,
		_w10241_,
		_w10242_
	);
	LUT2 #(
		.INIT('h2)
	) name9711 (
		\sa01_reg[1]/P0001 ,
		_w10242_,
		_w10243_
	);
	LUT2 #(
		.INIT('h1)
	) name9712 (
		_w10201_,
		_w10239_,
		_w10244_
	);
	LUT2 #(
		.INIT('h4)
	) name9713 (
		_w10243_,
		_w10244_,
		_w10245_
	);
	LUT2 #(
		.INIT('h4)
	) name9714 (
		_w10236_,
		_w10245_,
		_w10246_
	);
	LUT2 #(
		.INIT('h4)
	) name9715 (
		_w10225_,
		_w10246_,
		_w10247_
	);
	LUT2 #(
		.INIT('h4)
	) name9716 (
		_w10200_,
		_w10247_,
		_w10248_
	);
	LUT2 #(
		.INIT('h1)
	) name9717 (
		_w9783_,
		_w10248_,
		_w10249_
	);
	LUT2 #(
		.INIT('h8)
	) name9718 (
		_w9783_,
		_w10248_,
		_w10250_
	);
	LUT2 #(
		.INIT('h1)
	) name9719 (
		_w10249_,
		_w10250_,
		_w10251_
	);
	LUT2 #(
		.INIT('h2)
	) name9720 (
		_w10170_,
		_w10251_,
		_w10252_
	);
	LUT2 #(
		.INIT('h4)
	) name9721 (
		_w10170_,
		_w10251_,
		_w10253_
	);
	LUT2 #(
		.INIT('h1)
	) name9722 (
		_w10252_,
		_w10253_,
		_w10254_
	);
	LUT2 #(
		.INIT('h4)
	) name9723 (
		\sa30_reg[3]/P0001 ,
		_w8682_,
		_w10255_
	);
	LUT2 #(
		.INIT('h4)
	) name9724 (
		\sa30_reg[5]/P0001 ,
		_w10255_,
		_w10256_
	);
	LUT2 #(
		.INIT('h8)
	) name9725 (
		_w8741_,
		_w10256_,
		_w10257_
	);
	LUT2 #(
		.INIT('h1)
	) name9726 (
		_w8706_,
		_w8823_,
		_w10258_
	);
	LUT2 #(
		.INIT('h4)
	) name9727 (
		_w8951_,
		_w10258_,
		_w10259_
	);
	LUT2 #(
		.INIT('h2)
	) name9728 (
		\sa30_reg[2]/P0001 ,
		_w10259_,
		_w10260_
	);
	LUT2 #(
		.INIT('h2)
	) name9729 (
		\sa30_reg[5]/P0001 ,
		_w8682_,
		_w10261_
	);
	LUT2 #(
		.INIT('h2)
	) name9730 (
		_w8725_,
		_w10261_,
		_w10262_
	);
	LUT2 #(
		.INIT('h8)
	) name9731 (
		_w8698_,
		_w8756_,
		_w10263_
	);
	LUT2 #(
		.INIT('h1)
	) name9732 (
		_w10262_,
		_w10263_,
		_w10264_
	);
	LUT2 #(
		.INIT('h4)
	) name9733 (
		_w10257_,
		_w10264_,
		_w10265_
	);
	LUT2 #(
		.INIT('h4)
	) name9734 (
		_w10260_,
		_w10265_,
		_w10266_
	);
	LUT2 #(
		.INIT('h1)
	) name9735 (
		\sa30_reg[1]/P0001 ,
		_w10266_,
		_w10267_
	);
	LUT2 #(
		.INIT('h1)
	) name9736 (
		_w8697_,
		_w8950_,
		_w10268_
	);
	LUT2 #(
		.INIT('h1)
	) name9737 (
		\sa30_reg[2]/P0001 ,
		_w10268_,
		_w10269_
	);
	LUT2 #(
		.INIT('h1)
	) name9738 (
		_w8961_,
		_w10269_,
		_w10270_
	);
	LUT2 #(
		.INIT('h2)
	) name9739 (
		\sa30_reg[1]/P0001 ,
		_w10270_,
		_w10271_
	);
	LUT2 #(
		.INIT('h8)
	) name9740 (
		\sa30_reg[3]/P0001 ,
		_w8792_,
		_w10272_
	);
	LUT2 #(
		.INIT('h1)
	) name9741 (
		_w8838_,
		_w10272_,
		_w10273_
	);
	LUT2 #(
		.INIT('h1)
	) name9742 (
		\sa30_reg[2]/P0001 ,
		_w10273_,
		_w10274_
	);
	LUT2 #(
		.INIT('h8)
	) name9743 (
		\sa30_reg[6]/NET0131 ,
		_w8930_,
		_w10275_
	);
	LUT2 #(
		.INIT('h8)
	) name9744 (
		_w8721_,
		_w8756_,
		_w10276_
	);
	LUT2 #(
		.INIT('h1)
	) name9745 (
		_w10275_,
		_w10276_,
		_w10277_
	);
	LUT2 #(
		.INIT('h1)
	) name9746 (
		\sa30_reg[2]/P0001 ,
		_w10277_,
		_w10278_
	);
	LUT2 #(
		.INIT('h8)
	) name9747 (
		\sa30_reg[5]/P0001 ,
		_w8835_,
		_w10279_
	);
	LUT2 #(
		.INIT('h1)
	) name9748 (
		_w8786_,
		_w9543_,
		_w10280_
	);
	LUT2 #(
		.INIT('h8)
	) name9749 (
		_w8870_,
		_w10280_,
		_w10281_
	);
	LUT2 #(
		.INIT('h2)
	) name9750 (
		\sa30_reg[2]/P0001 ,
		_w10281_,
		_w10282_
	);
	LUT2 #(
		.INIT('h1)
	) name9751 (
		_w9608_,
		_w10279_,
		_w10283_
	);
	LUT2 #(
		.INIT('h4)
	) name9752 (
		_w10274_,
		_w10283_,
		_w10284_
	);
	LUT2 #(
		.INIT('h4)
	) name9753 (
		_w10278_,
		_w10284_,
		_w10285_
	);
	LUT2 #(
		.INIT('h4)
	) name9754 (
		_w10271_,
		_w10285_,
		_w10286_
	);
	LUT2 #(
		.INIT('h4)
	) name9755 (
		_w10282_,
		_w10286_,
		_w10287_
	);
	LUT2 #(
		.INIT('h4)
	) name9756 (
		_w10267_,
		_w10287_,
		_w10288_
	);
	LUT2 #(
		.INIT('h2)
	) name9757 (
		\sa30_reg[0]/P0002 ,
		_w10288_,
		_w10289_
	);
	LUT2 #(
		.INIT('h8)
	) name9758 (
		\sa30_reg[6]/NET0131 ,
		_w8704_,
		_w10290_
	);
	LUT2 #(
		.INIT('h1)
	) name9759 (
		_w8786_,
		_w10290_,
		_w10291_
	);
	LUT2 #(
		.INIT('h4)
	) name9760 (
		_w8916_,
		_w10291_,
		_w10292_
	);
	LUT2 #(
		.INIT('h1)
	) name9761 (
		\sa30_reg[2]/P0001 ,
		_w10292_,
		_w10293_
	);
	LUT2 #(
		.INIT('h4)
	) name9762 (
		\sa30_reg[1]/P0001 ,
		\sa30_reg[2]/P0001 ,
		_w10294_
	);
	LUT2 #(
		.INIT('h2)
	) name9763 (
		_w8694_,
		_w8758_,
		_w10295_
	);
	LUT2 #(
		.INIT('h8)
	) name9764 (
		_w10294_,
		_w10295_,
		_w10296_
	);
	LUT2 #(
		.INIT('h8)
	) name9765 (
		\sa30_reg[3]/P0001 ,
		_w9575_,
		_w10297_
	);
	LUT2 #(
		.INIT('h1)
	) name9766 (
		_w8792_,
		_w8845_,
		_w10298_
	);
	LUT2 #(
		.INIT('h2)
	) name9767 (
		_w10297_,
		_w10298_,
		_w10299_
	);
	LUT2 #(
		.INIT('h1)
	) name9768 (
		_w8767_,
		_w8952_,
		_w10300_
	);
	LUT2 #(
		.INIT('h1)
	) name9769 (
		\sa30_reg[3]/P0001 ,
		_w10300_,
		_w10301_
	);
	LUT2 #(
		.INIT('h1)
	) name9770 (
		_w9581_,
		_w10301_,
		_w10302_
	);
	LUT2 #(
		.INIT('h1)
	) name9771 (
		\sa30_reg[1]/P0001 ,
		_w10302_,
		_w10303_
	);
	LUT2 #(
		.INIT('h8)
	) name9772 (
		_w8705_,
		_w8844_,
		_w10304_
	);
	LUT2 #(
		.INIT('h8)
	) name9773 (
		_w8833_,
		_w8874_,
		_w10305_
	);
	LUT2 #(
		.INIT('h1)
	) name9774 (
		_w8724_,
		_w8733_,
		_w10306_
	);
	LUT2 #(
		.INIT('h1)
	) name9775 (
		_w9603_,
		_w10305_,
		_w10307_
	);
	LUT2 #(
		.INIT('h8)
	) name9776 (
		_w10306_,
		_w10307_,
		_w10308_
	);
	LUT2 #(
		.INIT('h4)
	) name9777 (
		_w10304_,
		_w10308_,
		_w10309_
	);
	LUT2 #(
		.INIT('h2)
	) name9778 (
		\sa30_reg[1]/P0001 ,
		_w10309_,
		_w10310_
	);
	LUT2 #(
		.INIT('h1)
	) name9779 (
		_w10296_,
		_w10299_,
		_w10311_
	);
	LUT2 #(
		.INIT('h4)
	) name9780 (
		_w10293_,
		_w10311_,
		_w10312_
	);
	LUT2 #(
		.INIT('h1)
	) name9781 (
		_w10303_,
		_w10310_,
		_w10313_
	);
	LUT2 #(
		.INIT('h8)
	) name9782 (
		_w10312_,
		_w10313_,
		_w10314_
	);
	LUT2 #(
		.INIT('h1)
	) name9783 (
		\sa30_reg[0]/P0002 ,
		_w10314_,
		_w10315_
	);
	LUT2 #(
		.INIT('h1)
	) name9784 (
		\sa30_reg[2]/P0001 ,
		_w8785_,
		_w10316_
	);
	LUT2 #(
		.INIT('h1)
	) name9785 (
		_w9592_,
		_w10316_,
		_w10317_
	);
	LUT2 #(
		.INIT('h8)
	) name9786 (
		_w8929_,
		_w9614_,
		_w10318_
	);
	LUT2 #(
		.INIT('h1)
	) name9787 (
		_w8916_,
		_w9620_,
		_w10319_
	);
	LUT2 #(
		.INIT('h4)
	) name9788 (
		_w10318_,
		_w10319_,
		_w10320_
	);
	LUT2 #(
		.INIT('h1)
	) name9789 (
		\sa30_reg[7]/P0001 ,
		_w10320_,
		_w10321_
	);
	LUT2 #(
		.INIT('h1)
	) name9790 (
		_w10317_,
		_w10321_,
		_w10322_
	);
	LUT2 #(
		.INIT('h2)
	) name9791 (
		\sa30_reg[1]/P0001 ,
		_w10322_,
		_w10323_
	);
	LUT2 #(
		.INIT('h4)
	) name9792 (
		\sa30_reg[2]/P0001 ,
		_w9603_,
		_w10324_
	);
	LUT2 #(
		.INIT('h8)
	) name9793 (
		_w9575_,
		_w10279_,
		_w10325_
	);
	LUT2 #(
		.INIT('h1)
	) name9794 (
		_w8735_,
		_w9565_,
		_w10326_
	);
	LUT2 #(
		.INIT('h1)
	) name9795 (
		\sa30_reg[7]/P0001 ,
		_w10326_,
		_w10327_
	);
	LUT2 #(
		.INIT('h4)
	) name9796 (
		\sa30_reg[3]/P0001 ,
		_w8814_,
		_w10328_
	);
	LUT2 #(
		.INIT('h1)
	) name9797 (
		_w10327_,
		_w10328_,
		_w10329_
	);
	LUT2 #(
		.INIT('h1)
	) name9798 (
		\sa30_reg[2]/P0001 ,
		_w10329_,
		_w10330_
	);
	LUT2 #(
		.INIT('h4)
	) name9799 (
		\sa30_reg[2]/P0001 ,
		_w8705_,
		_w10331_
	);
	LUT2 #(
		.INIT('h8)
	) name9800 (
		_w8725_,
		_w10331_,
		_w10332_
	);
	LUT2 #(
		.INIT('h8)
	) name9801 (
		\sa30_reg[7]/P0001 ,
		_w8916_,
		_w10333_
	);
	LUT2 #(
		.INIT('h1)
	) name9802 (
		_w8699_,
		_w10333_,
		_w10334_
	);
	LUT2 #(
		.INIT('h2)
	) name9803 (
		\sa30_reg[2]/P0001 ,
		_w10334_,
		_w10335_
	);
	LUT2 #(
		.INIT('h1)
	) name9804 (
		_w8847_,
		_w10332_,
		_w10336_
	);
	LUT2 #(
		.INIT('h4)
	) name9805 (
		_w10335_,
		_w10336_,
		_w10337_
	);
	LUT2 #(
		.INIT('h4)
	) name9806 (
		_w10330_,
		_w10337_,
		_w10338_
	);
	LUT2 #(
		.INIT('h1)
	) name9807 (
		\sa30_reg[1]/P0001 ,
		_w10338_,
		_w10339_
	);
	LUT2 #(
		.INIT('h1)
	) name9808 (
		_w10324_,
		_w10325_,
		_w10340_
	);
	LUT2 #(
		.INIT('h4)
	) name9809 (
		_w10323_,
		_w10340_,
		_w10341_
	);
	LUT2 #(
		.INIT('h4)
	) name9810 (
		_w10339_,
		_w10341_,
		_w10342_
	);
	LUT2 #(
		.INIT('h4)
	) name9811 (
		_w10315_,
		_w10342_,
		_w10343_
	);
	LUT2 #(
		.INIT('h4)
	) name9812 (
		_w10289_,
		_w10343_,
		_w10344_
	);
	LUT2 #(
		.INIT('h1)
	) name9813 (
		_w8773_,
		_w9582_,
		_w10345_
	);
	LUT2 #(
		.INIT('h2)
	) name9814 (
		\sa30_reg[7]/P0001 ,
		_w10345_,
		_w10346_
	);
	LUT2 #(
		.INIT('h8)
	) name9815 (
		_w8844_,
		_w9547_,
		_w10347_
	);
	LUT2 #(
		.INIT('h1)
	) name9816 (
		_w9553_,
		_w10347_,
		_w10348_
	);
	LUT2 #(
		.INIT('h4)
	) name9817 (
		_w10346_,
		_w10348_,
		_w10349_
	);
	LUT2 #(
		.INIT('h1)
	) name9818 (
		\sa30_reg[1]/P0001 ,
		_w10349_,
		_w10350_
	);
	LUT2 #(
		.INIT('h8)
	) name9819 (
		\sa30_reg[4]/P0001 ,
		_w8845_,
		_w10351_
	);
	LUT2 #(
		.INIT('h1)
	) name9820 (
		_w8749_,
		_w10275_,
		_w10352_
	);
	LUT2 #(
		.INIT('h4)
	) name9821 (
		_w10351_,
		_w10352_,
		_w10353_
	);
	LUT2 #(
		.INIT('h2)
	) name9822 (
		_w8844_,
		_w10353_,
		_w10354_
	);
	LUT2 #(
		.INIT('h4)
	) name9823 (
		\sa30_reg[3]/P0001 ,
		_w8816_,
		_w10355_
	);
	LUT2 #(
		.INIT('h1)
	) name9824 (
		_w10263_,
		_w10355_,
		_w10356_
	);
	LUT2 #(
		.INIT('h4)
	) name9825 (
		\sa30_reg[6]/NET0131 ,
		_w8774_,
		_w10357_
	);
	LUT2 #(
		.INIT('h1)
	) name9826 (
		_w8822_,
		_w10357_,
		_w10358_
	);
	LUT2 #(
		.INIT('h8)
	) name9827 (
		_w10356_,
		_w10358_,
		_w10359_
	);
	LUT2 #(
		.INIT('h1)
	) name9828 (
		\sa30_reg[2]/P0001 ,
		_w10359_,
		_w10360_
	);
	LUT2 #(
		.INIT('h1)
	) name9829 (
		_w9560_,
		_w9632_,
		_w10361_
	);
	LUT2 #(
		.INIT('h1)
	) name9830 (
		\sa30_reg[2]/P0001 ,
		_w10361_,
		_w10362_
	);
	LUT2 #(
		.INIT('h8)
	) name9831 (
		\sa30_reg[3]/P0001 ,
		_w8692_,
		_w10363_
	);
	LUT2 #(
		.INIT('h1)
	) name9832 (
		_w8915_,
		_w10318_,
		_w10364_
	);
	LUT2 #(
		.INIT('h4)
	) name9833 (
		_w10363_,
		_w10364_,
		_w10365_
	);
	LUT2 #(
		.INIT('h4)
	) name9834 (
		_w10362_,
		_w10365_,
		_w10366_
	);
	LUT2 #(
		.INIT('h2)
	) name9835 (
		\sa30_reg[1]/P0001 ,
		_w10366_,
		_w10367_
	);
	LUT2 #(
		.INIT('h1)
	) name9836 (
		_w10350_,
		_w10354_,
		_w10368_
	);
	LUT2 #(
		.INIT('h4)
	) name9837 (
		_w10360_,
		_w10368_,
		_w10369_
	);
	LUT2 #(
		.INIT('h4)
	) name9838 (
		_w10367_,
		_w10369_,
		_w10370_
	);
	LUT2 #(
		.INIT('h1)
	) name9839 (
		\sa30_reg[0]/P0002 ,
		_w10370_,
		_w10371_
	);
	LUT2 #(
		.INIT('h4)
	) name9840 (
		_w8684_,
		_w8741_,
		_w10372_
	);
	LUT2 #(
		.INIT('h4)
	) name9841 (
		_w8710_,
		_w10372_,
		_w10373_
	);
	LUT2 #(
		.INIT('h2)
	) name9842 (
		_w8835_,
		_w9575_,
		_w10374_
	);
	LUT2 #(
		.INIT('h4)
	) name9843 (
		\sa30_reg[4]/P0001 ,
		_w8874_,
		_w10375_
	);
	LUT2 #(
		.INIT('h8)
	) name9844 (
		_w8929_,
		_w10375_,
		_w10376_
	);
	LUT2 #(
		.INIT('h1)
	) name9845 (
		_w9620_,
		_w10331_,
		_w10377_
	);
	LUT2 #(
		.INIT('h1)
	) name9846 (
		_w10373_,
		_w10374_,
		_w10378_
	);
	LUT2 #(
		.INIT('h4)
	) name9847 (
		_w10376_,
		_w10378_,
		_w10379_
	);
	LUT2 #(
		.INIT('h8)
	) name9848 (
		_w10377_,
		_w10379_,
		_w10380_
	);
	LUT2 #(
		.INIT('h1)
	) name9849 (
		\sa30_reg[1]/P0001 ,
		_w10380_,
		_w10381_
	);
	LUT2 #(
		.INIT('h8)
	) name9850 (
		_w8682_,
		_w8871_,
		_w10382_
	);
	LUT2 #(
		.INIT('h1)
	) name9851 (
		_w9604_,
		_w10382_,
		_w10383_
	);
	LUT2 #(
		.INIT('h2)
	) name9852 (
		\sa30_reg[1]/P0001 ,
		_w10383_,
		_w10384_
	);
	LUT2 #(
		.INIT('h1)
	) name9853 (
		_w8685_,
		_w8743_,
		_w10385_
	);
	LUT2 #(
		.INIT('h1)
	) name9854 (
		\sa30_reg[3]/P0001 ,
		_w10385_,
		_w10386_
	);
	LUT2 #(
		.INIT('h1)
	) name9855 (
		_w8706_,
		_w10386_,
		_w10387_
	);
	LUT2 #(
		.INIT('h2)
	) name9856 (
		\sa30_reg[2]/P0001 ,
		_w10387_,
		_w10388_
	);
	LUT2 #(
		.INIT('h8)
	) name9857 (
		\sa30_reg[4]/P0001 ,
		_w8775_,
		_w10389_
	);
	LUT2 #(
		.INIT('h1)
	) name9858 (
		_w8724_,
		_w8766_,
		_w10390_
	);
	LUT2 #(
		.INIT('h1)
	) name9859 (
		_w8888_,
		_w10389_,
		_w10391_
	);
	LUT2 #(
		.INIT('h8)
	) name9860 (
		_w10390_,
		_w10391_,
		_w10392_
	);
	LUT2 #(
		.INIT('h2)
	) name9861 (
		_w8946_,
		_w10392_,
		_w10393_
	);
	LUT2 #(
		.INIT('h8)
	) name9862 (
		_w8792_,
		_w10297_,
		_w10394_
	);
	LUT2 #(
		.INIT('h8)
	) name9863 (
		_w8741_,
		_w8835_,
		_w10395_
	);
	LUT2 #(
		.INIT('h1)
	) name9864 (
		_w10276_,
		_w10394_,
		_w10396_
	);
	LUT2 #(
		.INIT('h4)
	) name9865 (
		_w10395_,
		_w10396_,
		_w10397_
	);
	LUT2 #(
		.INIT('h4)
	) name9866 (
		_w10384_,
		_w10397_,
		_w10398_
	);
	LUT2 #(
		.INIT('h4)
	) name9867 (
		_w10393_,
		_w10398_,
		_w10399_
	);
	LUT2 #(
		.INIT('h4)
	) name9868 (
		_w10388_,
		_w10399_,
		_w10400_
	);
	LUT2 #(
		.INIT('h4)
	) name9869 (
		_w10381_,
		_w10400_,
		_w10401_
	);
	LUT2 #(
		.INIT('h2)
	) name9870 (
		\sa30_reg[0]/P0002 ,
		_w10401_,
		_w10402_
	);
	LUT2 #(
		.INIT('h8)
	) name9871 (
		\sa30_reg[5]/P0001 ,
		_w8735_,
		_w10403_
	);
	LUT2 #(
		.INIT('h1)
	) name9872 (
		_w8703_,
		_w9604_,
		_w10404_
	);
	LUT2 #(
		.INIT('h4)
	) name9873 (
		_w10403_,
		_w10404_,
		_w10405_
	);
	LUT2 #(
		.INIT('h2)
	) name9874 (
		_w10294_,
		_w10405_,
		_w10406_
	);
	LUT2 #(
		.INIT('h1)
	) name9875 (
		_w8685_,
		_w8845_,
		_w10407_
	);
	LUT2 #(
		.INIT('h8)
	) name9876 (
		_w10300_,
		_w10407_,
		_w10408_
	);
	LUT2 #(
		.INIT('h8)
	) name9877 (
		\sa30_reg[1]/P0001 ,
		_w8940_,
		_w10409_
	);
	LUT2 #(
		.INIT('h4)
	) name9878 (
		_w10408_,
		_w10409_,
		_w10410_
	);
	LUT2 #(
		.INIT('h1)
	) name9879 (
		_w8700_,
		_w9561_,
		_w10411_
	);
	LUT2 #(
		.INIT('h1)
	) name9880 (
		\sa30_reg[2]/P0001 ,
		_w10411_,
		_w10412_
	);
	LUT2 #(
		.INIT('h2)
	) name9881 (
		\sa30_reg[2]/P0001 ,
		_w8785_,
		_w10413_
	);
	LUT2 #(
		.INIT('h1)
	) name9882 (
		_w8785_,
		_w8922_,
		_w10414_
	);
	LUT2 #(
		.INIT('h8)
	) name9883 (
		_w10356_,
		_w10414_,
		_w10415_
	);
	LUT2 #(
		.INIT('h1)
	) name9884 (
		\sa30_reg[1]/P0001 ,
		_w10413_,
		_w10416_
	);
	LUT2 #(
		.INIT('h4)
	) name9885 (
		_w10415_,
		_w10416_,
		_w10417_
	);
	LUT2 #(
		.INIT('h4)
	) name9886 (
		\sa30_reg[6]/NET0131 ,
		_w8757_,
		_w10418_
	);
	LUT2 #(
		.INIT('h1)
	) name9887 (
		_w8743_,
		_w9572_,
		_w10419_
	);
	LUT2 #(
		.INIT('h4)
	) name9888 (
		_w10418_,
		_w10419_,
		_w10420_
	);
	LUT2 #(
		.INIT('h1)
	) name9889 (
		\sa30_reg[3]/P0001 ,
		_w10420_,
		_w10421_
	);
	LUT2 #(
		.INIT('h1)
	) name9890 (
		_w8744_,
		_w8759_,
		_w10422_
	);
	LUT2 #(
		.INIT('h4)
	) name9891 (
		_w10421_,
		_w10422_,
		_w10423_
	);
	LUT2 #(
		.INIT('h2)
	) name9892 (
		_w8946_,
		_w10423_,
		_w10424_
	);
	LUT2 #(
		.INIT('h1)
	) name9893 (
		_w10410_,
		_w10412_,
		_w10425_
	);
	LUT2 #(
		.INIT('h4)
	) name9894 (
		_w10406_,
		_w10425_,
		_w10426_
	);
	LUT2 #(
		.INIT('h4)
	) name9895 (
		_w10417_,
		_w10426_,
		_w10427_
	);
	LUT2 #(
		.INIT('h4)
	) name9896 (
		_w10424_,
		_w10427_,
		_w10428_
	);
	LUT2 #(
		.INIT('h4)
	) name9897 (
		_w10371_,
		_w10428_,
		_w10429_
	);
	LUT2 #(
		.INIT('h4)
	) name9898 (
		_w10402_,
		_w10429_,
		_w10430_
	);
	LUT2 #(
		.INIT('h2)
	) name9899 (
		_w10344_,
		_w10430_,
		_w10431_
	);
	LUT2 #(
		.INIT('h4)
	) name9900 (
		_w10344_,
		_w10430_,
		_w10432_
	);
	LUT2 #(
		.INIT('h1)
	) name9901 (
		_w10431_,
		_w10432_,
		_w10433_
	);
	LUT2 #(
		.INIT('h4)
	) name9902 (
		_w8546_,
		_w8667_,
		_w10434_
	);
	LUT2 #(
		.INIT('h8)
	) name9903 (
		_w8509_,
		_w8519_,
		_w10435_
	);
	LUT2 #(
		.INIT('h8)
	) name9904 (
		\sa23_reg[4]/P0001 ,
		_w8618_,
		_w10436_
	);
	LUT2 #(
		.INIT('h2)
	) name9905 (
		_w8512_,
		_w9900_,
		_w10437_
	);
	LUT2 #(
		.INIT('h1)
	) name9906 (
		\sa23_reg[1]/P0001 ,
		_w9964_,
		_w10438_
	);
	LUT2 #(
		.INIT('h4)
	) name9907 (
		_w10435_,
		_w10438_,
		_w10439_
	);
	LUT2 #(
		.INIT('h1)
	) name9908 (
		_w10436_,
		_w10437_,
		_w10440_
	);
	LUT2 #(
		.INIT('h8)
	) name9909 (
		_w10439_,
		_w10440_,
		_w10441_
	);
	LUT2 #(
		.INIT('h8)
	) name9910 (
		_w8521_,
		_w9066_,
		_w10442_
	);
	LUT2 #(
		.INIT('h1)
	) name9911 (
		_w8563_,
		_w10442_,
		_w10443_
	);
	LUT2 #(
		.INIT('h1)
	) name9912 (
		_w9096_,
		_w9151_,
		_w10444_
	);
	LUT2 #(
		.INIT('h4)
	) name9913 (
		_w9453_,
		_w10444_,
		_w10445_
	);
	LUT2 #(
		.INIT('h2)
	) name9914 (
		\sa23_reg[2]/P0001 ,
		_w10445_,
		_w10446_
	);
	LUT2 #(
		.INIT('h8)
	) name9915 (
		\sa23_reg[1]/P0001 ,
		_w10443_,
		_w10447_
	);
	LUT2 #(
		.INIT('h4)
	) name9916 (
		_w10446_,
		_w10447_,
		_w10448_
	);
	LUT2 #(
		.INIT('h1)
	) name9917 (
		_w10441_,
		_w10448_,
		_w10449_
	);
	LUT2 #(
		.INIT('h1)
	) name9918 (
		_w9154_,
		_w9964_,
		_w10450_
	);
	LUT2 #(
		.INIT('h4)
	) name9919 (
		_w9492_,
		_w10450_,
		_w10451_
	);
	LUT2 #(
		.INIT('h1)
	) name9920 (
		\sa23_reg[2]/P0001 ,
		_w10451_,
		_w10452_
	);
	LUT2 #(
		.INIT('h2)
	) name9921 (
		_w8527_,
		_w9427_,
		_w10453_
	);
	LUT2 #(
		.INIT('h2)
	) name9922 (
		\sa23_reg[0]/P0001 ,
		_w10434_,
		_w10454_
	);
	LUT2 #(
		.INIT('h4)
	) name9923 (
		_w10453_,
		_w10454_,
		_w10455_
	);
	LUT2 #(
		.INIT('h4)
	) name9924 (
		_w10452_,
		_w10455_,
		_w10456_
	);
	LUT2 #(
		.INIT('h4)
	) name9925 (
		_w10449_,
		_w10456_,
		_w10457_
	);
	LUT2 #(
		.INIT('h4)
	) name9926 (
		_w9074_,
		_w9153_,
		_w10458_
	);
	LUT2 #(
		.INIT('h2)
	) name9927 (
		\sa23_reg[2]/P0001 ,
		_w9097_,
		_w10459_
	);
	LUT2 #(
		.INIT('h4)
	) name9928 (
		_w9492_,
		_w10459_,
		_w10460_
	);
	LUT2 #(
		.INIT('h1)
	) name9929 (
		_w10458_,
		_w10460_,
		_w10461_
	);
	LUT2 #(
		.INIT('h1)
	) name9930 (
		\sa23_reg[1]/P0001 ,
		_w9130_,
		_w10462_
	);
	LUT2 #(
		.INIT('h4)
	) name9931 (
		_w9476_,
		_w10462_,
		_w10463_
	);
	LUT2 #(
		.INIT('h4)
	) name9932 (
		_w10461_,
		_w10463_,
		_w10464_
	);
	LUT2 #(
		.INIT('h2)
	) name9933 (
		\sa23_reg[1]/P0001 ,
		_w8530_,
		_w10465_
	);
	LUT2 #(
		.INIT('h1)
	) name9934 (
		\sa23_reg[2]/P0001 ,
		_w8548_,
		_w10466_
	);
	LUT2 #(
		.INIT('h1)
	) name9935 (
		_w8550_,
		_w9129_,
		_w10467_
	);
	LUT2 #(
		.INIT('h8)
	) name9936 (
		_w10466_,
		_w10467_,
		_w10468_
	);
	LUT2 #(
		.INIT('h2)
	) name9937 (
		\sa23_reg[2]/P0001 ,
		_w9113_,
		_w10469_
	);
	LUT2 #(
		.INIT('h4)
	) name9938 (
		_w9942_,
		_w10469_,
		_w10470_
	);
	LUT2 #(
		.INIT('h1)
	) name9939 (
		_w10468_,
		_w10470_,
		_w10471_
	);
	LUT2 #(
		.INIT('h8)
	) name9940 (
		_w8592_,
		_w10465_,
		_w10472_
	);
	LUT2 #(
		.INIT('h4)
	) name9941 (
		_w10471_,
		_w10472_,
		_w10473_
	);
	LUT2 #(
		.INIT('h1)
	) name9942 (
		_w10464_,
		_w10473_,
		_w10474_
	);
	LUT2 #(
		.INIT('h2)
	) name9943 (
		\sa23_reg[2]/P0001 ,
		_w8523_,
		_w10475_
	);
	LUT2 #(
		.INIT('h4)
	) name9944 (
		_w9128_,
		_w10475_,
		_w10476_
	);
	LUT2 #(
		.INIT('h1)
	) name9945 (
		\sa23_reg[2]/P0001 ,
		_w8663_,
		_w10477_
	);
	LUT2 #(
		.INIT('h1)
	) name9946 (
		_w8633_,
		_w9476_,
		_w10478_
	);
	LUT2 #(
		.INIT('h8)
	) name9947 (
		_w10477_,
		_w10478_,
		_w10479_
	);
	LUT2 #(
		.INIT('h1)
	) name9948 (
		_w10476_,
		_w10479_,
		_w10480_
	);
	LUT2 #(
		.INIT('h1)
	) name9949 (
		\sa23_reg[0]/P0001 ,
		_w8668_,
		_w10481_
	);
	LUT2 #(
		.INIT('h4)
	) name9950 (
		_w10480_,
		_w10481_,
		_w10482_
	);
	LUT2 #(
		.INIT('h4)
	) name9951 (
		_w10474_,
		_w10482_,
		_w10483_
	);
	LUT2 #(
		.INIT('h1)
	) name9952 (
		_w10457_,
		_w10483_,
		_w10484_
	);
	LUT2 #(
		.INIT('h1)
	) name9953 (
		\sa23_reg[1]/P0001 ,
		_w8632_,
		_w10485_
	);
	LUT2 #(
		.INIT('h1)
	) name9954 (
		_w8641_,
		_w8663_,
		_w10486_
	);
	LUT2 #(
		.INIT('h4)
	) name9955 (
		_w9893_,
		_w10486_,
		_w10487_
	);
	LUT2 #(
		.INIT('h8)
	) name9956 (
		_w10485_,
		_w10487_,
		_w10488_
	);
	LUT2 #(
		.INIT('h1)
	) name9957 (
		_w8533_,
		_w8563_,
		_w10489_
	);
	LUT2 #(
		.INIT('h2)
	) name9958 (
		\sa23_reg[3]/P0001 ,
		_w10489_,
		_w10490_
	);
	LUT2 #(
		.INIT('h2)
	) name9959 (
		\sa23_reg[1]/P0001 ,
		_w9107_,
		_w10491_
	);
	LUT2 #(
		.INIT('h4)
	) name9960 (
		_w10490_,
		_w10491_,
		_w10492_
	);
	LUT2 #(
		.INIT('h1)
	) name9961 (
		_w10488_,
		_w10492_,
		_w10493_
	);
	LUT2 #(
		.INIT('h1)
	) name9962 (
		_w8670_,
		_w9467_,
		_w10494_
	);
	LUT2 #(
		.INIT('h4)
	) name9963 (
		_w10493_,
		_w10494_,
		_w10495_
	);
	LUT2 #(
		.INIT('h2)
	) name9964 (
		\sa23_reg[2]/P0001 ,
		_w10495_,
		_w10496_
	);
	LUT2 #(
		.INIT('h1)
	) name9965 (
		_w8509_,
		_w8568_,
		_w10497_
	);
	LUT2 #(
		.INIT('h1)
	) name9966 (
		_w8569_,
		_w10497_,
		_w10498_
	);
	LUT2 #(
		.INIT('h4)
	) name9967 (
		_w9085_,
		_w10465_,
		_w10499_
	);
	LUT2 #(
		.INIT('h4)
	) name9968 (
		_w10498_,
		_w10499_,
		_w10500_
	);
	LUT2 #(
		.INIT('h1)
	) name9969 (
		_w9078_,
		_w9927_,
		_w10501_
	);
	LUT2 #(
		.INIT('h4)
	) name9970 (
		_w8636_,
		_w10501_,
		_w10502_
	);
	LUT2 #(
		.INIT('h4)
	) name9971 (
		_w9467_,
		_w10502_,
		_w10503_
	);
	LUT2 #(
		.INIT('h8)
	) name9972 (
		_w10485_,
		_w10503_,
		_w10504_
	);
	LUT2 #(
		.INIT('h1)
	) name9973 (
		\sa23_reg[2]/P0001 ,
		_w10500_,
		_w10505_
	);
	LUT2 #(
		.INIT('h4)
	) name9974 (
		_w10504_,
		_w10505_,
		_w10506_
	);
	LUT2 #(
		.INIT('h1)
	) name9975 (
		_w10496_,
		_w10506_,
		_w10507_
	);
	LUT2 #(
		.INIT('h4)
	) name9976 (
		_w10484_,
		_w10507_,
		_w10508_
	);
	LUT2 #(
		.INIT('h2)
	) name9977 (
		\u0_w_reg[1][1]/P0001 ,
		_w10508_,
		_w10509_
	);
	LUT2 #(
		.INIT('h4)
	) name9978 (
		\u0_w_reg[1][1]/P0001 ,
		_w10508_,
		_w10510_
	);
	LUT2 #(
		.INIT('h1)
	) name9979 (
		_w10509_,
		_w10510_,
		_w10511_
	);
	LUT2 #(
		.INIT('h8)
	) name9980 (
		_w10433_,
		_w10511_,
		_w10512_
	);
	LUT2 #(
		.INIT('h1)
	) name9981 (
		_w10433_,
		_w10511_,
		_w10513_
	);
	LUT2 #(
		.INIT('h1)
	) name9982 (
		_w10512_,
		_w10513_,
		_w10514_
	);
	LUT2 #(
		.INIT('h1)
	) name9983 (
		_w10254_,
		_w10514_,
		_w10515_
	);
	LUT2 #(
		.INIT('h8)
	) name9984 (
		_w10254_,
		_w10514_,
		_w10516_
	);
	LUT2 #(
		.INIT('h1)
	) name9985 (
		\ld_r_reg/P0001 ,
		_w10515_,
		_w10517_
	);
	LUT2 #(
		.INIT('h4)
	) name9986 (
		_w10516_,
		_w10517_,
		_w10518_
	);
	LUT2 #(
		.INIT('h1)
	) name9987 (
		\text_in_r_reg[65]/P0001 ,
		\u0_w_reg[1][1]/P0001 ,
		_w10519_
	);
	LUT2 #(
		.INIT('h8)
	) name9988 (
		\text_in_r_reg[65]/P0001 ,
		\u0_w_reg[1][1]/P0001 ,
		_w10520_
	);
	LUT2 #(
		.INIT('h2)
	) name9989 (
		\ld_r_reg/P0001 ,
		_w10519_,
		_w10521_
	);
	LUT2 #(
		.INIT('h4)
	) name9990 (
		_w10520_,
		_w10521_,
		_w10522_
	);
	LUT2 #(
		.INIT('h1)
	) name9991 (
		_w10518_,
		_w10522_,
		_w10523_
	);
	LUT2 #(
		.INIT('h2)
	) name9992 (
		\u0_w_reg[1][28]/P0001 ,
		_w9639_,
		_w10524_
	);
	LUT2 #(
		.INIT('h4)
	) name9993 (
		\u0_w_reg[1][28]/P0001 ,
		_w9639_,
		_w10525_
	);
	LUT2 #(
		.INIT('h1)
	) name9994 (
		_w10524_,
		_w10525_,
		_w10526_
	);
	LUT2 #(
		.INIT('h8)
	) name9995 (
		_w9519_,
		_w10526_,
		_w10527_
	);
	LUT2 #(
		.INIT('h1)
	) name9996 (
		_w9519_,
		_w10526_,
		_w10528_
	);
	LUT2 #(
		.INIT('h1)
	) name9997 (
		_w10527_,
		_w10528_,
		_w10529_
	);
	LUT2 #(
		.INIT('h8)
	) name9998 (
		_w8228_,
		_w9197_,
		_w10530_
	);
	LUT2 #(
		.INIT('h8)
	) name9999 (
		_w8215_,
		_w8327_,
		_w10531_
	);
	LUT2 #(
		.INIT('h1)
	) name10000 (
		_w9710_,
		_w10531_,
		_w10532_
	);
	LUT2 #(
		.INIT('h4)
	) name10001 (
		_w9387_,
		_w10532_,
		_w10533_
	);
	LUT2 #(
		.INIT('h1)
	) name10002 (
		_w9389_,
		_w10530_,
		_w10534_
	);
	LUT2 #(
		.INIT('h8)
	) name10003 (
		_w10533_,
		_w10534_,
		_w10535_
	);
	LUT2 #(
		.INIT('h1)
	) name10004 (
		\sa01_reg[1]/P0001 ,
		_w10535_,
		_w10536_
	);
	LUT2 #(
		.INIT('h1)
	) name10005 (
		_w9216_,
		_w9357_,
		_w10537_
	);
	LUT2 #(
		.INIT('h2)
	) name10006 (
		\sa01_reg[2]/P0001 ,
		_w10537_,
		_w10538_
	);
	LUT2 #(
		.INIT('h8)
	) name10007 (
		_w8246_,
		_w8279_,
		_w10539_
	);
	LUT2 #(
		.INIT('h1)
	) name10008 (
		_w8255_,
		_w10083_,
		_w10540_
	);
	LUT2 #(
		.INIT('h4)
	) name10009 (
		_w10539_,
		_w10540_,
		_w10541_
	);
	LUT2 #(
		.INIT('h4)
	) name10010 (
		_w8322_,
		_w10541_,
		_w10542_
	);
	LUT2 #(
		.INIT('h4)
	) name10011 (
		_w10538_,
		_w10542_,
		_w10543_
	);
	LUT2 #(
		.INIT('h2)
	) name10012 (
		\sa01_reg[1]/P0001 ,
		_w10543_,
		_w10544_
	);
	LUT2 #(
		.INIT('h1)
	) name10013 (
		\sa01_reg[2]/P0001 ,
		_w9323_,
		_w10545_
	);
	LUT2 #(
		.INIT('h8)
	) name10014 (
		_w8329_,
		_w9216_,
		_w10546_
	);
	LUT2 #(
		.INIT('h1)
	) name10015 (
		_w9253_,
		_w9374_,
		_w10547_
	);
	LUT2 #(
		.INIT('h4)
	) name10016 (
		_w10546_,
		_w10547_,
		_w10548_
	);
	LUT2 #(
		.INIT('h4)
	) name10017 (
		_w10545_,
		_w10548_,
		_w10549_
	);
	LUT2 #(
		.INIT('h4)
	) name10018 (
		_w10536_,
		_w10549_,
		_w10550_
	);
	LUT2 #(
		.INIT('h4)
	) name10019 (
		_w10544_,
		_w10550_,
		_w10551_
	);
	LUT2 #(
		.INIT('h1)
	) name10020 (
		\sa01_reg[0]/P0001 ,
		_w10551_,
		_w10552_
	);
	LUT2 #(
		.INIT('h2)
	) name10021 (
		_w8353_,
		_w9741_,
		_w10553_
	);
	LUT2 #(
		.INIT('h2)
	) name10022 (
		\sa01_reg[2]/P0001 ,
		_w8277_,
		_w10554_
	);
	LUT2 #(
		.INIT('h4)
	) name10023 (
		_w9231_,
		_w10554_,
		_w10555_
	);
	LUT2 #(
		.INIT('h1)
	) name10024 (
		_w10553_,
		_w10555_,
		_w10556_
	);
	LUT2 #(
		.INIT('h1)
	) name10025 (
		_w8362_,
		_w9376_,
		_w10557_
	);
	LUT2 #(
		.INIT('h4)
	) name10026 (
		_w9322_,
		_w10557_,
		_w10558_
	);
	LUT2 #(
		.INIT('h4)
	) name10027 (
		_w10157_,
		_w10558_,
		_w10559_
	);
	LUT2 #(
		.INIT('h4)
	) name10028 (
		_w10556_,
		_w10559_,
		_w10560_
	);
	LUT2 #(
		.INIT('h1)
	) name10029 (
		\sa01_reg[1]/P0001 ,
		_w10560_,
		_w10561_
	);
	LUT2 #(
		.INIT('h4)
	) name10030 (
		_w9710_,
		_w10203_,
		_w10562_
	);
	LUT2 #(
		.INIT('h1)
	) name10031 (
		\sa01_reg[2]/P0001 ,
		_w10562_,
		_w10563_
	);
	LUT2 #(
		.INIT('h4)
	) name10032 (
		_w9183_,
		_w9263_,
		_w10564_
	);
	LUT2 #(
		.INIT('h2)
	) name10033 (
		_w8327_,
		_w10564_,
		_w10565_
	);
	LUT2 #(
		.INIT('h2)
	) name10034 (
		_w8240_,
		_w8242_,
		_w10566_
	);
	LUT2 #(
		.INIT('h1)
	) name10035 (
		_w9215_,
		_w10566_,
		_w10567_
	);
	LUT2 #(
		.INIT('h1)
	) name10036 (
		_w8264_,
		_w10567_,
		_w10568_
	);
	LUT2 #(
		.INIT('h1)
	) name10037 (
		_w8279_,
		_w8331_,
		_w10569_
	);
	LUT2 #(
		.INIT('h4)
	) name10038 (
		_w9184_,
		_w10569_,
		_w10570_
	);
	LUT2 #(
		.INIT('h2)
	) name10039 (
		\sa01_reg[2]/P0001 ,
		_w10570_,
		_w10571_
	);
	LUT2 #(
		.INIT('h1)
	) name10040 (
		_w8269_,
		_w10568_,
		_w10572_
	);
	LUT2 #(
		.INIT('h4)
	) name10041 (
		_w10571_,
		_w10572_,
		_w10573_
	);
	LUT2 #(
		.INIT('h2)
	) name10042 (
		\sa01_reg[1]/P0001 ,
		_w10573_,
		_w10574_
	);
	LUT2 #(
		.INIT('h1)
	) name10043 (
		_w9256_,
		_w10565_,
		_w10575_
	);
	LUT2 #(
		.INIT('h4)
	) name10044 (
		_w10563_,
		_w10575_,
		_w10576_
	);
	LUT2 #(
		.INIT('h4)
	) name10045 (
		_w10561_,
		_w10576_,
		_w10577_
	);
	LUT2 #(
		.INIT('h4)
	) name10046 (
		_w10574_,
		_w10577_,
		_w10578_
	);
	LUT2 #(
		.INIT('h2)
	) name10047 (
		\sa01_reg[0]/P0001 ,
		_w10578_,
		_w10579_
	);
	LUT2 #(
		.INIT('h8)
	) name10048 (
		_w8236_,
		_w10145_,
		_w10580_
	);
	LUT2 #(
		.INIT('h4)
	) name10049 (
		\sa01_reg[2]/P0001 ,
		_w8333_,
		_w10581_
	);
	LUT2 #(
		.INIT('h8)
	) name10050 (
		\sa01_reg[6]/NET0131 ,
		_w8265_,
		_w10582_
	);
	LUT2 #(
		.INIT('h1)
	) name10051 (
		_w9180_,
		_w9352_,
		_w10583_
	);
	LUT2 #(
		.INIT('h4)
	) name10052 (
		_w10582_,
		_w10583_,
		_w10584_
	);
	LUT2 #(
		.INIT('h2)
	) name10053 (
		_w9694_,
		_w10584_,
		_w10585_
	);
	LUT2 #(
		.INIT('h1)
	) name10054 (
		_w8244_,
		_w10581_,
		_w10586_
	);
	LUT2 #(
		.INIT('h4)
	) name10055 (
		_w10585_,
		_w10586_,
		_w10587_
	);
	LUT2 #(
		.INIT('h2)
	) name10056 (
		\sa01_reg[1]/P0001 ,
		_w10587_,
		_w10588_
	);
	LUT2 #(
		.INIT('h1)
	) name10057 (
		_w8217_,
		_w9253_,
		_w10589_
	);
	LUT2 #(
		.INIT('h2)
	) name10058 (
		_w9318_,
		_w10589_,
		_w10590_
	);
	LUT2 #(
		.INIT('h8)
	) name10059 (
		_w8218_,
		_w8257_,
		_w10591_
	);
	LUT2 #(
		.INIT('h1)
	) name10060 (
		_w8269_,
		_w10591_,
		_w10592_
	);
	LUT2 #(
		.INIT('h2)
	) name10061 (
		_w9388_,
		_w10592_,
		_w10593_
	);
	LUT2 #(
		.INIT('h8)
	) name10062 (
		\sa01_reg[7]/NET0131 ,
		_w9699_,
		_w10594_
	);
	LUT2 #(
		.INIT('h1)
	) name10063 (
		_w10116_,
		_w10144_,
		_w10595_
	);
	LUT2 #(
		.INIT('h4)
	) name10064 (
		_w10580_,
		_w10595_,
		_w10596_
	);
	LUT2 #(
		.INIT('h1)
	) name10065 (
		_w10593_,
		_w10594_,
		_w10597_
	);
	LUT2 #(
		.INIT('h8)
	) name10066 (
		_w10596_,
		_w10597_,
		_w10598_
	);
	LUT2 #(
		.INIT('h4)
	) name10067 (
		_w10590_,
		_w10598_,
		_w10599_
	);
	LUT2 #(
		.INIT('h4)
	) name10068 (
		_w10588_,
		_w10599_,
		_w10600_
	);
	LUT2 #(
		.INIT('h4)
	) name10069 (
		_w10552_,
		_w10600_,
		_w10601_
	);
	LUT2 #(
		.INIT('h4)
	) name10070 (
		_w10579_,
		_w10601_,
		_w10602_
	);
	LUT2 #(
		.INIT('h2)
	) name10071 (
		_w9783_,
		_w10602_,
		_w10603_
	);
	LUT2 #(
		.INIT('h4)
	) name10072 (
		_w9783_,
		_w10602_,
		_w10604_
	);
	LUT2 #(
		.INIT('h1)
	) name10073 (
		_w10603_,
		_w10604_,
		_w10605_
	);
	LUT2 #(
		.INIT('h4)
	) name10074 (
		\sa12_reg[4]/P0001 ,
		_w8413_,
		_w10606_
	);
	LUT2 #(
		.INIT('h1)
	) name10075 (
		_w8414_,
		_w8495_,
		_w10607_
	);
	LUT2 #(
		.INIT('h2)
	) name10076 (
		\sa12_reg[2]/P0001 ,
		_w10607_,
		_w10608_
	);
	LUT2 #(
		.INIT('h8)
	) name10077 (
		_w8077_,
		_w9846_,
		_w10609_
	);
	LUT2 #(
		.INIT('h2)
	) name10078 (
		\sa12_reg[1]/P0001 ,
		_w8127_,
		_w10610_
	);
	LUT2 #(
		.INIT('h4)
	) name10079 (
		_w8115_,
		_w10610_,
		_w10611_
	);
	LUT2 #(
		.INIT('h1)
	) name10080 (
		_w9996_,
		_w10609_,
		_w10612_
	);
	LUT2 #(
		.INIT('h8)
	) name10081 (
		_w10611_,
		_w10612_,
		_w10613_
	);
	LUT2 #(
		.INIT('h4)
	) name10082 (
		_w10608_,
		_w10613_,
		_w10614_
	);
	LUT2 #(
		.INIT('h4)
	) name10083 (
		_w8082_,
		_w8084_,
		_w10615_
	);
	LUT2 #(
		.INIT('h1)
	) name10084 (
		_w8156_,
		_w10615_,
		_w10616_
	);
	LUT2 #(
		.INIT('h2)
	) name10085 (
		\sa12_reg[2]/P0001 ,
		_w10616_,
		_w10617_
	);
	LUT2 #(
		.INIT('h1)
	) name10086 (
		\sa12_reg[1]/P0001 ,
		_w9801_,
		_w10618_
	);
	LUT2 #(
		.INIT('h4)
	) name10087 (
		_w9034_,
		_w10618_,
		_w10619_
	);
	LUT2 #(
		.INIT('h4)
	) name10088 (
		_w9041_,
		_w10619_,
		_w10620_
	);
	LUT2 #(
		.INIT('h4)
	) name10089 (
		_w10617_,
		_w10620_,
		_w10621_
	);
	LUT2 #(
		.INIT('h1)
	) name10090 (
		_w10614_,
		_w10621_,
		_w10622_
	);
	LUT2 #(
		.INIT('h1)
	) name10091 (
		\sa12_reg[2]/P0001 ,
		_w8993_,
		_w10623_
	);
	LUT2 #(
		.INIT('h8)
	) name10092 (
		_w8110_,
		_w8498_,
		_w10624_
	);
	LUT2 #(
		.INIT('h1)
	) name10093 (
		_w9044_,
		_w10624_,
		_w10625_
	);
	LUT2 #(
		.INIT('h2)
	) name10094 (
		\sa12_reg[2]/P0001 ,
		_w10625_,
		_w10626_
	);
	LUT2 #(
		.INIT('h1)
	) name10095 (
		_w10606_,
		_w10626_,
		_w10627_
	);
	LUT2 #(
		.INIT('h4)
	) name10096 (
		_w10623_,
		_w10627_,
		_w10628_
	);
	LUT2 #(
		.INIT('h4)
	) name10097 (
		_w10622_,
		_w10628_,
		_w10629_
	);
	LUT2 #(
		.INIT('h1)
	) name10098 (
		\sa12_reg[0]/P0001 ,
		_w10629_,
		_w10630_
	);
	LUT2 #(
		.INIT('h4)
	) name10099 (
		_w8077_,
		_w9841_,
		_w10631_
	);
	LUT2 #(
		.INIT('h1)
	) name10100 (
		_w8165_,
		_w10631_,
		_w10632_
	);
	LUT2 #(
		.INIT('h1)
	) name10101 (
		_w8075_,
		_w10632_,
		_w10633_
	);
	LUT2 #(
		.INIT('h1)
	) name10102 (
		_w8182_,
		_w8185_,
		_w10634_
	);
	LUT2 #(
		.INIT('h4)
	) name10103 (
		_w10055_,
		_w10634_,
		_w10635_
	);
	LUT2 #(
		.INIT('h2)
	) name10104 (
		\sa12_reg[2]/P0001 ,
		_w10635_,
		_w10636_
	);
	LUT2 #(
		.INIT('h1)
	) name10105 (
		_w8136_,
		_w10633_,
		_w10637_
	);
	LUT2 #(
		.INIT('h4)
	) name10106 (
		_w10636_,
		_w10637_,
		_w10638_
	);
	LUT2 #(
		.INIT('h2)
	) name10107 (
		\sa12_reg[1]/P0001 ,
		_w10638_,
		_w10639_
	);
	LUT2 #(
		.INIT('h8)
	) name10108 (
		\sa12_reg[6]/NET0131 ,
		_w8389_,
		_w10640_
	);
	LUT2 #(
		.INIT('h1)
	) name10109 (
		_w8461_,
		_w10640_,
		_w10641_
	);
	LUT2 #(
		.INIT('h4)
	) name10110 (
		_w9801_,
		_w10641_,
		_w10642_
	);
	LUT2 #(
		.INIT('h1)
	) name10111 (
		\sa12_reg[2]/P0001 ,
		_w10642_,
		_w10643_
	);
	LUT2 #(
		.INIT('h4)
	) name10112 (
		_w8381_,
		_w8482_,
		_w10644_
	);
	LUT2 #(
		.INIT('h2)
	) name10113 (
		_w8066_,
		_w10644_,
		_w10645_
	);
	LUT2 #(
		.INIT('h1)
	) name10114 (
		_w8096_,
		_w9042_,
		_w10646_
	);
	LUT2 #(
		.INIT('h1)
	) name10115 (
		\sa12_reg[2]/P0001 ,
		_w10646_,
		_w10647_
	);
	LUT2 #(
		.INIT('h1)
	) name10116 (
		_w8127_,
		_w8443_,
		_w10648_
	);
	LUT2 #(
		.INIT('h1)
	) name10117 (
		_w8162_,
		_w10648_,
		_w10649_
	);
	LUT2 #(
		.INIT('h1)
	) name10118 (
		_w8394_,
		_w8485_,
		_w10650_
	);
	LUT2 #(
		.INIT('h4)
	) name10119 (
		_w8189_,
		_w10650_,
		_w10651_
	);
	LUT2 #(
		.INIT('h4)
	) name10120 (
		_w10647_,
		_w10651_,
		_w10652_
	);
	LUT2 #(
		.INIT('h4)
	) name10121 (
		_w10649_,
		_w10652_,
		_w10653_
	);
	LUT2 #(
		.INIT('h1)
	) name10122 (
		\sa12_reg[1]/P0001 ,
		_w10653_,
		_w10654_
	);
	LUT2 #(
		.INIT('h1)
	) name10123 (
		_w8449_,
		_w10645_,
		_w10655_
	);
	LUT2 #(
		.INIT('h4)
	) name10124 (
		_w10643_,
		_w10655_,
		_w10656_
	);
	LUT2 #(
		.INIT('h4)
	) name10125 (
		_w10639_,
		_w10656_,
		_w10657_
	);
	LUT2 #(
		.INIT('h4)
	) name10126 (
		_w10654_,
		_w10657_,
		_w10658_
	);
	LUT2 #(
		.INIT('h2)
	) name10127 (
		\sa12_reg[0]/P0001 ,
		_w10658_,
		_w10659_
	);
	LUT2 #(
		.INIT('h8)
	) name10128 (
		\sa12_reg[2]/P0001 ,
		_w8136_,
		_w10660_
	);
	LUT2 #(
		.INIT('h8)
	) name10129 (
		_w8159_,
		_w10060_,
		_w10661_
	);
	LUT2 #(
		.INIT('h1)
	) name10130 (
		_w10660_,
		_w10661_,
		_w10662_
	);
	LUT2 #(
		.INIT('h1)
	) name10131 (
		\sa12_reg[4]/P0001 ,
		_w10662_,
		_w10663_
	);
	LUT2 #(
		.INIT('h1)
	) name10132 (
		_w8097_,
		_w8136_,
		_w10664_
	);
	LUT2 #(
		.INIT('h2)
	) name10133 (
		_w9033_,
		_w10664_,
		_w10665_
	);
	LUT2 #(
		.INIT('h8)
	) name10134 (
		_w8059_,
		_w9034_,
		_w10666_
	);
	LUT2 #(
		.INIT('h1)
	) name10135 (
		_w8448_,
		_w10666_,
		_w10667_
	);
	LUT2 #(
		.INIT('h1)
	) name10136 (
		\sa12_reg[1]/P0001 ,
		_w10667_,
		_w10668_
	);
	LUT2 #(
		.INIT('h1)
	) name10137 (
		_w8146_,
		_w8388_,
		_w10669_
	);
	LUT2 #(
		.INIT('h4)
	) name10138 (
		_w9025_,
		_w10669_,
		_w10670_
	);
	LUT2 #(
		.INIT('h2)
	) name10139 (
		_w8978_,
		_w10670_,
		_w10671_
	);
	LUT2 #(
		.INIT('h4)
	) name10140 (
		\sa12_reg[2]/P0001 ,
		_w8113_,
		_w10672_
	);
	LUT2 #(
		.INIT('h1)
	) name10141 (
		_w8167_,
		_w10672_,
		_w10673_
	);
	LUT2 #(
		.INIT('h4)
	) name10142 (
		_w10671_,
		_w10673_,
		_w10674_
	);
	LUT2 #(
		.INIT('h2)
	) name10143 (
		\sa12_reg[1]/P0001 ,
		_w10674_,
		_w10675_
	);
	LUT2 #(
		.INIT('h1)
	) name10144 (
		_w10024_,
		_w10063_,
		_w10676_
	);
	LUT2 #(
		.INIT('h4)
	) name10145 (
		_w10665_,
		_w10676_,
		_w10677_
	);
	LUT2 #(
		.INIT('h4)
	) name10146 (
		_w10663_,
		_w10677_,
		_w10678_
	);
	LUT2 #(
		.INIT('h4)
	) name10147 (
		_w10668_,
		_w10678_,
		_w10679_
	);
	LUT2 #(
		.INIT('h4)
	) name10148 (
		_w10675_,
		_w10679_,
		_w10680_
	);
	LUT2 #(
		.INIT('h4)
	) name10149 (
		_w10630_,
		_w10680_,
		_w10681_
	);
	LUT2 #(
		.INIT('h4)
	) name10150 (
		_w10659_,
		_w10681_,
		_w10682_
	);
	LUT2 #(
		.INIT('h2)
	) name10151 (
		_w9874_,
		_w10682_,
		_w10683_
	);
	LUT2 #(
		.INIT('h4)
	) name10152 (
		_w9874_,
		_w10682_,
		_w10684_
	);
	LUT2 #(
		.INIT('h1)
	) name10153 (
		_w10683_,
		_w10684_,
		_w10685_
	);
	LUT2 #(
		.INIT('h4)
	) name10154 (
		_w10605_,
		_w10685_,
		_w10686_
	);
	LUT2 #(
		.INIT('h2)
	) name10155 (
		_w10605_,
		_w10685_,
		_w10687_
	);
	LUT2 #(
		.INIT('h1)
	) name10156 (
		_w10686_,
		_w10687_,
		_w10688_
	);
	LUT2 #(
		.INIT('h2)
	) name10157 (
		_w10529_,
		_w10688_,
		_w10689_
	);
	LUT2 #(
		.INIT('h4)
	) name10158 (
		_w10529_,
		_w10688_,
		_w10690_
	);
	LUT2 #(
		.INIT('h1)
	) name10159 (
		\ld_r_reg/P0001 ,
		_w10689_,
		_w10691_
	);
	LUT2 #(
		.INIT('h4)
	) name10160 (
		_w10690_,
		_w10691_,
		_w10692_
	);
	LUT2 #(
		.INIT('h2)
	) name10161 (
		\text_in_r_reg[92]/P0001 ,
		\u0_w_reg[1][28]/P0001 ,
		_w10693_
	);
	LUT2 #(
		.INIT('h4)
	) name10162 (
		\text_in_r_reg[92]/P0001 ,
		\u0_w_reg[1][28]/P0001 ,
		_w10694_
	);
	LUT2 #(
		.INIT('h2)
	) name10163 (
		\ld_r_reg/P0001 ,
		_w10693_,
		_w10695_
	);
	LUT2 #(
		.INIT('h4)
	) name10164 (
		_w10694_,
		_w10695_,
		_w10696_
	);
	LUT2 #(
		.INIT('h1)
	) name10165 (
		_w10692_,
		_w10696_,
		_w10697_
	);
	LUT2 #(
		.INIT('h4)
	) name10166 (
		_w8588_,
		_w9113_,
		_w10698_
	);
	LUT2 #(
		.INIT('h1)
	) name10167 (
		_w8509_,
		_w9499_,
		_w10699_
	);
	LUT2 #(
		.INIT('h4)
	) name10168 (
		_w9920_,
		_w10699_,
		_w10700_
	);
	LUT2 #(
		.INIT('h2)
	) name10169 (
		\sa23_reg[2]/P0001 ,
		_w10700_,
		_w10701_
	);
	LUT2 #(
		.INIT('h4)
	) name10170 (
		\sa23_reg[2]/P0001 ,
		_w9489_,
		_w10702_
	);
	LUT2 #(
		.INIT('h8)
	) name10171 (
		_w8513_,
		_w9079_,
		_w10703_
	);
	LUT2 #(
		.INIT('h1)
	) name10172 (
		_w9097_,
		_w10703_,
		_w10704_
	);
	LUT2 #(
		.INIT('h1)
	) name10173 (
		_w10698_,
		_w10702_,
		_w10705_
	);
	LUT2 #(
		.INIT('h8)
	) name10174 (
		_w10704_,
		_w10705_,
		_w10706_
	);
	LUT2 #(
		.INIT('h4)
	) name10175 (
		_w10701_,
		_w10706_,
		_w10707_
	);
	LUT2 #(
		.INIT('h2)
	) name10176 (
		\sa23_reg[1]/P0001 ,
		_w10707_,
		_w10708_
	);
	LUT2 #(
		.INIT('h1)
	) name10177 (
		_w8598_,
		_w8615_,
		_w10709_
	);
	LUT2 #(
		.INIT('h8)
	) name10178 (
		_w9497_,
		_w10709_,
		_w10710_
	);
	LUT2 #(
		.INIT('h1)
	) name10179 (
		\sa23_reg[2]/P0001 ,
		_w8527_,
		_w10711_
	);
	LUT2 #(
		.INIT('h4)
	) name10180 (
		_w9927_,
		_w10711_,
		_w10712_
	);
	LUT2 #(
		.INIT('h1)
	) name10181 (
		_w10710_,
		_w10712_,
		_w10713_
	);
	LUT2 #(
		.INIT('h1)
	) name10182 (
		_w8663_,
		_w9158_,
		_w10714_
	);
	LUT2 #(
		.INIT('h4)
	) name10183 (
		_w9467_,
		_w10714_,
		_w10715_
	);
	LUT2 #(
		.INIT('h4)
	) name10184 (
		_w10713_,
		_w10715_,
		_w10716_
	);
	LUT2 #(
		.INIT('h1)
	) name10185 (
		\sa23_reg[1]/P0001 ,
		_w10716_,
		_w10717_
	);
	LUT2 #(
		.INIT('h8)
	) name10186 (
		\sa23_reg[6]/NET0131 ,
		_w8532_,
		_w10718_
	);
	LUT2 #(
		.INIT('h1)
	) name10187 (
		_w8633_,
		_w10718_,
		_w10719_
	);
	LUT2 #(
		.INIT('h4)
	) name10188 (
		_w9468_,
		_w10719_,
		_w10720_
	);
	LUT2 #(
		.INIT('h1)
	) name10189 (
		\sa23_reg[2]/P0001 ,
		_w10720_,
		_w10721_
	);
	LUT2 #(
		.INIT('h4)
	) name10190 (
		_w8512_,
		_w8656_,
		_w10722_
	);
	LUT2 #(
		.INIT('h2)
	) name10191 (
		_w9931_,
		_w10722_,
		_w10723_
	);
	LUT2 #(
		.INIT('h1)
	) name10192 (
		_w8647_,
		_w10723_,
		_w10724_
	);
	LUT2 #(
		.INIT('h4)
	) name10193 (
		_w10721_,
		_w10724_,
		_w10725_
	);
	LUT2 #(
		.INIT('h4)
	) name10194 (
		_w10708_,
		_w10725_,
		_w10726_
	);
	LUT2 #(
		.INIT('h4)
	) name10195 (
		_w10717_,
		_w10726_,
		_w10727_
	);
	LUT2 #(
		.INIT('h2)
	) name10196 (
		\sa23_reg[0]/P0001 ,
		_w10727_,
		_w10728_
	);
	LUT2 #(
		.INIT('h4)
	) name10197 (
		\sa23_reg[2]/P0001 ,
		_w9454_,
		_w10729_
	);
	LUT2 #(
		.INIT('h8)
	) name10198 (
		_w8521_,
		_w8572_,
		_w10730_
	);
	LUT2 #(
		.INIT('h1)
	) name10199 (
		_w9097_,
		_w10730_,
		_w10731_
	);
	LUT2 #(
		.INIT('h2)
	) name10200 (
		\sa23_reg[2]/P0001 ,
		_w10731_,
		_w10732_
	);
	LUT2 #(
		.INIT('h1)
	) name10201 (
		_w8514_,
		_w8520_,
		_w10733_
	);
	LUT2 #(
		.INIT('h4)
	) name10202 (
		_w9099_,
		_w10733_,
		_w10734_
	);
	LUT2 #(
		.INIT('h2)
	) name10203 (
		_w9079_,
		_w10734_,
		_w10735_
	);
	LUT2 #(
		.INIT('h1)
	) name10204 (
		_w9433_,
		_w10729_,
		_w10736_
	);
	LUT2 #(
		.INIT('h4)
	) name10205 (
		_w10732_,
		_w10736_,
		_w10737_
	);
	LUT2 #(
		.INIT('h4)
	) name10206 (
		_w10735_,
		_w10737_,
		_w10738_
	);
	LUT2 #(
		.INIT('h2)
	) name10207 (
		\sa23_reg[1]/P0001 ,
		_w10738_,
		_w10739_
	);
	LUT2 #(
		.INIT('h1)
	) name10208 (
		_w9125_,
		_w9964_,
		_w10740_
	);
	LUT2 #(
		.INIT('h2)
	) name10209 (
		_w9112_,
		_w10740_,
		_w10741_
	);
	LUT2 #(
		.INIT('h8)
	) name10210 (
		_w8588_,
		_w9922_,
		_w10742_
	);
	LUT2 #(
		.INIT('h1)
	) name10211 (
		_w10741_,
		_w10742_,
		_w10743_
	);
	LUT2 #(
		.INIT('h1)
	) name10212 (
		\sa23_reg[1]/P0001 ,
		_w10743_,
		_w10744_
	);
	LUT2 #(
		.INIT('h1)
	) name10213 (
		_w8563_,
		_w9420_,
		_w10745_
	);
	LUT2 #(
		.INIT('h2)
	) name10214 (
		_w8546_,
		_w10745_,
		_w10746_
	);
	LUT2 #(
		.INIT('h4)
	) name10215 (
		\sa23_reg[2]/P0001 ,
		_w9088_,
		_w10747_
	);
	LUT2 #(
		.INIT('h8)
	) name10216 (
		_w8529_,
		_w8577_,
		_w10748_
	);
	LUT2 #(
		.INIT('h1)
	) name10217 (
		_w9101_,
		_w9114_,
		_w10749_
	);
	LUT2 #(
		.INIT('h2)
	) name10218 (
		\sa23_reg[1]/P0001 ,
		_w10749_,
		_w10750_
	);
	LUT2 #(
		.INIT('h2)
	) name10219 (
		_w9148_,
		_w10748_,
		_w10751_
	);
	LUT2 #(
		.INIT('h4)
	) name10220 (
		_w10750_,
		_w10751_,
		_w10752_
	);
	LUT2 #(
		.INIT('h1)
	) name10221 (
		_w10747_,
		_w10752_,
		_w10753_
	);
	LUT2 #(
		.INIT('h8)
	) name10222 (
		\sa23_reg[2]/P0001 ,
		_w8526_,
		_w10754_
	);
	LUT2 #(
		.INIT('h4)
	) name10223 (
		_w8547_,
		_w10754_,
		_w10755_
	);
	LUT2 #(
		.INIT('h1)
	) name10224 (
		_w8547_,
		_w8660_,
		_w10756_
	);
	LUT2 #(
		.INIT('h2)
	) name10225 (
		_w8623_,
		_w10756_,
		_w10757_
	);
	LUT2 #(
		.INIT('h1)
	) name10226 (
		\sa23_reg[1]/P0001 ,
		_w9468_,
		_w10758_
	);
	LUT2 #(
		.INIT('h1)
	) name10227 (
		_w10755_,
		_w10757_,
		_w10759_
	);
	LUT2 #(
		.INIT('h8)
	) name10228 (
		_w10758_,
		_w10759_,
		_w10760_
	);
	LUT2 #(
		.INIT('h4)
	) name10229 (
		_w9134_,
		_w10760_,
		_w10761_
	);
	LUT2 #(
		.INIT('h8)
	) name10230 (
		_w8508_,
		_w9922_,
		_w10762_
	);
	LUT2 #(
		.INIT('h2)
	) name10231 (
		\sa23_reg[1]/P0001 ,
		_w8615_,
		_w10763_
	);
	LUT2 #(
		.INIT('h4)
	) name10232 (
		_w8558_,
		_w10763_,
		_w10764_
	);
	LUT2 #(
		.INIT('h1)
	) name10233 (
		_w10442_,
		_w10762_,
		_w10765_
	);
	LUT2 #(
		.INIT('h8)
	) name10234 (
		_w10764_,
		_w10765_,
		_w10766_
	);
	LUT2 #(
		.INIT('h1)
	) name10235 (
		_w10761_,
		_w10766_,
		_w10767_
	);
	LUT2 #(
		.INIT('h1)
	) name10236 (
		_w8643_,
		_w10753_,
		_w10768_
	);
	LUT2 #(
		.INIT('h4)
	) name10237 (
		_w10767_,
		_w10768_,
		_w10769_
	);
	LUT2 #(
		.INIT('h1)
	) name10238 (
		\sa23_reg[0]/P0001 ,
		_w10769_,
		_w10770_
	);
	LUT2 #(
		.INIT('h1)
	) name10239 (
		_w9130_,
		_w10746_,
		_w10771_
	);
	LUT2 #(
		.INIT('h4)
	) name10240 (
		_w10744_,
		_w10771_,
		_w10772_
	);
	LUT2 #(
		.INIT('h4)
	) name10241 (
		_w10739_,
		_w10772_,
		_w10773_
	);
	LUT2 #(
		.INIT('h4)
	) name10242 (
		_w10728_,
		_w10773_,
		_w10774_
	);
	LUT2 #(
		.INIT('h4)
	) name10243 (
		_w10770_,
		_w10774_,
		_w10775_
	);
	LUT2 #(
		.INIT('h2)
	) name10244 (
		_w8376_,
		_w10775_,
		_w10776_
	);
	LUT2 #(
		.INIT('h4)
	) name10245 (
		_w8376_,
		_w10775_,
		_w10777_
	);
	LUT2 #(
		.INIT('h1)
	) name10246 (
		_w10776_,
		_w10777_,
		_w10778_
	);
	LUT2 #(
		.INIT('h8)
	) name10247 (
		_w10685_,
		_w10778_,
		_w10779_
	);
	LUT2 #(
		.INIT('h1)
	) name10248 (
		_w10685_,
		_w10778_,
		_w10780_
	);
	LUT2 #(
		.INIT('h1)
	) name10249 (
		_w10779_,
		_w10780_,
		_w10781_
	);
	LUT2 #(
		.INIT('h1)
	) name10250 (
		_w9516_,
		_w9639_,
		_w10782_
	);
	LUT2 #(
		.INIT('h8)
	) name10251 (
		_w9516_,
		_w9639_,
		_w10783_
	);
	LUT2 #(
		.INIT('h1)
	) name10252 (
		_w10782_,
		_w10783_,
		_w10784_
	);
	LUT2 #(
		.INIT('h2)
	) name10253 (
		\u0_w_reg[1][20]/P0001 ,
		_w9980_,
		_w10785_
	);
	LUT2 #(
		.INIT('h4)
	) name10254 (
		\u0_w_reg[1][20]/P0001 ,
		_w9980_,
		_w10786_
	);
	LUT2 #(
		.INIT('h1)
	) name10255 (
		_w10785_,
		_w10786_,
		_w10787_
	);
	LUT2 #(
		.INIT('h8)
	) name10256 (
		_w10784_,
		_w10787_,
		_w10788_
	);
	LUT2 #(
		.INIT('h1)
	) name10257 (
		_w10784_,
		_w10787_,
		_w10789_
	);
	LUT2 #(
		.INIT('h1)
	) name10258 (
		_w10788_,
		_w10789_,
		_w10790_
	);
	LUT2 #(
		.INIT('h2)
	) name10259 (
		_w10781_,
		_w10790_,
		_w10791_
	);
	LUT2 #(
		.INIT('h4)
	) name10260 (
		_w10781_,
		_w10790_,
		_w10792_
	);
	LUT2 #(
		.INIT('h1)
	) name10261 (
		\ld_r_reg/P0001 ,
		_w10791_,
		_w10793_
	);
	LUT2 #(
		.INIT('h4)
	) name10262 (
		_w10792_,
		_w10793_,
		_w10794_
	);
	LUT2 #(
		.INIT('h2)
	) name10263 (
		\text_in_r_reg[84]/P0001 ,
		\u0_w_reg[1][20]/P0001 ,
		_w10795_
	);
	LUT2 #(
		.INIT('h4)
	) name10264 (
		\text_in_r_reg[84]/P0001 ,
		\u0_w_reg[1][20]/P0001 ,
		_w10796_
	);
	LUT2 #(
		.INIT('h2)
	) name10265 (
		\ld_r_reg/P0001 ,
		_w10795_,
		_w10797_
	);
	LUT2 #(
		.INIT('h4)
	) name10266 (
		_w10796_,
		_w10797_,
		_w10798_
	);
	LUT2 #(
		.INIT('h1)
	) name10267 (
		_w10794_,
		_w10798_,
		_w10799_
	);
	LUT2 #(
		.INIT('h1)
	) name10268 (
		_w8376_,
		_w9292_,
		_w10800_
	);
	LUT2 #(
		.INIT('h8)
	) name10269 (
		_w8376_,
		_w9292_,
		_w10801_
	);
	LUT2 #(
		.INIT('h1)
	) name10270 (
		_w10800_,
		_w10801_,
		_w10802_
	);
	LUT2 #(
		.INIT('h2)
	) name10271 (
		\u0_w_reg[1][5]/P0001 ,
		_w9639_,
		_w10803_
	);
	LUT2 #(
		.INIT('h4)
	) name10272 (
		\u0_w_reg[1][5]/P0001 ,
		_w9639_,
		_w10804_
	);
	LUT2 #(
		.INIT('h1)
	) name10273 (
		_w10803_,
		_w10804_,
		_w10805_
	);
	LUT2 #(
		.INIT('h8)
	) name10274 (
		_w8678_,
		_w10805_,
		_w10806_
	);
	LUT2 #(
		.INIT('h1)
	) name10275 (
		_w8678_,
		_w10805_,
		_w10807_
	);
	LUT2 #(
		.INIT('h1)
	) name10276 (
		_w10806_,
		_w10807_,
		_w10808_
	);
	LUT2 #(
		.INIT('h4)
	) name10277 (
		_w10802_,
		_w10808_,
		_w10809_
	);
	LUT2 #(
		.INIT('h2)
	) name10278 (
		_w10802_,
		_w10808_,
		_w10810_
	);
	LUT2 #(
		.INIT('h1)
	) name10279 (
		\ld_r_reg/P0001 ,
		_w10809_,
		_w10811_
	);
	LUT2 #(
		.INIT('h4)
	) name10280 (
		_w10810_,
		_w10811_,
		_w10812_
	);
	LUT2 #(
		.INIT('h1)
	) name10281 (
		\text_in_r_reg[69]/P0001 ,
		\u0_w_reg[1][5]/P0001 ,
		_w10813_
	);
	LUT2 #(
		.INIT('h8)
	) name10282 (
		\text_in_r_reg[69]/P0001 ,
		\u0_w_reg[1][5]/P0001 ,
		_w10814_
	);
	LUT2 #(
		.INIT('h2)
	) name10283 (
		\ld_r_reg/P0001 ,
		_w10813_,
		_w10815_
	);
	LUT2 #(
		.INIT('h4)
	) name10284 (
		_w10814_,
		_w10815_,
		_w10816_
	);
	LUT2 #(
		.INIT('h1)
	) name10285 (
		_w10812_,
		_w10816_,
		_w10817_
	);
	LUT2 #(
		.INIT('h1)
	) name10286 (
		_w9639_,
		_w10430_,
		_w10818_
	);
	LUT2 #(
		.INIT('h8)
	) name10287 (
		_w9639_,
		_w10430_,
		_w10819_
	);
	LUT2 #(
		.INIT('h1)
	) name10288 (
		_w10818_,
		_w10819_,
		_w10820_
	);
	LUT2 #(
		.INIT('h8)
	) name10289 (
		\sa30_reg[7]/P0001 ,
		_w8821_,
		_w10821_
	);
	LUT2 #(
		.INIT('h4)
	) name10290 (
		\sa30_reg[3]/P0001 ,
		_w8706_,
		_w10822_
	);
	LUT2 #(
		.INIT('h1)
	) name10291 (
		_w8748_,
		_w10822_,
		_w10823_
	);
	LUT2 #(
		.INIT('h2)
	) name10292 (
		\sa30_reg[2]/P0001 ,
		_w10823_,
		_w10824_
	);
	LUT2 #(
		.INIT('h8)
	) name10293 (
		_w8692_,
		_w9582_,
		_w10825_
	);
	LUT2 #(
		.INIT('h2)
	) name10294 (
		\sa30_reg[1]/P0001 ,
		_w8796_,
		_w10826_
	);
	LUT2 #(
		.INIT('h4)
	) name10295 (
		_w8720_,
		_w10826_,
		_w10827_
	);
	LUT2 #(
		.INIT('h1)
	) name10296 (
		_w10821_,
		_w10825_,
		_w10828_
	);
	LUT2 #(
		.INIT('h8)
	) name10297 (
		_w10827_,
		_w10828_,
		_w10829_
	);
	LUT2 #(
		.INIT('h4)
	) name10298 (
		_w10824_,
		_w10829_,
		_w10830_
	);
	LUT2 #(
		.INIT('h8)
	) name10299 (
		_w8701_,
		_w8811_,
		_w10831_
	);
	LUT2 #(
		.INIT('h2)
	) name10300 (
		\sa30_reg[7]/P0001 ,
		_w8775_,
		_w10832_
	);
	LUT2 #(
		.INIT('h8)
	) name10301 (
		_w8929_,
		_w10832_,
		_w10833_
	);
	LUT2 #(
		.INIT('h1)
	) name10302 (
		\sa30_reg[1]/P0001 ,
		_w8875_,
		_w10834_
	);
	LUT2 #(
		.INIT('h4)
	) name10303 (
		_w10831_,
		_w10834_,
		_w10835_
	);
	LUT2 #(
		.INIT('h1)
	) name10304 (
		_w10357_,
		_w10833_,
		_w10836_
	);
	LUT2 #(
		.INIT('h8)
	) name10305 (
		_w10835_,
		_w10836_,
		_w10837_
	);
	LUT2 #(
		.INIT('h4)
	) name10306 (
		_w8941_,
		_w10837_,
		_w10838_
	);
	LUT2 #(
		.INIT('h1)
	) name10307 (
		_w10830_,
		_w10838_,
		_w10839_
	);
	LUT2 #(
		.INIT('h1)
	) name10308 (
		\sa30_reg[2]/P0001 ,
		_w8890_,
		_w10840_
	);
	LUT2 #(
		.INIT('h1)
	) name10309 (
		_w8839_,
		_w8952_,
		_w10841_
	);
	LUT2 #(
		.INIT('h2)
	) name10310 (
		\sa30_reg[2]/P0001 ,
		_w10841_,
		_w10842_
	);
	LUT2 #(
		.INIT('h1)
	) name10311 (
		_w8768_,
		_w10840_,
		_w10843_
	);
	LUT2 #(
		.INIT('h4)
	) name10312 (
		_w10842_,
		_w10843_,
		_w10844_
	);
	LUT2 #(
		.INIT('h4)
	) name10313 (
		_w10839_,
		_w10844_,
		_w10845_
	);
	LUT2 #(
		.INIT('h1)
	) name10314 (
		\sa30_reg[0]/P0002 ,
		_w10845_,
		_w10846_
	);
	LUT2 #(
		.INIT('h1)
	) name10315 (
		_w8835_,
		_w8950_,
		_w10847_
	);
	LUT2 #(
		.INIT('h1)
	) name10316 (
		\sa30_reg[2]/P0001 ,
		_w10847_,
		_w10848_
	);
	LUT2 #(
		.INIT('h8)
	) name10317 (
		\sa30_reg[4]/P0001 ,
		_w10295_,
		_w10849_
	);
	LUT2 #(
		.INIT('h1)
	) name10318 (
		_w8692_,
		_w8884_,
		_w10850_
	);
	LUT2 #(
		.INIT('h4)
	) name10319 (
		_w9547_,
		_w10850_,
		_w10851_
	);
	LUT2 #(
		.INIT('h2)
	) name10320 (
		\sa30_reg[2]/P0001 ,
		_w10851_,
		_w10852_
	);
	LUT2 #(
		.INIT('h1)
	) name10321 (
		_w9596_,
		_w10849_,
		_w10853_
	);
	LUT2 #(
		.INIT('h4)
	) name10322 (
		_w10848_,
		_w10853_,
		_w10854_
	);
	LUT2 #(
		.INIT('h4)
	) name10323 (
		_w10852_,
		_w10854_,
		_w10855_
	);
	LUT2 #(
		.INIT('h2)
	) name10324 (
		\sa30_reg[1]/P0001 ,
		_w10855_,
		_w10856_
	);
	LUT2 #(
		.INIT('h4)
	) name10325 (
		_w8875_,
		_w10291_,
		_w10857_
	);
	LUT2 #(
		.INIT('h1)
	) name10326 (
		\sa30_reg[2]/P0001 ,
		_w10857_,
		_w10858_
	);
	LUT2 #(
		.INIT('h4)
	) name10327 (
		_w8683_,
		_w8815_,
		_w10859_
	);
	LUT2 #(
		.INIT('h2)
	) name10328 (
		_w8811_,
		_w10859_,
		_w10860_
	);
	LUT2 #(
		.INIT('h1)
	) name10329 (
		_w8705_,
		_w8757_,
		_w10861_
	);
	LUT2 #(
		.INIT('h8)
	) name10330 (
		_w9592_,
		_w10861_,
		_w10862_
	);
	LUT2 #(
		.INIT('h1)
	) name10331 (
		_w9633_,
		_w10862_,
		_w10863_
	);
	LUT2 #(
		.INIT('h8)
	) name10332 (
		_w8775_,
		_w8896_,
		_w10864_
	);
	LUT2 #(
		.INIT('h1)
	) name10333 (
		_w8699_,
		_w8810_,
		_w10865_
	);
	LUT2 #(
		.INIT('h4)
	) name10334 (
		_w8834_,
		_w10865_,
		_w10866_
	);
	LUT2 #(
		.INIT('h4)
	) name10335 (
		_w10864_,
		_w10866_,
		_w10867_
	);
	LUT2 #(
		.INIT('h4)
	) name10336 (
		_w10863_,
		_w10867_,
		_w10868_
	);
	LUT2 #(
		.INIT('h1)
	) name10337 (
		\sa30_reg[1]/P0001 ,
		_w10868_,
		_w10869_
	);
	LUT2 #(
		.INIT('h1)
	) name10338 (
		_w8764_,
		_w10860_,
		_w10870_
	);
	LUT2 #(
		.INIT('h4)
	) name10339 (
		_w10858_,
		_w10870_,
		_w10871_
	);
	LUT2 #(
		.INIT('h4)
	) name10340 (
		_w10856_,
		_w10871_,
		_w10872_
	);
	LUT2 #(
		.INIT('h4)
	) name10341 (
		_w10869_,
		_w10872_,
		_w10873_
	);
	LUT2 #(
		.INIT('h2)
	) name10342 (
		\sa30_reg[0]/P0002 ,
		_w10873_,
		_w10874_
	);
	LUT2 #(
		.INIT('h4)
	) name10343 (
		\sa30_reg[2]/P0001 ,
		_w9608_,
		_w10875_
	);
	LUT2 #(
		.INIT('h1)
	) name10344 (
		_w8687_,
		_w10389_,
		_w10876_
	);
	LUT2 #(
		.INIT('h4)
	) name10345 (
		_w8693_,
		_w10876_,
		_w10877_
	);
	LUT2 #(
		.INIT('h2)
	) name10346 (
		_w8833_,
		_w10877_,
		_w10878_
	);
	LUT2 #(
		.INIT('h8)
	) name10347 (
		_w8710_,
		_w8844_,
		_w10879_
	);
	LUT2 #(
		.INIT('h8)
	) name10348 (
		_w8697_,
		_w10297_,
		_w10880_
	);
	LUT2 #(
		.INIT('h1)
	) name10349 (
		_w9585_,
		_w10879_,
		_w10881_
	);
	LUT2 #(
		.INIT('h4)
	) name10350 (
		_w10880_,
		_w10881_,
		_w10882_
	);
	LUT2 #(
		.INIT('h4)
	) name10351 (
		_w10875_,
		_w10882_,
		_w10883_
	);
	LUT2 #(
		.INIT('h4)
	) name10352 (
		_w10878_,
		_w10883_,
		_w10884_
	);
	LUT2 #(
		.INIT('h2)
	) name10353 (
		\sa30_reg[1]/P0001 ,
		_w10884_,
		_w10885_
	);
	LUT2 #(
		.INIT('h1)
	) name10354 (
		_w8768_,
		_w8784_,
		_w10886_
	);
	LUT2 #(
		.INIT('h2)
	) name10355 (
		\sa30_reg[2]/P0001 ,
		_w10886_,
		_w10887_
	);
	LUT2 #(
		.INIT('h8)
	) name10356 (
		\sa30_reg[7]/P0001 ,
		_w8758_,
		_w10888_
	);
	LUT2 #(
		.INIT('h8)
	) name10357 (
		_w9582_,
		_w10888_,
		_w10889_
	);
	LUT2 #(
		.INIT('h1)
	) name10358 (
		_w10887_,
		_w10889_,
		_w10890_
	);
	LUT2 #(
		.INIT('h1)
	) name10359 (
		\sa30_reg[1]/P0001 ,
		_w10890_,
		_w10891_
	);
	LUT2 #(
		.INIT('h1)
	) name10360 (
		_w8744_,
		_w9572_,
		_w10892_
	);
	LUT2 #(
		.INIT('h2)
	) name10361 (
		_w8844_,
		_w10892_,
		_w10893_
	);
	LUT2 #(
		.INIT('h1)
	) name10362 (
		_w8956_,
		_w10893_,
		_w10894_
	);
	LUT2 #(
		.INIT('h4)
	) name10363 (
		_w10891_,
		_w10894_,
		_w10895_
	);
	LUT2 #(
		.INIT('h4)
	) name10364 (
		_w10885_,
		_w10895_,
		_w10896_
	);
	LUT2 #(
		.INIT('h4)
	) name10365 (
		_w10846_,
		_w10896_,
		_w10897_
	);
	LUT2 #(
		.INIT('h4)
	) name10366 (
		_w10874_,
		_w10897_,
		_w10898_
	);
	LUT2 #(
		.INIT('h2)
	) name10367 (
		\u0_w_reg[1][12]/P0001 ,
		_w10898_,
		_w10899_
	);
	LUT2 #(
		.INIT('h4)
	) name10368 (
		\u0_w_reg[1][12]/P0001 ,
		_w10898_,
		_w10900_
	);
	LUT2 #(
		.INIT('h1)
	) name10369 (
		_w10899_,
		_w10900_,
		_w10901_
	);
	LUT2 #(
		.INIT('h8)
	) name10370 (
		_w10820_,
		_w10901_,
		_w10902_
	);
	LUT2 #(
		.INIT('h1)
	) name10371 (
		_w10820_,
		_w10901_,
		_w10903_
	);
	LUT2 #(
		.INIT('h1)
	) name10372 (
		_w10902_,
		_w10903_,
		_w10904_
	);
	LUT2 #(
		.INIT('h2)
	) name10373 (
		_w9980_,
		_w10775_,
		_w10905_
	);
	LUT2 #(
		.INIT('h4)
	) name10374 (
		_w9980_,
		_w10775_,
		_w10906_
	);
	LUT2 #(
		.INIT('h1)
	) name10375 (
		_w10905_,
		_w10906_,
		_w10907_
	);
	LUT2 #(
		.INIT('h4)
	) name10376 (
		_w8379_,
		_w10907_,
		_w10908_
	);
	LUT2 #(
		.INIT('h2)
	) name10377 (
		_w8379_,
		_w10907_,
		_w10909_
	);
	LUT2 #(
		.INIT('h1)
	) name10378 (
		_w10908_,
		_w10909_,
		_w10910_
	);
	LUT2 #(
		.INIT('h1)
	) name10379 (
		_w10904_,
		_w10910_,
		_w10911_
	);
	LUT2 #(
		.INIT('h8)
	) name10380 (
		_w10904_,
		_w10910_,
		_w10912_
	);
	LUT2 #(
		.INIT('h1)
	) name10381 (
		\ld_r_reg/P0001 ,
		_w10911_,
		_w10913_
	);
	LUT2 #(
		.INIT('h4)
	) name10382 (
		_w10912_,
		_w10913_,
		_w10914_
	);
	LUT2 #(
		.INIT('h2)
	) name10383 (
		\text_in_r_reg[76]/P0001 ,
		\u0_w_reg[1][12]/P0001 ,
		_w10915_
	);
	LUT2 #(
		.INIT('h4)
	) name10384 (
		\text_in_r_reg[76]/P0001 ,
		\u0_w_reg[1][12]/P0001 ,
		_w10916_
	);
	LUT2 #(
		.INIT('h2)
	) name10385 (
		\ld_r_reg/P0001 ,
		_w10915_,
		_w10917_
	);
	LUT2 #(
		.INIT('h4)
	) name10386 (
		_w10916_,
		_w10917_,
		_w10918_
	);
	LUT2 #(
		.INIT('h1)
	) name10387 (
		_w10914_,
		_w10918_,
		_w10919_
	);
	LUT2 #(
		.INIT('h1)
	) name10388 (
		\sa12_reg[2]/P0001 ,
		_w8077_,
		_w10920_
	);
	LUT2 #(
		.INIT('h1)
	) name10389 (
		\sa12_reg[5]/P0001 ,
		_w8055_,
		_w10921_
	);
	LUT2 #(
		.INIT('h2)
	) name10390 (
		_w10920_,
		_w10921_,
		_w10922_
	);
	LUT2 #(
		.INIT('h1)
	) name10391 (
		_w9049_,
		_w10922_,
		_w10923_
	);
	LUT2 #(
		.INIT('h2)
	) name10392 (
		\sa12_reg[1]/P0001 ,
		_w10923_,
		_w10924_
	);
	LUT2 #(
		.INIT('h1)
	) name10393 (
		_w8093_,
		_w8498_,
		_w10925_
	);
	LUT2 #(
		.INIT('h2)
	) name10394 (
		\sa12_reg[3]/P0001 ,
		_w10925_,
		_w10926_
	);
	LUT2 #(
		.INIT('h1)
	) name10395 (
		_w8432_,
		_w8494_,
		_w10927_
	);
	LUT2 #(
		.INIT('h4)
	) name10396 (
		_w10926_,
		_w10927_,
		_w10928_
	);
	LUT2 #(
		.INIT('h1)
	) name10397 (
		\sa12_reg[2]/P0001 ,
		_w10928_,
		_w10929_
	);
	LUT2 #(
		.INIT('h1)
	) name10398 (
		_w8184_,
		_w8985_,
		_w10930_
	);
	LUT2 #(
		.INIT('h8)
	) name10399 (
		_w8462_,
		_w10930_,
		_w10931_
	);
	LUT2 #(
		.INIT('h2)
	) name10400 (
		\sa12_reg[2]/P0001 ,
		_w10931_,
		_w10932_
	);
	LUT2 #(
		.INIT('h8)
	) name10401 (
		_w8147_,
		_w8978_,
		_w10933_
	);
	LUT2 #(
		.INIT('h2)
	) name10402 (
		\sa12_reg[5]/P0001 ,
		_w8126_,
		_w10934_
	);
	LUT2 #(
		.INIT('h2)
	) name10403 (
		_w8078_,
		_w10934_,
		_w10935_
	);
	LUT2 #(
		.INIT('h8)
	) name10404 (
		_w8074_,
		_w8104_,
		_w10936_
	);
	LUT2 #(
		.INIT('h4)
	) name10405 (
		\sa12_reg[3]/P0001 ,
		_w8142_,
		_w10937_
	);
	LUT2 #(
		.INIT('h1)
	) name10406 (
		_w8391_,
		_w8452_,
		_w10938_
	);
	LUT2 #(
		.INIT('h4)
	) name10407 (
		_w10937_,
		_w10938_,
		_w10939_
	);
	LUT2 #(
		.INIT('h2)
	) name10408 (
		\sa12_reg[2]/P0001 ,
		_w10939_,
		_w10940_
	);
	LUT2 #(
		.INIT('h1)
	) name10409 (
		_w10933_,
		_w10936_,
		_w10941_
	);
	LUT2 #(
		.INIT('h4)
	) name10410 (
		_w10935_,
		_w10941_,
		_w10942_
	);
	LUT2 #(
		.INIT('h4)
	) name10411 (
		_w10940_,
		_w10942_,
		_w10943_
	);
	LUT2 #(
		.INIT('h1)
	) name10412 (
		\sa12_reg[1]/P0001 ,
		_w10943_,
		_w10944_
	);
	LUT2 #(
		.INIT('h1)
	) name10413 (
		_w8113_,
		_w8175_,
		_w10945_
	);
	LUT2 #(
		.INIT('h4)
	) name10414 (
		_w10924_,
		_w10945_,
		_w10946_
	);
	LUT2 #(
		.INIT('h4)
	) name10415 (
		_w10929_,
		_w10946_,
		_w10947_
	);
	LUT2 #(
		.INIT('h4)
	) name10416 (
		_w10932_,
		_w10947_,
		_w10948_
	);
	LUT2 #(
		.INIT('h4)
	) name10417 (
		_w10944_,
		_w10948_,
		_w10949_
	);
	LUT2 #(
		.INIT('h2)
	) name10418 (
		\sa12_reg[0]/P0001 ,
		_w10949_,
		_w10950_
	);
	LUT2 #(
		.INIT('h8)
	) name10419 (
		\sa12_reg[2]/P0001 ,
		_w8076_,
		_w10951_
	);
	LUT2 #(
		.INIT('h8)
	) name10420 (
		_w8075_,
		_w8080_,
		_w10952_
	);
	LUT2 #(
		.INIT('h2)
	) name10421 (
		\sa12_reg[1]/P0001 ,
		_w8417_,
		_w10953_
	);
	LUT2 #(
		.INIT('h1)
	) name10422 (
		_w9817_,
		_w9821_,
		_w10954_
	);
	LUT2 #(
		.INIT('h4)
	) name10423 (
		_w10952_,
		_w10954_,
		_w10955_
	);
	LUT2 #(
		.INIT('h4)
	) name10424 (
		_w10951_,
		_w10953_,
		_w10956_
	);
	LUT2 #(
		.INIT('h8)
	) name10425 (
		_w10955_,
		_w10956_,
		_w10957_
	);
	LUT2 #(
		.INIT('h2)
	) name10426 (
		\sa12_reg[2]/P0001 ,
		_w8075_,
		_w10958_
	);
	LUT2 #(
		.INIT('h8)
	) name10427 (
		_w8161_,
		_w10958_,
		_w10959_
	);
	LUT2 #(
		.INIT('h1)
	) name10428 (
		\sa12_reg[3]/P0001 ,
		_w9784_,
		_w10960_
	);
	LUT2 #(
		.INIT('h2)
	) name10429 (
		_w8158_,
		_w10959_,
		_w10961_
	);
	LUT2 #(
		.INIT('h4)
	) name10430 (
		_w10960_,
		_w10961_,
		_w10962_
	);
	LUT2 #(
		.INIT('h1)
	) name10431 (
		_w10957_,
		_w10962_,
		_w10963_
	);
	LUT2 #(
		.INIT('h1)
	) name10432 (
		_w8056_,
		_w8093_,
		_w10964_
	);
	LUT2 #(
		.INIT('h2)
	) name10433 (
		_w8078_,
		_w10964_,
		_w10965_
	);
	LUT2 #(
		.INIT('h2)
	) name10434 (
		\sa12_reg[2]/P0001 ,
		_w10965_,
		_w10966_
	);
	LUT2 #(
		.INIT('h1)
	) name10435 (
		\sa12_reg[2]/P0001 ,
		_w8117_,
		_w10967_
	);
	LUT2 #(
		.INIT('h8)
	) name10436 (
		_w10641_,
		_w10967_,
		_w10968_
	);
	LUT2 #(
		.INIT('h1)
	) name10437 (
		_w10966_,
		_w10968_,
		_w10969_
	);
	LUT2 #(
		.INIT('h1)
	) name10438 (
		_w10963_,
		_w10969_,
		_w10970_
	);
	LUT2 #(
		.INIT('h1)
	) name10439 (
		\sa12_reg[0]/P0001 ,
		_w10970_,
		_w10971_
	);
	LUT2 #(
		.INIT('h1)
	) name10440 (
		_w8086_,
		_w8394_,
		_w10972_
	);
	LUT2 #(
		.INIT('h2)
	) name10441 (
		_w10064_,
		_w10972_,
		_w10973_
	);
	LUT2 #(
		.INIT('h8)
	) name10442 (
		_w8059_,
		_w8174_,
		_w10974_
	);
	LUT2 #(
		.INIT('h1)
	) name10443 (
		_w10952_,
		_w10974_,
		_w10975_
	);
	LUT2 #(
		.INIT('h1)
	) name10444 (
		_w8066_,
		_w10975_,
		_w10976_
	);
	LUT2 #(
		.INIT('h1)
	) name10445 (
		\sa12_reg[2]/P0001 ,
		_w9865_,
		_w10977_
	);
	LUT2 #(
		.INIT('h1)
	) name10446 (
		_w8128_,
		_w10977_,
		_w10978_
	);
	LUT2 #(
		.INIT('h8)
	) name10447 (
		_w8066_,
		_w8413_,
		_w10979_
	);
	LUT2 #(
		.INIT('h1)
	) name10448 (
		_w8118_,
		_w8150_,
		_w10980_
	);
	LUT2 #(
		.INIT('h4)
	) name10449 (
		_w10978_,
		_w10980_,
		_w10981_
	);
	LUT2 #(
		.INIT('h4)
	) name10450 (
		_w10979_,
		_w10981_,
		_w10982_
	);
	LUT2 #(
		.INIT('h2)
	) name10451 (
		\sa12_reg[1]/P0001 ,
		_w10982_,
		_w10983_
	);
	LUT2 #(
		.INIT('h8)
	) name10452 (
		_w8074_,
		_w8155_,
		_w10984_
	);
	LUT2 #(
		.INIT('h8)
	) name10453 (
		_w8068_,
		_w10984_,
		_w10985_
	);
	LUT2 #(
		.INIT('h1)
	) name10454 (
		_w8061_,
		_w8412_,
		_w10986_
	);
	LUT2 #(
		.INIT('h4)
	) name10455 (
		_w9790_,
		_w10986_,
		_w10987_
	);
	LUT2 #(
		.INIT('h2)
	) name10456 (
		_w8978_,
		_w10987_,
		_w10988_
	);
	LUT2 #(
		.INIT('h1)
	) name10457 (
		_w8491_,
		_w10985_,
		_w10989_
	);
	LUT2 #(
		.INIT('h4)
	) name10458 (
		_w10988_,
		_w10989_,
		_w10990_
	);
	LUT2 #(
		.INIT('h1)
	) name10459 (
		\sa12_reg[1]/P0001 ,
		_w10990_,
		_w10991_
	);
	LUT2 #(
		.INIT('h1)
	) name10460 (
		_w10973_,
		_w10976_,
		_w10992_
	);
	LUT2 #(
		.INIT('h4)
	) name10461 (
		_w10983_,
		_w10992_,
		_w10993_
	);
	LUT2 #(
		.INIT('h4)
	) name10462 (
		_w10991_,
		_w10993_,
		_w10994_
	);
	LUT2 #(
		.INIT('h4)
	) name10463 (
		_w10971_,
		_w10994_,
		_w10995_
	);
	LUT2 #(
		.INIT('h4)
	) name10464 (
		_w10950_,
		_w10995_,
		_w10996_
	);
	LUT2 #(
		.INIT('h2)
	) name10465 (
		_w9874_,
		_w10996_,
		_w10997_
	);
	LUT2 #(
		.INIT('h4)
	) name10466 (
		_w9874_,
		_w10996_,
		_w10998_
	);
	LUT2 #(
		.INIT('h1)
	) name10467 (
		_w10997_,
		_w10998_,
		_w10999_
	);
	LUT2 #(
		.INIT('h1)
	) name10468 (
		_w8521_,
		_w9489_,
		_w11000_
	);
	LUT2 #(
		.INIT('h2)
	) name10469 (
		\sa23_reg[1]/P0001 ,
		_w11000_,
		_w11001_
	);
	LUT2 #(
		.INIT('h1)
	) name10470 (
		_w8525_,
		_w8577_,
		_w11002_
	);
	LUT2 #(
		.INIT('h2)
	) name10471 (
		\sa23_reg[3]/P0001 ,
		_w11002_,
		_w11003_
	);
	LUT2 #(
		.INIT('h1)
	) name10472 (
		_w9899_,
		_w9938_,
		_w11004_
	);
	LUT2 #(
		.INIT('h4)
	) name10473 (
		_w11003_,
		_w11004_,
		_w11005_
	);
	LUT2 #(
		.INIT('h4)
	) name10474 (
		_w11001_,
		_w11005_,
		_w11006_
	);
	LUT2 #(
		.INIT('h1)
	) name10475 (
		\sa23_reg[2]/P0001 ,
		_w11006_,
		_w11007_
	);
	LUT2 #(
		.INIT('h1)
	) name10476 (
		_w9078_,
		_w9498_,
		_w11008_
	);
	LUT2 #(
		.INIT('h8)
	) name10477 (
		_w8634_,
		_w11008_,
		_w11009_
	);
	LUT2 #(
		.INIT('h2)
	) name10478 (
		\sa23_reg[2]/P0001 ,
		_w11009_,
		_w11010_
	);
	LUT2 #(
		.INIT('h8)
	) name10479 (
		\sa23_reg[1]/P0001 ,
		_w9152_,
		_w11011_
	);
	LUT2 #(
		.INIT('h8)
	) name10480 (
		\sa23_reg[4]/P0001 ,
		_w9894_,
		_w11012_
	);
	LUT2 #(
		.INIT('h2)
	) name10481 (
		\sa23_reg[5]/P0001 ,
		_w8511_,
		_w11013_
	);
	LUT2 #(
		.INIT('h2)
	) name10482 (
		_w8572_,
		_w11013_,
		_w11014_
	);
	LUT2 #(
		.INIT('h1)
	) name10483 (
		_w8534_,
		_w8602_,
		_w11015_
	);
	LUT2 #(
		.INIT('h4)
	) name10484 (
		_w9128_,
		_w11015_,
		_w11016_
	);
	LUT2 #(
		.INIT('h2)
	) name10485 (
		\sa23_reg[2]/P0001 ,
		_w11016_,
		_w11017_
	);
	LUT2 #(
		.INIT('h1)
	) name10486 (
		_w9943_,
		_w11014_,
		_w11018_
	);
	LUT2 #(
		.INIT('h4)
	) name10487 (
		_w11012_,
		_w11018_,
		_w11019_
	);
	LUT2 #(
		.INIT('h4)
	) name10488 (
		_w11017_,
		_w11019_,
		_w11020_
	);
	LUT2 #(
		.INIT('h1)
	) name10489 (
		\sa23_reg[1]/P0001 ,
		_w11020_,
		_w11021_
	);
	LUT2 #(
		.INIT('h1)
	) name10490 (
		_w9454_,
		_w9492_,
		_w11022_
	);
	LUT2 #(
		.INIT('h4)
	) name10491 (
		_w11011_,
		_w11022_,
		_w11023_
	);
	LUT2 #(
		.INIT('h4)
	) name10492 (
		_w11010_,
		_w11023_,
		_w11024_
	);
	LUT2 #(
		.INIT('h4)
	) name10493 (
		_w11007_,
		_w11024_,
		_w11025_
	);
	LUT2 #(
		.INIT('h4)
	) name10494 (
		_w11021_,
		_w11025_,
		_w11026_
	);
	LUT2 #(
		.INIT('h2)
	) name10495 (
		\sa23_reg[0]/P0001 ,
		_w11026_,
		_w11027_
	);
	LUT2 #(
		.INIT('h4)
	) name10496 (
		_w9106_,
		_w10719_,
		_w11028_
	);
	LUT2 #(
		.INIT('h1)
	) name10497 (
		\sa23_reg[2]/P0001 ,
		_w11028_,
		_w11029_
	);
	LUT2 #(
		.INIT('h1)
	) name10498 (
		_w8525_,
		_w8631_,
		_w11030_
	);
	LUT2 #(
		.INIT('h2)
	) name10499 (
		_w9897_,
		_w11030_,
		_w11031_
	);
	LUT2 #(
		.INIT('h2)
	) name10500 (
		_w8531_,
		_w8588_,
		_w11032_
	);
	LUT2 #(
		.INIT('h8)
	) name10501 (
		_w9958_,
		_w11032_,
		_w11033_
	);
	LUT2 #(
		.INIT('h1)
	) name10502 (
		\sa23_reg[3]/P0001 ,
		_w9965_,
		_w11034_
	);
	LUT2 #(
		.INIT('h2)
	) name10503 (
		_w9432_,
		_w11034_,
		_w11035_
	);
	LUT2 #(
		.INIT('h8)
	) name10504 (
		_w8562_,
		_w9079_,
		_w11036_
	);
	LUT2 #(
		.INIT('h8)
	) name10505 (
		_w8569_,
		_w8588_,
		_w11037_
	);
	LUT2 #(
		.INIT('h8)
	) name10506 (
		_w8546_,
		_w8614_,
		_w11038_
	);
	LUT2 #(
		.INIT('h2)
	) name10507 (
		_w8528_,
		_w8537_,
		_w11039_
	);
	LUT2 #(
		.INIT('h2)
	) name10508 (
		\sa23_reg[1]/P0001 ,
		_w11036_,
		_w11040_
	);
	LUT2 #(
		.INIT('h1)
	) name10509 (
		_w11037_,
		_w11039_,
		_w11041_
	);
	LUT2 #(
		.INIT('h8)
	) name10510 (
		_w11040_,
		_w11041_,
		_w11042_
	);
	LUT2 #(
		.INIT('h4)
	) name10511 (
		_w11038_,
		_w11042_,
		_w11043_
	);
	LUT2 #(
		.INIT('h1)
	) name10512 (
		_w11035_,
		_w11043_,
		_w11044_
	);
	LUT2 #(
		.INIT('h1)
	) name10513 (
		_w11031_,
		_w11033_,
		_w11045_
	);
	LUT2 #(
		.INIT('h4)
	) name10514 (
		_w11029_,
		_w11045_,
		_w11046_
	);
	LUT2 #(
		.INIT('h4)
	) name10515 (
		_w11044_,
		_w11046_,
		_w11047_
	);
	LUT2 #(
		.INIT('h1)
	) name10516 (
		\sa23_reg[0]/P0001 ,
		_w11047_,
		_w11048_
	);
	LUT2 #(
		.INIT('h1)
	) name10517 (
		_w8574_,
		_w8642_,
		_w11049_
	);
	LUT2 #(
		.INIT('h4)
	) name10518 (
		_w10730_,
		_w11049_,
		_w11050_
	);
	LUT2 #(
		.INIT('h1)
	) name10519 (
		\sa23_reg[7]/NET0131 ,
		_w11050_,
		_w11051_
	);
	LUT2 #(
		.INIT('h1)
	) name10520 (
		_w9464_,
		_w11051_,
		_w11052_
	);
	LUT2 #(
		.INIT('h1)
	) name10521 (
		\sa23_reg[2]/P0001 ,
		_w11052_,
		_w11053_
	);
	LUT2 #(
		.INIT('h1)
	) name10522 (
		_w8521_,
		_w8654_,
		_w11054_
	);
	LUT2 #(
		.INIT('h8)
	) name10523 (
		\sa23_reg[2]/P0001 ,
		_w8522_,
		_w11055_
	);
	LUT2 #(
		.INIT('h4)
	) name10524 (
		_w11054_,
		_w11055_,
		_w11056_
	);
	LUT2 #(
		.INIT('h1)
	) name10525 (
		_w8668_,
		_w11056_,
		_w11057_
	);
	LUT2 #(
		.INIT('h4)
	) name10526 (
		_w11053_,
		_w11057_,
		_w11058_
	);
	LUT2 #(
		.INIT('h1)
	) name10527 (
		\sa23_reg[1]/P0001 ,
		_w11058_,
		_w11059_
	);
	LUT2 #(
		.INIT('h8)
	) name10528 (
		_w9112_,
		_w9152_,
		_w11060_
	);
	LUT2 #(
		.INIT('h1)
	) name10529 (
		\sa23_reg[2]/P0001 ,
		_w8619_,
		_w11061_
	);
	LUT2 #(
		.INIT('h1)
	) name10530 (
		_w9438_,
		_w11061_,
		_w11062_
	);
	LUT2 #(
		.INIT('h1)
	) name10531 (
		_w8609_,
		_w9137_,
		_w11063_
	);
	LUT2 #(
		.INIT('h4)
	) name10532 (
		_w11060_,
		_w11063_,
		_w11064_
	);
	LUT2 #(
		.INIT('h4)
	) name10533 (
		_w11062_,
		_w11064_,
		_w11065_
	);
	LUT2 #(
		.INIT('h2)
	) name10534 (
		\sa23_reg[1]/P0001 ,
		_w11065_,
		_w11066_
	);
	LUT2 #(
		.INIT('h8)
	) name10535 (
		\sa23_reg[2]/P0001 ,
		_w8524_,
		_w11067_
	);
	LUT2 #(
		.INIT('h4)
	) name10536 (
		\sa23_reg[2]/P0001 ,
		_w11037_,
		_w11068_
	);
	LUT2 #(
		.INIT('h1)
	) name10537 (
		_w11067_,
		_w11068_,
		_w11069_
	);
	LUT2 #(
		.INIT('h4)
	) name10538 (
		_w11066_,
		_w11069_,
		_w11070_
	);
	LUT2 #(
		.INIT('h4)
	) name10539 (
		_w11048_,
		_w11070_,
		_w11071_
	);
	LUT2 #(
		.INIT('h4)
	) name10540 (
		_w11059_,
		_w11071_,
		_w11072_
	);
	LUT2 #(
		.INIT('h4)
	) name10541 (
		_w11027_,
		_w11072_,
		_w11073_
	);
	LUT2 #(
		.INIT('h2)
	) name10542 (
		_w10167_,
		_w11073_,
		_w11074_
	);
	LUT2 #(
		.INIT('h4)
	) name10543 (
		_w10167_,
		_w11073_,
		_w11075_
	);
	LUT2 #(
		.INIT('h1)
	) name10544 (
		_w11074_,
		_w11075_,
		_w11076_
	);
	LUT2 #(
		.INIT('h8)
	) name10545 (
		_w10999_,
		_w11076_,
		_w11077_
	);
	LUT2 #(
		.INIT('h1)
	) name10546 (
		_w10999_,
		_w11076_,
		_w11078_
	);
	LUT2 #(
		.INIT('h1)
	) name10547 (
		_w11077_,
		_w11078_,
		_w11079_
	);
	LUT2 #(
		.INIT('h1)
	) name10548 (
		_w8744_,
		_w10821_,
		_w11080_
	);
	LUT2 #(
		.INIT('h1)
	) name10549 (
		_w9614_,
		_w10375_,
		_w11081_
	);
	LUT2 #(
		.INIT('h4)
	) name10550 (
		_w10888_,
		_w11081_,
		_w11082_
	);
	LUT2 #(
		.INIT('h2)
	) name10551 (
		\sa30_reg[2]/P0001 ,
		_w11082_,
		_w11083_
	);
	LUT2 #(
		.INIT('h2)
	) name10552 (
		_w11080_,
		_w11083_,
		_w11084_
	);
	LUT2 #(
		.INIT('h2)
	) name10553 (
		\sa30_reg[1]/P0001 ,
		_w11084_,
		_w11085_
	);
	LUT2 #(
		.INIT('h2)
	) name10554 (
		_w8710_,
		_w9582_,
		_w11086_
	);
	LUT2 #(
		.INIT('h1)
	) name10555 (
		_w10351_,
		_w11086_,
		_w11087_
	);
	LUT2 #(
		.INIT('h1)
	) name10556 (
		\sa30_reg[3]/P0001 ,
		_w11087_,
		_w11088_
	);
	LUT2 #(
		.INIT('h1)
	) name10557 (
		_w8767_,
		_w10279_,
		_w11089_
	);
	LUT2 #(
		.INIT('h1)
	) name10558 (
		_w10351_,
		_w10363_,
		_w11090_
	);
	LUT2 #(
		.INIT('h8)
	) name10559 (
		_w11089_,
		_w11090_,
		_w11091_
	);
	LUT2 #(
		.INIT('h1)
	) name10560 (
		\sa30_reg[2]/P0001 ,
		_w11091_,
		_w11092_
	);
	LUT2 #(
		.INIT('h2)
	) name10561 (
		_w8683_,
		_w9575_,
		_w11093_
	);
	LUT2 #(
		.INIT('h8)
	) name10562 (
		_w8692_,
		_w8698_,
		_w11094_
	);
	LUT2 #(
		.INIT('h1)
	) name10563 (
		_w8767_,
		_w8780_,
		_w11095_
	);
	LUT2 #(
		.INIT('h4)
	) name10564 (
		_w11093_,
		_w11095_,
		_w11096_
	);
	LUT2 #(
		.INIT('h4)
	) name10565 (
		_w11094_,
		_w11096_,
		_w11097_
	);
	LUT2 #(
		.INIT('h1)
	) name10566 (
		\sa30_reg[1]/P0001 ,
		_w11097_,
		_w11098_
	);
	LUT2 #(
		.INIT('h1)
	) name10567 (
		_w11088_,
		_w11092_,
		_w11099_
	);
	LUT2 #(
		.INIT('h4)
	) name10568 (
		_w11098_,
		_w11099_,
		_w11100_
	);
	LUT2 #(
		.INIT('h4)
	) name10569 (
		_w11085_,
		_w11100_,
		_w11101_
	);
	LUT2 #(
		.INIT('h2)
	) name10570 (
		\sa30_reg[0]/P0002 ,
		_w11101_,
		_w11102_
	);
	LUT2 #(
		.INIT('h2)
	) name10571 (
		_w8710_,
		_w9621_,
		_w11103_
	);
	LUT2 #(
		.INIT('h1)
	) name10572 (
		_w8821_,
		_w11103_,
		_w11104_
	);
	LUT2 #(
		.INIT('h2)
	) name10573 (
		_w8946_,
		_w11104_,
		_w11105_
	);
	LUT2 #(
		.INIT('h1)
	) name10574 (
		_w8749_,
		_w9572_,
		_w11106_
	);
	LUT2 #(
		.INIT('h2)
	) name10575 (
		_w8844_,
		_w11106_,
		_w11107_
	);
	LUT2 #(
		.INIT('h1)
	) name10576 (
		_w8769_,
		_w8810_,
		_w11108_
	);
	LUT2 #(
		.INIT('h4)
	) name10577 (
		_w10256_,
		_w11108_,
		_w11109_
	);
	LUT2 #(
		.INIT('h2)
	) name10578 (
		_w10294_,
		_w11109_,
		_w11110_
	);
	LUT2 #(
		.INIT('h1)
	) name10579 (
		_w8703_,
		_w8883_,
		_w11111_
	);
	LUT2 #(
		.INIT('h4)
	) name10580 (
		_w9565_,
		_w11111_,
		_w11112_
	);
	LUT2 #(
		.INIT('h1)
	) name10581 (
		_w8749_,
		_w8894_,
		_w11113_
	);
	LUT2 #(
		.INIT('h8)
	) name10582 (
		_w11112_,
		_w11113_,
		_w11114_
	);
	LUT2 #(
		.INIT('h2)
	) name10583 (
		_w8772_,
		_w11114_,
		_w11115_
	);
	LUT2 #(
		.INIT('h1)
	) name10584 (
		_w8869_,
		_w9632_,
		_w11116_
	);
	LUT2 #(
		.INIT('h4)
	) name10585 (
		_w8784_,
		_w11116_,
		_w11117_
	);
	LUT2 #(
		.INIT('h1)
	) name10586 (
		\sa30_reg[2]/P0001 ,
		_w11117_,
		_w11118_
	);
	LUT2 #(
		.INIT('h1)
	) name10587 (
		_w8781_,
		_w10864_,
		_w11119_
	);
	LUT2 #(
		.INIT('h4)
	) name10588 (
		_w11118_,
		_w11119_,
		_w11120_
	);
	LUT2 #(
		.INIT('h1)
	) name10589 (
		\sa30_reg[1]/P0001 ,
		_w11120_,
		_w11121_
	);
	LUT2 #(
		.INIT('h8)
	) name10590 (
		\sa30_reg[4]/P0001 ,
		_w10272_,
		_w11122_
	);
	LUT2 #(
		.INIT('h1)
	) name10591 (
		_w8776_,
		_w10255_,
		_w11123_
	);
	LUT2 #(
		.INIT('h4)
	) name10592 (
		_w11122_,
		_w11123_,
		_w11124_
	);
	LUT2 #(
		.INIT('h1)
	) name10593 (
		\sa30_reg[2]/P0001 ,
		_w11124_,
		_w11125_
	);
	LUT2 #(
		.INIT('h1)
	) name10594 (
		_w8930_,
		_w10355_,
		_w11126_
	);
	LUT2 #(
		.INIT('h2)
	) name10595 (
		\sa30_reg[2]/P0001 ,
		_w11126_,
		_w11127_
	);
	LUT2 #(
		.INIT('h2)
	) name10596 (
		\sa30_reg[1]/P0001 ,
		_w8703_,
		_w11128_
	);
	LUT2 #(
		.INIT('h8)
	) name10597 (
		_w8761_,
		_w11128_,
		_w11129_
	);
	LUT2 #(
		.INIT('h4)
	) name10598 (
		_w11125_,
		_w11129_,
		_w11130_
	);
	LUT2 #(
		.INIT('h4)
	) name10599 (
		_w11127_,
		_w11130_,
		_w11131_
	);
	LUT2 #(
		.INIT('h8)
	) name10600 (
		_w8686_,
		_w8929_,
		_w11132_
	);
	LUT2 #(
		.INIT('h8)
	) name10601 (
		\sa30_reg[5]/P0001 ,
		_w11132_,
		_w11133_
	);
	LUT2 #(
		.INIT('h1)
	) name10602 (
		_w8876_,
		_w8961_,
		_w11134_
	);
	LUT2 #(
		.INIT('h1)
	) name10603 (
		\sa30_reg[2]/P0001 ,
		_w11134_,
		_w11135_
	);
	LUT2 #(
		.INIT('h1)
	) name10604 (
		\sa30_reg[1]/P0001 ,
		_w8956_,
		_w11136_
	);
	LUT2 #(
		.INIT('h1)
	) name10605 (
		_w9617_,
		_w10879_,
		_w11137_
	);
	LUT2 #(
		.INIT('h4)
	) name10606 (
		_w11133_,
		_w11137_,
		_w11138_
	);
	LUT2 #(
		.INIT('h8)
	) name10607 (
		_w11136_,
		_w11138_,
		_w11139_
	);
	LUT2 #(
		.INIT('h4)
	) name10608 (
		_w11135_,
		_w11139_,
		_w11140_
	);
	LUT2 #(
		.INIT('h1)
	) name10609 (
		_w11131_,
		_w11140_,
		_w11141_
	);
	LUT2 #(
		.INIT('h4)
	) name10610 (
		_w8786_,
		_w9618_,
		_w11142_
	);
	LUT2 #(
		.INIT('h2)
	) name10611 (
		\sa30_reg[2]/P0001 ,
		_w8943_,
		_w11143_
	);
	LUT2 #(
		.INIT('h4)
	) name10612 (
		_w8951_,
		_w11143_,
		_w11144_
	);
	LUT2 #(
		.INIT('h1)
	) name10613 (
		_w11142_,
		_w11144_,
		_w11145_
	);
	LUT2 #(
		.INIT('h1)
	) name10614 (
		_w8810_,
		_w8847_,
		_w11146_
	);
	LUT2 #(
		.INIT('h4)
	) name10615 (
		_w11145_,
		_w11146_,
		_w11147_
	);
	LUT2 #(
		.INIT('h4)
	) name10616 (
		_w11141_,
		_w11147_,
		_w11148_
	);
	LUT2 #(
		.INIT('h1)
	) name10617 (
		\sa30_reg[0]/P0002 ,
		_w11148_,
		_w11149_
	);
	LUT2 #(
		.INIT('h1)
	) name10618 (
		_w11105_,
		_w11107_,
		_w11150_
	);
	LUT2 #(
		.INIT('h4)
	) name10619 (
		_w11110_,
		_w11150_,
		_w11151_
	);
	LUT2 #(
		.INIT('h4)
	) name10620 (
		_w11115_,
		_w11151_,
		_w11152_
	);
	LUT2 #(
		.INIT('h4)
	) name10621 (
		_w11121_,
		_w11152_,
		_w11153_
	);
	LUT2 #(
		.INIT('h4)
	) name10622 (
		_w11102_,
		_w11153_,
		_w11154_
	);
	LUT2 #(
		.INIT('h4)
	) name10623 (
		_w11149_,
		_w11154_,
		_w11155_
	);
	LUT2 #(
		.INIT('h1)
	) name10624 (
		\u0_w_reg[1][17]/P0001 ,
		_w11155_,
		_w11156_
	);
	LUT2 #(
		.INIT('h8)
	) name10625 (
		\u0_w_reg[1][17]/P0001 ,
		_w11155_,
		_w11157_
	);
	LUT2 #(
		.INIT('h1)
	) name10626 (
		_w11156_,
		_w11157_,
		_w11158_
	);
	LUT2 #(
		.INIT('h2)
	) name10627 (
		_w9980_,
		_w10508_,
		_w11159_
	);
	LUT2 #(
		.INIT('h4)
	) name10628 (
		_w9980_,
		_w10508_,
		_w11160_
	);
	LUT2 #(
		.INIT('h1)
	) name10629 (
		_w11159_,
		_w11160_,
		_w11161_
	);
	LUT2 #(
		.INIT('h8)
	) name10630 (
		_w11158_,
		_w11161_,
		_w11162_
	);
	LUT2 #(
		.INIT('h1)
	) name10631 (
		_w11158_,
		_w11161_,
		_w11163_
	);
	LUT2 #(
		.INIT('h1)
	) name10632 (
		_w11162_,
		_w11163_,
		_w11164_
	);
	LUT2 #(
		.INIT('h1)
	) name10633 (
		_w11079_,
		_w11164_,
		_w11165_
	);
	LUT2 #(
		.INIT('h8)
	) name10634 (
		_w11079_,
		_w11164_,
		_w11166_
	);
	LUT2 #(
		.INIT('h1)
	) name10635 (
		\ld_r_reg/P0001 ,
		_w11165_,
		_w11167_
	);
	LUT2 #(
		.INIT('h4)
	) name10636 (
		_w11166_,
		_w11167_,
		_w11168_
	);
	LUT2 #(
		.INIT('h1)
	) name10637 (
		\text_in_r_reg[81]/P0001 ,
		\u0_w_reg[1][17]/P0001 ,
		_w11169_
	);
	LUT2 #(
		.INIT('h8)
	) name10638 (
		\text_in_r_reg[81]/P0001 ,
		\u0_w_reg[1][17]/P0001 ,
		_w11170_
	);
	LUT2 #(
		.INIT('h2)
	) name10639 (
		\ld_r_reg/P0001 ,
		_w11169_,
		_w11171_
	);
	LUT2 #(
		.INIT('h4)
	) name10640 (
		_w11170_,
		_w11171_,
		_w11172_
	);
	LUT2 #(
		.INIT('h1)
	) name10641 (
		_w11168_,
		_w11172_,
		_w11173_
	);
	LUT2 #(
		.INIT('h8)
	) name10642 (
		_w10031_,
		_w10920_,
		_w11174_
	);
	LUT2 #(
		.INIT('h2)
	) name10643 (
		\sa12_reg[1]/P0001 ,
		_w9837_,
		_w11175_
	);
	LUT2 #(
		.INIT('h4)
	) name10644 (
		_w10985_,
		_w11175_,
		_w11176_
	);
	LUT2 #(
		.INIT('h4)
	) name10645 (
		_w11174_,
		_w11176_,
		_w11177_
	);
	LUT2 #(
		.INIT('h8)
	) name10646 (
		_w8059_,
		_w8060_,
		_w11178_
	);
	LUT2 #(
		.INIT('h8)
	) name10647 (
		_w8162_,
		_w9817_,
		_w11179_
	);
	LUT2 #(
		.INIT('h1)
	) name10648 (
		\sa12_reg[1]/P0001 ,
		_w8145_,
		_w11180_
	);
	LUT2 #(
		.INIT('h1)
	) name10649 (
		_w10936_,
		_w11178_,
		_w11181_
	);
	LUT2 #(
		.INIT('h8)
	) name10650 (
		_w11180_,
		_w11181_,
		_w11182_
	);
	LUT2 #(
		.INIT('h1)
	) name10651 (
		_w8087_,
		_w8160_,
		_w11183_
	);
	LUT2 #(
		.INIT('h1)
	) name10652 (
		_w8189_,
		_w8453_,
		_w11184_
	);
	LUT2 #(
		.INIT('h4)
	) name10653 (
		_w11179_,
		_w11184_,
		_w11185_
	);
	LUT2 #(
		.INIT('h8)
	) name10654 (
		_w11182_,
		_w11183_,
		_w11186_
	);
	LUT2 #(
		.INIT('h8)
	) name10655 (
		_w11185_,
		_w11186_,
		_w11187_
	);
	LUT2 #(
		.INIT('h1)
	) name10656 (
		_w11177_,
		_w11187_,
		_w11188_
	);
	LUT2 #(
		.INIT('h1)
	) name10657 (
		_w8130_,
		_w9049_,
		_w11189_
	);
	LUT2 #(
		.INIT('h4)
	) name10658 (
		_w8490_,
		_w11189_,
		_w11190_
	);
	LUT2 #(
		.INIT('h2)
	) name10659 (
		_w8057_,
		_w11190_,
		_w11191_
	);
	LUT2 #(
		.INIT('h1)
	) name10660 (
		_w8086_,
		_w8105_,
		_w11192_
	);
	LUT2 #(
		.INIT('h4)
	) name10661 (
		_w10974_,
		_w11192_,
		_w11193_
	);
	LUT2 #(
		.INIT('h4)
	) name10662 (
		_w11191_,
		_w11193_,
		_w11194_
	);
	LUT2 #(
		.INIT('h4)
	) name10663 (
		_w11188_,
		_w11194_,
		_w11195_
	);
	LUT2 #(
		.INIT('h2)
	) name10664 (
		\sa12_reg[0]/P0001 ,
		_w11195_,
		_w11196_
	);
	LUT2 #(
		.INIT('h2)
	) name10665 (
		_w8082_,
		_w8094_,
		_w11197_
	);
	LUT2 #(
		.INIT('h4)
	) name10666 (
		_w8498_,
		_w11197_,
		_w11198_
	);
	LUT2 #(
		.INIT('h1)
	) name10667 (
		_w9047_,
		_w9790_,
		_w11199_
	);
	LUT2 #(
		.INIT('h4)
	) name10668 (
		_w8103_,
		_w11199_,
		_w11200_
	);
	LUT2 #(
		.INIT('h8)
	) name10669 (
		_w8997_,
		_w11200_,
		_w11201_
	);
	LUT2 #(
		.INIT('h2)
	) name10670 (
		\sa12_reg[2]/P0001 ,
		_w8497_,
		_w11202_
	);
	LUT2 #(
		.INIT('h4)
	) name10671 (
		_w9865_,
		_w11202_,
		_w11203_
	);
	LUT2 #(
		.INIT('h4)
	) name10672 (
		_w8098_,
		_w11203_,
		_w11204_
	);
	LUT2 #(
		.INIT('h1)
	) name10673 (
		_w11201_,
		_w11204_,
		_w11205_
	);
	LUT2 #(
		.INIT('h1)
	) name10674 (
		\sa12_reg[1]/P0001 ,
		_w11198_,
		_w11206_
	);
	LUT2 #(
		.INIT('h4)
	) name10675 (
		_w11205_,
		_w11206_,
		_w11207_
	);
	LUT2 #(
		.INIT('h1)
	) name10676 (
		_w8084_,
		_w9042_,
		_w11208_
	);
	LUT2 #(
		.INIT('h1)
	) name10677 (
		\sa12_reg[4]/P0001 ,
		_w11208_,
		_w11209_
	);
	LUT2 #(
		.INIT('h2)
	) name10678 (
		\sa12_reg[2]/P0001 ,
		_w8452_,
		_w11210_
	);
	LUT2 #(
		.INIT('h4)
	) name10679 (
		_w11209_,
		_w11210_,
		_w11211_
	);
	LUT2 #(
		.INIT('h1)
	) name10680 (
		\sa12_reg[2]/P0001 ,
		_w8405_,
		_w11212_
	);
	LUT2 #(
		.INIT('h8)
	) name10681 (
		_w9997_,
		_w11212_,
		_w11213_
	);
	LUT2 #(
		.INIT('h1)
	) name10682 (
		_w11211_,
		_w11213_,
		_w11214_
	);
	LUT2 #(
		.INIT('h2)
	) name10683 (
		\sa12_reg[1]/P0001 ,
		_w8096_,
		_w11215_
	);
	LUT2 #(
		.INIT('h4)
	) name10684 (
		_w11214_,
		_w11215_,
		_w11216_
	);
	LUT2 #(
		.INIT('h1)
	) name10685 (
		_w11207_,
		_w11216_,
		_w11217_
	);
	LUT2 #(
		.INIT('h1)
	) name10686 (
		_w8056_,
		_w8135_,
		_w11218_
	);
	LUT2 #(
		.INIT('h2)
	) name10687 (
		_w8447_,
		_w11218_,
		_w11219_
	);
	LUT2 #(
		.INIT('h1)
	) name10688 (
		_w8138_,
		_w9817_,
		_w11220_
	);
	LUT2 #(
		.INIT('h2)
	) name10689 (
		\sa12_reg[2]/P0001 ,
		_w11220_,
		_w11221_
	);
	LUT2 #(
		.INIT('h1)
	) name10690 (
		_w9035_,
		_w11221_,
		_w11222_
	);
	LUT2 #(
		.INIT('h2)
	) name10691 (
		\sa12_reg[1]/P0001 ,
		_w11222_,
		_w11223_
	);
	LUT2 #(
		.INIT('h1)
	) name10692 (
		_w9865_,
		_w10984_,
		_w11224_
	);
	LUT2 #(
		.INIT('h1)
	) name10693 (
		\sa12_reg[1]/P0001 ,
		_w11224_,
		_w11225_
	);
	LUT2 #(
		.INIT('h1)
	) name10694 (
		_w8185_,
		_w10660_,
		_w11226_
	);
	LUT2 #(
		.INIT('h2)
	) name10695 (
		\sa12_reg[4]/P0001 ,
		_w11226_,
		_w11227_
	);
	LUT2 #(
		.INIT('h1)
	) name10696 (
		_w8075_,
		_w8498_,
		_w11228_
	);
	LUT2 #(
		.INIT('h2)
	) name10697 (
		\sa12_reg[1]/P0001 ,
		_w8074_,
		_w11229_
	);
	LUT2 #(
		.INIT('h4)
	) name10698 (
		_w11228_,
		_w11229_,
		_w11230_
	);
	LUT2 #(
		.INIT('h1)
	) name10699 (
		_w8150_,
		_w11230_,
		_w11231_
	);
	LUT2 #(
		.INIT('h1)
	) name10700 (
		\sa12_reg[2]/P0001 ,
		_w11231_,
		_w11232_
	);
	LUT2 #(
		.INIT('h1)
	) name10701 (
		_w11225_,
		_w11227_,
		_w11233_
	);
	LUT2 #(
		.INIT('h4)
	) name10702 (
		_w11232_,
		_w11233_,
		_w11234_
	);
	LUT2 #(
		.INIT('h4)
	) name10703 (
		_w11223_,
		_w11234_,
		_w11235_
	);
	LUT2 #(
		.INIT('h1)
	) name10704 (
		\sa12_reg[0]/P0001 ,
		_w11235_,
		_w11236_
	);
	LUT2 #(
		.INIT('h1)
	) name10705 (
		_w10672_,
		_w11219_,
		_w11237_
	);
	LUT2 #(
		.INIT('h4)
	) name10706 (
		_w11217_,
		_w11237_,
		_w11238_
	);
	LUT2 #(
		.INIT('h4)
	) name10707 (
		_w11196_,
		_w11238_,
		_w11239_
	);
	LUT2 #(
		.INIT('h4)
	) name10708 (
		_w11236_,
		_w11239_,
		_w11240_
	);
	LUT2 #(
		.INIT('h8)
	) name10709 (
		\sa01_reg[2]/P0001 ,
		_w8276_,
		_w11241_
	);
	LUT2 #(
		.INIT('h4)
	) name10710 (
		_w8318_,
		_w11241_,
		_w11242_
	);
	LUT2 #(
		.INIT('h1)
	) name10711 (
		\sa01_reg[5]/P0001 ,
		_w8246_,
		_w11243_
	);
	LUT2 #(
		.INIT('h2)
	) name10712 (
		_w8339_,
		_w11243_,
		_w11244_
	);
	LUT2 #(
		.INIT('h1)
	) name10713 (
		_w8223_,
		_w10185_,
		_w11245_
	);
	LUT2 #(
		.INIT('h8)
	) name10714 (
		_w8237_,
		_w11245_,
		_w11246_
	);
	LUT2 #(
		.INIT('h1)
	) name10715 (
		_w8312_,
		_w11242_,
		_w11247_
	);
	LUT2 #(
		.INIT('h4)
	) name10716 (
		_w11244_,
		_w11247_,
		_w11248_
	);
	LUT2 #(
		.INIT('h8)
	) name10717 (
		_w11246_,
		_w11248_,
		_w11249_
	);
	LUT2 #(
		.INIT('h1)
	) name10718 (
		_w8242_,
		_w8264_,
		_w11250_
	);
	LUT2 #(
		.INIT('h8)
	) name10719 (
		_w9209_,
		_w11250_,
		_w11251_
	);
	LUT2 #(
		.INIT('h2)
	) name10720 (
		\sa01_reg[1]/P0001 ,
		_w9208_,
		_w11252_
	);
	LUT2 #(
		.INIT('h4)
	) name10721 (
		_w11251_,
		_w11252_,
		_w11253_
	);
	LUT2 #(
		.INIT('h4)
	) name10722 (
		_w10229_,
		_w11253_,
		_w11254_
	);
	LUT2 #(
		.INIT('h1)
	) name10723 (
		_w11249_,
		_w11254_,
		_w11255_
	);
	LUT2 #(
		.INIT('h1)
	) name10724 (
		_w8278_,
		_w8309_,
		_w11256_
	);
	LUT2 #(
		.INIT('h4)
	) name10725 (
		_w8283_,
		_w11256_,
		_w11257_
	);
	LUT2 #(
		.INIT('h1)
	) name10726 (
		\sa01_reg[3]/P0001 ,
		_w11257_,
		_w11258_
	);
	LUT2 #(
		.INIT('h1)
	) name10727 (
		_w8258_,
		_w9276_,
		_w11259_
	);
	LUT2 #(
		.INIT('h4)
	) name10728 (
		_w9368_,
		_w11259_,
		_w11260_
	);
	LUT2 #(
		.INIT('h2)
	) name10729 (
		_w8329_,
		_w11260_,
		_w11261_
	);
	LUT2 #(
		.INIT('h1)
	) name10730 (
		_w11258_,
		_w11261_,
		_w11262_
	);
	LUT2 #(
		.INIT('h4)
	) name10731 (
		_w11255_,
		_w11262_,
		_w11263_
	);
	LUT2 #(
		.INIT('h2)
	) name10732 (
		\sa01_reg[0]/P0001 ,
		_w11263_,
		_w11264_
	);
	LUT2 #(
		.INIT('h4)
	) name10733 (
		_w9196_,
		_w10084_,
		_w11265_
	);
	LUT2 #(
		.INIT('h1)
	) name10734 (
		\sa01_reg[2]/P0001 ,
		_w11265_,
		_w11266_
	);
	LUT2 #(
		.INIT('h1)
	) name10735 (
		_w8352_,
		_w11266_,
		_w11267_
	);
	LUT2 #(
		.INIT('h2)
	) name10736 (
		\sa01_reg[1]/P0001 ,
		_w11267_,
		_w11268_
	);
	LUT2 #(
		.INIT('h1)
	) name10737 (
		_w8320_,
		_w9268_,
		_w11269_
	);
	LUT2 #(
		.INIT('h2)
	) name10738 (
		_w9388_,
		_w11269_,
		_w11270_
	);
	LUT2 #(
		.INIT('h8)
	) name10739 (
		\sa01_reg[1]/P0001 ,
		_w8329_,
		_w11271_
	);
	LUT2 #(
		.INIT('h8)
	) name10740 (
		_w8369_,
		_w11271_,
		_w11272_
	);
	LUT2 #(
		.INIT('h1)
	) name10741 (
		_w8219_,
		_w8254_,
		_w11273_
	);
	LUT2 #(
		.INIT('h2)
	) name10742 (
		_w10230_,
		_w11273_,
		_w11274_
	);
	LUT2 #(
		.INIT('h1)
	) name10743 (
		_w8227_,
		_w9373_,
		_w11275_
	);
	LUT2 #(
		.INIT('h2)
	) name10744 (
		\sa01_reg[3]/P0001 ,
		_w11275_,
		_w11276_
	);
	LUT2 #(
		.INIT('h1)
	) name10745 (
		_w9774_,
		_w11276_,
		_w11277_
	);
	LUT2 #(
		.INIT('h2)
	) name10746 (
		\sa01_reg[2]/P0001 ,
		_w11277_,
		_w11278_
	);
	LUT2 #(
		.INIT('h4)
	) name10747 (
		_w8214_,
		_w8227_,
		_w11279_
	);
	LUT2 #(
		.INIT('h4)
	) name10748 (
		_w8265_,
		_w11279_,
		_w11280_
	);
	LUT2 #(
		.INIT('h1)
	) name10749 (
		_w8309_,
		_w9375_,
		_w11281_
	);
	LUT2 #(
		.INIT('h4)
	) name10750 (
		_w8361_,
		_w11281_,
		_w11282_
	);
	LUT2 #(
		.INIT('h1)
	) name10751 (
		\sa01_reg[2]/P0001 ,
		_w11282_,
		_w11283_
	);
	LUT2 #(
		.INIT('h1)
	) name10752 (
		_w9305_,
		_w11280_,
		_w11284_
	);
	LUT2 #(
		.INIT('h4)
	) name10753 (
		_w11283_,
		_w11284_,
		_w11285_
	);
	LUT2 #(
		.INIT('h4)
	) name10754 (
		_w11278_,
		_w11285_,
		_w11286_
	);
	LUT2 #(
		.INIT('h1)
	) name10755 (
		\sa01_reg[1]/P0001 ,
		_w11286_,
		_w11287_
	);
	LUT2 #(
		.INIT('h1)
	) name10756 (
		_w8266_,
		_w8339_,
		_w11288_
	);
	LUT2 #(
		.INIT('h2)
	) name10757 (
		\sa01_reg[2]/P0001 ,
		_w11288_,
		_w11289_
	);
	LUT2 #(
		.INIT('h1)
	) name10758 (
		_w8264_,
		_w8265_,
		_w11290_
	);
	LUT2 #(
		.INIT('h1)
	) name10759 (
		\sa01_reg[2]/P0001 ,
		_w8342_,
		_w11291_
	);
	LUT2 #(
		.INIT('h4)
	) name10760 (
		_w11290_,
		_w11291_,
		_w11292_
	);
	LUT2 #(
		.INIT('h1)
	) name10761 (
		_w9369_,
		_w11292_,
		_w11293_
	);
	LUT2 #(
		.INIT('h4)
	) name10762 (
		_w11289_,
		_w11293_,
		_w11294_
	);
	LUT2 #(
		.INIT('h2)
	) name10763 (
		\sa01_reg[1]/P0001 ,
		_w11294_,
		_w11295_
	);
	LUT2 #(
		.INIT('h8)
	) name10764 (
		\sa01_reg[2]/P0001 ,
		_w8332_,
		_w11296_
	);
	LUT2 #(
		.INIT('h8)
	) name10765 (
		_w8342_,
		_w9386_,
		_w11297_
	);
	LUT2 #(
		.INIT('h1)
	) name10766 (
		_w9774_,
		_w11297_,
		_w11298_
	);
	LUT2 #(
		.INIT('h1)
	) name10767 (
		\sa01_reg[1]/P0001 ,
		_w11298_,
		_w11299_
	);
	LUT2 #(
		.INIT('h4)
	) name10768 (
		\sa01_reg[2]/P0001 ,
		_w8220_,
		_w11300_
	);
	LUT2 #(
		.INIT('h1)
	) name10769 (
		_w8243_,
		_w11296_,
		_w11301_
	);
	LUT2 #(
		.INIT('h1)
	) name10770 (
		_w11299_,
		_w11300_,
		_w11302_
	);
	LUT2 #(
		.INIT('h8)
	) name10771 (
		_w11301_,
		_w11302_,
		_w11303_
	);
	LUT2 #(
		.INIT('h4)
	) name10772 (
		_w11295_,
		_w11303_,
		_w11304_
	);
	LUT2 #(
		.INIT('h1)
	) name10773 (
		\sa01_reg[0]/P0001 ,
		_w11304_,
		_w11305_
	);
	LUT2 #(
		.INIT('h1)
	) name10774 (
		_w10581_,
		_w11272_,
		_w11306_
	);
	LUT2 #(
		.INIT('h4)
	) name10775 (
		_w11274_,
		_w11306_,
		_w11307_
	);
	LUT2 #(
		.INIT('h4)
	) name10776 (
		_w11270_,
		_w11307_,
		_w11308_
	);
	LUT2 #(
		.INIT('h4)
	) name10777 (
		_w11268_,
		_w11308_,
		_w11309_
	);
	LUT2 #(
		.INIT('h1)
	) name10778 (
		_w11287_,
		_w11305_,
		_w11310_
	);
	LUT2 #(
		.INIT('h8)
	) name10779 (
		_w11309_,
		_w11310_,
		_w11311_
	);
	LUT2 #(
		.INIT('h4)
	) name10780 (
		_w11264_,
		_w11311_,
		_w11312_
	);
	LUT2 #(
		.INIT('h2)
	) name10781 (
		_w11240_,
		_w11312_,
		_w11313_
	);
	LUT2 #(
		.INIT('h4)
	) name10782 (
		_w11240_,
		_w11312_,
		_w11314_
	);
	LUT2 #(
		.INIT('h1)
	) name10783 (
		_w11313_,
		_w11314_,
		_w11315_
	);
	LUT2 #(
		.INIT('h1)
	) name10784 (
		_w10167_,
		_w11315_,
		_w11316_
	);
	LUT2 #(
		.INIT('h8)
	) name10785 (
		_w10167_,
		_w11315_,
		_w11317_
	);
	LUT2 #(
		.INIT('h1)
	) name10786 (
		_w11316_,
		_w11317_,
		_w11318_
	);
	LUT2 #(
		.INIT('h4)
	) name10787 (
		_w8602_,
		_w10477_,
		_w11319_
	);
	LUT2 #(
		.INIT('h1)
	) name10788 (
		_w9497_,
		_w11319_,
		_w11320_
	);
	LUT2 #(
		.INIT('h1)
	) name10789 (
		_w9419_,
		_w9430_,
		_w11321_
	);
	LUT2 #(
		.INIT('h1)
	) name10790 (
		_w9451_,
		_w9943_,
		_w11322_
	);
	LUT2 #(
		.INIT('h8)
	) name10791 (
		_w11321_,
		_w11322_,
		_w11323_
	);
	LUT2 #(
		.INIT('h4)
	) name10792 (
		_w9064_,
		_w11323_,
		_w11324_
	);
	LUT2 #(
		.INIT('h4)
	) name10793 (
		_w11320_,
		_w11324_,
		_w11325_
	);
	LUT2 #(
		.INIT('h1)
	) name10794 (
		\sa23_reg[1]/P0001 ,
		_w11325_,
		_w11326_
	);
	LUT2 #(
		.INIT('h1)
	) name10795 (
		_w8653_,
		_w8667_,
		_w11327_
	);
	LUT2 #(
		.INIT('h4)
	) name10796 (
		_w9152_,
		_w11327_,
		_w11328_
	);
	LUT2 #(
		.INIT('h2)
	) name10797 (
		\sa23_reg[3]/P0001 ,
		_w11328_,
		_w11329_
	);
	LUT2 #(
		.INIT('h1)
	) name10798 (
		_w9492_,
		_w11329_,
		_w11330_
	);
	LUT2 #(
		.INIT('h2)
	) name10799 (
		\sa23_reg[2]/P0001 ,
		_w11330_,
		_w11331_
	);
	LUT2 #(
		.INIT('h2)
	) name10800 (
		\sa23_reg[2]/P0001 ,
		_w8578_,
		_w11332_
	);
	LUT2 #(
		.INIT('h1)
	) name10801 (
		\sa23_reg[2]/P0001 ,
		_w8574_,
		_w11333_
	);
	LUT2 #(
		.INIT('h4)
	) name10802 (
		_w9099_,
		_w11333_,
		_w11334_
	);
	LUT2 #(
		.INIT('h4)
	) name10803 (
		_w8647_,
		_w11334_,
		_w11335_
	);
	LUT2 #(
		.INIT('h2)
	) name10804 (
		\sa23_reg[1]/P0001 ,
		_w11332_,
		_w11336_
	);
	LUT2 #(
		.INIT('h4)
	) name10805 (
		_w11335_,
		_w11336_,
		_w11337_
	);
	LUT2 #(
		.INIT('h1)
	) name10806 (
		_w9464_,
		_w9469_,
		_w11338_
	);
	LUT2 #(
		.INIT('h4)
	) name10807 (
		_w11337_,
		_w11338_,
		_w11339_
	);
	LUT2 #(
		.INIT('h4)
	) name10808 (
		_w11326_,
		_w11339_,
		_w11340_
	);
	LUT2 #(
		.INIT('h4)
	) name10809 (
		_w11331_,
		_w11340_,
		_w11341_
	);
	LUT2 #(
		.INIT('h2)
	) name10810 (
		\sa23_reg[0]/P0001 ,
		_w11341_,
		_w11342_
	);
	LUT2 #(
		.INIT('h1)
	) name10811 (
		_w9159_,
		_w9482_,
		_w11343_
	);
	LUT2 #(
		.INIT('h4)
	) name10812 (
		_w9064_,
		_w11343_,
		_w11344_
	);
	LUT2 #(
		.INIT('h8)
	) name10813 (
		_w9474_,
		_w11344_,
		_w11345_
	);
	LUT2 #(
		.INIT('h8)
	) name10814 (
		\sa23_reg[3]/P0001 ,
		_w8547_,
		_w11346_
	);
	LUT2 #(
		.INIT('h1)
	) name10815 (
		_w9476_,
		_w11346_,
		_w11347_
	);
	LUT2 #(
		.INIT('h8)
	) name10816 (
		_w9953_,
		_w11347_,
		_w11348_
	);
	LUT2 #(
		.INIT('h1)
	) name10817 (
		_w11345_,
		_w11348_,
		_w11349_
	);
	LUT2 #(
		.INIT('h2)
	) name10818 (
		_w8547_,
		_w8573_,
		_w11350_
	);
	LUT2 #(
		.INIT('h4)
	) name10819 (
		_w8577_,
		_w11350_,
		_w11351_
	);
	LUT2 #(
		.INIT('h1)
	) name10820 (
		_w11349_,
		_w11351_,
		_w11352_
	);
	LUT2 #(
		.INIT('h1)
	) name10821 (
		\sa23_reg[1]/P0001 ,
		_w11352_,
		_w11353_
	);
	LUT2 #(
		.INIT('h1)
	) name10822 (
		_w8552_,
		_w8591_,
		_w11354_
	);
	LUT2 #(
		.INIT('h2)
	) name10823 (
		\sa23_reg[2]/P0001 ,
		_w11354_,
		_w11355_
	);
	LUT2 #(
		.INIT('h1)
	) name10824 (
		_w8577_,
		_w8588_,
		_w11356_
	);
	LUT2 #(
		.INIT('h1)
	) name10825 (
		\sa23_reg[2]/P0001 ,
		_w8589_,
		_w11357_
	);
	LUT2 #(
		.INIT('h4)
	) name10826 (
		_w11356_,
		_w11357_,
		_w11358_
	);
	LUT2 #(
		.INIT('h1)
	) name10827 (
		_w9154_,
		_w11358_,
		_w11359_
	);
	LUT2 #(
		.INIT('h4)
	) name10828 (
		_w11355_,
		_w11359_,
		_w11360_
	);
	LUT2 #(
		.INIT('h2)
	) name10829 (
		\sa23_reg[1]/P0001 ,
		_w11360_,
		_w11361_
	);
	LUT2 #(
		.INIT('h4)
	) name10830 (
		_w8620_,
		_w9954_,
		_w11362_
	);
	LUT2 #(
		.INIT('h8)
	) name10831 (
		_w8546_,
		_w8602_,
		_w11363_
	);
	LUT2 #(
		.INIT('h1)
	) name10832 (
		_w8570_,
		_w11363_,
		_w11364_
	);
	LUT2 #(
		.INIT('h4)
	) name10833 (
		_w9135_,
		_w11364_,
		_w11365_
	);
	LUT2 #(
		.INIT('h4)
	) name10834 (
		_w11362_,
		_w11365_,
		_w11366_
	);
	LUT2 #(
		.INIT('h4)
	) name10835 (
		_w11361_,
		_w11366_,
		_w11367_
	);
	LUT2 #(
		.INIT('h1)
	) name10836 (
		\sa23_reg[0]/P0001 ,
		_w11367_,
		_w11368_
	);
	LUT2 #(
		.INIT('h4)
	) name10837 (
		_w8551_,
		_w10443_,
		_w11369_
	);
	LUT2 #(
		.INIT('h1)
	) name10838 (
		\sa23_reg[2]/P0001 ,
		_w11369_,
		_w11370_
	);
	LUT2 #(
		.INIT('h1)
	) name10839 (
		_w8527_,
		_w11370_,
		_w11371_
	);
	LUT2 #(
		.INIT('h2)
	) name10840 (
		\sa23_reg[1]/P0001 ,
		_w11371_,
		_w11372_
	);
	LUT2 #(
		.INIT('h1)
	) name10841 (
		_w8562_,
		_w8631_,
		_w11373_
	);
	LUT2 #(
		.INIT('h2)
	) name10842 (
		_w8522_,
		_w11373_,
		_w11374_
	);
	LUT2 #(
		.INIT('h1)
	) name10843 (
		_w8602_,
		_w8603_,
		_w11375_
	);
	LUT2 #(
		.INIT('h4)
	) name10844 (
		_w9462_,
		_w11375_,
		_w11376_
	);
	LUT2 #(
		.INIT('h2)
	) name10845 (
		\sa23_reg[1]/P0001 ,
		_w11376_,
		_w11377_
	);
	LUT2 #(
		.INIT('h1)
	) name10846 (
		_w11374_,
		_w11377_,
		_w11378_
	);
	LUT2 #(
		.INIT('h2)
	) name10847 (
		\sa23_reg[2]/P0001 ,
		_w11378_,
		_w11379_
	);
	LUT2 #(
		.INIT('h1)
	) name10848 (
		_w10729_,
		_w11379_,
		_w11380_
	);
	LUT2 #(
		.INIT('h4)
	) name10849 (
		_w11353_,
		_w11380_,
		_w11381_
	);
	LUT2 #(
		.INIT('h1)
	) name10850 (
		_w11368_,
		_w11372_,
		_w11382_
	);
	LUT2 #(
		.INIT('h8)
	) name10851 (
		_w11381_,
		_w11382_,
		_w11383_
	);
	LUT2 #(
		.INIT('h4)
	) name10852 (
		_w11342_,
		_w11383_,
		_w11384_
	);
	LUT2 #(
		.INIT('h2)
	) name10853 (
		\u0_w_reg[1][2]/P0001 ,
		_w11384_,
		_w11385_
	);
	LUT2 #(
		.INIT('h4)
	) name10854 (
		\u0_w_reg[1][2]/P0001 ,
		_w11384_,
		_w11386_
	);
	LUT2 #(
		.INIT('h1)
	) name10855 (
		_w11385_,
		_w11386_,
		_w11387_
	);
	LUT2 #(
		.INIT('h8)
	) name10856 (
		_w11155_,
		_w11387_,
		_w11388_
	);
	LUT2 #(
		.INIT('h1)
	) name10857 (
		_w11155_,
		_w11387_,
		_w11389_
	);
	LUT2 #(
		.INIT('h1)
	) name10858 (
		_w11388_,
		_w11389_,
		_w11390_
	);
	LUT2 #(
		.INIT('h4)
	) name10859 (
		_w11318_,
		_w11390_,
		_w11391_
	);
	LUT2 #(
		.INIT('h2)
	) name10860 (
		_w11318_,
		_w11390_,
		_w11392_
	);
	LUT2 #(
		.INIT('h1)
	) name10861 (
		\ld_r_reg/P0001 ,
		_w11391_,
		_w11393_
	);
	LUT2 #(
		.INIT('h4)
	) name10862 (
		_w11392_,
		_w11393_,
		_w11394_
	);
	LUT2 #(
		.INIT('h1)
	) name10863 (
		\text_in_r_reg[66]/P0001 ,
		\u0_w_reg[1][2]/P0001 ,
		_w11395_
	);
	LUT2 #(
		.INIT('h8)
	) name10864 (
		\text_in_r_reg[66]/P0001 ,
		\u0_w_reg[1][2]/P0001 ,
		_w11396_
	);
	LUT2 #(
		.INIT('h2)
	) name10865 (
		\ld_r_reg/P0001 ,
		_w11395_,
		_w11397_
	);
	LUT2 #(
		.INIT('h4)
	) name10866 (
		_w11396_,
		_w11397_,
		_w11398_
	);
	LUT2 #(
		.INIT('h1)
	) name10867 (
		_w11394_,
		_w11398_,
		_w11399_
	);
	LUT2 #(
		.INIT('h2)
	) name10868 (
		_w10081_,
		_w10508_,
		_w11400_
	);
	LUT2 #(
		.INIT('h4)
	) name10869 (
		_w10081_,
		_w10508_,
		_w11401_
	);
	LUT2 #(
		.INIT('h1)
	) name10870 (
		_w11400_,
		_w11401_,
		_w11402_
	);
	LUT2 #(
		.INIT('h2)
	) name10871 (
		\u0_w_reg[1][25]/P0001 ,
		_w11155_,
		_w11403_
	);
	LUT2 #(
		.INIT('h4)
	) name10872 (
		\u0_w_reg[1][25]/P0001 ,
		_w11155_,
		_w11404_
	);
	LUT2 #(
		.INIT('h1)
	) name10873 (
		_w11403_,
		_w11404_,
		_w11405_
	);
	LUT2 #(
		.INIT('h8)
	) name10874 (
		_w11402_,
		_w11405_,
		_w11406_
	);
	LUT2 #(
		.INIT('h1)
	) name10875 (
		_w11402_,
		_w11405_,
		_w11407_
	);
	LUT2 #(
		.INIT('h1)
	) name10876 (
		_w11406_,
		_w11407_,
		_w11408_
	);
	LUT2 #(
		.INIT('h8)
	) name10877 (
		_w10251_,
		_w10999_,
		_w11409_
	);
	LUT2 #(
		.INIT('h1)
	) name10878 (
		_w10251_,
		_w10999_,
		_w11410_
	);
	LUT2 #(
		.INIT('h1)
	) name10879 (
		_w11409_,
		_w11410_,
		_w11411_
	);
	LUT2 #(
		.INIT('h1)
	) name10880 (
		_w11408_,
		_w11411_,
		_w11412_
	);
	LUT2 #(
		.INIT('h8)
	) name10881 (
		_w11408_,
		_w11411_,
		_w11413_
	);
	LUT2 #(
		.INIT('h1)
	) name10882 (
		\ld_r_reg/P0001 ,
		_w11412_,
		_w11414_
	);
	LUT2 #(
		.INIT('h4)
	) name10883 (
		_w11413_,
		_w11414_,
		_w11415_
	);
	LUT2 #(
		.INIT('h1)
	) name10884 (
		\text_in_r_reg[89]/P0001 ,
		\u0_w_reg[1][25]/P0001 ,
		_w11416_
	);
	LUT2 #(
		.INIT('h8)
	) name10885 (
		\text_in_r_reg[89]/P0001 ,
		\u0_w_reg[1][25]/P0001 ,
		_w11417_
	);
	LUT2 #(
		.INIT('h2)
	) name10886 (
		\ld_r_reg/P0001 ,
		_w11416_,
		_w11418_
	);
	LUT2 #(
		.INIT('h4)
	) name10887 (
		_w11417_,
		_w11418_,
		_w11419_
	);
	LUT2 #(
		.INIT('h1)
	) name10888 (
		_w11415_,
		_w11419_,
		_w11420_
	);
	LUT2 #(
		.INIT('h1)
	) name10889 (
		_w9169_,
		_w9877_,
		_w11421_
	);
	LUT2 #(
		.INIT('h8)
	) name10890 (
		_w9169_,
		_w9877_,
		_w11422_
	);
	LUT2 #(
		.INIT('h1)
	) name10891 (
		_w11421_,
		_w11422_,
		_w11423_
	);
	LUT2 #(
		.INIT('h2)
	) name10892 (
		\u0_w_reg[1][15]/P0001 ,
		_w10430_,
		_w11424_
	);
	LUT2 #(
		.INIT('h4)
	) name10893 (
		\u0_w_reg[1][15]/P0001 ,
		_w10430_,
		_w11425_
	);
	LUT2 #(
		.INIT('h1)
	) name10894 (
		_w11424_,
		_w11425_,
		_w11426_
	);
	LUT2 #(
		.INIT('h8)
	) name10895 (
		_w8974_,
		_w11426_,
		_w11427_
	);
	LUT2 #(
		.INIT('h1)
	) name10896 (
		_w8974_,
		_w11426_,
		_w11428_
	);
	LUT2 #(
		.INIT('h1)
	) name10897 (
		_w11427_,
		_w11428_,
		_w11429_
	);
	LUT2 #(
		.INIT('h4)
	) name10898 (
		_w11423_,
		_w11429_,
		_w11430_
	);
	LUT2 #(
		.INIT('h2)
	) name10899 (
		_w11423_,
		_w11429_,
		_w11431_
	);
	LUT2 #(
		.INIT('h1)
	) name10900 (
		\ld_r_reg/P0001 ,
		_w11430_,
		_w11432_
	);
	LUT2 #(
		.INIT('h4)
	) name10901 (
		_w11431_,
		_w11432_,
		_w11433_
	);
	LUT2 #(
		.INIT('h2)
	) name10902 (
		\text_in_r_reg[79]/P0001 ,
		\u0_w_reg[1][15]/P0001 ,
		_w11434_
	);
	LUT2 #(
		.INIT('h4)
	) name10903 (
		\text_in_r_reg[79]/P0001 ,
		\u0_w_reg[1][15]/P0001 ,
		_w11435_
	);
	LUT2 #(
		.INIT('h2)
	) name10904 (
		\ld_r_reg/P0001 ,
		_w11434_,
		_w11436_
	);
	LUT2 #(
		.INIT('h4)
	) name10905 (
		_w11435_,
		_w11436_,
		_w11437_
	);
	LUT2 #(
		.INIT('h1)
	) name10906 (
		_w11433_,
		_w11437_,
		_w11438_
	);
	LUT2 #(
		.INIT('h1)
	) name10907 (
		\u0_w_reg[1][27]/P0001 ,
		_w10898_,
		_w11439_
	);
	LUT2 #(
		.INIT('h8)
	) name10908 (
		\u0_w_reg[1][27]/P0001 ,
		_w10898_,
		_w11440_
	);
	LUT2 #(
		.INIT('h1)
	) name10909 (
		_w11439_,
		_w11440_,
		_w11441_
	);
	LUT2 #(
		.INIT('h2)
	) name10910 (
		_w10682_,
		_w10775_,
		_w11442_
	);
	LUT2 #(
		.INIT('h4)
	) name10911 (
		_w10682_,
		_w10775_,
		_w11443_
	);
	LUT2 #(
		.INIT('h1)
	) name10912 (
		_w11442_,
		_w11443_,
		_w11444_
	);
	LUT2 #(
		.INIT('h8)
	) name10913 (
		_w11441_,
		_w11444_,
		_w11445_
	);
	LUT2 #(
		.INIT('h1)
	) name10914 (
		_w11441_,
		_w11444_,
		_w11446_
	);
	LUT2 #(
		.INIT('h1)
	) name10915 (
		_w11445_,
		_w11446_,
		_w11447_
	);
	LUT2 #(
		.INIT('h2)
	) name10916 (
		_w9783_,
		_w11312_,
		_w11448_
	);
	LUT2 #(
		.INIT('h4)
	) name10917 (
		_w9783_,
		_w11312_,
		_w11449_
	);
	LUT2 #(
		.INIT('h1)
	) name10918 (
		_w11448_,
		_w11449_,
		_w11450_
	);
	LUT2 #(
		.INIT('h2)
	) name10919 (
		_w9874_,
		_w11240_,
		_w11451_
	);
	LUT2 #(
		.INIT('h4)
	) name10920 (
		_w9874_,
		_w11240_,
		_w11452_
	);
	LUT2 #(
		.INIT('h1)
	) name10921 (
		_w11451_,
		_w11452_,
		_w11453_
	);
	LUT2 #(
		.INIT('h2)
	) name10922 (
		_w11450_,
		_w11453_,
		_w11454_
	);
	LUT2 #(
		.INIT('h4)
	) name10923 (
		_w11450_,
		_w11453_,
		_w11455_
	);
	LUT2 #(
		.INIT('h1)
	) name10924 (
		_w11454_,
		_w11455_,
		_w11456_
	);
	LUT2 #(
		.INIT('h1)
	) name10925 (
		_w11447_,
		_w11456_,
		_w11457_
	);
	LUT2 #(
		.INIT('h8)
	) name10926 (
		_w11447_,
		_w11456_,
		_w11458_
	);
	LUT2 #(
		.INIT('h1)
	) name10927 (
		\ld_r_reg/P0001 ,
		_w11457_,
		_w11459_
	);
	LUT2 #(
		.INIT('h4)
	) name10928 (
		_w11458_,
		_w11459_,
		_w11460_
	);
	LUT2 #(
		.INIT('h2)
	) name10929 (
		\text_in_r_reg[91]/P0001 ,
		\u0_w_reg[1][27]/P0001 ,
		_w11461_
	);
	LUT2 #(
		.INIT('h4)
	) name10930 (
		\text_in_r_reg[91]/P0001 ,
		\u0_w_reg[1][27]/P0001 ,
		_w11462_
	);
	LUT2 #(
		.INIT('h2)
	) name10931 (
		\ld_r_reg/P0001 ,
		_w11461_,
		_w11463_
	);
	LUT2 #(
		.INIT('h4)
	) name10932 (
		_w11462_,
		_w11463_,
		_w11464_
	);
	LUT2 #(
		.INIT('h1)
	) name10933 (
		_w11460_,
		_w11464_,
		_w11465_
	);
	LUT2 #(
		.INIT('h2)
	) name10934 (
		\u0_w_reg[1][19]/P0001 ,
		_w10898_,
		_w11466_
	);
	LUT2 #(
		.INIT('h4)
	) name10935 (
		\u0_w_reg[1][19]/P0001 ,
		_w10898_,
		_w11467_
	);
	LUT2 #(
		.INIT('h1)
	) name10936 (
		_w11466_,
		_w11467_,
		_w11468_
	);
	LUT2 #(
		.INIT('h8)
	) name10937 (
		_w10907_,
		_w11468_,
		_w11469_
	);
	LUT2 #(
		.INIT('h1)
	) name10938 (
		_w10907_,
		_w11468_,
		_w11470_
	);
	LUT2 #(
		.INIT('h1)
	) name10939 (
		_w11469_,
		_w11470_,
		_w11471_
	);
	LUT2 #(
		.INIT('h2)
	) name10940 (
		_w10602_,
		_w11384_,
		_w11472_
	);
	LUT2 #(
		.INIT('h4)
	) name10941 (
		_w10602_,
		_w11384_,
		_w11473_
	);
	LUT2 #(
		.INIT('h1)
	) name10942 (
		_w11472_,
		_w11473_,
		_w11474_
	);
	LUT2 #(
		.INIT('h8)
	) name10943 (
		_w11453_,
		_w11474_,
		_w11475_
	);
	LUT2 #(
		.INIT('h1)
	) name10944 (
		_w11453_,
		_w11474_,
		_w11476_
	);
	LUT2 #(
		.INIT('h1)
	) name10945 (
		_w11475_,
		_w11476_,
		_w11477_
	);
	LUT2 #(
		.INIT('h1)
	) name10946 (
		_w11471_,
		_w11477_,
		_w11478_
	);
	LUT2 #(
		.INIT('h8)
	) name10947 (
		_w11471_,
		_w11477_,
		_w11479_
	);
	LUT2 #(
		.INIT('h1)
	) name10948 (
		\ld_r_reg/P0001 ,
		_w11478_,
		_w11480_
	);
	LUT2 #(
		.INIT('h4)
	) name10949 (
		_w11479_,
		_w11480_,
		_w11481_
	);
	LUT2 #(
		.INIT('h2)
	) name10950 (
		\text_in_r_reg[83]/P0001 ,
		\u0_w_reg[1][19]/P0001 ,
		_w11482_
	);
	LUT2 #(
		.INIT('h4)
	) name10951 (
		\text_in_r_reg[83]/P0001 ,
		\u0_w_reg[1][19]/P0001 ,
		_w11483_
	);
	LUT2 #(
		.INIT('h2)
	) name10952 (
		\ld_r_reg/P0001 ,
		_w11482_,
		_w11484_
	);
	LUT2 #(
		.INIT('h4)
	) name10953 (
		_w11483_,
		_w11484_,
		_w11485_
	);
	LUT2 #(
		.INIT('h1)
	) name10954 (
		_w11481_,
		_w11485_,
		_w11486_
	);
	LUT2 #(
		.INIT('h2)
	) name10955 (
		_w10602_,
		_w10682_,
		_w11487_
	);
	LUT2 #(
		.INIT('h4)
	) name10956 (
		_w10602_,
		_w10682_,
		_w11488_
	);
	LUT2 #(
		.INIT('h1)
	) name10957 (
		_w11487_,
		_w11488_,
		_w11489_
	);
	LUT2 #(
		.INIT('h2)
	) name10958 (
		_w9980_,
		_w11384_,
		_w11490_
	);
	LUT2 #(
		.INIT('h4)
	) name10959 (
		_w9980_,
		_w11384_,
		_w11491_
	);
	LUT2 #(
		.INIT('h1)
	) name10960 (
		_w11490_,
		_w11491_,
		_w11492_
	);
	LUT2 #(
		.INIT('h8)
	) name10961 (
		_w11489_,
		_w11492_,
		_w11493_
	);
	LUT2 #(
		.INIT('h1)
	) name10962 (
		_w11489_,
		_w11492_,
		_w11494_
	);
	LUT2 #(
		.INIT('h1)
	) name10963 (
		_w11493_,
		_w11494_,
		_w11495_
	);
	LUT2 #(
		.INIT('h1)
	) name10964 (
		_w8816_,
		_w8961_,
		_w11496_
	);
	LUT2 #(
		.INIT('h4)
	) name10965 (
		_w10351_,
		_w11496_,
		_w11497_
	);
	LUT2 #(
		.INIT('h2)
	) name10966 (
		_w8844_,
		_w11497_,
		_w11498_
	);
	LUT2 #(
		.INIT('h8)
	) name10967 (
		\sa30_reg[2]/P0001 ,
		_w8733_,
		_w11499_
	);
	LUT2 #(
		.INIT('h4)
	) name10968 (
		_w8758_,
		_w10372_,
		_w11500_
	);
	LUT2 #(
		.INIT('h2)
	) name10969 (
		\sa30_reg[1]/P0001 ,
		_w11499_,
		_w11501_
	);
	LUT2 #(
		.INIT('h4)
	) name10970 (
		_w11500_,
		_w11501_,
		_w11502_
	);
	LUT2 #(
		.INIT('h4)
	) name10971 (
		_w10332_,
		_w11502_,
		_w11503_
	);
	LUT2 #(
		.INIT('h8)
	) name10972 (
		_w8724_,
		_w9582_,
		_w11504_
	);
	LUT2 #(
		.INIT('h1)
	) name10973 (
		_w9576_,
		_w10263_,
		_w11505_
	);
	LUT2 #(
		.INIT('h4)
	) name10974 (
		_w11132_,
		_w11505_,
		_w11506_
	);
	LUT2 #(
		.INIT('h1)
	) name10975 (
		_w8765_,
		_w8894_,
		_w11507_
	);
	LUT2 #(
		.INIT('h1)
	) name10976 (
		_w9546_,
		_w11504_,
		_w11508_
	);
	LUT2 #(
		.INIT('h8)
	) name10977 (
		_w11507_,
		_w11508_,
		_w11509_
	);
	LUT2 #(
		.INIT('h8)
	) name10978 (
		_w9587_,
		_w11506_,
		_w11510_
	);
	LUT2 #(
		.INIT('h8)
	) name10979 (
		_w11509_,
		_w11510_,
		_w11511_
	);
	LUT2 #(
		.INIT('h1)
	) name10980 (
		_w11503_,
		_w11511_,
		_w11512_
	);
	LUT2 #(
		.INIT('h2)
	) name10981 (
		\sa30_reg[0]/P0002 ,
		_w9566_,
		_w11513_
	);
	LUT2 #(
		.INIT('h1)
	) name10982 (
		_w10333_,
		_w11133_,
		_w11514_
	);
	LUT2 #(
		.INIT('h8)
	) name10983 (
		_w11513_,
		_w11514_,
		_w11515_
	);
	LUT2 #(
		.INIT('h4)
	) name10984 (
		_w11498_,
		_w11515_,
		_w11516_
	);
	LUT2 #(
		.INIT('h4)
	) name10985 (
		_w11512_,
		_w11516_,
		_w11517_
	);
	LUT2 #(
		.INIT('h8)
	) name10986 (
		_w8756_,
		_w8940_,
		_w11518_
	);
	LUT2 #(
		.INIT('h1)
	) name10987 (
		\sa30_reg[1]/P0001 ,
		_w8785_,
		_w11519_
	);
	LUT2 #(
		.INIT('h4)
	) name10988 (
		_w11518_,
		_w11519_,
		_w11520_
	);
	LUT2 #(
		.INIT('h2)
	) name10989 (
		\sa30_reg[2]/P0001 ,
		_w8724_,
		_w11521_
	);
	LUT2 #(
		.INIT('h4)
	) name10990 (
		_w8760_,
		_w11521_,
		_w11522_
	);
	LUT2 #(
		.INIT('h4)
	) name10991 (
		_w8756_,
		_w8758_,
		_w11523_
	);
	LUT2 #(
		.INIT('h1)
	) name10992 (
		\sa30_reg[2]/P0001 ,
		_w8748_,
		_w11524_
	);
	LUT2 #(
		.INIT('h4)
	) name10993 (
		_w11523_,
		_w11524_,
		_w11525_
	);
	LUT2 #(
		.INIT('h1)
	) name10994 (
		_w11522_,
		_w11525_,
		_w11526_
	);
	LUT2 #(
		.INIT('h2)
	) name10995 (
		\sa30_reg[1]/P0001 ,
		_w10363_,
		_w11527_
	);
	LUT2 #(
		.INIT('h4)
	) name10996 (
		_w11526_,
		_w11527_,
		_w11528_
	);
	LUT2 #(
		.INIT('h1)
	) name10997 (
		_w11520_,
		_w11528_,
		_w11529_
	);
	LUT2 #(
		.INIT('h8)
	) name10998 (
		_w8811_,
		_w9596_,
		_w11530_
	);
	LUT2 #(
		.INIT('h1)
	) name10999 (
		\sa30_reg[0]/P0002 ,
		_w8899_,
		_w11531_
	);
	LUT2 #(
		.INIT('h4)
	) name11000 (
		_w11530_,
		_w11531_,
		_w11532_
	);
	LUT2 #(
		.INIT('h4)
	) name11001 (
		_w8832_,
		_w11532_,
		_w11533_
	);
	LUT2 #(
		.INIT('h4)
	) name11002 (
		_w11529_,
		_w11533_,
		_w11534_
	);
	LUT2 #(
		.INIT('h1)
	) name11003 (
		_w11517_,
		_w11534_,
		_w11535_
	);
	LUT2 #(
		.INIT('h1)
	) name11004 (
		_w8845_,
		_w8874_,
		_w11536_
	);
	LUT2 #(
		.INIT('h4)
	) name11005 (
		\sa30_reg[3]/P0001 ,
		_w9575_,
		_w11537_
	);
	LUT2 #(
		.INIT('h4)
	) name11006 (
		_w11536_,
		_w11537_,
		_w11538_
	);
	LUT2 #(
		.INIT('h1)
	) name11007 (
		_w8775_,
		_w8952_,
		_w11539_
	);
	LUT2 #(
		.INIT('h2)
	) name11008 (
		\sa30_reg[3]/P0001 ,
		_w11539_,
		_w11540_
	);
	LUT2 #(
		.INIT('h2)
	) name11009 (
		_w10413_,
		_w11540_,
		_w11541_
	);
	LUT2 #(
		.INIT('h1)
	) name11010 (
		\sa30_reg[2]/P0001 ,
		_w8964_,
		_w11542_
	);
	LUT2 #(
		.INIT('h4)
	) name11011 (
		_w8822_,
		_w11542_,
		_w11543_
	);
	LUT2 #(
		.INIT('h1)
	) name11012 (
		_w8894_,
		_w10418_,
		_w11544_
	);
	LUT2 #(
		.INIT('h8)
	) name11013 (
		_w11543_,
		_w11544_,
		_w11545_
	);
	LUT2 #(
		.INIT('h1)
	) name11014 (
		_w11541_,
		_w11545_,
		_w11546_
	);
	LUT2 #(
		.INIT('h8)
	) name11015 (
		_w8695_,
		_w8775_,
		_w11547_
	);
	LUT2 #(
		.INIT('h1)
	) name11016 (
		\sa30_reg[1]/P0001 ,
		_w11547_,
		_w11548_
	);
	LUT2 #(
		.INIT('h4)
	) name11017 (
		_w9543_,
		_w11548_,
		_w11549_
	);
	LUT2 #(
		.INIT('h4)
	) name11018 (
		_w11546_,
		_w11549_,
		_w11550_
	);
	LUT2 #(
		.INIT('h8)
	) name11019 (
		_w8723_,
		_w11080_,
		_w11551_
	);
	LUT2 #(
		.INIT('h8)
	) name11020 (
		_w8792_,
		_w8838_,
		_w11552_
	);
	LUT2 #(
		.INIT('h2)
	) name11021 (
		\sa30_reg[2]/P0001 ,
		_w8719_,
		_w11553_
	);
	LUT2 #(
		.INIT('h4)
	) name11022 (
		_w8823_,
		_w11553_,
		_w11554_
	);
	LUT2 #(
		.INIT('h4)
	) name11023 (
		_w11552_,
		_w11554_,
		_w11555_
	);
	LUT2 #(
		.INIT('h1)
	) name11024 (
		_w11551_,
		_w11555_,
		_w11556_
	);
	LUT2 #(
		.INIT('h2)
	) name11025 (
		\sa30_reg[1]/P0001 ,
		_w8711_,
		_w11557_
	);
	LUT2 #(
		.INIT('h4)
	) name11026 (
		_w11556_,
		_w11557_,
		_w11558_
	);
	LUT2 #(
		.INIT('h1)
	) name11027 (
		_w11550_,
		_w11558_,
		_w11559_
	);
	LUT2 #(
		.INIT('h1)
	) name11028 (
		_w10875_,
		_w11538_,
		_w11560_
	);
	LUT2 #(
		.INIT('h4)
	) name11029 (
		_w11559_,
		_w11560_,
		_w11561_
	);
	LUT2 #(
		.INIT('h4)
	) name11030 (
		_w11535_,
		_w11561_,
		_w11562_
	);
	LUT2 #(
		.INIT('h2)
	) name11031 (
		_w10430_,
		_w11562_,
		_w11563_
	);
	LUT2 #(
		.INIT('h4)
	) name11032 (
		_w10430_,
		_w11562_,
		_w11564_
	);
	LUT2 #(
		.INIT('h1)
	) name11033 (
		_w11563_,
		_w11564_,
		_w11565_
	);
	LUT2 #(
		.INIT('h2)
	) name11034 (
		\u0_w_reg[1][11]/P0001 ,
		_w10898_,
		_w11566_
	);
	LUT2 #(
		.INIT('h4)
	) name11035 (
		\u0_w_reg[1][11]/P0001 ,
		_w10898_,
		_w11567_
	);
	LUT2 #(
		.INIT('h1)
	) name11036 (
		_w11566_,
		_w11567_,
		_w11568_
	);
	LUT2 #(
		.INIT('h8)
	) name11037 (
		_w11565_,
		_w11568_,
		_w11569_
	);
	LUT2 #(
		.INIT('h1)
	) name11038 (
		_w11565_,
		_w11568_,
		_w11570_
	);
	LUT2 #(
		.INIT('h1)
	) name11039 (
		_w11569_,
		_w11570_,
		_w11571_
	);
	LUT2 #(
		.INIT('h1)
	) name11040 (
		_w11495_,
		_w11571_,
		_w11572_
	);
	LUT2 #(
		.INIT('h8)
	) name11041 (
		_w11495_,
		_w11571_,
		_w11573_
	);
	LUT2 #(
		.INIT('h1)
	) name11042 (
		\ld_r_reg/P0001 ,
		_w11572_,
		_w11574_
	);
	LUT2 #(
		.INIT('h4)
	) name11043 (
		_w11573_,
		_w11574_,
		_w11575_
	);
	LUT2 #(
		.INIT('h2)
	) name11044 (
		\text_in_r_reg[75]/P0001 ,
		\u0_w_reg[1][11]/P0001 ,
		_w11576_
	);
	LUT2 #(
		.INIT('h4)
	) name11045 (
		\text_in_r_reg[75]/P0001 ,
		\u0_w_reg[1][11]/P0001 ,
		_w11577_
	);
	LUT2 #(
		.INIT('h2)
	) name11046 (
		\ld_r_reg/P0001 ,
		_w11576_,
		_w11578_
	);
	LUT2 #(
		.INIT('h4)
	) name11047 (
		_w11577_,
		_w11578_,
		_w11579_
	);
	LUT2 #(
		.INIT('h1)
	) name11048 (
		_w11575_,
		_w11579_,
		_w11580_
	);
	LUT2 #(
		.INIT('h1)
	) name11049 (
		_w9516_,
		_w10430_,
		_w11581_
	);
	LUT2 #(
		.INIT('h8)
	) name11050 (
		_w9516_,
		_w10430_,
		_w11582_
	);
	LUT2 #(
		.INIT('h1)
	) name11051 (
		_w11581_,
		_w11582_,
		_w11583_
	);
	LUT2 #(
		.INIT('h2)
	) name11052 (
		\u0_w_reg[1][4]/P0001 ,
		_w10898_,
		_w11584_
	);
	LUT2 #(
		.INIT('h4)
	) name11053 (
		\u0_w_reg[1][4]/P0001 ,
		_w10898_,
		_w11585_
	);
	LUT2 #(
		.INIT('h1)
	) name11054 (
		_w11584_,
		_w11585_,
		_w11586_
	);
	LUT2 #(
		.INIT('h8)
	) name11055 (
		_w11583_,
		_w11586_,
		_w11587_
	);
	LUT2 #(
		.INIT('h1)
	) name11056 (
		_w11583_,
		_w11586_,
		_w11588_
	);
	LUT2 #(
		.INIT('h1)
	) name11057 (
		_w11587_,
		_w11588_,
		_w11589_
	);
	LUT2 #(
		.INIT('h4)
	) name11058 (
		_w8379_,
		_w10605_,
		_w11590_
	);
	LUT2 #(
		.INIT('h2)
	) name11059 (
		_w8379_,
		_w10605_,
		_w11591_
	);
	LUT2 #(
		.INIT('h1)
	) name11060 (
		_w11590_,
		_w11591_,
		_w11592_
	);
	LUT2 #(
		.INIT('h1)
	) name11061 (
		_w11589_,
		_w11592_,
		_w11593_
	);
	LUT2 #(
		.INIT('h8)
	) name11062 (
		_w11589_,
		_w11592_,
		_w11594_
	);
	LUT2 #(
		.INIT('h1)
	) name11063 (
		\ld_r_reg/P0001 ,
		_w11593_,
		_w11595_
	);
	LUT2 #(
		.INIT('h4)
	) name11064 (
		_w11594_,
		_w11595_,
		_w11596_
	);
	LUT2 #(
		.INIT('h2)
	) name11065 (
		\text_in_r_reg[68]/P0001 ,
		\u0_w_reg[1][4]/P0001 ,
		_w11597_
	);
	LUT2 #(
		.INIT('h4)
	) name11066 (
		\text_in_r_reg[68]/P0001 ,
		\u0_w_reg[1][4]/P0001 ,
		_w11598_
	);
	LUT2 #(
		.INIT('h2)
	) name11067 (
		\ld_r_reg/P0001 ,
		_w11597_,
		_w11599_
	);
	LUT2 #(
		.INIT('h4)
	) name11068 (
		_w11598_,
		_w11599_,
		_w11600_
	);
	LUT2 #(
		.INIT('h1)
	) name11069 (
		_w11596_,
		_w11600_,
		_w11601_
	);
	LUT2 #(
		.INIT('h1)
	) name11070 (
		\u0_w_reg[1][26]/P0001 ,
		_w11562_,
		_w11602_
	);
	LUT2 #(
		.INIT('h8)
	) name11071 (
		\u0_w_reg[1][26]/P0001 ,
		_w11562_,
		_w11603_
	);
	LUT2 #(
		.INIT('h1)
	) name11072 (
		_w11602_,
		_w11603_,
		_w11604_
	);
	LUT2 #(
		.INIT('h4)
	) name11073 (
		_w11240_,
		_w11384_,
		_w11605_
	);
	LUT2 #(
		.INIT('h2)
	) name11074 (
		_w11240_,
		_w11384_,
		_w11606_
	);
	LUT2 #(
		.INIT('h1)
	) name11075 (
		_w11605_,
		_w11606_,
		_w11607_
	);
	LUT2 #(
		.INIT('h8)
	) name11076 (
		_w11604_,
		_w11607_,
		_w11608_
	);
	LUT2 #(
		.INIT('h1)
	) name11077 (
		_w11604_,
		_w11607_,
		_w11609_
	);
	LUT2 #(
		.INIT('h1)
	) name11078 (
		_w11608_,
		_w11609_,
		_w11610_
	);
	LUT2 #(
		.INIT('h1)
	) name11079 (
		_w10170_,
		_w11610_,
		_w11611_
	);
	LUT2 #(
		.INIT('h8)
	) name11080 (
		_w10170_,
		_w11610_,
		_w11612_
	);
	LUT2 #(
		.INIT('h1)
	) name11081 (
		\ld_r_reg/P0001 ,
		_w11611_,
		_w11613_
	);
	LUT2 #(
		.INIT('h4)
	) name11082 (
		_w11612_,
		_w11613_,
		_w11614_
	);
	LUT2 #(
		.INIT('h1)
	) name11083 (
		\text_in_r_reg[90]/P0001 ,
		\u0_w_reg[1][26]/P0001 ,
		_w11615_
	);
	LUT2 #(
		.INIT('h8)
	) name11084 (
		\text_in_r_reg[90]/P0001 ,
		\u0_w_reg[1][26]/P0001 ,
		_w11616_
	);
	LUT2 #(
		.INIT('h2)
	) name11085 (
		\ld_r_reg/P0001 ,
		_w11615_,
		_w11617_
	);
	LUT2 #(
		.INIT('h4)
	) name11086 (
		_w11616_,
		_w11617_,
		_w11618_
	);
	LUT2 #(
		.INIT('h1)
	) name11087 (
		_w11614_,
		_w11618_,
		_w11619_
	);
	LUT2 #(
		.INIT('h2)
	) name11088 (
		\u0_w_reg[1][31]/P0001 ,
		_w10430_,
		_w11620_
	);
	LUT2 #(
		.INIT('h4)
	) name11089 (
		\u0_w_reg[1][31]/P0001 ,
		_w10430_,
		_w11621_
	);
	LUT2 #(
		.INIT('h1)
	) name11090 (
		_w11620_,
		_w11621_,
		_w11622_
	);
	LUT2 #(
		.INIT('h4)
	) name11091 (
		_w9874_,
		_w9980_,
		_w11623_
	);
	LUT2 #(
		.INIT('h2)
	) name11092 (
		_w9874_,
		_w9980_,
		_w11624_
	);
	LUT2 #(
		.INIT('h1)
	) name11093 (
		_w11623_,
		_w11624_,
		_w11625_
	);
	LUT2 #(
		.INIT('h8)
	) name11094 (
		_w9657_,
		_w11625_,
		_w11626_
	);
	LUT2 #(
		.INIT('h1)
	) name11095 (
		_w9657_,
		_w11625_,
		_w11627_
	);
	LUT2 #(
		.INIT('h1)
	) name11096 (
		_w11626_,
		_w11627_,
		_w11628_
	);
	LUT2 #(
		.INIT('h4)
	) name11097 (
		_w11622_,
		_w11628_,
		_w11629_
	);
	LUT2 #(
		.INIT('h2)
	) name11098 (
		_w11622_,
		_w11628_,
		_w11630_
	);
	LUT2 #(
		.INIT('h1)
	) name11099 (
		\ld_r_reg/P0001 ,
		_w11629_,
		_w11631_
	);
	LUT2 #(
		.INIT('h4)
	) name11100 (
		_w11630_,
		_w11631_,
		_w11632_
	);
	LUT2 #(
		.INIT('h2)
	) name11101 (
		\text_in_r_reg[95]/P0001 ,
		\u0_w_reg[1][31]/P0001 ,
		_w11633_
	);
	LUT2 #(
		.INIT('h4)
	) name11102 (
		\text_in_r_reg[95]/P0001 ,
		\u0_w_reg[1][31]/P0001 ,
		_w11634_
	);
	LUT2 #(
		.INIT('h2)
	) name11103 (
		\ld_r_reg/P0001 ,
		_w11633_,
		_w11635_
	);
	LUT2 #(
		.INIT('h4)
	) name11104 (
		_w11634_,
		_w11635_,
		_w11636_
	);
	LUT2 #(
		.INIT('h1)
	) name11105 (
		_w11632_,
		_w11636_,
		_w11637_
	);
	LUT2 #(
		.INIT('h1)
	) name11106 (
		\u0_w_reg[1][16]/P0001 ,
		_w10344_,
		_w11638_
	);
	LUT2 #(
		.INIT('h8)
	) name11107 (
		\u0_w_reg[1][16]/P0001 ,
		_w10344_,
		_w11639_
	);
	LUT2 #(
		.INIT('h1)
	) name11108 (
		_w11638_,
		_w11639_,
		_w11640_
	);
	LUT2 #(
		.INIT('h2)
	) name11109 (
		_w9980_,
		_w11073_,
		_w11641_
	);
	LUT2 #(
		.INIT('h4)
	) name11110 (
		_w9980_,
		_w11073_,
		_w11642_
	);
	LUT2 #(
		.INIT('h1)
	) name11111 (
		_w11641_,
		_w11642_,
		_w11643_
	);
	LUT2 #(
		.INIT('h2)
	) name11112 (
		_w9874_,
		_w10248_,
		_w11644_
	);
	LUT2 #(
		.INIT('h4)
	) name11113 (
		_w9874_,
		_w10248_,
		_w11645_
	);
	LUT2 #(
		.INIT('h1)
	) name11114 (
		_w11644_,
		_w11645_,
		_w11646_
	);
	LUT2 #(
		.INIT('h8)
	) name11115 (
		_w11643_,
		_w11646_,
		_w11647_
	);
	LUT2 #(
		.INIT('h1)
	) name11116 (
		_w11643_,
		_w11646_,
		_w11648_
	);
	LUT2 #(
		.INIT('h1)
	) name11117 (
		_w11647_,
		_w11648_,
		_w11649_
	);
	LUT2 #(
		.INIT('h4)
	) name11118 (
		_w11640_,
		_w11649_,
		_w11650_
	);
	LUT2 #(
		.INIT('h2)
	) name11119 (
		_w11640_,
		_w11649_,
		_w11651_
	);
	LUT2 #(
		.INIT('h1)
	) name11120 (
		\ld_r_reg/P0001 ,
		_w11650_,
		_w11652_
	);
	LUT2 #(
		.INIT('h4)
	) name11121 (
		_w11651_,
		_w11652_,
		_w11653_
	);
	LUT2 #(
		.INIT('h1)
	) name11122 (
		\text_in_r_reg[80]/P0001 ,
		\u0_w_reg[1][16]/P0001 ,
		_w11654_
	);
	LUT2 #(
		.INIT('h8)
	) name11123 (
		\text_in_r_reg[80]/P0001 ,
		\u0_w_reg[1][16]/P0001 ,
		_w11655_
	);
	LUT2 #(
		.INIT('h2)
	) name11124 (
		\ld_r_reg/P0001 ,
		_w11654_,
		_w11656_
	);
	LUT2 #(
		.INIT('h4)
	) name11125 (
		_w11655_,
		_w11656_,
		_w11657_
	);
	LUT2 #(
		.INIT('h1)
	) name11126 (
		_w11653_,
		_w11657_,
		_w11658_
	);
	LUT2 #(
		.INIT('h1)
	) name11127 (
		_w11312_,
		_w11402_,
		_w11659_
	);
	LUT2 #(
		.INIT('h8)
	) name11128 (
		_w11312_,
		_w11402_,
		_w11660_
	);
	LUT2 #(
		.INIT('h1)
	) name11129 (
		_w11659_,
		_w11660_,
		_w11661_
	);
	LUT2 #(
		.INIT('h2)
	) name11130 (
		\u0_w_reg[1][18]/P0001 ,
		_w11562_,
		_w11662_
	);
	LUT2 #(
		.INIT('h4)
	) name11131 (
		\u0_w_reg[1][18]/P0001 ,
		_w11562_,
		_w11663_
	);
	LUT2 #(
		.INIT('h1)
	) name11132 (
		_w11662_,
		_w11663_,
		_w11664_
	);
	LUT2 #(
		.INIT('h8)
	) name11133 (
		_w11384_,
		_w11664_,
		_w11665_
	);
	LUT2 #(
		.INIT('h1)
	) name11134 (
		_w11384_,
		_w11664_,
		_w11666_
	);
	LUT2 #(
		.INIT('h1)
	) name11135 (
		_w11665_,
		_w11666_,
		_w11667_
	);
	LUT2 #(
		.INIT('h1)
	) name11136 (
		_w11661_,
		_w11667_,
		_w11668_
	);
	LUT2 #(
		.INIT('h8)
	) name11137 (
		_w11661_,
		_w11667_,
		_w11669_
	);
	LUT2 #(
		.INIT('h1)
	) name11138 (
		\ld_r_reg/P0001 ,
		_w11668_,
		_w11670_
	);
	LUT2 #(
		.INIT('h4)
	) name11139 (
		_w11669_,
		_w11670_,
		_w11671_
	);
	LUT2 #(
		.INIT('h2)
	) name11140 (
		\text_in_r_reg[82]/P0001 ,
		\u0_w_reg[1][18]/P0001 ,
		_w11672_
	);
	LUT2 #(
		.INIT('h4)
	) name11141 (
		\text_in_r_reg[82]/P0001 ,
		\u0_w_reg[1][18]/P0001 ,
		_w11673_
	);
	LUT2 #(
		.INIT('h2)
	) name11142 (
		\ld_r_reg/P0001 ,
		_w11672_,
		_w11674_
	);
	LUT2 #(
		.INIT('h4)
	) name11143 (
		_w11673_,
		_w11674_,
		_w11675_
	);
	LUT2 #(
		.INIT('h1)
	) name11144 (
		_w11671_,
		_w11675_,
		_w11676_
	);
	LUT2 #(
		.INIT('h1)
	) name11145 (
		_w9172_,
		_w9783_,
		_w11677_
	);
	LUT2 #(
		.INIT('h8)
	) name11146 (
		_w9172_,
		_w9783_,
		_w11678_
	);
	LUT2 #(
		.INIT('h1)
	) name11147 (
		_w11677_,
		_w11678_,
		_w11679_
	);
	LUT2 #(
		.INIT('h2)
	) name11148 (
		_w9980_,
		_w10430_,
		_w11680_
	);
	LUT2 #(
		.INIT('h4)
	) name11149 (
		_w9980_,
		_w10430_,
		_w11681_
	);
	LUT2 #(
		.INIT('h1)
	) name11150 (
		_w11680_,
		_w11681_,
		_w11682_
	);
	LUT2 #(
		.INIT('h1)
	) name11151 (
		\u0_w_reg[1][23]/P0001 ,
		_w11682_,
		_w11683_
	);
	LUT2 #(
		.INIT('h8)
	) name11152 (
		\u0_w_reg[1][23]/P0001 ,
		_w11682_,
		_w11684_
	);
	LUT2 #(
		.INIT('h1)
	) name11153 (
		_w11683_,
		_w11684_,
		_w11685_
	);
	LUT2 #(
		.INIT('h1)
	) name11154 (
		_w11679_,
		_w11685_,
		_w11686_
	);
	LUT2 #(
		.INIT('h8)
	) name11155 (
		_w11679_,
		_w11685_,
		_w11687_
	);
	LUT2 #(
		.INIT('h1)
	) name11156 (
		\ld_r_reg/P0001 ,
		_w11686_,
		_w11688_
	);
	LUT2 #(
		.INIT('h4)
	) name11157 (
		_w11687_,
		_w11688_,
		_w11689_
	);
	LUT2 #(
		.INIT('h2)
	) name11158 (
		\text_in_r_reg[87]/P0001 ,
		\u0_w_reg[1][23]/P0001 ,
		_w11690_
	);
	LUT2 #(
		.INIT('h4)
	) name11159 (
		\text_in_r_reg[87]/P0001 ,
		\u0_w_reg[1][23]/P0001 ,
		_w11691_
	);
	LUT2 #(
		.INIT('h2)
	) name11160 (
		\ld_r_reg/P0001 ,
		_w11690_,
		_w11692_
	);
	LUT2 #(
		.INIT('h4)
	) name11161 (
		_w11691_,
		_w11692_,
		_w11693_
	);
	LUT2 #(
		.INIT('h1)
	) name11162 (
		_w11689_,
		_w11693_,
		_w11694_
	);
	LUT2 #(
		.INIT('h1)
	) name11163 (
		\u0_w_reg[1][24]/P0002 ,
		_w10344_,
		_w11695_
	);
	LUT2 #(
		.INIT('h8)
	) name11164 (
		\u0_w_reg[1][24]/P0002 ,
		_w10344_,
		_w11696_
	);
	LUT2 #(
		.INIT('h1)
	) name11165 (
		_w11695_,
		_w11696_,
		_w11697_
	);
	LUT2 #(
		.INIT('h2)
	) name11166 (
		_w10996_,
		_w11073_,
		_w11698_
	);
	LUT2 #(
		.INIT('h4)
	) name11167 (
		_w10996_,
		_w11073_,
		_w11699_
	);
	LUT2 #(
		.INIT('h1)
	) name11168 (
		_w11698_,
		_w11699_,
		_w11700_
	);
	LUT2 #(
		.INIT('h8)
	) name11169 (
		_w9877_,
		_w11700_,
		_w11701_
	);
	LUT2 #(
		.INIT('h1)
	) name11170 (
		_w9877_,
		_w11700_,
		_w11702_
	);
	LUT2 #(
		.INIT('h1)
	) name11171 (
		_w11701_,
		_w11702_,
		_w11703_
	);
	LUT2 #(
		.INIT('h1)
	) name11172 (
		_w11697_,
		_w11703_,
		_w11704_
	);
	LUT2 #(
		.INIT('h8)
	) name11173 (
		_w11697_,
		_w11703_,
		_w11705_
	);
	LUT2 #(
		.INIT('h1)
	) name11174 (
		\ld_r_reg/P0001 ,
		_w11704_,
		_w11706_
	);
	LUT2 #(
		.INIT('h4)
	) name11175 (
		_w11705_,
		_w11706_,
		_w11707_
	);
	LUT2 #(
		.INIT('h1)
	) name11176 (
		\text_in_r_reg[88]/P0001 ,
		\u0_w_reg[1][24]/P0002 ,
		_w11708_
	);
	LUT2 #(
		.INIT('h8)
	) name11177 (
		\text_in_r_reg[88]/P0001 ,
		\u0_w_reg[1][24]/P0002 ,
		_w11709_
	);
	LUT2 #(
		.INIT('h2)
	) name11178 (
		\ld_r_reg/P0001 ,
		_w11708_,
		_w11710_
	);
	LUT2 #(
		.INIT('h4)
	) name11179 (
		_w11709_,
		_w11710_,
		_w11711_
	);
	LUT2 #(
		.INIT('h1)
	) name11180 (
		_w11707_,
		_w11711_,
		_w11712_
	);
	LUT2 #(
		.INIT('h1)
	) name11181 (
		\u0_w_reg[1][8]/P0001 ,
		_w10344_,
		_w11713_
	);
	LUT2 #(
		.INIT('h8)
	) name11182 (
		\u0_w_reg[1][8]/P0001 ,
		_w10344_,
		_w11714_
	);
	LUT2 #(
		.INIT('h1)
	) name11183 (
		_w11713_,
		_w11714_,
		_w11715_
	);
	LUT2 #(
		.INIT('h2)
	) name11184 (
		_w10248_,
		_w10996_,
		_w11716_
	);
	LUT2 #(
		.INIT('h4)
	) name11185 (
		_w10248_,
		_w10996_,
		_w11717_
	);
	LUT2 #(
		.INIT('h1)
	) name11186 (
		_w11716_,
		_w11717_,
		_w11718_
	);
	LUT2 #(
		.INIT('h8)
	) name11187 (
		_w11682_,
		_w11718_,
		_w11719_
	);
	LUT2 #(
		.INIT('h1)
	) name11188 (
		_w11682_,
		_w11718_,
		_w11720_
	);
	LUT2 #(
		.INIT('h1)
	) name11189 (
		_w11719_,
		_w11720_,
		_w11721_
	);
	LUT2 #(
		.INIT('h1)
	) name11190 (
		_w11715_,
		_w11721_,
		_w11722_
	);
	LUT2 #(
		.INIT('h8)
	) name11191 (
		_w11715_,
		_w11721_,
		_w11723_
	);
	LUT2 #(
		.INIT('h1)
	) name11192 (
		\ld_r_reg/P0001 ,
		_w11722_,
		_w11724_
	);
	LUT2 #(
		.INIT('h4)
	) name11193 (
		_w11723_,
		_w11724_,
		_w11725_
	);
	LUT2 #(
		.INIT('h2)
	) name11194 (
		\text_in_r_reg[72]/P0001 ,
		\u0_w_reg[1][8]/P0001 ,
		_w11726_
	);
	LUT2 #(
		.INIT('h4)
	) name11195 (
		\text_in_r_reg[72]/P0001 ,
		\u0_w_reg[1][8]/P0001 ,
		_w11727_
	);
	LUT2 #(
		.INIT('h2)
	) name11196 (
		\ld_r_reg/P0001 ,
		_w11726_,
		_w11728_
	);
	LUT2 #(
		.INIT('h4)
	) name11197 (
		_w11727_,
		_w11728_,
		_w11729_
	);
	LUT2 #(
		.INIT('h1)
	) name11198 (
		_w11725_,
		_w11729_,
		_w11730_
	);
	LUT2 #(
		.INIT('h1)
	) name11199 (
		_w10508_,
		_w11315_,
		_w11731_
	);
	LUT2 #(
		.INIT('h8)
	) name11200 (
		_w10508_,
		_w11315_,
		_w11732_
	);
	LUT2 #(
		.INIT('h1)
	) name11201 (
		_w11731_,
		_w11732_,
		_w11733_
	);
	LUT2 #(
		.INIT('h2)
	) name11202 (
		\u0_w_reg[1][10]/P0001 ,
		_w11562_,
		_w11734_
	);
	LUT2 #(
		.INIT('h4)
	) name11203 (
		\u0_w_reg[1][10]/P0001 ,
		_w11562_,
		_w11735_
	);
	LUT2 #(
		.INIT('h1)
	) name11204 (
		_w11734_,
		_w11735_,
		_w11736_
	);
	LUT2 #(
		.INIT('h8)
	) name11205 (
		_w11155_,
		_w11736_,
		_w11737_
	);
	LUT2 #(
		.INIT('h1)
	) name11206 (
		_w11155_,
		_w11736_,
		_w11738_
	);
	LUT2 #(
		.INIT('h1)
	) name11207 (
		_w11737_,
		_w11738_,
		_w11739_
	);
	LUT2 #(
		.INIT('h1)
	) name11208 (
		_w11733_,
		_w11739_,
		_w11740_
	);
	LUT2 #(
		.INIT('h8)
	) name11209 (
		_w11733_,
		_w11739_,
		_w11741_
	);
	LUT2 #(
		.INIT('h1)
	) name11210 (
		\ld_r_reg/P0001 ,
		_w11740_,
		_w11742_
	);
	LUT2 #(
		.INIT('h4)
	) name11211 (
		_w11741_,
		_w11742_,
		_w11743_
	);
	LUT2 #(
		.INIT('h2)
	) name11212 (
		\text_in_r_reg[74]/P0001 ,
		\u0_w_reg[1][10]/P0001 ,
		_w11744_
	);
	LUT2 #(
		.INIT('h4)
	) name11213 (
		\text_in_r_reg[74]/P0001 ,
		\u0_w_reg[1][10]/P0001 ,
		_w11745_
	);
	LUT2 #(
		.INIT('h2)
	) name11214 (
		\ld_r_reg/P0001 ,
		_w11744_,
		_w11746_
	);
	LUT2 #(
		.INIT('h4)
	) name11215 (
		_w11745_,
		_w11746_,
		_w11747_
	);
	LUT2 #(
		.INIT('h1)
	) name11216 (
		_w11743_,
		_w11747_,
		_w11748_
	);
	LUT2 #(
		.INIT('h2)
	) name11217 (
		\u0_w_reg[1][3]/P0001 ,
		_w10775_,
		_w11749_
	);
	LUT2 #(
		.INIT('h4)
	) name11218 (
		\u0_w_reg[1][3]/P0001 ,
		_w10775_,
		_w11750_
	);
	LUT2 #(
		.INIT('h1)
	) name11219 (
		_w11749_,
		_w11750_,
		_w11751_
	);
	LUT2 #(
		.INIT('h8)
	) name11220 (
		_w11565_,
		_w11751_,
		_w11752_
	);
	LUT2 #(
		.INIT('h1)
	) name11221 (
		_w11565_,
		_w11751_,
		_w11753_
	);
	LUT2 #(
		.INIT('h1)
	) name11222 (
		_w11752_,
		_w11753_,
		_w11754_
	);
	LUT2 #(
		.INIT('h8)
	) name11223 (
		_w11450_,
		_w11489_,
		_w11755_
	);
	LUT2 #(
		.INIT('h1)
	) name11224 (
		_w11450_,
		_w11489_,
		_w11756_
	);
	LUT2 #(
		.INIT('h1)
	) name11225 (
		_w11755_,
		_w11756_,
		_w11757_
	);
	LUT2 #(
		.INIT('h1)
	) name11226 (
		_w11754_,
		_w11757_,
		_w11758_
	);
	LUT2 #(
		.INIT('h8)
	) name11227 (
		_w11754_,
		_w11757_,
		_w11759_
	);
	LUT2 #(
		.INIT('h1)
	) name11228 (
		\ld_r_reg/P0001 ,
		_w11758_,
		_w11760_
	);
	LUT2 #(
		.INIT('h4)
	) name11229 (
		_w11759_,
		_w11760_,
		_w11761_
	);
	LUT2 #(
		.INIT('h2)
	) name11230 (
		\text_in_r_reg[67]/P0001 ,
		\u0_w_reg[1][3]/P0001 ,
		_w11762_
	);
	LUT2 #(
		.INIT('h4)
	) name11231 (
		\text_in_r_reg[67]/P0001 ,
		\u0_w_reg[1][3]/P0001 ,
		_w11763_
	);
	LUT2 #(
		.INIT('h2)
	) name11232 (
		\ld_r_reg/P0001 ,
		_w11762_,
		_w11764_
	);
	LUT2 #(
		.INIT('h4)
	) name11233 (
		_w11763_,
		_w11764_,
		_w11765_
	);
	LUT2 #(
		.INIT('h1)
	) name11234 (
		_w11761_,
		_w11765_,
		_w11766_
	);
	LUT2 #(
		.INIT('h1)
	) name11235 (
		\u0_w_reg[1][5]/P0001 ,
		_w8853_,
		_w11767_
	);
	LUT2 #(
		.INIT('h8)
	) name11236 (
		\u0_w_reg[1][5]/P0001 ,
		_w8853_,
		_w11768_
	);
	LUT2 #(
		.INIT('h1)
	) name11237 (
		_w11767_,
		_w11768_,
		_w11769_
	);
	LUT2 #(
		.INIT('h1)
	) name11238 (
		\u0_w_reg[1][6]/P0001 ,
		_w8974_,
		_w11770_
	);
	LUT2 #(
		.INIT('h8)
	) name11239 (
		\u0_w_reg[1][6]/P0001 ,
		_w8974_,
		_w11771_
	);
	LUT2 #(
		.INIT('h1)
	) name11240 (
		_w11770_,
		_w11771_,
		_w11772_
	);
	LUT2 #(
		.INIT('h1)
	) name11241 (
		\u0_w_reg[1][4]/P0001 ,
		_w9639_,
		_w11773_
	);
	LUT2 #(
		.INIT('h8)
	) name11242 (
		\u0_w_reg[1][4]/P0001 ,
		_w9639_,
		_w11774_
	);
	LUT2 #(
		.INIT('h1)
	) name11243 (
		_w11773_,
		_w11774_,
		_w11775_
	);
	LUT2 #(
		.INIT('h1)
	) name11244 (
		\u0_w_reg[1][0]/P0001 ,
		_w10344_,
		_w11776_
	);
	LUT2 #(
		.INIT('h8)
	) name11245 (
		\u0_w_reg[1][0]/P0001 ,
		_w10344_,
		_w11777_
	);
	LUT2 #(
		.INIT('h1)
	) name11246 (
		_w11776_,
		_w11777_,
		_w11778_
	);
	LUT2 #(
		.INIT('h1)
	) name11247 (
		\u0_w_reg[1][3]/P0001 ,
		_w10898_,
		_w11779_
	);
	LUT2 #(
		.INIT('h8)
	) name11248 (
		\u0_w_reg[1][3]/P0001 ,
		_w10898_,
		_w11780_
	);
	LUT2 #(
		.INIT('h1)
	) name11249 (
		_w11779_,
		_w11780_,
		_w11781_
	);
	LUT2 #(
		.INIT('h1)
	) name11250 (
		\u0_w_reg[1][1]/P0001 ,
		_w11155_,
		_w11782_
	);
	LUT2 #(
		.INIT('h8)
	) name11251 (
		\u0_w_reg[1][1]/P0001 ,
		_w11155_,
		_w11783_
	);
	LUT2 #(
		.INIT('h1)
	) name11252 (
		_w11782_,
		_w11783_,
		_w11784_
	);
	LUT2 #(
		.INIT('h1)
	) name11253 (
		\u0_w_reg[1][2]/P0001 ,
		_w11562_,
		_w11785_
	);
	LUT2 #(
		.INIT('h8)
	) name11254 (
		\u0_w_reg[1][2]/P0001 ,
		_w11562_,
		_w11786_
	);
	LUT2 #(
		.INIT('h1)
	) name11255 (
		_w11785_,
		_w11786_,
		_w11787_
	);
	LUT2 #(
		.INIT('h1)
	) name11256 (
		\u0_w_reg[1][7]/P0001 ,
		_w10430_,
		_w11788_
	);
	LUT2 #(
		.INIT('h8)
	) name11257 (
		\u0_w_reg[1][7]/P0001 ,
		_w10430_,
		_w11789_
	);
	LUT2 #(
		.INIT('h1)
	) name11258 (
		_w11788_,
		_w11789_,
		_w11790_
	);
	LUT2 #(
		.INIT('h2)
	) name11259 (
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w11791_
	);
	LUT2 #(
		.INIT('h8)
	) name11260 (
		\sa11_reg[5]/P0001 ,
		_w11791_,
		_w11792_
	);
	LUT2 #(
		.INIT('h8)
	) name11261 (
		\sa11_reg[2]/P0001 ,
		_w11792_,
		_w11793_
	);
	LUT2 #(
		.INIT('h8)
	) name11262 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w11794_
	);
	LUT2 #(
		.INIT('h8)
	) name11263 (
		_w11791_,
		_w11794_,
		_w11795_
	);
	LUT2 #(
		.INIT('h2)
	) name11264 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w11796_
	);
	LUT2 #(
		.INIT('h2)
	) name11265 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w11797_
	);
	LUT2 #(
		.INIT('h8)
	) name11266 (
		\sa11_reg[7]/NET0131 ,
		_w11797_,
		_w11798_
	);
	LUT2 #(
		.INIT('h4)
	) name11267 (
		_w11796_,
		_w11798_,
		_w11799_
	);
	LUT2 #(
		.INIT('h1)
	) name11268 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w11800_
	);
	LUT2 #(
		.INIT('h4)
	) name11269 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w11801_
	);
	LUT2 #(
		.INIT('h8)
	) name11270 (
		_w11800_,
		_w11801_,
		_w11802_
	);
	LUT2 #(
		.INIT('h1)
	) name11271 (
		_w11799_,
		_w11802_,
		_w11803_
	);
	LUT2 #(
		.INIT('h1)
	) name11272 (
		\sa11_reg[2]/P0001 ,
		_w11803_,
		_w11804_
	);
	LUT2 #(
		.INIT('h2)
	) name11273 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w11805_
	);
	LUT2 #(
		.INIT('h8)
	) name11274 (
		\sa11_reg[4]/P0001 ,
		_w11801_,
		_w11806_
	);
	LUT2 #(
		.INIT('h8)
	) name11275 (
		_w11805_,
		_w11806_,
		_w11807_
	);
	LUT2 #(
		.INIT('h1)
	) name11276 (
		_w11793_,
		_w11795_,
		_w11808_
	);
	LUT2 #(
		.INIT('h4)
	) name11277 (
		_w11807_,
		_w11808_,
		_w11809_
	);
	LUT2 #(
		.INIT('h4)
	) name11278 (
		_w11804_,
		_w11809_,
		_w11810_
	);
	LUT2 #(
		.INIT('h2)
	) name11279 (
		\sa11_reg[1]/P0001 ,
		_w11810_,
		_w11811_
	);
	LUT2 #(
		.INIT('h1)
	) name11280 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w11812_
	);
	LUT2 #(
		.INIT('h8)
	) name11281 (
		\sa11_reg[4]/P0001 ,
		_w11812_,
		_w11813_
	);
	LUT2 #(
		.INIT('h8)
	) name11282 (
		\sa11_reg[3]/P0001 ,
		_w11813_,
		_w11814_
	);
	LUT2 #(
		.INIT('h4)
	) name11283 (
		\sa11_reg[6]/NET0131 ,
		_w11814_,
		_w11815_
	);
	LUT2 #(
		.INIT('h4)
	) name11284 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w11816_
	);
	LUT2 #(
		.INIT('h4)
	) name11285 (
		\sa11_reg[4]/P0001 ,
		_w11816_,
		_w11817_
	);
	LUT2 #(
		.INIT('h4)
	) name11286 (
		\sa11_reg[3]/P0001 ,
		_w11817_,
		_w11818_
	);
	LUT2 #(
		.INIT('h1)
	) name11287 (
		_w11815_,
		_w11818_,
		_w11819_
	);
	LUT2 #(
		.INIT('h2)
	) name11288 (
		\sa11_reg[2]/P0001 ,
		_w11819_,
		_w11820_
	);
	LUT2 #(
		.INIT('h8)
	) name11289 (
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w11821_
	);
	LUT2 #(
		.INIT('h4)
	) name11290 (
		\sa11_reg[5]/P0001 ,
		_w11821_,
		_w11822_
	);
	LUT2 #(
		.INIT('h4)
	) name11291 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w11823_
	);
	LUT2 #(
		.INIT('h8)
	) name11292 (
		_w11822_,
		_w11823_,
		_w11824_
	);
	LUT2 #(
		.INIT('h2)
	) name11293 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w11825_
	);
	LUT2 #(
		.INIT('h8)
	) name11294 (
		_w11800_,
		_w11825_,
		_w11826_
	);
	LUT2 #(
		.INIT('h1)
	) name11295 (
		_w11824_,
		_w11826_,
		_w11827_
	);
	LUT2 #(
		.INIT('h1)
	) name11296 (
		\sa11_reg[3]/P0001 ,
		_w11827_,
		_w11828_
	);
	LUT2 #(
		.INIT('h1)
	) name11297 (
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w11829_
	);
	LUT2 #(
		.INIT('h8)
	) name11298 (
		_w11796_,
		_w11829_,
		_w11830_
	);
	LUT2 #(
		.INIT('h2)
	) name11299 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w11831_
	);
	LUT2 #(
		.INIT('h8)
	) name11300 (
		_w11812_,
		_w11831_,
		_w11832_
	);
	LUT2 #(
		.INIT('h8)
	) name11301 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w11833_
	);
	LUT2 #(
		.INIT('h8)
	) name11302 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w11834_
	);
	LUT2 #(
		.INIT('h8)
	) name11303 (
		_w11833_,
		_w11834_,
		_w11835_
	);
	LUT2 #(
		.INIT('h4)
	) name11304 (
		\sa11_reg[3]/P0001 ,
		_w11792_,
		_w11836_
	);
	LUT2 #(
		.INIT('h4)
	) name11305 (
		\sa11_reg[2]/P0001 ,
		_w11836_,
		_w11837_
	);
	LUT2 #(
		.INIT('h1)
	) name11306 (
		_w11830_,
		_w11832_,
		_w11838_
	);
	LUT2 #(
		.INIT('h4)
	) name11307 (
		_w11835_,
		_w11838_,
		_w11839_
	);
	LUT2 #(
		.INIT('h4)
	) name11308 (
		_w11837_,
		_w11839_,
		_w11840_
	);
	LUT2 #(
		.INIT('h1)
	) name11309 (
		\sa11_reg[1]/P0001 ,
		_w11840_,
		_w11841_
	);
	LUT2 #(
		.INIT('h1)
	) name11310 (
		_w11820_,
		_w11828_,
		_w11842_
	);
	LUT2 #(
		.INIT('h4)
	) name11311 (
		_w11841_,
		_w11842_,
		_w11843_
	);
	LUT2 #(
		.INIT('h4)
	) name11312 (
		_w11811_,
		_w11843_,
		_w11844_
	);
	LUT2 #(
		.INIT('h1)
	) name11313 (
		\sa11_reg[0]/P0001 ,
		_w11844_,
		_w11845_
	);
	LUT2 #(
		.INIT('h8)
	) name11314 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w11846_
	);
	LUT2 #(
		.INIT('h8)
	) name11315 (
		\sa11_reg[5]/P0001 ,
		_w11829_,
		_w11847_
	);
	LUT2 #(
		.INIT('h8)
	) name11316 (
		_w11846_,
		_w11847_,
		_w11848_
	);
	LUT2 #(
		.INIT('h8)
	) name11317 (
		_w11791_,
		_w11805_,
		_w11849_
	);
	LUT2 #(
		.INIT('h8)
	) name11318 (
		\sa11_reg[4]/P0001 ,
		_w11849_,
		_w11850_
	);
	LUT2 #(
		.INIT('h1)
	) name11319 (
		_w11848_,
		_w11850_,
		_w11851_
	);
	LUT2 #(
		.INIT('h2)
	) name11320 (
		\sa11_reg[1]/P0001 ,
		_w11851_,
		_w11852_
	);
	LUT2 #(
		.INIT('h4)
	) name11321 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w11853_
	);
	LUT2 #(
		.INIT('h8)
	) name11322 (
		_w11812_,
		_w11853_,
		_w11854_
	);
	LUT2 #(
		.INIT('h4)
	) name11323 (
		\sa11_reg[2]/P0001 ,
		_w11854_,
		_w11855_
	);
	LUT2 #(
		.INIT('h1)
	) name11324 (
		_w11835_,
		_w11855_,
		_w11856_
	);
	LUT2 #(
		.INIT('h2)
	) name11325 (
		\sa11_reg[3]/P0001 ,
		_w11856_,
		_w11857_
	);
	LUT2 #(
		.INIT('h8)
	) name11326 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w11858_
	);
	LUT2 #(
		.INIT('h8)
	) name11327 (
		_w11806_,
		_w11858_,
		_w11859_
	);
	LUT2 #(
		.INIT('h1)
	) name11328 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w11860_
	);
	LUT2 #(
		.INIT('h8)
	) name11329 (
		\sa11_reg[7]/NET0131 ,
		_w11860_,
		_w11861_
	);
	LUT2 #(
		.INIT('h8)
	) name11330 (
		_w11833_,
		_w11861_,
		_w11862_
	);
	LUT2 #(
		.INIT('h2)
	) name11331 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		_w11863_
	);
	LUT2 #(
		.INIT('h4)
	) name11332 (
		_w11829_,
		_w11863_,
		_w11864_
	);
	LUT2 #(
		.INIT('h8)
	) name11333 (
		_w11829_,
		_w11860_,
		_w11865_
	);
	LUT2 #(
		.INIT('h4)
	) name11334 (
		\sa11_reg[5]/P0001 ,
		_w11865_,
		_w11866_
	);
	LUT2 #(
		.INIT('h1)
	) name11335 (
		_w11862_,
		_w11864_,
		_w11867_
	);
	LUT2 #(
		.INIT('h4)
	) name11336 (
		_w11866_,
		_w11867_,
		_w11868_
	);
	LUT2 #(
		.INIT('h1)
	) name11337 (
		\sa11_reg[2]/P0001 ,
		_w11868_,
		_w11869_
	);
	LUT2 #(
		.INIT('h4)
	) name11338 (
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w11870_
	);
	LUT2 #(
		.INIT('h4)
	) name11339 (
		\sa11_reg[5]/P0001 ,
		_w11870_,
		_w11871_
	);
	LUT2 #(
		.INIT('h8)
	) name11340 (
		_w11796_,
		_w11871_,
		_w11872_
	);
	LUT2 #(
		.INIT('h1)
	) name11341 (
		_w11859_,
		_w11872_,
		_w11873_
	);
	LUT2 #(
		.INIT('h4)
	) name11342 (
		_w11869_,
		_w11873_,
		_w11874_
	);
	LUT2 #(
		.INIT('h2)
	) name11343 (
		\sa11_reg[1]/P0001 ,
		_w11874_,
		_w11875_
	);
	LUT2 #(
		.INIT('h1)
	) name11344 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w11876_
	);
	LUT2 #(
		.INIT('h4)
	) name11345 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w11877_
	);
	LUT2 #(
		.INIT('h4)
	) name11346 (
		\sa11_reg[7]/NET0131 ,
		_w11877_,
		_w11878_
	);
	LUT2 #(
		.INIT('h8)
	) name11347 (
		_w11876_,
		_w11878_,
		_w11879_
	);
	LUT2 #(
		.INIT('h4)
	) name11348 (
		\sa11_reg[6]/NET0131 ,
		_w11796_,
		_w11880_
	);
	LUT2 #(
		.INIT('h8)
	) name11349 (
		_w11825_,
		_w11880_,
		_w11881_
	);
	LUT2 #(
		.INIT('h4)
	) name11350 (
		\sa11_reg[4]/P0001 ,
		_w11791_,
		_w11882_
	);
	LUT2 #(
		.INIT('h8)
	) name11351 (
		\sa11_reg[4]/P0001 ,
		_w11871_,
		_w11883_
	);
	LUT2 #(
		.INIT('h1)
	) name11352 (
		_w11882_,
		_w11883_,
		_w11884_
	);
	LUT2 #(
		.INIT('h1)
	) name11353 (
		\sa11_reg[2]/P0001 ,
		_w11884_,
		_w11885_
	);
	LUT2 #(
		.INIT('h4)
	) name11354 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w11886_
	);
	LUT2 #(
		.INIT('h8)
	) name11355 (
		_w11831_,
		_w11886_,
		_w11887_
	);
	LUT2 #(
		.INIT('h2)
	) name11356 (
		\sa11_reg[1]/P0001 ,
		_w11887_,
		_w11888_
	);
	LUT2 #(
		.INIT('h4)
	) name11357 (
		_w11879_,
		_w11888_,
		_w11889_
	);
	LUT2 #(
		.INIT('h4)
	) name11358 (
		_w11881_,
		_w11889_,
		_w11890_
	);
	LUT2 #(
		.INIT('h4)
	) name11359 (
		_w11885_,
		_w11890_,
		_w11891_
	);
	LUT2 #(
		.INIT('h8)
	) name11360 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w11892_
	);
	LUT2 #(
		.INIT('h1)
	) name11361 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w11893_
	);
	LUT2 #(
		.INIT('h1)
	) name11362 (
		\sa11_reg[3]/P0001 ,
		_w11893_,
		_w11894_
	);
	LUT2 #(
		.INIT('h2)
	) name11363 (
		_w11892_,
		_w11894_,
		_w11895_
	);
	LUT2 #(
		.INIT('h8)
	) name11364 (
		_w11858_,
		_w11886_,
		_w11896_
	);
	LUT2 #(
		.INIT('h1)
	) name11365 (
		\sa11_reg[1]/P0001 ,
		_w11896_,
		_w11897_
	);
	LUT2 #(
		.INIT('h8)
	) name11366 (
		\sa11_reg[4]/P0001 ,
		_w11798_,
		_w11898_
	);
	LUT2 #(
		.INIT('h8)
	) name11367 (
		\sa11_reg[2]/P0001 ,
		_w11898_,
		_w11899_
	);
	LUT2 #(
		.INIT('h4)
	) name11368 (
		\sa11_reg[6]/NET0131 ,
		_w11794_,
		_w11900_
	);
	LUT2 #(
		.INIT('h4)
	) name11369 (
		\sa11_reg[7]/NET0131 ,
		_w11900_,
		_w11901_
	);
	LUT2 #(
		.INIT('h4)
	) name11370 (
		\sa11_reg[2]/P0001 ,
		_w11901_,
		_w11902_
	);
	LUT2 #(
		.INIT('h4)
	) name11371 (
		_w11895_,
		_w11897_,
		_w11903_
	);
	LUT2 #(
		.INIT('h4)
	) name11372 (
		_w11899_,
		_w11903_,
		_w11904_
	);
	LUT2 #(
		.INIT('h4)
	) name11373 (
		_w11902_,
		_w11904_,
		_w11905_
	);
	LUT2 #(
		.INIT('h1)
	) name11374 (
		_w11891_,
		_w11905_,
		_w11906_
	);
	LUT2 #(
		.INIT('h8)
	) name11375 (
		_w11853_,
		_w11892_,
		_w11907_
	);
	LUT2 #(
		.INIT('h2)
	) name11376 (
		\sa11_reg[2]/P0001 ,
		_w11907_,
		_w11908_
	);
	LUT2 #(
		.INIT('h8)
	) name11377 (
		_w11863_,
		_w11870_,
		_w11909_
	);
	LUT2 #(
		.INIT('h1)
	) name11378 (
		_w11878_,
		_w11880_,
		_w11910_
	);
	LUT2 #(
		.INIT('h4)
	) name11379 (
		_w11909_,
		_w11910_,
		_w11911_
	);
	LUT2 #(
		.INIT('h8)
	) name11380 (
		_w11908_,
		_w11911_,
		_w11912_
	);
	LUT2 #(
		.INIT('h8)
	) name11381 (
		_w11801_,
		_w11858_,
		_w11913_
	);
	LUT2 #(
		.INIT('h1)
	) name11382 (
		\sa11_reg[2]/P0001 ,
		_w11913_,
		_w11914_
	);
	LUT2 #(
		.INIT('h8)
	) name11383 (
		_w11791_,
		_w11796_,
		_w11915_
	);
	LUT2 #(
		.INIT('h1)
	) name11384 (
		_w11866_,
		_w11915_,
		_w11916_
	);
	LUT2 #(
		.INIT('h8)
	) name11385 (
		_w11914_,
		_w11916_,
		_w11917_
	);
	LUT2 #(
		.INIT('h1)
	) name11386 (
		_w11912_,
		_w11917_,
		_w11918_
	);
	LUT2 #(
		.INIT('h1)
	) name11387 (
		_w11906_,
		_w11918_,
		_w11919_
	);
	LUT2 #(
		.INIT('h2)
	) name11388 (
		\sa11_reg[0]/P0001 ,
		_w11919_,
		_w11920_
	);
	LUT2 #(
		.INIT('h4)
	) name11389 (
		\sa11_reg[3]/P0001 ,
		_w11802_,
		_w11921_
	);
	LUT2 #(
		.INIT('h4)
	) name11390 (
		\sa11_reg[3]/P0001 ,
		_w11847_,
		_w11922_
	);
	LUT2 #(
		.INIT('h8)
	) name11391 (
		\sa11_reg[5]/P0001 ,
		_w11796_,
		_w11923_
	);
	LUT2 #(
		.INIT('h4)
	) name11392 (
		\sa11_reg[6]/NET0131 ,
		_w11923_,
		_w11924_
	);
	LUT2 #(
		.INIT('h8)
	) name11393 (
		_w11825_,
		_w11858_,
		_w11925_
	);
	LUT2 #(
		.INIT('h8)
	) name11394 (
		\sa11_reg[7]/NET0131 ,
		_w11794_,
		_w11926_
	);
	LUT2 #(
		.INIT('h8)
	) name11395 (
		_w11876_,
		_w11926_,
		_w11927_
	);
	LUT2 #(
		.INIT('h2)
	) name11396 (
		\sa11_reg[2]/P0001 ,
		_w11925_,
		_w11928_
	);
	LUT2 #(
		.INIT('h4)
	) name11397 (
		_w11921_,
		_w11928_,
		_w11929_
	);
	LUT2 #(
		.INIT('h1)
	) name11398 (
		_w11922_,
		_w11924_,
		_w11930_
	);
	LUT2 #(
		.INIT('h4)
	) name11399 (
		_w11927_,
		_w11930_,
		_w11931_
	);
	LUT2 #(
		.INIT('h8)
	) name11400 (
		_w11929_,
		_w11931_,
		_w11932_
	);
	LUT2 #(
		.INIT('h8)
	) name11401 (
		\sa11_reg[7]/NET0131 ,
		_w11833_,
		_w11933_
	);
	LUT2 #(
		.INIT('h8)
	) name11402 (
		_w11796_,
		_w11933_,
		_w11934_
	);
	LUT2 #(
		.INIT('h4)
	) name11403 (
		\sa11_reg[3]/P0001 ,
		_w11822_,
		_w11935_
	);
	LUT2 #(
		.INIT('h8)
	) name11404 (
		_w11816_,
		_w11877_,
		_w11936_
	);
	LUT2 #(
		.INIT('h1)
	) name11405 (
		\sa11_reg[2]/P0001 ,
		_w11936_,
		_w11937_
	);
	LUT2 #(
		.INIT('h4)
	) name11406 (
		_w11934_,
		_w11937_,
		_w11938_
	);
	LUT2 #(
		.INIT('h4)
	) name11407 (
		_w11935_,
		_w11938_,
		_w11939_
	);
	LUT2 #(
		.INIT('h1)
	) name11408 (
		_w11932_,
		_w11939_,
		_w11940_
	);
	LUT2 #(
		.INIT('h8)
	) name11409 (
		_w11792_,
		_w11794_,
		_w11941_
	);
	LUT2 #(
		.INIT('h8)
	) name11410 (
		_w11825_,
		_w11860_,
		_w11942_
	);
	LUT2 #(
		.INIT('h4)
	) name11411 (
		\sa11_reg[6]/NET0131 ,
		_w11942_,
		_w11943_
	);
	LUT2 #(
		.INIT('h1)
	) name11412 (
		_w11941_,
		_w11943_,
		_w11944_
	);
	LUT2 #(
		.INIT('h4)
	) name11413 (
		_w11940_,
		_w11944_,
		_w11945_
	);
	LUT2 #(
		.INIT('h1)
	) name11414 (
		\sa11_reg[1]/P0001 ,
		_w11945_,
		_w11946_
	);
	LUT2 #(
		.INIT('h1)
	) name11415 (
		_w11852_,
		_w11857_,
		_w11947_
	);
	LUT2 #(
		.INIT('h4)
	) name11416 (
		_w11875_,
		_w11947_,
		_w11948_
	);
	LUT2 #(
		.INIT('h4)
	) name11417 (
		_w11920_,
		_w11948_,
		_w11949_
	);
	LUT2 #(
		.INIT('h4)
	) name11418 (
		_w11946_,
		_w11949_,
		_w11950_
	);
	LUT2 #(
		.INIT('h4)
	) name11419 (
		_w11845_,
		_w11950_,
		_w11951_
	);
	LUT2 #(
		.INIT('h4)
	) name11420 (
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w11952_
	);
	LUT2 #(
		.INIT('h2)
	) name11421 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w11953_
	);
	LUT2 #(
		.INIT('h8)
	) name11422 (
		_w11952_,
		_w11953_,
		_w11954_
	);
	LUT2 #(
		.INIT('h4)
	) name11423 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w11955_
	);
	LUT2 #(
		.INIT('h1)
	) name11424 (
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w11956_
	);
	LUT2 #(
		.INIT('h4)
	) name11425 (
		\sa00_reg[5]/P0001 ,
		_w11956_,
		_w11957_
	);
	LUT2 #(
		.INIT('h8)
	) name11426 (
		_w11955_,
		_w11957_,
		_w11958_
	);
	LUT2 #(
		.INIT('h8)
	) name11427 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w11959_
	);
	LUT2 #(
		.INIT('h1)
	) name11428 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w11960_
	);
	LUT2 #(
		.INIT('h8)
	) name11429 (
		_w11959_,
		_w11960_,
		_w11961_
	);
	LUT2 #(
		.INIT('h2)
	) name11430 (
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w11962_
	);
	LUT2 #(
		.INIT('h4)
	) name11431 (
		\sa00_reg[4]/P0001 ,
		_w11962_,
		_w11963_
	);
	LUT2 #(
		.INIT('h1)
	) name11432 (
		_w11961_,
		_w11963_,
		_w11964_
	);
	LUT2 #(
		.INIT('h1)
	) name11433 (
		\sa00_reg[2]/P0001 ,
		_w11964_,
		_w11965_
	);
	LUT2 #(
		.INIT('h2)
	) name11434 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w11966_
	);
	LUT2 #(
		.INIT('h8)
	) name11435 (
		\sa00_reg[5]/P0001 ,
		_w11956_,
		_w11967_
	);
	LUT2 #(
		.INIT('h8)
	) name11436 (
		_w11966_,
		_w11967_,
		_w11968_
	);
	LUT2 #(
		.INIT('h2)
	) name11437 (
		\sa00_reg[1]/P0001 ,
		_w11954_,
		_w11969_
	);
	LUT2 #(
		.INIT('h4)
	) name11438 (
		_w11958_,
		_w11969_,
		_w11970_
	);
	LUT2 #(
		.INIT('h4)
	) name11439 (
		_w11968_,
		_w11970_,
		_w11971_
	);
	LUT2 #(
		.INIT('h4)
	) name11440 (
		_w11965_,
		_w11971_,
		_w11972_
	);
	LUT2 #(
		.INIT('h8)
	) name11441 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w11973_
	);
	LUT2 #(
		.INIT('h8)
	) name11442 (
		\sa00_reg[3]/P0001 ,
		_w11973_,
		_w11974_
	);
	LUT2 #(
		.INIT('h2)
	) name11443 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w11975_
	);
	LUT2 #(
		.INIT('h8)
	) name11444 (
		_w11959_,
		_w11975_,
		_w11976_
	);
	LUT2 #(
		.INIT('h8)
	) name11445 (
		\sa00_reg[2]/P0001 ,
		_w11976_,
		_w11977_
	);
	LUT2 #(
		.INIT('h4)
	) name11446 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w11978_
	);
	LUT2 #(
		.INIT('h8)
	) name11447 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w11979_
	);
	LUT2 #(
		.INIT('h8)
	) name11448 (
		_w11978_,
		_w11979_,
		_w11980_
	);
	LUT2 #(
		.INIT('h1)
	) name11449 (
		\sa00_reg[1]/P0001 ,
		_w11980_,
		_w11981_
	);
	LUT2 #(
		.INIT('h8)
	) name11450 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w11982_
	);
	LUT2 #(
		.INIT('h8)
	) name11451 (
		_w11956_,
		_w11982_,
		_w11983_
	);
	LUT2 #(
		.INIT('h4)
	) name11452 (
		\sa00_reg[2]/P0001 ,
		_w11983_,
		_w11984_
	);
	LUT2 #(
		.INIT('h4)
	) name11453 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w11985_
	);
	LUT2 #(
		.INIT('h8)
	) name11454 (
		_w11978_,
		_w11985_,
		_w11986_
	);
	LUT2 #(
		.INIT('h1)
	) name11455 (
		_w11974_,
		_w11986_,
		_w11987_
	);
	LUT2 #(
		.INIT('h4)
	) name11456 (
		_w11977_,
		_w11987_,
		_w11988_
	);
	LUT2 #(
		.INIT('h2)
	) name11457 (
		_w11981_,
		_w11984_,
		_w11989_
	);
	LUT2 #(
		.INIT('h8)
	) name11458 (
		_w11988_,
		_w11989_,
		_w11990_
	);
	LUT2 #(
		.INIT('h1)
	) name11459 (
		_w11972_,
		_w11990_,
		_w11991_
	);
	LUT2 #(
		.INIT('h2)
	) name11460 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w11992_
	);
	LUT2 #(
		.INIT('h8)
	) name11461 (
		_w11952_,
		_w11992_,
		_w11993_
	);
	LUT2 #(
		.INIT('h4)
	) name11462 (
		\sa00_reg[6]/NET0131 ,
		_w11966_,
		_w11994_
	);
	LUT2 #(
		.INIT('h8)
	) name11463 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w11995_
	);
	LUT2 #(
		.INIT('h8)
	) name11464 (
		\sa00_reg[7]/NET0131 ,
		_w11995_,
		_w11996_
	);
	LUT2 #(
		.INIT('h1)
	) name11465 (
		_w11955_,
		_w11996_,
		_w11997_
	);
	LUT2 #(
		.INIT('h1)
	) name11466 (
		_w11959_,
		_w11997_,
		_w11998_
	);
	LUT2 #(
		.INIT('h2)
	) name11467 (
		\sa00_reg[2]/P0001 ,
		_w11993_,
		_w11999_
	);
	LUT2 #(
		.INIT('h4)
	) name11468 (
		_w11994_,
		_w11999_,
		_w12000_
	);
	LUT2 #(
		.INIT('h4)
	) name11469 (
		_w11998_,
		_w12000_,
		_w12001_
	);
	LUT2 #(
		.INIT('h8)
	) name11470 (
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w12002_
	);
	LUT2 #(
		.INIT('h8)
	) name11471 (
		_w11992_,
		_w12002_,
		_w12003_
	);
	LUT2 #(
		.INIT('h1)
	) name11472 (
		\sa00_reg[2]/P0001 ,
		_w12003_,
		_w12004_
	);
	LUT2 #(
		.INIT('h1)
	) name11473 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w12005_
	);
	LUT2 #(
		.INIT('h8)
	) name11474 (
		_w11957_,
		_w12005_,
		_w12006_
	);
	LUT2 #(
		.INIT('h1)
	) name11475 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w12007_
	);
	LUT2 #(
		.INIT('h8)
	) name11476 (
		_w11979_,
		_w12007_,
		_w12008_
	);
	LUT2 #(
		.INIT('h2)
	) name11477 (
		_w12004_,
		_w12008_,
		_w12009_
	);
	LUT2 #(
		.INIT('h4)
	) name11478 (
		_w12006_,
		_w12009_,
		_w12010_
	);
	LUT2 #(
		.INIT('h1)
	) name11479 (
		_w12001_,
		_w12010_,
		_w12011_
	);
	LUT2 #(
		.INIT('h1)
	) name11480 (
		_w11991_,
		_w12011_,
		_w12012_
	);
	LUT2 #(
		.INIT('h2)
	) name11481 (
		\sa00_reg[0]/P0001 ,
		_w12012_,
		_w12013_
	);
	LUT2 #(
		.INIT('h4)
	) name11482 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w12014_
	);
	LUT2 #(
		.INIT('h4)
	) name11483 (
		\sa00_reg[3]/P0001 ,
		_w11956_,
		_w12015_
	);
	LUT2 #(
		.INIT('h8)
	) name11484 (
		_w12014_,
		_w12015_,
		_w12016_
	);
	LUT2 #(
		.INIT('h8)
	) name11485 (
		_w11962_,
		_w11982_,
		_w12017_
	);
	LUT2 #(
		.INIT('h8)
	) name11486 (
		\sa00_reg[5]/P0001 ,
		_w12017_,
		_w12018_
	);
	LUT2 #(
		.INIT('h8)
	) name11487 (
		_w11966_,
		_w11975_,
		_w12019_
	);
	LUT2 #(
		.INIT('h1)
	) name11488 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w12020_
	);
	LUT2 #(
		.INIT('h8)
	) name11489 (
		_w11978_,
		_w12020_,
		_w12021_
	);
	LUT2 #(
		.INIT('h4)
	) name11490 (
		\sa00_reg[6]/NET0131 ,
		_w12021_,
		_w12022_
	);
	LUT2 #(
		.INIT('h4)
	) name11491 (
		\sa00_reg[3]/P0001 ,
		_w11967_,
		_w12023_
	);
	LUT2 #(
		.INIT('h8)
	) name11492 (
		\sa00_reg[3]/P0001 ,
		_w11960_,
		_w12024_
	);
	LUT2 #(
		.INIT('h8)
	) name11493 (
		_w11959_,
		_w12024_,
		_w12025_
	);
	LUT2 #(
		.INIT('h2)
	) name11494 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w12026_
	);
	LUT2 #(
		.INIT('h8)
	) name11495 (
		_w11979_,
		_w12026_,
		_w12027_
	);
	LUT2 #(
		.INIT('h2)
	) name11496 (
		\sa00_reg[2]/P0001 ,
		_w12019_,
		_w12028_
	);
	LUT2 #(
		.INIT('h4)
	) name11497 (
		_w12027_,
		_w12028_,
		_w12029_
	);
	LUT2 #(
		.INIT('h1)
	) name11498 (
		_w12022_,
		_w12023_,
		_w12030_
	);
	LUT2 #(
		.INIT('h4)
	) name11499 (
		_w12025_,
		_w12030_,
		_w12031_
	);
	LUT2 #(
		.INIT('h8)
	) name11500 (
		_w12029_,
		_w12031_,
		_w12032_
	);
	LUT2 #(
		.INIT('h8)
	) name11501 (
		_w12002_,
		_w12020_,
		_w12033_
	);
	LUT2 #(
		.INIT('h8)
	) name11502 (
		_w11966_,
		_w11996_,
		_w12034_
	);
	LUT2 #(
		.INIT('h4)
	) name11503 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w12035_
	);
	LUT2 #(
		.INIT('h8)
	) name11504 (
		_w11955_,
		_w12035_,
		_w12036_
	);
	LUT2 #(
		.INIT('h1)
	) name11505 (
		\sa00_reg[2]/P0001 ,
		_w12033_,
		_w12037_
	);
	LUT2 #(
		.INIT('h4)
	) name11506 (
		_w12036_,
		_w12037_,
		_w12038_
	);
	LUT2 #(
		.INIT('h4)
	) name11507 (
		_w12034_,
		_w12038_,
		_w12039_
	);
	LUT2 #(
		.INIT('h1)
	) name11508 (
		_w12032_,
		_w12039_,
		_w12040_
	);
	LUT2 #(
		.INIT('h1)
	) name11509 (
		_w12016_,
		_w12018_,
		_w12041_
	);
	LUT2 #(
		.INIT('h4)
	) name11510 (
		_w12040_,
		_w12041_,
		_w12042_
	);
	LUT2 #(
		.INIT('h1)
	) name11511 (
		\sa00_reg[1]/P0001 ,
		_w12042_,
		_w12043_
	);
	LUT2 #(
		.INIT('h4)
	) name11512 (
		_w11956_,
		_w11992_,
		_w12044_
	);
	LUT2 #(
		.INIT('h8)
	) name11513 (
		_w12002_,
		_w12005_,
		_w12045_
	);
	LUT2 #(
		.INIT('h8)
	) name11514 (
		\sa00_reg[5]/P0001 ,
		_w12045_,
		_w12046_
	);
	LUT2 #(
		.INIT('h1)
	) name11515 (
		_w12006_,
		_w12044_,
		_w12047_
	);
	LUT2 #(
		.INIT('h4)
	) name11516 (
		_w12046_,
		_w12047_,
		_w12048_
	);
	LUT2 #(
		.INIT('h1)
	) name11517 (
		\sa00_reg[2]/P0001 ,
		_w12048_,
		_w12049_
	);
	LUT2 #(
		.INIT('h8)
	) name11518 (
		\sa00_reg[7]/NET0131 ,
		_w11982_,
		_w12050_
	);
	LUT2 #(
		.INIT('h8)
	) name11519 (
		_w12035_,
		_w12050_,
		_w12051_
	);
	LUT2 #(
		.INIT('h8)
	) name11520 (
		_w11978_,
		_w11992_,
		_w12052_
	);
	LUT2 #(
		.INIT('h4)
	) name11521 (
		\sa00_reg[6]/NET0131 ,
		_w12052_,
		_w12053_
	);
	LUT2 #(
		.INIT('h8)
	) name11522 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		_w12054_
	);
	LUT2 #(
		.INIT('h8)
	) name11523 (
		_w11967_,
		_w12054_,
		_w12055_
	);
	LUT2 #(
		.INIT('h2)
	) name11524 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		_w12056_
	);
	LUT2 #(
		.INIT('h8)
	) name11525 (
		\sa00_reg[4]/P0001 ,
		_w11962_,
		_w12057_
	);
	LUT2 #(
		.INIT('h8)
	) name11526 (
		_w12056_,
		_w12057_,
		_w12058_
	);
	LUT2 #(
		.INIT('h1)
	) name11527 (
		_w12051_,
		_w12053_,
		_w12059_
	);
	LUT2 #(
		.INIT('h1)
	) name11528 (
		_w12055_,
		_w12058_,
		_w12060_
	);
	LUT2 #(
		.INIT('h8)
	) name11529 (
		_w12059_,
		_w12060_,
		_w12061_
	);
	LUT2 #(
		.INIT('h4)
	) name11530 (
		_w12049_,
		_w12061_,
		_w12062_
	);
	LUT2 #(
		.INIT('h2)
	) name11531 (
		\sa00_reg[1]/P0001 ,
		_w12062_,
		_w12063_
	);
	LUT2 #(
		.INIT('h1)
	) name11532 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w12064_
	);
	LUT2 #(
		.INIT('h4)
	) name11533 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w12065_
	);
	LUT2 #(
		.INIT('h8)
	) name11534 (
		_w12064_,
		_w12065_,
		_w12066_
	);
	LUT2 #(
		.INIT('h1)
	) name11535 (
		\sa00_reg[2]/P0001 ,
		_w12066_,
		_w12067_
	);
	LUT2 #(
		.INIT('h8)
	) name11536 (
		\sa00_reg[4]/P0001 ,
		_w11995_,
		_w12068_
	);
	LUT2 #(
		.INIT('h2)
	) name11537 (
		\sa00_reg[2]/P0001 ,
		_w12068_,
		_w12069_
	);
	LUT2 #(
		.INIT('h2)
	) name11538 (
		\sa00_reg[3]/P0001 ,
		_w12067_,
		_w12070_
	);
	LUT2 #(
		.INIT('h4)
	) name11539 (
		_w12069_,
		_w12070_,
		_w12071_
	);
	LUT2 #(
		.INIT('h4)
	) name11540 (
		\sa00_reg[2]/P0001 ,
		_w11995_,
		_w12072_
	);
	LUT2 #(
		.INIT('h4)
	) name11541 (
		\sa00_reg[3]/P0001 ,
		_w12072_,
		_w12073_
	);
	LUT2 #(
		.INIT('h1)
	) name11542 (
		_w11994_,
		_w12073_,
		_w12074_
	);
	LUT2 #(
		.INIT('h1)
	) name11543 (
		\sa00_reg[7]/NET0131 ,
		_w12074_,
		_w12075_
	);
	LUT2 #(
		.INIT('h1)
	) name11544 (
		_w11957_,
		_w12068_,
		_w12076_
	);
	LUT2 #(
		.INIT('h2)
	) name11545 (
		\sa00_reg[2]/P0001 ,
		_w12076_,
		_w12077_
	);
	LUT2 #(
		.INIT('h1)
	) name11546 (
		_w12075_,
		_w12077_,
		_w12078_
	);
	LUT2 #(
		.INIT('h1)
	) name11547 (
		\sa00_reg[1]/P0001 ,
		_w12078_,
		_w12079_
	);
	LUT2 #(
		.INIT('h8)
	) name11548 (
		\sa00_reg[4]/P0001 ,
		_w11956_,
		_w12080_
	);
	LUT2 #(
		.INIT('h8)
	) name11549 (
		_w11992_,
		_w12080_,
		_w12081_
	);
	LUT2 #(
		.INIT('h4)
	) name11550 (
		\sa00_reg[4]/P0001 ,
		_w12035_,
		_w12082_
	);
	LUT2 #(
		.INIT('h4)
	) name11551 (
		\sa00_reg[3]/P0001 ,
		_w12082_,
		_w12083_
	);
	LUT2 #(
		.INIT('h1)
	) name11552 (
		_w12081_,
		_w12083_,
		_w12084_
	);
	LUT2 #(
		.INIT('h2)
	) name11553 (
		\sa00_reg[2]/P0001 ,
		_w12084_,
		_w12085_
	);
	LUT2 #(
		.INIT('h4)
	) name11554 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w12086_
	);
	LUT2 #(
		.INIT('h8)
	) name11555 (
		_w12033_,
		_w12086_,
		_w12087_
	);
	LUT2 #(
		.INIT('h8)
	) name11556 (
		\sa00_reg[5]/P0001 ,
		_w11952_,
		_w12088_
	);
	LUT2 #(
		.INIT('h4)
	) name11557 (
		_w11966_,
		_w12088_,
		_w12089_
	);
	LUT2 #(
		.INIT('h4)
	) name11558 (
		\sa00_reg[5]/P0001 ,
		_w11978_,
		_w12090_
	);
	LUT2 #(
		.INIT('h4)
	) name11559 (
		\sa00_reg[6]/NET0131 ,
		_w12090_,
		_w12091_
	);
	LUT2 #(
		.INIT('h1)
	) name11560 (
		_w12089_,
		_w12091_,
		_w12092_
	);
	LUT2 #(
		.INIT('h1)
	) name11561 (
		\sa00_reg[2]/P0001 ,
		_w12092_,
		_w12093_
	);
	LUT2 #(
		.INIT('h8)
	) name11562 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w12094_
	);
	LUT2 #(
		.INIT('h8)
	) name11563 (
		_w11962_,
		_w12094_,
		_w12095_
	);
	LUT2 #(
		.INIT('h4)
	) name11564 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w12096_
	);
	LUT2 #(
		.INIT('h8)
	) name11565 (
		\sa00_reg[2]/P0001 ,
		_w11955_,
		_w12097_
	);
	LUT2 #(
		.INIT('h8)
	) name11566 (
		_w12096_,
		_w12097_,
		_w12098_
	);
	LUT2 #(
		.INIT('h1)
	) name11567 (
		_w12017_,
		_w12095_,
		_w12099_
	);
	LUT2 #(
		.INIT('h4)
	) name11568 (
		_w12098_,
		_w12099_,
		_w12100_
	);
	LUT2 #(
		.INIT('h4)
	) name11569 (
		_w12093_,
		_w12100_,
		_w12101_
	);
	LUT2 #(
		.INIT('h2)
	) name11570 (
		\sa00_reg[1]/P0001 ,
		_w12101_,
		_w12102_
	);
	LUT2 #(
		.INIT('h1)
	) name11571 (
		_w12016_,
		_w12087_,
		_w12103_
	);
	LUT2 #(
		.INIT('h4)
	) name11572 (
		_w12085_,
		_w12103_,
		_w12104_
	);
	LUT2 #(
		.INIT('h4)
	) name11573 (
		_w12079_,
		_w12104_,
		_w12105_
	);
	LUT2 #(
		.INIT('h4)
	) name11574 (
		_w12102_,
		_w12105_,
		_w12106_
	);
	LUT2 #(
		.INIT('h1)
	) name11575 (
		\sa00_reg[0]/P0001 ,
		_w12106_,
		_w12107_
	);
	LUT2 #(
		.INIT('h1)
	) name11576 (
		_w12063_,
		_w12071_,
		_w12108_
	);
	LUT2 #(
		.INIT('h4)
	) name11577 (
		_w12013_,
		_w12108_,
		_w12109_
	);
	LUT2 #(
		.INIT('h4)
	) name11578 (
		_w12043_,
		_w12109_,
		_w12110_
	);
	LUT2 #(
		.INIT('h4)
	) name11579 (
		_w12107_,
		_w12110_,
		_w12111_
	);
	LUT2 #(
		.INIT('h2)
	) name11580 (
		_w11951_,
		_w12111_,
		_w12112_
	);
	LUT2 #(
		.INIT('h4)
	) name11581 (
		_w11951_,
		_w12111_,
		_w12113_
	);
	LUT2 #(
		.INIT('h1)
	) name11582 (
		_w12112_,
		_w12113_,
		_w12114_
	);
	LUT2 #(
		.INIT('h8)
	) name11583 (
		_w11797_,
		_w11877_,
		_w12115_
	);
	LUT2 #(
		.INIT('h4)
	) name11584 (
		\sa11_reg[3]/P0001 ,
		_w11882_,
		_w12116_
	);
	LUT2 #(
		.INIT('h1)
	) name11585 (
		_w12115_,
		_w12116_,
		_w12117_
	);
	LUT2 #(
		.INIT('h1)
	) name11586 (
		\sa11_reg[2]/P0001 ,
		_w12117_,
		_w12118_
	);
	LUT2 #(
		.INIT('h8)
	) name11587 (
		_w11829_,
		_w11863_,
		_w12119_
	);
	LUT2 #(
		.INIT('h8)
	) name11588 (
		\sa11_reg[3]/P0001 ,
		_w11870_,
		_w12120_
	);
	LUT2 #(
		.INIT('h4)
	) name11589 (
		\sa11_reg[2]/P0001 ,
		_w12120_,
		_w12121_
	);
	LUT2 #(
		.INIT('h1)
	) name11590 (
		_w11853_,
		_w11877_,
		_w12122_
	);
	LUT2 #(
		.INIT('h8)
	) name11591 (
		_w11892_,
		_w12122_,
		_w12123_
	);
	LUT2 #(
		.INIT('h8)
	) name11592 (
		_w11833_,
		_w11860_,
		_w12124_
	);
	LUT2 #(
		.INIT('h4)
	) name11593 (
		\sa11_reg[7]/NET0131 ,
		_w12124_,
		_w12125_
	);
	LUT2 #(
		.INIT('h8)
	) name11594 (
		\sa11_reg[3]/P0001 ,
		_w11892_,
		_w12126_
	);
	LUT2 #(
		.INIT('h8)
	) name11595 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w12127_
	);
	LUT2 #(
		.INIT('h8)
	) name11596 (
		\sa11_reg[5]/P0001 ,
		_w12127_,
		_w12128_
	);
	LUT2 #(
		.INIT('h4)
	) name11597 (
		\sa11_reg[7]/NET0131 ,
		_w12128_,
		_w12129_
	);
	LUT2 #(
		.INIT('h1)
	) name11598 (
		_w12126_,
		_w12129_,
		_w12130_
	);
	LUT2 #(
		.INIT('h2)
	) name11599 (
		\sa11_reg[2]/P0001 ,
		_w12130_,
		_w12131_
	);
	LUT2 #(
		.INIT('h1)
	) name11600 (
		_w11935_,
		_w12119_,
		_w12132_
	);
	LUT2 #(
		.INIT('h1)
	) name11601 (
		_w12121_,
		_w12123_,
		_w12133_
	);
	LUT2 #(
		.INIT('h4)
	) name11602 (
		_w12125_,
		_w12133_,
		_w12134_
	);
	LUT2 #(
		.INIT('h8)
	) name11603 (
		_w12132_,
		_w12134_,
		_w12135_
	);
	LUT2 #(
		.INIT('h1)
	) name11604 (
		_w12118_,
		_w12131_,
		_w12136_
	);
	LUT2 #(
		.INIT('h8)
	) name11605 (
		_w12135_,
		_w12136_,
		_w12137_
	);
	LUT2 #(
		.INIT('h2)
	) name11606 (
		\sa11_reg[1]/P0001 ,
		_w12137_,
		_w12138_
	);
	LUT2 #(
		.INIT('h8)
	) name11607 (
		_w11801_,
		_w11853_,
		_w12139_
	);
	LUT2 #(
		.INIT('h1)
	) name11608 (
		_w11814_,
		_w12139_,
		_w12140_
	);
	LUT2 #(
		.INIT('h1)
	) name11609 (
		\sa11_reg[2]/P0001 ,
		_w12140_,
		_w12141_
	);
	LUT2 #(
		.INIT('h8)
	) name11610 (
		_w11876_,
		_w11877_,
		_w12142_
	);
	LUT2 #(
		.INIT('h1)
	) name11611 (
		_w12124_,
		_w12142_,
		_w12143_
	);
	LUT2 #(
		.INIT('h2)
	) name11612 (
		\sa11_reg[7]/NET0131 ,
		_w12143_,
		_w12144_
	);
	LUT2 #(
		.INIT('h2)
	) name11613 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[5]/P0001 ,
		_w12145_
	);
	LUT2 #(
		.INIT('h4)
	) name11614 (
		\sa11_reg[3]/P0001 ,
		_w11829_,
		_w12146_
	);
	LUT2 #(
		.INIT('h1)
	) name11615 (
		_w11880_,
		_w12146_,
		_w12147_
	);
	LUT2 #(
		.INIT('h2)
	) name11616 (
		_w12145_,
		_w12147_,
		_w12148_
	);
	LUT2 #(
		.INIT('h1)
	) name11617 (
		_w12144_,
		_w12148_,
		_w12149_
	);
	LUT2 #(
		.INIT('h1)
	) name11618 (
		\sa11_reg[1]/P0001 ,
		_w12149_,
		_w12150_
	);
	LUT2 #(
		.INIT('h8)
	) name11619 (
		_w11800_,
		_w11812_,
		_w12151_
	);
	LUT2 #(
		.INIT('h8)
	) name11620 (
		\sa11_reg[4]/P0001 ,
		_w11892_,
		_w12152_
	);
	LUT2 #(
		.INIT('h4)
	) name11621 (
		\sa11_reg[4]/P0001 ,
		_w11812_,
		_w12153_
	);
	LUT2 #(
		.INIT('h1)
	) name11622 (
		_w12152_,
		_w12153_,
		_w12154_
	);
	LUT2 #(
		.INIT('h2)
	) name11623 (
		\sa11_reg[3]/P0001 ,
		_w12154_,
		_w12155_
	);
	LUT2 #(
		.INIT('h1)
	) name11624 (
		_w11800_,
		_w11936_,
		_w12156_
	);
	LUT2 #(
		.INIT('h1)
	) name11625 (
		\sa11_reg[7]/NET0131 ,
		_w12156_,
		_w12157_
	);
	LUT2 #(
		.INIT('h1)
	) name11626 (
		_w12155_,
		_w12157_,
		_w12158_
	);
	LUT2 #(
		.INIT('h2)
	) name11627 (
		\sa11_reg[2]/P0001 ,
		_w12158_,
		_w12159_
	);
	LUT2 #(
		.INIT('h8)
	) name11628 (
		_w11798_,
		_w11823_,
		_w12160_
	);
	LUT2 #(
		.INIT('h1)
	) name11629 (
		_w12151_,
		_w12160_,
		_w12161_
	);
	LUT2 #(
		.INIT('h4)
	) name11630 (
		_w12141_,
		_w12161_,
		_w12162_
	);
	LUT2 #(
		.INIT('h4)
	) name11631 (
		_w12150_,
		_w12162_,
		_w12163_
	);
	LUT2 #(
		.INIT('h4)
	) name11632 (
		_w12159_,
		_w12163_,
		_w12164_
	);
	LUT2 #(
		.INIT('h4)
	) name11633 (
		_w12138_,
		_w12164_,
		_w12165_
	);
	LUT2 #(
		.INIT('h1)
	) name11634 (
		\sa11_reg[0]/P0001 ,
		_w12165_,
		_w12166_
	);
	LUT2 #(
		.INIT('h1)
	) name11635 (
		_w11915_,
		_w11925_,
		_w12167_
	);
	LUT2 #(
		.INIT('h4)
	) name11636 (
		\sa11_reg[4]/P0001 ,
		_w11825_,
		_w12168_
	);
	LUT2 #(
		.INIT('h4)
	) name11637 (
		\sa11_reg[4]/P0001 ,
		_w11876_,
		_w12169_
	);
	LUT2 #(
		.INIT('h1)
	) name11638 (
		_w11813_,
		_w11923_,
		_w12170_
	);
	LUT2 #(
		.INIT('h4)
	) name11639 (
		_w12169_,
		_w12170_,
		_w12171_
	);
	LUT2 #(
		.INIT('h2)
	) name11640 (
		\sa11_reg[1]/P0001 ,
		_w12171_,
		_w12172_
	);
	LUT2 #(
		.INIT('h2)
	) name11641 (
		_w12167_,
		_w12168_,
		_w12173_
	);
	LUT2 #(
		.INIT('h4)
	) name11642 (
		_w12172_,
		_w12173_,
		_w12174_
	);
	LUT2 #(
		.INIT('h1)
	) name11643 (
		\sa11_reg[2]/P0001 ,
		_w12174_,
		_w12175_
	);
	LUT2 #(
		.INIT('h8)
	) name11644 (
		_w11798_,
		_w11877_,
		_w12176_
	);
	LUT2 #(
		.INIT('h8)
	) name11645 (
		_w11794_,
		_w11847_,
		_w12177_
	);
	LUT2 #(
		.INIT('h1)
	) name11646 (
		_w12176_,
		_w12177_,
		_w12178_
	);
	LUT2 #(
		.INIT('h8)
	) name11647 (
		_w11796_,
		_w11870_,
		_w12179_
	);
	LUT2 #(
		.INIT('h1)
	) name11648 (
		_w11879_,
		_w12179_,
		_w12180_
	);
	LUT2 #(
		.INIT('h8)
	) name11649 (
		_w12178_,
		_w12180_,
		_w12181_
	);
	LUT2 #(
		.INIT('h2)
	) name11650 (
		\sa11_reg[1]/P0001 ,
		_w12181_,
		_w12182_
	);
	LUT2 #(
		.INIT('h1)
	) name11651 (
		_w11817_,
		_w11901_,
		_w12183_
	);
	LUT2 #(
		.INIT('h2)
	) name11652 (
		\sa11_reg[2]/P0001 ,
		_w12183_,
		_w12184_
	);
	LUT2 #(
		.INIT('h8)
	) name11653 (
		_w11892_,
		_w12127_,
		_w12185_
	);
	LUT2 #(
		.INIT('h4)
	) name11654 (
		\sa11_reg[3]/P0001 ,
		_w12185_,
		_w12186_
	);
	LUT2 #(
		.INIT('h2)
	) name11655 (
		_w11792_,
		_w11805_,
		_w12187_
	);
	LUT2 #(
		.INIT('h4)
	) name11656 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w12188_
	);
	LUT2 #(
		.INIT('h8)
	) name11657 (
		_w11871_,
		_w12188_,
		_w12189_
	);
	LUT2 #(
		.INIT('h1)
	) name11658 (
		_w12186_,
		_w12187_,
		_w12190_
	);
	LUT2 #(
		.INIT('h4)
	) name11659 (
		_w12189_,
		_w12190_,
		_w12191_
	);
	LUT2 #(
		.INIT('h4)
	) name11660 (
		_w12184_,
		_w12191_,
		_w12192_
	);
	LUT2 #(
		.INIT('h1)
	) name11661 (
		\sa11_reg[1]/P0001 ,
		_w12192_,
		_w12193_
	);
	LUT2 #(
		.INIT('h4)
	) name11662 (
		\sa11_reg[5]/P0001 ,
		_w11791_,
		_w12194_
	);
	LUT2 #(
		.INIT('h8)
	) name11663 (
		_w11860_,
		_w12194_,
		_w12195_
	);
	LUT2 #(
		.INIT('h1)
	) name11664 (
		_w12186_,
		_w12195_,
		_w12196_
	);
	LUT2 #(
		.INIT('h2)
	) name11665 (
		\sa11_reg[2]/P0001 ,
		_w12196_,
		_w12197_
	);
	LUT2 #(
		.INIT('h8)
	) name11666 (
		_w11792_,
		_w11796_,
		_w12198_
	);
	LUT2 #(
		.INIT('h1)
	) name11667 (
		_w11824_,
		_w12198_,
		_w12199_
	);
	LUT2 #(
		.INIT('h4)
	) name11668 (
		_w12197_,
		_w12199_,
		_w12200_
	);
	LUT2 #(
		.INIT('h4)
	) name11669 (
		_w12182_,
		_w12200_,
		_w12201_
	);
	LUT2 #(
		.INIT('h4)
	) name11670 (
		_w12175_,
		_w12201_,
		_w12202_
	);
	LUT2 #(
		.INIT('h4)
	) name11671 (
		_w12193_,
		_w12202_,
		_w12203_
	);
	LUT2 #(
		.INIT('h2)
	) name11672 (
		\sa11_reg[0]/P0001 ,
		_w12203_,
		_w12204_
	);
	LUT2 #(
		.INIT('h8)
	) name11673 (
		\sa11_reg[4]/P0001 ,
		_w11848_,
		_w12205_
	);
	LUT2 #(
		.INIT('h8)
	) name11674 (
		\sa11_reg[2]/P0001 ,
		_w11877_,
		_w12206_
	);
	LUT2 #(
		.INIT('h1)
	) name11675 (
		_w11871_,
		_w12194_,
		_w12207_
	);
	LUT2 #(
		.INIT('h4)
	) name11676 (
		_w11933_,
		_w12207_,
		_w12208_
	);
	LUT2 #(
		.INIT('h2)
	) name11677 (
		_w12206_,
		_w12208_,
		_w12209_
	);
	LUT2 #(
		.INIT('h8)
	) name11678 (
		\sa11_reg[5]/P0001 ,
		_w11794_,
		_w12210_
	);
	LUT2 #(
		.INIT('h8)
	) name11679 (
		_w11831_,
		_w12210_,
		_w12211_
	);
	LUT2 #(
		.INIT('h1)
	) name11680 (
		_w11865_,
		_w12211_,
		_w12212_
	);
	LUT2 #(
		.INIT('h4)
	) name11681 (
		_w12209_,
		_w12212_,
		_w12213_
	);
	LUT2 #(
		.INIT('h1)
	) name11682 (
		\sa11_reg[1]/P0001 ,
		_w12213_,
		_w12214_
	);
	LUT2 #(
		.INIT('h1)
	) name11683 (
		_w11881_,
		_w11935_,
		_w12215_
	);
	LUT2 #(
		.INIT('h1)
	) name11684 (
		\sa11_reg[2]/P0001 ,
		_w12215_,
		_w12216_
	);
	LUT2 #(
		.INIT('h8)
	) name11685 (
		\sa11_reg[3]/P0001 ,
		_w12151_,
		_w12217_
	);
	LUT2 #(
		.INIT('h8)
	) name11686 (
		_w11792_,
		_w12206_,
		_w12218_
	);
	LUT2 #(
		.INIT('h1)
	) name11687 (
		_w12160_,
		_w12217_,
		_w12219_
	);
	LUT2 #(
		.INIT('h4)
	) name11688 (
		_w12218_,
		_w12219_,
		_w12220_
	);
	LUT2 #(
		.INIT('h2)
	) name11689 (
		\sa11_reg[1]/P0001 ,
		_w12220_,
		_w12221_
	);
	LUT2 #(
		.INIT('h1)
	) name11690 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[2]/P0001 ,
		_w12222_
	);
	LUT2 #(
		.INIT('h8)
	) name11691 (
		_w11801_,
		_w12127_,
		_w12223_
	);
	LUT2 #(
		.INIT('h8)
	) name11692 (
		\sa11_reg[5]/P0001 ,
		_w11861_,
		_w12224_
	);
	LUT2 #(
		.INIT('h1)
	) name11693 (
		_w11941_,
		_w12223_,
		_w12225_
	);
	LUT2 #(
		.INIT('h4)
	) name11694 (
		_w12224_,
		_w12225_,
		_w12226_
	);
	LUT2 #(
		.INIT('h2)
	) name11695 (
		_w12222_,
		_w12226_,
		_w12227_
	);
	LUT2 #(
		.INIT('h1)
	) name11696 (
		_w12205_,
		_w12216_,
		_w12228_
	);
	LUT2 #(
		.INIT('h4)
	) name11697 (
		_w12221_,
		_w12228_,
		_w12229_
	);
	LUT2 #(
		.INIT('h4)
	) name11698 (
		_w12227_,
		_w12229_,
		_w12230_
	);
	LUT2 #(
		.INIT('h4)
	) name11699 (
		_w12214_,
		_w12230_,
		_w12231_
	);
	LUT2 #(
		.INIT('h4)
	) name11700 (
		_w12166_,
		_w12231_,
		_w12232_
	);
	LUT2 #(
		.INIT('h4)
	) name11701 (
		_w12204_,
		_w12232_,
		_w12233_
	);
	LUT2 #(
		.INIT('h1)
	) name11702 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w12234_
	);
	LUT2 #(
		.INIT('h8)
	) name11703 (
		\sa22_reg[3]/P0001 ,
		_w12234_,
		_w12235_
	);
	LUT2 #(
		.INIT('h4)
	) name11704 (
		\sa22_reg[7]/NET0131 ,
		_w12235_,
		_w12236_
	);
	LUT2 #(
		.INIT('h2)
	) name11705 (
		\sa22_reg[1]/P0001 ,
		_w12236_,
		_w12237_
	);
	LUT2 #(
		.INIT('h1)
	) name11706 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w12238_
	);
	LUT2 #(
		.INIT('h8)
	) name11707 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w12239_
	);
	LUT2 #(
		.INIT('h8)
	) name11708 (
		_w12238_,
		_w12239_,
		_w12240_
	);
	LUT2 #(
		.INIT('h4)
	) name11709 (
		\sa22_reg[7]/NET0131 ,
		_w12240_,
		_w12241_
	);
	LUT2 #(
		.INIT('h4)
	) name11710 (
		\sa22_reg[7]/NET0131 ,
		_w12238_,
		_w12242_
	);
	LUT2 #(
		.INIT('h8)
	) name11711 (
		\sa22_reg[6]/NET0131 ,
		_w12242_,
		_w12243_
	);
	LUT2 #(
		.INIT('h4)
	) name11712 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w12244_
	);
	LUT2 #(
		.INIT('h2)
	) name11713 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w12245_
	);
	LUT2 #(
		.INIT('h8)
	) name11714 (
		_w12244_,
		_w12245_,
		_w12246_
	);
	LUT2 #(
		.INIT('h1)
	) name11715 (
		\sa22_reg[2]/P0001 ,
		_w12246_,
		_w12247_
	);
	LUT2 #(
		.INIT('h4)
	) name11716 (
		_w12243_,
		_w12247_,
		_w12248_
	);
	LUT2 #(
		.INIT('h8)
	) name11717 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w12249_
	);
	LUT2 #(
		.INIT('h8)
	) name11718 (
		\sa22_reg[3]/P0001 ,
		_w12249_,
		_w12250_
	);
	LUT2 #(
		.INIT('h2)
	) name11719 (
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w12251_
	);
	LUT2 #(
		.INIT('h8)
	) name11720 (
		\sa22_reg[4]/P0001 ,
		_w12251_,
		_w12252_
	);
	LUT2 #(
		.INIT('h8)
	) name11721 (
		\sa22_reg[5]/P0001 ,
		_w12252_,
		_w12253_
	);
	LUT2 #(
		.INIT('h2)
	) name11722 (
		\sa22_reg[2]/P0001 ,
		_w12250_,
		_w12254_
	);
	LUT2 #(
		.INIT('h4)
	) name11723 (
		_w12253_,
		_w12254_,
		_w12255_
	);
	LUT2 #(
		.INIT('h1)
	) name11724 (
		_w12248_,
		_w12255_,
		_w12256_
	);
	LUT2 #(
		.INIT('h4)
	) name11725 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w12257_
	);
	LUT2 #(
		.INIT('h4)
	) name11726 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w12258_
	);
	LUT2 #(
		.INIT('h8)
	) name11727 (
		_w12257_,
		_w12258_,
		_w12259_
	);
	LUT2 #(
		.INIT('h8)
	) name11728 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w12260_
	);
	LUT2 #(
		.INIT('h8)
	) name11729 (
		\sa22_reg[5]/P0001 ,
		_w12260_,
		_w12261_
	);
	LUT2 #(
		.INIT('h8)
	) name11730 (
		\sa22_reg[7]/NET0131 ,
		_w12261_,
		_w12262_
	);
	LUT2 #(
		.INIT('h2)
	) name11731 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w12263_
	);
	LUT2 #(
		.INIT('h8)
	) name11732 (
		\sa22_reg[7]/NET0131 ,
		_w12263_,
		_w12264_
	);
	LUT2 #(
		.INIT('h4)
	) name11733 (
		\sa22_reg[2]/P0001 ,
		_w12264_,
		_w12265_
	);
	LUT2 #(
		.INIT('h4)
	) name11734 (
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w12266_
	);
	LUT2 #(
		.INIT('h4)
	) name11735 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		_w12267_
	);
	LUT2 #(
		.INIT('h8)
	) name11736 (
		_w12266_,
		_w12267_,
		_w12268_
	);
	LUT2 #(
		.INIT('h1)
	) name11737 (
		_w12259_,
		_w12268_,
		_w12269_
	);
	LUT2 #(
		.INIT('h4)
	) name11738 (
		_w12241_,
		_w12269_,
		_w12270_
	);
	LUT2 #(
		.INIT('h1)
	) name11739 (
		_w12262_,
		_w12265_,
		_w12271_
	);
	LUT2 #(
		.INIT('h8)
	) name11740 (
		_w12270_,
		_w12271_,
		_w12272_
	);
	LUT2 #(
		.INIT('h8)
	) name11741 (
		_w12237_,
		_w12272_,
		_w12273_
	);
	LUT2 #(
		.INIT('h4)
	) name11742 (
		_w12256_,
		_w12273_,
		_w12274_
	);
	LUT2 #(
		.INIT('h8)
	) name11743 (
		_w12234_,
		_w12258_,
		_w12275_
	);
	LUT2 #(
		.INIT('h8)
	) name11744 (
		\sa22_reg[4]/P0001 ,
		_w12275_,
		_w12276_
	);
	LUT2 #(
		.INIT('h1)
	) name11745 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w12277_
	);
	LUT2 #(
		.INIT('h2)
	) name11746 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w12278_
	);
	LUT2 #(
		.INIT('h8)
	) name11747 (
		_w12277_,
		_w12278_,
		_w12279_
	);
	LUT2 #(
		.INIT('h4)
	) name11748 (
		\sa22_reg[3]/P0001 ,
		_w12279_,
		_w12280_
	);
	LUT2 #(
		.INIT('h8)
	) name11749 (
		\sa22_reg[7]/NET0131 ,
		_w12240_,
		_w12281_
	);
	LUT2 #(
		.INIT('h2)
	) name11750 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w12282_
	);
	LUT2 #(
		.INIT('h8)
	) name11751 (
		_w12235_,
		_w12282_,
		_w12283_
	);
	LUT2 #(
		.INIT('h1)
	) name11752 (
		\sa22_reg[1]/P0001 ,
		_w12276_,
		_w12284_
	);
	LUT2 #(
		.INIT('h1)
	) name11753 (
		_w12280_,
		_w12281_,
		_w12285_
	);
	LUT2 #(
		.INIT('h4)
	) name11754 (
		_w12283_,
		_w12285_,
		_w12286_
	);
	LUT2 #(
		.INIT('h8)
	) name11755 (
		_w12284_,
		_w12286_,
		_w12287_
	);
	LUT2 #(
		.INIT('h1)
	) name11756 (
		_w12274_,
		_w12287_,
		_w12288_
	);
	LUT2 #(
		.INIT('h8)
	) name11757 (
		_w12260_,
		_w12277_,
		_w12289_
	);
	LUT2 #(
		.INIT('h4)
	) name11758 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w12290_
	);
	LUT2 #(
		.INIT('h4)
	) name11759 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w12291_
	);
	LUT2 #(
		.INIT('h8)
	) name11760 (
		_w12290_,
		_w12291_,
		_w12292_
	);
	LUT2 #(
		.INIT('h1)
	) name11761 (
		_w12289_,
		_w12292_,
		_w12293_
	);
	LUT2 #(
		.INIT('h1)
	) name11762 (
		\sa22_reg[2]/P0001 ,
		_w12293_,
		_w12294_
	);
	LUT2 #(
		.INIT('h4)
	) name11763 (
		\sa22_reg[4]/P0001 ,
		_w12234_,
		_w12295_
	);
	LUT2 #(
		.INIT('h4)
	) name11764 (
		\sa22_reg[7]/NET0131 ,
		_w12295_,
		_w12296_
	);
	LUT2 #(
		.INIT('h8)
	) name11765 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w12297_
	);
	LUT2 #(
		.INIT('h8)
	) name11766 (
		_w12245_,
		_w12297_,
		_w12298_
	);
	LUT2 #(
		.INIT('h4)
	) name11767 (
		\sa22_reg[2]/P0001 ,
		_w12298_,
		_w12299_
	);
	LUT2 #(
		.INIT('h1)
	) name11768 (
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w12300_
	);
	LUT2 #(
		.INIT('h4)
	) name11769 (
		\sa22_reg[4]/P0001 ,
		_w12300_,
		_w12301_
	);
	LUT2 #(
		.INIT('h8)
	) name11770 (
		\sa22_reg[6]/NET0131 ,
		_w12244_,
		_w12302_
	);
	LUT2 #(
		.INIT('h2)
	) name11771 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w12303_
	);
	LUT2 #(
		.INIT('h1)
	) name11772 (
		_w12302_,
		_w12303_,
		_w12304_
	);
	LUT2 #(
		.INIT('h2)
	) name11773 (
		_w12277_,
		_w12304_,
		_w12305_
	);
	LUT2 #(
		.INIT('h1)
	) name11774 (
		_w12262_,
		_w12301_,
		_w12306_
	);
	LUT2 #(
		.INIT('h4)
	) name11775 (
		_w12305_,
		_w12306_,
		_w12307_
	);
	LUT2 #(
		.INIT('h2)
	) name11776 (
		\sa22_reg[2]/P0001 ,
		_w12307_,
		_w12308_
	);
	LUT2 #(
		.INIT('h1)
	) name11777 (
		_w12296_,
		_w12299_,
		_w12309_
	);
	LUT2 #(
		.INIT('h4)
	) name11778 (
		_w12294_,
		_w12309_,
		_w12310_
	);
	LUT2 #(
		.INIT('h4)
	) name11779 (
		_w12308_,
		_w12310_,
		_w12311_
	);
	LUT2 #(
		.INIT('h4)
	) name11780 (
		_w12288_,
		_w12311_,
		_w12312_
	);
	LUT2 #(
		.INIT('h1)
	) name11781 (
		\sa22_reg[0]/P0001 ,
		_w12312_,
		_w12313_
	);
	LUT2 #(
		.INIT('h4)
	) name11782 (
		\sa22_reg[4]/P0001 ,
		_w12257_,
		_w12314_
	);
	LUT2 #(
		.INIT('h4)
	) name11783 (
		\sa22_reg[6]/NET0131 ,
		_w12260_,
		_w12315_
	);
	LUT2 #(
		.INIT('h4)
	) name11784 (
		\sa22_reg[7]/NET0131 ,
		_w12315_,
		_w12316_
	);
	LUT2 #(
		.INIT('h1)
	) name11785 (
		_w12314_,
		_w12316_,
		_w12317_
	);
	LUT2 #(
		.INIT('h2)
	) name11786 (
		\sa22_reg[2]/P0001 ,
		_w12317_,
		_w12318_
	);
	LUT2 #(
		.INIT('h8)
	) name11787 (
		\sa22_reg[7]/NET0131 ,
		_w12239_,
		_w12319_
	);
	LUT2 #(
		.INIT('h8)
	) name11788 (
		_w12244_,
		_w12319_,
		_w12320_
	);
	LUT2 #(
		.INIT('h8)
	) name11789 (
		\sa22_reg[5]/P0001 ,
		_w12251_,
		_w12321_
	);
	LUT2 #(
		.INIT('h2)
	) name11790 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		_w12322_
	);
	LUT2 #(
		.INIT('h2)
	) name11791 (
		_w12321_,
		_w12322_,
		_w12323_
	);
	LUT2 #(
		.INIT('h8)
	) name11792 (
		_w12263_,
		_w12291_,
		_w12324_
	);
	LUT2 #(
		.INIT('h4)
	) name11793 (
		\sa22_reg[2]/P0001 ,
		_w12324_,
		_w12325_
	);
	LUT2 #(
		.INIT('h1)
	) name11794 (
		_w12320_,
		_w12323_,
		_w12326_
	);
	LUT2 #(
		.INIT('h4)
	) name11795 (
		_w12325_,
		_w12326_,
		_w12327_
	);
	LUT2 #(
		.INIT('h4)
	) name11796 (
		_w12318_,
		_w12327_,
		_w12328_
	);
	LUT2 #(
		.INIT('h1)
	) name11797 (
		\sa22_reg[1]/P0001 ,
		_w12328_,
		_w12329_
	);
	LUT2 #(
		.INIT('h4)
	) name11798 (
		\sa22_reg[3]/P0001 ,
		_w12245_,
		_w12330_
	);
	LUT2 #(
		.INIT('h8)
	) name11799 (
		_w12297_,
		_w12330_,
		_w12331_
	);
	LUT2 #(
		.INIT('h8)
	) name11800 (
		\sa22_reg[5]/P0001 ,
		_w12300_,
		_w12332_
	);
	LUT2 #(
		.INIT('h8)
	) name11801 (
		_w12260_,
		_w12332_,
		_w12333_
	);
	LUT2 #(
		.INIT('h4)
	) name11802 (
		\sa22_reg[7]/NET0131 ,
		_w12244_,
		_w12334_
	);
	LUT2 #(
		.INIT('h8)
	) name11803 (
		_w12234_,
		_w12334_,
		_w12335_
	);
	LUT2 #(
		.INIT('h4)
	) name11804 (
		\sa22_reg[4]/P0001 ,
		_w12263_,
		_w12336_
	);
	LUT2 #(
		.INIT('h8)
	) name11805 (
		\sa22_reg[7]/NET0131 ,
		_w12336_,
		_w12337_
	);
	LUT2 #(
		.INIT('h1)
	) name11806 (
		_w12331_,
		_w12333_,
		_w12338_
	);
	LUT2 #(
		.INIT('h1)
	) name11807 (
		_w12335_,
		_w12337_,
		_w12339_
	);
	LUT2 #(
		.INIT('h8)
	) name11808 (
		_w12338_,
		_w12339_,
		_w12340_
	);
	LUT2 #(
		.INIT('h2)
	) name11809 (
		\sa22_reg[1]/P0001 ,
		_w12340_,
		_w12341_
	);
	LUT2 #(
		.INIT('h8)
	) name11810 (
		\sa22_reg[2]/P0001 ,
		_w12320_,
		_w12342_
	);
	LUT2 #(
		.INIT('h8)
	) name11811 (
		_w12303_,
		_w12321_,
		_w12343_
	);
	LUT2 #(
		.INIT('h8)
	) name11812 (
		\sa22_reg[4]/P0001 ,
		_w12291_,
		_w12344_
	);
	LUT2 #(
		.INIT('h8)
	) name11813 (
		\sa22_reg[6]/NET0131 ,
		_w12344_,
		_w12345_
	);
	LUT2 #(
		.INIT('h4)
	) name11814 (
		\sa22_reg[2]/P0001 ,
		_w12345_,
		_w12346_
	);
	LUT2 #(
		.INIT('h8)
	) name11815 (
		_w12277_,
		_w12290_,
		_w12347_
	);
	LUT2 #(
		.INIT('h8)
	) name11816 (
		_w12322_,
		_w12347_,
		_w12348_
	);
	LUT2 #(
		.INIT('h2)
	) name11817 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w12349_
	);
	LUT2 #(
		.INIT('h8)
	) name11818 (
		\sa22_reg[3]/P0001 ,
		_w12349_,
		_w12350_
	);
	LUT2 #(
		.INIT('h8)
	) name11819 (
		\sa22_reg[6]/NET0131 ,
		_w12350_,
		_w12351_
	);
	LUT2 #(
		.INIT('h8)
	) name11820 (
		\sa22_reg[3]/P0001 ,
		_w12251_,
		_w12352_
	);
	LUT2 #(
		.INIT('h4)
	) name11821 (
		\sa22_reg[4]/P0001 ,
		_w12352_,
		_w12353_
	);
	LUT2 #(
		.INIT('h1)
	) name11822 (
		_w12351_,
		_w12353_,
		_w12354_
	);
	LUT2 #(
		.INIT('h8)
	) name11823 (
		\sa22_reg[5]/P0001 ,
		_w12303_,
		_w12355_
	);
	LUT2 #(
		.INIT('h1)
	) name11824 (
		\sa22_reg[5]/P0001 ,
		_w12290_,
		_w12356_
	);
	LUT2 #(
		.INIT('h4)
	) name11825 (
		_w12297_,
		_w12356_,
		_w12357_
	);
	LUT2 #(
		.INIT('h1)
	) name11826 (
		_w12355_,
		_w12357_,
		_w12358_
	);
	LUT2 #(
		.INIT('h2)
	) name11827 (
		\sa22_reg[1]/P0001 ,
		_w12358_,
		_w12359_
	);
	LUT2 #(
		.INIT('h4)
	) name11828 (
		\sa22_reg[4]/P0001 ,
		_w12349_,
		_w12360_
	);
	LUT2 #(
		.INIT('h2)
	) name11829 (
		_w12354_,
		_w12360_,
		_w12361_
	);
	LUT2 #(
		.INIT('h4)
	) name11830 (
		_w12359_,
		_w12361_,
		_w12362_
	);
	LUT2 #(
		.INIT('h1)
	) name11831 (
		\sa22_reg[2]/P0001 ,
		_w12362_,
		_w12363_
	);
	LUT2 #(
		.INIT('h1)
	) name11832 (
		_w12343_,
		_w12348_,
		_w12364_
	);
	LUT2 #(
		.INIT('h4)
	) name11833 (
		_w12342_,
		_w12364_,
		_w12365_
	);
	LUT2 #(
		.INIT('h4)
	) name11834 (
		_w12346_,
		_w12365_,
		_w12366_
	);
	LUT2 #(
		.INIT('h4)
	) name11835 (
		_w12341_,
		_w12366_,
		_w12367_
	);
	LUT2 #(
		.INIT('h4)
	) name11836 (
		_w12329_,
		_w12367_,
		_w12368_
	);
	LUT2 #(
		.INIT('h4)
	) name11837 (
		_w12363_,
		_w12368_,
		_w12369_
	);
	LUT2 #(
		.INIT('h2)
	) name11838 (
		\sa22_reg[0]/P0001 ,
		_w12369_,
		_w12370_
	);
	LUT2 #(
		.INIT('h4)
	) name11839 (
		\sa22_reg[6]/NET0131 ,
		_w12242_,
		_w12371_
	);
	LUT2 #(
		.INIT('h8)
	) name11840 (
		_w12261_,
		_w12278_,
		_w12372_
	);
	LUT2 #(
		.INIT('h1)
	) name11841 (
		_w12251_,
		_w12266_,
		_w12373_
	);
	LUT2 #(
		.INIT('h1)
	) name11842 (
		\sa22_reg[5]/P0001 ,
		_w12373_,
		_w12374_
	);
	LUT2 #(
		.INIT('h1)
	) name11843 (
		_w12319_,
		_w12374_,
		_w12375_
	);
	LUT2 #(
		.INIT('h8)
	) name11844 (
		\sa22_reg[2]/P0001 ,
		_w12244_,
		_w12376_
	);
	LUT2 #(
		.INIT('h4)
	) name11845 (
		_w12375_,
		_w12376_,
		_w12377_
	);
	LUT2 #(
		.INIT('h1)
	) name11846 (
		_w12371_,
		_w12372_,
		_w12378_
	);
	LUT2 #(
		.INIT('h4)
	) name11847 (
		_w12377_,
		_w12378_,
		_w12379_
	);
	LUT2 #(
		.INIT('h1)
	) name11848 (
		\sa22_reg[1]/P0001 ,
		_w12379_,
		_w12380_
	);
	LUT2 #(
		.INIT('h4)
	) name11849 (
		\sa22_reg[7]/NET0131 ,
		_w12261_,
		_w12381_
	);
	LUT2 #(
		.INIT('h8)
	) name11850 (
		_w12278_,
		_w12381_,
		_w12382_
	);
	LUT2 #(
		.INIT('h1)
	) name11851 (
		\sa22_reg[1]/P0001 ,
		\sa22_reg[2]/P0001 ,
		_w12383_
	);
	LUT2 #(
		.INIT('h8)
	) name11852 (
		_w12251_,
		_w12261_,
		_w12384_
	);
	LUT2 #(
		.INIT('h4)
	) name11853 (
		\sa22_reg[4]/P0001 ,
		_w12258_,
		_w12385_
	);
	LUT2 #(
		.INIT('h8)
	) name11854 (
		\sa22_reg[5]/P0001 ,
		_w12385_,
		_w12386_
	);
	LUT2 #(
		.INIT('h1)
	) name11855 (
		_w12345_,
		_w12384_,
		_w12387_
	);
	LUT2 #(
		.INIT('h4)
	) name11856 (
		_w12386_,
		_w12387_,
		_w12388_
	);
	LUT2 #(
		.INIT('h2)
	) name11857 (
		_w12383_,
		_w12388_,
		_w12389_
	);
	LUT2 #(
		.INIT('h8)
	) name11858 (
		_w12303_,
		_w12332_,
		_w12390_
	);
	LUT2 #(
		.INIT('h1)
	) name11859 (
		_w12259_,
		_w12390_,
		_w12391_
	);
	LUT2 #(
		.INIT('h1)
	) name11860 (
		\sa22_reg[2]/P0001 ,
		_w12391_,
		_w12392_
	);
	LUT2 #(
		.INIT('h8)
	) name11861 (
		_w12239_,
		_w12334_,
		_w12393_
	);
	LUT2 #(
		.INIT('h8)
	) name11862 (
		\sa22_reg[2]/P0001 ,
		_w12393_,
		_w12394_
	);
	LUT2 #(
		.INIT('h4)
	) name11863 (
		\sa22_reg[4]/P0001 ,
		_w12277_,
		_w12395_
	);
	LUT2 #(
		.INIT('h8)
	) name11864 (
		_w12263_,
		_w12395_,
		_w12396_
	);
	LUT2 #(
		.INIT('h1)
	) name11865 (
		_w12299_,
		_w12396_,
		_w12397_
	);
	LUT2 #(
		.INIT('h4)
	) name11866 (
		_w12394_,
		_w12397_,
		_w12398_
	);
	LUT2 #(
		.INIT('h2)
	) name11867 (
		\sa22_reg[1]/P0001 ,
		_w12398_,
		_w12399_
	);
	LUT2 #(
		.INIT('h1)
	) name11868 (
		_w12382_,
		_w12392_,
		_w12400_
	);
	LUT2 #(
		.INIT('h4)
	) name11869 (
		_w12389_,
		_w12400_,
		_w12401_
	);
	LUT2 #(
		.INIT('h4)
	) name11870 (
		_w12399_,
		_w12401_,
		_w12402_
	);
	LUT2 #(
		.INIT('h4)
	) name11871 (
		_w12380_,
		_w12402_,
		_w12403_
	);
	LUT2 #(
		.INIT('h4)
	) name11872 (
		_w12313_,
		_w12403_,
		_w12404_
	);
	LUT2 #(
		.INIT('h4)
	) name11873 (
		_w12370_,
		_w12404_,
		_w12405_
	);
	LUT2 #(
		.INIT('h2)
	) name11874 (
		_w12233_,
		_w12405_,
		_w12406_
	);
	LUT2 #(
		.INIT('h4)
	) name11875 (
		_w12233_,
		_w12405_,
		_w12407_
	);
	LUT2 #(
		.INIT('h1)
	) name11876 (
		_w12406_,
		_w12407_,
		_w12408_
	);
	LUT2 #(
		.INIT('h4)
	) name11877 (
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w12409_
	);
	LUT2 #(
		.INIT('h4)
	) name11878 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		_w12410_
	);
	LUT2 #(
		.INIT('h8)
	) name11879 (
		_w12409_,
		_w12410_,
		_w12411_
	);
	LUT2 #(
		.INIT('h8)
	) name11880 (
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w12412_
	);
	LUT2 #(
		.INIT('h4)
	) name11881 (
		\sa33_reg[5]/P0001 ,
		_w12412_,
		_w12413_
	);
	LUT2 #(
		.INIT('h2)
	) name11882 (
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w12414_
	);
	LUT2 #(
		.INIT('h8)
	) name11883 (
		_w12410_,
		_w12414_,
		_w12415_
	);
	LUT2 #(
		.INIT('h1)
	) name11884 (
		_w12413_,
		_w12415_,
		_w12416_
	);
	LUT2 #(
		.INIT('h1)
	) name11885 (
		\sa33_reg[3]/P0001 ,
		_w12416_,
		_w12417_
	);
	LUT2 #(
		.INIT('h8)
	) name11886 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w12418_
	);
	LUT2 #(
		.INIT('h8)
	) name11887 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w12419_
	);
	LUT2 #(
		.INIT('h8)
	) name11888 (
		_w12418_,
		_w12419_,
		_w12420_
	);
	LUT2 #(
		.INIT('h8)
	) name11889 (
		\sa33_reg[3]/P0001 ,
		_w12418_,
		_w12421_
	);
	LUT2 #(
		.INIT('h8)
	) name11890 (
		\sa33_reg[4]/P0001 ,
		_w12414_,
		_w12422_
	);
	LUT2 #(
		.INIT('h8)
	) name11891 (
		\sa33_reg[5]/P0001 ,
		_w12422_,
		_w12423_
	);
	LUT2 #(
		.INIT('h1)
	) name11892 (
		_w12421_,
		_w12423_,
		_w12424_
	);
	LUT2 #(
		.INIT('h2)
	) name11893 (
		\sa33_reg[2]/P0001 ,
		_w12424_,
		_w12425_
	);
	LUT2 #(
		.INIT('h2)
	) name11894 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		_w12426_
	);
	LUT2 #(
		.INIT('h4)
	) name11895 (
		\sa33_reg[6]/P0001 ,
		_w12426_,
		_w12427_
	);
	LUT2 #(
		.INIT('h4)
	) name11896 (
		\sa33_reg[7]/NET0131 ,
		_w12427_,
		_w12428_
	);
	LUT2 #(
		.INIT('h2)
	) name11897 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w12429_
	);
	LUT2 #(
		.INIT('h4)
	) name11898 (
		\sa33_reg[3]/P0001 ,
		_w12429_,
		_w12430_
	);
	LUT2 #(
		.INIT('h8)
	) name11899 (
		\sa33_reg[4]/P0001 ,
		_w12430_,
		_w12431_
	);
	LUT2 #(
		.INIT('h8)
	) name11900 (
		\sa33_reg[3]/P0001 ,
		_w12409_,
		_w12432_
	);
	LUT2 #(
		.INIT('h4)
	) name11901 (
		\sa33_reg[3]/P0001 ,
		_w12414_,
		_w12433_
	);
	LUT2 #(
		.INIT('h4)
	) name11902 (
		\sa33_reg[4]/P0001 ,
		_w12433_,
		_w12434_
	);
	LUT2 #(
		.INIT('h1)
	) name11903 (
		_w12431_,
		_w12432_,
		_w12435_
	);
	LUT2 #(
		.INIT('h4)
	) name11904 (
		_w12434_,
		_w12435_,
		_w12436_
	);
	LUT2 #(
		.INIT('h1)
	) name11905 (
		\sa33_reg[2]/P0001 ,
		_w12436_,
		_w12437_
	);
	LUT2 #(
		.INIT('h1)
	) name11906 (
		_w12411_,
		_w12420_,
		_w12438_
	);
	LUT2 #(
		.INIT('h4)
	) name11907 (
		_w12428_,
		_w12438_,
		_w12439_
	);
	LUT2 #(
		.INIT('h4)
	) name11908 (
		_w12417_,
		_w12439_,
		_w12440_
	);
	LUT2 #(
		.INIT('h4)
	) name11909 (
		_w12425_,
		_w12440_,
		_w12441_
	);
	LUT2 #(
		.INIT('h4)
	) name11910 (
		_w12437_,
		_w12441_,
		_w12442_
	);
	LUT2 #(
		.INIT('h2)
	) name11911 (
		\sa33_reg[1]/P0001 ,
		_w12442_,
		_w12443_
	);
	LUT2 #(
		.INIT('h1)
	) name11912 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w12444_
	);
	LUT2 #(
		.INIT('h4)
	) name11913 (
		\sa33_reg[6]/P0001 ,
		_w12444_,
		_w12445_
	);
	LUT2 #(
		.INIT('h1)
	) name11914 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		_w12446_
	);
	LUT2 #(
		.INIT('h8)
	) name11915 (
		\sa33_reg[3]/P0001 ,
		_w12446_,
		_w12447_
	);
	LUT2 #(
		.INIT('h4)
	) name11916 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w12448_
	);
	LUT2 #(
		.INIT('h8)
	) name11917 (
		\sa33_reg[6]/P0001 ,
		_w12448_,
		_w12449_
	);
	LUT2 #(
		.INIT('h4)
	) name11918 (
		\sa33_reg[5]/P0001 ,
		_w12449_,
		_w12450_
	);
	LUT2 #(
		.INIT('h1)
	) name11919 (
		_w12447_,
		_w12450_,
		_w12451_
	);
	LUT2 #(
		.INIT('h1)
	) name11920 (
		\sa33_reg[7]/NET0131 ,
		_w12451_,
		_w12452_
	);
	LUT2 #(
		.INIT('h1)
	) name11921 (
		_w12420_,
		_w12445_,
		_w12453_
	);
	LUT2 #(
		.INIT('h4)
	) name11922 (
		_w12452_,
		_w12453_,
		_w12454_
	);
	LUT2 #(
		.INIT('h2)
	) name11923 (
		\sa33_reg[2]/P0001 ,
		_w12454_,
		_w12455_
	);
	LUT2 #(
		.INIT('h4)
	) name11924 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		_w12456_
	);
	LUT2 #(
		.INIT('h2)
	) name11925 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		_w12457_
	);
	LUT2 #(
		.INIT('h4)
	) name11926 (
		\sa33_reg[7]/NET0131 ,
		_w12457_,
		_w12458_
	);
	LUT2 #(
		.INIT('h8)
	) name11927 (
		_w12456_,
		_w12458_,
		_w12459_
	);
	LUT2 #(
		.INIT('h4)
	) name11928 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w12460_
	);
	LUT2 #(
		.INIT('h4)
	) name11929 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w12461_
	);
	LUT2 #(
		.INIT('h8)
	) name11930 (
		_w12460_,
		_w12461_,
		_w12462_
	);
	LUT2 #(
		.INIT('h4)
	) name11931 (
		\sa33_reg[2]/P0001 ,
		_w12462_,
		_w12463_
	);
	LUT2 #(
		.INIT('h1)
	) name11932 (
		_w12459_,
		_w12463_,
		_w12464_
	);
	LUT2 #(
		.INIT('h1)
	) name11933 (
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w12465_
	);
	LUT2 #(
		.INIT('h8)
	) name11934 (
		_w12446_,
		_w12465_,
		_w12466_
	);
	LUT2 #(
		.INIT('h8)
	) name11935 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w12467_
	);
	LUT2 #(
		.INIT('h8)
	) name11936 (
		_w12429_,
		_w12467_,
		_w12468_
	);
	LUT2 #(
		.INIT('h4)
	) name11937 (
		\sa33_reg[2]/P0001 ,
		_w12468_,
		_w12469_
	);
	LUT2 #(
		.INIT('h4)
	) name11938 (
		\sa33_reg[3]/P0001 ,
		_w12409_,
		_w12470_
	);
	LUT2 #(
		.INIT('h8)
	) name11939 (
		_w12457_,
		_w12470_,
		_w12471_
	);
	LUT2 #(
		.INIT('h2)
	) name11940 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		_w12472_
	);
	LUT2 #(
		.INIT('h4)
	) name11941 (
		\sa33_reg[5]/P0001 ,
		_w12465_,
		_w12473_
	);
	LUT2 #(
		.INIT('h8)
	) name11942 (
		_w12472_,
		_w12473_,
		_w12474_
	);
	LUT2 #(
		.INIT('h1)
	) name11943 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w12475_
	);
	LUT2 #(
		.INIT('h2)
	) name11944 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w12476_
	);
	LUT2 #(
		.INIT('h8)
	) name11945 (
		\sa33_reg[2]/P0001 ,
		_w12476_,
		_w12477_
	);
	LUT2 #(
		.INIT('h8)
	) name11946 (
		_w12475_,
		_w12477_,
		_w12478_
	);
	LUT2 #(
		.INIT('h1)
	) name11947 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w12479_
	);
	LUT2 #(
		.INIT('h8)
	) name11948 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w12480_
	);
	LUT2 #(
		.INIT('h8)
	) name11949 (
		\sa33_reg[7]/NET0131 ,
		_w12480_,
		_w12481_
	);
	LUT2 #(
		.INIT('h8)
	) name11950 (
		_w12479_,
		_w12481_,
		_w12482_
	);
	LUT2 #(
		.INIT('h1)
	) name11951 (
		_w12471_,
		_w12474_,
		_w12483_
	);
	LUT2 #(
		.INIT('h1)
	) name11952 (
		_w12478_,
		_w12482_,
		_w12484_
	);
	LUT2 #(
		.INIT('h8)
	) name11953 (
		_w12483_,
		_w12484_,
		_w12485_
	);
	LUT2 #(
		.INIT('h1)
	) name11954 (
		\sa33_reg[1]/P0001 ,
		_w12485_,
		_w12486_
	);
	LUT2 #(
		.INIT('h1)
	) name11955 (
		_w12466_,
		_w12469_,
		_w12487_
	);
	LUT2 #(
		.INIT('h8)
	) name11956 (
		_w12464_,
		_w12487_,
		_w12488_
	);
	LUT2 #(
		.INIT('h4)
	) name11957 (
		_w12486_,
		_w12488_,
		_w12489_
	);
	LUT2 #(
		.INIT('h4)
	) name11958 (
		_w12455_,
		_w12489_,
		_w12490_
	);
	LUT2 #(
		.INIT('h4)
	) name11959 (
		_w12443_,
		_w12490_,
		_w12491_
	);
	LUT2 #(
		.INIT('h1)
	) name11960 (
		\sa33_reg[0]/P0001 ,
		_w12491_,
		_w12492_
	);
	LUT2 #(
		.INIT('h8)
	) name11961 (
		_w12409_,
		_w12426_,
		_w12493_
	);
	LUT2 #(
		.INIT('h4)
	) name11962 (
		\sa33_reg[2]/P0001 ,
		_w12493_,
		_w12494_
	);
	LUT2 #(
		.INIT('h8)
	) name11963 (
		_w12419_,
		_w12465_,
		_w12495_
	);
	LUT2 #(
		.INIT('h8)
	) name11964 (
		\sa33_reg[6]/P0001 ,
		_w12446_,
		_w12496_
	);
	LUT2 #(
		.INIT('h1)
	) name11965 (
		_w12495_,
		_w12496_,
		_w12497_
	);
	LUT2 #(
		.INIT('h2)
	) name11966 (
		\sa33_reg[2]/P0001 ,
		_w12497_,
		_w12498_
	);
	LUT2 #(
		.INIT('h8)
	) name11967 (
		\sa33_reg[5]/P0001 ,
		_w12414_,
		_w12499_
	);
	LUT2 #(
		.INIT('h4)
	) name11968 (
		_w12472_,
		_w12499_,
		_w12500_
	);
	LUT2 #(
		.INIT('h8)
	) name11969 (
		_w12418_,
		_w12449_,
		_w12501_
	);
	LUT2 #(
		.INIT('h1)
	) name11970 (
		_w12494_,
		_w12500_,
		_w12502_
	);
	LUT2 #(
		.INIT('h4)
	) name11971 (
		_w12501_,
		_w12502_,
		_w12503_
	);
	LUT2 #(
		.INIT('h4)
	) name11972 (
		_w12498_,
		_w12503_,
		_w12504_
	);
	LUT2 #(
		.INIT('h1)
	) name11973 (
		\sa33_reg[1]/P0001 ,
		_w12504_,
		_w12505_
	);
	LUT2 #(
		.INIT('h8)
	) name11974 (
		_w12418_,
		_w12448_,
		_w12506_
	);
	LUT2 #(
		.INIT('h4)
	) name11975 (
		\sa33_reg[6]/P0001 ,
		_w12506_,
		_w12507_
	);
	LUT2 #(
		.INIT('h8)
	) name11976 (
		_w12448_,
		_w12473_,
		_w12508_
	);
	LUT2 #(
		.INIT('h8)
	) name11977 (
		_w12409_,
		_w12476_,
		_w12509_
	);
	LUT2 #(
		.INIT('h2)
	) name11978 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w12510_
	);
	LUT2 #(
		.INIT('h8)
	) name11979 (
		_w12419_,
		_w12510_,
		_w12511_
	);
	LUT2 #(
		.INIT('h4)
	) name11980 (
		\sa33_reg[6]/P0001 ,
		_w12511_,
		_w12512_
	);
	LUT2 #(
		.INIT('h1)
	) name11981 (
		_w12507_,
		_w12509_,
		_w12513_
	);
	LUT2 #(
		.INIT('h1)
	) name11982 (
		_w12508_,
		_w12512_,
		_w12514_
	);
	LUT2 #(
		.INIT('h8)
	) name11983 (
		_w12513_,
		_w12514_,
		_w12515_
	);
	LUT2 #(
		.INIT('h2)
	) name11984 (
		\sa33_reg[1]/P0001 ,
		_w12515_,
		_w12516_
	);
	LUT2 #(
		.INIT('h4)
	) name11985 (
		\sa33_reg[5]/P0001 ,
		_w12414_,
		_w12517_
	);
	LUT2 #(
		.INIT('h8)
	) name11986 (
		_w12479_,
		_w12517_,
		_w12518_
	);
	LUT2 #(
		.INIT('h1)
	) name11987 (
		_w12501_,
		_w12518_,
		_w12519_
	);
	LUT2 #(
		.INIT('h2)
	) name11988 (
		\sa33_reg[2]/P0001 ,
		_w12519_,
		_w12520_
	);
	LUT2 #(
		.INIT('h4)
	) name11989 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w12521_
	);
	LUT2 #(
		.INIT('h8)
	) name11990 (
		_w12467_,
		_w12521_,
		_w12522_
	);
	LUT2 #(
		.INIT('h4)
	) name11991 (
		\sa33_reg[2]/P0001 ,
		_w12522_,
		_w12523_
	);
	LUT2 #(
		.INIT('h8)
	) name11992 (
		_w12476_,
		_w12499_,
		_w12524_
	);
	LUT2 #(
		.INIT('h4)
	) name11993 (
		\sa33_reg[4]/P0001 ,
		_w12510_,
		_w12525_
	);
	LUT2 #(
		.INIT('h8)
	) name11994 (
		\sa33_reg[5]/P0001 ,
		_w12476_,
		_w12526_
	);
	LUT2 #(
		.INIT('h1)
	) name11995 (
		_w12460_,
		_w12467_,
		_w12527_
	);
	LUT2 #(
		.INIT('h4)
	) name11996 (
		\sa33_reg[5]/P0001 ,
		_w12527_,
		_w12528_
	);
	LUT2 #(
		.INIT('h1)
	) name11997 (
		_w12526_,
		_w12528_,
		_w12529_
	);
	LUT2 #(
		.INIT('h2)
	) name11998 (
		\sa33_reg[1]/P0001 ,
		_w12529_,
		_w12530_
	);
	LUT2 #(
		.INIT('h8)
	) name11999 (
		\sa33_reg[3]/P0001 ,
		_w12414_,
		_w12531_
	);
	LUT2 #(
		.INIT('h4)
	) name12000 (
		_w12457_,
		_w12531_,
		_w12532_
	);
	LUT2 #(
		.INIT('h1)
	) name12001 (
		_w12525_,
		_w12532_,
		_w12533_
	);
	LUT2 #(
		.INIT('h4)
	) name12002 (
		_w12530_,
		_w12533_,
		_w12534_
	);
	LUT2 #(
		.INIT('h1)
	) name12003 (
		\sa33_reg[2]/P0001 ,
		_w12534_,
		_w12535_
	);
	LUT2 #(
		.INIT('h1)
	) name12004 (
		_w12523_,
		_w12524_,
		_w12536_
	);
	LUT2 #(
		.INIT('h4)
	) name12005 (
		_w12520_,
		_w12536_,
		_w12537_
	);
	LUT2 #(
		.INIT('h4)
	) name12006 (
		_w12516_,
		_w12537_,
		_w12538_
	);
	LUT2 #(
		.INIT('h4)
	) name12007 (
		_w12505_,
		_w12538_,
		_w12539_
	);
	LUT2 #(
		.INIT('h4)
	) name12008 (
		_w12535_,
		_w12539_,
		_w12540_
	);
	LUT2 #(
		.INIT('h2)
	) name12009 (
		\sa33_reg[0]/P0001 ,
		_w12540_,
		_w12541_
	);
	LUT2 #(
		.INIT('h8)
	) name12010 (
		\sa33_reg[2]/P0001 ,
		_w12419_,
		_w12542_
	);
	LUT2 #(
		.INIT('h8)
	) name12011 (
		_w12429_,
		_w12542_,
		_w12543_
	);
	LUT2 #(
		.INIT('h4)
	) name12012 (
		\sa33_reg[5]/P0001 ,
		_w12409_,
		_w12544_
	);
	LUT2 #(
		.INIT('h1)
	) name12013 (
		_w12517_,
		_w12544_,
		_w12545_
	);
	LUT2 #(
		.INIT('h4)
	) name12014 (
		_w12481_,
		_w12545_,
		_w12546_
	);
	LUT2 #(
		.INIT('h8)
	) name12015 (
		\sa33_reg[4]/P0001 ,
		_w12472_,
		_w12547_
	);
	LUT2 #(
		.INIT('h4)
	) name12016 (
		_w12546_,
		_w12547_,
		_w12548_
	);
	LUT2 #(
		.INIT('h8)
	) name12017 (
		_w12465_,
		_w12479_,
		_w12549_
	);
	LUT2 #(
		.INIT('h8)
	) name12018 (
		\sa33_reg[6]/P0001 ,
		_w12511_,
		_w12550_
	);
	LUT2 #(
		.INIT('h8)
	) name12019 (
		\sa33_reg[7]/NET0131 ,
		_w12479_,
		_w12551_
	);
	LUT2 #(
		.INIT('h8)
	) name12020 (
		\sa33_reg[5]/P0001 ,
		_w12551_,
		_w12552_
	);
	LUT2 #(
		.INIT('h1)
	) name12021 (
		_w12522_,
		_w12550_,
		_w12553_
	);
	LUT2 #(
		.INIT('h4)
	) name12022 (
		_w12552_,
		_w12553_,
		_w12554_
	);
	LUT2 #(
		.INIT('h1)
	) name12023 (
		\sa33_reg[2]/P0001 ,
		_w12554_,
		_w12555_
	);
	LUT2 #(
		.INIT('h1)
	) name12024 (
		_w12543_,
		_w12549_,
		_w12556_
	);
	LUT2 #(
		.INIT('h4)
	) name12025 (
		_w12548_,
		_w12556_,
		_w12557_
	);
	LUT2 #(
		.INIT('h4)
	) name12026 (
		_w12555_,
		_w12557_,
		_w12558_
	);
	LUT2 #(
		.INIT('h1)
	) name12027 (
		\sa33_reg[1]/P0001 ,
		_w12558_,
		_w12559_
	);
	LUT2 #(
		.INIT('h8)
	) name12028 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		_w12560_
	);
	LUT2 #(
		.INIT('h8)
	) name12029 (
		\sa33_reg[5]/P0001 ,
		_w12465_,
		_w12561_
	);
	LUT2 #(
		.INIT('h8)
	) name12030 (
		_w12560_,
		_w12561_,
		_w12562_
	);
	LUT2 #(
		.INIT('h8)
	) name12031 (
		\sa33_reg[4]/P0001 ,
		_w12562_,
		_w12563_
	);
	LUT2 #(
		.INIT('h4)
	) name12032 (
		\sa33_reg[3]/P0001 ,
		_w12413_,
		_w12564_
	);
	LUT2 #(
		.INIT('h8)
	) name12033 (
		_w12429_,
		_w12476_,
		_w12565_
	);
	LUT2 #(
		.INIT('h4)
	) name12034 (
		\sa33_reg[7]/NET0131 ,
		_w12565_,
		_w12566_
	);
	LUT2 #(
		.INIT('h1)
	) name12035 (
		_w12564_,
		_w12566_,
		_w12567_
	);
	LUT2 #(
		.INIT('h1)
	) name12036 (
		\sa33_reg[2]/P0001 ,
		_w12567_,
		_w12568_
	);
	LUT2 #(
		.INIT('h8)
	) name12037 (
		_w12448_,
		_w12510_,
		_w12569_
	);
	LUT2 #(
		.INIT('h8)
	) name12038 (
		\sa33_reg[6]/P0001 ,
		_w12569_,
		_w12570_
	);
	LUT2 #(
		.INIT('h8)
	) name12039 (
		\sa33_reg[2]/P0001 ,
		_w12570_,
		_w12571_
	);
	LUT2 #(
		.INIT('h8)
	) name12040 (
		_w12427_,
		_w12444_,
		_w12572_
	);
	LUT2 #(
		.INIT('h1)
	) name12041 (
		_w12469_,
		_w12572_,
		_w12573_
	);
	LUT2 #(
		.INIT('h4)
	) name12042 (
		_w12571_,
		_w12573_,
		_w12574_
	);
	LUT2 #(
		.INIT('h2)
	) name12043 (
		\sa33_reg[1]/P0001 ,
		_w12574_,
		_w12575_
	);
	LUT2 #(
		.INIT('h1)
	) name12044 (
		_w12563_,
		_w12568_,
		_w12576_
	);
	LUT2 #(
		.INIT('h4)
	) name12045 (
		_w12575_,
		_w12576_,
		_w12577_
	);
	LUT2 #(
		.INIT('h4)
	) name12046 (
		_w12559_,
		_w12577_,
		_w12578_
	);
	LUT2 #(
		.INIT('h4)
	) name12047 (
		_w12492_,
		_w12578_,
		_w12579_
	);
	LUT2 #(
		.INIT('h4)
	) name12048 (
		_w12541_,
		_w12579_,
		_w12580_
	);
	LUT2 #(
		.INIT('h2)
	) name12049 (
		\u0_w_reg[0][29]/P0001 ,
		_w12580_,
		_w12581_
	);
	LUT2 #(
		.INIT('h4)
	) name12050 (
		\u0_w_reg[0][29]/P0001 ,
		_w12580_,
		_w12582_
	);
	LUT2 #(
		.INIT('h1)
	) name12051 (
		_w12581_,
		_w12582_,
		_w12583_
	);
	LUT2 #(
		.INIT('h8)
	) name12052 (
		_w12408_,
		_w12583_,
		_w12584_
	);
	LUT2 #(
		.INIT('h1)
	) name12053 (
		_w12408_,
		_w12583_,
		_w12585_
	);
	LUT2 #(
		.INIT('h1)
	) name12054 (
		_w12584_,
		_w12585_,
		_w12586_
	);
	LUT2 #(
		.INIT('h1)
	) name12055 (
		_w12114_,
		_w12586_,
		_w12587_
	);
	LUT2 #(
		.INIT('h8)
	) name12056 (
		_w12114_,
		_w12586_,
		_w12588_
	);
	LUT2 #(
		.INIT('h1)
	) name12057 (
		\ld_r_reg/P0001 ,
		_w12587_,
		_w12589_
	);
	LUT2 #(
		.INIT('h4)
	) name12058 (
		_w12588_,
		_w12589_,
		_w12590_
	);
	LUT2 #(
		.INIT('h1)
	) name12059 (
		\text_in_r_reg[125]/P0001 ,
		\u0_w_reg[0][29]/P0001 ,
		_w12591_
	);
	LUT2 #(
		.INIT('h8)
	) name12060 (
		\text_in_r_reg[125]/P0001 ,
		\u0_w_reg[0][29]/P0001 ,
		_w12592_
	);
	LUT2 #(
		.INIT('h2)
	) name12061 (
		\ld_r_reg/P0001 ,
		_w12591_,
		_w12593_
	);
	LUT2 #(
		.INIT('h4)
	) name12062 (
		_w12592_,
		_w12593_,
		_w12594_
	);
	LUT2 #(
		.INIT('h1)
	) name12063 (
		_w12590_,
		_w12594_,
		_w12595_
	);
	LUT2 #(
		.INIT('h8)
	) name12064 (
		\sa00_reg[2]/P0001 ,
		_w11966_,
		_w12596_
	);
	LUT2 #(
		.INIT('h4)
	) name12065 (
		\sa00_reg[7]/NET0131 ,
		_w12056_,
		_w12597_
	);
	LUT2 #(
		.INIT('h1)
	) name12066 (
		_w12596_,
		_w12597_,
		_w12598_
	);
	LUT2 #(
		.INIT('h1)
	) name12067 (
		\sa00_reg[6]/NET0131 ,
		_w12598_,
		_w12599_
	);
	LUT2 #(
		.INIT('h8)
	) name12068 (
		_w11952_,
		_w11955_,
		_w12600_
	);
	LUT2 #(
		.INIT('h1)
	) name12069 (
		_w12599_,
		_w12600_,
		_w12601_
	);
	LUT2 #(
		.INIT('h1)
	) name12070 (
		\sa00_reg[5]/P0001 ,
		_w12601_,
		_w12602_
	);
	LUT2 #(
		.INIT('h1)
	) name12071 (
		_w12046_,
		_w12602_,
		_w12603_
	);
	LUT2 #(
		.INIT('h1)
	) name12072 (
		\sa00_reg[1]/P0001 ,
		_w12603_,
		_w12604_
	);
	LUT2 #(
		.INIT('h8)
	) name12073 (
		\sa00_reg[5]/P0001 ,
		_w12057_,
		_w12605_
	);
	LUT2 #(
		.INIT('h1)
	) name12074 (
		_w11974_,
		_w12605_,
		_w12606_
	);
	LUT2 #(
		.INIT('h2)
	) name12075 (
		\sa00_reg[2]/P0001 ,
		_w12606_,
		_w12607_
	);
	LUT2 #(
		.INIT('h8)
	) name12076 (
		_w11962_,
		_w12005_,
		_w12608_
	);
	LUT2 #(
		.INIT('h1)
	) name12077 (
		_w12050_,
		_w12608_,
		_w12609_
	);
	LUT2 #(
		.INIT('h2)
	) name12078 (
		\sa00_reg[5]/P0001 ,
		_w12609_,
		_w12610_
	);
	LUT2 #(
		.INIT('h8)
	) name12079 (
		_w11956_,
		_w11992_,
		_w12611_
	);
	LUT2 #(
		.INIT('h8)
	) name12080 (
		_w11952_,
		_w12014_,
		_w12612_
	);
	LUT2 #(
		.INIT('h8)
	) name12081 (
		\sa00_reg[3]/P0001 ,
		_w11952_,
		_w12613_
	);
	LUT2 #(
		.INIT('h8)
	) name12082 (
		_w11955_,
		_w11975_,
		_w12614_
	);
	LUT2 #(
		.INIT('h1)
	) name12083 (
		_w12608_,
		_w12613_,
		_w12615_
	);
	LUT2 #(
		.INIT('h4)
	) name12084 (
		_w12614_,
		_w12615_,
		_w12616_
	);
	LUT2 #(
		.INIT('h1)
	) name12085 (
		\sa00_reg[2]/P0001 ,
		_w12616_,
		_w12617_
	);
	LUT2 #(
		.INIT('h1)
	) name12086 (
		_w12033_,
		_w12611_,
		_w12618_
	);
	LUT2 #(
		.INIT('h4)
	) name12087 (
		_w12612_,
		_w12618_,
		_w12619_
	);
	LUT2 #(
		.INIT('h4)
	) name12088 (
		_w12610_,
		_w12619_,
		_w12620_
	);
	LUT2 #(
		.INIT('h4)
	) name12089 (
		_w12607_,
		_w12620_,
		_w12621_
	);
	LUT2 #(
		.INIT('h4)
	) name12090 (
		_w12617_,
		_w12621_,
		_w12622_
	);
	LUT2 #(
		.INIT('h2)
	) name12091 (
		\sa00_reg[1]/P0001 ,
		_w12622_,
		_w12623_
	);
	LUT2 #(
		.INIT('h8)
	) name12092 (
		_w11978_,
		_w12035_,
		_w12624_
	);
	LUT2 #(
		.INIT('h8)
	) name12093 (
		\sa00_reg[4]/P0001 ,
		_w12064_,
		_w12625_
	);
	LUT2 #(
		.INIT('h8)
	) name12094 (
		\sa00_reg[3]/P0001 ,
		_w12625_,
		_w12626_
	);
	LUT2 #(
		.INIT('h1)
	) name12095 (
		_w12624_,
		_w12626_,
		_w12627_
	);
	LUT2 #(
		.INIT('h1)
	) name12096 (
		\sa00_reg[2]/P0001 ,
		_w12627_,
		_w12628_
	);
	LUT2 #(
		.INIT('h4)
	) name12097 (
		\sa00_reg[4]/P0001 ,
		_w11960_,
		_w12629_
	);
	LUT2 #(
		.INIT('h4)
	) name12098 (
		\sa00_reg[7]/NET0131 ,
		_w12629_,
		_w12630_
	);
	LUT2 #(
		.INIT('h8)
	) name12099 (
		_w12086_,
		_w12088_,
		_w12631_
	);
	LUT2 #(
		.INIT('h8)
	) name12100 (
		\sa00_reg[4]/P0001 ,
		_w11973_,
		_w12632_
	);
	LUT2 #(
		.INIT('h4)
	) name12101 (
		\sa00_reg[4]/P0001 ,
		_w12064_,
		_w12633_
	);
	LUT2 #(
		.INIT('h1)
	) name12102 (
		_w12632_,
		_w12633_,
		_w12634_
	);
	LUT2 #(
		.INIT('h2)
	) name12103 (
		\sa00_reg[3]/P0001 ,
		_w12634_,
		_w12635_
	);
	LUT2 #(
		.INIT('h4)
	) name12104 (
		\sa00_reg[4]/P0001 ,
		_w11956_,
		_w12636_
	);
	LUT2 #(
		.INIT('h4)
	) name12105 (
		\sa00_reg[7]/NET0131 ,
		_w12036_,
		_w12637_
	);
	LUT2 #(
		.INIT('h1)
	) name12106 (
		_w12636_,
		_w12637_,
		_w12638_
	);
	LUT2 #(
		.INIT('h4)
	) name12107 (
		_w12635_,
		_w12638_,
		_w12639_
	);
	LUT2 #(
		.INIT('h2)
	) name12108 (
		\sa00_reg[2]/P0001 ,
		_w12639_,
		_w12640_
	);
	LUT2 #(
		.INIT('h1)
	) name12109 (
		_w12630_,
		_w12631_,
		_w12641_
	);
	LUT2 #(
		.INIT('h4)
	) name12110 (
		_w12628_,
		_w12641_,
		_w12642_
	);
	LUT2 #(
		.INIT('h4)
	) name12111 (
		_w12640_,
		_w12642_,
		_w12643_
	);
	LUT2 #(
		.INIT('h4)
	) name12112 (
		_w12604_,
		_w12643_,
		_w12644_
	);
	LUT2 #(
		.INIT('h4)
	) name12113 (
		_w12623_,
		_w12644_,
		_w12645_
	);
	LUT2 #(
		.INIT('h1)
	) name12114 (
		\sa00_reg[0]/P0001 ,
		_w12645_,
		_w12646_
	);
	LUT2 #(
		.INIT('h8)
	) name12115 (
		_w11955_,
		_w11996_,
		_w12647_
	);
	LUT2 #(
		.INIT('h4)
	) name12116 (
		\sa00_reg[5]/P0001 ,
		_w12608_,
		_w12648_
	);
	LUT2 #(
		.INIT('h1)
	) name12117 (
		_w12647_,
		_w12648_,
		_w12649_
	);
	LUT2 #(
		.INIT('h2)
	) name12118 (
		\sa00_reg[2]/P0001 ,
		_w12649_,
		_w12650_
	);
	LUT2 #(
		.INIT('h8)
	) name12119 (
		\sa00_reg[5]/P0001 ,
		_w11962_,
		_w12651_
	);
	LUT2 #(
		.INIT('h8)
	) name12120 (
		_w11966_,
		_w12651_,
		_w12652_
	);
	LUT2 #(
		.INIT('h1)
	) name12121 (
		_w12008_,
		_w12027_,
		_w12653_
	);
	LUT2 #(
		.INIT('h1)
	) name12122 (
		_w12007_,
		_w12035_,
		_w12654_
	);
	LUT2 #(
		.INIT('h1)
	) name12123 (
		\sa00_reg[5]/P0001 ,
		_w11959_,
		_w12655_
	);
	LUT2 #(
		.INIT('h1)
	) name12124 (
		_w12654_,
		_w12655_,
		_w12656_
	);
	LUT2 #(
		.INIT('h2)
	) name12125 (
		_w12653_,
		_w12656_,
		_w12657_
	);
	LUT2 #(
		.INIT('h1)
	) name12126 (
		\sa00_reg[2]/P0001 ,
		_w12657_,
		_w12658_
	);
	LUT2 #(
		.INIT('h2)
	) name12127 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[2]/P0001 ,
		_w12659_
	);
	LUT2 #(
		.INIT('h8)
	) name12128 (
		\sa00_reg[5]/P0001 ,
		_w11966_,
		_w12660_
	);
	LUT2 #(
		.INIT('h1)
	) name12129 (
		_w12625_,
		_w12629_,
		_w12661_
	);
	LUT2 #(
		.INIT('h4)
	) name12130 (
		_w12660_,
		_w12661_,
		_w12662_
	);
	LUT2 #(
		.INIT('h2)
	) name12131 (
		_w12659_,
		_w12662_,
		_w12663_
	);
	LUT2 #(
		.INIT('h1)
	) name12132 (
		_w11994_,
		_w12614_,
		_w12664_
	);
	LUT2 #(
		.INIT('h2)
	) name12133 (
		\sa00_reg[7]/NET0131 ,
		_w12664_,
		_w12665_
	);
	LUT2 #(
		.INIT('h4)
	) name12134 (
		\sa00_reg[6]/NET0131 ,
		_w11982_,
		_w12666_
	);
	LUT2 #(
		.INIT('h8)
	) name12135 (
		_w12026_,
		_w12666_,
		_w12667_
	);
	LUT2 #(
		.INIT('h1)
	) name12136 (
		_w11958_,
		_w12667_,
		_w12668_
	);
	LUT2 #(
		.INIT('h4)
	) name12137 (
		_w12665_,
		_w12668_,
		_w12669_
	);
	LUT2 #(
		.INIT('h2)
	) name12138 (
		\sa00_reg[1]/P0001 ,
		_w12669_,
		_w12670_
	);
	LUT2 #(
		.INIT('h4)
	) name12139 (
		_w12056_,
		_w12651_,
		_w12671_
	);
	LUT2 #(
		.INIT('h4)
	) name12140 (
		\sa00_reg[2]/P0001 ,
		_w11993_,
		_w12672_
	);
	LUT2 #(
		.INIT('h1)
	) name12141 (
		_w11983_,
		_w12082_,
		_w12673_
	);
	LUT2 #(
		.INIT('h2)
	) name12142 (
		\sa00_reg[2]/P0001 ,
		_w12673_,
		_w12674_
	);
	LUT2 #(
		.INIT('h1)
	) name12143 (
		_w12647_,
		_w12671_,
		_w12675_
	);
	LUT2 #(
		.INIT('h4)
	) name12144 (
		_w12672_,
		_w12675_,
		_w12676_
	);
	LUT2 #(
		.INIT('h4)
	) name12145 (
		_w12674_,
		_w12676_,
		_w12677_
	);
	LUT2 #(
		.INIT('h1)
	) name12146 (
		\sa00_reg[1]/P0001 ,
		_w12677_,
		_w12678_
	);
	LUT2 #(
		.INIT('h1)
	) name12147 (
		_w12650_,
		_w12652_,
		_w12679_
	);
	LUT2 #(
		.INIT('h1)
	) name12148 (
		_w12658_,
		_w12663_,
		_w12680_
	);
	LUT2 #(
		.INIT('h8)
	) name12149 (
		_w12679_,
		_w12680_,
		_w12681_
	);
	LUT2 #(
		.INIT('h4)
	) name12150 (
		_w12670_,
		_w12681_,
		_w12682_
	);
	LUT2 #(
		.INIT('h4)
	) name12151 (
		_w12678_,
		_w12682_,
		_w12683_
	);
	LUT2 #(
		.INIT('h2)
	) name12152 (
		\sa00_reg[0]/P0001 ,
		_w12683_,
		_w12684_
	);
	LUT2 #(
		.INIT('h4)
	) name12153 (
		\sa00_reg[5]/P0001 ,
		_w11952_,
		_w12685_
	);
	LUT2 #(
		.INIT('h4)
	) name12154 (
		\sa00_reg[5]/P0001 ,
		_w11962_,
		_w12686_
	);
	LUT2 #(
		.INIT('h1)
	) name12155 (
		_w12685_,
		_w12686_,
		_w12687_
	);
	LUT2 #(
		.INIT('h4)
	) name12156 (
		_w11996_,
		_w12687_,
		_w12688_
	);
	LUT2 #(
		.INIT('h2)
	) name12157 (
		_w12097_,
		_w12688_,
		_w12689_
	);
	LUT2 #(
		.INIT('h8)
	) name12158 (
		_w12094_,
		_w12666_,
		_w12690_
	);
	LUT2 #(
		.INIT('h8)
	) name12159 (
		_w11956_,
		_w12005_,
		_w12691_
	);
	LUT2 #(
		.INIT('h8)
	) name12160 (
		_w11959_,
		_w12035_,
		_w12692_
	);
	LUT2 #(
		.INIT('h4)
	) name12161 (
		\sa00_reg[3]/P0001 ,
		_w12014_,
		_w12693_
	);
	LUT2 #(
		.INIT('h8)
	) name12162 (
		\sa00_reg[7]/NET0131 ,
		_w12693_,
		_w12694_
	);
	LUT2 #(
		.INIT('h1)
	) name12163 (
		_w12018_,
		_w12692_,
		_w12695_
	);
	LUT2 #(
		.INIT('h4)
	) name12164 (
		_w12694_,
		_w12695_,
		_w12696_
	);
	LUT2 #(
		.INIT('h1)
	) name12165 (
		\sa00_reg[2]/P0001 ,
		_w12696_,
		_w12697_
	);
	LUT2 #(
		.INIT('h1)
	) name12166 (
		_w12690_,
		_w12691_,
		_w12698_
	);
	LUT2 #(
		.INIT('h4)
	) name12167 (
		_w12689_,
		_w12698_,
		_w12699_
	);
	LUT2 #(
		.INIT('h4)
	) name12168 (
		_w12697_,
		_w12699_,
		_w12700_
	);
	LUT2 #(
		.INIT('h1)
	) name12169 (
		\sa00_reg[1]/P0001 ,
		_w12700_,
		_w12701_
	);
	LUT2 #(
		.INIT('h4)
	) name12170 (
		\sa00_reg[7]/NET0131 ,
		_w12690_,
		_w12702_
	);
	LUT2 #(
		.INIT('h1)
	) name12171 (
		_w11968_,
		_w12033_,
		_w12703_
	);
	LUT2 #(
		.INIT('h1)
	) name12172 (
		\sa00_reg[2]/P0001 ,
		_w12703_,
		_w12704_
	);
	LUT2 #(
		.INIT('h8)
	) name12173 (
		_w11994_,
		_w12064_,
		_w12705_
	);
	LUT2 #(
		.INIT('h8)
	) name12174 (
		_w12056_,
		_w12605_,
		_w12706_
	);
	LUT2 #(
		.INIT('h1)
	) name12175 (
		_w12631_,
		_w12705_,
		_w12707_
	);
	LUT2 #(
		.INIT('h4)
	) name12176 (
		_w12706_,
		_w12707_,
		_w12708_
	);
	LUT2 #(
		.INIT('h2)
	) name12177 (
		\sa00_reg[1]/P0001 ,
		_w12708_,
		_w12709_
	);
	LUT2 #(
		.INIT('h1)
	) name12178 (
		_w12702_,
		_w12704_,
		_w12710_
	);
	LUT2 #(
		.INIT('h4)
	) name12179 (
		_w12709_,
		_w12710_,
		_w12711_
	);
	LUT2 #(
		.INIT('h4)
	) name12180 (
		_w12701_,
		_w12711_,
		_w12712_
	);
	LUT2 #(
		.INIT('h4)
	) name12181 (
		_w12684_,
		_w12712_,
		_w12713_
	);
	LUT2 #(
		.INIT('h4)
	) name12182 (
		_w12646_,
		_w12713_,
		_w12714_
	);
	LUT2 #(
		.INIT('h1)
	) name12183 (
		\sa22_reg[5]/P0001 ,
		_w12300_,
		_w12715_
	);
	LUT2 #(
		.INIT('h8)
	) name12184 (
		\sa22_reg[3]/P0001 ,
		_w12715_,
		_w12716_
	);
	LUT2 #(
		.INIT('h4)
	) name12185 (
		\sa22_reg[3]/P0001 ,
		_w12296_,
		_w12717_
	);
	LUT2 #(
		.INIT('h1)
	) name12186 (
		_w12281_,
		_w12716_,
		_w12718_
	);
	LUT2 #(
		.INIT('h4)
	) name12187 (
		_w12717_,
		_w12718_,
		_w12719_
	);
	LUT2 #(
		.INIT('h1)
	) name12188 (
		\sa22_reg[2]/P0001 ,
		_w12719_,
		_w12720_
	);
	LUT2 #(
		.INIT('h8)
	) name12189 (
		\sa22_reg[3]/P0001 ,
		_w12257_,
		_w12721_
	);
	LUT2 #(
		.INIT('h8)
	) name12190 (
		_w12297_,
		_w12721_,
		_w12722_
	);
	LUT2 #(
		.INIT('h8)
	) name12191 (
		_w12278_,
		_w12350_,
		_w12723_
	);
	LUT2 #(
		.INIT('h4)
	) name12192 (
		\sa22_reg[4]/P0001 ,
		_w12324_,
		_w12724_
	);
	LUT2 #(
		.INIT('h8)
	) name12193 (
		_w12252_,
		_w12322_,
		_w12725_
	);
	LUT2 #(
		.INIT('h1)
	) name12194 (
		_w12722_,
		_w12723_,
		_w12726_
	);
	LUT2 #(
		.INIT('h1)
	) name12195 (
		_w12724_,
		_w12725_,
		_w12727_
	);
	LUT2 #(
		.INIT('h8)
	) name12196 (
		_w12726_,
		_w12727_,
		_w12728_
	);
	LUT2 #(
		.INIT('h4)
	) name12197 (
		_w12720_,
		_w12728_,
		_w12729_
	);
	LUT2 #(
		.INIT('h2)
	) name12198 (
		\sa22_reg[1]/P0001 ,
		_w12729_,
		_w12730_
	);
	LUT2 #(
		.INIT('h1)
	) name12199 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w12731_
	);
	LUT2 #(
		.INIT('h8)
	) name12200 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w12732_
	);
	LUT2 #(
		.INIT('h8)
	) name12201 (
		_w12277_,
		_w12732_,
		_w12733_
	);
	LUT2 #(
		.INIT('h8)
	) name12202 (
		_w12731_,
		_w12733_,
		_w12734_
	);
	LUT2 #(
		.INIT('h8)
	) name12203 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		_w12735_
	);
	LUT2 #(
		.INIT('h8)
	) name12204 (
		\sa22_reg[4]/P0001 ,
		_w12239_,
		_w12736_
	);
	LUT2 #(
		.INIT('h8)
	) name12205 (
		_w12735_,
		_w12736_,
		_w12737_
	);
	LUT2 #(
		.INIT('h8)
	) name12206 (
		_w12267_,
		_w12300_,
		_w12738_
	);
	LUT2 #(
		.INIT('h1)
	) name12207 (
		_w12346_,
		_w12738_,
		_w12739_
	);
	LUT2 #(
		.INIT('h1)
	) name12208 (
		\sa22_reg[3]/P0001 ,
		_w12739_,
		_w12740_
	);
	LUT2 #(
		.INIT('h4)
	) name12209 (
		\sa22_reg[3]/P0001 ,
		_w12314_,
		_w12741_
	);
	LUT2 #(
		.INIT('h4)
	) name12210 (
		\sa22_reg[6]/NET0131 ,
		_w12289_,
		_w12742_
	);
	LUT2 #(
		.INIT('h1)
	) name12211 (
		_w12741_,
		_w12742_,
		_w12743_
	);
	LUT2 #(
		.INIT('h2)
	) name12212 (
		\sa22_reg[2]/P0001 ,
		_w12743_,
		_w12744_
	);
	LUT2 #(
		.INIT('h4)
	) name12213 (
		\sa22_reg[7]/NET0131 ,
		_w12336_,
		_w12745_
	);
	LUT2 #(
		.INIT('h8)
	) name12214 (
		\sa22_reg[2]/P0001 ,
		_w12736_,
		_w12746_
	);
	LUT2 #(
		.INIT('h4)
	) name12215 (
		\sa22_reg[3]/P0001 ,
		_w12321_,
		_w12747_
	);
	LUT2 #(
		.INIT('h4)
	) name12216 (
		\sa22_reg[2]/P0001 ,
		_w12747_,
		_w12748_
	);
	LUT2 #(
		.INIT('h1)
	) name12217 (
		_w12279_,
		_w12745_,
		_w12749_
	);
	LUT2 #(
		.INIT('h4)
	) name12218 (
		_w12746_,
		_w12749_,
		_w12750_
	);
	LUT2 #(
		.INIT('h4)
	) name12219 (
		_w12748_,
		_w12750_,
		_w12751_
	);
	LUT2 #(
		.INIT('h1)
	) name12220 (
		\sa22_reg[1]/P0001 ,
		_w12751_,
		_w12752_
	);
	LUT2 #(
		.INIT('h8)
	) name12221 (
		\sa22_reg[5]/P0001 ,
		_w12266_,
		_w12753_
	);
	LUT2 #(
		.INIT('h4)
	) name12222 (
		_w12303_,
		_w12753_,
		_w12754_
	);
	LUT2 #(
		.INIT('h4)
	) name12223 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w12755_
	);
	LUT2 #(
		.INIT('h8)
	) name12224 (
		_w12234_,
		_w12755_,
		_w12756_
	);
	LUT2 #(
		.INIT('h1)
	) name12225 (
		_w12754_,
		_w12756_,
		_w12757_
	);
	LUT2 #(
		.INIT('h1)
	) name12226 (
		\sa22_reg[2]/P0001 ,
		_w12757_,
		_w12758_
	);
	LUT2 #(
		.INIT('h8)
	) name12227 (
		_w12251_,
		_w12260_,
		_w12759_
	);
	LUT2 #(
		.INIT('h8)
	) name12228 (
		\sa22_reg[2]/P0001 ,
		_w12321_,
		_w12760_
	);
	LUT2 #(
		.INIT('h8)
	) name12229 (
		_w12322_,
		_w12344_,
		_w12761_
	);
	LUT2 #(
		.INIT('h1)
	) name12230 (
		_w12759_,
		_w12760_,
		_w12762_
	);
	LUT2 #(
		.INIT('h4)
	) name12231 (
		_w12761_,
		_w12762_,
		_w12763_
	);
	LUT2 #(
		.INIT('h4)
	) name12232 (
		_w12758_,
		_w12763_,
		_w12764_
	);
	LUT2 #(
		.INIT('h2)
	) name12233 (
		\sa22_reg[1]/P0001 ,
		_w12764_,
		_w12765_
	);
	LUT2 #(
		.INIT('h1)
	) name12234 (
		_w12740_,
		_w12744_,
		_w12766_
	);
	LUT2 #(
		.INIT('h4)
	) name12235 (
		_w12752_,
		_w12766_,
		_w12767_
	);
	LUT2 #(
		.INIT('h4)
	) name12236 (
		_w12765_,
		_w12767_,
		_w12768_
	);
	LUT2 #(
		.INIT('h1)
	) name12237 (
		\sa22_reg[0]/P0001 ,
		_w12768_,
		_w12769_
	);
	LUT2 #(
		.INIT('h2)
	) name12238 (
		\sa22_reg[1]/P0001 ,
		_w12390_,
		_w12770_
	);
	LUT2 #(
		.INIT('h8)
	) name12239 (
		_w12278_,
		_w12755_,
		_w12771_
	);
	LUT2 #(
		.INIT('h4)
	) name12240 (
		\sa22_reg[4]/P0001 ,
		_w12251_,
		_w12772_
	);
	LUT2 #(
		.INIT('h8)
	) name12241 (
		_w12234_,
		_w12297_,
		_w12773_
	);
	LUT2 #(
		.INIT('h1)
	) name12242 (
		_w12772_,
		_w12773_,
		_w12774_
	);
	LUT2 #(
		.INIT('h1)
	) name12243 (
		\sa22_reg[2]/P0001 ,
		_w12774_,
		_w12775_
	);
	LUT2 #(
		.INIT('h1)
	) name12244 (
		_w12335_,
		_w12771_,
		_w12776_
	);
	LUT2 #(
		.INIT('h8)
	) name12245 (
		_w12770_,
		_w12776_,
		_w12777_
	);
	LUT2 #(
		.INIT('h4)
	) name12246 (
		_w12775_,
		_w12777_,
		_w12778_
	);
	LUT2 #(
		.INIT('h1)
	) name12247 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w12779_
	);
	LUT2 #(
		.INIT('h8)
	) name12248 (
		_w12315_,
		_w12779_,
		_w12780_
	);
	LUT2 #(
		.INIT('h1)
	) name12249 (
		\sa22_reg[1]/P0001 ,
		_w12780_,
		_w12781_
	);
	LUT2 #(
		.INIT('h8)
	) name12250 (
		_w12732_,
		_w12755_,
		_w12782_
	);
	LUT2 #(
		.INIT('h1)
	) name12251 (
		\sa22_reg[3]/P0001 ,
		_w12731_,
		_w12783_
	);
	LUT2 #(
		.INIT('h2)
	) name12252 (
		_w12249_,
		_w12783_,
		_w12784_
	);
	LUT2 #(
		.INIT('h8)
	) name12253 (
		\sa22_reg[2]/P0001 ,
		_w12298_,
		_w12785_
	);
	LUT2 #(
		.INIT('h1)
	) name12254 (
		_w12782_,
		_w12784_,
		_w12786_
	);
	LUT2 #(
		.INIT('h4)
	) name12255 (
		_w12785_,
		_w12786_,
		_w12787_
	);
	LUT2 #(
		.INIT('h8)
	) name12256 (
		_w12781_,
		_w12787_,
		_w12788_
	);
	LUT2 #(
		.INIT('h1)
	) name12257 (
		_w12778_,
		_w12788_,
		_w12789_
	);
	LUT2 #(
		.INIT('h8)
	) name12258 (
		_w12291_,
		_w12732_,
		_w12790_
	);
	LUT2 #(
		.INIT('h1)
	) name12259 (
		\sa22_reg[2]/P0001 ,
		_w12790_,
		_w12791_
	);
	LUT2 #(
		.INIT('h4)
	) name12260 (
		_w12353_,
		_w12791_,
		_w12792_
	);
	LUT2 #(
		.INIT('h4)
	) name12261 (
		_w12717_,
		_w12792_,
		_w12793_
	);
	LUT2 #(
		.INIT('h2)
	) name12262 (
		\sa22_reg[2]/P0001 ,
		_w12324_,
		_w12794_
	);
	LUT2 #(
		.INIT('h8)
	) name12263 (
		_w12249_,
		_w12290_,
		_w12795_
	);
	LUT2 #(
		.INIT('h1)
	) name12264 (
		_w12334_,
		_w12336_,
		_w12796_
	);
	LUT2 #(
		.INIT('h4)
	) name12265 (
		_w12795_,
		_w12796_,
		_w12797_
	);
	LUT2 #(
		.INIT('h8)
	) name12266 (
		_w12794_,
		_w12797_,
		_w12798_
	);
	LUT2 #(
		.INIT('h1)
	) name12267 (
		_w12793_,
		_w12798_,
		_w12799_
	);
	LUT2 #(
		.INIT('h1)
	) name12268 (
		_w12789_,
		_w12799_,
		_w12800_
	);
	LUT2 #(
		.INIT('h2)
	) name12269 (
		\sa22_reg[0]/P0001 ,
		_w12800_,
		_w12801_
	);
	LUT2 #(
		.INIT('h4)
	) name12270 (
		\sa22_reg[3]/P0001 ,
		_w12738_,
		_w12802_
	);
	LUT2 #(
		.INIT('h1)
	) name12271 (
		_w12244_,
		_w12258_,
		_w12803_
	);
	LUT2 #(
		.INIT('h2)
	) name12272 (
		_w12257_,
		_w12803_,
		_w12804_
	);
	LUT2 #(
		.INIT('h8)
	) name12273 (
		\sa22_reg[7]/NET0131 ,
		_w12732_,
		_w12805_
	);
	LUT2 #(
		.INIT('h8)
	) name12274 (
		_w12267_,
		_w12805_,
		_w12806_
	);
	LUT2 #(
		.INIT('h1)
	) name12275 (
		\sa22_reg[2]/P0001 ,
		_w12806_,
		_w12807_
	);
	LUT2 #(
		.INIT('h4)
	) name12276 (
		_w12804_,
		_w12807_,
		_w12808_
	);
	LUT2 #(
		.INIT('h8)
	) name12277 (
		_w12234_,
		_w12385_,
		_w12809_
	);
	LUT2 #(
		.INIT('h2)
	) name12278 (
		\sa22_reg[2]/P0001 ,
		_w12809_,
		_w12810_
	);
	LUT2 #(
		.INIT('h8)
	) name12279 (
		\sa22_reg[3]/P0001 ,
		_w12297_,
		_w12811_
	);
	LUT2 #(
		.INIT('h8)
	) name12280 (
		_w12234_,
		_w12811_,
		_w12812_
	);
	LUT2 #(
		.INIT('h4)
	) name12281 (
		\sa22_reg[3]/P0001 ,
		_w12332_,
		_w12813_
	);
	LUT2 #(
		.INIT('h8)
	) name12282 (
		_w12263_,
		_w12267_,
		_w12814_
	);
	LUT2 #(
		.INIT('h1)
	) name12283 (
		_w12351_,
		_w12814_,
		_w12815_
	);
	LUT2 #(
		.INIT('h1)
	) name12284 (
		_w12812_,
		_w12813_,
		_w12816_
	);
	LUT2 #(
		.INIT('h8)
	) name12285 (
		_w12815_,
		_w12816_,
		_w12817_
	);
	LUT2 #(
		.INIT('h8)
	) name12286 (
		_w12810_,
		_w12817_,
		_w12818_
	);
	LUT2 #(
		.INIT('h1)
	) name12287 (
		_w12808_,
		_w12818_,
		_w12819_
	);
	LUT2 #(
		.INIT('h1)
	) name12288 (
		_w12384_,
		_w12802_,
		_w12820_
	);
	LUT2 #(
		.INIT('h4)
	) name12289 (
		_w12819_,
		_w12820_,
		_w12821_
	);
	LUT2 #(
		.INIT('h1)
	) name12290 (
		\sa22_reg[1]/P0001 ,
		_w12821_,
		_w12822_
	);
	LUT2 #(
		.INIT('h1)
	) name12291 (
		_w12734_,
		_w12737_,
		_w12823_
	);
	LUT2 #(
		.INIT('h4)
	) name12292 (
		_w12730_,
		_w12823_,
		_w12824_
	);
	LUT2 #(
		.INIT('h4)
	) name12293 (
		_w12801_,
		_w12824_,
		_w12825_
	);
	LUT2 #(
		.INIT('h4)
	) name12294 (
		_w12822_,
		_w12825_,
		_w12826_
	);
	LUT2 #(
		.INIT('h4)
	) name12295 (
		_w12769_,
		_w12826_,
		_w12827_
	);
	LUT2 #(
		.INIT('h2)
	) name12296 (
		_w11951_,
		_w12827_,
		_w12828_
	);
	LUT2 #(
		.INIT('h4)
	) name12297 (
		_w11951_,
		_w12827_,
		_w12829_
	);
	LUT2 #(
		.INIT('h1)
	) name12298 (
		_w12828_,
		_w12829_,
		_w12830_
	);
	LUT2 #(
		.INIT('h1)
	) name12299 (
		_w12714_,
		_w12830_,
		_w12831_
	);
	LUT2 #(
		.INIT('h8)
	) name12300 (
		_w12714_,
		_w12830_,
		_w12832_
	);
	LUT2 #(
		.INIT('h1)
	) name12301 (
		_w12831_,
		_w12832_,
		_w12833_
	);
	LUT2 #(
		.INIT('h2)
	) name12302 (
		\u0_w_reg[0][21]/P0001 ,
		_w12580_,
		_w12834_
	);
	LUT2 #(
		.INIT('h4)
	) name12303 (
		\u0_w_reg[0][21]/P0001 ,
		_w12580_,
		_w12835_
	);
	LUT2 #(
		.INIT('h1)
	) name12304 (
		_w12834_,
		_w12835_,
		_w12836_
	);
	LUT2 #(
		.INIT('h8)
	) name12305 (
		_w12405_,
		_w12836_,
		_w12837_
	);
	LUT2 #(
		.INIT('h1)
	) name12306 (
		_w12405_,
		_w12836_,
		_w12838_
	);
	LUT2 #(
		.INIT('h1)
	) name12307 (
		_w12837_,
		_w12838_,
		_w12839_
	);
	LUT2 #(
		.INIT('h1)
	) name12308 (
		_w12833_,
		_w12839_,
		_w12840_
	);
	LUT2 #(
		.INIT('h8)
	) name12309 (
		_w12833_,
		_w12839_,
		_w12841_
	);
	LUT2 #(
		.INIT('h1)
	) name12310 (
		\ld_r_reg/P0001 ,
		_w12840_,
		_w12842_
	);
	LUT2 #(
		.INIT('h4)
	) name12311 (
		_w12841_,
		_w12842_,
		_w12843_
	);
	LUT2 #(
		.INIT('h2)
	) name12312 (
		\text_in_r_reg[117]/P0001 ,
		\u0_w_reg[0][21]/P0001 ,
		_w12844_
	);
	LUT2 #(
		.INIT('h4)
	) name12313 (
		\text_in_r_reg[117]/P0001 ,
		\u0_w_reg[0][21]/P0001 ,
		_w12845_
	);
	LUT2 #(
		.INIT('h2)
	) name12314 (
		\ld_r_reg/P0001 ,
		_w12844_,
		_w12846_
	);
	LUT2 #(
		.INIT('h4)
	) name12315 (
		_w12845_,
		_w12846_,
		_w12847_
	);
	LUT2 #(
		.INIT('h1)
	) name12316 (
		_w12843_,
		_w12847_,
		_w12848_
	);
	LUT2 #(
		.INIT('h2)
	) name12317 (
		_w12233_,
		_w12714_,
		_w12849_
	);
	LUT2 #(
		.INIT('h4)
	) name12318 (
		_w12233_,
		_w12714_,
		_w12850_
	);
	LUT2 #(
		.INIT('h1)
	) name12319 (
		_w12849_,
		_w12850_,
		_w12851_
	);
	LUT2 #(
		.INIT('h1)
	) name12320 (
		_w12827_,
		_w12851_,
		_w12852_
	);
	LUT2 #(
		.INIT('h8)
	) name12321 (
		_w12827_,
		_w12851_,
		_w12853_
	);
	LUT2 #(
		.INIT('h1)
	) name12322 (
		_w12852_,
		_w12853_,
		_w12854_
	);
	LUT2 #(
		.INIT('h2)
	) name12323 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w12855_
	);
	LUT2 #(
		.INIT('h8)
	) name12324 (
		_w12481_,
		_w12855_,
		_w12856_
	);
	LUT2 #(
		.INIT('h1)
	) name12325 (
		_w12419_,
		_w12479_,
		_w12857_
	);
	LUT2 #(
		.INIT('h8)
	) name12326 (
		_w12527_,
		_w12857_,
		_w12858_
	);
	LUT2 #(
		.INIT('h2)
	) name12327 (
		\sa33_reg[2]/P0001 ,
		_w12493_,
		_w12859_
	);
	LUT2 #(
		.INIT('h4)
	) name12328 (
		_w12858_,
		_w12859_,
		_w12860_
	);
	LUT2 #(
		.INIT('h8)
	) name12329 (
		_w12412_,
		_w12426_,
		_w12861_
	);
	LUT2 #(
		.INIT('h1)
	) name12330 (
		\sa33_reg[2]/P0001 ,
		_w12861_,
		_w12862_
	);
	LUT2 #(
		.INIT('h4)
	) name12331 (
		\sa33_reg[5]/P0001 ,
		_w12549_,
		_w12863_
	);
	LUT2 #(
		.INIT('h8)
	) name12332 (
		_w12414_,
		_w12476_,
		_w12864_
	);
	LUT2 #(
		.INIT('h2)
	) name12333 (
		_w12862_,
		_w12864_,
		_w12865_
	);
	LUT2 #(
		.INIT('h4)
	) name12334 (
		_w12863_,
		_w12865_,
		_w12866_
	);
	LUT2 #(
		.INIT('h1)
	) name12335 (
		_w12860_,
		_w12866_,
		_w12867_
	);
	LUT2 #(
		.INIT('h2)
	) name12336 (
		\sa33_reg[7]/NET0131 ,
		_w12475_,
		_w12868_
	);
	LUT2 #(
		.INIT('h1)
	) name12337 (
		\sa33_reg[2]/P0001 ,
		_w12527_,
		_w12869_
	);
	LUT2 #(
		.INIT('h4)
	) name12338 (
		_w12868_,
		_w12869_,
		_w12870_
	);
	LUT2 #(
		.INIT('h2)
	) name12339 (
		\sa33_reg[1]/P0001 ,
		_w12566_,
		_w12871_
	);
	LUT2 #(
		.INIT('h8)
	) name12340 (
		_w12409_,
		_w12855_,
		_w12872_
	);
	LUT2 #(
		.INIT('h1)
	) name12341 (
		_w12508_,
		_w12872_,
		_w12873_
	);
	LUT2 #(
		.INIT('h4)
	) name12342 (
		_w12870_,
		_w12873_,
		_w12874_
	);
	LUT2 #(
		.INIT('h8)
	) name12343 (
		_w12871_,
		_w12874_,
		_w12875_
	);
	LUT2 #(
		.INIT('h4)
	) name12344 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w12876_
	);
	LUT2 #(
		.INIT('h8)
	) name12345 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w12877_
	);
	LUT2 #(
		.INIT('h8)
	) name12346 (
		_w12876_,
		_w12877_,
		_w12878_
	);
	LUT2 #(
		.INIT('h1)
	) name12347 (
		\sa33_reg[1]/P0001 ,
		_w12878_,
		_w12879_
	);
	LUT2 #(
		.INIT('h4)
	) name12348 (
		\sa33_reg[6]/P0001 ,
		_w12419_,
		_w12880_
	);
	LUT2 #(
		.INIT('h1)
	) name12349 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w12881_
	);
	LUT2 #(
		.INIT('h8)
	) name12350 (
		_w12880_,
		_w12881_,
		_w12882_
	);
	LUT2 #(
		.INIT('h8)
	) name12351 (
		\sa33_reg[2]/P0001 ,
		_w12468_,
		_w12883_
	);
	LUT2 #(
		.INIT('h1)
	) name12352 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w12884_
	);
	LUT2 #(
		.INIT('h1)
	) name12353 (
		\sa33_reg[3]/P0001 ,
		_w12884_,
		_w12885_
	);
	LUT2 #(
		.INIT('h2)
	) name12354 (
		_w12418_,
		_w12885_,
		_w12886_
	);
	LUT2 #(
		.INIT('h2)
	) name12355 (
		_w12879_,
		_w12882_,
		_w12887_
	);
	LUT2 #(
		.INIT('h1)
	) name12356 (
		_w12883_,
		_w12886_,
		_w12888_
	);
	LUT2 #(
		.INIT('h8)
	) name12357 (
		_w12887_,
		_w12888_,
		_w12889_
	);
	LUT2 #(
		.INIT('h1)
	) name12358 (
		_w12875_,
		_w12889_,
		_w12890_
	);
	LUT2 #(
		.INIT('h1)
	) name12359 (
		_w12856_,
		_w12867_,
		_w12891_
	);
	LUT2 #(
		.INIT('h4)
	) name12360 (
		_w12890_,
		_w12891_,
		_w12892_
	);
	LUT2 #(
		.INIT('h2)
	) name12361 (
		\sa33_reg[0]/P0001 ,
		_w12892_,
		_w12893_
	);
	LUT2 #(
		.INIT('h2)
	) name12362 (
		_w12426_,
		_w12465_,
		_w12894_
	);
	LUT2 #(
		.INIT('h1)
	) name12363 (
		_w12482_,
		_w12894_,
		_w12895_
	);
	LUT2 #(
		.INIT('h4)
	) name12364 (
		_w12863_,
		_w12895_,
		_w12896_
	);
	LUT2 #(
		.INIT('h1)
	) name12365 (
		\sa33_reg[2]/P0001 ,
		_w12896_,
		_w12897_
	);
	LUT2 #(
		.INIT('h8)
	) name12366 (
		_w12422_,
		_w12472_,
		_w12898_
	);
	LUT2 #(
		.INIT('h8)
	) name12367 (
		_w12476_,
		_w12544_,
		_w12899_
	);
	LUT2 #(
		.INIT('h8)
	) name12368 (
		_w12413_,
		_w12419_,
		_w12900_
	);
	LUT2 #(
		.INIT('h1)
	) name12369 (
		_w12562_,
		_w12898_,
		_w12901_
	);
	LUT2 #(
		.INIT('h1)
	) name12370 (
		_w12899_,
		_w12900_,
		_w12902_
	);
	LUT2 #(
		.INIT('h8)
	) name12371 (
		_w12901_,
		_w12902_,
		_w12903_
	);
	LUT2 #(
		.INIT('h4)
	) name12372 (
		_w12897_,
		_w12903_,
		_w12904_
	);
	LUT2 #(
		.INIT('h2)
	) name12373 (
		\sa33_reg[1]/P0001 ,
		_w12904_,
		_w12905_
	);
	LUT2 #(
		.INIT('h8)
	) name12374 (
		_w12414_,
		_w12446_,
		_w12906_
	);
	LUT2 #(
		.INIT('h8)
	) name12375 (
		_w12456_,
		_w12906_,
		_w12907_
	);
	LUT2 #(
		.INIT('h8)
	) name12376 (
		_w12480_,
		_w12542_,
		_w12908_
	);
	LUT2 #(
		.INIT('h8)
	) name12377 (
		_w12479_,
		_w12561_,
		_w12909_
	);
	LUT2 #(
		.INIT('h8)
	) name12378 (
		_w12475_,
		_w12551_,
		_w12910_
	);
	LUT2 #(
		.INIT('h2)
	) name12379 (
		\sa33_reg[2]/P0001 ,
		_w12910_,
		_w12911_
	);
	LUT2 #(
		.INIT('h4)
	) name12380 (
		\sa33_reg[3]/P0001 ,
		_w12561_,
		_w12912_
	);
	LUT2 #(
		.INIT('h8)
	) name12381 (
		\sa33_reg[5]/P0001 ,
		_w12531_,
		_w12913_
	);
	LUT2 #(
		.INIT('h8)
	) name12382 (
		_w12432_,
		_w12457_,
		_w12914_
	);
	LUT2 #(
		.INIT('h1)
	) name12383 (
		_w12565_,
		_w12912_,
		_w12915_
	);
	LUT2 #(
		.INIT('h1)
	) name12384 (
		_w12913_,
		_w12914_,
		_w12916_
	);
	LUT2 #(
		.INIT('h8)
	) name12385 (
		_w12915_,
		_w12916_,
		_w12917_
	);
	LUT2 #(
		.INIT('h8)
	) name12386 (
		_w12911_,
		_w12917_,
		_w12918_
	);
	LUT2 #(
		.INIT('h8)
	) name12387 (
		_w12476_,
		_w12481_,
		_w12919_
	);
	LUT2 #(
		.INIT('h1)
	) name12388 (
		\sa33_reg[2]/P0001 ,
		_w12450_,
		_w12920_
	);
	LUT2 #(
		.INIT('h1)
	) name12389 (
		_w12564_,
		_w12919_,
		_w12921_
	);
	LUT2 #(
		.INIT('h8)
	) name12390 (
		_w12920_,
		_w12921_,
		_w12922_
	);
	LUT2 #(
		.INIT('h1)
	) name12391 (
		_w12918_,
		_w12922_,
		_w12923_
	);
	LUT2 #(
		.INIT('h1)
	) name12392 (
		_w12550_,
		_w12909_,
		_w12924_
	);
	LUT2 #(
		.INIT('h4)
	) name12393 (
		_w12923_,
		_w12924_,
		_w12925_
	);
	LUT2 #(
		.INIT('h1)
	) name12394 (
		\sa33_reg[1]/P0001 ,
		_w12925_,
		_w12926_
	);
	LUT2 #(
		.INIT('h4)
	) name12395 (
		\sa33_reg[3]/P0001 ,
		_w12499_,
		_w12927_
	);
	LUT2 #(
		.INIT('h4)
	) name12396 (
		\sa33_reg[1]/P0001 ,
		_w12927_,
		_w12928_
	);
	LUT2 #(
		.INIT('h8)
	) name12397 (
		\sa33_reg[4]/P0001 ,
		_w12564_,
		_w12929_
	);
	LUT2 #(
		.INIT('h1)
	) name12398 (
		_w12928_,
		_w12929_,
		_w12930_
	);
	LUT2 #(
		.INIT('h1)
	) name12399 (
		\sa33_reg[2]/P0001 ,
		_w12930_,
		_w12931_
	);
	LUT2 #(
		.INIT('h8)
	) name12400 (
		\sa33_reg[4]/P0001 ,
		_w12480_,
		_w12932_
	);
	LUT2 #(
		.INIT('h1)
	) name12401 (
		_w12473_,
		_w12932_,
		_w12933_
	);
	LUT2 #(
		.INIT('h2)
	) name12402 (
		\sa33_reg[2]/P0001 ,
		_w12933_,
		_w12934_
	);
	LUT2 #(
		.INIT('h8)
	) name12403 (
		_w12465_,
		_w12476_,
		_w12935_
	);
	LUT2 #(
		.INIT('h1)
	) name12404 (
		_w12934_,
		_w12935_,
		_w12936_
	);
	LUT2 #(
		.INIT('h1)
	) name12405 (
		\sa33_reg[1]/P0001 ,
		_w12936_,
		_w12937_
	);
	LUT2 #(
		.INIT('h8)
	) name12406 (
		_w12479_,
		_w12521_,
		_w12938_
	);
	LUT2 #(
		.INIT('h8)
	) name12407 (
		_w12419_,
		_w12473_,
		_w12939_
	);
	LUT2 #(
		.INIT('h1)
	) name12408 (
		_w12938_,
		_w12939_,
		_w12940_
	);
	LUT2 #(
		.INIT('h2)
	) name12409 (
		\sa33_reg[2]/P0001 ,
		_w12940_,
		_w12941_
	);
	LUT2 #(
		.INIT('h4)
	) name12410 (
		\sa33_reg[2]/P0001 ,
		_w12409_,
		_w12942_
	);
	LUT2 #(
		.INIT('h1)
	) name12411 (
		_w12457_,
		_w12526_,
		_w12943_
	);
	LUT2 #(
		.INIT('h8)
	) name12412 (
		_w12942_,
		_w12943_,
		_w12944_
	);
	LUT2 #(
		.INIT('h8)
	) name12413 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w12945_
	);
	LUT2 #(
		.INIT('h8)
	) name12414 (
		_w12510_,
		_w12945_,
		_w12946_
	);
	LUT2 #(
		.INIT('h8)
	) name12415 (
		_w12461_,
		_w12547_,
		_w12947_
	);
	LUT2 #(
		.INIT('h8)
	) name12416 (
		\sa33_reg[4]/P0001 ,
		_w12531_,
		_w12948_
	);
	LUT2 #(
		.INIT('h1)
	) name12417 (
		_w12946_,
		_w12947_,
		_w12949_
	);
	LUT2 #(
		.INIT('h4)
	) name12418 (
		_w12948_,
		_w12949_,
		_w12950_
	);
	LUT2 #(
		.INIT('h4)
	) name12419 (
		_w12944_,
		_w12950_,
		_w12951_
	);
	LUT2 #(
		.INIT('h2)
	) name12420 (
		\sa33_reg[1]/P0001 ,
		_w12951_,
		_w12952_
	);
	LUT2 #(
		.INIT('h1)
	) name12421 (
		_w12909_,
		_w12941_,
		_w12953_
	);
	LUT2 #(
		.INIT('h4)
	) name12422 (
		_w12931_,
		_w12953_,
		_w12954_
	);
	LUT2 #(
		.INIT('h4)
	) name12423 (
		_w12937_,
		_w12954_,
		_w12955_
	);
	LUT2 #(
		.INIT('h4)
	) name12424 (
		_w12952_,
		_w12955_,
		_w12956_
	);
	LUT2 #(
		.INIT('h1)
	) name12425 (
		\sa33_reg[0]/P0001 ,
		_w12956_,
		_w12957_
	);
	LUT2 #(
		.INIT('h1)
	) name12426 (
		_w12907_,
		_w12908_,
		_w12958_
	);
	LUT2 #(
		.INIT('h4)
	) name12427 (
		_w12905_,
		_w12958_,
		_w12959_
	);
	LUT2 #(
		.INIT('h4)
	) name12428 (
		_w12893_,
		_w12959_,
		_w12960_
	);
	LUT2 #(
		.INIT('h4)
	) name12429 (
		_w12926_,
		_w12960_,
		_w12961_
	);
	LUT2 #(
		.INIT('h4)
	) name12430 (
		_w12957_,
		_w12961_,
		_w12962_
	);
	LUT2 #(
		.INIT('h2)
	) name12431 (
		\u0_w_reg[0][13]/P0001 ,
		_w12962_,
		_w12963_
	);
	LUT2 #(
		.INIT('h4)
	) name12432 (
		\u0_w_reg[0][13]/P0001 ,
		_w12962_,
		_w12964_
	);
	LUT2 #(
		.INIT('h1)
	) name12433 (
		_w12963_,
		_w12964_,
		_w12965_
	);
	LUT2 #(
		.INIT('h8)
	) name12434 (
		_w12580_,
		_w12965_,
		_w12966_
	);
	LUT2 #(
		.INIT('h1)
	) name12435 (
		_w12580_,
		_w12965_,
		_w12967_
	);
	LUT2 #(
		.INIT('h1)
	) name12436 (
		_w12966_,
		_w12967_,
		_w12968_
	);
	LUT2 #(
		.INIT('h4)
	) name12437 (
		_w12854_,
		_w12968_,
		_w12969_
	);
	LUT2 #(
		.INIT('h2)
	) name12438 (
		_w12854_,
		_w12968_,
		_w12970_
	);
	LUT2 #(
		.INIT('h1)
	) name12439 (
		\ld_r_reg/P0001 ,
		_w12969_,
		_w12971_
	);
	LUT2 #(
		.INIT('h4)
	) name12440 (
		_w12970_,
		_w12971_,
		_w12972_
	);
	LUT2 #(
		.INIT('h1)
	) name12441 (
		\text_in_r_reg[109]/P0001 ,
		\u0_w_reg[0][13]/P0001 ,
		_w12973_
	);
	LUT2 #(
		.INIT('h8)
	) name12442 (
		\text_in_r_reg[109]/P0001 ,
		\u0_w_reg[0][13]/P0001 ,
		_w12974_
	);
	LUT2 #(
		.INIT('h2)
	) name12443 (
		\ld_r_reg/P0001 ,
		_w12973_,
		_w12975_
	);
	LUT2 #(
		.INIT('h4)
	) name12444 (
		_w12974_,
		_w12975_,
		_w12976_
	);
	LUT2 #(
		.INIT('h1)
	) name12445 (
		_w12972_,
		_w12976_,
		_w12977_
	);
	LUT2 #(
		.INIT('h1)
	) name12446 (
		_w12111_,
		_w12851_,
		_w12978_
	);
	LUT2 #(
		.INIT('h8)
	) name12447 (
		_w12111_,
		_w12851_,
		_w12979_
	);
	LUT2 #(
		.INIT('h1)
	) name12448 (
		_w12978_,
		_w12979_,
		_w12980_
	);
	LUT2 #(
		.INIT('h2)
	) name12449 (
		\u0_w_reg[0][5]/P0001 ,
		_w12962_,
		_w12981_
	);
	LUT2 #(
		.INIT('h4)
	) name12450 (
		\u0_w_reg[0][5]/P0001 ,
		_w12962_,
		_w12982_
	);
	LUT2 #(
		.INIT('h1)
	) name12451 (
		_w12981_,
		_w12982_,
		_w12983_
	);
	LUT2 #(
		.INIT('h8)
	) name12452 (
		_w12405_,
		_w12983_,
		_w12984_
	);
	LUT2 #(
		.INIT('h1)
	) name12453 (
		_w12405_,
		_w12983_,
		_w12985_
	);
	LUT2 #(
		.INIT('h1)
	) name12454 (
		_w12984_,
		_w12985_,
		_w12986_
	);
	LUT2 #(
		.INIT('h4)
	) name12455 (
		_w12980_,
		_w12986_,
		_w12987_
	);
	LUT2 #(
		.INIT('h2)
	) name12456 (
		_w12980_,
		_w12986_,
		_w12988_
	);
	LUT2 #(
		.INIT('h1)
	) name12457 (
		\ld_r_reg/P0001 ,
		_w12987_,
		_w12989_
	);
	LUT2 #(
		.INIT('h4)
	) name12458 (
		_w12988_,
		_w12989_,
		_w12990_
	);
	LUT2 #(
		.INIT('h1)
	) name12459 (
		\text_in_r_reg[101]/P0001 ,
		\u0_w_reg[0][5]/P0001 ,
		_w12991_
	);
	LUT2 #(
		.INIT('h8)
	) name12460 (
		\text_in_r_reg[101]/P0001 ,
		\u0_w_reg[0][5]/P0001 ,
		_w12992_
	);
	LUT2 #(
		.INIT('h2)
	) name12461 (
		\ld_r_reg/P0001 ,
		_w12991_,
		_w12993_
	);
	LUT2 #(
		.INIT('h4)
	) name12462 (
		_w12992_,
		_w12993_,
		_w12994_
	);
	LUT2 #(
		.INIT('h1)
	) name12463 (
		_w12990_,
		_w12994_,
		_w12995_
	);
	LUT2 #(
		.INIT('h1)
	) name12464 (
		_w12017_,
		_w12647_,
		_w12996_
	);
	LUT2 #(
		.INIT('h4)
	) name12465 (
		\sa00_reg[4]/P0001 ,
		_w12033_,
		_w12997_
	);
	LUT2 #(
		.INIT('h1)
	) name12466 (
		_w12057_,
		_w12612_,
		_w12998_
	);
	LUT2 #(
		.INIT('h4)
	) name12467 (
		_w12997_,
		_w12998_,
		_w12999_
	);
	LUT2 #(
		.INIT('h2)
	) name12468 (
		\sa00_reg[1]/P0001 ,
		_w12999_,
		_w13000_
	);
	LUT2 #(
		.INIT('h4)
	) name12469 (
		_w12630_,
		_w12996_,
		_w13001_
	);
	LUT2 #(
		.INIT('h4)
	) name12470 (
		_w13000_,
		_w13001_,
		_w13002_
	);
	LUT2 #(
		.INIT('h2)
	) name12471 (
		\sa00_reg[2]/P0001 ,
		_w13002_,
		_w13003_
	);
	LUT2 #(
		.INIT('h2)
	) name12472 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w13004_
	);
	LUT2 #(
		.INIT('h8)
	) name12473 (
		_w12613_,
		_w13004_,
		_w13005_
	);
	LUT2 #(
		.INIT('h8)
	) name12474 (
		_w11962_,
		_w12014_,
		_w13006_
	);
	LUT2 #(
		.INIT('h8)
	) name12475 (
		\sa00_reg[1]/P0001 ,
		_w12020_,
		_w13007_
	);
	LUT2 #(
		.INIT('h4)
	) name12476 (
		_w12065_,
		_w13007_,
		_w13008_
	);
	LUT2 #(
		.INIT('h1)
	) name12477 (
		_w12614_,
		_w13006_,
		_w13009_
	);
	LUT2 #(
		.INIT('h4)
	) name12478 (
		_w13008_,
		_w13009_,
		_w13010_
	);
	LUT2 #(
		.INIT('h1)
	) name12479 (
		\sa00_reg[2]/P0001 ,
		_w13010_,
		_w13011_
	);
	LUT2 #(
		.INIT('h4)
	) name12480 (
		\sa00_reg[4]/P0001 ,
		_w11974_,
		_w13012_
	);
	LUT2 #(
		.INIT('h1)
	) name12481 (
		_w12667_,
		_w13012_,
		_w13013_
	);
	LUT2 #(
		.INIT('h2)
	) name12482 (
		\sa00_reg[1]/P0001 ,
		_w13013_,
		_w13014_
	);
	LUT2 #(
		.INIT('h4)
	) name12483 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[2]/P0001 ,
		_w13015_
	);
	LUT2 #(
		.INIT('h1)
	) name12484 (
		_w12050_,
		_w12686_,
		_w13016_
	);
	LUT2 #(
		.INIT('h2)
	) name12485 (
		_w13015_,
		_w13016_,
		_w13017_
	);
	LUT2 #(
		.INIT('h8)
	) name12486 (
		_w11985_,
		_w12015_,
		_w13018_
	);
	LUT2 #(
		.INIT('h1)
	) name12487 (
		_w11976_,
		_w13018_,
		_w13019_
	);
	LUT2 #(
		.INIT('h4)
	) name12488 (
		_w12628_,
		_w13019_,
		_w13020_
	);
	LUT2 #(
		.INIT('h1)
	) name12489 (
		\sa00_reg[1]/P0001 ,
		_w13020_,
		_w13021_
	);
	LUT2 #(
		.INIT('h1)
	) name12490 (
		_w13005_,
		_w13017_,
		_w13022_
	);
	LUT2 #(
		.INIT('h4)
	) name12491 (
		_w13011_,
		_w13022_,
		_w13023_
	);
	LUT2 #(
		.INIT('h4)
	) name12492 (
		_w13014_,
		_w13023_,
		_w13024_
	);
	LUT2 #(
		.INIT('h4)
	) name12493 (
		_w13003_,
		_w13024_,
		_w13025_
	);
	LUT2 #(
		.INIT('h4)
	) name12494 (
		_w13021_,
		_w13025_,
		_w13026_
	);
	LUT2 #(
		.INIT('h2)
	) name12495 (
		\sa00_reg[0]/P0001 ,
		_w13026_,
		_w13027_
	);
	LUT2 #(
		.INIT('h8)
	) name12496 (
		\sa00_reg[4]/P0001 ,
		_w11960_,
		_w13028_
	);
	LUT2 #(
		.INIT('h4)
	) name12497 (
		\sa00_reg[3]/P0001 ,
		_w13028_,
		_w13029_
	);
	LUT2 #(
		.INIT('h4)
	) name12498 (
		\sa00_reg[4]/P0001 ,
		_w12044_,
		_w13030_
	);
	LUT2 #(
		.INIT('h8)
	) name12499 (
		_w11955_,
		_w12026_,
		_w13031_
	);
	LUT2 #(
		.INIT('h8)
	) name12500 (
		\sa00_reg[6]/NET0131 ,
		_w13031_,
		_w13032_
	);
	LUT2 #(
		.INIT('h2)
	) name12501 (
		_w12004_,
		_w13029_,
		_w13033_
	);
	LUT2 #(
		.INIT('h1)
	) name12502 (
		_w13030_,
		_w13032_,
		_w13034_
	);
	LUT2 #(
		.INIT('h8)
	) name12503 (
		_w13033_,
		_w13034_,
		_w13035_
	);
	LUT2 #(
		.INIT('h8)
	) name12504 (
		\sa00_reg[6]/NET0131 ,
		_w11955_,
		_w13036_
	);
	LUT2 #(
		.INIT('h8)
	) name12505 (
		_w12096_,
		_w13036_,
		_w13037_
	);
	LUT2 #(
		.INIT('h4)
	) name12506 (
		\sa00_reg[3]/P0001 ,
		_w12629_,
		_w13038_
	);
	LUT2 #(
		.INIT('h2)
	) name12507 (
		\sa00_reg[2]/P0001 ,
		_w13037_,
		_w13039_
	);
	LUT2 #(
		.INIT('h4)
	) name12508 (
		_w13038_,
		_w13039_,
		_w13040_
	);
	LUT2 #(
		.INIT('h1)
	) name12509 (
		_w13035_,
		_w13040_,
		_w13041_
	);
	LUT2 #(
		.INIT('h4)
	) name12510 (
		\sa00_reg[3]/P0001 ,
		_w11952_,
		_w13042_
	);
	LUT2 #(
		.INIT('h4)
	) name12511 (
		\sa00_reg[4]/P0001 ,
		_w13042_,
		_w13043_
	);
	LUT2 #(
		.INIT('h4)
	) name12512 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		_w13044_
	);
	LUT2 #(
		.INIT('h8)
	) name12513 (
		_w11959_,
		_w13044_,
		_w13045_
	);
	LUT2 #(
		.INIT('h1)
	) name12514 (
		\sa00_reg[1]/P0001 ,
		_w12052_,
		_w13046_
	);
	LUT2 #(
		.INIT('h1)
	) name12515 (
		_w13006_,
		_w13045_,
		_w13047_
	);
	LUT2 #(
		.INIT('h8)
	) name12516 (
		_w13046_,
		_w13047_,
		_w13048_
	);
	LUT2 #(
		.INIT('h1)
	) name12517 (
		_w12055_,
		_w13037_,
		_w13049_
	);
	LUT2 #(
		.INIT('h4)
	) name12518 (
		_w13043_,
		_w13049_,
		_w13050_
	);
	LUT2 #(
		.INIT('h8)
	) name12519 (
		_w13048_,
		_w13050_,
		_w13051_
	);
	LUT2 #(
		.INIT('h2)
	) name12520 (
		_w12056_,
		_w12634_,
		_w13052_
	);
	LUT2 #(
		.INIT('h4)
	) name12521 (
		\sa00_reg[2]/P0001 ,
		_w12630_,
		_w13053_
	);
	LUT2 #(
		.INIT('h2)
	) name12522 (
		\sa00_reg[1]/P0001 ,
		_w12018_,
		_w13054_
	);
	LUT2 #(
		.INIT('h4)
	) name12523 (
		_w13052_,
		_w13054_,
		_w13055_
	);
	LUT2 #(
		.INIT('h4)
	) name12524 (
		_w13053_,
		_w13055_,
		_w13056_
	);
	LUT2 #(
		.INIT('h1)
	) name12525 (
		_w13051_,
		_w13056_,
		_w13057_
	);
	LUT2 #(
		.INIT('h1)
	) name12526 (
		_w13041_,
		_w13057_,
		_w13058_
	);
	LUT2 #(
		.INIT('h1)
	) name12527 (
		\sa00_reg[0]/P0001 ,
		_w13058_,
		_w13059_
	);
	LUT2 #(
		.INIT('h4)
	) name12528 (
		\sa00_reg[2]/P0001 ,
		_w11968_,
		_w13060_
	);
	LUT2 #(
		.INIT('h8)
	) name12529 (
		_w11973_,
		_w11994_,
		_w13061_
	);
	LUT2 #(
		.INIT('h4)
	) name12530 (
		\sa00_reg[6]/NET0131 ,
		_w12625_,
		_w13062_
	);
	LUT2 #(
		.INIT('h1)
	) name12531 (
		_w12691_,
		_w13061_,
		_w13063_
	);
	LUT2 #(
		.INIT('h4)
	) name12532 (
		_w13062_,
		_w13063_,
		_w13064_
	);
	LUT2 #(
		.INIT('h2)
	) name12533 (
		\sa00_reg[2]/P0001 ,
		_w13064_,
		_w13065_
	);
	LUT2 #(
		.INIT('h1)
	) name12534 (
		_w13060_,
		_w13065_,
		_w13066_
	);
	LUT2 #(
		.INIT('h2)
	) name12535 (
		\sa00_reg[1]/P0001 ,
		_w13066_,
		_w13067_
	);
	LUT2 #(
		.INIT('h4)
	) name12536 (
		\sa00_reg[5]/P0001 ,
		_w12057_,
		_w13068_
	);
	LUT2 #(
		.INIT('h4)
	) name12537 (
		\sa00_reg[6]/NET0131 ,
		_w11974_,
		_w13069_
	);
	LUT2 #(
		.INIT('h1)
	) name12538 (
		_w11976_,
		_w13068_,
		_w13070_
	);
	LUT2 #(
		.INIT('h4)
	) name12539 (
		_w13069_,
		_w13070_,
		_w13071_
	);
	LUT2 #(
		.INIT('h1)
	) name12540 (
		\sa00_reg[2]/P0001 ,
		_w13071_,
		_w13072_
	);
	LUT2 #(
		.INIT('h8)
	) name12541 (
		_w11995_,
		_w12005_,
		_w13073_
	);
	LUT2 #(
		.INIT('h4)
	) name12542 (
		\sa00_reg[4]/P0001 ,
		_w12002_,
		_w13074_
	);
	LUT2 #(
		.INIT('h8)
	) name12543 (
		_w12094_,
		_w13074_,
		_w13075_
	);
	LUT2 #(
		.INIT('h8)
	) name12544 (
		_w12054_,
		_w12636_,
		_w13076_
	);
	LUT2 #(
		.INIT('h4)
	) name12545 (
		\sa00_reg[6]/NET0131 ,
		_w12050_,
		_w13077_
	);
	LUT2 #(
		.INIT('h1)
	) name12546 (
		_w13073_,
		_w13075_,
		_w13078_
	);
	LUT2 #(
		.INIT('h1)
	) name12547 (
		_w13076_,
		_w13077_,
		_w13079_
	);
	LUT2 #(
		.INIT('h8)
	) name12548 (
		_w13078_,
		_w13079_,
		_w13080_
	);
	LUT2 #(
		.INIT('h4)
	) name12549 (
		_w13072_,
		_w13080_,
		_w13081_
	);
	LUT2 #(
		.INIT('h1)
	) name12550 (
		\sa00_reg[1]/P0001 ,
		_w13081_,
		_w13082_
	);
	LUT2 #(
		.INIT('h1)
	) name12551 (
		_w12015_,
		_w12017_,
		_w13083_
	);
	LUT2 #(
		.INIT('h2)
	) name12552 (
		_w13004_,
		_w13083_,
		_w13084_
	);
	LUT2 #(
		.INIT('h8)
	) name12553 (
		_w11976_,
		_w13044_,
		_w13085_
	);
	LUT2 #(
		.INIT('h1)
	) name12554 (
		_w12006_,
		_w13085_,
		_w13086_
	);
	LUT2 #(
		.INIT('h4)
	) name12555 (
		_w13084_,
		_w13086_,
		_w13087_
	);
	LUT2 #(
		.INIT('h4)
	) name12556 (
		_w13067_,
		_w13087_,
		_w13088_
	);
	LUT2 #(
		.INIT('h4)
	) name12557 (
		_w13082_,
		_w13088_,
		_w13089_
	);
	LUT2 #(
		.INIT('h4)
	) name12558 (
		_w13059_,
		_w13089_,
		_w13090_
	);
	LUT2 #(
		.INIT('h4)
	) name12559 (
		_w13027_,
		_w13090_,
		_w13091_
	);
	LUT2 #(
		.INIT('h1)
	) name12560 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w13092_
	);
	LUT2 #(
		.INIT('h8)
	) name12561 (
		_w11833_,
		_w13092_,
		_w13093_
	);
	LUT2 #(
		.INIT('h1)
	) name12562 (
		_w12115_,
		_w13093_,
		_w13094_
	);
	LUT2 #(
		.INIT('h1)
	) name12563 (
		\sa11_reg[2]/P0001 ,
		_w13094_,
		_w13095_
	);
	LUT2 #(
		.INIT('h1)
	) name12564 (
		_w11795_,
		_w12186_,
		_w13096_
	);
	LUT2 #(
		.INIT('h1)
	) name12565 (
		_w11909_,
		_w12151_,
		_w13097_
	);
	LUT2 #(
		.INIT('h8)
	) name12566 (
		_w13096_,
		_w13097_,
		_w13098_
	);
	LUT2 #(
		.INIT('h2)
	) name12567 (
		\sa11_reg[2]/P0001 ,
		_w13098_,
		_w13099_
	);
	LUT2 #(
		.INIT('h4)
	) name12568 (
		\sa11_reg[7]/NET0131 ,
		_w12127_,
		_w13100_
	);
	LUT2 #(
		.INIT('h4)
	) name12569 (
		\sa11_reg[3]/P0001 ,
		_w12139_,
		_w13101_
	);
	LUT2 #(
		.INIT('h8)
	) name12570 (
		_w11800_,
		_w11892_,
		_w13102_
	);
	LUT2 #(
		.INIT('h1)
	) name12571 (
		_w13100_,
		_w13102_,
		_w13103_
	);
	LUT2 #(
		.INIT('h4)
	) name12572 (
		_w13101_,
		_w13103_,
		_w13104_
	);
	LUT2 #(
		.INIT('h2)
	) name12573 (
		\sa11_reg[2]/P0001 ,
		_w13104_,
		_w13105_
	);
	LUT2 #(
		.INIT('h1)
	) name12574 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w13106_
	);
	LUT2 #(
		.INIT('h4)
	) name12575 (
		\sa11_reg[5]/P0001 ,
		_w13106_,
		_w13107_
	);
	LUT2 #(
		.INIT('h4)
	) name12576 (
		_w11853_,
		_w13107_,
		_w13108_
	);
	LUT2 #(
		.INIT('h8)
	) name12577 (
		_w11796_,
		_w11892_,
		_w13109_
	);
	LUT2 #(
		.INIT('h1)
	) name12578 (
		_w12177_,
		_w13109_,
		_w13110_
	);
	LUT2 #(
		.INIT('h4)
	) name12579 (
		_w13108_,
		_w13110_,
		_w13111_
	);
	LUT2 #(
		.INIT('h4)
	) name12580 (
		_w13105_,
		_w13111_,
		_w13112_
	);
	LUT2 #(
		.INIT('h2)
	) name12581 (
		\sa11_reg[1]/P0001 ,
		_w13112_,
		_w13113_
	);
	LUT2 #(
		.INIT('h1)
	) name12582 (
		_w11926_,
		_w12194_,
		_w13114_
	);
	LUT2 #(
		.INIT('h2)
	) name12583 (
		\sa11_reg[2]/P0001 ,
		_w13114_,
		_w13115_
	);
	LUT2 #(
		.INIT('h4)
	) name12584 (
		\sa11_reg[2]/P0001 ,
		_w11922_,
		_w13116_
	);
	LUT2 #(
		.INIT('h1)
	) name12585 (
		_w11898_,
		_w13115_,
		_w13117_
	);
	LUT2 #(
		.INIT('h4)
	) name12586 (
		_w13116_,
		_w13117_,
		_w13118_
	);
	LUT2 #(
		.INIT('h4)
	) name12587 (
		_w12141_,
		_w13118_,
		_w13119_
	);
	LUT2 #(
		.INIT('h1)
	) name12588 (
		\sa11_reg[1]/P0001 ,
		_w13119_,
		_w13120_
	);
	LUT2 #(
		.INIT('h1)
	) name12589 (
		_w13095_,
		_w13099_,
		_w13121_
	);
	LUT2 #(
		.INIT('h4)
	) name12590 (
		_w13113_,
		_w13121_,
		_w13122_
	);
	LUT2 #(
		.INIT('h4)
	) name12591 (
		_w13120_,
		_w13122_,
		_w13123_
	);
	LUT2 #(
		.INIT('h2)
	) name12592 (
		\sa11_reg[0]/P0001 ,
		_w13123_,
		_w13124_
	);
	LUT2 #(
		.INIT('h4)
	) name12593 (
		\sa11_reg[4]/P0001 ,
		_w11864_,
		_w13125_
	);
	LUT2 #(
		.INIT('h8)
	) name12594 (
		_w11825_,
		_w11877_,
		_w13126_
	);
	LUT2 #(
		.INIT('h8)
	) name12595 (
		\sa11_reg[6]/NET0131 ,
		_w13126_,
		_w13127_
	);
	LUT2 #(
		.INIT('h2)
	) name12596 (
		_w11914_,
		_w12142_,
		_w13128_
	);
	LUT2 #(
		.INIT('h1)
	) name12597 (
		_w13125_,
		_w13127_,
		_w13129_
	);
	LUT2 #(
		.INIT('h8)
	) name12598 (
		_w13128_,
		_w13129_,
		_w13130_
	);
	LUT2 #(
		.INIT('h8)
	) name12599 (
		\sa11_reg[6]/NET0131 ,
		_w11877_,
		_w13131_
	);
	LUT2 #(
		.INIT('h8)
	) name12600 (
		_w11801_,
		_w13131_,
		_w13132_
	);
	LUT2 #(
		.INIT('h8)
	) name12601 (
		_w11860_,
		_w11876_,
		_w13133_
	);
	LUT2 #(
		.INIT('h2)
	) name12602 (
		\sa11_reg[2]/P0001 ,
		_w13133_,
		_w13134_
	);
	LUT2 #(
		.INIT('h4)
	) name12603 (
		_w13132_,
		_w13134_,
		_w13135_
	);
	LUT2 #(
		.INIT('h1)
	) name12604 (
		_w13130_,
		_w13135_,
		_w13136_
	);
	LUT2 #(
		.INIT('h4)
	) name12605 (
		\sa11_reg[2]/P0001 ,
		_w11926_,
		_w13137_
	);
	LUT2 #(
		.INIT('h8)
	) name12606 (
		_w11796_,
		_w11801_,
		_w13138_
	);
	LUT2 #(
		.INIT('h4)
	) name12607 (
		\sa11_reg[3]/P0001 ,
		_w11870_,
		_w13139_
	);
	LUT2 #(
		.INIT('h4)
	) name12608 (
		\sa11_reg[4]/P0001 ,
		_w13139_,
		_w13140_
	);
	LUT2 #(
		.INIT('h1)
	) name12609 (
		\sa11_reg[1]/P0001 ,
		_w13093_,
		_w13141_
	);
	LUT2 #(
		.INIT('h4)
	) name12610 (
		_w13138_,
		_w13141_,
		_w13142_
	);
	LUT2 #(
		.INIT('h1)
	) name12611 (
		_w11848_,
		_w13132_,
		_w13143_
	);
	LUT2 #(
		.INIT('h1)
	) name12612 (
		_w13137_,
		_w13140_,
		_w13144_
	);
	LUT2 #(
		.INIT('h8)
	) name12613 (
		_w13143_,
		_w13144_,
		_w13145_
	);
	LUT2 #(
		.INIT('h8)
	) name12614 (
		_w13142_,
		_w13145_,
		_w13146_
	);
	LUT2 #(
		.INIT('h2)
	) name12615 (
		_w11805_,
		_w12154_,
		_w13147_
	);
	LUT2 #(
		.INIT('h4)
	) name12616 (
		\sa11_reg[2]/P0001 ,
		_w12151_,
		_w13148_
	);
	LUT2 #(
		.INIT('h2)
	) name12617 (
		\sa11_reg[1]/P0001 ,
		_w11941_,
		_w13149_
	);
	LUT2 #(
		.INIT('h4)
	) name12618 (
		_w13148_,
		_w13149_,
		_w13150_
	);
	LUT2 #(
		.INIT('h4)
	) name12619 (
		_w13147_,
		_w13150_,
		_w13151_
	);
	LUT2 #(
		.INIT('h1)
	) name12620 (
		_w13146_,
		_w13151_,
		_w13152_
	);
	LUT2 #(
		.INIT('h1)
	) name12621 (
		_w13136_,
		_w13152_,
		_w13153_
	);
	LUT2 #(
		.INIT('h1)
	) name12622 (
		\sa11_reg[0]/P0001 ,
		_w13153_,
		_w13154_
	);
	LUT2 #(
		.INIT('h4)
	) name12623 (
		\sa11_reg[6]/NET0131 ,
		_w11926_,
		_w13155_
	);
	LUT2 #(
		.INIT('h1)
	) name12624 (
		_w11830_,
		_w11907_,
		_w13156_
	);
	LUT2 #(
		.INIT('h2)
	) name12625 (
		\sa11_reg[2]/P0001 ,
		_w13156_,
		_w13157_
	);
	LUT2 #(
		.INIT('h2)
	) name12626 (
		_w11798_,
		_w11860_,
		_w13158_
	);
	LUT2 #(
		.INIT('h4)
	) name12627 (
		\sa11_reg[5]/P0001 ,
		_w13100_,
		_w13159_
	);
	LUT2 #(
		.INIT('h1)
	) name12628 (
		_w13158_,
		_w13159_,
		_w13160_
	);
	LUT2 #(
		.INIT('h1)
	) name12629 (
		\sa11_reg[2]/P0001 ,
		_w13160_,
		_w13161_
	);
	LUT2 #(
		.INIT('h1)
	) name12630 (
		_w12124_,
		_w13155_,
		_w13162_
	);
	LUT2 #(
		.INIT('h4)
	) name12631 (
		_w13157_,
		_w13162_,
		_w13163_
	);
	LUT2 #(
		.INIT('h4)
	) name12632 (
		_w13161_,
		_w13163_,
		_w13164_
	);
	LUT2 #(
		.INIT('h1)
	) name12633 (
		\sa11_reg[1]/P0001 ,
		_w13164_,
		_w13165_
	);
	LUT2 #(
		.INIT('h2)
	) name12634 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[2]/P0001 ,
		_w13166_
	);
	LUT2 #(
		.INIT('h8)
	) name12635 (
		_w11881_,
		_w13166_,
		_w13167_
	);
	LUT2 #(
		.INIT('h1)
	) name12636 (
		_w11795_,
		_w12146_,
		_w13168_
	);
	LUT2 #(
		.INIT('h2)
	) name12637 (
		_w12145_,
		_w13168_,
		_w13169_
	);
	LUT2 #(
		.INIT('h8)
	) name12638 (
		\sa11_reg[3]/P0001 ,
		_w12160_,
		_w13170_
	);
	LUT2 #(
		.INIT('h8)
	) name12639 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[2]/P0001 ,
		_w13171_
	);
	LUT2 #(
		.INIT('h4)
	) name12640 (
		\sa11_reg[6]/NET0131 ,
		_w11813_,
		_w13172_
	);
	LUT2 #(
		.INIT('h8)
	) name12641 (
		\sa11_reg[3]/P0001 ,
		_w13102_,
		_w13173_
	);
	LUT2 #(
		.INIT('h1)
	) name12642 (
		_w11865_,
		_w13172_,
		_w13174_
	);
	LUT2 #(
		.INIT('h4)
	) name12643 (
		_w13173_,
		_w13174_,
		_w13175_
	);
	LUT2 #(
		.INIT('h2)
	) name12644 (
		_w13171_,
		_w13175_,
		_w13176_
	);
	LUT2 #(
		.INIT('h1)
	) name12645 (
		_w11866_,
		_w13167_,
		_w13177_
	);
	LUT2 #(
		.INIT('h1)
	) name12646 (
		_w13169_,
		_w13170_,
		_w13178_
	);
	LUT2 #(
		.INIT('h8)
	) name12647 (
		_w13177_,
		_w13178_,
		_w13179_
	);
	LUT2 #(
		.INIT('h4)
	) name12648 (
		_w13176_,
		_w13179_,
		_w13180_
	);
	LUT2 #(
		.INIT('h4)
	) name12649 (
		_w13165_,
		_w13180_,
		_w13181_
	);
	LUT2 #(
		.INIT('h4)
	) name12650 (
		_w13154_,
		_w13181_,
		_w13182_
	);
	LUT2 #(
		.INIT('h4)
	) name12651 (
		_w13124_,
		_w13182_,
		_w13183_
	);
	LUT2 #(
		.INIT('h2)
	) name12652 (
		_w13091_,
		_w13183_,
		_w13184_
	);
	LUT2 #(
		.INIT('h4)
	) name12653 (
		_w13091_,
		_w13183_,
		_w13185_
	);
	LUT2 #(
		.INIT('h1)
	) name12654 (
		_w13184_,
		_w13185_,
		_w13186_
	);
	LUT2 #(
		.INIT('h1)
	) name12655 (
		_w12714_,
		_w13186_,
		_w13187_
	);
	LUT2 #(
		.INIT('h8)
	) name12656 (
		_w12714_,
		_w13186_,
		_w13188_
	);
	LUT2 #(
		.INIT('h1)
	) name12657 (
		_w13187_,
		_w13188_,
		_w13189_
	);
	LUT2 #(
		.INIT('h8)
	) name12658 (
		_w12251_,
		_w12267_,
		_w13190_
	);
	LUT2 #(
		.INIT('h1)
	) name12659 (
		_w12246_,
		_w13190_,
		_w13191_
	);
	LUT2 #(
		.INIT('h1)
	) name12660 (
		\sa22_reg[2]/P0001 ,
		_w13191_,
		_w13192_
	);
	LUT2 #(
		.INIT('h1)
	) name12661 (
		_w12320_,
		_w12759_,
		_w13193_
	);
	LUT2 #(
		.INIT('h1)
	) name12662 (
		_w12296_,
		_w12324_,
		_w13194_
	);
	LUT2 #(
		.INIT('h8)
	) name12663 (
		_w13193_,
		_w13194_,
		_w13195_
	);
	LUT2 #(
		.INIT('h2)
	) name12664 (
		\sa22_reg[2]/P0001 ,
		_w13195_,
		_w13196_
	);
	LUT2 #(
		.INIT('h4)
	) name12665 (
		\sa22_reg[7]/NET0131 ,
		_w12257_,
		_w13197_
	);
	LUT2 #(
		.INIT('h1)
	) name12666 (
		_w12811_,
		_w13197_,
		_w13198_
	);
	LUT2 #(
		.INIT('h2)
	) name12667 (
		\sa22_reg[2]/P0001 ,
		_w13198_,
		_w13199_
	);
	LUT2 #(
		.INIT('h1)
	) name12668 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		_w13200_
	);
	LUT2 #(
		.INIT('h8)
	) name12669 (
		_w12332_,
		_w13200_,
		_w13201_
	);
	LUT2 #(
		.INIT('h1)
	) name12670 (
		_w12298_,
		_w13201_,
		_w13202_
	);
	LUT2 #(
		.INIT('h4)
	) name12671 (
		_w12294_,
		_w13202_,
		_w13203_
	);
	LUT2 #(
		.INIT('h4)
	) name12672 (
		_w13199_,
		_w13203_,
		_w13204_
	);
	LUT2 #(
		.INIT('h1)
	) name12673 (
		\sa22_reg[1]/P0001 ,
		_w13204_,
		_w13205_
	);
	LUT2 #(
		.INIT('h8)
	) name12674 (
		_w12249_,
		_w12303_,
		_w13206_
	);
	LUT2 #(
		.INIT('h1)
	) name12675 (
		_w12333_,
		_w13206_,
		_w13207_
	);
	LUT2 #(
		.INIT('h8)
	) name12676 (
		_w12356_,
		_w13200_,
		_w13208_
	);
	LUT2 #(
		.INIT('h8)
	) name12677 (
		_w12257_,
		_w12385_,
		_w13209_
	);
	LUT2 #(
		.INIT('h1)
	) name12678 (
		_w12252_,
		_w12268_,
		_w13210_
	);
	LUT2 #(
		.INIT('h4)
	) name12679 (
		_w13209_,
		_w13210_,
		_w13211_
	);
	LUT2 #(
		.INIT('h2)
	) name12680 (
		\sa22_reg[2]/P0001 ,
		_w13211_,
		_w13212_
	);
	LUT2 #(
		.INIT('h2)
	) name12681 (
		_w13207_,
		_w13208_,
		_w13213_
	);
	LUT2 #(
		.INIT('h4)
	) name12682 (
		_w13212_,
		_w13213_,
		_w13214_
	);
	LUT2 #(
		.INIT('h2)
	) name12683 (
		\sa22_reg[1]/P0001 ,
		_w13214_,
		_w13215_
	);
	LUT2 #(
		.INIT('h1)
	) name12684 (
		_w13192_,
		_w13196_,
		_w13216_
	);
	LUT2 #(
		.INIT('h4)
	) name12685 (
		_w13205_,
		_w13216_,
		_w13217_
	);
	LUT2 #(
		.INIT('h4)
	) name12686 (
		_w13215_,
		_w13217_,
		_w13218_
	);
	LUT2 #(
		.INIT('h2)
	) name12687 (
		\sa22_reg[0]/P0001 ,
		_w13218_,
		_w13219_
	);
	LUT2 #(
		.INIT('h8)
	) name12688 (
		\sa22_reg[4]/P0001 ,
		_w12249_,
		_w13220_
	);
	LUT2 #(
		.INIT('h1)
	) name12689 (
		_w12395_,
		_w13220_,
		_w13221_
	);
	LUT2 #(
		.INIT('h2)
	) name12690 (
		_w12322_,
		_w13221_,
		_w13222_
	);
	LUT2 #(
		.INIT('h8)
	) name12691 (
		_w12295_,
		_w12779_,
		_w13223_
	);
	LUT2 #(
		.INIT('h2)
	) name12692 (
		\sa22_reg[1]/P0001 ,
		_w12384_,
		_w13224_
	);
	LUT2 #(
		.INIT('h4)
	) name12693 (
		_w13223_,
		_w13224_,
		_w13225_
	);
	LUT2 #(
		.INIT('h4)
	) name12694 (
		_w13222_,
		_w13225_,
		_w13226_
	);
	LUT2 #(
		.INIT('h4)
	) name12695 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		_w13227_
	);
	LUT2 #(
		.INIT('h8)
	) name12696 (
		_w12297_,
		_w13227_,
		_w13228_
	);
	LUT2 #(
		.INIT('h8)
	) name12697 (
		_w12291_,
		_w12303_,
		_w13229_
	);
	LUT2 #(
		.INIT('h8)
	) name12698 (
		\sa22_reg[4]/P0001 ,
		_w12259_,
		_w13230_
	);
	LUT2 #(
		.INIT('h4)
	) name12699 (
		\sa22_reg[6]/NET0131 ,
		_w12258_,
		_w13231_
	);
	LUT2 #(
		.INIT('h1)
	) name12700 (
		_w12321_,
		_w13231_,
		_w13232_
	);
	LUT2 #(
		.INIT('h1)
	) name12701 (
		\sa22_reg[4]/P0001 ,
		_w13232_,
		_w13233_
	);
	LUT2 #(
		.INIT('h1)
	) name12702 (
		\sa22_reg[1]/P0001 ,
		_w13228_,
		_w13234_
	);
	LUT2 #(
		.INIT('h4)
	) name12703 (
		_w13229_,
		_w13234_,
		_w13235_
	);
	LUT2 #(
		.INIT('h1)
	) name12704 (
		_w12723_,
		_w13230_,
		_w13236_
	);
	LUT2 #(
		.INIT('h8)
	) name12705 (
		_w13235_,
		_w13236_,
		_w13237_
	);
	LUT2 #(
		.INIT('h4)
	) name12706 (
		_w13233_,
		_w13237_,
		_w13238_
	);
	LUT2 #(
		.INIT('h1)
	) name12707 (
		_w13226_,
		_w13238_,
		_w13239_
	);
	LUT2 #(
		.INIT('h8)
	) name12708 (
		\sa22_reg[4]/P0001 ,
		_w12234_,
		_w13240_
	);
	LUT2 #(
		.INIT('h1)
	) name12709 (
		_w12716_,
		_w13240_,
		_w13241_
	);
	LUT2 #(
		.INIT('h1)
	) name12710 (
		_w12260_,
		_w13241_,
		_w13242_
	);
	LUT2 #(
		.INIT('h4)
	) name12711 (
		_w12393_,
		_w12791_,
		_w13243_
	);
	LUT2 #(
		.INIT('h4)
	) name12712 (
		_w13242_,
		_w13243_,
		_w13244_
	);
	LUT2 #(
		.INIT('h4)
	) name12713 (
		\sa22_reg[3]/P0001 ,
		_w12295_,
		_w13245_
	);
	LUT2 #(
		.INIT('h2)
	) name12714 (
		\sa22_reg[2]/P0001 ,
		_w13230_,
		_w13246_
	);
	LUT2 #(
		.INIT('h4)
	) name12715 (
		_w13245_,
		_w13246_,
		_w13247_
	);
	LUT2 #(
		.INIT('h1)
	) name12716 (
		_w13244_,
		_w13247_,
		_w13248_
	);
	LUT2 #(
		.INIT('h1)
	) name12717 (
		_w13239_,
		_w13248_,
		_w13249_
	);
	LUT2 #(
		.INIT('h1)
	) name12718 (
		\sa22_reg[0]/P0001 ,
		_w13249_,
		_w13250_
	);
	LUT2 #(
		.INIT('h8)
	) name12719 (
		\sa22_reg[4]/P0001 ,
		_w13197_,
		_w13251_
	);
	LUT2 #(
		.INIT('h4)
	) name12720 (
		\sa22_reg[6]/NET0131 ,
		_w12250_,
		_w13252_
	);
	LUT2 #(
		.INIT('h1)
	) name12721 (
		_w12298_,
		_w13251_,
		_w13253_
	);
	LUT2 #(
		.INIT('h4)
	) name12722 (
		_w13252_,
		_w13253_,
		_w13254_
	);
	LUT2 #(
		.INIT('h1)
	) name12723 (
		\sa22_reg[2]/P0001 ,
		_w13254_,
		_w13255_
	);
	LUT2 #(
		.INIT('h8)
	) name12724 (
		_w12301_,
		_w12735_,
		_w13256_
	);
	LUT2 #(
		.INIT('h8)
	) name12725 (
		_w12263_,
		_w12297_,
		_w13257_
	);
	LUT2 #(
		.INIT('h8)
	) name12726 (
		_w12282_,
		_w12319_,
		_w13258_
	);
	LUT2 #(
		.INIT('h1)
	) name12727 (
		_w12240_,
		_w13257_,
		_w13259_
	);
	LUT2 #(
		.INIT('h4)
	) name12728 (
		_w13256_,
		_w13259_,
		_w13260_
	);
	LUT2 #(
		.INIT('h4)
	) name12729 (
		_w13258_,
		_w13260_,
		_w13261_
	);
	LUT2 #(
		.INIT('h4)
	) name12730 (
		_w13255_,
		_w13261_,
		_w13262_
	);
	LUT2 #(
		.INIT('h1)
	) name12731 (
		\sa22_reg[1]/P0001 ,
		_w13262_,
		_w13263_
	);
	LUT2 #(
		.INIT('h8)
	) name12732 (
		\sa22_reg[1]/P0001 ,
		\sa22_reg[2]/P0001 ,
		_w13264_
	);
	LUT2 #(
		.INIT('h4)
	) name12733 (
		\sa22_reg[3]/P0001 ,
		_w12300_,
		_w13265_
	);
	LUT2 #(
		.INIT('h1)
	) name12734 (
		_w13252_,
		_w13265_,
		_w13266_
	);
	LUT2 #(
		.INIT('h1)
	) name12735 (
		\sa22_reg[4]/P0001 ,
		_w13266_,
		_w13267_
	);
	LUT2 #(
		.INIT('h8)
	) name12736 (
		\sa22_reg[4]/P0001 ,
		_w12300_,
		_w13268_
	);
	LUT2 #(
		.INIT('h4)
	) name12737 (
		\sa22_reg[5]/P0001 ,
		_w13268_,
		_w13269_
	);
	LUT2 #(
		.INIT('h1)
	) name12738 (
		_w13267_,
		_w13269_,
		_w13270_
	);
	LUT2 #(
		.INIT('h2)
	) name12739 (
		_w13264_,
		_w13270_,
		_w13271_
	);
	LUT2 #(
		.INIT('h8)
	) name12740 (
		_w12298_,
		_w13227_,
		_w13272_
	);
	LUT2 #(
		.INIT('h8)
	) name12741 (
		_w12738_,
		_w13227_,
		_w13273_
	);
	LUT2 #(
		.INIT('h8)
	) name12742 (
		\sa22_reg[1]/P0001 ,
		_w13273_,
		_w13274_
	);
	LUT2 #(
		.INIT('h8)
	) name12743 (
		_w12260_,
		_w13197_,
		_w13275_
	);
	LUT2 #(
		.INIT('h8)
	) name12744 (
		\sa22_reg[2]/P0001 ,
		_w13275_,
		_w13276_
	);
	LUT2 #(
		.INIT('h1)
	) name12745 (
		_w12280_,
		_w13272_,
		_w13277_
	);
	LUT2 #(
		.INIT('h4)
	) name12746 (
		_w12717_,
		_w13277_,
		_w13278_
	);
	LUT2 #(
		.INIT('h1)
	) name12747 (
		_w13274_,
		_w13276_,
		_w13279_
	);
	LUT2 #(
		.INIT('h8)
	) name12748 (
		_w13278_,
		_w13279_,
		_w13280_
	);
	LUT2 #(
		.INIT('h4)
	) name12749 (
		_w13271_,
		_w13280_,
		_w13281_
	);
	LUT2 #(
		.INIT('h4)
	) name12750 (
		_w13263_,
		_w13281_,
		_w13282_
	);
	LUT2 #(
		.INIT('h4)
	) name12751 (
		_w13250_,
		_w13282_,
		_w13283_
	);
	LUT2 #(
		.INIT('h4)
	) name12752 (
		_w13219_,
		_w13283_,
		_w13284_
	);
	LUT2 #(
		.INIT('h2)
	) name12753 (
		\u0_w_reg[0][6]/P0001 ,
		_w13284_,
		_w13285_
	);
	LUT2 #(
		.INIT('h4)
	) name12754 (
		\u0_w_reg[0][6]/P0001 ,
		_w13284_,
		_w13286_
	);
	LUT2 #(
		.INIT('h1)
	) name12755 (
		_w13285_,
		_w13286_,
		_w13287_
	);
	LUT2 #(
		.INIT('h8)
	) name12756 (
		_w12580_,
		_w13287_,
		_w13288_
	);
	LUT2 #(
		.INIT('h1)
	) name12757 (
		_w12580_,
		_w13287_,
		_w13289_
	);
	LUT2 #(
		.INIT('h1)
	) name12758 (
		_w13288_,
		_w13289_,
		_w13290_
	);
	LUT2 #(
		.INIT('h4)
	) name12759 (
		_w13189_,
		_w13290_,
		_w13291_
	);
	LUT2 #(
		.INIT('h2)
	) name12760 (
		_w13189_,
		_w13290_,
		_w13292_
	);
	LUT2 #(
		.INIT('h1)
	) name12761 (
		\ld_r_reg/P0001 ,
		_w13291_,
		_w13293_
	);
	LUT2 #(
		.INIT('h4)
	) name12762 (
		_w13292_,
		_w13293_,
		_w13294_
	);
	LUT2 #(
		.INIT('h1)
	) name12763 (
		\text_in_r_reg[102]/P0001 ,
		\u0_w_reg[0][6]/P0001 ,
		_w13295_
	);
	LUT2 #(
		.INIT('h8)
	) name12764 (
		\text_in_r_reg[102]/P0001 ,
		\u0_w_reg[0][6]/P0001 ,
		_w13296_
	);
	LUT2 #(
		.INIT('h2)
	) name12765 (
		\ld_r_reg/P0001 ,
		_w13295_,
		_w13297_
	);
	LUT2 #(
		.INIT('h4)
	) name12766 (
		_w13296_,
		_w13297_,
		_w13298_
	);
	LUT2 #(
		.INIT('h1)
	) name12767 (
		_w13294_,
		_w13298_,
		_w13299_
	);
	LUT2 #(
		.INIT('h2)
	) name12768 (
		\sa22_reg[5]/P0001 ,
		_w12266_,
		_w13300_
	);
	LUT2 #(
		.INIT('h2)
	) name12769 (
		_w12303_,
		_w13300_,
		_w13301_
	);
	LUT2 #(
		.INIT('h8)
	) name12770 (
		_w12773_,
		_w13200_,
		_w13302_
	);
	LUT2 #(
		.INIT('h8)
	) name12771 (
		_w12238_,
		_w12349_,
		_w13303_
	);
	LUT2 #(
		.INIT('h4)
	) name12772 (
		\sa22_reg[5]/P0001 ,
		_w13265_,
		_w13304_
	);
	LUT2 #(
		.INIT('h1)
	) name12773 (
		_w12253_,
		_w12345_,
		_w13305_
	);
	LUT2 #(
		.INIT('h4)
	) name12774 (
		_w13304_,
		_w13305_,
		_w13306_
	);
	LUT2 #(
		.INIT('h2)
	) name12775 (
		\sa22_reg[2]/P0001 ,
		_w13306_,
		_w13307_
	);
	LUT2 #(
		.INIT('h1)
	) name12776 (
		_w13301_,
		_w13303_,
		_w13308_
	);
	LUT2 #(
		.INIT('h4)
	) name12777 (
		_w13302_,
		_w13308_,
		_w13309_
	);
	LUT2 #(
		.INIT('h4)
	) name12778 (
		_w13307_,
		_w13309_,
		_w13310_
	);
	LUT2 #(
		.INIT('h1)
	) name12779 (
		\sa22_reg[1]/P0001 ,
		_w13310_,
		_w13311_
	);
	LUT2 #(
		.INIT('h1)
	) name12780 (
		\sa22_reg[2]/P0001 ,
		_w12245_,
		_w13312_
	);
	LUT2 #(
		.INIT('h4)
	) name12781 (
		_w12715_,
		_w13312_,
		_w13313_
	);
	LUT2 #(
		.INIT('h1)
	) name12782 (
		_w13251_,
		_w13313_,
		_w13314_
	);
	LUT2 #(
		.INIT('h2)
	) name12783 (
		\sa22_reg[1]/P0001 ,
		_w13314_,
		_w13315_
	);
	LUT2 #(
		.INIT('h8)
	) name12784 (
		_w12244_,
		_w12349_,
		_w13316_
	);
	LUT2 #(
		.INIT('h1)
	) name12785 (
		_w12303_,
		_w12319_,
		_w13317_
	);
	LUT2 #(
		.INIT('h1)
	) name12786 (
		_w12755_,
		_w13317_,
		_w13318_
	);
	LUT2 #(
		.INIT('h1)
	) name12787 (
		\sa22_reg[2]/P0001 ,
		_w12721_,
		_w13319_
	);
	LUT2 #(
		.INIT('h4)
	) name12788 (
		_w13316_,
		_w13319_,
		_w13320_
	);
	LUT2 #(
		.INIT('h4)
	) name12789 (
		_w13318_,
		_w13320_,
		_w13321_
	);
	LUT2 #(
		.INIT('h2)
	) name12790 (
		\sa22_reg[2]/P0001 ,
		_w12756_,
		_w13322_
	);
	LUT2 #(
		.INIT('h4)
	) name12791 (
		_w12331_,
		_w13322_,
		_w13323_
	);
	LUT2 #(
		.INIT('h8)
	) name12792 (
		_w13207_,
		_w13323_,
		_w13324_
	);
	LUT2 #(
		.INIT('h1)
	) name12793 (
		_w13321_,
		_w13324_,
		_w13325_
	);
	LUT2 #(
		.INIT('h1)
	) name12794 (
		_w12724_,
		_w12747_,
		_w13326_
	);
	LUT2 #(
		.INIT('h4)
	) name12795 (
		_w13315_,
		_w13326_,
		_w13327_
	);
	LUT2 #(
		.INIT('h4)
	) name12796 (
		_w13325_,
		_w13327_,
		_w13328_
	);
	LUT2 #(
		.INIT('h4)
	) name12797 (
		_w13311_,
		_w13328_,
		_w13329_
	);
	LUT2 #(
		.INIT('h2)
	) name12798 (
		\sa22_reg[0]/P0001 ,
		_w13329_,
		_w13330_
	);
	LUT2 #(
		.INIT('h8)
	) name12799 (
		_w12282_,
		_w12747_,
		_w13331_
	);
	LUT2 #(
		.INIT('h1)
	) name12800 (
		_w12347_,
		_w12795_,
		_w13332_
	);
	LUT2 #(
		.INIT('h1)
	) name12801 (
		\sa22_reg[3]/P0001 ,
		_w13332_,
		_w13333_
	);
	LUT2 #(
		.INIT('h2)
	) name12802 (
		_w12781_,
		_w13333_,
		_w13334_
	);
	LUT2 #(
		.INIT('h1)
	) name12803 (
		_w12300_,
		_w12811_,
		_w13335_
	);
	LUT2 #(
		.INIT('h1)
	) name12804 (
		_w12263_,
		_w13335_,
		_w13336_
	);
	LUT2 #(
		.INIT('h8)
	) name12805 (
		_w12321_,
		_w12735_,
		_w13337_
	);
	LUT2 #(
		.INIT('h8)
	) name12806 (
		_w12291_,
		_w13200_,
		_w13338_
	);
	LUT2 #(
		.INIT('h2)
	) name12807 (
		\sa22_reg[1]/P0001 ,
		_w12301_,
		_w13339_
	);
	LUT2 #(
		.INIT('h4)
	) name12808 (
		_w13338_,
		_w13339_,
		_w13340_
	);
	LUT2 #(
		.INIT('h4)
	) name12809 (
		_w13337_,
		_w13340_,
		_w13341_
	);
	LUT2 #(
		.INIT('h4)
	) name12810 (
		_w13336_,
		_w13341_,
		_w13342_
	);
	LUT2 #(
		.INIT('h1)
	) name12811 (
		_w13334_,
		_w13342_,
		_w13343_
	);
	LUT2 #(
		.INIT('h4)
	) name12812 (
		\sa22_reg[1]/P0001 ,
		_w12249_,
		_w13344_
	);
	LUT2 #(
		.INIT('h4)
	) name12813 (
		_w12732_,
		_w13344_,
		_w13345_
	);
	LUT2 #(
		.INIT('h1)
	) name12814 (
		_w12257_,
		_w12332_,
		_w13346_
	);
	LUT2 #(
		.INIT('h2)
	) name12815 (
		_w12303_,
		_w13346_,
		_w13347_
	);
	LUT2 #(
		.INIT('h2)
	) name12816 (
		\sa22_reg[2]/P0001 ,
		_w13345_,
		_w13348_
	);
	LUT2 #(
		.INIT('h4)
	) name12817 (
		_w13347_,
		_w13348_,
		_w13349_
	);
	LUT2 #(
		.INIT('h8)
	) name12818 (
		_w12249_,
		_w12732_,
		_w13350_
	);
	LUT2 #(
		.INIT('h1)
	) name12819 (
		_w12331_,
		_w13350_,
		_w13351_
	);
	LUT2 #(
		.INIT('h1)
	) name12820 (
		\sa22_reg[2]/P0001 ,
		_w13245_,
		_w13352_
	);
	LUT2 #(
		.INIT('h8)
	) name12821 (
		_w13351_,
		_w13352_,
		_w13353_
	);
	LUT2 #(
		.INIT('h1)
	) name12822 (
		_w13349_,
		_w13353_,
		_w13354_
	);
	LUT2 #(
		.INIT('h1)
	) name12823 (
		_w13343_,
		_w13354_,
		_w13355_
	);
	LUT2 #(
		.INIT('h1)
	) name12824 (
		\sa22_reg[0]/P0001 ,
		_w13355_,
		_w13356_
	);
	LUT2 #(
		.INIT('h8)
	) name12825 (
		\sa22_reg[6]/NET0131 ,
		_w13228_,
		_w13357_
	);
	LUT2 #(
		.INIT('h8)
	) name12826 (
		_w12244_,
		_w12249_,
		_w13358_
	);
	LUT2 #(
		.INIT('h4)
	) name12827 (
		\sa22_reg[2]/P0001 ,
		_w13358_,
		_w13359_
	);
	LUT2 #(
		.INIT('h8)
	) name12828 (
		_w12244_,
		_w13197_,
		_w13360_
	);
	LUT2 #(
		.INIT('h1)
	) name12829 (
		_w12324_,
		_w13360_,
		_w13361_
	);
	LUT2 #(
		.INIT('h2)
	) name12830 (
		\sa22_reg[2]/P0001 ,
		_w13361_,
		_w13362_
	);
	LUT2 #(
		.INIT('h1)
	) name12831 (
		_w12717_,
		_w13359_,
		_w13363_
	);
	LUT2 #(
		.INIT('h8)
	) name12832 (
		_w12770_,
		_w13363_,
		_w13364_
	);
	LUT2 #(
		.INIT('h4)
	) name12833 (
		_w13362_,
		_w13364_,
		_w13365_
	);
	LUT2 #(
		.INIT('h4)
	) name12834 (
		_w12240_,
		_w12810_,
		_w13366_
	);
	LUT2 #(
		.INIT('h1)
	) name12835 (
		\sa22_reg[2]/P0001 ,
		_w12343_,
		_w13367_
	);
	LUT2 #(
		.INIT('h4)
	) name12836 (
		\sa22_reg[3]/P0001 ,
		_w12251_,
		_w13368_
	);
	LUT2 #(
		.INIT('h4)
	) name12837 (
		_w12267_,
		_w13368_,
		_w13369_
	);
	LUT2 #(
		.INIT('h1)
	) name12838 (
		_w12802_,
		_w13369_,
		_w13370_
	);
	LUT2 #(
		.INIT('h8)
	) name12839 (
		_w13367_,
		_w13370_,
		_w13371_
	);
	LUT2 #(
		.INIT('h1)
	) name12840 (
		_w13366_,
		_w13371_,
		_w13372_
	);
	LUT2 #(
		.INIT('h1)
	) name12841 (
		\sa22_reg[1]/P0001 ,
		_w12382_,
		_w13373_
	);
	LUT2 #(
		.INIT('h4)
	) name12842 (
		_w13372_,
		_w13373_,
		_w13374_
	);
	LUT2 #(
		.INIT('h1)
	) name12843 (
		_w13365_,
		_w13374_,
		_w13375_
	);
	LUT2 #(
		.INIT('h1)
	) name12844 (
		_w13331_,
		_w13357_,
		_w13376_
	);
	LUT2 #(
		.INIT('h4)
	) name12845 (
		_w13375_,
		_w13376_,
		_w13377_
	);
	LUT2 #(
		.INIT('h4)
	) name12846 (
		_w13356_,
		_w13377_,
		_w13378_
	);
	LUT2 #(
		.INIT('h4)
	) name12847 (
		_w13330_,
		_w13378_,
		_w13379_
	);
	LUT2 #(
		.INIT('h1)
	) name12848 (
		_w11802_,
		_w13109_,
		_w13380_
	);
	LUT2 #(
		.INIT('h8)
	) name12849 (
		_w12178_,
		_w13380_,
		_w13381_
	);
	LUT2 #(
		.INIT('h2)
	) name12850 (
		\sa11_reg[2]/P0001 ,
		_w13381_,
		_w13382_
	);
	LUT2 #(
		.INIT('h1)
	) name12851 (
		_w11816_,
		_w13092_,
		_w13383_
	);
	LUT2 #(
		.INIT('h2)
	) name12852 (
		\sa11_reg[3]/P0001 ,
		_w13383_,
		_w13384_
	);
	LUT2 #(
		.INIT('h1)
	) name12853 (
		_w12185_,
		_w13126_,
		_w13385_
	);
	LUT2 #(
		.INIT('h4)
	) name12854 (
		_w13384_,
		_w13385_,
		_w13386_
	);
	LUT2 #(
		.INIT('h1)
	) name12855 (
		\sa11_reg[2]/P0001 ,
		_w13386_,
		_w13387_
	);
	LUT2 #(
		.INIT('h4)
	) name12856 (
		\sa11_reg[2]/P0001 ,
		_w11833_,
		_w13388_
	);
	LUT2 #(
		.INIT('h4)
	) name12857 (
		\sa11_reg[5]/P0001 ,
		_w11829_,
		_w13389_
	);
	LUT2 #(
		.INIT('h4)
	) name12858 (
		\sa11_reg[2]/P0001 ,
		_w13389_,
		_w13390_
	);
	LUT2 #(
		.INIT('h1)
	) name12859 (
		_w13159_,
		_w13388_,
		_w13391_
	);
	LUT2 #(
		.INIT('h4)
	) name12860 (
		_w13390_,
		_w13391_,
		_w13392_
	);
	LUT2 #(
		.INIT('h2)
	) name12861 (
		\sa11_reg[1]/P0001 ,
		_w13392_,
		_w13393_
	);
	LUT2 #(
		.INIT('h4)
	) name12862 (
		\sa11_reg[5]/P0001 ,
		_w13139_,
		_w13394_
	);
	LUT2 #(
		.INIT('h8)
	) name12863 (
		_w11823_,
		_w13394_,
		_w13395_
	);
	LUT2 #(
		.INIT('h2)
	) name12864 (
		\sa11_reg[5]/P0001 ,
		_w11870_,
		_w13396_
	);
	LUT2 #(
		.INIT('h2)
	) name12865 (
		_w11796_,
		_w13396_,
		_w13397_
	);
	LUT2 #(
		.INIT('h4)
	) name12866 (
		\sa11_reg[3]/P0001 ,
		_w13389_,
		_w13398_
	);
	LUT2 #(
		.INIT('h1)
	) name12867 (
		_w12129_,
		_w12223_,
		_w13399_
	);
	LUT2 #(
		.INIT('h4)
	) name12868 (
		_w13398_,
		_w13399_,
		_w13400_
	);
	LUT2 #(
		.INIT('h2)
	) name12869 (
		\sa11_reg[2]/P0001 ,
		_w13400_,
		_w13401_
	);
	LUT2 #(
		.INIT('h1)
	) name12870 (
		_w11942_,
		_w13397_,
		_w13402_
	);
	LUT2 #(
		.INIT('h4)
	) name12871 (
		_w13395_,
		_w13402_,
		_w13403_
	);
	LUT2 #(
		.INIT('h4)
	) name12872 (
		_w13401_,
		_w13403_,
		_w13404_
	);
	LUT2 #(
		.INIT('h1)
	) name12873 (
		\sa11_reg[1]/P0001 ,
		_w13404_,
		_w13405_
	);
	LUT2 #(
		.INIT('h1)
	) name12874 (
		_w11836_,
		_w11872_,
		_w13406_
	);
	LUT2 #(
		.INIT('h4)
	) name12875 (
		_w13387_,
		_w13406_,
		_w13407_
	);
	LUT2 #(
		.INIT('h4)
	) name12876 (
		_w13382_,
		_w13407_,
		_w13408_
	);
	LUT2 #(
		.INIT('h4)
	) name12877 (
		_w13393_,
		_w13408_,
		_w13409_
	);
	LUT2 #(
		.INIT('h4)
	) name12878 (
		_w13405_,
		_w13409_,
		_w13410_
	);
	LUT2 #(
		.INIT('h2)
	) name12879 (
		\sa11_reg[0]/P0001 ,
		_w13410_,
		_w13411_
	);
	LUT2 #(
		.INIT('h8)
	) name12880 (
		\sa11_reg[3]/P0001 ,
		_w11793_,
		_w13412_
	);
	LUT2 #(
		.INIT('h8)
	) name12881 (
		\sa11_reg[4]/P0001 ,
		_w11858_,
		_w13413_
	);
	LUT2 #(
		.INIT('h1)
	) name12882 (
		_w13107_,
		_w13413_,
		_w13414_
	);
	LUT2 #(
		.INIT('h2)
	) name12883 (
		\sa11_reg[7]/NET0131 ,
		_w13414_,
		_w13415_
	);
	LUT2 #(
		.INIT('h4)
	) name12884 (
		_w11794_,
		_w11829_,
		_w13416_
	);
	LUT2 #(
		.INIT('h1)
	) name12885 (
		_w13412_,
		_w13416_,
		_w13417_
	);
	LUT2 #(
		.INIT('h4)
	) name12886 (
		_w13415_,
		_w13417_,
		_w13418_
	);
	LUT2 #(
		.INIT('h2)
	) name12887 (
		\sa11_reg[1]/P0001 ,
		_w13418_,
		_w13419_
	);
	LUT2 #(
		.INIT('h8)
	) name12888 (
		\sa11_reg[6]/NET0131 ,
		_w12126_,
		_w13420_
	);
	LUT2 #(
		.INIT('h1)
	) name12889 (
		_w12176_,
		_w13420_,
		_w13421_
	);
	LUT2 #(
		.INIT('h4)
	) name12890 (
		_w13133_,
		_w13421_,
		_w13422_
	);
	LUT2 #(
		.INIT('h1)
	) name12891 (
		\sa11_reg[2]/P0001 ,
		_w13422_,
		_w13423_
	);
	LUT2 #(
		.INIT('h1)
	) name12892 (
		_w11816_,
		_w11847_,
		_w13424_
	);
	LUT2 #(
		.INIT('h2)
	) name12893 (
		_w11796_,
		_w13424_,
		_w13425_
	);
	LUT2 #(
		.INIT('h1)
	) name12894 (
		\sa11_reg[1]/P0001 ,
		_w11858_,
		_w13426_
	);
	LUT2 #(
		.INIT('h8)
	) name12895 (
		_w11892_,
		_w13426_,
		_w13427_
	);
	LUT2 #(
		.INIT('h1)
	) name12896 (
		_w13425_,
		_w13427_,
		_w13428_
	);
	LUT2 #(
		.INIT('h2)
	) name12897 (
		\sa11_reg[2]/P0001 ,
		_w13428_,
		_w13429_
	);
	LUT2 #(
		.INIT('h1)
	) name12898 (
		_w11854_,
		_w11907_,
		_w13430_
	);
	LUT2 #(
		.INIT('h1)
	) name12899 (
		\sa11_reg[3]/P0001 ,
		_w13430_,
		_w13431_
	);
	LUT2 #(
		.INIT('h1)
	) name12900 (
		_w11902_,
		_w13431_,
		_w13432_
	);
	LUT2 #(
		.INIT('h1)
	) name12901 (
		\sa11_reg[1]/P0001 ,
		_w13432_,
		_w13433_
	);
	LUT2 #(
		.INIT('h1)
	) name12902 (
		_w13423_,
		_w13429_,
		_w13434_
	);
	LUT2 #(
		.INIT('h4)
	) name12903 (
		_w13433_,
		_w13434_,
		_w13435_
	);
	LUT2 #(
		.INIT('h4)
	) name12904 (
		_w13419_,
		_w13435_,
		_w13436_
	);
	LUT2 #(
		.INIT('h1)
	) name12905 (
		\sa11_reg[0]/P0001 ,
		_w13436_,
		_w13437_
	);
	LUT2 #(
		.INIT('h8)
	) name12906 (
		\sa11_reg[6]/NET0131 ,
		_w13137_,
		_w13438_
	);
	LUT2 #(
		.INIT('h8)
	) name12907 (
		_w11825_,
		_w12188_,
		_w13439_
	);
	LUT2 #(
		.INIT('h8)
	) name12908 (
		_w11853_,
		_w13439_,
		_w13440_
	);
	LUT2 #(
		.INIT('h1)
	) name12909 (
		_w11826_,
		_w12194_,
		_w13441_
	);
	LUT2 #(
		.INIT('h4)
	) name12910 (
		_w13100_,
		_w13441_,
		_w13442_
	);
	LUT2 #(
		.INIT('h2)
	) name12911 (
		_w13106_,
		_w13442_,
		_w13443_
	);
	LUT2 #(
		.INIT('h1)
	) name12912 (
		_w12205_,
		_w13440_,
		_w13444_
	);
	LUT2 #(
		.INIT('h4)
	) name12913 (
		_w13443_,
		_w13444_,
		_w13445_
	);
	LUT2 #(
		.INIT('h1)
	) name12914 (
		\sa11_reg[1]/P0001 ,
		_w13445_,
		_w13446_
	);
	LUT2 #(
		.INIT('h4)
	) name12915 (
		\sa11_reg[3]/P0001 ,
		_w12152_,
		_w13447_
	);
	LUT2 #(
		.INIT('h4)
	) name12916 (
		\sa11_reg[2]/P0001 ,
		_w13447_,
		_w13448_
	);
	LUT2 #(
		.INIT('h8)
	) name12917 (
		_w12194_,
		_w12206_,
		_w13449_
	);
	LUT2 #(
		.INIT('h8)
	) name12918 (
		_w11846_,
		_w11871_,
		_w13450_
	);
	LUT2 #(
		.INIT('h1)
	) name12919 (
		_w11866_,
		_w11881_,
		_w13451_
	);
	LUT2 #(
		.INIT('h1)
	) name12920 (
		_w13449_,
		_w13450_,
		_w13452_
	);
	LUT2 #(
		.INIT('h8)
	) name12921 (
		_w13451_,
		_w13452_,
		_w13453_
	);
	LUT2 #(
		.INIT('h4)
	) name12922 (
		_w13448_,
		_w13453_,
		_w13454_
	);
	LUT2 #(
		.INIT('h2)
	) name12923 (
		\sa11_reg[1]/P0001 ,
		_w13454_,
		_w13455_
	);
	LUT2 #(
		.INIT('h2)
	) name12924 (
		\sa11_reg[1]/P0001 ,
		_w12125_,
		_w13456_
	);
	LUT2 #(
		.INIT('h8)
	) name12925 (
		\sa11_reg[2]/P0001 ,
		_w11860_,
		_w13457_
	);
	LUT2 #(
		.INIT('h1)
	) name12926 (
		_w11833_,
		_w11871_,
		_w13458_
	);
	LUT2 #(
		.INIT('h2)
	) name12927 (
		_w13457_,
		_w13458_,
		_w13459_
	);
	LUT2 #(
		.INIT('h4)
	) name12928 (
		_w13456_,
		_w13459_,
		_w13460_
	);
	LUT2 #(
		.INIT('h1)
	) name12929 (
		_w13438_,
		_w13460_,
		_w13461_
	);
	LUT2 #(
		.INIT('h4)
	) name12930 (
		_w13446_,
		_w13461_,
		_w13462_
	);
	LUT2 #(
		.INIT('h4)
	) name12931 (
		_w13455_,
		_w13462_,
		_w13463_
	);
	LUT2 #(
		.INIT('h4)
	) name12932 (
		_w13411_,
		_w13463_,
		_w13464_
	);
	LUT2 #(
		.INIT('h4)
	) name12933 (
		_w13437_,
		_w13464_,
		_w13465_
	);
	LUT2 #(
		.INIT('h2)
	) name12934 (
		_w13379_,
		_w13465_,
		_w13466_
	);
	LUT2 #(
		.INIT('h4)
	) name12935 (
		_w13379_,
		_w13465_,
		_w13467_
	);
	LUT2 #(
		.INIT('h1)
	) name12936 (
		_w13466_,
		_w13467_,
		_w13468_
	);
	LUT2 #(
		.INIT('h1)
	) name12937 (
		_w13131_,
		_w13388_,
		_w13469_
	);
	LUT2 #(
		.INIT('h1)
	) name12938 (
		\sa11_reg[7]/NET0131 ,
		_w13469_,
		_w13470_
	);
	LUT2 #(
		.INIT('h4)
	) name12939 (
		_w11797_,
		_w11823_,
		_w13471_
	);
	LUT2 #(
		.INIT('h4)
	) name12940 (
		_w11822_,
		_w13471_,
		_w13472_
	);
	LUT2 #(
		.INIT('h8)
	) name12941 (
		_w11791_,
		_w13106_,
		_w13473_
	);
	LUT2 #(
		.INIT('h8)
	) name12942 (
		_w11801_,
		_w13457_,
		_w13474_
	);
	LUT2 #(
		.INIT('h1)
	) name12943 (
		_w11924_,
		_w13473_,
		_w13475_
	);
	LUT2 #(
		.INIT('h1)
	) name12944 (
		_w13472_,
		_w13474_,
		_w13476_
	);
	LUT2 #(
		.INIT('h8)
	) name12945 (
		_w13475_,
		_w13476_,
		_w13477_
	);
	LUT2 #(
		.INIT('h4)
	) name12946 (
		_w13470_,
		_w13477_,
		_w13478_
	);
	LUT2 #(
		.INIT('h1)
	) name12947 (
		\sa11_reg[1]/P0001 ,
		_w13478_,
		_w13479_
	);
	LUT2 #(
		.INIT('h8)
	) name12948 (
		_w13100_,
		_w13106_,
		_w13480_
	);
	LUT2 #(
		.INIT('h4)
	) name12949 (
		\sa11_reg[5]/P0001 ,
		_w11796_,
		_w13481_
	);
	LUT2 #(
		.INIT('h1)
	) name12950 (
		_w11861_,
		_w13481_,
		_w13482_
	);
	LUT2 #(
		.INIT('h2)
	) name12951 (
		\sa11_reg[6]/NET0131 ,
		_w13482_,
		_w13483_
	);
	LUT2 #(
		.INIT('h1)
	) name12952 (
		_w12115_,
		_w12129_,
		_w13484_
	);
	LUT2 #(
		.INIT('h4)
	) name12953 (
		_w13483_,
		_w13484_,
		_w13485_
	);
	LUT2 #(
		.INIT('h2)
	) name12954 (
		\sa11_reg[2]/P0001 ,
		_w13485_,
		_w13486_
	);
	LUT2 #(
		.INIT('h8)
	) name12955 (
		_w11870_,
		_w13107_,
		_w13487_
	);
	LUT2 #(
		.INIT('h8)
	) name12956 (
		\sa11_reg[3]/P0001 ,
		_w11791_,
		_w13488_
	);
	LUT2 #(
		.INIT('h8)
	) name12957 (
		\sa11_reg[4]/P0001 ,
		_w11876_,
		_w13489_
	);
	LUT2 #(
		.INIT('h1)
	) name12958 (
		_w11853_,
		_w12146_,
		_w13490_
	);
	LUT2 #(
		.INIT('h1)
	) name12959 (
		_w13488_,
		_w13489_,
		_w13491_
	);
	LUT2 #(
		.INIT('h8)
	) name12960 (
		_w13490_,
		_w13491_,
		_w13492_
	);
	LUT2 #(
		.INIT('h2)
	) name12961 (
		\sa11_reg[2]/P0001 ,
		_w13492_,
		_w13493_
	);
	LUT2 #(
		.INIT('h1)
	) name12962 (
		_w11859_,
		_w13487_,
		_w13494_
	);
	LUT2 #(
		.INIT('h4)
	) name12963 (
		_w13493_,
		_w13494_,
		_w13495_
	);
	LUT2 #(
		.INIT('h2)
	) name12964 (
		\sa11_reg[1]/P0001 ,
		_w13495_,
		_w13496_
	);
	LUT2 #(
		.INIT('h1)
	) name12965 (
		_w13126_,
		_w13480_,
		_w13497_
	);
	LUT2 #(
		.INIT('h4)
	) name12966 (
		_w13486_,
		_w13497_,
		_w13498_
	);
	LUT2 #(
		.INIT('h4)
	) name12967 (
		_w13479_,
		_w13498_,
		_w13499_
	);
	LUT2 #(
		.INIT('h4)
	) name12968 (
		_w13496_,
		_w13499_,
		_w13500_
	);
	LUT2 #(
		.INIT('h2)
	) name12969 (
		\sa11_reg[0]/P0001 ,
		_w13500_,
		_w13501_
	);
	LUT2 #(
		.INIT('h4)
	) name12970 (
		\sa11_reg[2]/P0001 ,
		_w11886_,
		_w13502_
	);
	LUT2 #(
		.INIT('h8)
	) name12971 (
		_w11806_,
		_w11846_,
		_w13503_
	);
	LUT2 #(
		.INIT('h1)
	) name12972 (
		\sa11_reg[1]/P0001 ,
		_w11832_,
		_w13504_
	);
	LUT2 #(
		.INIT('h1)
	) name12973 (
		_w13109_,
		_w13502_,
		_w13505_
	);
	LUT2 #(
		.INIT('h8)
	) name12974 (
		_w13504_,
		_w13505_,
		_w13506_
	);
	LUT2 #(
		.INIT('h4)
	) name12975 (
		_w13503_,
		_w13506_,
		_w13507_
	);
	LUT2 #(
		.INIT('h2)
	) name12976 (
		\sa11_reg[2]/P0001 ,
		_w11936_,
		_w13508_
	);
	LUT2 #(
		.INIT('h8)
	) name12977 (
		_w11791_,
		_w11863_,
		_w13509_
	);
	LUT2 #(
		.INIT('h1)
	) name12978 (
		\sa11_reg[2]/P0001 ,
		_w11900_,
		_w13510_
	);
	LUT2 #(
		.INIT('h4)
	) name12979 (
		_w13509_,
		_w13510_,
		_w13511_
	);
	LUT2 #(
		.INIT('h1)
	) name12980 (
		_w13508_,
		_w13511_,
		_w13512_
	);
	LUT2 #(
		.INIT('h8)
	) name12981 (
		\sa11_reg[3]/P0001 ,
		_w11798_,
		_w13513_
	);
	LUT2 #(
		.INIT('h2)
	) name12982 (
		\sa11_reg[1]/P0001 ,
		_w13132_,
		_w13514_
	);
	LUT2 #(
		.INIT('h4)
	) name12983 (
		_w13513_,
		_w13514_,
		_w13515_
	);
	LUT2 #(
		.INIT('h4)
	) name12984 (
		_w13512_,
		_w13515_,
		_w13516_
	);
	LUT2 #(
		.INIT('h1)
	) name12985 (
		_w13507_,
		_w13516_,
		_w13517_
	);
	LUT2 #(
		.INIT('h4)
	) name12986 (
		_w11791_,
		_w11794_,
		_w13518_
	);
	LUT2 #(
		.INIT('h8)
	) name12987 (
		_w13396_,
		_w13518_,
		_w13519_
	);
	LUT2 #(
		.INIT('h2)
	) name12988 (
		\sa11_reg[2]/P0001 ,
		_w12217_,
		_w13520_
	);
	LUT2 #(
		.INIT('h4)
	) name12989 (
		_w13519_,
		_w13520_,
		_w13521_
	);
	LUT2 #(
		.INIT('h4)
	) name12990 (
		\sa11_reg[3]/P0001 ,
		_w11933_,
		_w13522_
	);
	LUT2 #(
		.INIT('h1)
	) name12991 (
		_w11942_,
		_w13522_,
		_w13523_
	);
	LUT2 #(
		.INIT('h1)
	) name12992 (
		\sa11_reg[2]/P0001 ,
		_w11941_,
		_w13524_
	);
	LUT2 #(
		.INIT('h4)
	) name12993 (
		_w13172_,
		_w13523_,
		_w13525_
	);
	LUT2 #(
		.INIT('h8)
	) name12994 (
		_w13524_,
		_w13525_,
		_w13526_
	);
	LUT2 #(
		.INIT('h1)
	) name12995 (
		_w13521_,
		_w13526_,
		_w13527_
	);
	LUT2 #(
		.INIT('h1)
	) name12996 (
		_w13517_,
		_w13527_,
		_w13528_
	);
	LUT2 #(
		.INIT('h1)
	) name12997 (
		\sa11_reg[0]/P0001 ,
		_w13528_,
		_w13529_
	);
	LUT2 #(
		.INIT('h2)
	) name12998 (
		_w11797_,
		_w11886_,
		_w13530_
	);
	LUT2 #(
		.INIT('h2)
	) name12999 (
		_w13430_,
		_w13530_,
		_w13531_
	);
	LUT2 #(
		.INIT('h2)
	) name13000 (
		_w12188_,
		_w13531_,
		_w13532_
	);
	LUT2 #(
		.INIT('h8)
	) name13001 (
		\sa11_reg[7]/NET0131 ,
		_w11853_,
		_w13533_
	);
	LUT2 #(
		.INIT('h1)
	) name13002 (
		_w11826_,
		_w13533_,
		_w13534_
	);
	LUT2 #(
		.INIT('h4)
	) name13003 (
		_w11883_,
		_w13534_,
		_w13535_
	);
	LUT2 #(
		.INIT('h1)
	) name13004 (
		\sa11_reg[3]/P0001 ,
		_w13535_,
		_w13536_
	);
	LUT2 #(
		.INIT('h1)
	) name13005 (
		_w11925_,
		_w12139_,
		_w13537_
	);
	LUT2 #(
		.INIT('h4)
	) name13006 (
		_w13536_,
		_w13537_,
		_w13538_
	);
	LUT2 #(
		.INIT('h2)
	) name13007 (
		\sa11_reg[2]/P0001 ,
		_w13538_,
		_w13539_
	);
	LUT2 #(
		.INIT('h1)
	) name13008 (
		_w13532_,
		_w13539_,
		_w13540_
	);
	LUT2 #(
		.INIT('h2)
	) name13009 (
		\sa11_reg[1]/P0001 ,
		_w13540_,
		_w13541_
	);
	LUT2 #(
		.INIT('h1)
	) name13010 (
		_w11815_,
		_w12125_,
		_w13542_
	);
	LUT2 #(
		.INIT('h1)
	) name13011 (
		\sa11_reg[2]/P0001 ,
		_w13542_,
		_w13543_
	);
	LUT2 #(
		.INIT('h4)
	) name13012 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[2]/P0001 ,
		_w13544_
	);
	LUT2 #(
		.INIT('h8)
	) name13013 (
		\sa11_reg[5]/P0001 ,
		_w13131_,
		_w13545_
	);
	LUT2 #(
		.INIT('h1)
	) name13014 (
		_w11859_,
		_w12119_,
		_w13546_
	);
	LUT2 #(
		.INIT('h4)
	) name13015 (
		_w13545_,
		_w13546_,
		_w13547_
	);
	LUT2 #(
		.INIT('h2)
	) name13016 (
		_w13544_,
		_w13547_,
		_w13548_
	);
	LUT2 #(
		.INIT('h2)
	) name13017 (
		\sa11_reg[2]/P0001 ,
		_w13447_,
		_w13549_
	);
	LUT2 #(
		.INIT('h1)
	) name13018 (
		_w13138_,
		_w13447_,
		_w13550_
	);
	LUT2 #(
		.INIT('h8)
	) name13019 (
		_w13523_,
		_w13550_,
		_w13551_
	);
	LUT2 #(
		.INIT('h1)
	) name13020 (
		\sa11_reg[1]/P0001 ,
		_w13549_,
		_w13552_
	);
	LUT2 #(
		.INIT('h4)
	) name13021 (
		_w13551_,
		_w13552_,
		_w13553_
	);
	LUT2 #(
		.INIT('h1)
	) name13022 (
		_w13543_,
		_w13548_,
		_w13554_
	);
	LUT2 #(
		.INIT('h4)
	) name13023 (
		_w13553_,
		_w13554_,
		_w13555_
	);
	LUT2 #(
		.INIT('h4)
	) name13024 (
		_w13529_,
		_w13555_,
		_w13556_
	);
	LUT2 #(
		.INIT('h4)
	) name13025 (
		_w13541_,
		_w13556_,
		_w13557_
	);
	LUT2 #(
		.INIT('h4)
	) name13026 (
		_w13501_,
		_w13557_,
		_w13558_
	);
	LUT2 #(
		.INIT('h8)
	) name13027 (
		\sa00_reg[4]/P0001 ,
		_w12035_,
		_w13559_
	);
	LUT2 #(
		.INIT('h8)
	) name13028 (
		\sa00_reg[3]/P0001 ,
		_w13559_,
		_w13560_
	);
	LUT2 #(
		.INIT('h1)
	) name13029 (
		_w12629_,
		_w13042_,
		_w13561_
	);
	LUT2 #(
		.INIT('h4)
	) name13030 (
		_w13560_,
		_w13561_,
		_w13562_
	);
	LUT2 #(
		.INIT('h1)
	) name13031 (
		\sa00_reg[2]/P0001 ,
		_w13562_,
		_w13563_
	);
	LUT2 #(
		.INIT('h4)
	) name13032 (
		_w12611_,
		_w12653_,
		_w13564_
	);
	LUT2 #(
		.INIT('h4)
	) name13033 (
		_w13563_,
		_w13564_,
		_w13565_
	);
	LUT2 #(
		.INIT('h2)
	) name13034 (
		\sa00_reg[1]/P0001 ,
		_w13565_,
		_w13566_
	);
	LUT2 #(
		.INIT('h1)
	) name13035 (
		_w11957_,
		_w12007_,
		_w13567_
	);
	LUT2 #(
		.INIT('h2)
	) name13036 (
		_w12056_,
		_w13567_,
		_w13568_
	);
	LUT2 #(
		.INIT('h1)
	) name13037 (
		_w11980_,
		_w12600_,
		_w13569_
	);
	LUT2 #(
		.INIT('h2)
	) name13038 (
		_w11985_,
		_w13569_,
		_w13570_
	);
	LUT2 #(
		.INIT('h8)
	) name13039 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[2]/P0001 ,
		_w13571_
	);
	LUT2 #(
		.INIT('h4)
	) name13040 (
		\sa00_reg[3]/P0001 ,
		_w11996_,
		_w13572_
	);
	LUT2 #(
		.INIT('h1)
	) name13041 (
		_w12632_,
		_w13572_,
		_w13573_
	);
	LUT2 #(
		.INIT('h2)
	) name13042 (
		_w13571_,
		_w13573_,
		_w13574_
	);
	LUT2 #(
		.INIT('h4)
	) name13043 (
		\sa00_reg[3]/P0001 ,
		_w12651_,
		_w13575_
	);
	LUT2 #(
		.INIT('h1)
	) name13044 (
		_w12003_,
		_w13575_,
		_w13576_
	);
	LUT2 #(
		.INIT('h2)
	) name13045 (
		_w13015_,
		_w13576_,
		_w13577_
	);
	LUT2 #(
		.INIT('h1)
	) name13046 (
		_w12997_,
		_w13068_,
		_w13578_
	);
	LUT2 #(
		.INIT('h1)
	) name13047 (
		\sa00_reg[2]/P0001 ,
		_w13578_,
		_w13579_
	);
	LUT2 #(
		.INIT('h8)
	) name13048 (
		_w11979_,
		_w12064_,
		_w13580_
	);
	LUT2 #(
		.INIT('h8)
	) name13049 (
		\sa00_reg[4]/P0001 ,
		_w13580_,
		_w13581_
	);
	LUT2 #(
		.INIT('h1)
	) name13050 (
		_w12034_,
		_w13581_,
		_w13582_
	);
	LUT2 #(
		.INIT('h4)
	) name13051 (
		_w13579_,
		_w13582_,
		_w13583_
	);
	LUT2 #(
		.INIT('h1)
	) name13052 (
		\sa00_reg[1]/P0001 ,
		_w13583_,
		_w13584_
	);
	LUT2 #(
		.INIT('h1)
	) name13053 (
		_w12691_,
		_w12702_,
		_w13585_
	);
	LUT2 #(
		.INIT('h1)
	) name13054 (
		_w13568_,
		_w13570_,
		_w13586_
	);
	LUT2 #(
		.INIT('h8)
	) name13055 (
		_w13585_,
		_w13586_,
		_w13587_
	);
	LUT2 #(
		.INIT('h1)
	) name13056 (
		_w13574_,
		_w13577_,
		_w13588_
	);
	LUT2 #(
		.INIT('h8)
	) name13057 (
		_w13587_,
		_w13588_,
		_w13589_
	);
	LUT2 #(
		.INIT('h4)
	) name13058 (
		_w13566_,
		_w13589_,
		_w13590_
	);
	LUT2 #(
		.INIT('h4)
	) name13059 (
		_w13584_,
		_w13590_,
		_w13591_
	);
	LUT2 #(
		.INIT('h1)
	) name13060 (
		\sa00_reg[0]/P0001 ,
		_w13591_,
		_w13592_
	);
	LUT2 #(
		.INIT('h8)
	) name13061 (
		_w11982_,
		_w11996_,
		_w13593_
	);
	LUT2 #(
		.INIT('h1)
	) name13062 (
		_w12624_,
		_w13593_,
		_w13594_
	);
	LUT2 #(
		.INIT('h8)
	) name13063 (
		\sa00_reg[7]/NET0131 ,
		_w11979_,
		_w13595_
	);
	LUT2 #(
		.INIT('h1)
	) name13064 (
		_w12090_,
		_w13559_,
		_w13596_
	);
	LUT2 #(
		.INIT('h4)
	) name13065 (
		_w13595_,
		_w13596_,
		_w13597_
	);
	LUT2 #(
		.INIT('h2)
	) name13066 (
		\sa00_reg[2]/P0001 ,
		_w13597_,
		_w13598_
	);
	LUT2 #(
		.INIT('h2)
	) name13067 (
		_w13594_,
		_w13598_,
		_w13599_
	);
	LUT2 #(
		.INIT('h2)
	) name13068 (
		\sa00_reg[1]/P0001 ,
		_w13599_,
		_w13600_
	);
	LUT2 #(
		.INIT('h1)
	) name13069 (
		_w12693_,
		_w13044_,
		_w13601_
	);
	LUT2 #(
		.INIT('h2)
	) name13070 (
		_w11952_,
		_w13601_,
		_w13602_
	);
	LUT2 #(
		.INIT('h2)
	) name13071 (
		_w11982_,
		_w12002_,
		_w13603_
	);
	LUT2 #(
		.INIT('h4)
	) name13072 (
		_w12064_,
		_w13603_,
		_w13604_
	);
	LUT2 #(
		.INIT('h1)
	) name13073 (
		_w12066_,
		_w13604_,
		_w13605_
	);
	LUT2 #(
		.INIT('h4)
	) name13074 (
		_w13602_,
		_w13605_,
		_w13606_
	);
	LUT2 #(
		.INIT('h1)
	) name13075 (
		\sa00_reg[1]/P0001 ,
		_w13606_,
		_w13607_
	);
	LUT2 #(
		.INIT('h4)
	) name13076 (
		\sa00_reg[6]/NET0131 ,
		_w13031_,
		_w13608_
	);
	LUT2 #(
		.INIT('h8)
	) name13077 (
		\sa00_reg[2]/P0001 ,
		_w12033_,
		_w13609_
	);
	LUT2 #(
		.INIT('h8)
	) name13078 (
		\sa00_reg[4]/P0001 ,
		_w11967_,
		_w13610_
	);
	LUT2 #(
		.INIT('h1)
	) name13079 (
		_w12066_,
		_w13069_,
		_w13611_
	);
	LUT2 #(
		.INIT('h1)
	) name13080 (
		_w13575_,
		_w13610_,
		_w13612_
	);
	LUT2 #(
		.INIT('h8)
	) name13081 (
		_w13611_,
		_w13612_,
		_w13613_
	);
	LUT2 #(
		.INIT('h1)
	) name13082 (
		\sa00_reg[2]/P0001 ,
		_w13613_,
		_w13614_
	);
	LUT2 #(
		.INIT('h1)
	) name13083 (
		_w13037_,
		_w13608_,
		_w13615_
	);
	LUT2 #(
		.INIT('h4)
	) name13084 (
		_w13609_,
		_w13615_,
		_w13616_
	);
	LUT2 #(
		.INIT('h4)
	) name13085 (
		_w13607_,
		_w13616_,
		_w13617_
	);
	LUT2 #(
		.INIT('h4)
	) name13086 (
		_w13614_,
		_w13617_,
		_w13618_
	);
	LUT2 #(
		.INIT('h4)
	) name13087 (
		_w13600_,
		_w13618_,
		_w13619_
	);
	LUT2 #(
		.INIT('h2)
	) name13088 (
		\sa00_reg[0]/P0001 ,
		_w13619_,
		_w13620_
	);
	LUT2 #(
		.INIT('h1)
	) name13089 (
		_w12068_,
		_w12624_,
		_w13621_
	);
	LUT2 #(
		.INIT('h2)
	) name13090 (
		\sa00_reg[3]/P0001 ,
		_w13621_,
		_w13622_
	);
	LUT2 #(
		.INIT('h1)
	) name13091 (
		_w13037_,
		_w13622_,
		_w13623_
	);
	LUT2 #(
		.INIT('h2)
	) name13092 (
		_w13571_,
		_w13623_,
		_w13624_
	);
	LUT2 #(
		.INIT('h8)
	) name13093 (
		\sa00_reg[2]/P0001 ,
		_w12025_,
		_w13625_
	);
	LUT2 #(
		.INIT('h1)
	) name13094 (
		_w12630_,
		_w13625_,
		_w13626_
	);
	LUT2 #(
		.INIT('h2)
	) name13095 (
		_w12054_,
		_w13626_,
		_w13627_
	);
	LUT2 #(
		.INIT('h1)
	) name13096 (
		_w12659_,
		_w13627_,
		_w13628_
	);
	LUT2 #(
		.INIT('h4)
	) name13097 (
		\sa00_reg[3]/P0001 ,
		_w11975_,
		_w13629_
	);
	LUT2 #(
		.INIT('h4)
	) name13098 (
		_w11959_,
		_w13629_,
		_w13630_
	);
	LUT2 #(
		.INIT('h1)
	) name13099 (
		_w12611_,
		_w13006_,
		_w13631_
	);
	LUT2 #(
		.INIT('h4)
	) name13100 (
		_w13630_,
		_w13631_,
		_w13632_
	);
	LUT2 #(
		.INIT('h8)
	) name13101 (
		_w13626_,
		_w13632_,
		_w13633_
	);
	LUT2 #(
		.INIT('h1)
	) name13102 (
		_w13628_,
		_w13633_,
		_w13634_
	);
	LUT2 #(
		.INIT('h4)
	) name13103 (
		\sa00_reg[5]/P0001 ,
		_w13042_,
		_w13635_
	);
	LUT2 #(
		.INIT('h2)
	) name13104 (
		\sa00_reg[2]/P0001 ,
		_w12691_,
		_w13636_
	);
	LUT2 #(
		.INIT('h4)
	) name13105 (
		_w12647_,
		_w13636_,
		_w13637_
	);
	LUT2 #(
		.INIT('h4)
	) name13106 (
		_w13635_,
		_w13637_,
		_w13638_
	);
	LUT2 #(
		.INIT('h1)
	) name13107 (
		\sa00_reg[2]/P0001 ,
		_w13580_,
		_w13639_
	);
	LUT2 #(
		.INIT('h1)
	) name13108 (
		_w11958_,
		_w13012_,
		_w13640_
	);
	LUT2 #(
		.INIT('h8)
	) name13109 (
		_w13639_,
		_w13640_,
		_w13641_
	);
	LUT2 #(
		.INIT('h1)
	) name13110 (
		_w13638_,
		_w13641_,
		_w13642_
	);
	LUT2 #(
		.INIT('h1)
	) name13111 (
		_w12025_,
		_w12667_,
		_w13643_
	);
	LUT2 #(
		.INIT('h4)
	) name13112 (
		_w13642_,
		_w13643_,
		_w13644_
	);
	LUT2 #(
		.INIT('h1)
	) name13113 (
		\sa00_reg[1]/P0001 ,
		_w13644_,
		_w13645_
	);
	LUT2 #(
		.INIT('h1)
	) name13114 (
		_w13624_,
		_w13634_,
		_w13646_
	);
	LUT2 #(
		.INIT('h4)
	) name13115 (
		_w13645_,
		_w13646_,
		_w13647_
	);
	LUT2 #(
		.INIT('h4)
	) name13116 (
		_w13592_,
		_w13647_,
		_w13648_
	);
	LUT2 #(
		.INIT('h4)
	) name13117 (
		_w13620_,
		_w13648_,
		_w13649_
	);
	LUT2 #(
		.INIT('h2)
	) name13118 (
		_w13558_,
		_w13649_,
		_w13650_
	);
	LUT2 #(
		.INIT('h4)
	) name13119 (
		_w13558_,
		_w13649_,
		_w13651_
	);
	LUT2 #(
		.INIT('h1)
	) name13120 (
		_w13650_,
		_w13651_,
		_w13652_
	);
	LUT2 #(
		.INIT('h8)
	) name13121 (
		_w13468_,
		_w13652_,
		_w13653_
	);
	LUT2 #(
		.INIT('h1)
	) name13122 (
		_w13468_,
		_w13652_,
		_w13654_
	);
	LUT2 #(
		.INIT('h1)
	) name13123 (
		_w13653_,
		_w13654_,
		_w13655_
	);
	LUT2 #(
		.INIT('h2)
	) name13124 (
		_w12564_,
		_w12884_,
		_w13656_
	);
	LUT2 #(
		.INIT('h8)
	) name13125 (
		\sa33_reg[6]/P0001 ,
		_w12457_,
		_w13657_
	);
	LUT2 #(
		.INIT('h1)
	) name13126 (
		_w12446_,
		_w12877_,
		_w13658_
	);
	LUT2 #(
		.INIT('h2)
	) name13127 (
		\sa33_reg[7]/NET0131 ,
		_w13658_,
		_w13659_
	);
	LUT2 #(
		.INIT('h1)
	) name13128 (
		_w13657_,
		_w13659_,
		_w13660_
	);
	LUT2 #(
		.INIT('h2)
	) name13129 (
		\sa33_reg[2]/P0001 ,
		_w13660_,
		_w13661_
	);
	LUT2 #(
		.INIT('h8)
	) name13130 (
		_w12418_,
		_w12877_,
		_w13662_
	);
	LUT2 #(
		.INIT('h8)
	) name13131 (
		\sa33_reg[4]/P0001 ,
		_w13662_,
		_w13663_
	);
	LUT2 #(
		.INIT('h1)
	) name13132 (
		_w12462_,
		_w13663_,
		_w13664_
	);
	LUT2 #(
		.INIT('h4)
	) name13133 (
		_w13661_,
		_w13664_,
		_w13665_
	);
	LUT2 #(
		.INIT('h2)
	) name13134 (
		\sa33_reg[1]/P0001 ,
		_w13665_,
		_w13666_
	);
	LUT2 #(
		.INIT('h8)
	) name13135 (
		\sa33_reg[4]/P0001 ,
		_w12561_,
		_w13667_
	);
	LUT2 #(
		.INIT('h4)
	) name13136 (
		\sa33_reg[6]/P0001 ,
		_w12421_,
		_w13668_
	);
	LUT2 #(
		.INIT('h1)
	) name13137 (
		_w12906_,
		_w12927_,
		_w13669_
	);
	LUT2 #(
		.INIT('h1)
	) name13138 (
		_w13667_,
		_w13668_,
		_w13670_
	);
	LUT2 #(
		.INIT('h8)
	) name13139 (
		_w13669_,
		_w13670_,
		_w13671_
	);
	LUT2 #(
		.INIT('h1)
	) name13140 (
		\sa33_reg[2]/P0001 ,
		_w13671_,
		_w13672_
	);
	LUT2 #(
		.INIT('h8)
	) name13141 (
		_w12448_,
		_w12561_,
		_w13673_
	);
	LUT2 #(
		.INIT('h2)
	) name13142 (
		_w12432_,
		_w12855_,
		_w13674_
	);
	LUT2 #(
		.INIT('h8)
	) name13143 (
		_w12410_,
		_w12470_,
		_w13675_
	);
	LUT2 #(
		.INIT('h1)
	) name13144 (
		_w12511_,
		_w12906_,
		_w13676_
	);
	LUT2 #(
		.INIT('h4)
	) name13145 (
		_w13674_,
		_w13676_,
		_w13677_
	);
	LUT2 #(
		.INIT('h4)
	) name13146 (
		_w13675_,
		_w13677_,
		_w13678_
	);
	LUT2 #(
		.INIT('h1)
	) name13147 (
		\sa33_reg[1]/P0001 ,
		_w13678_,
		_w13679_
	);
	LUT2 #(
		.INIT('h1)
	) name13148 (
		_w13656_,
		_w13673_,
		_w13680_
	);
	LUT2 #(
		.INIT('h4)
	) name13149 (
		_w13672_,
		_w13680_,
		_w13681_
	);
	LUT2 #(
		.INIT('h4)
	) name13150 (
		_w13679_,
		_w13681_,
		_w13682_
	);
	LUT2 #(
		.INIT('h4)
	) name13151 (
		_w13666_,
		_w13682_,
		_w13683_
	);
	LUT2 #(
		.INIT('h2)
	) name13152 (
		\sa33_reg[0]/P0001 ,
		_w13683_,
		_w13684_
	);
	LUT2 #(
		.INIT('h8)
	) name13153 (
		\sa33_reg[4]/P0001 ,
		_w12418_,
		_w13685_
	);
	LUT2 #(
		.INIT('h4)
	) name13154 (
		\sa33_reg[3]/P0001 ,
		_w12481_,
		_w13686_
	);
	LUT2 #(
		.INIT('h1)
	) name13155 (
		_w13685_,
		_w13686_,
		_w13687_
	);
	LUT2 #(
		.INIT('h2)
	) name13156 (
		\sa33_reg[2]/P0001 ,
		_w13687_,
		_w13688_
	);
	LUT2 #(
		.INIT('h1)
	) name13157 (
		\sa33_reg[5]/P0001 ,
		_w12460_,
		_w13689_
	);
	LUT2 #(
		.INIT('h2)
	) name13158 (
		\sa33_reg[4]/P0001 ,
		_w12877_,
		_w13690_
	);
	LUT2 #(
		.INIT('h2)
	) name13159 (
		_w13689_,
		_w13690_,
		_w13691_
	);
	LUT2 #(
		.INIT('h1)
	) name13160 (
		_w12470_,
		_w13691_,
		_w13692_
	);
	LUT2 #(
		.INIT('h1)
	) name13161 (
		\sa33_reg[2]/P0001 ,
		_w13692_,
		_w13693_
	);
	LUT2 #(
		.INIT('h1)
	) name13162 (
		_w12428_,
		_w12532_,
		_w13694_
	);
	LUT2 #(
		.INIT('h4)
	) name13163 (
		_w13688_,
		_w13694_,
		_w13695_
	);
	LUT2 #(
		.INIT('h4)
	) name13164 (
		_w13693_,
		_w13695_,
		_w13696_
	);
	LUT2 #(
		.INIT('h2)
	) name13165 (
		\sa33_reg[1]/P0001 ,
		_w13696_,
		_w13697_
	);
	LUT2 #(
		.INIT('h8)
	) name13166 (
		_w12414_,
		_w12457_,
		_w13698_
	);
	LUT2 #(
		.INIT('h8)
	) name13167 (
		_w12521_,
		_w12551_,
		_w13699_
	);
	LUT2 #(
		.INIT('h1)
	) name13168 (
		_w13698_,
		_w13699_,
		_w13700_
	);
	LUT2 #(
		.INIT('h1)
	) name13169 (
		\sa33_reg[2]/P0001 ,
		_w13700_,
		_w13701_
	);
	LUT2 #(
		.INIT('h8)
	) name13170 (
		_w12472_,
		_w12499_,
		_w13702_
	);
	LUT2 #(
		.INIT('h8)
	) name13171 (
		_w12413_,
		_w12560_,
		_w13703_
	);
	LUT2 #(
		.INIT('h8)
	) name13172 (
		_w12458_,
		_w12877_,
		_w13704_
	);
	LUT2 #(
		.INIT('h1)
	) name13173 (
		_w12919_,
		_w13702_,
		_w13705_
	);
	LUT2 #(
		.INIT('h1)
	) name13174 (
		_w13703_,
		_w13704_,
		_w13706_
	);
	LUT2 #(
		.INIT('h8)
	) name13175 (
		_w13705_,
		_w13706_,
		_w13707_
	);
	LUT2 #(
		.INIT('h4)
	) name13176 (
		_w13701_,
		_w13707_,
		_w13708_
	);
	LUT2 #(
		.INIT('h1)
	) name13177 (
		\sa33_reg[1]/P0001 ,
		_w13708_,
		_w13709_
	);
	LUT2 #(
		.INIT('h1)
	) name13178 (
		_w12444_,
		_w12473_,
		_w13710_
	);
	LUT2 #(
		.INIT('h2)
	) name13179 (
		_w12472_,
		_w13710_,
		_w13711_
	);
	LUT2 #(
		.INIT('h1)
	) name13180 (
		_w12507_,
		_w12919_,
		_w13712_
	);
	LUT2 #(
		.INIT('h1)
	) name13181 (
		\sa33_reg[2]/P0001 ,
		_w13712_,
		_w13713_
	);
	LUT2 #(
		.INIT('h1)
	) name13182 (
		_w12549_,
		_w12563_,
		_w13714_
	);
	LUT2 #(
		.INIT('h4)
	) name13183 (
		_w13711_,
		_w13714_,
		_w13715_
	);
	LUT2 #(
		.INIT('h4)
	) name13184 (
		_w13713_,
		_w13715_,
		_w13716_
	);
	LUT2 #(
		.INIT('h4)
	) name13185 (
		_w13709_,
		_w13716_,
		_w13717_
	);
	LUT2 #(
		.INIT('h4)
	) name13186 (
		_w13697_,
		_w13717_,
		_w13718_
	);
	LUT2 #(
		.INIT('h1)
	) name13187 (
		\sa33_reg[0]/P0001 ,
		_w13718_,
		_w13719_
	);
	LUT2 #(
		.INIT('h8)
	) name13188 (
		_w12414_,
		_w12426_,
		_w13720_
	);
	LUT2 #(
		.INIT('h4)
	) name13189 (
		\sa33_reg[4]/P0001 ,
		_w12421_,
		_w13721_
	);
	LUT2 #(
		.INIT('h1)
	) name13190 (
		_w12508_,
		_w13720_,
		_w13722_
	);
	LUT2 #(
		.INIT('h4)
	) name13191 (
		_w13721_,
		_w13722_,
		_w13723_
	);
	LUT2 #(
		.INIT('h1)
	) name13192 (
		\sa33_reg[2]/P0001 ,
		_w13723_,
		_w13724_
	);
	LUT2 #(
		.INIT('h1)
	) name13193 (
		_w12512_,
		_w12914_,
		_w13725_
	);
	LUT2 #(
		.INIT('h4)
	) name13194 (
		_w13724_,
		_w13725_,
		_w13726_
	);
	LUT2 #(
		.INIT('h1)
	) name13195 (
		\sa33_reg[1]/P0001 ,
		_w13726_,
		_w13727_
	);
	LUT2 #(
		.INIT('h2)
	) name13196 (
		_w12430_,
		_w12467_,
		_w13728_
	);
	LUT2 #(
		.INIT('h4)
	) name13197 (
		_w12448_,
		_w12473_,
		_w13729_
	);
	LUT2 #(
		.INIT('h1)
	) name13198 (
		\sa33_reg[2]/P0001 ,
		_w12415_,
		_w13730_
	);
	LUT2 #(
		.INIT('h4)
	) name13199 (
		_w13728_,
		_w13730_,
		_w13731_
	);
	LUT2 #(
		.INIT('h4)
	) name13200 (
		_w13729_,
		_w13731_,
		_w13732_
	);
	LUT2 #(
		.INIT('h1)
	) name13201 (
		_w12462_,
		_w12932_,
		_w13733_
	);
	LUT2 #(
		.INIT('h2)
	) name13202 (
		\sa33_reg[3]/P0001 ,
		_w13733_,
		_w13734_
	);
	LUT2 #(
		.INIT('h2)
	) name13203 (
		\sa33_reg[2]/P0001 ,
		_w12929_,
		_w13735_
	);
	LUT2 #(
		.INIT('h4)
	) name13204 (
		_w13734_,
		_w13735_,
		_w13736_
	);
	LUT2 #(
		.INIT('h2)
	) name13205 (
		\sa33_reg[1]/P0001 ,
		_w13732_,
		_w13737_
	);
	LUT2 #(
		.INIT('h4)
	) name13206 (
		_w13736_,
		_w13737_,
		_w13738_
	);
	LUT2 #(
		.INIT('h8)
	) name13207 (
		_w12544_,
		_w12560_,
		_w13739_
	);
	LUT2 #(
		.INIT('h8)
	) name13208 (
		\sa33_reg[4]/P0001 ,
		_w13739_,
		_w13740_
	);
	LUT2 #(
		.INIT('h4)
	) name13209 (
		\sa33_reg[1]/P0001 ,
		\sa33_reg[2]/P0001 ,
		_w13741_
	);
	LUT2 #(
		.INIT('h1)
	) name13210 (
		_w12445_,
		_w12544_,
		_w13742_
	);
	LUT2 #(
		.INIT('h1)
	) name13211 (
		\sa33_reg[3]/P0001 ,
		_w13742_,
		_w13743_
	);
	LUT2 #(
		.INIT('h1)
	) name13212 (
		_w12501_,
		_w13743_,
		_w13744_
	);
	LUT2 #(
		.INIT('h2)
	) name13213 (
		_w13741_,
		_w13744_,
		_w13745_
	);
	LUT2 #(
		.INIT('h4)
	) name13214 (
		\sa33_reg[7]/NET0131 ,
		_w12478_,
		_w13746_
	);
	LUT2 #(
		.INIT('h1)
	) name13215 (
		_w13740_,
		_w13746_,
		_w13747_
	);
	LUT2 #(
		.INIT('h4)
	) name13216 (
		_w13745_,
		_w13747_,
		_w13748_
	);
	LUT2 #(
		.INIT('h4)
	) name13217 (
		_w13738_,
		_w13748_,
		_w13749_
	);
	LUT2 #(
		.INIT('h4)
	) name13218 (
		_w13727_,
		_w13749_,
		_w13750_
	);
	LUT2 #(
		.INIT('h4)
	) name13219 (
		_w13684_,
		_w13750_,
		_w13751_
	);
	LUT2 #(
		.INIT('h4)
	) name13220 (
		_w13719_,
		_w13751_,
		_w13752_
	);
	LUT2 #(
		.INIT('h8)
	) name13221 (
		\sa22_reg[2]/P0001 ,
		_w12790_,
		_w13753_
	);
	LUT2 #(
		.INIT('h4)
	) name13222 (
		\sa22_reg[3]/P0001 ,
		_w12760_,
		_w13754_
	);
	LUT2 #(
		.INIT('h1)
	) name13223 (
		_w13209_,
		_w13251_,
		_w13755_
	);
	LUT2 #(
		.INIT('h1)
	) name13224 (
		\sa22_reg[2]/P0001 ,
		_w13755_,
		_w13756_
	);
	LUT2 #(
		.INIT('h1)
	) name13225 (
		\sa22_reg[1]/P0001 ,
		_w12806_,
		_w13757_
	);
	LUT2 #(
		.INIT('h1)
	) name13226 (
		_w13275_,
		_w13753_,
		_w13758_
	);
	LUT2 #(
		.INIT('h8)
	) name13227 (
		_w13757_,
		_w13758_,
		_w13759_
	);
	LUT2 #(
		.INIT('h4)
	) name13228 (
		_w13754_,
		_w13759_,
		_w13760_
	);
	LUT2 #(
		.INIT('h4)
	) name13229 (
		_w13756_,
		_w13760_,
		_w13761_
	);
	LUT2 #(
		.INIT('h8)
	) name13230 (
		\sa22_reg[4]/P0001 ,
		_w12721_,
		_w13762_
	);
	LUT2 #(
		.INIT('h1)
	) name13231 (
		_w12295_,
		_w13231_,
		_w13763_
	);
	LUT2 #(
		.INIT('h4)
	) name13232 (
		_w13762_,
		_w13763_,
		_w13764_
	);
	LUT2 #(
		.INIT('h1)
	) name13233 (
		\sa22_reg[2]/P0001 ,
		_w13764_,
		_w13765_
	);
	LUT2 #(
		.INIT('h4)
	) name13234 (
		\sa22_reg[3]/P0001 ,
		_w12319_,
		_w13766_
	);
	LUT2 #(
		.INIT('h1)
	) name13235 (
		_w13220_,
		_w13766_,
		_w13767_
	);
	LUT2 #(
		.INIT('h2)
	) name13236 (
		\sa22_reg[2]/P0001 ,
		_w13767_,
		_w13768_
	);
	LUT2 #(
		.INIT('h8)
	) name13237 (
		_w12237_,
		_w12354_,
		_w13769_
	);
	LUT2 #(
		.INIT('h4)
	) name13238 (
		_w13765_,
		_w13769_,
		_w13770_
	);
	LUT2 #(
		.INIT('h4)
	) name13239 (
		_w13768_,
		_w13770_,
		_w13771_
	);
	LUT2 #(
		.INIT('h1)
	) name13240 (
		_w13761_,
		_w13771_,
		_w13772_
	);
	LUT2 #(
		.INIT('h1)
	) name13241 (
		_w12331_,
		_w12371_,
		_w13773_
	);
	LUT2 #(
		.INIT('h8)
	) name13242 (
		_w12807_,
		_w13773_,
		_w13774_
	);
	LUT2 #(
		.INIT('h2)
	) name13243 (
		\sa22_reg[2]/P0001 ,
		_w12242_,
		_w13775_
	);
	LUT2 #(
		.INIT('h4)
	) name13244 (
		_w13304_,
		_w13775_,
		_w13776_
	);
	LUT2 #(
		.INIT('h1)
	) name13245 (
		_w13774_,
		_w13776_,
		_w13777_
	);
	LUT2 #(
		.INIT('h1)
	) name13246 (
		_w12382_,
		_w13777_,
		_w13778_
	);
	LUT2 #(
		.INIT('h4)
	) name13247 (
		_w13772_,
		_w13778_,
		_w13779_
	);
	LUT2 #(
		.INIT('h1)
	) name13248 (
		\sa22_reg[0]/P0001 ,
		_w13779_,
		_w13780_
	);
	LUT2 #(
		.INIT('h8)
	) name13249 (
		\sa22_reg[4]/P0001 ,
		_w12813_,
		_w13781_
	);
	LUT2 #(
		.INIT('h8)
	) name13250 (
		\sa22_reg[5]/P0001 ,
		_w13268_,
		_w13782_
	);
	LUT2 #(
		.INIT('h1)
	) name13251 (
		_w12747_,
		_w13252_,
		_w13783_
	);
	LUT2 #(
		.INIT('h4)
	) name13252 (
		_w13782_,
		_w13783_,
		_w13784_
	);
	LUT2 #(
		.INIT('h1)
	) name13253 (
		\sa22_reg[2]/P0001 ,
		_w13784_,
		_w13785_
	);
	LUT2 #(
		.INIT('h8)
	) name13254 (
		_w12238_,
		_w12753_,
		_w13786_
	);
	LUT2 #(
		.INIT('h2)
	) name13255 (
		_w12264_,
		_w12282_,
		_w13787_
	);
	LUT2 #(
		.INIT('h1)
	) name13256 (
		_w12381_,
		_w13786_,
		_w13788_
	);
	LUT2 #(
		.INIT('h4)
	) name13257 (
		_w13787_,
		_w13788_,
		_w13789_
	);
	LUT2 #(
		.INIT('h1)
	) name13258 (
		\sa22_reg[1]/P0001 ,
		_w13789_,
		_w13790_
	);
	LUT2 #(
		.INIT('h2)
	) name13259 (
		_w12347_,
		_w13264_,
		_w13791_
	);
	LUT2 #(
		.INIT('h2)
	) name13260 (
		_w12259_,
		_w12731_,
		_w13792_
	);
	LUT2 #(
		.INIT('h1)
	) name13261 (
		_w13791_,
		_w13792_,
		_w13793_
	);
	LUT2 #(
		.INIT('h4)
	) name13262 (
		_w13781_,
		_w13793_,
		_w13794_
	);
	LUT2 #(
		.INIT('h4)
	) name13263 (
		_w13785_,
		_w13794_,
		_w13795_
	);
	LUT2 #(
		.INIT('h4)
	) name13264 (
		_w13790_,
		_w13795_,
		_w13796_
	);
	LUT2 #(
		.INIT('h2)
	) name13265 (
		\sa22_reg[0]/P0001 ,
		_w13796_,
		_w13797_
	);
	LUT2 #(
		.INIT('h1)
	) name13266 (
		_w12296_,
		_w12330_,
		_w13798_
	);
	LUT2 #(
		.INIT('h1)
	) name13267 (
		_w12297_,
		_w13798_,
		_w13799_
	);
	LUT2 #(
		.INIT('h1)
	) name13268 (
		_w12236_,
		_w13190_,
		_w13800_
	);
	LUT2 #(
		.INIT('h4)
	) name13269 (
		_w13799_,
		_w13800_,
		_w13801_
	);
	LUT2 #(
		.INIT('h1)
	) name13270 (
		\sa22_reg[2]/P0001 ,
		_w13801_,
		_w13802_
	);
	LUT2 #(
		.INIT('h8)
	) name13271 (
		\sa22_reg[6]/NET0131 ,
		_w12262_,
		_w13803_
	);
	LUT2 #(
		.INIT('h1)
	) name13272 (
		_w12292_,
		_w13803_,
		_w13804_
	);
	LUT2 #(
		.INIT('h4)
	) name13273 (
		\sa22_reg[5]/P0001 ,
		_w12755_,
		_w13805_
	);
	LUT2 #(
		.INIT('h8)
	) name13274 (
		\sa22_reg[4]/P0001 ,
		_w12257_,
		_w13806_
	);
	LUT2 #(
		.INIT('h1)
	) name13275 (
		_w12805_,
		_w13805_,
		_w13807_
	);
	LUT2 #(
		.INIT('h4)
	) name13276 (
		_w13806_,
		_w13807_,
		_w13808_
	);
	LUT2 #(
		.INIT('h2)
	) name13277 (
		\sa22_reg[2]/P0001 ,
		_w13808_,
		_w13809_
	);
	LUT2 #(
		.INIT('h2)
	) name13278 (
		_w13804_,
		_w13809_,
		_w13810_
	);
	LUT2 #(
		.INIT('h2)
	) name13279 (
		\sa22_reg[0]/P0001 ,
		_w13810_,
		_w13811_
	);
	LUT2 #(
		.INIT('h1)
	) name13280 (
		_w13802_,
		_w13811_,
		_w13812_
	);
	LUT2 #(
		.INIT('h2)
	) name13281 (
		\sa22_reg[1]/P0001 ,
		_w13812_,
		_w13813_
	);
	LUT2 #(
		.INIT('h1)
	) name13282 (
		_w12292_,
		_w12736_,
		_w13814_
	);
	LUT2 #(
		.INIT('h2)
	) name13283 (
		\sa22_reg[3]/P0001 ,
		_w13814_,
		_w13815_
	);
	LUT2 #(
		.INIT('h1)
	) name13284 (
		_w13230_,
		_w13815_,
		_w13816_
	);
	LUT2 #(
		.INIT('h2)
	) name13285 (
		_w13264_,
		_w13816_,
		_w13817_
	);
	LUT2 #(
		.INIT('h1)
	) name13286 (
		_w12396_,
		_w12812_,
		_w13818_
	);
	LUT2 #(
		.INIT('h2)
	) name13287 (
		\sa22_reg[2]/P0001 ,
		_w13818_,
		_w13819_
	);
	LUT2 #(
		.INIT('h4)
	) name13288 (
		\sa22_reg[1]/P0001 ,
		\sa22_reg[2]/P0001 ,
		_w13820_
	);
	LUT2 #(
		.INIT('h1)
	) name13289 (
		_w12275_,
		_w12320_,
		_w13821_
	);
	LUT2 #(
		.INIT('h4)
	) name13290 (
		_w12371_,
		_w13821_,
		_w13822_
	);
	LUT2 #(
		.INIT('h2)
	) name13291 (
		_w13820_,
		_w13822_,
		_w13823_
	);
	LUT2 #(
		.INIT('h1)
	) name13292 (
		_w12733_,
		_w13206_,
		_w13824_
	);
	LUT2 #(
		.INIT('h4)
	) name13293 (
		_w12335_,
		_w13824_,
		_w13825_
	);
	LUT2 #(
		.INIT('h1)
	) name13294 (
		\sa22_reg[2]/P0001 ,
		_w13825_,
		_w13826_
	);
	LUT2 #(
		.INIT('h1)
	) name13295 (
		_w12333_,
		_w12812_,
		_w13827_
	);
	LUT2 #(
		.INIT('h4)
	) name13296 (
		_w13826_,
		_w13827_,
		_w13828_
	);
	LUT2 #(
		.INIT('h1)
	) name13297 (
		\sa22_reg[1]/P0001 ,
		_w13828_,
		_w13829_
	);
	LUT2 #(
		.INIT('h1)
	) name13298 (
		_w13817_,
		_w13819_,
		_w13830_
	);
	LUT2 #(
		.INIT('h4)
	) name13299 (
		_w13823_,
		_w13830_,
		_w13831_
	);
	LUT2 #(
		.INIT('h4)
	) name13300 (
		_w13829_,
		_w13831_,
		_w13832_
	);
	LUT2 #(
		.INIT('h4)
	) name13301 (
		_w13797_,
		_w13832_,
		_w13833_
	);
	LUT2 #(
		.INIT('h4)
	) name13302 (
		_w13813_,
		_w13833_,
		_w13834_
	);
	LUT2 #(
		.INIT('h4)
	) name13303 (
		_w13780_,
		_w13834_,
		_w13835_
	);
	LUT2 #(
		.INIT('h2)
	) name13304 (
		_w13752_,
		_w13835_,
		_w13836_
	);
	LUT2 #(
		.INIT('h4)
	) name13305 (
		_w13752_,
		_w13835_,
		_w13837_
	);
	LUT2 #(
		.INIT('h1)
	) name13306 (
		_w13836_,
		_w13837_,
		_w13838_
	);
	LUT2 #(
		.INIT('h8)
	) name13307 (
		_w12239_,
		_w12297_,
		_w13839_
	);
	LUT2 #(
		.INIT('h1)
	) name13308 (
		_w13782_,
		_w13839_,
		_w13840_
	);
	LUT2 #(
		.INIT('h2)
	) name13309 (
		\sa22_reg[3]/P0001 ,
		_w13840_,
		_w13841_
	);
	LUT2 #(
		.INIT('h1)
	) name13310 (
		_w12396_,
		_w13841_,
		_w13842_
	);
	LUT2 #(
		.INIT('h2)
	) name13311 (
		\sa22_reg[2]/P0001 ,
		_w13842_,
		_w13843_
	);
	LUT2 #(
		.INIT('h8)
	) name13312 (
		_w12244_,
		_w12257_,
		_w13844_
	);
	LUT2 #(
		.INIT('h4)
	) name13313 (
		_w12779_,
		_w13844_,
		_w13845_
	);
	LUT2 #(
		.INIT('h1)
	) name13314 (
		_w12315_,
		_w12733_,
		_w13846_
	);
	LUT2 #(
		.INIT('h1)
	) name13315 (
		\sa22_reg[2]/P0001 ,
		_w13846_,
		_w13847_
	);
	LUT2 #(
		.INIT('h2)
	) name13316 (
		\sa22_reg[1]/P0001 ,
		_w13252_,
		_w13848_
	);
	LUT2 #(
		.INIT('h4)
	) name13317 (
		_w13845_,
		_w13848_,
		_w13849_
	);
	LUT2 #(
		.INIT('h4)
	) name13318 (
		_w13847_,
		_w13849_,
		_w13850_
	);
	LUT2 #(
		.INIT('h8)
	) name13319 (
		_w12344_,
		_w12735_,
		_w13851_
	);
	LUT2 #(
		.INIT('h4)
	) name13320 (
		\sa22_reg[2]/P0001 ,
		_w12755_,
		_w13852_
	);
	LUT2 #(
		.INIT('h1)
	) name13321 (
		\sa22_reg[1]/P0001 ,
		_w12279_,
		_w13853_
	);
	LUT2 #(
		.INIT('h1)
	) name13322 (
		_w13206_,
		_w13852_,
		_w13854_
	);
	LUT2 #(
		.INIT('h8)
	) name13323 (
		_w13853_,
		_w13854_,
		_w13855_
	);
	LUT2 #(
		.INIT('h4)
	) name13324 (
		_w13851_,
		_w13855_,
		_w13856_
	);
	LUT2 #(
		.INIT('h1)
	) name13325 (
		_w13850_,
		_w13856_,
		_w13857_
	);
	LUT2 #(
		.INIT('h1)
	) name13326 (
		_w13303_,
		_w13766_,
		_w13858_
	);
	LUT2 #(
		.INIT('h1)
	) name13327 (
		_w12384_,
		_w13269_,
		_w13859_
	);
	LUT2 #(
		.INIT('h8)
	) name13328 (
		_w13858_,
		_w13859_,
		_w13860_
	);
	LUT2 #(
		.INIT('h1)
	) name13329 (
		\sa22_reg[2]/P0001 ,
		_w13860_,
		_w13861_
	);
	LUT2 #(
		.INIT('h1)
	) name13330 (
		_w13843_,
		_w13861_,
		_w13862_
	);
	LUT2 #(
		.INIT('h4)
	) name13331 (
		_w13857_,
		_w13862_,
		_w13863_
	);
	LUT2 #(
		.INIT('h1)
	) name13332 (
		\sa22_reg[0]/P0001 ,
		_w13863_,
		_w13864_
	);
	LUT2 #(
		.INIT('h8)
	) name13333 (
		_w12322_,
		_w13805_,
		_w13865_
	);
	LUT2 #(
		.INIT('h2)
	) name13334 (
		_w12239_,
		_w12755_,
		_w13866_
	);
	LUT2 #(
		.INIT('h1)
	) name13335 (
		_w12252_,
		_w13240_,
		_w13867_
	);
	LUT2 #(
		.INIT('h4)
	) name13336 (
		_w13866_,
		_w13867_,
		_w13868_
	);
	LUT2 #(
		.INIT('h1)
	) name13337 (
		\sa22_reg[2]/P0001 ,
		_w13868_,
		_w13869_
	);
	LUT2 #(
		.INIT('h4)
	) name13338 (
		_w12282_,
		_w13368_,
		_w13870_
	);
	LUT2 #(
		.INIT('h1)
	) name13339 (
		_w12814_,
		_w13865_,
		_w13871_
	);
	LUT2 #(
		.INIT('h4)
	) name13340 (
		_w13870_,
		_w13871_,
		_w13872_
	);
	LUT2 #(
		.INIT('h4)
	) name13341 (
		_w13869_,
		_w13872_,
		_w13873_
	);
	LUT2 #(
		.INIT('h1)
	) name13342 (
		\sa22_reg[1]/P0001 ,
		_w13873_,
		_w13874_
	);
	LUT2 #(
		.INIT('h1)
	) name13343 (
		_w12290_,
		_w12352_,
		_w13875_
	);
	LUT2 #(
		.INIT('h1)
	) name13344 (
		_w13240_,
		_w13265_,
		_w13876_
	);
	LUT2 #(
		.INIT('h8)
	) name13345 (
		_w13875_,
		_w13876_,
		_w13877_
	);
	LUT2 #(
		.INIT('h2)
	) name13346 (
		\sa22_reg[2]/P0001 ,
		_w13877_,
		_w13878_
	);
	LUT2 #(
		.INIT('h4)
	) name13347 (
		\sa22_reg[2]/P0001 ,
		_w12275_,
		_w13879_
	);
	LUT2 #(
		.INIT('h1)
	) name13348 (
		_w12722_,
		_w13879_,
		_w13880_
	);
	LUT2 #(
		.INIT('h4)
	) name13349 (
		_w13878_,
		_w13880_,
		_w13881_
	);
	LUT2 #(
		.INIT('h2)
	) name13350 (
		\sa22_reg[1]/P0001 ,
		_w13881_,
		_w13882_
	);
	LUT2 #(
		.INIT('h8)
	) name13351 (
		\sa22_reg[6]/NET0131 ,
		_w12385_,
		_w13883_
	);
	LUT2 #(
		.INIT('h8)
	) name13352 (
		_w12257_,
		_w12303_,
		_w13884_
	);
	LUT2 #(
		.INIT('h1)
	) name13353 (
		_w12246_,
		_w13884_,
		_w13885_
	);
	LUT2 #(
		.INIT('h4)
	) name13354 (
		_w12253_,
		_w13885_,
		_w13886_
	);
	LUT2 #(
		.INIT('h4)
	) name13355 (
		_w13883_,
		_w13886_,
		_w13887_
	);
	LUT2 #(
		.INIT('h2)
	) name13356 (
		\sa22_reg[2]/P0001 ,
		_w13887_,
		_w13888_
	);
	LUT2 #(
		.INIT('h8)
	) name13357 (
		_w12252_,
		_w13200_,
		_w13889_
	);
	LUT2 #(
		.INIT('h1)
	) name13358 (
		_w13316_,
		_w13889_,
		_w13890_
	);
	LUT2 #(
		.INIT('h4)
	) name13359 (
		_w13888_,
		_w13890_,
		_w13891_
	);
	LUT2 #(
		.INIT('h4)
	) name13360 (
		_w13874_,
		_w13891_,
		_w13892_
	);
	LUT2 #(
		.INIT('h4)
	) name13361 (
		_w13882_,
		_w13892_,
		_w13893_
	);
	LUT2 #(
		.INIT('h2)
	) name13362 (
		\sa22_reg[0]/P0001 ,
		_w13893_,
		_w13894_
	);
	LUT2 #(
		.INIT('h2)
	) name13363 (
		_w12245_,
		_w12755_,
		_w13895_
	);
	LUT2 #(
		.INIT('h2)
	) name13364 (
		_w13332_,
		_w13895_,
		_w13896_
	);
	LUT2 #(
		.INIT('h2)
	) name13365 (
		_w13227_,
		_w13896_,
		_w13897_
	);
	LUT2 #(
		.INIT('h8)
	) name13366 (
		\sa22_reg[7]/NET0131 ,
		_w12290_,
		_w13898_
	);
	LUT2 #(
		.INIT('h1)
	) name13367 (
		_w12738_,
		_w12773_,
		_w13899_
	);
	LUT2 #(
		.INIT('h4)
	) name13368 (
		_w13898_,
		_w13899_,
		_w13900_
	);
	LUT2 #(
		.INIT('h1)
	) name13369 (
		\sa22_reg[3]/P0001 ,
		_w13900_,
		_w13901_
	);
	LUT2 #(
		.INIT('h1)
	) name13370 (
		_w12292_,
		_w12351_,
		_w13902_
	);
	LUT2 #(
		.INIT('h4)
	) name13371 (
		_w13901_,
		_w13902_,
		_w13903_
	);
	LUT2 #(
		.INIT('h2)
	) name13372 (
		\sa22_reg[2]/P0001 ,
		_w13903_,
		_w13904_
	);
	LUT2 #(
		.INIT('h1)
	) name13373 (
		_w13897_,
		_w13904_,
		_w13905_
	);
	LUT2 #(
		.INIT('h2)
	) name13374 (
		\sa22_reg[1]/P0001 ,
		_w13905_,
		_w13906_
	);
	LUT2 #(
		.INIT('h4)
	) name13375 (
		_w13229_,
		_w13858_,
		_w13907_
	);
	LUT2 #(
		.INIT('h1)
	) name13376 (
		\sa22_reg[2]/P0001 ,
		_w13907_,
		_w13908_
	);
	LUT2 #(
		.INIT('h1)
	) name13377 (
		_w13358_,
		_w13908_,
		_w13909_
	);
	LUT2 #(
		.INIT('h1)
	) name13378 (
		\sa22_reg[1]/P0001 ,
		_w13909_,
		_w13910_
	);
	LUT2 #(
		.INIT('h8)
	) name13379 (
		_w12234_,
		_w12260_,
		_w13911_
	);
	LUT2 #(
		.INIT('h1)
	) name13380 (
		_w12240_,
		_w13911_,
		_w13912_
	);
	LUT2 #(
		.INIT('h2)
	) name13381 (
		_w12779_,
		_w13912_,
		_w13913_
	);
	LUT2 #(
		.INIT('h8)
	) name13382 (
		_w12239_,
		_w12244_,
		_w13914_
	);
	LUT2 #(
		.INIT('h1)
	) name13383 (
		_w12236_,
		_w13914_,
		_w13915_
	);
	LUT2 #(
		.INIT('h4)
	) name13384 (
		_w12722_,
		_w13915_,
		_w13916_
	);
	LUT2 #(
		.INIT('h2)
	) name13385 (
		_w13820_,
		_w13916_,
		_w13917_
	);
	LUT2 #(
		.INIT('h1)
	) name13386 (
		_w13913_,
		_w13917_,
		_w13918_
	);
	LUT2 #(
		.INIT('h4)
	) name13387 (
		_w13910_,
		_w13918_,
		_w13919_
	);
	LUT2 #(
		.INIT('h4)
	) name13388 (
		_w13906_,
		_w13919_,
		_w13920_
	);
	LUT2 #(
		.INIT('h4)
	) name13389 (
		_w13864_,
		_w13920_,
		_w13921_
	);
	LUT2 #(
		.INIT('h4)
	) name13390 (
		_w13894_,
		_w13921_,
		_w13922_
	);
	LUT2 #(
		.INIT('h2)
	) name13391 (
		\u0_w_reg[0][17]/P0001 ,
		_w13922_,
		_w13923_
	);
	LUT2 #(
		.INIT('h4)
	) name13392 (
		\u0_w_reg[0][17]/P0001 ,
		_w13922_,
		_w13924_
	);
	LUT2 #(
		.INIT('h1)
	) name13393 (
		_w13923_,
		_w13924_,
		_w13925_
	);
	LUT2 #(
		.INIT('h8)
	) name13394 (
		_w13838_,
		_w13925_,
		_w13926_
	);
	LUT2 #(
		.INIT('h1)
	) name13395 (
		_w13838_,
		_w13925_,
		_w13927_
	);
	LUT2 #(
		.INIT('h1)
	) name13396 (
		_w13926_,
		_w13927_,
		_w13928_
	);
	LUT2 #(
		.INIT('h2)
	) name13397 (
		_w13655_,
		_w13928_,
		_w13929_
	);
	LUT2 #(
		.INIT('h4)
	) name13398 (
		_w13655_,
		_w13928_,
		_w13930_
	);
	LUT2 #(
		.INIT('h1)
	) name13399 (
		\ld_r_reg/P0001 ,
		_w13929_,
		_w13931_
	);
	LUT2 #(
		.INIT('h4)
	) name13400 (
		_w13930_,
		_w13931_,
		_w13932_
	);
	LUT2 #(
		.INIT('h1)
	) name13401 (
		\text_in_r_reg[113]/P0001 ,
		\u0_w_reg[0][17]/P0001 ,
		_w13933_
	);
	LUT2 #(
		.INIT('h8)
	) name13402 (
		\text_in_r_reg[113]/P0001 ,
		\u0_w_reg[0][17]/P0001 ,
		_w13934_
	);
	LUT2 #(
		.INIT('h2)
	) name13403 (
		\ld_r_reg/P0001 ,
		_w13933_,
		_w13935_
	);
	LUT2 #(
		.INIT('h4)
	) name13404 (
		_w13934_,
		_w13935_,
		_w13936_
	);
	LUT2 #(
		.INIT('h1)
	) name13405 (
		_w13932_,
		_w13936_,
		_w13937_
	);
	LUT2 #(
		.INIT('h2)
	) name13406 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[5]/P0001 ,
		_w13938_
	);
	LUT2 #(
		.INIT('h8)
	) name13407 (
		\sa33_reg[3]/P0001 ,
		_w12467_,
		_w13939_
	);
	LUT2 #(
		.INIT('h1)
	) name13408 (
		_w12465_,
		_w13939_,
		_w13940_
	);
	LUT2 #(
		.INIT('h2)
	) name13409 (
		_w13938_,
		_w13940_,
		_w13941_
	);
	LUT2 #(
		.INIT('h1)
	) name13410 (
		_w13721_,
		_w13941_,
		_w13942_
	);
	LUT2 #(
		.INIT('h1)
	) name13411 (
		\sa33_reg[1]/P0001 ,
		_w13942_,
		_w13943_
	);
	LUT2 #(
		.INIT('h8)
	) name13412 (
		\sa33_reg[7]/NET0131 ,
		_w12932_,
		_w13944_
	);
	LUT2 #(
		.INIT('h1)
	) name13413 (
		_w13667_,
		_w13944_,
		_w13945_
	);
	LUT2 #(
		.INIT('h2)
	) name13414 (
		_w12560_,
		_w13945_,
		_w13946_
	);
	LUT2 #(
		.INIT('h1)
	) name13415 (
		\sa33_reg[1]/P0001 ,
		\sa33_reg[2]/P0001 ,
		_w13947_
	);
	LUT2 #(
		.INIT('h8)
	) name13416 (
		_w12876_,
		_w13947_,
		_w13948_
	);
	LUT2 #(
		.INIT('h8)
	) name13417 (
		_w12457_,
		_w12465_,
		_w13949_
	);
	LUT2 #(
		.INIT('h1)
	) name13418 (
		_w12550_,
		_w13949_,
		_w13950_
	);
	LUT2 #(
		.INIT('h1)
	) name13419 (
		\sa33_reg[2]/P0001 ,
		_w13950_,
		_w13951_
	);
	LUT2 #(
		.INIT('h1)
	) name13420 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		_w13952_
	);
	LUT2 #(
		.INIT('h1)
	) name13421 (
		_w12481_,
		_w12525_,
		_w13953_
	);
	LUT2 #(
		.INIT('h2)
	) name13422 (
		_w13952_,
		_w13953_,
		_w13954_
	);
	LUT2 #(
		.INIT('h2)
	) name13423 (
		_w12450_,
		_w12881_,
		_w13955_
	);
	LUT2 #(
		.INIT('h1)
	) name13424 (
		_w12880_,
		_w13720_,
		_w13956_
	);
	LUT2 #(
		.INIT('h1)
	) name13425 (
		\sa33_reg[2]/P0001 ,
		_w13956_,
		_w13957_
	);
	LUT2 #(
		.INIT('h1)
	) name13426 (
		_w13668_,
		_w13955_,
		_w13958_
	);
	LUT2 #(
		.INIT('h4)
	) name13427 (
		_w13957_,
		_w13958_,
		_w13959_
	);
	LUT2 #(
		.INIT('h2)
	) name13428 (
		\sa33_reg[1]/P0001 ,
		_w13959_,
		_w13960_
	);
	LUT2 #(
		.INIT('h1)
	) name13429 (
		_w13746_,
		_w13948_,
		_w13961_
	);
	LUT2 #(
		.INIT('h4)
	) name13430 (
		_w13954_,
		_w13961_,
		_w13962_
	);
	LUT2 #(
		.INIT('h1)
	) name13431 (
		_w13946_,
		_w13951_,
		_w13963_
	);
	LUT2 #(
		.INIT('h8)
	) name13432 (
		_w13962_,
		_w13963_,
		_w13964_
	);
	LUT2 #(
		.INIT('h4)
	) name13433 (
		_w13943_,
		_w13964_,
		_w13965_
	);
	LUT2 #(
		.INIT('h4)
	) name13434 (
		_w13960_,
		_w13965_,
		_w13966_
	);
	LUT2 #(
		.INIT('h1)
	) name13435 (
		\sa33_reg[0]/P0001 ,
		_w13966_,
		_w13967_
	);
	LUT2 #(
		.INIT('h2)
	) name13436 (
		_w12433_,
		_w12855_,
		_w13968_
	);
	LUT2 #(
		.INIT('h8)
	) name13437 (
		_w12551_,
		_w13938_,
		_w13969_
	);
	LUT2 #(
		.INIT('h8)
	) name13438 (
		\sa33_reg[4]/P0001 ,
		_w12475_,
		_w13970_
	);
	LUT2 #(
		.INIT('h2)
	) name13439 (
		_w12480_,
		_w12876_,
		_w13971_
	);
	LUT2 #(
		.INIT('h1)
	) name13440 (
		_w12422_,
		_w13970_,
		_w13972_
	);
	LUT2 #(
		.INIT('h4)
	) name13441 (
		_w13971_,
		_w13972_,
		_w13973_
	);
	LUT2 #(
		.INIT('h1)
	) name13442 (
		\sa33_reg[2]/P0001 ,
		_w13973_,
		_w13974_
	);
	LUT2 #(
		.INIT('h1)
	) name13443 (
		_w12565_,
		_w13968_,
		_w13975_
	);
	LUT2 #(
		.INIT('h4)
	) name13444 (
		_w13969_,
		_w13975_,
		_w13976_
	);
	LUT2 #(
		.INIT('h4)
	) name13445 (
		_w13974_,
		_w13976_,
		_w13977_
	);
	LUT2 #(
		.INIT('h1)
	) name13446 (
		\sa33_reg[1]/P0001 ,
		_w13977_,
		_w13978_
	);
	LUT2 #(
		.INIT('h8)
	) name13447 (
		_w12422_,
		_w13952_,
		_w13979_
	);
	LUT2 #(
		.INIT('h8)
	) name13448 (
		_w12461_,
		_w13952_,
		_w13980_
	);
	LUT2 #(
		.INIT('h4)
	) name13449 (
		\sa33_reg[6]/P0001 ,
		_w13980_,
		_w13981_
	);
	LUT2 #(
		.INIT('h1)
	) name13450 (
		_w12900_,
		_w13981_,
		_w13982_
	);
	LUT2 #(
		.INIT('h2)
	) name13451 (
		\sa33_reg[1]/P0001 ,
		_w13982_,
		_w13983_
	);
	LUT2 #(
		.INIT('h8)
	) name13452 (
		_w12477_,
		_w12521_,
		_w13984_
	);
	LUT2 #(
		.INIT('h1)
	) name13453 (
		_w12460_,
		_w13970_,
		_w13985_
	);
	LUT2 #(
		.INIT('h4)
	) name13454 (
		\sa33_reg[3]/P0001 ,
		_w12465_,
		_w13986_
	);
	LUT2 #(
		.INIT('h1)
	) name13455 (
		_w12531_,
		_w13986_,
		_w13987_
	);
	LUT2 #(
		.INIT('h8)
	) name13456 (
		_w13985_,
		_w13987_,
		_w13988_
	);
	LUT2 #(
		.INIT('h2)
	) name13457 (
		\sa33_reg[1]/P0001 ,
		_w13988_,
		_w13989_
	);
	LUT2 #(
		.INIT('h8)
	) name13458 (
		\sa33_reg[6]/P0001 ,
		_w12551_,
		_w13990_
	);
	LUT2 #(
		.INIT('h1)
	) name13459 (
		_w12423_,
		_w12431_,
		_w13991_
	);
	LUT2 #(
		.INIT('h4)
	) name13460 (
		_w13990_,
		_w13991_,
		_w13992_
	);
	LUT2 #(
		.INIT('h4)
	) name13461 (
		_w13989_,
		_w13992_,
		_w13993_
	);
	LUT2 #(
		.INIT('h2)
	) name13462 (
		\sa33_reg[2]/P0001 ,
		_w13993_,
		_w13994_
	);
	LUT2 #(
		.INIT('h1)
	) name13463 (
		_w12569_,
		_w13979_,
		_w13995_
	);
	LUT2 #(
		.INIT('h4)
	) name13464 (
		_w13984_,
		_w13995_,
		_w13996_
	);
	LUT2 #(
		.INIT('h4)
	) name13465 (
		_w13983_,
		_w13996_,
		_w13997_
	);
	LUT2 #(
		.INIT('h4)
	) name13466 (
		_w13978_,
		_w13997_,
		_w13998_
	);
	LUT2 #(
		.INIT('h4)
	) name13467 (
		_w13994_,
		_w13998_,
		_w13999_
	);
	LUT2 #(
		.INIT('h2)
	) name13468 (
		\sa33_reg[0]/P0001 ,
		_w13999_,
		_w14000_
	);
	LUT2 #(
		.INIT('h8)
	) name13469 (
		_w12448_,
		_w12480_,
		_w14001_
	);
	LUT2 #(
		.INIT('h1)
	) name13470 (
		_w12428_,
		_w14001_,
		_w14002_
	);
	LUT2 #(
		.INIT('h4)
	) name13471 (
		_w12900_,
		_w14002_,
		_w14003_
	);
	LUT2 #(
		.INIT('h2)
	) name13472 (
		\sa33_reg[2]/P0001 ,
		_w14003_,
		_w14004_
	);
	LUT2 #(
		.INIT('h8)
	) name13473 (
		\sa33_reg[3]/P0001 ,
		_w12461_,
		_w14005_
	);
	LUT2 #(
		.INIT('h8)
	) name13474 (
		_w12884_,
		_w14005_,
		_w14006_
	);
	LUT2 #(
		.INIT('h1)
	) name13475 (
		_w12506_,
		_w14006_,
		_w14007_
	);
	LUT2 #(
		.INIT('h4)
	) name13476 (
		_w13954_,
		_w14007_,
		_w14008_
	);
	LUT2 #(
		.INIT('h4)
	) name13477 (
		_w14004_,
		_w14008_,
		_w14009_
	);
	LUT2 #(
		.INIT('h1)
	) name13478 (
		\sa33_reg[1]/P0001 ,
		_w14009_,
		_w14010_
	);
	LUT2 #(
		.INIT('h8)
	) name13479 (
		_w12479_,
		_w12480_,
		_w14011_
	);
	LUT2 #(
		.INIT('h8)
	) name13480 (
		_w12419_,
		_w12475_,
		_w14012_
	);
	LUT2 #(
		.INIT('h1)
	) name13481 (
		_w14011_,
		_w14012_,
		_w14013_
	);
	LUT2 #(
		.INIT('h2)
	) name13482 (
		_w12881_,
		_w14013_,
		_w14014_
	);
	LUT2 #(
		.INIT('h2)
	) name13483 (
		_w12429_,
		_w12876_,
		_w14015_
	);
	LUT2 #(
		.INIT('h8)
	) name13484 (
		_w12480_,
		_w12876_,
		_w14016_
	);
	LUT2 #(
		.INIT('h1)
	) name13485 (
		_w12906_,
		_w14016_,
		_w14017_
	);
	LUT2 #(
		.INIT('h4)
	) name13486 (
		_w14015_,
		_w14017_,
		_w14018_
	);
	LUT2 #(
		.INIT('h8)
	) name13487 (
		\sa33_reg[1]/P0001 ,
		_w12456_,
		_w14019_
	);
	LUT2 #(
		.INIT('h4)
	) name13488 (
		_w14018_,
		_w14019_,
		_w14020_
	);
	LUT2 #(
		.INIT('h8)
	) name13489 (
		\sa33_reg[1]/P0001 ,
		\sa33_reg[2]/P0001 ,
		_w14021_
	);
	LUT2 #(
		.INIT('h2)
	) name13490 (
		\sa33_reg[7]/NET0131 ,
		_w13985_,
		_w14022_
	);
	LUT2 #(
		.INIT('h8)
	) name13491 (
		_w12429_,
		_w12444_,
		_w14023_
	);
	LUT2 #(
		.INIT('h1)
	) name13492 (
		_w14022_,
		_w14023_,
		_w14024_
	);
	LUT2 #(
		.INIT('h1)
	) name13493 (
		\sa33_reg[3]/P0001 ,
		_w14024_,
		_w14025_
	);
	LUT2 #(
		.INIT('h1)
	) name13494 (
		_w12462_,
		_w12913_,
		_w14026_
	);
	LUT2 #(
		.INIT('h4)
	) name13495 (
		_w14025_,
		_w14026_,
		_w14027_
	);
	LUT2 #(
		.INIT('h2)
	) name13496 (
		_w14021_,
		_w14027_,
		_w14028_
	);
	LUT2 #(
		.INIT('h1)
	) name13497 (
		_w14014_,
		_w14020_,
		_w14029_
	);
	LUT2 #(
		.INIT('h4)
	) name13498 (
		_w14010_,
		_w14029_,
		_w14030_
	);
	LUT2 #(
		.INIT('h4)
	) name13499 (
		_w14028_,
		_w14030_,
		_w14031_
	);
	LUT2 #(
		.INIT('h4)
	) name13500 (
		_w13967_,
		_w14031_,
		_w14032_
	);
	LUT2 #(
		.INIT('h4)
	) name13501 (
		_w14000_,
		_w14032_,
		_w14033_
	);
	LUT2 #(
		.INIT('h1)
	) name13502 (
		\sa33_reg[2]/P0001 ,
		_w12429_,
		_w14034_
	);
	LUT2 #(
		.INIT('h1)
	) name13503 (
		\sa33_reg[5]/P0001 ,
		_w12465_,
		_w14035_
	);
	LUT2 #(
		.INIT('h2)
	) name13504 (
		_w14034_,
		_w14035_,
		_w14036_
	);
	LUT2 #(
		.INIT('h1)
	) name13505 (
		_w13698_,
		_w14036_,
		_w14037_
	);
	LUT2 #(
		.INIT('h2)
	) name13506 (
		\sa33_reg[1]/P0001 ,
		_w14037_,
		_w14038_
	);
	LUT2 #(
		.INIT('h1)
	) name13507 (
		_w12444_,
		_w12521_,
		_w14039_
	);
	LUT2 #(
		.INIT('h2)
	) name13508 (
		_w12456_,
		_w14039_,
		_w14040_
	);
	LUT2 #(
		.INIT('h1)
	) name13509 (
		_w12569_,
		_w13944_,
		_w14041_
	);
	LUT2 #(
		.INIT('h1)
	) name13510 (
		\sa33_reg[2]/P0001 ,
		_w14041_,
		_w14042_
	);
	LUT2 #(
		.INIT('h1)
	) name13511 (
		_w12512_,
		_w13721_,
		_w14043_
	);
	LUT2 #(
		.INIT('h8)
	) name13512 (
		_w12475_,
		_w12876_,
		_w14044_
	);
	LUT2 #(
		.INIT('h1)
	) name13513 (
		_w12507_,
		_w14044_,
		_w14045_
	);
	LUT2 #(
		.INIT('h8)
	) name13514 (
		_w14043_,
		_w14045_,
		_w14046_
	);
	LUT2 #(
		.INIT('h2)
	) name13515 (
		\sa33_reg[2]/P0001 ,
		_w14046_,
		_w14047_
	);
	LUT2 #(
		.INIT('h8)
	) name13516 (
		_w12448_,
		_w12942_,
		_w14048_
	);
	LUT2 #(
		.INIT('h8)
	) name13517 (
		\sa33_reg[2]/P0001 ,
		_w13986_,
		_w14049_
	);
	LUT2 #(
		.INIT('h1)
	) name13518 (
		_w14048_,
		_w14049_,
		_w14050_
	);
	LUT2 #(
		.INIT('h1)
	) name13519 (
		\sa33_reg[5]/P0001 ,
		_w14050_,
		_w14051_
	);
	LUT2 #(
		.INIT('h8)
	) name13520 (
		_w12479_,
		_w12510_,
		_w14052_
	);
	LUT2 #(
		.INIT('h1)
	) name13521 (
		_w12423_,
		_w12522_,
		_w14053_
	);
	LUT2 #(
		.INIT('h2)
	) name13522 (
		\sa33_reg[2]/P0001 ,
		_w14053_,
		_w14054_
	);
	LUT2 #(
		.INIT('h1)
	) name13523 (
		_w12447_,
		_w12509_,
		_w14055_
	);
	LUT2 #(
		.INIT('h4)
	) name13524 (
		_w14052_,
		_w14055_,
		_w14056_
	);
	LUT2 #(
		.INIT('h4)
	) name13525 (
		_w14051_,
		_w14056_,
		_w14057_
	);
	LUT2 #(
		.INIT('h4)
	) name13526 (
		_w14054_,
		_w14057_,
		_w14058_
	);
	LUT2 #(
		.INIT('h1)
	) name13527 (
		\sa33_reg[1]/P0001 ,
		_w14058_,
		_w14059_
	);
	LUT2 #(
		.INIT('h1)
	) name13528 (
		_w12899_,
		_w12927_,
		_w14060_
	);
	LUT2 #(
		.INIT('h4)
	) name13529 (
		_w14040_,
		_w14060_,
		_w14061_
	);
	LUT2 #(
		.INIT('h4)
	) name13530 (
		_w14038_,
		_w14061_,
		_w14062_
	);
	LUT2 #(
		.INIT('h4)
	) name13531 (
		_w14042_,
		_w14062_,
		_w14063_
	);
	LUT2 #(
		.INIT('h4)
	) name13532 (
		_w14047_,
		_w14063_,
		_w14064_
	);
	LUT2 #(
		.INIT('h4)
	) name13533 (
		_w14059_,
		_w14064_,
		_w14065_
	);
	LUT2 #(
		.INIT('h2)
	) name13534 (
		\sa33_reg[0]/P0001 ,
		_w14065_,
		_w14066_
	);
	LUT2 #(
		.INIT('h1)
	) name13535 (
		_w12521_,
		_w12561_,
		_w14067_
	);
	LUT2 #(
		.INIT('h2)
	) name13536 (
		_w12476_,
		_w14067_,
		_w14068_
	);
	LUT2 #(
		.INIT('h4)
	) name13537 (
		\sa33_reg[1]/P0001 ,
		_w12418_,
		_w14069_
	);
	LUT2 #(
		.INIT('h4)
	) name13538 (
		_w12877_,
		_w14069_,
		_w14070_
	);
	LUT2 #(
		.INIT('h1)
	) name13539 (
		_w14068_,
		_w14070_,
		_w14071_
	);
	LUT2 #(
		.INIT('h2)
	) name13540 (
		\sa33_reg[2]/P0001 ,
		_w14071_,
		_w14072_
	);
	LUT2 #(
		.INIT('h8)
	) name13541 (
		_w12475_,
		_w12479_,
		_w14073_
	);
	LUT2 #(
		.INIT('h1)
	) name13542 (
		_w12507_,
		_w13662_,
		_w14074_
	);
	LUT2 #(
		.INIT('h4)
	) name13543 (
		_w14073_,
		_w14074_,
		_w14075_
	);
	LUT2 #(
		.INIT('h1)
	) name13544 (
		\sa33_reg[2]/P0001 ,
		_w14075_,
		_w14076_
	);
	LUT2 #(
		.INIT('h8)
	) name13545 (
		_w12412_,
		_w12419_,
		_w14077_
	);
	LUT2 #(
		.INIT('h4)
	) name13546 (
		_w12419_,
		_w12465_,
		_w14078_
	);
	LUT2 #(
		.INIT('h8)
	) name13547 (
		\sa33_reg[2]/P0001 ,
		_w12913_,
		_w14079_
	);
	LUT2 #(
		.INIT('h2)
	) name13548 (
		\sa33_reg[1]/P0001 ,
		_w13980_,
		_w14080_
	);
	LUT2 #(
		.INIT('h1)
	) name13549 (
		_w14077_,
		_w14078_,
		_w14081_
	);
	LUT2 #(
		.INIT('h8)
	) name13550 (
		_w14080_,
		_w14081_,
		_w14082_
	);
	LUT2 #(
		.INIT('h4)
	) name13551 (
		_w14079_,
		_w14082_,
		_w14083_
	);
	LUT2 #(
		.INIT('h1)
	) name13552 (
		\sa33_reg[3]/P0001 ,
		_w14017_,
		_w14084_
	);
	LUT2 #(
		.INIT('h1)
	) name13553 (
		\sa33_reg[1]/P0001 ,
		_w12882_,
		_w14085_
	);
	LUT2 #(
		.INIT('h4)
	) name13554 (
		_w14084_,
		_w14085_,
		_w14086_
	);
	LUT2 #(
		.INIT('h1)
	) name13555 (
		_w14083_,
		_w14086_,
		_w14087_
	);
	LUT2 #(
		.INIT('h1)
	) name13556 (
		_w14072_,
		_w14076_,
		_w14088_
	);
	LUT2 #(
		.INIT('h4)
	) name13557 (
		_w14087_,
		_w14088_,
		_w14089_
	);
	LUT2 #(
		.INIT('h1)
	) name13558 (
		\sa33_reg[0]/P0001 ,
		_w14089_,
		_w14090_
	);
	LUT2 #(
		.INIT('h4)
	) name13559 (
		\sa33_reg[2]/P0001 ,
		_w13939_,
		_w14091_
	);
	LUT2 #(
		.INIT('h8)
	) name13560 (
		_w12472_,
		_w12525_,
		_w14092_
	);
	LUT2 #(
		.INIT('h1)
	) name13561 (
		_w14091_,
		_w14092_,
		_w14093_
	);
	LUT2 #(
		.INIT('h2)
	) name13562 (
		\sa33_reg[6]/P0001 ,
		_w14093_,
		_w14094_
	);
	LUT2 #(
		.INIT('h8)
	) name13563 (
		_w13685_,
		_w13952_,
		_w14095_
	);
	LUT2 #(
		.INIT('h4)
	) name13564 (
		\sa33_reg[5]/P0001 ,
		_w12898_,
		_w14096_
	);
	LUT2 #(
		.INIT('h1)
	) name13565 (
		_w12863_,
		_w13739_,
		_w14097_
	);
	LUT2 #(
		.INIT('h4)
	) name13566 (
		_w14095_,
		_w14097_,
		_w14098_
	);
	LUT2 #(
		.INIT('h2)
	) name13567 (
		_w12871_,
		_w14096_,
		_w14099_
	);
	LUT2 #(
		.INIT('h8)
	) name13568 (
		_w14098_,
		_w14099_,
		_w14100_
	);
	LUT2 #(
		.INIT('h2)
	) name13569 (
		_w12911_,
		_w14011_,
		_w14101_
	);
	LUT2 #(
		.INIT('h4)
	) name13570 (
		_w12410_,
		_w12433_,
		_w14102_
	);
	LUT2 #(
		.INIT('h1)
	) name13571 (
		\sa33_reg[2]/P0001 ,
		_w12909_,
		_w14103_
	);
	LUT2 #(
		.INIT('h4)
	) name13572 (
		_w14102_,
		_w14103_,
		_w14104_
	);
	LUT2 #(
		.INIT('h1)
	) name13573 (
		_w14101_,
		_w14104_,
		_w14105_
	);
	LUT2 #(
		.INIT('h8)
	) name13574 (
		_w12415_,
		_w12456_,
		_w14106_
	);
	LUT2 #(
		.INIT('h1)
	) name13575 (
		\sa33_reg[1]/P0001 ,
		_w14106_,
		_w14107_
	);
	LUT2 #(
		.INIT('h4)
	) name13576 (
		_w12563_,
		_w14107_,
		_w14108_
	);
	LUT2 #(
		.INIT('h4)
	) name13577 (
		_w14105_,
		_w14108_,
		_w14109_
	);
	LUT2 #(
		.INIT('h1)
	) name13578 (
		_w14100_,
		_w14109_,
		_w14110_
	);
	LUT2 #(
		.INIT('h1)
	) name13579 (
		_w14094_,
		_w14110_,
		_w14111_
	);
	LUT2 #(
		.INIT('h4)
	) name13580 (
		_w14090_,
		_w14111_,
		_w14112_
	);
	LUT2 #(
		.INIT('h4)
	) name13581 (
		_w14066_,
		_w14112_,
		_w14113_
	);
	LUT2 #(
		.INIT('h2)
	) name13582 (
		_w14033_,
		_w14113_,
		_w14114_
	);
	LUT2 #(
		.INIT('h4)
	) name13583 (
		_w14033_,
		_w14113_,
		_w14115_
	);
	LUT2 #(
		.INIT('h1)
	) name13584 (
		_w14114_,
		_w14115_,
		_w14116_
	);
	LUT2 #(
		.INIT('h2)
	) name13585 (
		\u0_w_reg[0][9]/P0001 ,
		_w13752_,
		_w14117_
	);
	LUT2 #(
		.INIT('h4)
	) name13586 (
		\u0_w_reg[0][9]/P0001 ,
		_w13752_,
		_w14118_
	);
	LUT2 #(
		.INIT('h1)
	) name13587 (
		_w14117_,
		_w14118_,
		_w14119_
	);
	LUT2 #(
		.INIT('h8)
	) name13588 (
		_w14116_,
		_w14119_,
		_w14120_
	);
	LUT2 #(
		.INIT('h1)
	) name13589 (
		_w14116_,
		_w14119_,
		_w14121_
	);
	LUT2 #(
		.INIT('h1)
	) name13590 (
		_w14120_,
		_w14121_,
		_w14122_
	);
	LUT2 #(
		.INIT('h2)
	) name13591 (
		_w13379_,
		_w13922_,
		_w14123_
	);
	LUT2 #(
		.INIT('h4)
	) name13592 (
		_w13379_,
		_w13922_,
		_w14124_
	);
	LUT2 #(
		.INIT('h1)
	) name13593 (
		_w14123_,
		_w14124_,
		_w14125_
	);
	LUT2 #(
		.INIT('h1)
	) name13594 (
		_w12152_,
		_w13522_,
		_w14126_
	);
	LUT2 #(
		.INIT('h2)
	) name13595 (
		\sa11_reg[2]/P0001 ,
		_w14126_,
		_w14127_
	);
	LUT2 #(
		.INIT('h8)
	) name13596 (
		_w11794_,
		_w11816_,
		_w14128_
	);
	LUT2 #(
		.INIT('h1)
	) name13597 (
		_w12169_,
		_w13139_,
		_w14129_
	);
	LUT2 #(
		.INIT('h4)
	) name13598 (
		_w14128_,
		_w14129_,
		_w14130_
	);
	LUT2 #(
		.INIT('h1)
	) name13599 (
		\sa11_reg[2]/P0001 ,
		_w14130_,
		_w14131_
	);
	LUT2 #(
		.INIT('h4)
	) name13600 (
		_w12119_,
		_w12167_,
		_w14132_
	);
	LUT2 #(
		.INIT('h4)
	) name13601 (
		_w14127_,
		_w14132_,
		_w14133_
	);
	LUT2 #(
		.INIT('h4)
	) name13602 (
		_w14131_,
		_w14133_,
		_w14134_
	);
	LUT2 #(
		.INIT('h2)
	) name13603 (
		\sa11_reg[1]/P0001 ,
		_w14134_,
		_w14135_
	);
	LUT2 #(
		.INIT('h1)
	) name13604 (
		_w11836_,
		_w11913_,
		_w14136_
	);
	LUT2 #(
		.INIT('h2)
	) name13605 (
		\sa11_reg[2]/P0001 ,
		_w14136_,
		_w14137_
	);
	LUT2 #(
		.INIT('h8)
	) name13606 (
		_w11813_,
		_w11858_,
		_w14138_
	);
	LUT2 #(
		.INIT('h1)
	) name13607 (
		_w13101_,
		_w13159_,
		_w14139_
	);
	LUT2 #(
		.INIT('h1)
	) name13608 (
		\sa11_reg[2]/P0001 ,
		_w14139_,
		_w14140_
	);
	LUT2 #(
		.INIT('h1)
	) name13609 (
		_w11934_,
		_w14138_,
		_w14141_
	);
	LUT2 #(
		.INIT('h4)
	) name13610 (
		_w14137_,
		_w14141_,
		_w14142_
	);
	LUT2 #(
		.INIT('h4)
	) name13611 (
		_w14140_,
		_w14142_,
		_w14143_
	);
	LUT2 #(
		.INIT('h1)
	) name13612 (
		\sa11_reg[1]/P0001 ,
		_w14143_,
		_w14144_
	);
	LUT2 #(
		.INIT('h1)
	) name13613 (
		_w11934_,
		_w12176_,
		_w14145_
	);
	LUT2 #(
		.INIT('h1)
	) name13614 (
		\sa11_reg[2]/P0001 ,
		_w14145_,
		_w14146_
	);
	LUT2 #(
		.INIT('h1)
	) name13615 (
		_w13092_,
		_w13389_,
		_w14147_
	);
	LUT2 #(
		.INIT('h2)
	) name13616 (
		_w11805_,
		_w14147_,
		_w14148_
	);
	LUT2 #(
		.INIT('h1)
	) name13617 (
		_w11865_,
		_w12205_,
		_w14149_
	);
	LUT2 #(
		.INIT('h4)
	) name13618 (
		_w14148_,
		_w14149_,
		_w14150_
	);
	LUT2 #(
		.INIT('h4)
	) name13619 (
		_w14146_,
		_w14150_,
		_w14151_
	);
	LUT2 #(
		.INIT('h4)
	) name13620 (
		_w14135_,
		_w14151_,
		_w14152_
	);
	LUT2 #(
		.INIT('h4)
	) name13621 (
		_w14144_,
		_w14152_,
		_w14153_
	);
	LUT2 #(
		.INIT('h1)
	) name13622 (
		\sa11_reg[0]/P0001 ,
		_w14153_,
		_w14154_
	);
	LUT2 #(
		.INIT('h8)
	) name13623 (
		_w12126_,
		_w12127_,
		_w14155_
	);
	LUT2 #(
		.INIT('h1)
	) name13624 (
		_w12139_,
		_w14155_,
		_w14156_
	);
	LUT2 #(
		.INIT('h1)
	) name13625 (
		_w11886_,
		_w12127_,
		_w14157_
	);
	LUT2 #(
		.INIT('h1)
	) name13626 (
		\sa11_reg[5]/P0001 ,
		_w14157_,
		_w14158_
	);
	LUT2 #(
		.INIT('h8)
	) name13627 (
		\sa11_reg[3]/P0001 ,
		_w11821_,
		_w14159_
	);
	LUT2 #(
		.INIT('h1)
	) name13628 (
		_w14158_,
		_w14159_,
		_w14160_
	);
	LUT2 #(
		.INIT('h2)
	) name13629 (
		\sa11_reg[2]/P0001 ,
		_w14160_,
		_w14161_
	);
	LUT2 #(
		.INIT('h2)
	) name13630 (
		_w14156_,
		_w14161_,
		_w14162_
	);
	LUT2 #(
		.INIT('h2)
	) name13631 (
		\sa11_reg[1]/P0001 ,
		_w14162_,
		_w14163_
	);
	LUT2 #(
		.INIT('h8)
	) name13632 (
		\sa11_reg[4]/P0001 ,
		_w11847_,
		_w14164_
	);
	LUT2 #(
		.INIT('h1)
	) name13633 (
		_w11836_,
		_w11854_,
		_w14165_
	);
	LUT2 #(
		.INIT('h1)
	) name13634 (
		_w13513_,
		_w14164_,
		_w14166_
	);
	LUT2 #(
		.INIT('h8)
	) name13635 (
		_w14165_,
		_w14166_,
		_w14167_
	);
	LUT2 #(
		.INIT('h1)
	) name13636 (
		\sa11_reg[2]/P0001 ,
		_w14167_,
		_w14168_
	);
	LUT2 #(
		.INIT('h2)
	) name13637 (
		_w11822_,
		_w11893_,
		_w14169_
	);
	LUT2 #(
		.INIT('h4)
	) name13638 (
		\sa11_reg[1]/P0001 ,
		_w13102_,
		_w14170_
	);
	LUT2 #(
		.INIT('h1)
	) name13639 (
		_w14164_,
		_w14169_,
		_w14171_
	);
	LUT2 #(
		.INIT('h4)
	) name13640 (
		_w14170_,
		_w14171_,
		_w14172_
	);
	LUT2 #(
		.INIT('h1)
	) name13641 (
		\sa11_reg[3]/P0001 ,
		_w14172_,
		_w14173_
	);
	LUT2 #(
		.INIT('h2)
	) name13642 (
		_w11794_,
		_w11812_,
		_w14174_
	);
	LUT2 #(
		.INIT('h4)
	) name13643 (
		_w11821_,
		_w14174_,
		_w14175_
	);
	LUT2 #(
		.INIT('h1)
	) name13644 (
		_w11854_,
		_w12121_,
		_w14176_
	);
	LUT2 #(
		.INIT('h4)
	) name13645 (
		_w14175_,
		_w14176_,
		_w14177_
	);
	LUT2 #(
		.INIT('h1)
	) name13646 (
		\sa11_reg[1]/P0001 ,
		_w14177_,
		_w14178_
	);
	LUT2 #(
		.INIT('h1)
	) name13647 (
		_w14168_,
		_w14173_,
		_w14179_
	);
	LUT2 #(
		.INIT('h4)
	) name13648 (
		_w14178_,
		_w14179_,
		_w14180_
	);
	LUT2 #(
		.INIT('h4)
	) name13649 (
		_w14163_,
		_w14180_,
		_w14181_
	);
	LUT2 #(
		.INIT('h2)
	) name13650 (
		\sa11_reg[0]/P0001 ,
		_w14181_,
		_w14182_
	);
	LUT2 #(
		.INIT('h1)
	) name13651 (
		_w13109_,
		_w13509_,
		_w14183_
	);
	LUT2 #(
		.INIT('h4)
	) name13652 (
		_w11879_,
		_w14183_,
		_w14184_
	);
	LUT2 #(
		.INIT('h1)
	) name13653 (
		\sa11_reg[2]/P0001 ,
		_w14184_,
		_w14185_
	);
	LUT2 #(
		.INIT('h1)
	) name13654 (
		_w11927_,
		_w12177_,
		_w14186_
	);
	LUT2 #(
		.INIT('h4)
	) name13655 (
		_w14185_,
		_w14186_,
		_w14187_
	);
	LUT2 #(
		.INIT('h1)
	) name13656 (
		\sa11_reg[1]/P0001 ,
		_w14187_,
		_w14188_
	);
	LUT2 #(
		.INIT('h8)
	) name13657 (
		\sa11_reg[4]/P0001 ,
		_w13450_,
		_w14189_
	);
	LUT2 #(
		.INIT('h1)
	) name13658 (
		_w12128_,
		_w12139_,
		_w14190_
	);
	LUT2 #(
		.INIT('h2)
	) name13659 (
		\sa11_reg[3]/P0001 ,
		_w14190_,
		_w14191_
	);
	LUT2 #(
		.INIT('h1)
	) name13660 (
		_w13132_,
		_w14191_,
		_w14192_
	);
	LUT2 #(
		.INIT('h2)
	) name13661 (
		_w13171_,
		_w14192_,
		_w14193_
	);
	LUT2 #(
		.INIT('h8)
	) name13662 (
		_w11797_,
		_w11860_,
		_w14194_
	);
	LUT2 #(
		.INIT('h1)
	) name13663 (
		_w12151_,
		_w13093_,
		_w14195_
	);
	LUT2 #(
		.INIT('h4)
	) name13664 (
		_w14194_,
		_w14195_,
		_w14196_
	);
	LUT2 #(
		.INIT('h4)
	) name13665 (
		_w11922_,
		_w14196_,
		_w14197_
	);
	LUT2 #(
		.INIT('h2)
	) name13666 (
		_w13166_,
		_w14197_,
		_w14198_
	);
	LUT2 #(
		.INIT('h1)
	) name13667 (
		_w11834_,
		_w12222_,
		_w14199_
	);
	LUT2 #(
		.INIT('h8)
	) name13668 (
		_w12119_,
		_w14199_,
		_w14200_
	);
	LUT2 #(
		.INIT('h1)
	) name13669 (
		_w11865_,
		_w12186_,
		_w14201_
	);
	LUT2 #(
		.INIT('h4)
	) name13670 (
		_w13394_,
		_w14201_,
		_w14202_
	);
	LUT2 #(
		.INIT('h2)
	) name13671 (
		_w13544_,
		_w14202_,
		_w14203_
	);
	LUT2 #(
		.INIT('h1)
	) name13672 (
		_w14189_,
		_w14200_,
		_w14204_
	);
	LUT2 #(
		.INIT('h4)
	) name13673 (
		_w14193_,
		_w14204_,
		_w14205_
	);
	LUT2 #(
		.INIT('h1)
	) name13674 (
		_w14198_,
		_w14203_,
		_w14206_
	);
	LUT2 #(
		.INIT('h8)
	) name13675 (
		_w14205_,
		_w14206_,
		_w14207_
	);
	LUT2 #(
		.INIT('h4)
	) name13676 (
		_w14188_,
		_w14207_,
		_w14208_
	);
	LUT2 #(
		.INIT('h4)
	) name13677 (
		_w14182_,
		_w14208_,
		_w14209_
	);
	LUT2 #(
		.INIT('h4)
	) name13678 (
		_w14154_,
		_w14209_,
		_w14210_
	);
	LUT2 #(
		.INIT('h2)
	) name13679 (
		_w13649_,
		_w14210_,
		_w14211_
	);
	LUT2 #(
		.INIT('h4)
	) name13680 (
		_w13649_,
		_w14210_,
		_w14212_
	);
	LUT2 #(
		.INIT('h1)
	) name13681 (
		_w14211_,
		_w14212_,
		_w14213_
	);
	LUT2 #(
		.INIT('h4)
	) name13682 (
		_w14125_,
		_w14213_,
		_w14214_
	);
	LUT2 #(
		.INIT('h2)
	) name13683 (
		_w14125_,
		_w14213_,
		_w14215_
	);
	LUT2 #(
		.INIT('h1)
	) name13684 (
		_w14214_,
		_w14215_,
		_w14216_
	);
	LUT2 #(
		.INIT('h1)
	) name13685 (
		_w14122_,
		_w14216_,
		_w14217_
	);
	LUT2 #(
		.INIT('h8)
	) name13686 (
		_w14122_,
		_w14216_,
		_w14218_
	);
	LUT2 #(
		.INIT('h1)
	) name13687 (
		\ld_r_reg/P0001 ,
		_w14217_,
		_w14219_
	);
	LUT2 #(
		.INIT('h4)
	) name13688 (
		_w14218_,
		_w14219_,
		_w14220_
	);
	LUT2 #(
		.INIT('h1)
	) name13689 (
		\text_in_r_reg[105]/P0001 ,
		\u0_w_reg[0][9]/P0001 ,
		_w14221_
	);
	LUT2 #(
		.INIT('h8)
	) name13690 (
		\text_in_r_reg[105]/P0001 ,
		\u0_w_reg[0][9]/P0001 ,
		_w14222_
	);
	LUT2 #(
		.INIT('h2)
	) name13691 (
		\ld_r_reg/P0001 ,
		_w14221_,
		_w14223_
	);
	LUT2 #(
		.INIT('h4)
	) name13692 (
		_w14222_,
		_w14223_,
		_w14224_
	);
	LUT2 #(
		.INIT('h1)
	) name13693 (
		_w14220_,
		_w14224_,
		_w14225_
	);
	LUT2 #(
		.INIT('h2)
	) name13694 (
		\u0_w_reg[0][1]/P0001 ,
		_w13835_,
		_w14226_
	);
	LUT2 #(
		.INIT('h4)
	) name13695 (
		\u0_w_reg[0][1]/P0001 ,
		_w13835_,
		_w14227_
	);
	LUT2 #(
		.INIT('h1)
	) name13696 (
		_w14226_,
		_w14227_,
		_w14228_
	);
	LUT2 #(
		.INIT('h8)
	) name13697 (
		_w14116_,
		_w14228_,
		_w14229_
	);
	LUT2 #(
		.INIT('h1)
	) name13698 (
		_w14116_,
		_w14228_,
		_w14230_
	);
	LUT2 #(
		.INIT('h1)
	) name13699 (
		_w14229_,
		_w14230_,
		_w14231_
	);
	LUT2 #(
		.INIT('h4)
	) name13700 (
		\sa00_reg[2]/P0001 ,
		_w11957_,
		_w14232_
	);
	LUT2 #(
		.INIT('h1)
	) name13701 (
		_w12072_,
		_w13068_,
		_w14233_
	);
	LUT2 #(
		.INIT('h4)
	) name13702 (
		_w14232_,
		_w14233_,
		_w14234_
	);
	LUT2 #(
		.INIT('h2)
	) name13703 (
		\sa00_reg[1]/P0001 ,
		_w14234_,
		_w14235_
	);
	LUT2 #(
		.INIT('h4)
	) name13704 (
		_w12654_,
		_w13044_,
		_w14236_
	);
	LUT2 #(
		.INIT('h8)
	) name13705 (
		_w11959_,
		_w11995_,
		_w14237_
	);
	LUT2 #(
		.INIT('h1)
	) name13706 (
		_w13031_,
		_w14237_,
		_w14238_
	);
	LUT2 #(
		.INIT('h1)
	) name13707 (
		\sa00_reg[2]/P0001 ,
		_w14238_,
		_w14239_
	);
	LUT2 #(
		.INIT('h8)
	) name13708 (
		_w11959_,
		_w13629_,
		_w14240_
	);
	LUT2 #(
		.INIT('h1)
	) name13709 (
		_w12091_,
		_w14240_,
		_w14241_
	);
	LUT2 #(
		.INIT('h8)
	) name13710 (
		_w13013_,
		_w14241_,
		_w14242_
	);
	LUT2 #(
		.INIT('h2)
	) name13711 (
		\sa00_reg[2]/P0001 ,
		_w14242_,
		_w14243_
	);
	LUT2 #(
		.INIT('h2)
	) name13712 (
		\sa00_reg[5]/P0001 ,
		_w11952_,
		_w14244_
	);
	LUT2 #(
		.INIT('h2)
	) name13713 (
		_w11966_,
		_w14244_,
		_w14245_
	);
	LUT2 #(
		.INIT('h1)
	) name13714 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		_w14246_
	);
	LUT2 #(
		.INIT('h8)
	) name13715 (
		_w11961_,
		_w14246_,
		_w14247_
	);
	LUT2 #(
		.INIT('h8)
	) name13716 (
		_w12005_,
		_w12026_,
		_w14248_
	);
	LUT2 #(
		.INIT('h4)
	) name13717 (
		\sa00_reg[5]/P0001 ,
		_w12015_,
		_w14249_
	);
	LUT2 #(
		.INIT('h1)
	) name13718 (
		_w12605_,
		_w12692_,
		_w14250_
	);
	LUT2 #(
		.INIT('h4)
	) name13719 (
		_w14249_,
		_w14250_,
		_w14251_
	);
	LUT2 #(
		.INIT('h2)
	) name13720 (
		\sa00_reg[2]/P0001 ,
		_w14251_,
		_w14252_
	);
	LUT2 #(
		.INIT('h1)
	) name13721 (
		_w14245_,
		_w14248_,
		_w14253_
	);
	LUT2 #(
		.INIT('h4)
	) name13722 (
		_w14247_,
		_w14253_,
		_w14254_
	);
	LUT2 #(
		.INIT('h4)
	) name13723 (
		_w14252_,
		_w14254_,
		_w14255_
	);
	LUT2 #(
		.INIT('h1)
	) name13724 (
		\sa00_reg[1]/P0001 ,
		_w14255_,
		_w14256_
	);
	LUT2 #(
		.INIT('h1)
	) name13725 (
		_w12053_,
		_w13575_,
		_w14257_
	);
	LUT2 #(
		.INIT('h4)
	) name13726 (
		_w14236_,
		_w14257_,
		_w14258_
	);
	LUT2 #(
		.INIT('h4)
	) name13727 (
		_w14239_,
		_w14258_,
		_w14259_
	);
	LUT2 #(
		.INIT('h4)
	) name13728 (
		_w14235_,
		_w14259_,
		_w14260_
	);
	LUT2 #(
		.INIT('h4)
	) name13729 (
		_w14243_,
		_w14260_,
		_w14261_
	);
	LUT2 #(
		.INIT('h4)
	) name13730 (
		_w14256_,
		_w14261_,
		_w14262_
	);
	LUT2 #(
		.INIT('h2)
	) name13731 (
		\sa00_reg[0]/P0001 ,
		_w14262_,
		_w14263_
	);
	LUT2 #(
		.INIT('h4)
	) name13732 (
		\sa00_reg[4]/P0001 ,
		_w11996_,
		_w14264_
	);
	LUT2 #(
		.INIT('h1)
	) name13733 (
		_w12066_,
		_w14264_,
		_w14265_
	);
	LUT2 #(
		.INIT('h1)
	) name13734 (
		\sa00_reg[3]/P0001 ,
		_w14265_,
		_w14266_
	);
	LUT2 #(
		.INIT('h1)
	) name13735 (
		_w11984_,
		_w14266_,
		_w14267_
	);
	LUT2 #(
		.INIT('h1)
	) name13736 (
		\sa00_reg[1]/P0001 ,
		_w14267_,
		_w14268_
	);
	LUT2 #(
		.INIT('h8)
	) name13737 (
		\sa00_reg[6]/NET0131 ,
		_w11974_,
		_w14269_
	);
	LUT2 #(
		.INIT('h1)
	) name13738 (
		_w14240_,
		_w14269_,
		_w14270_
	);
	LUT2 #(
		.INIT('h4)
	) name13739 (
		_w13038_,
		_w14270_,
		_w14271_
	);
	LUT2 #(
		.INIT('h1)
	) name13740 (
		\sa00_reg[2]/P0001 ,
		_w14271_,
		_w14272_
	);
	LUT2 #(
		.INIT('h1)
	) name13741 (
		_w11967_,
		_w12035_,
		_w14273_
	);
	LUT2 #(
		.INIT('h2)
	) name13742 (
		_w12596_,
		_w14273_,
		_w14274_
	);
	LUT2 #(
		.INIT('h2)
	) name13743 (
		_w11973_,
		_w11979_,
		_w14275_
	);
	LUT2 #(
		.INIT('h8)
	) name13744 (
		_w13015_,
		_w14275_,
		_w14276_
	);
	LUT2 #(
		.INIT('h8)
	) name13745 (
		_w12096_,
		_w14246_,
		_w14277_
	);
	LUT2 #(
		.INIT('h8)
	) name13746 (
		\sa00_reg[3]/P0001 ,
		_w12095_,
		_w14278_
	);
	LUT2 #(
		.INIT('h8)
	) name13747 (
		_w11982_,
		_w12002_,
		_w14279_
	);
	LUT2 #(
		.INIT('h1)
	) name13748 (
		_w12015_,
		_w12636_,
		_w14280_
	);
	LUT2 #(
		.INIT('h1)
	) name13749 (
		_w14277_,
		_w14279_,
		_w14281_
	);
	LUT2 #(
		.INIT('h8)
	) name13750 (
		_w14280_,
		_w14281_,
		_w14282_
	);
	LUT2 #(
		.INIT('h4)
	) name13751 (
		_w14278_,
		_w14282_,
		_w14283_
	);
	LUT2 #(
		.INIT('h2)
	) name13752 (
		\sa00_reg[1]/P0001 ,
		_w14283_,
		_w14284_
	);
	LUT2 #(
		.INIT('h1)
	) name13753 (
		_w14274_,
		_w14276_,
		_w14285_
	);
	LUT2 #(
		.INIT('h4)
	) name13754 (
		_w14272_,
		_w14285_,
		_w14286_
	);
	LUT2 #(
		.INIT('h4)
	) name13755 (
		_w14284_,
		_w14286_,
		_w14287_
	);
	LUT2 #(
		.INIT('h4)
	) name13756 (
		_w14268_,
		_w14287_,
		_w14288_
	);
	LUT2 #(
		.INIT('h1)
	) name13757 (
		\sa00_reg[0]/P0001 ,
		_w14288_,
		_w14289_
	);
	LUT2 #(
		.INIT('h4)
	) name13758 (
		\sa00_reg[4]/P0001 ,
		_w12026_,
		_w14290_
	);
	LUT2 #(
		.INIT('h8)
	) name13759 (
		_w12056_,
		_w14290_,
		_w14291_
	);
	LUT2 #(
		.INIT('h1)
	) name13760 (
		_w13045_,
		_w14291_,
		_w14292_
	);
	LUT2 #(
		.INIT('h2)
	) name13761 (
		\sa00_reg[6]/NET0131 ,
		_w14292_,
		_w14293_
	);
	LUT2 #(
		.INIT('h1)
	) name13762 (
		_w11993_,
		_w12637_,
		_w14294_
	);
	LUT2 #(
		.INIT('h2)
	) name13763 (
		\sa00_reg[2]/P0001 ,
		_w14294_,
		_w14295_
	);
	LUT2 #(
		.INIT('h8)
	) name13764 (
		_w12632_,
		_w14246_,
		_w14296_
	);
	LUT2 #(
		.INIT('h1)
	) name13765 (
		_w11968_,
		_w12006_,
		_w14297_
	);
	LUT2 #(
		.INIT('h4)
	) name13766 (
		_w14296_,
		_w14297_,
		_w14298_
	);
	LUT2 #(
		.INIT('h4)
	) name13767 (
		_w14295_,
		_w14298_,
		_w14299_
	);
	LUT2 #(
		.INIT('h2)
	) name13768 (
		\sa00_reg[1]/P0001 ,
		_w14299_,
		_w14300_
	);
	LUT2 #(
		.INIT('h4)
	) name13769 (
		\sa00_reg[3]/P0001 ,
		_w11962_,
		_w14301_
	);
	LUT2 #(
		.INIT('h4)
	) name13770 (
		_w12014_,
		_w14301_,
		_w14302_
	);
	LUT2 #(
		.INIT('h1)
	) name13771 (
		_w12016_,
		_w14302_,
		_w14303_
	);
	LUT2 #(
		.INIT('h1)
	) name13772 (
		\sa00_reg[2]/P0001 ,
		_w14303_,
		_w14304_
	);
	LUT2 #(
		.INIT('h8)
	) name13773 (
		\sa00_reg[2]/P0001 ,
		_w12005_,
		_w14305_
	);
	LUT2 #(
		.INIT('h1)
	) name13774 (
		_w11995_,
		_w12685_,
		_w14306_
	);
	LUT2 #(
		.INIT('h2)
	) name13775 (
		_w14305_,
		_w14306_,
		_w14307_
	);
	LUT2 #(
		.INIT('h8)
	) name13776 (
		_w13006_,
		_w13044_,
		_w14308_
	);
	LUT2 #(
		.INIT('h1)
	) name13777 (
		_w12702_,
		_w14308_,
		_w14309_
	);
	LUT2 #(
		.INIT('h4)
	) name13778 (
		_w14307_,
		_w14309_,
		_w14310_
	);
	LUT2 #(
		.INIT('h4)
	) name13779 (
		_w14304_,
		_w14310_,
		_w14311_
	);
	LUT2 #(
		.INIT('h1)
	) name13780 (
		\sa00_reg[1]/P0001 ,
		_w14311_,
		_w14312_
	);
	LUT2 #(
		.INIT('h1)
	) name13781 (
		_w14293_,
		_w14300_,
		_w14313_
	);
	LUT2 #(
		.INIT('h4)
	) name13782 (
		_w14312_,
		_w14313_,
		_w14314_
	);
	LUT2 #(
		.INIT('h4)
	) name13783 (
		_w14263_,
		_w14314_,
		_w14315_
	);
	LUT2 #(
		.INIT('h4)
	) name13784 (
		_w14289_,
		_w14315_,
		_w14316_
	);
	LUT2 #(
		.INIT('h1)
	) name13785 (
		_w12630_,
		_w14237_,
		_w14317_
	);
	LUT2 #(
		.INIT('h4)
	) name13786 (
		_w13610_,
		_w14317_,
		_w14318_
	);
	LUT2 #(
		.INIT('h2)
	) name13787 (
		_w12054_,
		_w14318_,
		_w14319_
	);
	LUT2 #(
		.INIT('h1)
	) name13788 (
		_w11956_,
		_w12050_,
		_w14320_
	);
	LUT2 #(
		.INIT('h2)
	) name13789 (
		_w13004_,
		_w14320_,
		_w14321_
	);
	LUT2 #(
		.INIT('h4)
	) name13790 (
		\sa00_reg[2]/P0001 ,
		_w11978_,
		_w14322_
	);
	LUT2 #(
		.INIT('h1)
	) name13791 (
		_w13012_,
		_w14322_,
		_w14323_
	);
	LUT2 #(
		.INIT('h4)
	) name13792 (
		_w14321_,
		_w14323_,
		_w14324_
	);
	LUT2 #(
		.INIT('h1)
	) name13793 (
		\sa00_reg[1]/P0001 ,
		_w14324_,
		_w14325_
	);
	LUT2 #(
		.INIT('h1)
	) name13794 (
		_w13572_,
		_w14248_,
		_w14326_
	);
	LUT2 #(
		.INIT('h1)
	) name13795 (
		_w12018_,
		_w13062_,
		_w14327_
	);
	LUT2 #(
		.INIT('h8)
	) name13796 (
		_w14326_,
		_w14327_,
		_w14328_
	);
	LUT2 #(
		.INIT('h1)
	) name13797 (
		\sa00_reg[2]/P0001 ,
		_w14328_,
		_w14329_
	);
	LUT2 #(
		.INIT('h2)
	) name13798 (
		\sa00_reg[2]/P0001 ,
		_w12036_,
		_w14330_
	);
	LUT2 #(
		.INIT('h4)
	) name13799 (
		_w12666_,
		_w13639_,
		_w14331_
	);
	LUT2 #(
		.INIT('h1)
	) name13800 (
		_w14330_,
		_w14331_,
		_w14332_
	);
	LUT2 #(
		.INIT('h1)
	) name13801 (
		_w13037_,
		_w13069_,
		_w14333_
	);
	LUT2 #(
		.INIT('h4)
	) name13802 (
		_w14332_,
		_w14333_,
		_w14334_
	);
	LUT2 #(
		.INIT('h2)
	) name13803 (
		\sa00_reg[1]/P0001 ,
		_w14334_,
		_w14335_
	);
	LUT2 #(
		.INIT('h1)
	) name13804 (
		_w14319_,
		_w14325_,
		_w14336_
	);
	LUT2 #(
		.INIT('h4)
	) name13805 (
		_w14329_,
		_w14336_,
		_w14337_
	);
	LUT2 #(
		.INIT('h4)
	) name13806 (
		_w14335_,
		_w14337_,
		_w14338_
	);
	LUT2 #(
		.INIT('h1)
	) name13807 (
		\sa00_reg[0]/P0001 ,
		_w14338_,
		_w14339_
	);
	LUT2 #(
		.INIT('h8)
	) name13808 (
		\sa00_reg[3]/P0001 ,
		_w11962_,
		_w14340_
	);
	LUT2 #(
		.INIT('h1)
	) name13809 (
		_w12015_,
		_w12065_,
		_w14341_
	);
	LUT2 #(
		.INIT('h1)
	) name13810 (
		_w13028_,
		_w14340_,
		_w14342_
	);
	LUT2 #(
		.INIT('h8)
	) name13811 (
		_w14341_,
		_w14342_,
		_w14343_
	);
	LUT2 #(
		.INIT('h2)
	) name13812 (
		\sa00_reg[1]/P0001 ,
		_w14343_,
		_w14344_
	);
	LUT2 #(
		.INIT('h1)
	) name13813 (
		_w12045_,
		_w12614_,
		_w14345_
	);
	LUT2 #(
		.INIT('h4)
	) name13814 (
		_w12605_,
		_w14345_,
		_w14346_
	);
	LUT2 #(
		.INIT('h4)
	) name13815 (
		_w14344_,
		_w14346_,
		_w14347_
	);
	LUT2 #(
		.INIT('h2)
	) name13816 (
		\sa00_reg[2]/P0001 ,
		_w14347_,
		_w14348_
	);
	LUT2 #(
		.INIT('h8)
	) name13817 (
		_w12054_,
		_w12082_,
		_w14349_
	);
	LUT2 #(
		.INIT('h8)
	) name13818 (
		_w12685_,
		_w14246_,
		_w14350_
	);
	LUT2 #(
		.INIT('h1)
	) name13819 (
		_w12051_,
		_w14350_,
		_w14351_
	);
	LUT2 #(
		.INIT('h2)
	) name13820 (
		\sa00_reg[1]/P0001 ,
		_w14351_,
		_w14352_
	);
	LUT2 #(
		.INIT('h8)
	) name13821 (
		_w12086_,
		_w14301_,
		_w14353_
	);
	LUT2 #(
		.INIT('h1)
	) name13822 (
		_w12057_,
		_w12068_,
		_w14354_
	);
	LUT2 #(
		.INIT('h1)
	) name13823 (
		_w13028_,
		_w14301_,
		_w14355_
	);
	LUT2 #(
		.INIT('h8)
	) name13824 (
		_w14354_,
		_w14355_,
		_w14356_
	);
	LUT2 #(
		.INIT('h1)
	) name13825 (
		\sa00_reg[2]/P0001 ,
		_w14356_,
		_w14357_
	);
	LUT2 #(
		.INIT('h1)
	) name13826 (
		_w12072_,
		_w13036_,
		_w14358_
	);
	LUT2 #(
		.INIT('h1)
	) name13827 (
		\sa00_reg[7]/NET0131 ,
		_w14358_,
		_w14359_
	);
	LUT2 #(
		.INIT('h8)
	) name13828 (
		_w12056_,
		_w12090_,
		_w14360_
	);
	LUT2 #(
		.INIT('h1)
	) name13829 (
		_w12019_,
		_w14360_,
		_w14361_
	);
	LUT2 #(
		.INIT('h4)
	) name13830 (
		_w14359_,
		_w14361_,
		_w14362_
	);
	LUT2 #(
		.INIT('h4)
	) name13831 (
		_w14357_,
		_w14362_,
		_w14363_
	);
	LUT2 #(
		.INIT('h1)
	) name13832 (
		\sa00_reg[1]/P0001 ,
		_w14363_,
		_w14364_
	);
	LUT2 #(
		.INIT('h1)
	) name13833 (
		_w13031_,
		_w14349_,
		_w14365_
	);
	LUT2 #(
		.INIT('h4)
	) name13834 (
		_w14353_,
		_w14365_,
		_w14366_
	);
	LUT2 #(
		.INIT('h4)
	) name13835 (
		_w14352_,
		_w14366_,
		_w14367_
	);
	LUT2 #(
		.INIT('h4)
	) name13836 (
		_w14348_,
		_w14367_,
		_w14368_
	);
	LUT2 #(
		.INIT('h4)
	) name13837 (
		_w14364_,
		_w14368_,
		_w14369_
	);
	LUT2 #(
		.INIT('h2)
	) name13838 (
		\sa00_reg[0]/P0001 ,
		_w14369_,
		_w14370_
	);
	LUT2 #(
		.INIT('h8)
	) name13839 (
		_w11956_,
		_w12014_,
		_w14371_
	);
	LUT2 #(
		.INIT('h1)
	) name13840 (
		_w11961_,
		_w13074_,
		_w14372_
	);
	LUT2 #(
		.INIT('h4)
	) name13841 (
		_w14371_,
		_w14372_,
		_w14373_
	);
	LUT2 #(
		.INIT('h1)
	) name13842 (
		\sa00_reg[3]/P0001 ,
		_w14373_,
		_w14374_
	);
	LUT2 #(
		.INIT('h1)
	) name13843 (
		_w12027_,
		_w12624_,
		_w14375_
	);
	LUT2 #(
		.INIT('h4)
	) name13844 (
		_w14374_,
		_w14375_,
		_w14376_
	);
	LUT2 #(
		.INIT('h2)
	) name13845 (
		\sa00_reg[2]/P0001 ,
		_w14376_,
		_w14377_
	);
	LUT2 #(
		.INIT('h2)
	) name13846 (
		_w11975_,
		_w11978_,
		_w14378_
	);
	LUT2 #(
		.INIT('h2)
	) name13847 (
		_w14265_,
		_w14378_,
		_w14379_
	);
	LUT2 #(
		.INIT('h2)
	) name13848 (
		_w13044_,
		_w14379_,
		_w14380_
	);
	LUT2 #(
		.INIT('h1)
	) name13849 (
		_w14377_,
		_w14380_,
		_w14381_
	);
	LUT2 #(
		.INIT('h2)
	) name13850 (
		\sa00_reg[1]/P0001 ,
		_w14381_,
		_w14382_
	);
	LUT2 #(
		.INIT('h8)
	) name13851 (
		_w11962_,
		_w12693_,
		_w14383_
	);
	LUT2 #(
		.INIT('h1)
	) name13852 (
		_w12081_,
		_w14383_,
		_w14384_
	);
	LUT2 #(
		.INIT('h1)
	) name13853 (
		\sa00_reg[2]/P0001 ,
		_w14384_,
		_w14385_
	);
	LUT2 #(
		.INIT('h8)
	) name13854 (
		\sa00_reg[5]/P0001 ,
		_w13036_,
		_w14386_
	);
	LUT2 #(
		.INIT('h1)
	) name13855 (
		_w12051_,
		_w12611_,
		_w14387_
	);
	LUT2 #(
		.INIT('h4)
	) name13856 (
		_w14386_,
		_w14387_,
		_w14388_
	);
	LUT2 #(
		.INIT('h2)
	) name13857 (
		_w13015_,
		_w14388_,
		_w14389_
	);
	LUT2 #(
		.INIT('h8)
	) name13858 (
		_w11955_,
		_w11973_,
		_w14390_
	);
	LUT2 #(
		.INIT('h2)
	) name13859 (
		\sa00_reg[2]/P0001 ,
		_w14390_,
		_w14391_
	);
	LUT2 #(
		.INIT('h1)
	) name13860 (
		_w12052_,
		_w14390_,
		_w14392_
	);
	LUT2 #(
		.INIT('h8)
	) name13861 (
		_w14326_,
		_w14392_,
		_w14393_
	);
	LUT2 #(
		.INIT('h1)
	) name13862 (
		\sa00_reg[1]/P0001 ,
		_w14391_,
		_w14394_
	);
	LUT2 #(
		.INIT('h4)
	) name13863 (
		_w14393_,
		_w14394_,
		_w14395_
	);
	LUT2 #(
		.INIT('h1)
	) name13864 (
		_w14385_,
		_w14389_,
		_w14396_
	);
	LUT2 #(
		.INIT('h4)
	) name13865 (
		_w14395_,
		_w14396_,
		_w14397_
	);
	LUT2 #(
		.INIT('h4)
	) name13866 (
		_w14382_,
		_w14397_,
		_w14398_
	);
	LUT2 #(
		.INIT('h4)
	) name13867 (
		_w14339_,
		_w14398_,
		_w14399_
	);
	LUT2 #(
		.INIT('h4)
	) name13868 (
		_w14370_,
		_w14399_,
		_w14400_
	);
	LUT2 #(
		.INIT('h2)
	) name13869 (
		_w14316_,
		_w14400_,
		_w14401_
	);
	LUT2 #(
		.INIT('h4)
	) name13870 (
		_w14316_,
		_w14400_,
		_w14402_
	);
	LUT2 #(
		.INIT('h1)
	) name13871 (
		_w14401_,
		_w14402_,
		_w14403_
	);
	LUT2 #(
		.INIT('h4)
	) name13872 (
		_w14213_,
		_w14403_,
		_w14404_
	);
	LUT2 #(
		.INIT('h2)
	) name13873 (
		_w14213_,
		_w14403_,
		_w14405_
	);
	LUT2 #(
		.INIT('h1)
	) name13874 (
		_w14404_,
		_w14405_,
		_w14406_
	);
	LUT2 #(
		.INIT('h1)
	) name13875 (
		_w14231_,
		_w14406_,
		_w14407_
	);
	LUT2 #(
		.INIT('h8)
	) name13876 (
		_w14231_,
		_w14406_,
		_w14408_
	);
	LUT2 #(
		.INIT('h1)
	) name13877 (
		\ld_r_reg/P0001 ,
		_w14407_,
		_w14409_
	);
	LUT2 #(
		.INIT('h4)
	) name13878 (
		_w14408_,
		_w14409_,
		_w14410_
	);
	LUT2 #(
		.INIT('h1)
	) name13879 (
		\text_in_r_reg[97]/P0001 ,
		\u0_w_reg[0][1]/P0001 ,
		_w14411_
	);
	LUT2 #(
		.INIT('h8)
	) name13880 (
		\text_in_r_reg[97]/P0001 ,
		\u0_w_reg[0][1]/P0001 ,
		_w14412_
	);
	LUT2 #(
		.INIT('h2)
	) name13881 (
		\ld_r_reg/P0001 ,
		_w14411_,
		_w14413_
	);
	LUT2 #(
		.INIT('h4)
	) name13882 (
		_w14412_,
		_w14413_,
		_w14414_
	);
	LUT2 #(
		.INIT('h1)
	) name13883 (
		_w14410_,
		_w14414_,
		_w14415_
	);
	LUT2 #(
		.INIT('h1)
	) name13884 (
		_w11935_,
		_w13509_,
		_w14416_
	);
	LUT2 #(
		.INIT('h1)
	) name13885 (
		\sa11_reg[2]/P0001 ,
		_w14416_,
		_w14417_
	);
	LUT2 #(
		.INIT('h1)
	) name13886 (
		_w11792_,
		_w12168_,
		_w14418_
	);
	LUT2 #(
		.INIT('h2)
	) name13887 (
		\sa11_reg[2]/P0001 ,
		_w14418_,
		_w14419_
	);
	LUT2 #(
		.INIT('h1)
	) name13888 (
		_w11865_,
		_w12124_,
		_w14420_
	);
	LUT2 #(
		.INIT('h4)
	) name13889 (
		_w11927_,
		_w14420_,
		_w14421_
	);
	LUT2 #(
		.INIT('h4)
	) name13890 (
		_w13450_,
		_w14421_,
		_w14422_
	);
	LUT2 #(
		.INIT('h4)
	) name13891 (
		_w14419_,
		_w14422_,
		_w14423_
	);
	LUT2 #(
		.INIT('h4)
	) name13892 (
		_w14417_,
		_w14423_,
		_w14424_
	);
	LUT2 #(
		.INIT('h1)
	) name13893 (
		\sa11_reg[1]/P0001 ,
		_w14424_,
		_w14425_
	);
	LUT2 #(
		.INIT('h2)
	) name13894 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w14426_
	);
	LUT2 #(
		.INIT('h2)
	) name13895 (
		_w11797_,
		_w14426_,
		_w14427_
	);
	LUT2 #(
		.INIT('h1)
	) name13896 (
		_w11806_,
		_w14427_,
		_w14428_
	);
	LUT2 #(
		.INIT('h2)
	) name13897 (
		\sa11_reg[2]/P0001 ,
		_w14428_,
		_w14429_
	);
	LUT2 #(
		.INIT('h1)
	) name13898 (
		_w11913_,
		_w13473_,
		_w14430_
	);
	LUT2 #(
		.INIT('h4)
	) name13899 (
		_w11898_,
		_w14430_,
		_w14431_
	);
	LUT2 #(
		.INIT('h1)
	) name13900 (
		_w13390_,
		_w13447_,
		_w14432_
	);
	LUT2 #(
		.INIT('h8)
	) name13901 (
		_w14431_,
		_w14432_,
		_w14433_
	);
	LUT2 #(
		.INIT('h4)
	) name13902 (
		_w14429_,
		_w14433_,
		_w14434_
	);
	LUT2 #(
		.INIT('h2)
	) name13903 (
		\sa11_reg[1]/P0001 ,
		_w14434_,
		_w14435_
	);
	LUT2 #(
		.INIT('h8)
	) name13904 (
		_w11801_,
		_w11860_,
		_w14436_
	);
	LUT2 #(
		.INIT('h2)
	) name13905 (
		_w13421_,
		_w14436_,
		_w14437_
	);
	LUT2 #(
		.INIT('h1)
	) name13906 (
		\sa11_reg[2]/P0001 ,
		_w14437_,
		_w14438_
	);
	LUT2 #(
		.INIT('h4)
	) name13907 (
		_w12120_,
		_w12207_,
		_w14439_
	);
	LUT2 #(
		.INIT('h2)
	) name13908 (
		_w11834_,
		_w14439_,
		_w14440_
	);
	LUT2 #(
		.INIT('h1)
	) name13909 (
		_w12198_,
		_w14440_,
		_w14441_
	);
	LUT2 #(
		.INIT('h4)
	) name13910 (
		_w14438_,
		_w14441_,
		_w14442_
	);
	LUT2 #(
		.INIT('h4)
	) name13911 (
		_w14435_,
		_w14442_,
		_w14443_
	);
	LUT2 #(
		.INIT('h4)
	) name13912 (
		_w14425_,
		_w14443_,
		_w14444_
	);
	LUT2 #(
		.INIT('h2)
	) name13913 (
		\sa11_reg[0]/P0001 ,
		_w14444_,
		_w14445_
	);
	LUT2 #(
		.INIT('h8)
	) name13914 (
		_w11893_,
		_w11909_,
		_w14446_
	);
	LUT2 #(
		.INIT('h1)
	) name13915 (
		_w11882_,
		_w13102_,
		_w14447_
	);
	LUT2 #(
		.INIT('h4)
	) name13916 (
		_w13489_,
		_w14447_,
		_w14448_
	);
	LUT2 #(
		.INIT('h2)
	) name13917 (
		_w13106_,
		_w14448_,
		_w14449_
	);
	LUT2 #(
		.INIT('h1)
	) name13918 (
		_w11899_,
		_w14446_,
		_w14450_
	);
	LUT2 #(
		.INIT('h4)
	) name13919 (
		_w14449_,
		_w14450_,
		_w14451_
	);
	LUT2 #(
		.INIT('h2)
	) name13920 (
		\sa11_reg[1]/P0001 ,
		_w14451_,
		_w14452_
	);
	LUT2 #(
		.INIT('h1)
	) name13921 (
		_w11879_,
		_w12195_,
		_w14453_
	);
	LUT2 #(
		.INIT('h2)
	) name13922 (
		_w13544_,
		_w14453_,
		_w14454_
	);
	LUT2 #(
		.INIT('h1)
	) name13923 (
		_w11883_,
		_w12139_,
		_w14455_
	);
	LUT2 #(
		.INIT('h2)
	) name13924 (
		_w11846_,
		_w14455_,
		_w14456_
	);
	LUT2 #(
		.INIT('h8)
	) name13925 (
		_w11896_,
		_w12222_,
		_w14457_
	);
	LUT2 #(
		.INIT('h8)
	) name13926 (
		\sa11_reg[6]/NET0131 ,
		_w11923_,
		_w14458_
	);
	LUT2 #(
		.INIT('h1)
	) name13927 (
		_w11913_,
		_w14458_,
		_w14459_
	);
	LUT2 #(
		.INIT('h2)
	) name13928 (
		_w13171_,
		_w14459_,
		_w14460_
	);
	LUT2 #(
		.INIT('h4)
	) name13929 (
		\sa11_reg[2]/P0001 ,
		_w13096_,
		_w14461_
	);
	LUT2 #(
		.INIT('h8)
	) name13930 (
		_w11863_,
		_w13092_,
		_w14462_
	);
	LUT2 #(
		.INIT('h2)
	) name13931 (
		_w11908_,
		_w14462_,
		_w14463_
	);
	LUT2 #(
		.INIT('h1)
	) name13932 (
		_w14461_,
		_w14463_,
		_w14464_
	);
	LUT2 #(
		.INIT('h8)
	) name13933 (
		_w11797_,
		_w13502_,
		_w14465_
	);
	LUT2 #(
		.INIT('h1)
	) name13934 (
		_w12153_,
		_w13127_,
		_w14466_
	);
	LUT2 #(
		.INIT('h2)
	) name13935 (
		\sa11_reg[2]/P0001 ,
		_w14466_,
		_w14467_
	);
	LUT2 #(
		.INIT('h2)
	) name13936 (
		\sa11_reg[1]/P0001 ,
		_w11909_,
		_w14468_
	);
	LUT2 #(
		.INIT('h4)
	) name13937 (
		_w11862_,
		_w14468_,
		_w14469_
	);
	LUT2 #(
		.INIT('h1)
	) name13938 (
		_w14155_,
		_w14465_,
		_w14470_
	);
	LUT2 #(
		.INIT('h8)
	) name13939 (
		_w14469_,
		_w14470_,
		_w14471_
	);
	LUT2 #(
		.INIT('h4)
	) name13940 (
		_w14467_,
		_w14471_,
		_w14472_
	);
	LUT2 #(
		.INIT('h8)
	) name13941 (
		\sa11_reg[7]/NET0131 ,
		_w11805_,
		_w14473_
	);
	LUT2 #(
		.INIT('h4)
	) name13942 (
		_w11876_,
		_w14473_,
		_w14474_
	);
	LUT2 #(
		.INIT('h8)
	) name13943 (
		_w11829_,
		_w11834_,
		_w14475_
	);
	LUT2 #(
		.INIT('h1)
	) name13944 (
		\sa11_reg[1]/P0001 ,
		_w14436_,
		_w14476_
	);
	LUT2 #(
		.INIT('h4)
	) name13945 (
		_w14475_,
		_w14476_,
		_w14477_
	);
	LUT2 #(
		.INIT('h1)
	) name13946 (
		_w13172_,
		_w14474_,
		_w14478_
	);
	LUT2 #(
		.INIT('h8)
	) name13947 (
		_w14477_,
		_w14478_,
		_w14479_
	);
	LUT2 #(
		.INIT('h4)
	) name13948 (
		_w13170_,
		_w14479_,
		_w14480_
	);
	LUT2 #(
		.INIT('h1)
	) name13949 (
		_w14472_,
		_w14480_,
		_w14481_
	);
	LUT2 #(
		.INIT('h1)
	) name13950 (
		_w12195_,
		_w14464_,
		_w14482_
	);
	LUT2 #(
		.INIT('h4)
	) name13951 (
		_w14481_,
		_w14482_,
		_w14483_
	);
	LUT2 #(
		.INIT('h1)
	) name13952 (
		\sa11_reg[0]/P0001 ,
		_w14483_,
		_w14484_
	);
	LUT2 #(
		.INIT('h1)
	) name13953 (
		_w14138_,
		_w14457_,
		_w14485_
	);
	LUT2 #(
		.INIT('h4)
	) name13954 (
		_w14454_,
		_w14485_,
		_w14486_
	);
	LUT2 #(
		.INIT('h1)
	) name13955 (
		_w14456_,
		_w14460_,
		_w14487_
	);
	LUT2 #(
		.INIT('h8)
	) name13956 (
		_w14486_,
		_w14487_,
		_w14488_
	);
	LUT2 #(
		.INIT('h4)
	) name13957 (
		_w14452_,
		_w14488_,
		_w14489_
	);
	LUT2 #(
		.INIT('h4)
	) name13958 (
		_w14484_,
		_w14489_,
		_w14490_
	);
	LUT2 #(
		.INIT('h4)
	) name13959 (
		_w14445_,
		_w14490_,
		_w14491_
	);
	LUT2 #(
		.INIT('h4)
	) name13960 (
		_w12234_,
		_w12258_,
		_w14492_
	);
	LUT2 #(
		.INIT('h1)
	) name13961 (
		_w13268_,
		_w14492_,
		_w14493_
	);
	LUT2 #(
		.INIT('h2)
	) name13962 (
		\sa22_reg[2]/P0001 ,
		_w14493_,
		_w14494_
	);
	LUT2 #(
		.INIT('h8)
	) name13963 (
		_w12238_,
		_w12291_,
		_w14495_
	);
	LUT2 #(
		.INIT('h1)
	) name13964 (
		_w13269_,
		_w14495_,
		_w14496_
	);
	LUT2 #(
		.INIT('h4)
	) name13965 (
		_w13272_,
		_w14496_,
		_w14497_
	);
	LUT2 #(
		.INIT('h4)
	) name13966 (
		_w14494_,
		_w14497_,
		_w14498_
	);
	LUT2 #(
		.INIT('h1)
	) name13967 (
		\sa22_reg[1]/P0001 ,
		_w14498_,
		_w14499_
	);
	LUT2 #(
		.INIT('h4)
	) name13968 (
		\sa22_reg[2]/P0001 ,
		_w12268_,
		_w14500_
	);
	LUT2 #(
		.INIT('h1)
	) name13969 (
		_w12393_,
		_w12395_,
		_w14501_
	);
	LUT2 #(
		.INIT('h2)
	) name13970 (
		\sa22_reg[2]/P0001 ,
		_w14501_,
		_w14502_
	);
	LUT2 #(
		.INIT('h1)
	) name13971 (
		_w12281_,
		_w12324_,
		_w14503_
	);
	LUT2 #(
		.INIT('h4)
	) name13972 (
		_w14500_,
		_w14503_,
		_w14504_
	);
	LUT2 #(
		.INIT('h4)
	) name13973 (
		_w13803_,
		_w14504_,
		_w14505_
	);
	LUT2 #(
		.INIT('h4)
	) name13974 (
		_w14502_,
		_w14505_,
		_w14506_
	);
	LUT2 #(
		.INIT('h2)
	) name13975 (
		\sa22_reg[1]/P0001 ,
		_w14506_,
		_w14507_
	);
	LUT2 #(
		.INIT('h8)
	) name13976 (
		_w12238_,
		_w13197_,
		_w14508_
	);
	LUT2 #(
		.INIT('h1)
	) name13977 (
		\sa22_reg[2]/P0001 ,
		_w13193_,
		_w14509_
	);
	LUT2 #(
		.INIT('h8)
	) name13978 (
		_w12395_,
		_w12735_,
		_w14510_
	);
	LUT2 #(
		.INIT('h1)
	) name13979 (
		_w13258_,
		_w14508_,
		_w14511_
	);
	LUT2 #(
		.INIT('h4)
	) name13980 (
		_w14510_,
		_w14511_,
		_w14512_
	);
	LUT2 #(
		.INIT('h4)
	) name13981 (
		_w14509_,
		_w14512_,
		_w14513_
	);
	LUT2 #(
		.INIT('h4)
	) name13982 (
		_w14499_,
		_w14513_,
		_w14514_
	);
	LUT2 #(
		.INIT('h4)
	) name13983 (
		_w14507_,
		_w14514_,
		_w14515_
	);
	LUT2 #(
		.INIT('h1)
	) name13984 (
		\sa22_reg[0]/P0001 ,
		_w14515_,
		_w14516_
	);
	LUT2 #(
		.INIT('h1)
	) name13985 (
		_w12321_,
		_w12360_,
		_w14517_
	);
	LUT2 #(
		.INIT('h8)
	) name13986 (
		_w12794_,
		_w14517_,
		_w14518_
	);
	LUT2 #(
		.INIT('h1)
	) name13987 (
		\sa22_reg[2]/P0001 ,
		_w12259_,
		_w14519_
	);
	LUT2 #(
		.INIT('h4)
	) name13988 (
		_w12733_,
		_w14519_,
		_w14520_
	);
	LUT2 #(
		.INIT('h1)
	) name13989 (
		_w14518_,
		_w14520_,
		_w14521_
	);
	LUT2 #(
		.INIT('h1)
	) name13990 (
		_w12240_,
		_w12371_,
		_w14522_
	);
	LUT2 #(
		.INIT('h4)
	) name13991 (
		_w12812_,
		_w14522_,
		_w14523_
	);
	LUT2 #(
		.INIT('h4)
	) name13992 (
		_w14521_,
		_w14523_,
		_w14524_
	);
	LUT2 #(
		.INIT('h1)
	) name13993 (
		\sa22_reg[1]/P0001 ,
		_w14524_,
		_w14525_
	);
	LUT2 #(
		.INIT('h1)
	) name13994 (
		_w12330_,
		_w12344_,
		_w14526_
	);
	LUT2 #(
		.INIT('h4)
	) name13995 (
		_w12753_,
		_w14526_,
		_w14527_
	);
	LUT2 #(
		.INIT('h2)
	) name13996 (
		\sa22_reg[2]/P0001 ,
		_w14527_,
		_w14528_
	);
	LUT2 #(
		.INIT('h8)
	) name13997 (
		_w12234_,
		_w12779_,
		_w14529_
	);
	LUT2 #(
		.INIT('h1)
	) name13998 (
		_w12298_,
		_w12790_,
		_w14530_
	);
	LUT2 #(
		.INIT('h8)
	) name13999 (
		_w12251_,
		_w13200_,
		_w14531_
	);
	LUT2 #(
		.INIT('h1)
	) name14000 (
		_w13358_,
		_w14529_,
		_w14532_
	);
	LUT2 #(
		.INIT('h4)
	) name14001 (
		_w14531_,
		_w14532_,
		_w14533_
	);
	LUT2 #(
		.INIT('h8)
	) name14002 (
		_w14530_,
		_w14533_,
		_w14534_
	);
	LUT2 #(
		.INIT('h4)
	) name14003 (
		_w14528_,
		_w14534_,
		_w14535_
	);
	LUT2 #(
		.INIT('h2)
	) name14004 (
		\sa22_reg[1]/P0001 ,
		_w14535_,
		_w14536_
	);
	LUT2 #(
		.INIT('h2)
	) name14005 (
		_w13351_,
		_w14495_,
		_w14537_
	);
	LUT2 #(
		.INIT('h1)
	) name14006 (
		\sa22_reg[2]/P0001 ,
		_w14537_,
		_w14538_
	);
	LUT2 #(
		.INIT('h1)
	) name14007 (
		_w12264_,
		_w12374_,
		_w14539_
	);
	LUT2 #(
		.INIT('h8)
	) name14008 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w14540_
	);
	LUT2 #(
		.INIT('h4)
	) name14009 (
		_w14539_,
		_w14540_,
		_w14541_
	);
	LUT2 #(
		.INIT('h1)
	) name14010 (
		_w12343_,
		_w14541_,
		_w14542_
	);
	LUT2 #(
		.INIT('h4)
	) name14011 (
		_w14538_,
		_w14542_,
		_w14543_
	);
	LUT2 #(
		.INIT('h4)
	) name14012 (
		_w14525_,
		_w14543_,
		_w14544_
	);
	LUT2 #(
		.INIT('h4)
	) name14013 (
		_w14536_,
		_w14544_,
		_w14545_
	);
	LUT2 #(
		.INIT('h2)
	) name14014 (
		\sa22_reg[0]/P0001 ,
		_w14545_,
		_w14546_
	);
	LUT2 #(
		.INIT('h8)
	) name14015 (
		_w12756_,
		_w13227_,
		_w14547_
	);
	LUT2 #(
		.INIT('h8)
	) name14016 (
		\sa22_reg[6]/NET0131 ,
		_w12355_,
		_w14548_
	);
	LUT2 #(
		.INIT('h2)
	) name14017 (
		_w14530_,
		_w14548_,
		_w14549_
	);
	LUT2 #(
		.INIT('h2)
	) name14018 (
		\sa22_reg[2]/P0001 ,
		_w14549_,
		_w14550_
	);
	LUT2 #(
		.INIT('h1)
	) name14019 (
		_w12268_,
		_w12772_,
		_w14551_
	);
	LUT2 #(
		.INIT('h4)
	) name14020 (
		_w13240_,
		_w14551_,
		_w14552_
	);
	LUT2 #(
		.INIT('h2)
	) name14021 (
		_w13200_,
		_w14552_,
		_w14553_
	);
	LUT2 #(
		.INIT('h1)
	) name14022 (
		_w14547_,
		_w14550_,
		_w14554_
	);
	LUT2 #(
		.INIT('h4)
	) name14023 (
		_w14553_,
		_w14554_,
		_w14555_
	);
	LUT2 #(
		.INIT('h2)
	) name14024 (
		\sa22_reg[1]/P0001 ,
		_w14555_,
		_w14556_
	);
	LUT2 #(
		.INIT('h1)
	) name14025 (
		_w12335_,
		_w14508_,
		_w14557_
	);
	LUT2 #(
		.INIT('h2)
	) name14026 (
		_w13820_,
		_w14557_,
		_w14558_
	);
	LUT2 #(
		.INIT('h1)
	) name14027 (
		_w12292_,
		_w12773_,
		_w14559_
	);
	LUT2 #(
		.INIT('h2)
	) name14028 (
		_w12735_,
		_w14559_,
		_w14560_
	);
	LUT2 #(
		.INIT('h8)
	) name14029 (
		_w12383_,
		_w12782_,
		_w14561_
	);
	LUT2 #(
		.INIT('h1)
	) name14030 (
		_w13275_,
		_w14561_,
		_w14562_
	);
	LUT2 #(
		.INIT('h4)
	) name14031 (
		_w14560_,
		_w14562_,
		_w14563_
	);
	LUT2 #(
		.INIT('h4)
	) name14032 (
		_w14558_,
		_w14563_,
		_w14564_
	);
	LUT2 #(
		.INIT('h4)
	) name14033 (
		_w14556_,
		_w14564_,
		_w14565_
	);
	LUT2 #(
		.INIT('h4)
	) name14034 (
		_w14516_,
		_w14565_,
		_w14566_
	);
	LUT2 #(
		.INIT('h4)
	) name14035 (
		_w14546_,
		_w14566_,
		_w14567_
	);
	LUT2 #(
		.INIT('h2)
	) name14036 (
		_w14491_,
		_w14567_,
		_w14568_
	);
	LUT2 #(
		.INIT('h4)
	) name14037 (
		_w14491_,
		_w14567_,
		_w14569_
	);
	LUT2 #(
		.INIT('h1)
	) name14038 (
		_w14568_,
		_w14569_,
		_w14570_
	);
	LUT2 #(
		.INIT('h8)
	) name14039 (
		\sa33_reg[2]/P0001 ,
		_w12525_,
		_w14571_
	);
	LUT2 #(
		.INIT('h1)
	) name14040 (
		_w12564_,
		_w13720_,
		_w14572_
	);
	LUT2 #(
		.INIT('h1)
	) name14041 (
		\sa33_reg[2]/P0001 ,
		_w14572_,
		_w14573_
	);
	LUT2 #(
		.INIT('h1)
	) name14042 (
		_w12549_,
		_w12946_,
		_w14574_
	);
	LUT2 #(
		.INIT('h4)
	) name14043 (
		_w14011_,
		_w14574_,
		_w14575_
	);
	LUT2 #(
		.INIT('h1)
	) name14044 (
		_w12914_,
		_w13739_,
		_w14576_
	);
	LUT2 #(
		.INIT('h4)
	) name14045 (
		_w14571_,
		_w14576_,
		_w14577_
	);
	LUT2 #(
		.INIT('h8)
	) name14046 (
		_w14575_,
		_w14577_,
		_w14578_
	);
	LUT2 #(
		.INIT('h4)
	) name14047 (
		_w14573_,
		_w14578_,
		_w14579_
	);
	LUT2 #(
		.INIT('h1)
	) name14048 (
		\sa33_reg[1]/P0001 ,
		_w14579_,
		_w14580_
	);
	LUT2 #(
		.INIT('h8)
	) name14049 (
		_w12418_,
		_w13690_,
		_w14581_
	);
	LUT2 #(
		.INIT('h2)
	) name14050 (
		\sa33_reg[7]/NET0131 ,
		_w12446_,
		_w14582_
	);
	LUT2 #(
		.INIT('h4)
	) name14051 (
		_w12480_,
		_w14582_,
		_w14583_
	);
	LUT2 #(
		.INIT('h1)
	) name14052 (
		_w12430_,
		_w14583_,
		_w14584_
	);
	LUT2 #(
		.INIT('h2)
	) name14053 (
		\sa33_reg[2]/P0001 ,
		_w14584_,
		_w14585_
	);
	LUT2 #(
		.INIT('h1)
	) name14054 (
		_w12433_,
		_w12473_,
		_w14586_
	);
	LUT2 #(
		.INIT('h1)
	) name14055 (
		\sa33_reg[2]/P0001 ,
		_w14586_,
		_w14587_
	);
	LUT2 #(
		.INIT('h1)
	) name14056 (
		_w12861_,
		_w14581_,
		_w14588_
	);
	LUT2 #(
		.INIT('h4)
	) name14057 (
		_w14587_,
		_w14588_,
		_w14589_
	);
	LUT2 #(
		.INIT('h4)
	) name14058 (
		_w14585_,
		_w14589_,
		_w14590_
	);
	LUT2 #(
		.INIT('h2)
	) name14059 (
		\sa33_reg[1]/P0001 ,
		_w14590_,
		_w14591_
	);
	LUT2 #(
		.INIT('h8)
	) name14060 (
		_w12461_,
		_w12479_,
		_w14592_
	);
	LUT2 #(
		.INIT('h2)
	) name14061 (
		_w14074_,
		_w14592_,
		_w14593_
	);
	LUT2 #(
		.INIT('h1)
	) name14062 (
		\sa33_reg[2]/P0001 ,
		_w14593_,
		_w14594_
	);
	LUT2 #(
		.INIT('h8)
	) name14063 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w14595_
	);
	LUT2 #(
		.INIT('h4)
	) name14064 (
		_w12432_,
		_w12545_,
		_w14596_
	);
	LUT2 #(
		.INIT('h2)
	) name14065 (
		_w14595_,
		_w14596_,
		_w14597_
	);
	LUT2 #(
		.INIT('h1)
	) name14066 (
		_w12524_,
		_w14597_,
		_w14598_
	);
	LUT2 #(
		.INIT('h4)
	) name14067 (
		_w14594_,
		_w14598_,
		_w14599_
	);
	LUT2 #(
		.INIT('h4)
	) name14068 (
		_w14591_,
		_w14599_,
		_w14600_
	);
	LUT2 #(
		.INIT('h4)
	) name14069 (
		_w14580_,
		_w14600_,
		_w14601_
	);
	LUT2 #(
		.INIT('h2)
	) name14070 (
		\sa33_reg[0]/P0001 ,
		_w14601_,
		_w14602_
	);
	LUT2 #(
		.INIT('h4)
	) name14071 (
		\sa33_reg[7]/NET0131 ,
		_w12446_,
		_w14603_
	);
	LUT2 #(
		.INIT('h1)
	) name14072 (
		_w12570_,
		_w14603_,
		_w14604_
	);
	LUT2 #(
		.INIT('h2)
	) name14073 (
		\sa33_reg[2]/P0001 ,
		_w14604_,
		_w14605_
	);
	LUT2 #(
		.INIT('h2)
	) name14074 (
		_w12481_,
		_w12857_,
		_w14606_
	);
	LUT2 #(
		.INIT('h4)
	) name14075 (
		\sa33_reg[2]/P0001 ,
		_w12411_,
		_w14607_
	);
	LUT2 #(
		.INIT('h2)
	) name14076 (
		\sa33_reg[1]/P0001 ,
		_w12493_,
		_w14608_
	);
	LUT2 #(
		.INIT('h4)
	) name14077 (
		_w14606_,
		_w14608_,
		_w14609_
	);
	LUT2 #(
		.INIT('h4)
	) name14078 (
		_w14607_,
		_w14609_,
		_w14610_
	);
	LUT2 #(
		.INIT('h4)
	) name14079 (
		_w14605_,
		_w14610_,
		_w14611_
	);
	LUT2 #(
		.INIT('h8)
	) name14080 (
		_w12456_,
		_w12468_,
		_w14612_
	);
	LUT2 #(
		.INIT('h8)
	) name14081 (
		_w12472_,
		_w12868_,
		_w14613_
	);
	LUT2 #(
		.INIT('h1)
	) name14082 (
		_w12457_,
		_w14595_,
		_w14614_
	);
	LUT2 #(
		.INIT('h2)
	) name14083 (
		_w12465_,
		_w14614_,
		_w14615_
	);
	LUT2 #(
		.INIT('h1)
	) name14084 (
		\sa33_reg[1]/P0001 ,
		_w14592_,
		_w14616_
	);
	LUT2 #(
		.INIT('h4)
	) name14085 (
		_w14612_,
		_w14616_,
		_w14617_
	);
	LUT2 #(
		.INIT('h1)
	) name14086 (
		_w14613_,
		_w14615_,
		_w14618_
	);
	LUT2 #(
		.INIT('h8)
	) name14087 (
		_w14617_,
		_w14618_,
		_w14619_
	);
	LUT2 #(
		.INIT('h1)
	) name14088 (
		_w14611_,
		_w14619_,
		_w14620_
	);
	LUT2 #(
		.INIT('h1)
	) name14089 (
		_w12501_,
		_w12948_,
		_w14621_
	);
	LUT2 #(
		.INIT('h1)
	) name14090 (
		\sa33_reg[2]/P0001 ,
		_w14621_,
		_w14622_
	);
	LUT2 #(
		.INIT('h4)
	) name14091 (
		\sa33_reg[7]/NET0131 ,
		_w12476_,
		_w14623_
	);
	LUT2 #(
		.INIT('h8)
	) name14092 (
		_w13938_,
		_w14623_,
		_w14624_
	);
	LUT2 #(
		.INIT('h1)
	) name14093 (
		_w12518_,
		_w12856_,
		_w14625_
	);
	LUT2 #(
		.INIT('h4)
	) name14094 (
		_w14624_,
		_w14625_,
		_w14626_
	);
	LUT2 #(
		.INIT('h4)
	) name14095 (
		_w14622_,
		_w14626_,
		_w14627_
	);
	LUT2 #(
		.INIT('h4)
	) name14096 (
		_w14620_,
		_w14627_,
		_w14628_
	);
	LUT2 #(
		.INIT('h1)
	) name14097 (
		\sa33_reg[0]/P0001 ,
		_w14628_,
		_w14629_
	);
	LUT2 #(
		.INIT('h1)
	) name14098 (
		_w12526_,
		_w14005_,
		_w14630_
	);
	LUT2 #(
		.INIT('h2)
	) name14099 (
		_w12945_,
		_w14630_,
		_w14631_
	);
	LUT2 #(
		.INIT('h8)
	) name14100 (
		_w12456_,
		_w14044_,
		_w14632_
	);
	LUT2 #(
		.INIT('h8)
	) name14101 (
		\sa33_reg[6]/P0001 ,
		_w12444_,
		_w14633_
	);
	LUT2 #(
		.INIT('h1)
	) name14102 (
		_w12411_,
		_w13970_,
		_w14634_
	);
	LUT2 #(
		.INIT('h4)
	) name14103 (
		_w14633_,
		_w14634_,
		_w14635_
	);
	LUT2 #(
		.INIT('h2)
	) name14104 (
		_w13952_,
		_w14635_,
		_w14636_
	);
	LUT2 #(
		.INIT('h1)
	) name14105 (
		_w12883_,
		_w14632_,
		_w14637_
	);
	LUT2 #(
		.INIT('h4)
	) name14106 (
		_w14631_,
		_w14637_,
		_w14638_
	);
	LUT2 #(
		.INIT('h4)
	) name14107 (
		_w14636_,
		_w14638_,
		_w14639_
	);
	LUT2 #(
		.INIT('h2)
	) name14108 (
		\sa33_reg[1]/P0001 ,
		_w14639_,
		_w14640_
	);
	LUT2 #(
		.INIT('h1)
	) name14109 (
		_w12508_,
		_w12518_,
		_w14641_
	);
	LUT2 #(
		.INIT('h2)
	) name14110 (
		_w13741_,
		_w14641_,
		_w14642_
	);
	LUT2 #(
		.INIT('h1)
	) name14111 (
		_w12458_,
		_w13948_,
		_w14643_
	);
	LUT2 #(
		.INIT('h2)
	) name14112 (
		_w12877_,
		_w14643_,
		_w14644_
	);
	LUT2 #(
		.INIT('h8)
	) name14113 (
		_w12462_,
		_w12560_,
		_w14645_
	);
	LUT2 #(
		.INIT('h1)
	) name14114 (
		_w13740_,
		_w14645_,
		_w14646_
	);
	LUT2 #(
		.INIT('h4)
	) name14115 (
		_w14644_,
		_w14646_,
		_w14647_
	);
	LUT2 #(
		.INIT('h4)
	) name14116 (
		_w14642_,
		_w14647_,
		_w14648_
	);
	LUT2 #(
		.INIT('h4)
	) name14117 (
		_w14640_,
		_w14648_,
		_w14649_
	);
	LUT2 #(
		.INIT('h4)
	) name14118 (
		_w14629_,
		_w14649_,
		_w14650_
	);
	LUT2 #(
		.INIT('h4)
	) name14119 (
		_w14602_,
		_w14650_,
		_w14651_
	);
	LUT2 #(
		.INIT('h2)
	) name14120 (
		\u0_w_reg[0][27]/P0001 ,
		_w14651_,
		_w14652_
	);
	LUT2 #(
		.INIT('h4)
	) name14121 (
		\u0_w_reg[0][27]/P0001 ,
		_w14651_,
		_w14653_
	);
	LUT2 #(
		.INIT('h1)
	) name14122 (
		_w14652_,
		_w14653_,
		_w14654_
	);
	LUT2 #(
		.INIT('h8)
	) name14123 (
		_w14570_,
		_w14654_,
		_w14655_
	);
	LUT2 #(
		.INIT('h1)
	) name14124 (
		_w14570_,
		_w14654_,
		_w14656_
	);
	LUT2 #(
		.INIT('h1)
	) name14125 (
		_w14655_,
		_w14656_,
		_w14657_
	);
	LUT2 #(
		.INIT('h2)
	) name14126 (
		_w13558_,
		_w14400_,
		_w14658_
	);
	LUT2 #(
		.INIT('h4)
	) name14127 (
		_w13558_,
		_w14400_,
		_w14659_
	);
	LUT2 #(
		.INIT('h1)
	) name14128 (
		_w14658_,
		_w14659_,
		_w14660_
	);
	LUT2 #(
		.INIT('h8)
	) name14129 (
		\sa11_reg[4]/P0001 ,
		_w13139_,
		_w14661_
	);
	LUT2 #(
		.INIT('h2)
	) name14130 (
		_w14156_,
		_w14661_,
		_w14662_
	);
	LUT2 #(
		.INIT('h1)
	) name14131 (
		\sa11_reg[2]/P0001 ,
		_w14662_,
		_w14663_
	);
	LUT2 #(
		.INIT('h1)
	) name14132 (
		_w11935_,
		_w14663_,
		_w14664_
	);
	LUT2 #(
		.INIT('h2)
	) name14133 (
		\sa11_reg[1]/P0001 ,
		_w14664_,
		_w14665_
	);
	LUT2 #(
		.INIT('h1)
	) name14134 (
		_w11826_,
		_w11922_,
		_w14666_
	);
	LUT2 #(
		.INIT('h4)
	) name14135 (
		_w13155_,
		_w14666_,
		_w14667_
	);
	LUT2 #(
		.INIT('h8)
	) name14136 (
		_w13524_,
		_w14667_,
		_w14668_
	);
	LUT2 #(
		.INIT('h8)
	) name14137 (
		\sa11_reg[3]/P0001 ,
		_w11876_,
		_w14669_
	);
	LUT2 #(
		.INIT('h1)
	) name14138 (
		_w11934_,
		_w14669_,
		_w14670_
	);
	LUT2 #(
		.INIT('h8)
	) name14139 (
		_w13549_,
		_w14670_,
		_w14671_
	);
	LUT2 #(
		.INIT('h1)
	) name14140 (
		_w14668_,
		_w14671_,
		_w14672_
	);
	LUT2 #(
		.INIT('h2)
	) name14141 (
		_w11876_,
		_w11877_,
		_w14673_
	);
	LUT2 #(
		.INIT('h4)
	) name14142 (
		_w13092_,
		_w14673_,
		_w14674_
	);
	LUT2 #(
		.INIT('h1)
	) name14143 (
		_w14672_,
		_w14674_,
		_w14675_
	);
	LUT2 #(
		.INIT('h1)
	) name14144 (
		\sa11_reg[1]/P0001 ,
		_w14675_,
		_w14676_
	);
	LUT2 #(
		.INIT('h8)
	) name14145 (
		_w11796_,
		_w12194_,
		_w14677_
	);
	LUT2 #(
		.INIT('h1)
	) name14146 (
		_w11861_,
		_w12223_,
		_w14678_
	);
	LUT2 #(
		.INIT('h4)
	) name14147 (
		_w14677_,
		_w14678_,
		_w14679_
	);
	LUT2 #(
		.INIT('h2)
	) name14148 (
		_w13171_,
		_w14679_,
		_w14680_
	);
	LUT2 #(
		.INIT('h1)
	) name14149 (
		_w11801_,
		_w11847_,
		_w14681_
	);
	LUT2 #(
		.INIT('h2)
	) name14150 (
		_w13457_,
		_w14681_,
		_w14682_
	);
	LUT2 #(
		.INIT('h1)
	) name14151 (
		_w11933_,
		_w13159_,
		_w14683_
	);
	LUT2 #(
		.INIT('h4)
	) name14152 (
		_w14164_,
		_w14683_,
		_w14684_
	);
	LUT2 #(
		.INIT('h2)
	) name14153 (
		_w11846_,
		_w14684_,
		_w14685_
	);
	LUT2 #(
		.INIT('h1)
	) name14154 (
		\sa11_reg[5]/P0001 ,
		_w11893_,
		_w14686_
	);
	LUT2 #(
		.INIT('h2)
	) name14155 (
		_w12146_,
		_w14686_,
		_w14687_
	);
	LUT2 #(
		.INIT('h1)
	) name14156 (
		_w11849_,
		_w11887_,
		_w14688_
	);
	LUT2 #(
		.INIT('h4)
	) name14157 (
		_w11942_,
		_w14688_,
		_w14689_
	);
	LUT2 #(
		.INIT('h1)
	) name14158 (
		_w11793_,
		_w11824_,
		_w14690_
	);
	LUT2 #(
		.INIT('h2)
	) name14159 (
		_w11897_,
		_w14687_,
		_w14691_
	);
	LUT2 #(
		.INIT('h8)
	) name14160 (
		_w14690_,
		_w14691_,
		_w14692_
	);
	LUT2 #(
		.INIT('h8)
	) name14161 (
		_w14689_,
		_w14692_,
		_w14693_
	);
	LUT2 #(
		.INIT('h8)
	) name14162 (
		_w11831_,
		_w13092_,
		_w14694_
	);
	LUT2 #(
		.INIT('h1)
	) name14163 (
		_w13131_,
		_w13489_,
		_w14695_
	);
	LUT2 #(
		.INIT('h1)
	) name14164 (
		\sa11_reg[2]/P0001 ,
		_w14695_,
		_w14696_
	);
	LUT2 #(
		.INIT('h2)
	) name14165 (
		\sa11_reg[1]/P0001 ,
		_w14694_,
		_w14697_
	);
	LUT2 #(
		.INIT('h4)
	) name14166 (
		_w13440_,
		_w14697_,
		_w14698_
	);
	LUT2 #(
		.INIT('h4)
	) name14167 (
		_w14696_,
		_w14698_,
		_w14699_
	);
	LUT2 #(
		.INIT('h1)
	) name14168 (
		_w14693_,
		_w14699_,
		_w14700_
	);
	LUT2 #(
		.INIT('h1)
	) name14169 (
		_w11849_,
		_w11865_,
		_w14701_
	);
	LUT2 #(
		.INIT('h2)
	) name14170 (
		\sa11_reg[5]/P0001 ,
		_w14701_,
		_w14702_
	);
	LUT2 #(
		.INIT('h2)
	) name14171 (
		\sa11_reg[0]/P0001 ,
		_w11921_,
		_w14703_
	);
	LUT2 #(
		.INIT('h4)
	) name14172 (
		_w14702_,
		_w14703_,
		_w14704_
	);
	LUT2 #(
		.INIT('h4)
	) name14173 (
		_w14685_,
		_w14704_,
		_w14705_
	);
	LUT2 #(
		.INIT('h4)
	) name14174 (
		_w14700_,
		_w14705_,
		_w14706_
	);
	LUT2 #(
		.INIT('h8)
	) name14175 (
		_w11846_,
		_w12223_,
		_w14707_
	);
	LUT2 #(
		.INIT('h1)
	) name14176 (
		_w11915_,
		_w12146_,
		_w14708_
	);
	LUT2 #(
		.INIT('h2)
	) name14177 (
		\sa11_reg[2]/P0001 ,
		_w14708_,
		_w14709_
	);
	LUT2 #(
		.INIT('h1)
	) name14178 (
		_w13513_,
		_w14709_,
		_w14710_
	);
	LUT2 #(
		.INIT('h2)
	) name14179 (
		\sa11_reg[1]/P0001 ,
		_w14710_,
		_w14711_
	);
	LUT2 #(
		.INIT('h1)
	) name14180 (
		_w11858_,
		_w13092_,
		_w14712_
	);
	LUT2 #(
		.INIT('h2)
	) name14181 (
		\sa11_reg[1]/P0001 ,
		_w11825_,
		_w14713_
	);
	LUT2 #(
		.INIT('h4)
	) name14182 (
		_w14712_,
		_w14713_,
		_w14714_
	);
	LUT2 #(
		.INIT('h1)
	) name14183 (
		_w11881_,
		_w14714_,
		_w14715_
	);
	LUT2 #(
		.INIT('h1)
	) name14184 (
		\sa11_reg[2]/P0001 ,
		_w14715_,
		_w14716_
	);
	LUT2 #(
		.INIT('h1)
	) name14185 (
		_w13439_,
		_w13447_,
		_w14717_
	);
	LUT2 #(
		.INIT('h1)
	) name14186 (
		\sa11_reg[1]/P0001 ,
		_w14717_,
		_w14718_
	);
	LUT2 #(
		.INIT('h1)
	) name14187 (
		\sa11_reg[0]/P0001 ,
		_w11898_,
		_w14719_
	);
	LUT2 #(
		.INIT('h4)
	) name14188 (
		_w14707_,
		_w14719_,
		_w14720_
	);
	LUT2 #(
		.INIT('h4)
	) name14189 (
		_w14716_,
		_w14720_,
		_w14721_
	);
	LUT2 #(
		.INIT('h4)
	) name14190 (
		_w14718_,
		_w14721_,
		_w14722_
	);
	LUT2 #(
		.INIT('h4)
	) name14191 (
		_w14711_,
		_w14722_,
		_w14723_
	);
	LUT2 #(
		.INIT('h1)
	) name14192 (
		_w14706_,
		_w14723_,
		_w14724_
	);
	LUT2 #(
		.INIT('h1)
	) name14193 (
		_w14446_,
		_w14682_,
		_w14725_
	);
	LUT2 #(
		.INIT('h4)
	) name14194 (
		_w14680_,
		_w14725_,
		_w14726_
	);
	LUT2 #(
		.INIT('h4)
	) name14195 (
		_w14665_,
		_w14726_,
		_w14727_
	);
	LUT2 #(
		.INIT('h4)
	) name14196 (
		_w14676_,
		_w14727_,
		_w14728_
	);
	LUT2 #(
		.INIT('h4)
	) name14197 (
		_w14724_,
		_w14728_,
		_w14729_
	);
	LUT2 #(
		.INIT('h1)
	) name14198 (
		_w12008_,
		_w12015_,
		_w14730_
	);
	LUT2 #(
		.INIT('h2)
	) name14199 (
		\sa00_reg[2]/P0001 ,
		_w14730_,
		_w14731_
	);
	LUT2 #(
		.INIT('h1)
	) name14200 (
		_w11979_,
		_w12007_,
		_w14732_
	);
	LUT2 #(
		.INIT('h1)
	) name14201 (
		\sa00_reg[2]/P0001 ,
		_w12026_,
		_w14733_
	);
	LUT2 #(
		.INIT('h4)
	) name14202 (
		_w14732_,
		_w14733_,
		_w14734_
	);
	LUT2 #(
		.INIT('h1)
	) name14203 (
		_w13069_,
		_w14734_,
		_w14735_
	);
	LUT2 #(
		.INIT('h4)
	) name14204 (
		_w14731_,
		_w14735_,
		_w14736_
	);
	LUT2 #(
		.INIT('h2)
	) name14205 (
		\sa00_reg[1]/P0001 ,
		_w14736_,
		_w14737_
	);
	LUT2 #(
		.INIT('h8)
	) name14206 (
		_w13004_,
		_w14279_,
		_w14738_
	);
	LUT2 #(
		.INIT('h8)
	) name14207 (
		_w12026_,
		_w13044_,
		_w14739_
	);
	LUT2 #(
		.INIT('h1)
	) name14208 (
		_w14390_,
		_w14739_,
		_w14740_
	);
	LUT2 #(
		.INIT('h1)
	) name14209 (
		\sa00_reg[1]/P0001 ,
		_w14740_,
		_w14741_
	);
	LUT2 #(
		.INIT('h1)
	) name14210 (
		_w11976_,
		_w14738_,
		_w14742_
	);
	LUT2 #(
		.INIT('h4)
	) name14211 (
		_w13060_,
		_w14742_,
		_w14743_
	);
	LUT2 #(
		.INIT('h4)
	) name14212 (
		_w14741_,
		_w14743_,
		_w14744_
	);
	LUT2 #(
		.INIT('h4)
	) name14213 (
		_w14737_,
		_w14744_,
		_w14745_
	);
	LUT2 #(
		.INIT('h1)
	) name14214 (
		\sa00_reg[0]/P0001 ,
		_w14745_,
		_w14746_
	);
	LUT2 #(
		.INIT('h8)
	) name14215 (
		\sa00_reg[1]/P0001 ,
		_w12054_,
		_w14747_
	);
	LUT2 #(
		.INIT('h8)
	) name14216 (
		_w12066_,
		_w14747_,
		_w14748_
	);
	LUT2 #(
		.INIT('h1)
	) name14217 (
		_w11967_,
		_w12096_,
		_w14749_
	);
	LUT2 #(
		.INIT('h2)
	) name14218 (
		_w14305_,
		_w14749_,
		_w14750_
	);
	LUT2 #(
		.INIT('h8)
	) name14219 (
		_w12091_,
		_w13044_,
		_w14751_
	);
	LUT2 #(
		.INIT('h1)
	) name14220 (
		_w12005_,
		_w13559_,
		_w14752_
	);
	LUT2 #(
		.INIT('h8)
	) name14221 (
		\sa00_reg[7]/NET0131 ,
		_w13571_,
		_w14753_
	);
	LUT2 #(
		.INIT('h4)
	) name14222 (
		_w14752_,
		_w14753_,
		_w14754_
	);
	LUT2 #(
		.INIT('h1)
	) name14223 (
		_w12024_,
		_w12034_,
		_w14755_
	);
	LUT2 #(
		.INIT('h8)
	) name14224 (
		_w14391_,
		_w14755_,
		_w14756_
	);
	LUT2 #(
		.INIT('h1)
	) name14225 (
		\sa00_reg[2]/P0001 ,
		_w14371_,
		_w14757_
	);
	LUT2 #(
		.INIT('h4)
	) name14226 (
		_w12018_,
		_w14757_,
		_w14758_
	);
	LUT2 #(
		.INIT('h4)
	) name14227 (
		_w13077_,
		_w14758_,
		_w14759_
	);
	LUT2 #(
		.INIT('h1)
	) name14228 (
		_w14756_,
		_w14759_,
		_w14760_
	);
	LUT2 #(
		.INIT('h4)
	) name14229 (
		_w11955_,
		_w11960_,
		_w14761_
	);
	LUT2 #(
		.INIT('h4)
	) name14230 (
		_w12007_,
		_w14761_,
		_w14762_
	);
	LUT2 #(
		.INIT('h1)
	) name14231 (
		\sa00_reg[1]/P0001 ,
		_w13018_,
		_w14763_
	);
	LUT2 #(
		.INIT('h4)
	) name14232 (
		_w14762_,
		_w14763_,
		_w14764_
	);
	LUT2 #(
		.INIT('h4)
	) name14233 (
		_w14760_,
		_w14764_,
		_w14765_
	);
	LUT2 #(
		.INIT('h4)
	) name14234 (
		_w12600_,
		_w13594_,
		_w14766_
	);
	LUT2 #(
		.INIT('h1)
	) name14235 (
		\sa00_reg[2]/P0001 ,
		_w14766_,
		_w14767_
	);
	LUT2 #(
		.INIT('h2)
	) name14236 (
		\sa00_reg[1]/P0001 ,
		_w12033_,
		_w14768_
	);
	LUT2 #(
		.INIT('h4)
	) name14237 (
		_w14767_,
		_w14768_,
		_w14769_
	);
	LUT2 #(
		.INIT('h1)
	) name14238 (
		_w14765_,
		_w14769_,
		_w14770_
	);
	LUT2 #(
		.INIT('h1)
	) name14239 (
		_w12691_,
		_w12692_,
		_w14771_
	);
	LUT2 #(
		.INIT('h1)
	) name14240 (
		\sa00_reg[2]/P0001 ,
		_w14771_,
		_w14772_
	);
	LUT2 #(
		.INIT('h8)
	) name14241 (
		_w11962_,
		_w12056_,
		_w14773_
	);
	LUT2 #(
		.INIT('h1)
	) name14242 (
		_w11954_,
		_w12095_,
		_w14774_
	);
	LUT2 #(
		.INIT('h1)
	) name14243 (
		_w14248_,
		_w14773_,
		_w14775_
	);
	LUT2 #(
		.INIT('h8)
	) name14244 (
		_w14774_,
		_w14775_,
		_w14776_
	);
	LUT2 #(
		.INIT('h2)
	) name14245 (
		_w11981_,
		_w12023_,
		_w14777_
	);
	LUT2 #(
		.INIT('h8)
	) name14246 (
		_w14776_,
		_w14777_,
		_w14778_
	);
	LUT2 #(
		.INIT('h4)
	) name14247 (
		_w14772_,
		_w14778_,
		_w14779_
	);
	LUT2 #(
		.INIT('h8)
	) name14248 (
		\sa00_reg[2]/P0001 ,
		_w12636_,
		_w14780_
	);
	LUT2 #(
		.INIT('h1)
	) name14249 (
		_w13028_,
		_w13036_,
		_w14781_
	);
	LUT2 #(
		.INIT('h1)
	) name14250 (
		\sa00_reg[2]/P0001 ,
		_w14781_,
		_w14782_
	);
	LUT2 #(
		.INIT('h2)
	) name14251 (
		\sa00_reg[1]/P0001 ,
		_w14308_,
		_w14783_
	);
	LUT2 #(
		.INIT('h4)
	) name14252 (
		_w14780_,
		_w14783_,
		_w14784_
	);
	LUT2 #(
		.INIT('h4)
	) name14253 (
		_w14782_,
		_w14784_,
		_w14785_
	);
	LUT2 #(
		.INIT('h1)
	) name14254 (
		_w14779_,
		_w14785_,
		_w14786_
	);
	LUT2 #(
		.INIT('h8)
	) name14255 (
		_w12056_,
		_w12651_,
		_w14787_
	);
	LUT2 #(
		.INIT('h1)
	) name14256 (
		_w11996_,
		_w13068_,
		_w14788_
	);
	LUT2 #(
		.INIT('h4)
	) name14257 (
		_w13610_,
		_w14788_,
		_w14789_
	);
	LUT2 #(
		.INIT('h2)
	) name14258 (
		_w12054_,
		_w14789_,
		_w14790_
	);
	LUT2 #(
		.INIT('h1)
	) name14259 (
		_w12016_,
		_w12022_,
		_w14791_
	);
	LUT2 #(
		.INIT('h4)
	) name14260 (
		_w14787_,
		_w14791_,
		_w14792_
	);
	LUT2 #(
		.INIT('h4)
	) name14261 (
		_w14790_,
		_w14792_,
		_w14793_
	);
	LUT2 #(
		.INIT('h4)
	) name14262 (
		_w14786_,
		_w14793_,
		_w14794_
	);
	LUT2 #(
		.INIT('h2)
	) name14263 (
		\sa00_reg[0]/P0001 ,
		_w14794_,
		_w14795_
	);
	LUT2 #(
		.INIT('h1)
	) name14264 (
		_w14748_,
		_w14750_,
		_w14796_
	);
	LUT2 #(
		.INIT('h1)
	) name14265 (
		_w14751_,
		_w14754_,
		_w14797_
	);
	LUT2 #(
		.INIT('h8)
	) name14266 (
		_w14796_,
		_w14797_,
		_w14798_
	);
	LUT2 #(
		.INIT('h4)
	) name14267 (
		_w14746_,
		_w14798_,
		_w14799_
	);
	LUT2 #(
		.INIT('h4)
	) name14268 (
		_w14770_,
		_w14799_,
		_w14800_
	);
	LUT2 #(
		.INIT('h4)
	) name14269 (
		_w14795_,
		_w14800_,
		_w14801_
	);
	LUT2 #(
		.INIT('h2)
	) name14270 (
		_w14729_,
		_w14801_,
		_w14802_
	);
	LUT2 #(
		.INIT('h4)
	) name14271 (
		_w14729_,
		_w14801_,
		_w14803_
	);
	LUT2 #(
		.INIT('h1)
	) name14272 (
		_w14802_,
		_w14803_,
		_w14804_
	);
	LUT2 #(
		.INIT('h4)
	) name14273 (
		_w14660_,
		_w14804_,
		_w14805_
	);
	LUT2 #(
		.INIT('h2)
	) name14274 (
		_w14660_,
		_w14804_,
		_w14806_
	);
	LUT2 #(
		.INIT('h1)
	) name14275 (
		_w14805_,
		_w14806_,
		_w14807_
	);
	LUT2 #(
		.INIT('h2)
	) name14276 (
		_w14657_,
		_w14807_,
		_w14808_
	);
	LUT2 #(
		.INIT('h4)
	) name14277 (
		_w14657_,
		_w14807_,
		_w14809_
	);
	LUT2 #(
		.INIT('h1)
	) name14278 (
		\ld_r_reg/P0001 ,
		_w14808_,
		_w14810_
	);
	LUT2 #(
		.INIT('h4)
	) name14279 (
		_w14809_,
		_w14810_,
		_w14811_
	);
	LUT2 #(
		.INIT('h2)
	) name14280 (
		\text_in_r_reg[123]/P0001 ,
		\u0_w_reg[0][27]/P0001 ,
		_w14812_
	);
	LUT2 #(
		.INIT('h4)
	) name14281 (
		\text_in_r_reg[123]/P0001 ,
		\u0_w_reg[0][27]/P0001 ,
		_w14813_
	);
	LUT2 #(
		.INIT('h2)
	) name14282 (
		\ld_r_reg/P0001 ,
		_w14812_,
		_w14814_
	);
	LUT2 #(
		.INIT('h4)
	) name14283 (
		_w14813_,
		_w14814_,
		_w14815_
	);
	LUT2 #(
		.INIT('h1)
	) name14284 (
		_w14811_,
		_w14815_,
		_w14816_
	);
	LUT2 #(
		.INIT('h2)
	) name14285 (
		_w13922_,
		_w14567_,
		_w14817_
	);
	LUT2 #(
		.INIT('h4)
	) name14286 (
		_w13922_,
		_w14567_,
		_w14818_
	);
	LUT2 #(
		.INIT('h1)
	) name14287 (
		_w14817_,
		_w14818_,
		_w14819_
	);
	LUT2 #(
		.INIT('h2)
	) name14288 (
		\u0_w_reg[0][19]/P0001 ,
		_w14651_,
		_w14820_
	);
	LUT2 #(
		.INIT('h4)
	) name14289 (
		\u0_w_reg[0][19]/P0001 ,
		_w14651_,
		_w14821_
	);
	LUT2 #(
		.INIT('h1)
	) name14290 (
		_w14820_,
		_w14821_,
		_w14822_
	);
	LUT2 #(
		.INIT('h8)
	) name14291 (
		_w14819_,
		_w14822_,
		_w14823_
	);
	LUT2 #(
		.INIT('h1)
	) name14292 (
		_w14819_,
		_w14822_,
		_w14824_
	);
	LUT2 #(
		.INIT('h1)
	) name14293 (
		_w14823_,
		_w14824_,
		_w14825_
	);
	LUT2 #(
		.INIT('h8)
	) name14294 (
		_w12244_,
		_w12266_,
		_w14826_
	);
	LUT2 #(
		.INIT('h2)
	) name14295 (
		_w13804_,
		_w14826_,
		_w14827_
	);
	LUT2 #(
		.INIT('h1)
	) name14296 (
		\sa22_reg[2]/P0001 ,
		_w14827_,
		_w14828_
	);
	LUT2 #(
		.INIT('h1)
	) name14297 (
		_w12259_,
		_w14828_,
		_w14829_
	);
	LUT2 #(
		.INIT('h2)
	) name14298 (
		\sa22_reg[1]/P0001 ,
		_w14829_,
		_w14830_
	);
	LUT2 #(
		.INIT('h1)
	) name14299 (
		_w12235_,
		_w13358_,
		_w14831_
	);
	LUT2 #(
		.INIT('h4)
	) name14300 (
		_w12806_,
		_w14831_,
		_w14832_
	);
	LUT2 #(
		.INIT('h2)
	) name14301 (
		\sa22_reg[2]/P0001 ,
		_w14832_,
		_w14833_
	);
	LUT2 #(
		.INIT('h1)
	) name14302 (
		_w12738_,
		_w13257_,
		_w14834_
	);
	LUT2 #(
		.INIT('h4)
	) name14303 (
		_w12384_,
		_w14834_,
		_w14835_
	);
	LUT2 #(
		.INIT('h1)
	) name14304 (
		\sa22_reg[2]/P0001 ,
		_w14835_,
		_w14836_
	);
	LUT2 #(
		.INIT('h1)
	) name14305 (
		_w12756_,
		_w13911_,
		_w14837_
	);
	LUT2 #(
		.INIT('h4)
	) name14306 (
		_w13201_,
		_w14837_,
		_w14838_
	);
	LUT2 #(
		.INIT('h4)
	) name14307 (
		_w14833_,
		_w14838_,
		_w14839_
	);
	LUT2 #(
		.INIT('h4)
	) name14308 (
		_w14836_,
		_w14839_,
		_w14840_
	);
	LUT2 #(
		.INIT('h1)
	) name14309 (
		\sa22_reg[1]/P0001 ,
		_w14840_,
		_w14841_
	);
	LUT2 #(
		.INIT('h8)
	) name14310 (
		_w12303_,
		_w13197_,
		_w14842_
	);
	LUT2 #(
		.INIT('h1)
	) name14311 (
		_w12345_,
		_w12385_,
		_w14843_
	);
	LUT2 #(
		.INIT('h4)
	) name14312 (
		_w14842_,
		_w14843_,
		_w14844_
	);
	LUT2 #(
		.INIT('h2)
	) name14313 (
		_w13264_,
		_w14844_,
		_w14845_
	);
	LUT2 #(
		.INIT('h1)
	) name14314 (
		_w12291_,
		_w12332_,
		_w14846_
	);
	LUT2 #(
		.INIT('h8)
	) name14315 (
		\sa22_reg[2]/P0001 ,
		_w12238_,
		_w14847_
	);
	LUT2 #(
		.INIT('h4)
	) name14316 (
		_w14846_,
		_w14847_,
		_w14848_
	);
	LUT2 #(
		.INIT('h1)
	) name14317 (
		_w12395_,
		_w12805_,
		_w14849_
	);
	LUT2 #(
		.INIT('h8)
	) name14318 (
		_w13319_,
		_w14849_,
		_w14850_
	);
	LUT2 #(
		.INIT('h2)
	) name14319 (
		\sa22_reg[2]/P0001 ,
		_w13265_,
		_w14851_
	);
	LUT2 #(
		.INIT('h4)
	) name14320 (
		_w12353_,
		_w14851_,
		_w14852_
	);
	LUT2 #(
		.INIT('h1)
	) name14321 (
		_w14850_,
		_w14852_,
		_w14853_
	);
	LUT2 #(
		.INIT('h1)
	) name14322 (
		_w13252_,
		_w14853_,
		_w14854_
	);
	LUT2 #(
		.INIT('h2)
	) name14323 (
		\sa22_reg[1]/P0001 ,
		_w14854_,
		_w14855_
	);
	LUT2 #(
		.INIT('h8)
	) name14324 (
		\sa22_reg[2]/P0001 ,
		_w12722_,
		_w14856_
	);
	LUT2 #(
		.INIT('h8)
	) name14325 (
		_w12349_,
		_w13227_,
		_w14857_
	);
	LUT2 #(
		.INIT('h1)
	) name14326 (
		_w13358_,
		_w14857_,
		_w14858_
	);
	LUT2 #(
		.INIT('h1)
	) name14327 (
		\sa22_reg[1]/P0001 ,
		_w14858_,
		_w14859_
	);
	LUT2 #(
		.INIT('h1)
	) name14328 (
		_w12298_,
		_w13273_,
		_w14860_
	);
	LUT2 #(
		.INIT('h4)
	) name14329 (
		_w14856_,
		_w14860_,
		_w14861_
	);
	LUT2 #(
		.INIT('h4)
	) name14330 (
		_w14859_,
		_w14861_,
		_w14862_
	);
	LUT2 #(
		.INIT('h4)
	) name14331 (
		_w14855_,
		_w14862_,
		_w14863_
	);
	LUT2 #(
		.INIT('h1)
	) name14332 (
		\sa22_reg[0]/P0001 ,
		_w14863_,
		_w14864_
	);
	LUT2 #(
		.INIT('h8)
	) name14333 (
		_w12251_,
		_w12322_,
		_w14865_
	);
	LUT2 #(
		.INIT('h8)
	) name14334 (
		_w12301_,
		_w13200_,
		_w14866_
	);
	LUT2 #(
		.INIT('h1)
	) name14335 (
		_w12771_,
		_w12782_,
		_w14867_
	);
	LUT2 #(
		.INIT('h1)
	) name14336 (
		_w13303_,
		_w14865_,
		_w14868_
	);
	LUT2 #(
		.INIT('h8)
	) name14337 (
		_w14867_,
		_w14868_,
		_w14869_
	);
	LUT2 #(
		.INIT('h1)
	) name14338 (
		_w12760_,
		_w12813_,
		_w14870_
	);
	LUT2 #(
		.INIT('h4)
	) name14339 (
		_w14866_,
		_w14870_,
		_w14871_
	);
	LUT2 #(
		.INIT('h4)
	) name14340 (
		_w12346_,
		_w14869_,
		_w14872_
	);
	LUT2 #(
		.INIT('h8)
	) name14341 (
		_w14871_,
		_w14872_,
		_w14873_
	);
	LUT2 #(
		.INIT('h1)
	) name14342 (
		\sa22_reg[1]/P0001 ,
		_w14873_,
		_w14874_
	);
	LUT2 #(
		.INIT('h1)
	) name14343 (
		_w12302_,
		_w13240_,
		_w14875_
	);
	LUT2 #(
		.INIT('h8)
	) name14344 (
		_w13367_,
		_w14875_,
		_w14876_
	);
	LUT2 #(
		.INIT('h2)
	) name14345 (
		\sa22_reg[2]/P0001 ,
		_w12301_,
		_w14877_
	);
	LUT2 #(
		.INIT('h2)
	) name14346 (
		\sa22_reg[1]/P0001 ,
		_w14877_,
		_w14878_
	);
	LUT2 #(
		.INIT('h4)
	) name14347 (
		_w14876_,
		_w14878_,
		_w14879_
	);
	LUT2 #(
		.INIT('h1)
	) name14348 (
		_w12319_,
		_w13251_,
		_w14880_
	);
	LUT2 #(
		.INIT('h4)
	) name14349 (
		_w13782_,
		_w14880_,
		_w14881_
	);
	LUT2 #(
		.INIT('h2)
	) name14350 (
		_w12735_,
		_w14881_,
		_w14882_
	);
	LUT2 #(
		.INIT('h1)
	) name14351 (
		_w12802_,
		_w12809_,
		_w14883_
	);
	LUT2 #(
		.INIT('h4)
	) name14352 (
		_w13754_,
		_w14883_,
		_w14884_
	);
	LUT2 #(
		.INIT('h4)
	) name14353 (
		_w14879_,
		_w14884_,
		_w14885_
	);
	LUT2 #(
		.INIT('h4)
	) name14354 (
		_w14882_,
		_w14885_,
		_w14886_
	);
	LUT2 #(
		.INIT('h4)
	) name14355 (
		_w14874_,
		_w14886_,
		_w14887_
	);
	LUT2 #(
		.INIT('h2)
	) name14356 (
		\sa22_reg[0]/P0001 ,
		_w14887_,
		_w14888_
	);
	LUT2 #(
		.INIT('h1)
	) name14357 (
		_w14547_,
		_w14848_,
		_w14889_
	);
	LUT2 #(
		.INIT('h4)
	) name14358 (
		_w14845_,
		_w14889_,
		_w14890_
	);
	LUT2 #(
		.INIT('h4)
	) name14359 (
		_w14841_,
		_w14890_,
		_w14891_
	);
	LUT2 #(
		.INIT('h4)
	) name14360 (
		_w14830_,
		_w14891_,
		_w14892_
	);
	LUT2 #(
		.INIT('h4)
	) name14361 (
		_w14864_,
		_w14892_,
		_w14893_
	);
	LUT2 #(
		.INIT('h4)
	) name14362 (
		_w14888_,
		_w14893_,
		_w14894_
	);
	LUT2 #(
		.INIT('h2)
	) name14363 (
		_w14729_,
		_w14894_,
		_w14895_
	);
	LUT2 #(
		.INIT('h4)
	) name14364 (
		_w14729_,
		_w14894_,
		_w14896_
	);
	LUT2 #(
		.INIT('h1)
	) name14365 (
		_w14895_,
		_w14896_,
		_w14897_
	);
	LUT2 #(
		.INIT('h4)
	) name14366 (
		\sa00_reg[2]/P0001 ,
		_w12612_,
		_w14898_
	);
	LUT2 #(
		.INIT('h1)
	) name14367 (
		_w12633_,
		_w13032_,
		_w14899_
	);
	LUT2 #(
		.INIT('h2)
	) name14368 (
		\sa00_reg[2]/P0001 ,
		_w14899_,
		_w14900_
	);
	LUT2 #(
		.INIT('h1)
	) name14369 (
		_w11993_,
		_w12046_,
		_w14901_
	);
	LUT2 #(
		.INIT('h1)
	) name14370 (
		_w13593_,
		_w14898_,
		_w14902_
	);
	LUT2 #(
		.INIT('h8)
	) name14371 (
		_w14901_,
		_w14902_,
		_w14903_
	);
	LUT2 #(
		.INIT('h4)
	) name14372 (
		_w14900_,
		_w14903_,
		_w14904_
	);
	LUT2 #(
		.INIT('h2)
	) name14373 (
		\sa00_reg[1]/P0001 ,
		_w14904_,
		_w14905_
	);
	LUT2 #(
		.INIT('h8)
	) name14374 (
		_w12054_,
		_w12633_,
		_w14906_
	);
	LUT2 #(
		.INIT('h1)
	) name14375 (
		\sa00_reg[2]/P0001 ,
		_w12996_,
		_w14907_
	);
	LUT2 #(
		.INIT('h4)
	) name14376 (
		_w11985_,
		_w12080_,
		_w14908_
	);
	LUT2 #(
		.INIT('h2)
	) name14377 (
		\sa00_reg[7]/NET0131 ,
		_w11960_,
		_w14909_
	);
	LUT2 #(
		.INIT('h8)
	) name14378 (
		_w12056_,
		_w14909_,
		_w14910_
	);
	LUT2 #(
		.INIT('h1)
	) name14379 (
		_w12021_,
		_w13085_,
		_w14911_
	);
	LUT2 #(
		.INIT('h1)
	) name14380 (
		_w14908_,
		_w14910_,
		_w14912_
	);
	LUT2 #(
		.INIT('h8)
	) name14381 (
		_w14911_,
		_w14912_,
		_w14913_
	);
	LUT2 #(
		.INIT('h1)
	) name14382 (
		\sa00_reg[1]/P0001 ,
		_w14913_,
		_w14914_
	);
	LUT2 #(
		.INIT('h1)
	) name14383 (
		_w12648_,
		_w13075_,
		_w14915_
	);
	LUT2 #(
		.INIT('h4)
	) name14384 (
		_w14906_,
		_w14915_,
		_w14916_
	);
	LUT2 #(
		.INIT('h4)
	) name14385 (
		_w14907_,
		_w14916_,
		_w14917_
	);
	LUT2 #(
		.INIT('h4)
	) name14386 (
		_w14914_,
		_w14917_,
		_w14918_
	);
	LUT2 #(
		.INIT('h4)
	) name14387 (
		_w14905_,
		_w14918_,
		_w14919_
	);
	LUT2 #(
		.INIT('h1)
	) name14388 (
		\sa00_reg[0]/P0001 ,
		_w14919_,
		_w14920_
	);
	LUT2 #(
		.INIT('h1)
	) name14389 (
		_w12033_,
		_w13580_,
		_w14921_
	);
	LUT2 #(
		.INIT('h1)
	) name14390 (
		\sa00_reg[2]/P0001 ,
		_w14921_,
		_w14922_
	);
	LUT2 #(
		.INIT('h1)
	) name14391 (
		_w11993_,
		_w12651_,
		_w14923_
	);
	LUT2 #(
		.INIT('h4)
	) name14392 (
		_w14290_,
		_w14923_,
		_w14924_
	);
	LUT2 #(
		.INIT('h2)
	) name14393 (
		\sa00_reg[2]/P0001 ,
		_w14924_,
		_w14925_
	);
	LUT2 #(
		.INIT('h1)
	) name14394 (
		_w12691_,
		_w13073_,
		_w14926_
	);
	LUT2 #(
		.INIT('h4)
	) name14395 (
		_w12025_,
		_w14926_,
		_w14927_
	);
	LUT2 #(
		.INIT('h4)
	) name14396 (
		_w14922_,
		_w14927_,
		_w14928_
	);
	LUT2 #(
		.INIT('h4)
	) name14397 (
		_w14925_,
		_w14928_,
		_w14929_
	);
	LUT2 #(
		.INIT('h1)
	) name14398 (
		\sa00_reg[1]/P0001 ,
		_w14929_,
		_w14930_
	);
	LUT2 #(
		.INIT('h1)
	) name14399 (
		_w12655_,
		_w14244_,
		_w14931_
	);
	LUT2 #(
		.INIT('h1)
	) name14400 (
		_w13629_,
		_w14931_,
		_w14932_
	);
	LUT2 #(
		.INIT('h2)
	) name14401 (
		\sa00_reg[2]/P0001 ,
		_w14932_,
		_w14933_
	);
	LUT2 #(
		.INIT('h4)
	) name14402 (
		\sa00_reg[2]/P0001 ,
		_w14301_,
		_w14934_
	);
	LUT2 #(
		.INIT('h1)
	) name14403 (
		_w11976_,
		_w12003_,
		_w14935_
	);
	LUT2 #(
		.INIT('h4)
	) name14404 (
		_w14390_,
		_w14935_,
		_w14936_
	);
	LUT2 #(
		.INIT('h1)
	) name14405 (
		_w14232_,
		_w14934_,
		_w14937_
	);
	LUT2 #(
		.INIT('h8)
	) name14406 (
		_w14936_,
		_w14937_,
		_w14938_
	);
	LUT2 #(
		.INIT('h4)
	) name14407 (
		_w14933_,
		_w14938_,
		_w14939_
	);
	LUT2 #(
		.INIT('h2)
	) name14408 (
		\sa00_reg[1]/P0001 ,
		_w14939_,
		_w14940_
	);
	LUT2 #(
		.INIT('h4)
	) name14409 (
		_w12021_,
		_w14270_,
		_w14941_
	);
	LUT2 #(
		.INIT('h1)
	) name14410 (
		\sa00_reg[2]/P0001 ,
		_w14941_,
		_w14942_
	);
	LUT2 #(
		.INIT('h4)
	) name14411 (
		_w12613_,
		_w12687_,
		_w14943_
	);
	LUT2 #(
		.INIT('h8)
	) name14412 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w14944_
	);
	LUT2 #(
		.INIT('h4)
	) name14413 (
		_w14943_,
		_w14944_,
		_w14945_
	);
	LUT2 #(
		.INIT('h1)
	) name14414 (
		_w12652_,
		_w14945_,
		_w14946_
	);
	LUT2 #(
		.INIT('h4)
	) name14415 (
		_w14942_,
		_w14946_,
		_w14947_
	);
	LUT2 #(
		.INIT('h4)
	) name14416 (
		_w14930_,
		_w14947_,
		_w14948_
	);
	LUT2 #(
		.INIT('h4)
	) name14417 (
		_w14940_,
		_w14948_,
		_w14949_
	);
	LUT2 #(
		.INIT('h2)
	) name14418 (
		\sa00_reg[0]/P0001 ,
		_w14949_,
		_w14950_
	);
	LUT2 #(
		.INIT('h1)
	) name14419 (
		_w11963_,
		_w12612_,
		_w14951_
	);
	LUT2 #(
		.INIT('h4)
	) name14420 (
		_w13028_,
		_w14951_,
		_w14952_
	);
	LUT2 #(
		.INIT('h2)
	) name14421 (
		_w14246_,
		_w14952_,
		_w14953_
	);
	LUT2 #(
		.INIT('h1)
	) name14422 (
		_w11977_,
		_w14751_,
		_w14954_
	);
	LUT2 #(
		.INIT('h4)
	) name14423 (
		_w14953_,
		_w14954_,
		_w14955_
	);
	LUT2 #(
		.INIT('h2)
	) name14424 (
		\sa00_reg[1]/P0001 ,
		_w14955_,
		_w14956_
	);
	LUT2 #(
		.INIT('h1)
	) name14425 (
		_w11958_,
		_w12648_,
		_w14957_
	);
	LUT2 #(
		.INIT('h2)
	) name14426 (
		_w13015_,
		_w14957_,
		_w14958_
	);
	LUT2 #(
		.INIT('h1)
	) name14427 (
		_w12094_,
		_w12659_,
		_w14959_
	);
	LUT2 #(
		.INIT('h8)
	) name14428 (
		_w11980_,
		_w14959_,
		_w14960_
	);
	LUT2 #(
		.INIT('h8)
	) name14429 (
		\sa00_reg[6]/NET0131 ,
		_w12660_,
		_w14961_
	);
	LUT2 #(
		.INIT('h1)
	) name14430 (
		_w12003_,
		_w14961_,
		_w14962_
	);
	LUT2 #(
		.INIT('h2)
	) name14431 (
		_w13571_,
		_w14962_,
		_w14963_
	);
	LUT2 #(
		.INIT('h1)
	) name14432 (
		_w13581_,
		_w14960_,
		_w14964_
	);
	LUT2 #(
		.INIT('h4)
	) name14433 (
		_w13625_,
		_w14964_,
		_w14965_
	);
	LUT2 #(
		.INIT('h4)
	) name14434 (
		_w14958_,
		_w14965_,
		_w14966_
	);
	LUT2 #(
		.INIT('h4)
	) name14435 (
		_w14963_,
		_w14966_,
		_w14967_
	);
	LUT2 #(
		.INIT('h4)
	) name14436 (
		_w14956_,
		_w14967_,
		_w14968_
	);
	LUT2 #(
		.INIT('h4)
	) name14437 (
		_w14920_,
		_w14968_,
		_w14969_
	);
	LUT2 #(
		.INIT('h4)
	) name14438 (
		_w14950_,
		_w14969_,
		_w14970_
	);
	LUT2 #(
		.INIT('h2)
	) name14439 (
		_w13558_,
		_w14970_,
		_w14971_
	);
	LUT2 #(
		.INIT('h4)
	) name14440 (
		_w13558_,
		_w14970_,
		_w14972_
	);
	LUT2 #(
		.INIT('h1)
	) name14441 (
		_w14971_,
		_w14972_,
		_w14973_
	);
	LUT2 #(
		.INIT('h8)
	) name14442 (
		_w14897_,
		_w14973_,
		_w14974_
	);
	LUT2 #(
		.INIT('h1)
	) name14443 (
		_w14897_,
		_w14973_,
		_w14975_
	);
	LUT2 #(
		.INIT('h1)
	) name14444 (
		_w14974_,
		_w14975_,
		_w14976_
	);
	LUT2 #(
		.INIT('h1)
	) name14445 (
		_w14825_,
		_w14976_,
		_w14977_
	);
	LUT2 #(
		.INIT('h8)
	) name14446 (
		_w14825_,
		_w14976_,
		_w14978_
	);
	LUT2 #(
		.INIT('h1)
	) name14447 (
		\ld_r_reg/P0001 ,
		_w14977_,
		_w14979_
	);
	LUT2 #(
		.INIT('h4)
	) name14448 (
		_w14978_,
		_w14979_,
		_w14980_
	);
	LUT2 #(
		.INIT('h2)
	) name14449 (
		\text_in_r_reg[115]/P0001 ,
		\u0_w_reg[0][19]/P0001 ,
		_w14981_
	);
	LUT2 #(
		.INIT('h4)
	) name14450 (
		\text_in_r_reg[115]/P0001 ,
		\u0_w_reg[0][19]/P0001 ,
		_w14982_
	);
	LUT2 #(
		.INIT('h2)
	) name14451 (
		\ld_r_reg/P0001 ,
		_w14981_,
		_w14983_
	);
	LUT2 #(
		.INIT('h4)
	) name14452 (
		_w14982_,
		_w14983_,
		_w14984_
	);
	LUT2 #(
		.INIT('h1)
	) name14453 (
		_w14980_,
		_w14984_,
		_w14985_
	);
	LUT2 #(
		.INIT('h2)
	) name14454 (
		_w14491_,
		_w14970_,
		_w14986_
	);
	LUT2 #(
		.INIT('h4)
	) name14455 (
		_w14491_,
		_w14970_,
		_w14987_
	);
	LUT2 #(
		.INIT('h1)
	) name14456 (
		_w14986_,
		_w14987_,
		_w14988_
	);
	LUT2 #(
		.INIT('h2)
	) name14457 (
		_w13922_,
		_w14894_,
		_w14989_
	);
	LUT2 #(
		.INIT('h4)
	) name14458 (
		_w13922_,
		_w14894_,
		_w14990_
	);
	LUT2 #(
		.INIT('h1)
	) name14459 (
		_w14989_,
		_w14990_,
		_w14991_
	);
	LUT2 #(
		.INIT('h8)
	) name14460 (
		_w14988_,
		_w14991_,
		_w14992_
	);
	LUT2 #(
		.INIT('h1)
	) name14461 (
		_w14988_,
		_w14991_,
		_w14993_
	);
	LUT2 #(
		.INIT('h1)
	) name14462 (
		_w14992_,
		_w14993_,
		_w14994_
	);
	LUT2 #(
		.INIT('h2)
	) name14463 (
		_w14033_,
		_w14651_,
		_w14995_
	);
	LUT2 #(
		.INIT('h4)
	) name14464 (
		_w14033_,
		_w14651_,
		_w14996_
	);
	LUT2 #(
		.INIT('h1)
	) name14465 (
		_w14995_,
		_w14996_,
		_w14997_
	);
	LUT2 #(
		.INIT('h8)
	) name14466 (
		\sa33_reg[2]/P0001 ,
		_w12445_,
		_w14998_
	);
	LUT2 #(
		.INIT('h8)
	) name14467 (
		_w13690_,
		_w14034_,
		_w14999_
	);
	LUT2 #(
		.INIT('h2)
	) name14468 (
		\sa33_reg[1]/P0001 ,
		_w14106_,
		_w15000_
	);
	LUT2 #(
		.INIT('h1)
	) name14469 (
		_w14998_,
		_w14999_,
		_w15001_
	);
	LUT2 #(
		.INIT('h8)
	) name14470 (
		_w15000_,
		_w15001_,
		_w15002_
	);
	LUT2 #(
		.INIT('h8)
	) name14471 (
		\sa33_reg[2]/P0001 ,
		_w12414_,
		_w15003_
	);
	LUT2 #(
		.INIT('h4)
	) name14472 (
		_w12426_,
		_w15003_,
		_w15004_
	);
	LUT2 #(
		.INIT('h8)
	) name14473 (
		_w12884_,
		_w13986_,
		_w15005_
	);
	LUT2 #(
		.INIT('h1)
	) name14474 (
		_w12872_,
		_w14052_,
		_w15006_
	);
	LUT2 #(
		.INIT('h4)
	) name14475 (
		_w12523_,
		_w15006_,
		_w15007_
	);
	LUT2 #(
		.INIT('h2)
	) name14476 (
		_w12879_,
		_w12912_,
		_w15008_
	);
	LUT2 #(
		.INIT('h1)
	) name14477 (
		_w15004_,
		_w15005_,
		_w15009_
	);
	LUT2 #(
		.INIT('h8)
	) name14478 (
		_w15008_,
		_w15009_,
		_w15010_
	);
	LUT2 #(
		.INIT('h8)
	) name14479 (
		_w15007_,
		_w15010_,
		_w15011_
	);
	LUT2 #(
		.INIT('h1)
	) name14480 (
		_w15002_,
		_w15011_,
		_w15012_
	);
	LUT2 #(
		.INIT('h1)
	) name14481 (
		_w12481_,
		_w13698_,
		_w15013_
	);
	LUT2 #(
		.INIT('h4)
	) name14482 (
		_w13667_,
		_w15013_,
		_w15014_
	);
	LUT2 #(
		.INIT('h2)
	) name14483 (
		_w12560_,
		_w15014_,
		_w15015_
	);
	LUT2 #(
		.INIT('h2)
	) name14484 (
		\sa33_reg[0]/P0001 ,
		_w12909_,
		_w15016_
	);
	LUT2 #(
		.INIT('h1)
	) name14485 (
		_w12910_,
		_w13702_,
		_w15017_
	);
	LUT2 #(
		.INIT('h8)
	) name14486 (
		_w15016_,
		_w15017_,
		_w15018_
	);
	LUT2 #(
		.INIT('h4)
	) name14487 (
		_w15015_,
		_w15018_,
		_w15019_
	);
	LUT2 #(
		.INIT('h4)
	) name14488 (
		_w15012_,
		_w15019_,
		_w15020_
	);
	LUT2 #(
		.INIT('h1)
	) name14489 (
		_w12444_,
		_w12877_,
		_w15021_
	);
	LUT2 #(
		.INIT('h1)
	) name14490 (
		\sa33_reg[2]/P0001 ,
		_w12510_,
		_w15022_
	);
	LUT2 #(
		.INIT('h4)
	) name14491 (
		_w15021_,
		_w15022_,
		_w15023_
	);
	LUT2 #(
		.INIT('h1)
	) name14492 (
		_w12864_,
		_w13986_,
		_w15024_
	);
	LUT2 #(
		.INIT('h2)
	) name14493 (
		\sa33_reg[2]/P0001 ,
		_w15024_,
		_w15025_
	);
	LUT2 #(
		.INIT('h2)
	) name14494 (
		\sa33_reg[1]/P0001 ,
		_w13668_,
		_w15026_
	);
	LUT2 #(
		.INIT('h4)
	) name14495 (
		_w15023_,
		_w15026_,
		_w15027_
	);
	LUT2 #(
		.INIT('h4)
	) name14496 (
		_w15025_,
		_w15027_,
		_w15028_
	);
	LUT2 #(
		.INIT('h8)
	) name14497 (
		_w12456_,
		_w12510_,
		_w15029_
	);
	LUT2 #(
		.INIT('h1)
	) name14498 (
		\sa33_reg[1]/P0001 ,
		_w12506_,
		_w15030_
	);
	LUT2 #(
		.INIT('h4)
	) name14499 (
		_w15029_,
		_w15030_,
		_w15031_
	);
	LUT2 #(
		.INIT('h1)
	) name14500 (
		_w15028_,
		_w15031_,
		_w15032_
	);
	LUT2 #(
		.INIT('h8)
	) name14501 (
		_w12565_,
		_w12881_,
		_w15033_
	);
	LUT2 #(
		.INIT('h8)
	) name14502 (
		_w12861_,
		_w14595_,
		_w15034_
	);
	LUT2 #(
		.INIT('h1)
	) name14503 (
		\sa33_reg[0]/P0001 ,
		_w12468_,
		_w15035_
	);
	LUT2 #(
		.INIT('h4)
	) name14504 (
		_w15033_,
		_w15035_,
		_w15036_
	);
	LUT2 #(
		.INIT('h4)
	) name14505 (
		_w15034_,
		_w15036_,
		_w15037_
	);
	LUT2 #(
		.INIT('h4)
	) name14506 (
		_w15032_,
		_w15037_,
		_w15038_
	);
	LUT2 #(
		.INIT('h1)
	) name14507 (
		_w15020_,
		_w15038_,
		_w15039_
	);
	LUT2 #(
		.INIT('h1)
	) name14508 (
		_w12461_,
		_w12561_,
		_w15040_
	);
	LUT2 #(
		.INIT('h8)
	) name14509 (
		\sa33_reg[2]/P0001 ,
		_w12479_,
		_w15041_
	);
	LUT2 #(
		.INIT('h4)
	) name14510 (
		_w15040_,
		_w15041_,
		_w15042_
	);
	LUT2 #(
		.INIT('h8)
	) name14511 (
		_w12409_,
		_w12419_,
		_w15043_
	);
	LUT2 #(
		.INIT('h1)
	) name14512 (
		\sa33_reg[2]/P0001 ,
		_w14023_,
		_w15044_
	);
	LUT2 #(
		.INIT('h4)
	) name14513 (
		_w15043_,
		_w15044_,
		_w15045_
	);
	LUT2 #(
		.INIT('h1)
	) name14514 (
		_w12550_,
		_w12912_,
		_w15046_
	);
	LUT2 #(
		.INIT('h8)
	) name14515 (
		_w15045_,
		_w15046_,
		_w15047_
	);
	LUT2 #(
		.INIT('h2)
	) name14516 (
		\sa33_reg[2]/P0001 ,
		_w12427_,
		_w15048_
	);
	LUT2 #(
		.INIT('h4)
	) name14517 (
		_w12506_,
		_w15048_,
		_w15049_
	);
	LUT2 #(
		.INIT('h4)
	) name14518 (
		_w12919_,
		_w15049_,
		_w15050_
	);
	LUT2 #(
		.INIT('h1)
	) name14519 (
		_w15047_,
		_w15050_,
		_w15051_
	);
	LUT2 #(
		.INIT('h1)
	) name14520 (
		\sa33_reg[1]/P0001 ,
		_w14012_,
		_w15052_
	);
	LUT2 #(
		.INIT('h4)
	) name14521 (
		_w14044_,
		_w15052_,
		_w15053_
	);
	LUT2 #(
		.INIT('h4)
	) name14522 (
		_w15051_,
		_w15053_,
		_w15054_
	);
	LUT2 #(
		.INIT('h8)
	) name14523 (
		\sa33_reg[5]/P0001 ,
		_w14091_,
		_w15055_
	);
	LUT2 #(
		.INIT('h1)
	) name14524 (
		_w14624_,
		_w15055_,
		_w15056_
	);
	LUT2 #(
		.INIT('h2)
	) name14525 (
		\sa33_reg[6]/P0001 ,
		_w15056_,
		_w15057_
	);
	LUT2 #(
		.INIT('h1)
	) name14526 (
		_w12522_,
		_w12551_,
		_w15058_
	);
	LUT2 #(
		.INIT('h2)
	) name14527 (
		\sa33_reg[2]/P0001 ,
		_w15058_,
		_w15059_
	);
	LUT2 #(
		.INIT('h2)
	) name14528 (
		\sa33_reg[1]/P0001 ,
		_w12463_,
		_w15060_
	);
	LUT2 #(
		.INIT('h1)
	) name14529 (
		_w12564_,
		_w14048_,
		_w15061_
	);
	LUT2 #(
		.INIT('h8)
	) name14530 (
		_w15060_,
		_w15061_,
		_w15062_
	);
	LUT2 #(
		.INIT('h4)
	) name14531 (
		_w15059_,
		_w15062_,
		_w15063_
	);
	LUT2 #(
		.INIT('h4)
	) name14532 (
		_w15057_,
		_w15063_,
		_w15064_
	);
	LUT2 #(
		.INIT('h1)
	) name14533 (
		_w15054_,
		_w15064_,
		_w15065_
	);
	LUT2 #(
		.INIT('h1)
	) name14534 (
		_w14632_,
		_w15042_,
		_w15066_
	);
	LUT2 #(
		.INIT('h4)
	) name14535 (
		_w15065_,
		_w15066_,
		_w15067_
	);
	LUT2 #(
		.INIT('h4)
	) name14536 (
		_w15039_,
		_w15067_,
		_w15068_
	);
	LUT2 #(
		.INIT('h2)
	) name14537 (
		\u0_w_reg[0][11]/P0001 ,
		_w15068_,
		_w15069_
	);
	LUT2 #(
		.INIT('h4)
	) name14538 (
		\u0_w_reg[0][11]/P0001 ,
		_w15068_,
		_w15070_
	);
	LUT2 #(
		.INIT('h1)
	) name14539 (
		_w15069_,
		_w15070_,
		_w15071_
	);
	LUT2 #(
		.INIT('h8)
	) name14540 (
		_w14997_,
		_w15071_,
		_w15072_
	);
	LUT2 #(
		.INIT('h1)
	) name14541 (
		_w14997_,
		_w15071_,
		_w15073_
	);
	LUT2 #(
		.INIT('h1)
	) name14542 (
		_w15072_,
		_w15073_,
		_w15074_
	);
	LUT2 #(
		.INIT('h1)
	) name14543 (
		_w14994_,
		_w15074_,
		_w15075_
	);
	LUT2 #(
		.INIT('h8)
	) name14544 (
		_w14994_,
		_w15074_,
		_w15076_
	);
	LUT2 #(
		.INIT('h1)
	) name14545 (
		\ld_r_reg/P0001 ,
		_w15075_,
		_w15077_
	);
	LUT2 #(
		.INIT('h4)
	) name14546 (
		_w15076_,
		_w15077_,
		_w15078_
	);
	LUT2 #(
		.INIT('h2)
	) name14547 (
		\text_in_r_reg[107]/P0001 ,
		\u0_w_reg[0][11]/P0001 ,
		_w15079_
	);
	LUT2 #(
		.INIT('h4)
	) name14548 (
		\text_in_r_reg[107]/P0001 ,
		\u0_w_reg[0][11]/P0001 ,
		_w15080_
	);
	LUT2 #(
		.INIT('h2)
	) name14549 (
		\ld_r_reg/P0001 ,
		_w15079_,
		_w15081_
	);
	LUT2 #(
		.INIT('h4)
	) name14550 (
		_w15080_,
		_w15081_,
		_w15082_
	);
	LUT2 #(
		.INIT('h1)
	) name14551 (
		_w15078_,
		_w15082_,
		_w15083_
	);
	LUT2 #(
		.INIT('h2)
	) name14552 (
		\u0_w_reg[0][12]/P0001 ,
		_w12962_,
		_w15084_
	);
	LUT2 #(
		.INIT('h4)
	) name14553 (
		\u0_w_reg[0][12]/P0001 ,
		_w12962_,
		_w15085_
	);
	LUT2 #(
		.INIT('h1)
	) name14554 (
		_w15084_,
		_w15085_,
		_w15086_
	);
	LUT2 #(
		.INIT('h8)
	) name14555 (
		_w14997_,
		_w15086_,
		_w15087_
	);
	LUT2 #(
		.INIT('h1)
	) name14556 (
		_w14997_,
		_w15086_,
		_w15088_
	);
	LUT2 #(
		.INIT('h1)
	) name14557 (
		_w15087_,
		_w15088_,
		_w15089_
	);
	LUT2 #(
		.INIT('h8)
	) name14558 (
		_w12114_,
		_w14819_,
		_w15090_
	);
	LUT2 #(
		.INIT('h1)
	) name14559 (
		_w12114_,
		_w14819_,
		_w15091_
	);
	LUT2 #(
		.INIT('h1)
	) name14560 (
		_w15090_,
		_w15091_,
		_w15092_
	);
	LUT2 #(
		.INIT('h1)
	) name14561 (
		_w15089_,
		_w15092_,
		_w15093_
	);
	LUT2 #(
		.INIT('h8)
	) name14562 (
		_w15089_,
		_w15092_,
		_w15094_
	);
	LUT2 #(
		.INIT('h1)
	) name14563 (
		\ld_r_reg/P0001 ,
		_w15093_,
		_w15095_
	);
	LUT2 #(
		.INIT('h4)
	) name14564 (
		_w15094_,
		_w15095_,
		_w15096_
	);
	LUT2 #(
		.INIT('h2)
	) name14565 (
		\text_in_r_reg[108]/P0001 ,
		\u0_w_reg[0][12]/P0001 ,
		_w15097_
	);
	LUT2 #(
		.INIT('h4)
	) name14566 (
		\text_in_r_reg[108]/P0001 ,
		\u0_w_reg[0][12]/P0001 ,
		_w15098_
	);
	LUT2 #(
		.INIT('h2)
	) name14567 (
		\ld_r_reg/P0001 ,
		_w15097_,
		_w15099_
	);
	LUT2 #(
		.INIT('h4)
	) name14568 (
		_w15098_,
		_w15099_,
		_w15100_
	);
	LUT2 #(
		.INIT('h1)
	) name14569 (
		_w15096_,
		_w15100_,
		_w15101_
	);
	LUT2 #(
		.INIT('h2)
	) name14570 (
		\u0_w_reg[0][4]/P0001 ,
		_w12827_,
		_w15102_
	);
	LUT2 #(
		.INIT('h4)
	) name14571 (
		\u0_w_reg[0][4]/P0001 ,
		_w12827_,
		_w15103_
	);
	LUT2 #(
		.INIT('h1)
	) name14572 (
		_w15102_,
		_w15103_,
		_w15104_
	);
	LUT2 #(
		.INIT('h8)
	) name14573 (
		_w14997_,
		_w15104_,
		_w15105_
	);
	LUT2 #(
		.INIT('h1)
	) name14574 (
		_w14997_,
		_w15104_,
		_w15106_
	);
	LUT2 #(
		.INIT('h1)
	) name14575 (
		_w15105_,
		_w15106_,
		_w15107_
	);
	LUT2 #(
		.INIT('h2)
	) name14576 (
		_w14400_,
		_w14970_,
		_w15108_
	);
	LUT2 #(
		.INIT('h4)
	) name14577 (
		_w14400_,
		_w14970_,
		_w15109_
	);
	LUT2 #(
		.INIT('h1)
	) name14578 (
		_w15108_,
		_w15109_,
		_w15110_
	);
	LUT2 #(
		.INIT('h8)
	) name14579 (
		_w12114_,
		_w15110_,
		_w15111_
	);
	LUT2 #(
		.INIT('h1)
	) name14580 (
		_w12114_,
		_w15110_,
		_w15112_
	);
	LUT2 #(
		.INIT('h1)
	) name14581 (
		_w15111_,
		_w15112_,
		_w15113_
	);
	LUT2 #(
		.INIT('h1)
	) name14582 (
		_w15107_,
		_w15113_,
		_w15114_
	);
	LUT2 #(
		.INIT('h8)
	) name14583 (
		_w15107_,
		_w15113_,
		_w15115_
	);
	LUT2 #(
		.INIT('h1)
	) name14584 (
		\ld_r_reg/P0001 ,
		_w15114_,
		_w15116_
	);
	LUT2 #(
		.INIT('h4)
	) name14585 (
		_w15115_,
		_w15116_,
		_w15117_
	);
	LUT2 #(
		.INIT('h2)
	) name14586 (
		\text_in_r_reg[100]/P0001 ,
		\u0_w_reg[0][4]/P0001 ,
		_w15118_
	);
	LUT2 #(
		.INIT('h4)
	) name14587 (
		\text_in_r_reg[100]/P0001 ,
		\u0_w_reg[0][4]/P0001 ,
		_w15119_
	);
	LUT2 #(
		.INIT('h2)
	) name14588 (
		\ld_r_reg/P0001 ,
		_w15118_,
		_w15120_
	);
	LUT2 #(
		.INIT('h4)
	) name14589 (
		_w15119_,
		_w15120_,
		_w15121_
	);
	LUT2 #(
		.INIT('h1)
	) name14590 (
		_w15117_,
		_w15121_,
		_w15122_
	);
	LUT2 #(
		.INIT('h2)
	) name14591 (
		\u0_w_reg[0][25]/P0001 ,
		_w14210_,
		_w15123_
	);
	LUT2 #(
		.INIT('h4)
	) name14592 (
		\u0_w_reg[0][25]/P0001 ,
		_w14210_,
		_w15124_
	);
	LUT2 #(
		.INIT('h1)
	) name14593 (
		_w15123_,
		_w15124_,
		_w15125_
	);
	LUT2 #(
		.INIT('h8)
	) name14594 (
		_w13838_,
		_w15125_,
		_w15126_
	);
	LUT2 #(
		.INIT('h1)
	) name14595 (
		_w13838_,
		_w15125_,
		_w15127_
	);
	LUT2 #(
		.INIT('h1)
	) name14596 (
		_w15126_,
		_w15127_,
		_w15128_
	);
	LUT2 #(
		.INIT('h2)
	) name14597 (
		_w13465_,
		_w14316_,
		_w15129_
	);
	LUT2 #(
		.INIT('h4)
	) name14598 (
		_w13465_,
		_w14316_,
		_w15130_
	);
	LUT2 #(
		.INIT('h1)
	) name14599 (
		_w15129_,
		_w15130_,
		_w15131_
	);
	LUT2 #(
		.INIT('h2)
	) name14600 (
		_w14660_,
		_w15131_,
		_w15132_
	);
	LUT2 #(
		.INIT('h4)
	) name14601 (
		_w14660_,
		_w15131_,
		_w15133_
	);
	LUT2 #(
		.INIT('h1)
	) name14602 (
		_w15132_,
		_w15133_,
		_w15134_
	);
	LUT2 #(
		.INIT('h1)
	) name14603 (
		_w15128_,
		_w15134_,
		_w15135_
	);
	LUT2 #(
		.INIT('h8)
	) name14604 (
		_w15128_,
		_w15134_,
		_w15136_
	);
	LUT2 #(
		.INIT('h1)
	) name14605 (
		\ld_r_reg/P0001 ,
		_w15135_,
		_w15137_
	);
	LUT2 #(
		.INIT('h4)
	) name14606 (
		_w15136_,
		_w15137_,
		_w15138_
	);
	LUT2 #(
		.INIT('h1)
	) name14607 (
		\text_in_r_reg[121]/P0001 ,
		\u0_w_reg[0][25]/P0001 ,
		_w15139_
	);
	LUT2 #(
		.INIT('h8)
	) name14608 (
		\text_in_r_reg[121]/P0001 ,
		\u0_w_reg[0][25]/P0001 ,
		_w15140_
	);
	LUT2 #(
		.INIT('h2)
	) name14609 (
		\ld_r_reg/P0001 ,
		_w15139_,
		_w15141_
	);
	LUT2 #(
		.INIT('h4)
	) name14610 (
		_w15140_,
		_w15141_,
		_w15142_
	);
	LUT2 #(
		.INIT('h1)
	) name14611 (
		_w15138_,
		_w15142_,
		_w15143_
	);
	LUT2 #(
		.INIT('h2)
	) name14612 (
		\u0_w_reg[0][28]/P0001 ,
		_w12962_,
		_w15144_
	);
	LUT2 #(
		.INIT('h4)
	) name14613 (
		\u0_w_reg[0][28]/P0001 ,
		_w12962_,
		_w15145_
	);
	LUT2 #(
		.INIT('h1)
	) name14614 (
		_w15144_,
		_w15145_,
		_w15146_
	);
	LUT2 #(
		.INIT('h8)
	) name14615 (
		_w12830_,
		_w15146_,
		_w15147_
	);
	LUT2 #(
		.INIT('h1)
	) name14616 (
		_w12830_,
		_w15146_,
		_w15148_
	);
	LUT2 #(
		.INIT('h1)
	) name14617 (
		_w15147_,
		_w15148_,
		_w15149_
	);
	LUT2 #(
		.INIT('h4)
	) name14618 (
		_w14660_,
		_w14988_,
		_w15150_
	);
	LUT2 #(
		.INIT('h2)
	) name14619 (
		_w14660_,
		_w14988_,
		_w15151_
	);
	LUT2 #(
		.INIT('h1)
	) name14620 (
		_w15150_,
		_w15151_,
		_w15152_
	);
	LUT2 #(
		.INIT('h2)
	) name14621 (
		_w15149_,
		_w15152_,
		_w15153_
	);
	LUT2 #(
		.INIT('h4)
	) name14622 (
		_w15149_,
		_w15152_,
		_w15154_
	);
	LUT2 #(
		.INIT('h1)
	) name14623 (
		\ld_r_reg/P0001 ,
		_w15153_,
		_w15155_
	);
	LUT2 #(
		.INIT('h4)
	) name14624 (
		_w15154_,
		_w15155_,
		_w15156_
	);
	LUT2 #(
		.INIT('h2)
	) name14625 (
		\text_in_r_reg[124]/P0001 ,
		\u0_w_reg[0][28]/P0001 ,
		_w15157_
	);
	LUT2 #(
		.INIT('h4)
	) name14626 (
		\text_in_r_reg[124]/P0001 ,
		\u0_w_reg[0][28]/P0001 ,
		_w15158_
	);
	LUT2 #(
		.INIT('h2)
	) name14627 (
		\ld_r_reg/P0001 ,
		_w15157_,
		_w15159_
	);
	LUT2 #(
		.INIT('h4)
	) name14628 (
		_w15158_,
		_w15159_,
		_w15160_
	);
	LUT2 #(
		.INIT('h1)
	) name14629 (
		_w15156_,
		_w15160_,
		_w15161_
	);
	LUT2 #(
		.INIT('h1)
	) name14630 (
		\u0_w_reg[0][24]/P0001 ,
		_w14113_,
		_w15162_
	);
	LUT2 #(
		.INIT('h8)
	) name14631 (
		\u0_w_reg[0][24]/P0001 ,
		_w14113_,
		_w15163_
	);
	LUT2 #(
		.INIT('h1)
	) name14632 (
		_w15162_,
		_w15163_,
		_w15164_
	);
	LUT2 #(
		.INIT('h4)
	) name14633 (
		_w13468_,
		_w14660_,
		_w15165_
	);
	LUT2 #(
		.INIT('h2)
	) name14634 (
		_w13468_,
		_w14660_,
		_w15166_
	);
	LUT2 #(
		.INIT('h1)
	) name14635 (
		_w15165_,
		_w15166_,
		_w15167_
	);
	LUT2 #(
		.INIT('h1)
	) name14636 (
		_w15164_,
		_w15167_,
		_w15168_
	);
	LUT2 #(
		.INIT('h8)
	) name14637 (
		_w15164_,
		_w15167_,
		_w15169_
	);
	LUT2 #(
		.INIT('h1)
	) name14638 (
		\ld_r_reg/P0001 ,
		_w15168_,
		_w15170_
	);
	LUT2 #(
		.INIT('h4)
	) name14639 (
		_w15169_,
		_w15170_,
		_w15171_
	);
	LUT2 #(
		.INIT('h1)
	) name14640 (
		\text_in_r_reg[120]/P0001 ,
		\u0_w_reg[0][24]/P0001 ,
		_w15172_
	);
	LUT2 #(
		.INIT('h8)
	) name14641 (
		\text_in_r_reg[120]/P0001 ,
		\u0_w_reg[0][24]/P0001 ,
		_w15173_
	);
	LUT2 #(
		.INIT('h2)
	) name14642 (
		\ld_r_reg/P0001 ,
		_w15172_,
		_w15174_
	);
	LUT2 #(
		.INIT('h4)
	) name14643 (
		_w15173_,
		_w15174_,
		_w15175_
	);
	LUT2 #(
		.INIT('h1)
	) name14644 (
		_w15171_,
		_w15175_,
		_w15176_
	);
	LUT2 #(
		.INIT('h1)
	) name14645 (
		\u0_w_reg[0][16]/P0001 ,
		_w14113_,
		_w15177_
	);
	LUT2 #(
		.INIT('h8)
	) name14646 (
		\u0_w_reg[0][16]/P0001 ,
		_w14113_,
		_w15178_
	);
	LUT2 #(
		.INIT('h1)
	) name14647 (
		_w15177_,
		_w15178_,
		_w15179_
	);
	LUT2 #(
		.INIT('h2)
	) name14648 (
		_w13558_,
		_w14316_,
		_w15180_
	);
	LUT2 #(
		.INIT('h4)
	) name14649 (
		_w13558_,
		_w14316_,
		_w15181_
	);
	LUT2 #(
		.INIT('h1)
	) name14650 (
		_w15180_,
		_w15181_,
		_w15182_
	);
	LUT2 #(
		.INIT('h8)
	) name14651 (
		_w14125_,
		_w15182_,
		_w15183_
	);
	LUT2 #(
		.INIT('h1)
	) name14652 (
		_w14125_,
		_w15182_,
		_w15184_
	);
	LUT2 #(
		.INIT('h1)
	) name14653 (
		_w15183_,
		_w15184_,
		_w15185_
	);
	LUT2 #(
		.INIT('h4)
	) name14654 (
		_w15179_,
		_w15185_,
		_w15186_
	);
	LUT2 #(
		.INIT('h2)
	) name14655 (
		_w15179_,
		_w15185_,
		_w15187_
	);
	LUT2 #(
		.INIT('h1)
	) name14656 (
		\ld_r_reg/P0001 ,
		_w15186_,
		_w15188_
	);
	LUT2 #(
		.INIT('h4)
	) name14657 (
		_w15187_,
		_w15188_,
		_w15189_
	);
	LUT2 #(
		.INIT('h1)
	) name14658 (
		\text_in_r_reg[112]/P0001 ,
		\u0_w_reg[0][16]/P0001 ,
		_w15190_
	);
	LUT2 #(
		.INIT('h8)
	) name14659 (
		\text_in_r_reg[112]/P0001 ,
		\u0_w_reg[0][16]/P0001 ,
		_w15191_
	);
	LUT2 #(
		.INIT('h2)
	) name14660 (
		\ld_r_reg/P0001 ,
		_w15190_,
		_w15192_
	);
	LUT2 #(
		.INIT('h4)
	) name14661 (
		_w15191_,
		_w15192_,
		_w15193_
	);
	LUT2 #(
		.INIT('h1)
	) name14662 (
		_w15189_,
		_w15193_,
		_w15194_
	);
	LUT2 #(
		.INIT('h2)
	) name14663 (
		_w12111_,
		_w13558_,
		_w15195_
	);
	LUT2 #(
		.INIT('h4)
	) name14664 (
		_w12111_,
		_w13558_,
		_w15196_
	);
	LUT2 #(
		.INIT('h1)
	) name14665 (
		_w15195_,
		_w15196_,
		_w15197_
	);
	LUT2 #(
		.INIT('h8)
	) name14666 (
		_w14570_,
		_w15197_,
		_w15198_
	);
	LUT2 #(
		.INIT('h1)
	) name14667 (
		_w14570_,
		_w15197_,
		_w15199_
	);
	LUT2 #(
		.INIT('h1)
	) name14668 (
		_w15198_,
		_w15199_,
		_w15200_
	);
	LUT2 #(
		.INIT('h1)
	) name14669 (
		_w12827_,
		_w12962_,
		_w15201_
	);
	LUT2 #(
		.INIT('h8)
	) name14670 (
		_w12827_,
		_w12962_,
		_w15202_
	);
	LUT2 #(
		.INIT('h1)
	) name14671 (
		_w15201_,
		_w15202_,
		_w15203_
	);
	LUT2 #(
		.INIT('h2)
	) name14672 (
		\u0_w_reg[0][20]/P0001 ,
		_w13922_,
		_w15204_
	);
	LUT2 #(
		.INIT('h4)
	) name14673 (
		\u0_w_reg[0][20]/P0001 ,
		_w13922_,
		_w15205_
	);
	LUT2 #(
		.INIT('h1)
	) name14674 (
		_w15204_,
		_w15205_,
		_w15206_
	);
	LUT2 #(
		.INIT('h8)
	) name14675 (
		_w15203_,
		_w15206_,
		_w15207_
	);
	LUT2 #(
		.INIT('h1)
	) name14676 (
		_w15203_,
		_w15206_,
		_w15208_
	);
	LUT2 #(
		.INIT('h1)
	) name14677 (
		_w15207_,
		_w15208_,
		_w15209_
	);
	LUT2 #(
		.INIT('h2)
	) name14678 (
		_w15200_,
		_w15209_,
		_w15210_
	);
	LUT2 #(
		.INIT('h4)
	) name14679 (
		_w15200_,
		_w15209_,
		_w15211_
	);
	LUT2 #(
		.INIT('h1)
	) name14680 (
		\ld_r_reg/P0001 ,
		_w15210_,
		_w15212_
	);
	LUT2 #(
		.INIT('h4)
	) name14681 (
		_w15211_,
		_w15212_,
		_w15213_
	);
	LUT2 #(
		.INIT('h2)
	) name14682 (
		\text_in_r_reg[116]/P0001 ,
		\u0_w_reg[0][20]/P0001 ,
		_w15214_
	);
	LUT2 #(
		.INIT('h4)
	) name14683 (
		\text_in_r_reg[116]/P0001 ,
		\u0_w_reg[0][20]/P0001 ,
		_w15215_
	);
	LUT2 #(
		.INIT('h2)
	) name14684 (
		\ld_r_reg/P0001 ,
		_w15214_,
		_w15216_
	);
	LUT2 #(
		.INIT('h4)
	) name14685 (
		_w15215_,
		_w15216_,
		_w15217_
	);
	LUT2 #(
		.INIT('h1)
	) name14686 (
		_w15213_,
		_w15217_,
		_w15218_
	);
	LUT2 #(
		.INIT('h1)
	) name14687 (
		_w12408_,
		_w13091_,
		_w15219_
	);
	LUT2 #(
		.INIT('h8)
	) name14688 (
		_w12408_,
		_w13091_,
		_w15220_
	);
	LUT2 #(
		.INIT('h1)
	) name14689 (
		_w15219_,
		_w15220_,
		_w15221_
	);
	LUT2 #(
		.INIT('h1)
	) name14690 (
		_w12415_,
		_w12431_,
		_w15222_
	);
	LUT2 #(
		.INIT('h1)
	) name14691 (
		\sa33_reg[2]/P0001 ,
		_w15222_,
		_w15223_
	);
	LUT2 #(
		.INIT('h1)
	) name14692 (
		_w12466_,
		_w12493_,
		_w15224_
	);
	LUT2 #(
		.INIT('h8)
	) name14693 (
		_w14621_,
		_w15224_,
		_w15225_
	);
	LUT2 #(
		.INIT('h2)
	) name14694 (
		\sa33_reg[2]/P0001 ,
		_w15225_,
		_w15226_
	);
	LUT2 #(
		.INIT('h1)
	) name14695 (
		_w12517_,
		_w13939_,
		_w15227_
	);
	LUT2 #(
		.INIT('h2)
	) name14696 (
		\sa33_reg[2]/P0001 ,
		_w15227_,
		_w15228_
	);
	LUT2 #(
		.INIT('h8)
	) name14697 (
		_w12430_,
		_w12881_,
		_w15229_
	);
	LUT2 #(
		.INIT('h1)
	) name14698 (
		_w12468_,
		_w15229_,
		_w15230_
	);
	LUT2 #(
		.INIT('h8)
	) name14699 (
		_w12464_,
		_w15230_,
		_w15231_
	);
	LUT2 #(
		.INIT('h4)
	) name14700 (
		_w15228_,
		_w15231_,
		_w15232_
	);
	LUT2 #(
		.INIT('h1)
	) name14701 (
		\sa33_reg[1]/P0001 ,
		_w15232_,
		_w15233_
	);
	LUT2 #(
		.INIT('h8)
	) name14702 (
		_w13689_,
		_w13952_,
		_w15234_
	);
	LUT2 #(
		.INIT('h1)
	) name14703 (
		_w12411_,
		_w12422_,
		_w15235_
	);
	LUT2 #(
		.INIT('h4)
	) name14704 (
		_w13699_,
		_w15235_,
		_w15236_
	);
	LUT2 #(
		.INIT('h2)
	) name14705 (
		\sa33_reg[2]/P0001 ,
		_w15236_,
		_w15237_
	);
	LUT2 #(
		.INIT('h2)
	) name14706 (
		_w14043_,
		_w15234_,
		_w15238_
	);
	LUT2 #(
		.INIT('h4)
	) name14707 (
		_w15237_,
		_w15238_,
		_w15239_
	);
	LUT2 #(
		.INIT('h2)
	) name14708 (
		\sa33_reg[1]/P0001 ,
		_w15239_,
		_w15240_
	);
	LUT2 #(
		.INIT('h1)
	) name14709 (
		_w15223_,
		_w15226_,
		_w15241_
	);
	LUT2 #(
		.INIT('h4)
	) name14710 (
		_w15233_,
		_w15241_,
		_w15242_
	);
	LUT2 #(
		.INIT('h4)
	) name14711 (
		_w15240_,
		_w15242_,
		_w15243_
	);
	LUT2 #(
		.INIT('h2)
	) name14712 (
		\sa33_reg[0]/P0001 ,
		_w15243_,
		_w15244_
	);
	LUT2 #(
		.INIT('h1)
	) name14713 (
		_w12470_,
		_w14005_,
		_w15245_
	);
	LUT2 #(
		.INIT('h1)
	) name14714 (
		\sa33_reg[4]/P0001 ,
		_w15245_,
		_w15246_
	);
	LUT2 #(
		.INIT('h1)
	) name14715 (
		\sa33_reg[1]/P0001 ,
		_w12415_,
		_w15247_
	);
	LUT2 #(
		.INIT('h4)
	) name14716 (
		_w12562_,
		_w15247_,
		_w15248_
	);
	LUT2 #(
		.INIT('h4)
	) name14717 (
		_w14091_,
		_w15248_,
		_w15249_
	);
	LUT2 #(
		.INIT('h1)
	) name14718 (
		_w12929_,
		_w15246_,
		_w15250_
	);
	LUT2 #(
		.INIT('h8)
	) name14719 (
		_w15249_,
		_w15250_,
		_w15251_
	);
	LUT2 #(
		.INIT('h8)
	) name14720 (
		_w12473_,
		_w12884_,
		_w15252_
	);
	LUT2 #(
		.INIT('h1)
	) name14721 (
		_w13685_,
		_w14603_,
		_w15253_
	);
	LUT2 #(
		.INIT('h2)
	) name14722 (
		_w12472_,
		_w15253_,
		_w15254_
	);
	LUT2 #(
		.INIT('h2)
	) name14723 (
		\sa33_reg[1]/P0001 ,
		_w12550_,
		_w15255_
	);
	LUT2 #(
		.INIT('h4)
	) name14724 (
		_w15252_,
		_w15255_,
		_w15256_
	);
	LUT2 #(
		.INIT('h4)
	) name14725 (
		_w15254_,
		_w15256_,
		_w15257_
	);
	LUT2 #(
		.INIT('h1)
	) name14726 (
		_w15251_,
		_w15257_,
		_w15258_
	);
	LUT2 #(
		.INIT('h2)
	) name14727 (
		_w13735_,
		_w14073_,
		_w15259_
	);
	LUT2 #(
		.INIT('h1)
	) name14728 (
		_w12894_,
		_w13970_,
		_w15260_
	);
	LUT2 #(
		.INIT('h1)
	) name14729 (
		_w12419_,
		_w15260_,
		_w15261_
	);
	LUT2 #(
		.INIT('h4)
	) name14730 (
		_w12570_,
		_w12862_,
		_w15262_
	);
	LUT2 #(
		.INIT('h4)
	) name14731 (
		_w15261_,
		_w15262_,
		_w15263_
	);
	LUT2 #(
		.INIT('h1)
	) name14732 (
		_w15259_,
		_w15263_,
		_w15264_
	);
	LUT2 #(
		.INIT('h1)
	) name14733 (
		_w15258_,
		_w15264_,
		_w15265_
	);
	LUT2 #(
		.INIT('h1)
	) name14734 (
		\sa33_reg[0]/P0001 ,
		_w15265_,
		_w15266_
	);
	LUT2 #(
		.INIT('h2)
	) name14735 (
		\sa33_reg[2]/P0001 ,
		_w12935_,
		_w15267_
	);
	LUT2 #(
		.INIT('h4)
	) name14736 (
		_w14016_,
		_w15267_,
		_w15268_
	);
	LUT2 #(
		.INIT('h1)
	) name14737 (
		\sa33_reg[2]/P0001 ,
		_w12468_,
		_w15269_
	);
	LUT2 #(
		.INIT('h4)
	) name14738 (
		_w13698_,
		_w15269_,
		_w15270_
	);
	LUT2 #(
		.INIT('h4)
	) name14739 (
		_w13668_,
		_w15270_,
		_w15271_
	);
	LUT2 #(
		.INIT('h1)
	) name14740 (
		_w15268_,
		_w15271_,
		_w15272_
	);
	LUT2 #(
		.INIT('h1)
	) name14741 (
		_w14011_,
		_w15043_,
		_w15273_
	);
	LUT2 #(
		.INIT('h4)
	) name14742 (
		_w15272_,
		_w15273_,
		_w15274_
	);
	LUT2 #(
		.INIT('h1)
	) name14743 (
		\sa33_reg[1]/P0001 ,
		_w15274_,
		_w15275_
	);
	LUT2 #(
		.INIT('h1)
	) name14744 (
		_w13668_,
		_w13986_,
		_w15276_
	);
	LUT2 #(
		.INIT('h1)
	) name14745 (
		\sa33_reg[4]/P0001 ,
		_w15276_,
		_w15277_
	);
	LUT2 #(
		.INIT('h1)
	) name14746 (
		_w13949_,
		_w15277_,
		_w15278_
	);
	LUT2 #(
		.INIT('h2)
	) name14747 (
		_w14021_,
		_w15278_,
		_w15279_
	);
	LUT2 #(
		.INIT('h8)
	) name14748 (
		\sa33_reg[1]/P0001 ,
		_w15033_,
		_w15280_
	);
	LUT2 #(
		.INIT('h8)
	) name14749 (
		_w13720_,
		_w14595_,
		_w15281_
	);
	LUT2 #(
		.INIT('h1)
	) name14750 (
		_w12474_,
		_w12863_,
		_w15282_
	);
	LUT2 #(
		.INIT('h1)
	) name14751 (
		_w14612_,
		_w15281_,
		_w15283_
	);
	LUT2 #(
		.INIT('h8)
	) name14752 (
		_w15282_,
		_w15283_,
		_w15284_
	);
	LUT2 #(
		.INIT('h4)
	) name14753 (
		_w15280_,
		_w15284_,
		_w15285_
	);
	LUT2 #(
		.INIT('h4)
	) name14754 (
		_w15279_,
		_w15285_,
		_w15286_
	);
	LUT2 #(
		.INIT('h4)
	) name14755 (
		_w15275_,
		_w15286_,
		_w15287_
	);
	LUT2 #(
		.INIT('h4)
	) name14756 (
		_w15266_,
		_w15287_,
		_w15288_
	);
	LUT2 #(
		.INIT('h4)
	) name14757 (
		_w15244_,
		_w15288_,
		_w15289_
	);
	LUT2 #(
		.INIT('h2)
	) name14758 (
		\u0_w_reg[0][22]/P0001 ,
		_w15289_,
		_w15290_
	);
	LUT2 #(
		.INIT('h4)
	) name14759 (
		\u0_w_reg[0][22]/P0001 ,
		_w15289_,
		_w15291_
	);
	LUT2 #(
		.INIT('h1)
	) name14760 (
		_w15290_,
		_w15291_,
		_w15292_
	);
	LUT2 #(
		.INIT('h8)
	) name14761 (
		_w13284_,
		_w15292_,
		_w15293_
	);
	LUT2 #(
		.INIT('h1)
	) name14762 (
		_w13284_,
		_w15292_,
		_w15294_
	);
	LUT2 #(
		.INIT('h1)
	) name14763 (
		_w15293_,
		_w15294_,
		_w15295_
	);
	LUT2 #(
		.INIT('h1)
	) name14764 (
		_w15221_,
		_w15295_,
		_w15296_
	);
	LUT2 #(
		.INIT('h8)
	) name14765 (
		_w15221_,
		_w15295_,
		_w15297_
	);
	LUT2 #(
		.INIT('h1)
	) name14766 (
		\ld_r_reg/P0001 ,
		_w15296_,
		_w15298_
	);
	LUT2 #(
		.INIT('h4)
	) name14767 (
		_w15297_,
		_w15298_,
		_w15299_
	);
	LUT2 #(
		.INIT('h2)
	) name14768 (
		\text_in_r_reg[118]/P0001 ,
		\u0_w_reg[0][22]/P0001 ,
		_w15300_
	);
	LUT2 #(
		.INIT('h4)
	) name14769 (
		\text_in_r_reg[118]/P0001 ,
		\u0_w_reg[0][22]/P0001 ,
		_w15301_
	);
	LUT2 #(
		.INIT('h2)
	) name14770 (
		\ld_r_reg/P0001 ,
		_w15300_,
		_w15302_
	);
	LUT2 #(
		.INIT('h4)
	) name14771 (
		_w15301_,
		_w15302_,
		_w15303_
	);
	LUT2 #(
		.INIT('h1)
	) name14772 (
		_w15299_,
		_w15303_,
		_w15304_
	);
	LUT2 #(
		.INIT('h1)
	) name14773 (
		\u0_w_reg[0][8]/P0001 ,
		_w14113_,
		_w15305_
	);
	LUT2 #(
		.INIT('h8)
	) name14774 (
		\u0_w_reg[0][8]/P0001 ,
		_w14113_,
		_w15306_
	);
	LUT2 #(
		.INIT('h1)
	) name14775 (
		_w15305_,
		_w15306_,
		_w15307_
	);
	LUT2 #(
		.INIT('h2)
	) name14776 (
		_w13922_,
		_w14033_,
		_w15308_
	);
	LUT2 #(
		.INIT('h4)
	) name14777 (
		_w13922_,
		_w14033_,
		_w15309_
	);
	LUT2 #(
		.INIT('h1)
	) name14778 (
		_w15308_,
		_w15309_,
		_w15310_
	);
	LUT2 #(
		.INIT('h2)
	) name14779 (
		_w15131_,
		_w15310_,
		_w15311_
	);
	LUT2 #(
		.INIT('h4)
	) name14780 (
		_w15131_,
		_w15310_,
		_w15312_
	);
	LUT2 #(
		.INIT('h1)
	) name14781 (
		_w15311_,
		_w15312_,
		_w15313_
	);
	LUT2 #(
		.INIT('h4)
	) name14782 (
		_w15307_,
		_w15313_,
		_w15314_
	);
	LUT2 #(
		.INIT('h2)
	) name14783 (
		_w15307_,
		_w15313_,
		_w15315_
	);
	LUT2 #(
		.INIT('h1)
	) name14784 (
		\ld_r_reg/P0001 ,
		_w15314_,
		_w15316_
	);
	LUT2 #(
		.INIT('h4)
	) name14785 (
		_w15315_,
		_w15316_,
		_w15317_
	);
	LUT2 #(
		.INIT('h2)
	) name14786 (
		\text_in_r_reg[104]/P0001 ,
		\u0_w_reg[0][8]/P0001 ,
		_w15318_
	);
	LUT2 #(
		.INIT('h4)
	) name14787 (
		\text_in_r_reg[104]/P0001 ,
		\u0_w_reg[0][8]/P0001 ,
		_w15319_
	);
	LUT2 #(
		.INIT('h2)
	) name14788 (
		\ld_r_reg/P0001 ,
		_w15318_,
		_w15320_
	);
	LUT2 #(
		.INIT('h4)
	) name14789 (
		_w15319_,
		_w15320_,
		_w15321_
	);
	LUT2 #(
		.INIT('h1)
	) name14790 (
		_w15317_,
		_w15321_,
		_w15322_
	);
	LUT2 #(
		.INIT('h2)
	) name14791 (
		_w14491_,
		_w14801_,
		_w15323_
	);
	LUT2 #(
		.INIT('h4)
	) name14792 (
		_w14491_,
		_w14801_,
		_w15324_
	);
	LUT2 #(
		.INIT('h1)
	) name14793 (
		_w15323_,
		_w15324_,
		_w15325_
	);
	LUT2 #(
		.INIT('h8)
	) name14794 (
		_w15110_,
		_w15325_,
		_w15326_
	);
	LUT2 #(
		.INIT('h1)
	) name14795 (
		_w15110_,
		_w15325_,
		_w15327_
	);
	LUT2 #(
		.INIT('h1)
	) name14796 (
		_w15326_,
		_w15327_,
		_w15328_
	);
	LUT2 #(
		.INIT('h1)
	) name14797 (
		_w14033_,
		_w14567_,
		_w15329_
	);
	LUT2 #(
		.INIT('h8)
	) name14798 (
		_w14033_,
		_w14567_,
		_w15330_
	);
	LUT2 #(
		.INIT('h1)
	) name14799 (
		_w15329_,
		_w15330_,
		_w15331_
	);
	LUT2 #(
		.INIT('h2)
	) name14800 (
		\u0_w_reg[0][3]/P0001 ,
		_w15068_,
		_w15332_
	);
	LUT2 #(
		.INIT('h4)
	) name14801 (
		\u0_w_reg[0][3]/P0001 ,
		_w15068_,
		_w15333_
	);
	LUT2 #(
		.INIT('h1)
	) name14802 (
		_w15332_,
		_w15333_,
		_w15334_
	);
	LUT2 #(
		.INIT('h8)
	) name14803 (
		_w15331_,
		_w15334_,
		_w15335_
	);
	LUT2 #(
		.INIT('h1)
	) name14804 (
		_w15331_,
		_w15334_,
		_w15336_
	);
	LUT2 #(
		.INIT('h1)
	) name14805 (
		_w15335_,
		_w15336_,
		_w15337_
	);
	LUT2 #(
		.INIT('h2)
	) name14806 (
		_w15328_,
		_w15337_,
		_w15338_
	);
	LUT2 #(
		.INIT('h4)
	) name14807 (
		_w15328_,
		_w15337_,
		_w15339_
	);
	LUT2 #(
		.INIT('h1)
	) name14808 (
		\ld_r_reg/P0001 ,
		_w15338_,
		_w15340_
	);
	LUT2 #(
		.INIT('h4)
	) name14809 (
		_w15339_,
		_w15340_,
		_w15341_
	);
	LUT2 #(
		.INIT('h2)
	) name14810 (
		\text_in_r_reg[99]/P0001 ,
		\u0_w_reg[0][3]/P0001 ,
		_w15342_
	);
	LUT2 #(
		.INIT('h4)
	) name14811 (
		\text_in_r_reg[99]/P0001 ,
		\u0_w_reg[0][3]/P0001 ,
		_w15343_
	);
	LUT2 #(
		.INIT('h2)
	) name14812 (
		\ld_r_reg/P0001 ,
		_w15342_,
		_w15344_
	);
	LUT2 #(
		.INIT('h4)
	) name14813 (
		_w15343_,
		_w15344_,
		_w15345_
	);
	LUT2 #(
		.INIT('h1)
	) name14814 (
		_w15341_,
		_w15345_,
		_w15346_
	);
	LUT2 #(
		.INIT('h2)
	) name14815 (
		\u0_w_reg[0][26]/P0001 ,
		_w15068_,
		_w15347_
	);
	LUT2 #(
		.INIT('h4)
	) name14816 (
		\u0_w_reg[0][26]/P0001 ,
		_w15068_,
		_w15348_
	);
	LUT2 #(
		.INIT('h1)
	) name14817 (
		_w15347_,
		_w15348_,
		_w15349_
	);
	LUT2 #(
		.INIT('h8)
	) name14818 (
		_w14897_,
		_w15349_,
		_w15350_
	);
	LUT2 #(
		.INIT('h1)
	) name14819 (
		_w14897_,
		_w15349_,
		_w15351_
	);
	LUT2 #(
		.INIT('h1)
	) name14820 (
		_w15350_,
		_w15351_,
		_w15352_
	);
	LUT2 #(
		.INIT('h1)
	) name14821 (
		_w14213_,
		_w15352_,
		_w15353_
	);
	LUT2 #(
		.INIT('h8)
	) name14822 (
		_w14213_,
		_w15352_,
		_w15354_
	);
	LUT2 #(
		.INIT('h1)
	) name14823 (
		\ld_r_reg/P0001 ,
		_w15353_,
		_w15355_
	);
	LUT2 #(
		.INIT('h4)
	) name14824 (
		_w15354_,
		_w15355_,
		_w15356_
	);
	LUT2 #(
		.INIT('h1)
	) name14825 (
		\text_in_r_reg[122]/P0001 ,
		\u0_w_reg[0][26]/P0001 ,
		_w15357_
	);
	LUT2 #(
		.INIT('h8)
	) name14826 (
		\text_in_r_reg[122]/P0001 ,
		\u0_w_reg[0][26]/P0001 ,
		_w15358_
	);
	LUT2 #(
		.INIT('h2)
	) name14827 (
		\ld_r_reg/P0001 ,
		_w15357_,
		_w15359_
	);
	LUT2 #(
		.INIT('h4)
	) name14828 (
		_w15358_,
		_w15359_,
		_w15360_
	);
	LUT2 #(
		.INIT('h1)
	) name14829 (
		_w15356_,
		_w15360_,
		_w15361_
	);
	LUT2 #(
		.INIT('h1)
	) name14830 (
		_w13649_,
		_w14804_,
		_w15362_
	);
	LUT2 #(
		.INIT('h8)
	) name14831 (
		_w13649_,
		_w14804_,
		_w15363_
	);
	LUT2 #(
		.INIT('h1)
	) name14832 (
		_w15362_,
		_w15363_,
		_w15364_
	);
	LUT2 #(
		.INIT('h2)
	) name14833 (
		\u0_w_reg[0][2]/P0001 ,
		_w14894_,
		_w15365_
	);
	LUT2 #(
		.INIT('h4)
	) name14834 (
		\u0_w_reg[0][2]/P0001 ,
		_w14894_,
		_w15366_
	);
	LUT2 #(
		.INIT('h1)
	) name14835 (
		_w15365_,
		_w15366_,
		_w15367_
	);
	LUT2 #(
		.INIT('h8)
	) name14836 (
		_w13752_,
		_w15367_,
		_w15368_
	);
	LUT2 #(
		.INIT('h1)
	) name14837 (
		_w13752_,
		_w15367_,
		_w15369_
	);
	LUT2 #(
		.INIT('h1)
	) name14838 (
		_w15368_,
		_w15369_,
		_w15370_
	);
	LUT2 #(
		.INIT('h1)
	) name14839 (
		_w15364_,
		_w15370_,
		_w15371_
	);
	LUT2 #(
		.INIT('h8)
	) name14840 (
		_w15364_,
		_w15370_,
		_w15372_
	);
	LUT2 #(
		.INIT('h1)
	) name14841 (
		\ld_r_reg/P0001 ,
		_w15371_,
		_w15373_
	);
	LUT2 #(
		.INIT('h4)
	) name14842 (
		_w15372_,
		_w15373_,
		_w15374_
	);
	LUT2 #(
		.INIT('h2)
	) name14843 (
		\text_in_r_reg[98]/P0001 ,
		\u0_w_reg[0][2]/P0001 ,
		_w15375_
	);
	LUT2 #(
		.INIT('h4)
	) name14844 (
		\text_in_r_reg[98]/P0001 ,
		\u0_w_reg[0][2]/P0001 ,
		_w15376_
	);
	LUT2 #(
		.INIT('h2)
	) name14845 (
		\ld_r_reg/P0001 ,
		_w15375_,
		_w15377_
	);
	LUT2 #(
		.INIT('h4)
	) name14846 (
		_w15376_,
		_w15377_,
		_w15378_
	);
	LUT2 #(
		.INIT('h1)
	) name14847 (
		_w15374_,
		_w15378_,
		_w15379_
	);
	LUT2 #(
		.INIT('h2)
	) name14848 (
		_w13183_,
		_w13284_,
		_w15380_
	);
	LUT2 #(
		.INIT('h4)
	) name14849 (
		_w13183_,
		_w13284_,
		_w15381_
	);
	LUT2 #(
		.INIT('h1)
	) name14850 (
		_w15380_,
		_w15381_,
		_w15382_
	);
	LUT2 #(
		.INIT('h2)
	) name14851 (
		\u0_w_reg[0][30]/P0001 ,
		_w15289_,
		_w15383_
	);
	LUT2 #(
		.INIT('h4)
	) name14852 (
		\u0_w_reg[0][30]/P0001 ,
		_w15289_,
		_w15384_
	);
	LUT2 #(
		.INIT('h1)
	) name14853 (
		_w15383_,
		_w15384_,
		_w15385_
	);
	LUT2 #(
		.INIT('h8)
	) name14854 (
		_w15382_,
		_w15385_,
		_w15386_
	);
	LUT2 #(
		.INIT('h1)
	) name14855 (
		_w15382_,
		_w15385_,
		_w15387_
	);
	LUT2 #(
		.INIT('h1)
	) name14856 (
		_w15386_,
		_w15387_,
		_w15388_
	);
	LUT2 #(
		.INIT('h1)
	) name14857 (
		_w12851_,
		_w15388_,
		_w15389_
	);
	LUT2 #(
		.INIT('h8)
	) name14858 (
		_w12851_,
		_w15388_,
		_w15390_
	);
	LUT2 #(
		.INIT('h1)
	) name14859 (
		\ld_r_reg/P0001 ,
		_w15389_,
		_w15391_
	);
	LUT2 #(
		.INIT('h4)
	) name14860 (
		_w15390_,
		_w15391_,
		_w15392_
	);
	LUT2 #(
		.INIT('h1)
	) name14861 (
		\text_in_r_reg[126]/P0001 ,
		\u0_w_reg[0][30]/P0001 ,
		_w15393_
	);
	LUT2 #(
		.INIT('h8)
	) name14862 (
		\text_in_r_reg[126]/P0001 ,
		\u0_w_reg[0][30]/P0001 ,
		_w15394_
	);
	LUT2 #(
		.INIT('h2)
	) name14863 (
		\ld_r_reg/P0001 ,
		_w15393_,
		_w15395_
	);
	LUT2 #(
		.INIT('h4)
	) name14864 (
		_w15394_,
		_w15395_,
		_w15396_
	);
	LUT2 #(
		.INIT('h1)
	) name14865 (
		_w15392_,
		_w15396_,
		_w15397_
	);
	LUT2 #(
		.INIT('h2)
	) name14866 (
		\u0_w_reg[0][31]/P0001 ,
		_w13558_,
		_w15398_
	);
	LUT2 #(
		.INIT('h4)
	) name14867 (
		\u0_w_reg[0][31]/P0001 ,
		_w13558_,
		_w15399_
	);
	LUT2 #(
		.INIT('h1)
	) name14868 (
		_w15398_,
		_w15399_,
		_w15400_
	);
	LUT2 #(
		.INIT('h8)
	) name14869 (
		_w13186_,
		_w15310_,
		_w15401_
	);
	LUT2 #(
		.INIT('h1)
	) name14870 (
		_w13186_,
		_w15310_,
		_w15402_
	);
	LUT2 #(
		.INIT('h1)
	) name14871 (
		_w15401_,
		_w15402_,
		_w15403_
	);
	LUT2 #(
		.INIT('h4)
	) name14872 (
		_w15400_,
		_w15403_,
		_w15404_
	);
	LUT2 #(
		.INIT('h2)
	) name14873 (
		_w15400_,
		_w15403_,
		_w15405_
	);
	LUT2 #(
		.INIT('h1)
	) name14874 (
		\ld_r_reg/P0001 ,
		_w15404_,
		_w15406_
	);
	LUT2 #(
		.INIT('h4)
	) name14875 (
		_w15405_,
		_w15406_,
		_w15407_
	);
	LUT2 #(
		.INIT('h2)
	) name14876 (
		\text_in_r_reg[127]/P0001 ,
		\u0_w_reg[0][31]/P0001 ,
		_w15408_
	);
	LUT2 #(
		.INIT('h4)
	) name14877 (
		\text_in_r_reg[127]/P0001 ,
		\u0_w_reg[0][31]/P0001 ,
		_w15409_
	);
	LUT2 #(
		.INIT('h2)
	) name14878 (
		\ld_r_reg/P0001 ,
		_w15408_,
		_w15410_
	);
	LUT2 #(
		.INIT('h4)
	) name14879 (
		_w15409_,
		_w15410_,
		_w15411_
	);
	LUT2 #(
		.INIT('h1)
	) name14880 (
		_w15407_,
		_w15411_,
		_w15412_
	);
	LUT2 #(
		.INIT('h1)
	) name14881 (
		_w13835_,
		_w14801_,
		_w15413_
	);
	LUT2 #(
		.INIT('h8)
	) name14882 (
		_w13835_,
		_w14801_,
		_w15414_
	);
	LUT2 #(
		.INIT('h1)
	) name14883 (
		_w15413_,
		_w15414_,
		_w15415_
	);
	LUT2 #(
		.INIT('h1)
	) name14884 (
		_w14210_,
		_w15415_,
		_w15416_
	);
	LUT2 #(
		.INIT('h8)
	) name14885 (
		_w14210_,
		_w15415_,
		_w15417_
	);
	LUT2 #(
		.INIT('h1)
	) name14886 (
		_w15416_,
		_w15417_,
		_w15418_
	);
	LUT2 #(
		.INIT('h2)
	) name14887 (
		\u0_w_reg[0][18]/P0001 ,
		_w15068_,
		_w15419_
	);
	LUT2 #(
		.INIT('h4)
	) name14888 (
		\u0_w_reg[0][18]/P0001 ,
		_w15068_,
		_w15420_
	);
	LUT2 #(
		.INIT('h1)
	) name14889 (
		_w15419_,
		_w15420_,
		_w15421_
	);
	LUT2 #(
		.INIT('h8)
	) name14890 (
		_w14894_,
		_w15421_,
		_w15422_
	);
	LUT2 #(
		.INIT('h1)
	) name14891 (
		_w14894_,
		_w15421_,
		_w15423_
	);
	LUT2 #(
		.INIT('h1)
	) name14892 (
		_w15422_,
		_w15423_,
		_w15424_
	);
	LUT2 #(
		.INIT('h4)
	) name14893 (
		_w15418_,
		_w15424_,
		_w15425_
	);
	LUT2 #(
		.INIT('h2)
	) name14894 (
		_w15418_,
		_w15424_,
		_w15426_
	);
	LUT2 #(
		.INIT('h1)
	) name14895 (
		\ld_r_reg/P0001 ,
		_w15425_,
		_w15427_
	);
	LUT2 #(
		.INIT('h4)
	) name14896 (
		_w15426_,
		_w15427_,
		_w15428_
	);
	LUT2 #(
		.INIT('h2)
	) name14897 (
		\text_in_r_reg[114]/P0001 ,
		\u0_w_reg[0][18]/P0001 ,
		_w15429_
	);
	LUT2 #(
		.INIT('h4)
	) name14898 (
		\text_in_r_reg[114]/P0001 ,
		\u0_w_reg[0][18]/P0001 ,
		_w15430_
	);
	LUT2 #(
		.INIT('h2)
	) name14899 (
		\ld_r_reg/P0001 ,
		_w15429_,
		_w15431_
	);
	LUT2 #(
		.INIT('h4)
	) name14900 (
		_w15430_,
		_w15431_,
		_w15432_
	);
	LUT2 #(
		.INIT('h1)
	) name14901 (
		_w15428_,
		_w15432_,
		_w15433_
	);
	LUT2 #(
		.INIT('h1)
	) name14902 (
		_w14400_,
		_w15382_,
		_w15434_
	);
	LUT2 #(
		.INIT('h8)
	) name14903 (
		_w14400_,
		_w15382_,
		_w15435_
	);
	LUT2 #(
		.INIT('h1)
	) name14904 (
		_w15434_,
		_w15435_,
		_w15436_
	);
	LUT2 #(
		.INIT('h1)
	) name14905 (
		\u0_w_reg[0][23]/P0001 ,
		_w15310_,
		_w15437_
	);
	LUT2 #(
		.INIT('h8)
	) name14906 (
		\u0_w_reg[0][23]/P0001 ,
		_w15310_,
		_w15438_
	);
	LUT2 #(
		.INIT('h1)
	) name14907 (
		_w15437_,
		_w15438_,
		_w15439_
	);
	LUT2 #(
		.INIT('h1)
	) name14908 (
		_w15436_,
		_w15439_,
		_w15440_
	);
	LUT2 #(
		.INIT('h8)
	) name14909 (
		_w15436_,
		_w15439_,
		_w15441_
	);
	LUT2 #(
		.INIT('h1)
	) name14910 (
		\ld_r_reg/P0001 ,
		_w15440_,
		_w15442_
	);
	LUT2 #(
		.INIT('h4)
	) name14911 (
		_w15441_,
		_w15442_,
		_w15443_
	);
	LUT2 #(
		.INIT('h2)
	) name14912 (
		\text_in_r_reg[119]/P0001 ,
		\u0_w_reg[0][23]/P0001 ,
		_w15444_
	);
	LUT2 #(
		.INIT('h4)
	) name14913 (
		\text_in_r_reg[119]/P0001 ,
		\u0_w_reg[0][23]/P0001 ,
		_w15445_
	);
	LUT2 #(
		.INIT('h2)
	) name14914 (
		\ld_r_reg/P0001 ,
		_w15444_,
		_w15446_
	);
	LUT2 #(
		.INIT('h4)
	) name14915 (
		_w15445_,
		_w15446_,
		_w15447_
	);
	LUT2 #(
		.INIT('h1)
	) name14916 (
		_w15443_,
		_w15447_,
		_w15448_
	);
	LUT2 #(
		.INIT('h1)
	) name14917 (
		_w12405_,
		_w13186_,
		_w15449_
	);
	LUT2 #(
		.INIT('h8)
	) name14918 (
		_w12405_,
		_w13186_,
		_w15450_
	);
	LUT2 #(
		.INIT('h1)
	) name14919 (
		_w15449_,
		_w15450_,
		_w15451_
	);
	LUT2 #(
		.INIT('h2)
	) name14920 (
		\u0_w_reg[0][14]/P0001 ,
		_w15289_,
		_w15452_
	);
	LUT2 #(
		.INIT('h4)
	) name14921 (
		\u0_w_reg[0][14]/P0001 ,
		_w15289_,
		_w15453_
	);
	LUT2 #(
		.INIT('h1)
	) name14922 (
		_w15452_,
		_w15453_,
		_w15454_
	);
	LUT2 #(
		.INIT('h8)
	) name14923 (
		_w12580_,
		_w15454_,
		_w15455_
	);
	LUT2 #(
		.INIT('h1)
	) name14924 (
		_w12580_,
		_w15454_,
		_w15456_
	);
	LUT2 #(
		.INIT('h1)
	) name14925 (
		_w15455_,
		_w15456_,
		_w15457_
	);
	LUT2 #(
		.INIT('h1)
	) name14926 (
		_w15451_,
		_w15457_,
		_w15458_
	);
	LUT2 #(
		.INIT('h8)
	) name14927 (
		_w15451_,
		_w15457_,
		_w15459_
	);
	LUT2 #(
		.INIT('h1)
	) name14928 (
		\ld_r_reg/P0001 ,
		_w15458_,
		_w15460_
	);
	LUT2 #(
		.INIT('h4)
	) name14929 (
		_w15459_,
		_w15460_,
		_w15461_
	);
	LUT2 #(
		.INIT('h2)
	) name14930 (
		\text_in_r_reg[110]/P0001 ,
		\u0_w_reg[0][14]/P0001 ,
		_w15462_
	);
	LUT2 #(
		.INIT('h4)
	) name14931 (
		\text_in_r_reg[110]/P0001 ,
		\u0_w_reg[0][14]/P0001 ,
		_w15463_
	);
	LUT2 #(
		.INIT('h2)
	) name14932 (
		\ld_r_reg/P0001 ,
		_w15462_,
		_w15464_
	);
	LUT2 #(
		.INIT('h4)
	) name14933 (
		_w15463_,
		_w15464_,
		_w15465_
	);
	LUT2 #(
		.INIT('h1)
	) name14934 (
		_w15461_,
		_w15465_,
		_w15466_
	);
	LUT2 #(
		.INIT('h1)
	) name14935 (
		_w13284_,
		_w14660_,
		_w15467_
	);
	LUT2 #(
		.INIT('h8)
	) name14936 (
		_w13284_,
		_w14660_,
		_w15468_
	);
	LUT2 #(
		.INIT('h1)
	) name14937 (
		_w15467_,
		_w15468_,
		_w15469_
	);
	LUT2 #(
		.INIT('h2)
	) name14938 (
		\u0_w_reg[0][15]/P0001 ,
		_w14033_,
		_w15470_
	);
	LUT2 #(
		.INIT('h4)
	) name14939 (
		\u0_w_reg[0][15]/P0001 ,
		_w14033_,
		_w15471_
	);
	LUT2 #(
		.INIT('h1)
	) name14940 (
		_w15470_,
		_w15471_,
		_w15472_
	);
	LUT2 #(
		.INIT('h8)
	) name14941 (
		_w15289_,
		_w15472_,
		_w15473_
	);
	LUT2 #(
		.INIT('h1)
	) name14942 (
		_w15289_,
		_w15472_,
		_w15474_
	);
	LUT2 #(
		.INIT('h1)
	) name14943 (
		_w15473_,
		_w15474_,
		_w15475_
	);
	LUT2 #(
		.INIT('h1)
	) name14944 (
		_w15469_,
		_w15475_,
		_w15476_
	);
	LUT2 #(
		.INIT('h8)
	) name14945 (
		_w15469_,
		_w15475_,
		_w15477_
	);
	LUT2 #(
		.INIT('h1)
	) name14946 (
		\ld_r_reg/P0001 ,
		_w15476_,
		_w15478_
	);
	LUT2 #(
		.INIT('h4)
	) name14947 (
		_w15477_,
		_w15478_,
		_w15479_
	);
	LUT2 #(
		.INIT('h2)
	) name14948 (
		\text_in_r_reg[111]/P0001 ,
		\u0_w_reg[0][15]/P0001 ,
		_w15480_
	);
	LUT2 #(
		.INIT('h4)
	) name14949 (
		\text_in_r_reg[111]/P0001 ,
		\u0_w_reg[0][15]/P0001 ,
		_w15481_
	);
	LUT2 #(
		.INIT('h2)
	) name14950 (
		\ld_r_reg/P0001 ,
		_w15480_,
		_w15482_
	);
	LUT2 #(
		.INIT('h4)
	) name14951 (
		_w15481_,
		_w15482_,
		_w15483_
	);
	LUT2 #(
		.INIT('h1)
	) name14952 (
		_w15479_,
		_w15483_,
		_w15484_
	);
	LUT2 #(
		.INIT('h1)
	) name14953 (
		_w13091_,
		_w14660_,
		_w15485_
	);
	LUT2 #(
		.INIT('h8)
	) name14954 (
		_w13091_,
		_w14660_,
		_w15486_
	);
	LUT2 #(
		.INIT('h1)
	) name14955 (
		_w15485_,
		_w15486_,
		_w15487_
	);
	LUT2 #(
		.INIT('h2)
	) name14956 (
		\u0_w_reg[0][7]/P0001 ,
		_w15289_,
		_w15488_
	);
	LUT2 #(
		.INIT('h4)
	) name14957 (
		\u0_w_reg[0][7]/P0001 ,
		_w15289_,
		_w15489_
	);
	LUT2 #(
		.INIT('h1)
	) name14958 (
		_w15488_,
		_w15489_,
		_w15490_
	);
	LUT2 #(
		.INIT('h8)
	) name14959 (
		_w13922_,
		_w15490_,
		_w15491_
	);
	LUT2 #(
		.INIT('h1)
	) name14960 (
		_w13922_,
		_w15490_,
		_w15492_
	);
	LUT2 #(
		.INIT('h1)
	) name14961 (
		_w15491_,
		_w15492_,
		_w15493_
	);
	LUT2 #(
		.INIT('h1)
	) name14962 (
		_w15487_,
		_w15493_,
		_w15494_
	);
	LUT2 #(
		.INIT('h8)
	) name14963 (
		_w15487_,
		_w15493_,
		_w15495_
	);
	LUT2 #(
		.INIT('h1)
	) name14964 (
		\ld_r_reg/P0001 ,
		_w15494_,
		_w15496_
	);
	LUT2 #(
		.INIT('h4)
	) name14965 (
		_w15495_,
		_w15496_,
		_w15497_
	);
	LUT2 #(
		.INIT('h2)
	) name14966 (
		\text_in_r_reg[103]/P0001 ,
		\u0_w_reg[0][7]/P0001 ,
		_w15498_
	);
	LUT2 #(
		.INIT('h4)
	) name14967 (
		\text_in_r_reg[103]/P0001 ,
		\u0_w_reg[0][7]/P0001 ,
		_w15499_
	);
	LUT2 #(
		.INIT('h2)
	) name14968 (
		\ld_r_reg/P0001 ,
		_w15498_,
		_w15500_
	);
	LUT2 #(
		.INIT('h4)
	) name14969 (
		_w15499_,
		_w15500_,
		_w15501_
	);
	LUT2 #(
		.INIT('h1)
	) name14970 (
		_w15497_,
		_w15501_,
		_w15502_
	);
	LUT2 #(
		.INIT('h2)
	) name14971 (
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w15503_
	);
	LUT2 #(
		.INIT('h2)
	) name14972 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w15504_
	);
	LUT2 #(
		.INIT('h8)
	) name14973 (
		\u0_w_reg[3][21]/P0001 ,
		_w15504_,
		_w15505_
	);
	LUT2 #(
		.INIT('h1)
	) name14974 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w15506_
	);
	LUT2 #(
		.INIT('h8)
	) name14975 (
		\u0_w_reg[3][18]/P0001 ,
		_w15506_,
		_w15507_
	);
	LUT2 #(
		.INIT('h4)
	) name14976 (
		\u0_w_reg[3][21]/P0001 ,
		_w15507_,
		_w15508_
	);
	LUT2 #(
		.INIT('h1)
	) name14977 (
		_w15505_,
		_w15508_,
		_w15509_
	);
	LUT2 #(
		.INIT('h2)
	) name14978 (
		_w15503_,
		_w15509_,
		_w15510_
	);
	LUT2 #(
		.INIT('h2)
	) name14979 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w15511_
	);
	LUT2 #(
		.INIT('h8)
	) name14980 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w15512_
	);
	LUT2 #(
		.INIT('h8)
	) name14981 (
		\u0_w_reg[3][20]/P0001 ,
		_w15512_,
		_w15513_
	);
	LUT2 #(
		.INIT('h8)
	) name14982 (
		\u0_w_reg[3][23]/P0001 ,
		_w15513_,
		_w15514_
	);
	LUT2 #(
		.INIT('h8)
	) name14983 (
		_w15511_,
		_w15514_,
		_w15515_
	);
	LUT2 #(
		.INIT('h8)
	) name14984 (
		\u0_w_reg[3][21]/P0001 ,
		_w15503_,
		_w15516_
	);
	LUT2 #(
		.INIT('h4)
	) name14985 (
		_w15511_,
		_w15516_,
		_w15517_
	);
	LUT2 #(
		.INIT('h4)
	) name14986 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w15518_
	);
	LUT2 #(
		.INIT('h4)
	) name14987 (
		\u0_w_reg[3][20]/P0001 ,
		_w15518_,
		_w15519_
	);
	LUT2 #(
		.INIT('h1)
	) name14988 (
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w15520_
	);
	LUT2 #(
		.INIT('h8)
	) name14989 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w15521_
	);
	LUT2 #(
		.INIT('h8)
	) name14990 (
		_w15520_,
		_w15521_,
		_w15522_
	);
	LUT2 #(
		.INIT('h1)
	) name14991 (
		_w15519_,
		_w15522_,
		_w15523_
	);
	LUT2 #(
		.INIT('h2)
	) name14992 (
		\u0_w_reg[3][18]/P0001 ,
		_w15523_,
		_w15524_
	);
	LUT2 #(
		.INIT('h4)
	) name14993 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w15525_
	);
	LUT2 #(
		.INIT('h8)
	) name14994 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w15526_
	);
	LUT2 #(
		.INIT('h8)
	) name14995 (
		_w15525_,
		_w15526_,
		_w15527_
	);
	LUT2 #(
		.INIT('h8)
	) name14996 (
		\u0_w_reg[3][22]/P0001 ,
		_w15527_,
		_w15528_
	);
	LUT2 #(
		.INIT('h4)
	) name14997 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w15529_
	);
	LUT2 #(
		.INIT('h4)
	) name14998 (
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w15530_
	);
	LUT2 #(
		.INIT('h4)
	) name14999 (
		\u0_w_reg[3][21]/P0001 ,
		_w15530_,
		_w15531_
	);
	LUT2 #(
		.INIT('h8)
	) name15000 (
		_w15529_,
		_w15531_,
		_w15532_
	);
	LUT2 #(
		.INIT('h1)
	) name15001 (
		_w15517_,
		_w15528_,
		_w15533_
	);
	LUT2 #(
		.INIT('h4)
	) name15002 (
		_w15532_,
		_w15533_,
		_w15534_
	);
	LUT2 #(
		.INIT('h4)
	) name15003 (
		_w15524_,
		_w15534_,
		_w15535_
	);
	LUT2 #(
		.INIT('h1)
	) name15004 (
		\u0_w_reg[3][17]/P0001 ,
		_w15535_,
		_w15536_
	);
	LUT2 #(
		.INIT('h2)
	) name15005 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w15537_
	);
	LUT2 #(
		.INIT('h8)
	) name15006 (
		_w15512_,
		_w15537_,
		_w15538_
	);
	LUT2 #(
		.INIT('h4)
	) name15007 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w15539_
	);
	LUT2 #(
		.INIT('h8)
	) name15008 (
		_w15537_,
		_w15539_,
		_w15540_
	);
	LUT2 #(
		.INIT('h1)
	) name15009 (
		_w15538_,
		_w15540_,
		_w15541_
	);
	LUT2 #(
		.INIT('h2)
	) name15010 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w15542_
	);
	LUT2 #(
		.INIT('h4)
	) name15011 (
		\u0_w_reg[3][20]/P0001 ,
		_w15542_,
		_w15543_
	);
	LUT2 #(
		.INIT('h8)
	) name15012 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w15544_
	);
	LUT2 #(
		.INIT('h8)
	) name15013 (
		_w15518_,
		_w15544_,
		_w15545_
	);
	LUT2 #(
		.INIT('h1)
	) name15014 (
		_w15543_,
		_w15545_,
		_w15546_
	);
	LUT2 #(
		.INIT('h8)
	) name15015 (
		_w15541_,
		_w15546_,
		_w15547_
	);
	LUT2 #(
		.INIT('h1)
	) name15016 (
		\u0_w_reg[3][18]/P0001 ,
		_w15547_,
		_w15548_
	);
	LUT2 #(
		.INIT('h1)
	) name15017 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w15549_
	);
	LUT2 #(
		.INIT('h4)
	) name15018 (
		\u0_w_reg[3][20]/P0001 ,
		_w15549_,
		_w15550_
	);
	LUT2 #(
		.INIT('h2)
	) name15019 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w15551_
	);
	LUT2 #(
		.INIT('h4)
	) name15020 (
		\u0_w_reg[3][21]/P0001 ,
		_w15551_,
		_w15552_
	);
	LUT2 #(
		.INIT('h1)
	) name15021 (
		_w15505_,
		_w15550_,
		_w15553_
	);
	LUT2 #(
		.INIT('h4)
	) name15022 (
		_w15552_,
		_w15553_,
		_w15554_
	);
	LUT2 #(
		.INIT('h1)
	) name15023 (
		\u0_w_reg[3][18]/P0001 ,
		_w15554_,
		_w15555_
	);
	LUT2 #(
		.INIT('h8)
	) name15024 (
		_w15504_,
		_w15530_,
		_w15556_
	);
	LUT2 #(
		.INIT('h4)
	) name15025 (
		\u0_w_reg[3][21]/P0001 ,
		_w15520_,
		_w15557_
	);
	LUT2 #(
		.INIT('h8)
	) name15026 (
		_w15525_,
		_w15557_,
		_w15558_
	);
	LUT2 #(
		.INIT('h2)
	) name15027 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w15559_
	);
	LUT2 #(
		.INIT('h4)
	) name15028 (
		\u0_w_reg[3][19]/P0001 ,
		_w15559_,
		_w15560_
	);
	LUT2 #(
		.INIT('h8)
	) name15029 (
		_w15544_,
		_w15560_,
		_w15561_
	);
	LUT2 #(
		.INIT('h4)
	) name15030 (
		\u0_w_reg[3][22]/P0001 ,
		_w15521_,
		_w15562_
	);
	LUT2 #(
		.INIT('h8)
	) name15031 (
		_w15542_,
		_w15562_,
		_w15563_
	);
	LUT2 #(
		.INIT('h1)
	) name15032 (
		_w15556_,
		_w15558_,
		_w15564_
	);
	LUT2 #(
		.INIT('h1)
	) name15033 (
		_w15561_,
		_w15563_,
		_w15565_
	);
	LUT2 #(
		.INIT('h8)
	) name15034 (
		_w15564_,
		_w15565_,
		_w15566_
	);
	LUT2 #(
		.INIT('h4)
	) name15035 (
		_w15555_,
		_w15566_,
		_w15567_
	);
	LUT2 #(
		.INIT('h2)
	) name15036 (
		\u0_w_reg[3][17]/P0001 ,
		_w15567_,
		_w15568_
	);
	LUT2 #(
		.INIT('h1)
	) name15037 (
		_w15510_,
		_w15515_,
		_w15569_
	);
	LUT2 #(
		.INIT('h4)
	) name15038 (
		_w15548_,
		_w15569_,
		_w15570_
	);
	LUT2 #(
		.INIT('h4)
	) name15039 (
		_w15536_,
		_w15570_,
		_w15571_
	);
	LUT2 #(
		.INIT('h4)
	) name15040 (
		_w15568_,
		_w15571_,
		_w15572_
	);
	LUT2 #(
		.INIT('h2)
	) name15041 (
		\u0_w_reg[3][16]/P0001 ,
		_w15572_,
		_w15573_
	);
	LUT2 #(
		.INIT('h8)
	) name15042 (
		_w15503_,
		_w15506_,
		_w15574_
	);
	LUT2 #(
		.INIT('h8)
	) name15043 (
		\u0_w_reg[3][19]/P0001 ,
		_w15530_,
		_w15575_
	);
	LUT2 #(
		.INIT('h8)
	) name15044 (
		_w15525_,
		_w15559_,
		_w15576_
	);
	LUT2 #(
		.INIT('h1)
	) name15045 (
		_w15574_,
		_w15575_,
		_w15577_
	);
	LUT2 #(
		.INIT('h4)
	) name15046 (
		_w15576_,
		_w15577_,
		_w15578_
	);
	LUT2 #(
		.INIT('h1)
	) name15047 (
		\u0_w_reg[3][18]/P0001 ,
		_w15578_,
		_w15579_
	);
	LUT2 #(
		.INIT('h8)
	) name15048 (
		_w15506_,
		_w15512_,
		_w15580_
	);
	LUT2 #(
		.INIT('h4)
	) name15049 (
		\u0_w_reg[3][23]/P0001 ,
		_w15580_,
		_w15581_
	);
	LUT2 #(
		.INIT('h4)
	) name15050 (
		\u0_w_reg[3][20]/P0001 ,
		_w15526_,
		_w15582_
	);
	LUT2 #(
		.INIT('h4)
	) name15051 (
		\u0_w_reg[3][22]/P0001 ,
		_w15582_,
		_w15583_
	);
	LUT2 #(
		.INIT('h8)
	) name15052 (
		_w15537_,
		_w15549_,
		_w15584_
	);
	LUT2 #(
		.INIT('h8)
	) name15053 (
		_w15512_,
		_w15551_,
		_w15585_
	);
	LUT2 #(
		.INIT('h8)
	) name15054 (
		\u0_w_reg[3][18]/P0001 ,
		_w15585_,
		_w15586_
	);
	LUT2 #(
		.INIT('h8)
	) name15055 (
		\u0_w_reg[3][19]/P0001 ,
		_w15526_,
		_w15587_
	);
	LUT2 #(
		.INIT('h1)
	) name15056 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w15588_
	);
	LUT2 #(
		.INIT('h2)
	) name15057 (
		_w15587_,
		_w15588_,
		_w15589_
	);
	LUT2 #(
		.INIT('h8)
	) name15058 (
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w15590_
	);
	LUT2 #(
		.INIT('h4)
	) name15059 (
		\u0_w_reg[3][21]/P0001 ,
		_w15590_,
		_w15591_
	);
	LUT2 #(
		.INIT('h4)
	) name15060 (
		\u0_w_reg[3][19]/P0001 ,
		_w15591_,
		_w15592_
	);
	LUT2 #(
		.INIT('h1)
	) name15061 (
		_w15581_,
		_w15584_,
		_w15593_
	);
	LUT2 #(
		.INIT('h1)
	) name15062 (
		_w15583_,
		_w15586_,
		_w15594_
	);
	LUT2 #(
		.INIT('h1)
	) name15063 (
		_w15589_,
		_w15592_,
		_w15595_
	);
	LUT2 #(
		.INIT('h8)
	) name15064 (
		_w15594_,
		_w15595_,
		_w15596_
	);
	LUT2 #(
		.INIT('h8)
	) name15065 (
		_w15593_,
		_w15596_,
		_w15597_
	);
	LUT2 #(
		.INIT('h4)
	) name15066 (
		_w15579_,
		_w15597_,
		_w15598_
	);
	LUT2 #(
		.INIT('h2)
	) name15067 (
		\u0_w_reg[3][17]/P0001 ,
		_w15598_,
		_w15599_
	);
	LUT2 #(
		.INIT('h8)
	) name15068 (
		\u0_w_reg[3][18]/P0001 ,
		_w15557_,
		_w15600_
	);
	LUT2 #(
		.INIT('h4)
	) name15069 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w15601_
	);
	LUT2 #(
		.INIT('h8)
	) name15070 (
		\u0_w_reg[3][20]/P0001 ,
		_w15601_,
		_w15602_
	);
	LUT2 #(
		.INIT('h4)
	) name15071 (
		\u0_w_reg[3][22]/P0001 ,
		_w15602_,
		_w15603_
	);
	LUT2 #(
		.INIT('h1)
	) name15072 (
		_w15600_,
		_w15603_,
		_w15604_
	);
	LUT2 #(
		.INIT('h1)
	) name15073 (
		\u0_w_reg[3][19]/P0001 ,
		_w15604_,
		_w15605_
	);
	LUT2 #(
		.INIT('h8)
	) name15074 (
		\u0_w_reg[3][21]/P0001 ,
		_w15590_,
		_w15606_
	);
	LUT2 #(
		.INIT('h8)
	) name15075 (
		_w15506_,
		_w15606_,
		_w15607_
	);
	LUT2 #(
		.INIT('h8)
	) name15076 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w15608_
	);
	LUT2 #(
		.INIT('h8)
	) name15077 (
		_w15550_,
		_w15608_,
		_w15609_
	);
	LUT2 #(
		.INIT('h1)
	) name15078 (
		_w15607_,
		_w15609_,
		_w15610_
	);
	LUT2 #(
		.INIT('h4)
	) name15079 (
		_w15605_,
		_w15610_,
		_w15611_
	);
	LUT2 #(
		.INIT('h1)
	) name15080 (
		\u0_w_reg[3][17]/P0001 ,
		_w15611_,
		_w15612_
	);
	LUT2 #(
		.INIT('h1)
	) name15081 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w15613_
	);
	LUT2 #(
		.INIT('h4)
	) name15082 (
		\u0_w_reg[3][21]/P0001 ,
		_w15613_,
		_w15614_
	);
	LUT2 #(
		.INIT('h8)
	) name15083 (
		\u0_w_reg[3][20]/P0001 ,
		_w15526_,
		_w15615_
	);
	LUT2 #(
		.INIT('h1)
	) name15084 (
		_w15614_,
		_w15615_,
		_w15616_
	);
	LUT2 #(
		.INIT('h2)
	) name15085 (
		\u0_w_reg[3][19]/P0001 ,
		_w15616_,
		_w15617_
	);
	LUT2 #(
		.INIT('h8)
	) name15086 (
		_w15518_,
		_w15551_,
		_w15618_
	);
	LUT2 #(
		.INIT('h4)
	) name15087 (
		\u0_w_reg[3][19]/P0001 ,
		_w15618_,
		_w15619_
	);
	LUT2 #(
		.INIT('h4)
	) name15088 (
		\u0_w_reg[3][20]/P0001 ,
		_w15520_,
		_w15620_
	);
	LUT2 #(
		.INIT('h1)
	) name15089 (
		_w15619_,
		_w15620_,
		_w15621_
	);
	LUT2 #(
		.INIT('h4)
	) name15090 (
		_w15617_,
		_w15621_,
		_w15622_
	);
	LUT2 #(
		.INIT('h2)
	) name15091 (
		\u0_w_reg[3][18]/P0001 ,
		_w15622_,
		_w15623_
	);
	LUT2 #(
		.INIT('h8)
	) name15092 (
		\u0_w_reg[3][19]/P0001 ,
		_w15552_,
		_w15624_
	);
	LUT2 #(
		.INIT('h8)
	) name15093 (
		_w15539_,
		_w15601_,
		_w15625_
	);
	LUT2 #(
		.INIT('h1)
	) name15094 (
		_w15624_,
		_w15625_,
		_w15626_
	);
	LUT2 #(
		.INIT('h1)
	) name15095 (
		\u0_w_reg[3][18]/P0001 ,
		_w15626_,
		_w15627_
	);
	LUT2 #(
		.INIT('h8)
	) name15096 (
		_w15544_,
		_w15559_,
		_w15628_
	);
	LUT2 #(
		.INIT('h4)
	) name15097 (
		\u0_w_reg[3][18]/P0001 ,
		_w15628_,
		_w15629_
	);
	LUT2 #(
		.INIT('h8)
	) name15098 (
		_w15549_,
		_w15613_,
		_w15630_
	);
	LUT2 #(
		.INIT('h1)
	) name15099 (
		_w15629_,
		_w15630_,
		_w15631_
	);
	LUT2 #(
		.INIT('h4)
	) name15100 (
		_w15627_,
		_w15631_,
		_w15632_
	);
	LUT2 #(
		.INIT('h4)
	) name15101 (
		_w15623_,
		_w15632_,
		_w15633_
	);
	LUT2 #(
		.INIT('h4)
	) name15102 (
		_w15612_,
		_w15633_,
		_w15634_
	);
	LUT2 #(
		.INIT('h4)
	) name15103 (
		_w15599_,
		_w15634_,
		_w15635_
	);
	LUT2 #(
		.INIT('h1)
	) name15104 (
		\u0_w_reg[3][16]/P0001 ,
		_w15635_,
		_w15636_
	);
	LUT2 #(
		.INIT('h8)
	) name15105 (
		_w15506_,
		_w15520_,
		_w15637_
	);
	LUT2 #(
		.INIT('h4)
	) name15106 (
		\u0_w_reg[3][21]/P0001 ,
		_w15503_,
		_w15638_
	);
	LUT2 #(
		.INIT('h1)
	) name15107 (
		_w15531_,
		_w15638_,
		_w15639_
	);
	LUT2 #(
		.INIT('h2)
	) name15108 (
		_w15525_,
		_w15639_,
		_w15640_
	);
	LUT2 #(
		.INIT('h8)
	) name15109 (
		_w15521_,
		_w15559_,
		_w15641_
	);
	LUT2 #(
		.INIT('h1)
	) name15110 (
		_w15528_,
		_w15641_,
		_w15642_
	);
	LUT2 #(
		.INIT('h4)
	) name15111 (
		_w15640_,
		_w15642_,
		_w15643_
	);
	LUT2 #(
		.INIT('h2)
	) name15112 (
		\u0_w_reg[3][18]/P0001 ,
		_w15643_,
		_w15644_
	);
	LUT2 #(
		.INIT('h1)
	) name15113 (
		_w15637_,
		_w15644_,
		_w15645_
	);
	LUT2 #(
		.INIT('h1)
	) name15114 (
		\u0_w_reg[3][17]/P0001 ,
		_w15645_,
		_w15646_
	);
	LUT2 #(
		.INIT('h4)
	) name15115 (
		\u0_w_reg[3][18]/P0001 ,
		_w15545_,
		_w15647_
	);
	LUT2 #(
		.INIT('h1)
	) name15116 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w15648_
	);
	LUT2 #(
		.INIT('h8)
	) name15117 (
		_w15582_,
		_w15648_,
		_w15649_
	);
	LUT2 #(
		.INIT('h8)
	) name15118 (
		_w15513_,
		_w15537_,
		_w15650_
	);
	LUT2 #(
		.INIT('h4)
	) name15119 (
		\u0_w_reg[3][18]/P0001 ,
		_w15650_,
		_w15651_
	);
	LUT2 #(
		.INIT('h1)
	) name15120 (
		_w15647_,
		_w15649_,
		_w15652_
	);
	LUT2 #(
		.INIT('h4)
	) name15121 (
		_w15651_,
		_w15652_,
		_w15653_
	);
	LUT2 #(
		.INIT('h1)
	) name15122 (
		\u0_w_reg[3][17]/P0001 ,
		_w15653_,
		_w15654_
	);
	LUT2 #(
		.INIT('h8)
	) name15123 (
		_w15551_,
		_w15559_,
		_w15655_
	);
	LUT2 #(
		.INIT('h8)
	) name15124 (
		_w15608_,
		_w15655_,
		_w15656_
	);
	LUT2 #(
		.INIT('h8)
	) name15125 (
		_w15504_,
		_w15559_,
		_w15657_
	);
	LUT2 #(
		.INIT('h4)
	) name15126 (
		\u0_w_reg[3][23]/P0001 ,
		_w15657_,
		_w15658_
	);
	LUT2 #(
		.INIT('h4)
	) name15127 (
		\u0_w_reg[3][18]/P0001 ,
		_w15658_,
		_w15659_
	);
	LUT2 #(
		.INIT('h4)
	) name15128 (
		\u0_w_reg[3][21]/P0001 ,
		_w15648_,
		_w15660_
	);
	LUT2 #(
		.INIT('h8)
	) name15129 (
		_w15590_,
		_w15660_,
		_w15661_
	);
	LUT2 #(
		.INIT('h4)
	) name15130 (
		\u0_w_reg[3][21]/P0001 ,
		_w15504_,
		_w15662_
	);
	LUT2 #(
		.INIT('h8)
	) name15131 (
		_w15520_,
		_w15662_,
		_w15663_
	);
	LUT2 #(
		.INIT('h8)
	) name15132 (
		_w15511_,
		_w15585_,
		_w15664_
	);
	LUT2 #(
		.INIT('h1)
	) name15133 (
		_w15629_,
		_w15663_,
		_w15665_
	);
	LUT2 #(
		.INIT('h4)
	) name15134 (
		_w15664_,
		_w15665_,
		_w15666_
	);
	LUT2 #(
		.INIT('h2)
	) name15135 (
		\u0_w_reg[3][17]/P0001 ,
		_w15666_,
		_w15667_
	);
	LUT2 #(
		.INIT('h1)
	) name15136 (
		_w15656_,
		_w15661_,
		_w15668_
	);
	LUT2 #(
		.INIT('h4)
	) name15137 (
		_w15659_,
		_w15668_,
		_w15669_
	);
	LUT2 #(
		.INIT('h4)
	) name15138 (
		_w15654_,
		_w15669_,
		_w15670_
	);
	LUT2 #(
		.INIT('h4)
	) name15139 (
		_w15667_,
		_w15670_,
		_w15671_
	);
	LUT2 #(
		.INIT('h4)
	) name15140 (
		_w15646_,
		_w15671_,
		_w15672_
	);
	LUT2 #(
		.INIT('h4)
	) name15141 (
		_w15573_,
		_w15672_,
		_w15673_
	);
	LUT2 #(
		.INIT('h4)
	) name15142 (
		_w15636_,
		_w15673_,
		_w15674_
	);
	LUT2 #(
		.INIT('h2)
	) name15143 (
		\u0_r0_out_reg[29]/P0001 ,
		_w15674_,
		_w15675_
	);
	LUT2 #(
		.INIT('h4)
	) name15144 (
		\u0_r0_out_reg[29]/P0001 ,
		_w15674_,
		_w15676_
	);
	LUT2 #(
		.INIT('h1)
	) name15145 (
		_w15675_,
		_w15676_,
		_w15677_
	);
	LUT2 #(
		.INIT('h1)
	) name15146 (
		\u0_w_reg[0][29]/P0001 ,
		_w15677_,
		_w15678_
	);
	LUT2 #(
		.INIT('h8)
	) name15147 (
		\u0_w_reg[0][29]/P0001 ,
		_w15677_,
		_w15679_
	);
	LUT2 #(
		.INIT('h1)
	) name15148 (
		ld_pad,
		_w15678_,
		_w15680_
	);
	LUT2 #(
		.INIT('h4)
	) name15149 (
		_w15679_,
		_w15680_,
		_w15681_
	);
	LUT2 #(
		.INIT('h8)
	) name15150 (
		\key[125]_pad ,
		ld_pad,
		_w15682_
	);
	LUT2 #(
		.INIT('h1)
	) name15151 (
		_w15681_,
		_w15682_,
		_w15683_
	);
	LUT2 #(
		.INIT('h4)
	) name15152 (
		\key[61]_pad ,
		ld_pad,
		_w15684_
	);
	LUT2 #(
		.INIT('h2)
	) name15153 (
		\u0_w_reg[0][29]/P0001 ,
		\u0_w_reg[1][29]/P0002 ,
		_w15685_
	);
	LUT2 #(
		.INIT('h4)
	) name15154 (
		\u0_w_reg[0][29]/P0001 ,
		\u0_w_reg[1][29]/P0002 ,
		_w15686_
	);
	LUT2 #(
		.INIT('h1)
	) name15155 (
		_w15685_,
		_w15686_,
		_w15687_
	);
	LUT2 #(
		.INIT('h8)
	) name15156 (
		\u0_w_reg[2][29]/P0001 ,
		_w15687_,
		_w15688_
	);
	LUT2 #(
		.INIT('h1)
	) name15157 (
		\u0_w_reg[2][29]/P0001 ,
		_w15687_,
		_w15689_
	);
	LUT2 #(
		.INIT('h1)
	) name15158 (
		_w15688_,
		_w15689_,
		_w15690_
	);
	LUT2 #(
		.INIT('h8)
	) name15159 (
		_w15677_,
		_w15690_,
		_w15691_
	);
	LUT2 #(
		.INIT('h1)
	) name15160 (
		_w15677_,
		_w15690_,
		_w15692_
	);
	LUT2 #(
		.INIT('h1)
	) name15161 (
		_w15691_,
		_w15692_,
		_w15693_
	);
	LUT2 #(
		.INIT('h4)
	) name15162 (
		ld_pad,
		_w15693_,
		_w15694_
	);
	LUT2 #(
		.INIT('h1)
	) name15163 (
		_w15684_,
		_w15694_,
		_w15695_
	);
	LUT2 #(
		.INIT('h4)
	) name15164 (
		\u0_w_reg[3][29]/P0001 ,
		_w15693_,
		_w15696_
	);
	LUT2 #(
		.INIT('h2)
	) name15165 (
		\u0_w_reg[3][29]/P0001 ,
		_w15693_,
		_w15697_
	);
	LUT2 #(
		.INIT('h1)
	) name15166 (
		ld_pad,
		_w15696_,
		_w15698_
	);
	LUT2 #(
		.INIT('h4)
	) name15167 (
		_w15697_,
		_w15698_,
		_w15699_
	);
	LUT2 #(
		.INIT('h8)
	) name15168 (
		\key[29]_pad ,
		ld_pad,
		_w15700_
	);
	LUT2 #(
		.INIT('h1)
	) name15169 (
		_w15699_,
		_w15700_,
		_w15701_
	);
	LUT2 #(
		.INIT('h4)
	) name15170 (
		\key[53]_pad ,
		ld_pad,
		_w15702_
	);
	LUT2 #(
		.INIT('h8)
	) name15171 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w15703_
	);
	LUT2 #(
		.INIT('h8)
	) name15172 (
		\u0_w_reg[3][14]/P0001 ,
		_w15703_,
		_w15704_
	);
	LUT2 #(
		.INIT('h8)
	) name15173 (
		\u0_w_reg[3][13]/P0001 ,
		_w15704_,
		_w15705_
	);
	LUT2 #(
		.INIT('h4)
	) name15174 (
		\u0_w_reg[3][11]/P0001 ,
		_w15705_,
		_w15706_
	);
	LUT2 #(
		.INIT('h2)
	) name15175 (
		\u0_w_reg[3][10]/P0001 ,
		_w15706_,
		_w15707_
	);
	LUT2 #(
		.INIT('h4)
	) name15176 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w15708_
	);
	LUT2 #(
		.INIT('h1)
	) name15177 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		_w15709_
	);
	LUT2 #(
		.INIT('h8)
	) name15178 (
		_w15708_,
		_w15709_,
		_w15710_
	);
	LUT2 #(
		.INIT('h4)
	) name15179 (
		\u0_w_reg[3][15]/P0001 ,
		_w15710_,
		_w15711_
	);
	LUT2 #(
		.INIT('h2)
	) name15180 (
		_w15707_,
		_w15711_,
		_w15712_
	);
	LUT2 #(
		.INIT('h8)
	) name15181 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w15713_
	);
	LUT2 #(
		.INIT('h2)
	) name15182 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w15714_
	);
	LUT2 #(
		.INIT('h8)
	) name15183 (
		_w15713_,
		_w15714_,
		_w15715_
	);
	LUT2 #(
		.INIT('h4)
	) name15184 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w15716_
	);
	LUT2 #(
		.INIT('h8)
	) name15185 (
		_w15714_,
		_w15716_,
		_w15717_
	);
	LUT2 #(
		.INIT('h1)
	) name15186 (
		_w15715_,
		_w15717_,
		_w15718_
	);
	LUT2 #(
		.INIT('h2)
	) name15187 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w15719_
	);
	LUT2 #(
		.INIT('h4)
	) name15188 (
		\u0_w_reg[3][12]/P0001 ,
		_w15719_,
		_w15720_
	);
	LUT2 #(
		.INIT('h1)
	) name15189 (
		\u0_w_reg[3][10]/P0001 ,
		_w15720_,
		_w15721_
	);
	LUT2 #(
		.INIT('h8)
	) name15190 (
		_w15718_,
		_w15721_,
		_w15722_
	);
	LUT2 #(
		.INIT('h1)
	) name15191 (
		_w15712_,
		_w15722_,
		_w15723_
	);
	LUT2 #(
		.INIT('h2)
	) name15192 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		_w15724_
	);
	LUT2 #(
		.INIT('h2)
	) name15193 (
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w15725_
	);
	LUT2 #(
		.INIT('h4)
	) name15194 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w15726_
	);
	LUT2 #(
		.INIT('h1)
	) name15195 (
		_w15725_,
		_w15726_,
		_w15727_
	);
	LUT2 #(
		.INIT('h8)
	) name15196 (
		\u0_w_reg[3][13]/P0001 ,
		_w15724_,
		_w15728_
	);
	LUT2 #(
		.INIT('h4)
	) name15197 (
		_w15727_,
		_w15728_,
		_w15729_
	);
	LUT2 #(
		.INIT('h4)
	) name15198 (
		\u0_w_reg[3][10]/P0001 ,
		_w15708_,
		_w15730_
	);
	LUT2 #(
		.INIT('h8)
	) name15199 (
		_w15703_,
		_w15730_,
		_w15731_
	);
	LUT2 #(
		.INIT('h1)
	) name15200 (
		\u0_w_reg[3][13]/P0001 ,
		_w15716_,
		_w15732_
	);
	LUT2 #(
		.INIT('h4)
	) name15201 (
		_w15703_,
		_w15726_,
		_w15733_
	);
	LUT2 #(
		.INIT('h8)
	) name15202 (
		_w15732_,
		_w15733_,
		_w15734_
	);
	LUT2 #(
		.INIT('h8)
	) name15203 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		_w15735_
	);
	LUT2 #(
		.INIT('h1)
	) name15204 (
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w15736_
	);
	LUT2 #(
		.INIT('h8)
	) name15205 (
		_w15735_,
		_w15736_,
		_w15737_
	);
	LUT2 #(
		.INIT('h4)
	) name15206 (
		\u0_w_reg[3][12]/P0001 ,
		_w15708_,
		_w15738_
	);
	LUT2 #(
		.INIT('h1)
	) name15207 (
		_w15737_,
		_w15738_,
		_w15739_
	);
	LUT2 #(
		.INIT('h2)
	) name15208 (
		\u0_w_reg[3][10]/P0001 ,
		_w15739_,
		_w15740_
	);
	LUT2 #(
		.INIT('h8)
	) name15209 (
		\u0_w_reg[3][13]/P0001 ,
		_w15725_,
		_w15741_
	);
	LUT2 #(
		.INIT('h4)
	) name15210 (
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w15742_
	);
	LUT2 #(
		.INIT('h8)
	) name15211 (
		\u0_w_reg[3][11]/P0001 ,
		_w15742_,
		_w15743_
	);
	LUT2 #(
		.INIT('h4)
	) name15212 (
		\u0_w_reg[3][13]/P0001 ,
		_w15743_,
		_w15744_
	);
	LUT2 #(
		.INIT('h1)
	) name15213 (
		_w15741_,
		_w15744_,
		_w15745_
	);
	LUT2 #(
		.INIT('h1)
	) name15214 (
		\u0_w_reg[3][10]/P0001 ,
		_w15745_,
		_w15746_
	);
	LUT2 #(
		.INIT('h1)
	) name15215 (
		\u0_w_reg[3][9]/P0001 ,
		_w15715_,
		_w15747_
	);
	LUT2 #(
		.INIT('h4)
	) name15216 (
		_w15706_,
		_w15747_,
		_w15748_
	);
	LUT2 #(
		.INIT('h4)
	) name15217 (
		_w15740_,
		_w15748_,
		_w15749_
	);
	LUT2 #(
		.INIT('h4)
	) name15218 (
		_w15746_,
		_w15749_,
		_w15750_
	);
	LUT2 #(
		.INIT('h4)
	) name15219 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		_w15751_
	);
	LUT2 #(
		.INIT('h8)
	) name15220 (
		_w15742_,
		_w15751_,
		_w15752_
	);
	LUT2 #(
		.INIT('h8)
	) name15221 (
		\u0_w_reg[3][13]/P0001 ,
		_w15752_,
		_w15753_
	);
	LUT2 #(
		.INIT('h4)
	) name15222 (
		\u0_w_reg[3][14]/P0001 ,
		_w15735_,
		_w15754_
	);
	LUT2 #(
		.INIT('h8)
	) name15223 (
		_w15719_,
		_w15754_,
		_w15755_
	);
	LUT2 #(
		.INIT('h1)
	) name15224 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w15756_
	);
	LUT2 #(
		.INIT('h2)
	) name15225 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w15757_
	);
	LUT2 #(
		.INIT('h8)
	) name15226 (
		_w15756_,
		_w15757_,
		_w15758_
	);
	LUT2 #(
		.INIT('h4)
	) name15227 (
		\u0_w_reg[3][11]/P0001 ,
		_w15758_,
		_w15759_
	);
	LUT2 #(
		.INIT('h2)
	) name15228 (
		\u0_w_reg[3][9]/P0001 ,
		_w15759_,
		_w15760_
	);
	LUT2 #(
		.INIT('h4)
	) name15229 (
		\u0_w_reg[3][12]/P0001 ,
		_w15743_,
		_w15761_
	);
	LUT2 #(
		.INIT('h1)
	) name15230 (
		_w15753_,
		_w15755_,
		_w15762_
	);
	LUT2 #(
		.INIT('h4)
	) name15231 (
		_w15761_,
		_w15762_,
		_w15763_
	);
	LUT2 #(
		.INIT('h8)
	) name15232 (
		_w15760_,
		_w15763_,
		_w15764_
	);
	LUT2 #(
		.INIT('h1)
	) name15233 (
		_w15750_,
		_w15764_,
		_w15765_
	);
	LUT2 #(
		.INIT('h2)
	) name15234 (
		\u0_w_reg[3][8]/P0001 ,
		_w15729_,
		_w15766_
	);
	LUT2 #(
		.INIT('h1)
	) name15235 (
		_w15731_,
		_w15734_,
		_w15767_
	);
	LUT2 #(
		.INIT('h8)
	) name15236 (
		_w15766_,
		_w15767_,
		_w15768_
	);
	LUT2 #(
		.INIT('h4)
	) name15237 (
		_w15723_,
		_w15768_,
		_w15769_
	);
	LUT2 #(
		.INIT('h4)
	) name15238 (
		_w15765_,
		_w15769_,
		_w15770_
	);
	LUT2 #(
		.INIT('h4)
	) name15239 (
		\u0_w_reg[3][12]/P0001 ,
		_w15725_,
		_w15771_
	);
	LUT2 #(
		.INIT('h4)
	) name15240 (
		\u0_w_reg[3][11]/P0001 ,
		_w15771_,
		_w15772_
	);
	LUT2 #(
		.INIT('h2)
	) name15241 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w15773_
	);
	LUT2 #(
		.INIT('h8)
	) name15242 (
		_w15751_,
		_w15773_,
		_w15774_
	);
	LUT2 #(
		.INIT('h1)
	) name15243 (
		_w15743_,
		_w15774_,
		_w15775_
	);
	LUT2 #(
		.INIT('h4)
	) name15244 (
		_w15772_,
		_w15775_,
		_w15776_
	);
	LUT2 #(
		.INIT('h1)
	) name15245 (
		\u0_w_reg[3][10]/P0001 ,
		_w15776_,
		_w15777_
	);
	LUT2 #(
		.INIT('h4)
	) name15246 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w15778_
	);
	LUT2 #(
		.INIT('h8)
	) name15247 (
		_w15773_,
		_w15778_,
		_w15779_
	);
	LUT2 #(
		.INIT('h8)
	) name15248 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w15780_
	);
	LUT2 #(
		.INIT('h8)
	) name15249 (
		\u0_w_reg[3][11]/P0001 ,
		_w15780_,
		_w15781_
	);
	LUT2 #(
		.INIT('h1)
	) name15250 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		_w15782_
	);
	LUT2 #(
		.INIT('h2)
	) name15251 (
		_w15781_,
		_w15782_,
		_w15783_
	);
	LUT2 #(
		.INIT('h4)
	) name15252 (
		\u0_w_reg[3][11]/P0001 ,
		_w15741_,
		_w15784_
	);
	LUT2 #(
		.INIT('h4)
	) name15253 (
		\u0_w_reg[3][12]/P0001 ,
		_w15784_,
		_w15785_
	);
	LUT2 #(
		.INIT('h8)
	) name15254 (
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w15786_
	);
	LUT2 #(
		.INIT('h4)
	) name15255 (
		\u0_w_reg[3][13]/P0001 ,
		_w15786_,
		_w15787_
	);
	LUT2 #(
		.INIT('h4)
	) name15256 (
		\u0_w_reg[3][11]/P0001 ,
		_w15787_,
		_w15788_
	);
	LUT2 #(
		.INIT('h8)
	) name15257 (
		_w15714_,
		_w15756_,
		_w15789_
	);
	LUT2 #(
		.INIT('h2)
	) name15258 (
		\u0_w_reg[3][9]/P0001 ,
		_w15789_,
		_w15790_
	);
	LUT2 #(
		.INIT('h8)
	) name15259 (
		\u0_w_reg[3][10]/P0001 ,
		_w15713_,
		_w15791_
	);
	LUT2 #(
		.INIT('h8)
	) name15260 (
		_w15757_,
		_w15791_,
		_w15792_
	);
	LUT2 #(
		.INIT('h1)
	) name15261 (
		_w15779_,
		_w15783_,
		_w15793_
	);
	LUT2 #(
		.INIT('h4)
	) name15262 (
		_w15788_,
		_w15790_,
		_w15794_
	);
	LUT2 #(
		.INIT('h4)
	) name15263 (
		_w15792_,
		_w15794_,
		_w15795_
	);
	LUT2 #(
		.INIT('h4)
	) name15264 (
		_w15785_,
		_w15793_,
		_w15796_
	);
	LUT2 #(
		.INIT('h8)
	) name15265 (
		_w15795_,
		_w15796_,
		_w15797_
	);
	LUT2 #(
		.INIT('h4)
	) name15266 (
		_w15777_,
		_w15797_,
		_w15798_
	);
	LUT2 #(
		.INIT('h8)
	) name15267 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w15799_
	);
	LUT2 #(
		.INIT('h4)
	) name15268 (
		\u0_w_reg[3][12]/P0001 ,
		_w15799_,
		_w15800_
	);
	LUT2 #(
		.INIT('h8)
	) name15269 (
		_w15756_,
		_w15800_,
		_w15801_
	);
	LUT2 #(
		.INIT('h8)
	) name15270 (
		_w15703_,
		_w15756_,
		_w15802_
	);
	LUT2 #(
		.INIT('h2)
	) name15271 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		_w15803_
	);
	LUT2 #(
		.INIT('h8)
	) name15272 (
		_w15736_,
		_w15803_,
		_w15804_
	);
	LUT2 #(
		.INIT('h8)
	) name15273 (
		_w15716_,
		_w15780_,
		_w15805_
	);
	LUT2 #(
		.INIT('h1)
	) name15274 (
		_w15802_,
		_w15804_,
		_w15806_
	);
	LUT2 #(
		.INIT('h4)
	) name15275 (
		_w15805_,
		_w15806_,
		_w15807_
	);
	LUT2 #(
		.INIT('h1)
	) name15276 (
		\u0_w_reg[3][11]/P0001 ,
		_w15807_,
		_w15808_
	);
	LUT2 #(
		.INIT('h1)
	) name15277 (
		\u0_w_reg[3][9]/P0001 ,
		_w15801_,
		_w15809_
	);
	LUT2 #(
		.INIT('h4)
	) name15278 (
		_w15808_,
		_w15809_,
		_w15810_
	);
	LUT2 #(
		.INIT('h1)
	) name15279 (
		_w15798_,
		_w15810_,
		_w15811_
	);
	LUT2 #(
		.INIT('h4)
	) name15280 (
		\u0_w_reg[3][13]/P0001 ,
		_w15757_,
		_w15812_
	);
	LUT2 #(
		.INIT('h8)
	) name15281 (
		\u0_w_reg[3][11]/P0001 ,
		_w15812_,
		_w15813_
	);
	LUT2 #(
		.INIT('h4)
	) name15282 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w15814_
	);
	LUT2 #(
		.INIT('h8)
	) name15283 (
		_w15716_,
		_w15814_,
		_w15815_
	);
	LUT2 #(
		.INIT('h1)
	) name15284 (
		_w15813_,
		_w15815_,
		_w15816_
	);
	LUT2 #(
		.INIT('h8)
	) name15285 (
		_w15703_,
		_w15773_,
		_w15817_
	);
	LUT2 #(
		.INIT('h1)
	) name15286 (
		\u0_w_reg[3][10]/P0001 ,
		_w15817_,
		_w15818_
	);
	LUT2 #(
		.INIT('h8)
	) name15287 (
		_w15816_,
		_w15818_,
		_w15819_
	);
	LUT2 #(
		.INIT('h4)
	) name15288 (
		\u0_w_reg[3][12]/P0001 ,
		_w15736_,
		_w15820_
	);
	LUT2 #(
		.INIT('h8)
	) name15289 (
		\u0_w_reg[3][12]/P0001 ,
		_w15780_,
		_w15821_
	);
	LUT2 #(
		.INIT('h1)
	) name15290 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w15822_
	);
	LUT2 #(
		.INIT('h4)
	) name15291 (
		\u0_w_reg[3][13]/P0001 ,
		_w15822_,
		_w15823_
	);
	LUT2 #(
		.INIT('h1)
	) name15292 (
		_w15821_,
		_w15823_,
		_w15824_
	);
	LUT2 #(
		.INIT('h2)
	) name15293 (
		\u0_w_reg[3][11]/P0001 ,
		_w15824_,
		_w15825_
	);
	LUT2 #(
		.INIT('h8)
	) name15294 (
		_w15708_,
		_w15757_,
		_w15826_
	);
	LUT2 #(
		.INIT('h4)
	) name15295 (
		\u0_w_reg[3][11]/P0001 ,
		_w15826_,
		_w15827_
	);
	LUT2 #(
		.INIT('h2)
	) name15296 (
		\u0_w_reg[3][10]/P0001 ,
		_w15820_,
		_w15828_
	);
	LUT2 #(
		.INIT('h4)
	) name15297 (
		_w15827_,
		_w15828_,
		_w15829_
	);
	LUT2 #(
		.INIT('h4)
	) name15298 (
		_w15825_,
		_w15829_,
		_w15830_
	);
	LUT2 #(
		.INIT('h1)
	) name15299 (
		_w15819_,
		_w15830_,
		_w15831_
	);
	LUT2 #(
		.INIT('h8)
	) name15300 (
		_w15756_,
		_w15822_,
		_w15832_
	);
	LUT2 #(
		.INIT('h1)
	) name15301 (
		\u0_w_reg[3][8]/P0001 ,
		_w15832_,
		_w15833_
	);
	LUT2 #(
		.INIT('h4)
	) name15302 (
		_w15831_,
		_w15833_,
		_w15834_
	);
	LUT2 #(
		.INIT('h4)
	) name15303 (
		_w15811_,
		_w15834_,
		_w15835_
	);
	LUT2 #(
		.INIT('h1)
	) name15304 (
		_w15770_,
		_w15835_,
		_w15836_
	);
	LUT2 #(
		.INIT('h8)
	) name15305 (
		_w15735_,
		_w15773_,
		_w15837_
	);
	LUT2 #(
		.INIT('h4)
	) name15306 (
		\u0_w_reg[3][13]/P0001 ,
		_w15725_,
		_w15838_
	);
	LUT2 #(
		.INIT('h4)
	) name15307 (
		\u0_w_reg[3][13]/P0001 ,
		_w15742_,
		_w15839_
	);
	LUT2 #(
		.INIT('h8)
	) name15308 (
		\u0_w_reg[3][13]/P0001 ,
		_w15786_,
		_w15840_
	);
	LUT2 #(
		.INIT('h1)
	) name15309 (
		_w15838_,
		_w15839_,
		_w15841_
	);
	LUT2 #(
		.INIT('h4)
	) name15310 (
		_w15840_,
		_w15841_,
		_w15842_
	);
	LUT2 #(
		.INIT('h2)
	) name15311 (
		_w15751_,
		_w15842_,
		_w15843_
	);
	LUT2 #(
		.INIT('h1)
	) name15312 (
		_w15837_,
		_w15843_,
		_w15844_
	);
	LUT2 #(
		.INIT('h2)
	) name15313 (
		\u0_w_reg[3][10]/P0001 ,
		_w15844_,
		_w15845_
	);
	LUT2 #(
		.INIT('h4)
	) name15314 (
		\u0_w_reg[3][12]/P0001 ,
		_w15780_,
		_w15846_
	);
	LUT2 #(
		.INIT('h1)
	) name15315 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w15847_
	);
	LUT2 #(
		.INIT('h8)
	) name15316 (
		_w15846_,
		_w15847_,
		_w15848_
	);
	LUT2 #(
		.INIT('h4)
	) name15317 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w15849_
	);
	LUT2 #(
		.INIT('h8)
	) name15318 (
		\u0_w_reg[3][12]/P0001 ,
		_w15725_,
		_w15850_
	);
	LUT2 #(
		.INIT('h8)
	) name15319 (
		\u0_w_reg[3][13]/P0001 ,
		_w15850_,
		_w15851_
	);
	LUT2 #(
		.INIT('h8)
	) name15320 (
		_w15849_,
		_w15851_,
		_w15852_
	);
	LUT2 #(
		.INIT('h8)
	) name15321 (
		_w15709_,
		_w15736_,
		_w15853_
	);
	LUT2 #(
		.INIT('h1)
	) name15322 (
		_w15731_,
		_w15853_,
		_w15854_
	);
	LUT2 #(
		.INIT('h4)
	) name15323 (
		_w15848_,
		_w15854_,
		_w15855_
	);
	LUT2 #(
		.INIT('h4)
	) name15324 (
		_w15852_,
		_w15855_,
		_w15856_
	);
	LUT2 #(
		.INIT('h4)
	) name15325 (
		_w15845_,
		_w15856_,
		_w15857_
	);
	LUT2 #(
		.INIT('h1)
	) name15326 (
		\u0_w_reg[3][9]/P0001 ,
		_w15857_,
		_w15858_
	);
	LUT2 #(
		.INIT('h8)
	) name15327 (
		_w15719_,
		_w15735_,
		_w15859_
	);
	LUT2 #(
		.INIT('h2)
	) name15328 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w15860_
	);
	LUT2 #(
		.INIT('h8)
	) name15329 (
		_w15859_,
		_w15860_,
		_w15861_
	);
	LUT2 #(
		.INIT('h4)
	) name15330 (
		\u0_w_reg[3][14]/P0001 ,
		_w15724_,
		_w15862_
	);
	LUT2 #(
		.INIT('h8)
	) name15331 (
		_w15719_,
		_w15862_,
		_w15863_
	);
	LUT2 #(
		.INIT('h4)
	) name15332 (
		\u0_w_reg[3][10]/P0001 ,
		_w15863_,
		_w15864_
	);
	LUT2 #(
		.INIT('h8)
	) name15333 (
		_w15724_,
		_w15736_,
		_w15865_
	);
	LUT2 #(
		.INIT('h4)
	) name15334 (
		\u0_w_reg[3][13]/P0001 ,
		_w15865_,
		_w15866_
	);
	LUT2 #(
		.INIT('h4)
	) name15335 (
		\u0_w_reg[3][10]/P0001 ,
		_w15817_,
		_w15867_
	);
	LUT2 #(
		.INIT('h4)
	) name15336 (
		\u0_w_reg[3][11]/P0001 ,
		_w15792_,
		_w15868_
	);
	LUT2 #(
		.INIT('h1)
	) name15337 (
		_w15866_,
		_w15867_,
		_w15869_
	);
	LUT2 #(
		.INIT('h4)
	) name15338 (
		_w15868_,
		_w15869_,
		_w15870_
	);
	LUT2 #(
		.INIT('h2)
	) name15339 (
		\u0_w_reg[3][9]/P0001 ,
		_w15870_,
		_w15871_
	);
	LUT2 #(
		.INIT('h4)
	) name15340 (
		\u0_w_reg[3][10]/P0001 ,
		_w15788_,
		_w15872_
	);
	LUT2 #(
		.INIT('h1)
	) name15341 (
		_w15861_,
		_w15864_,
		_w15873_
	);
	LUT2 #(
		.INIT('h4)
	) name15342 (
		_w15872_,
		_w15873_,
		_w15874_
	);
	LUT2 #(
		.INIT('h4)
	) name15343 (
		_w15871_,
		_w15874_,
		_w15875_
	);
	LUT2 #(
		.INIT('h4)
	) name15344 (
		_w15858_,
		_w15875_,
		_w15876_
	);
	LUT2 #(
		.INIT('h4)
	) name15345 (
		_w15836_,
		_w15876_,
		_w15877_
	);
	LUT2 #(
		.INIT('h2)
	) name15346 (
		\u0_w_reg[0][21]/P0001 ,
		_w15877_,
		_w15878_
	);
	LUT2 #(
		.INIT('h4)
	) name15347 (
		\u0_w_reg[0][21]/P0001 ,
		_w15877_,
		_w15879_
	);
	LUT2 #(
		.INIT('h1)
	) name15348 (
		_w15878_,
		_w15879_,
		_w15880_
	);
	LUT2 #(
		.INIT('h2)
	) name15349 (
		\u0_w_reg[1][21]/P0001 ,
		\u0_w_reg[2][21]/P0001 ,
		_w15881_
	);
	LUT2 #(
		.INIT('h4)
	) name15350 (
		\u0_w_reg[1][21]/P0001 ,
		\u0_w_reg[2][21]/P0001 ,
		_w15882_
	);
	LUT2 #(
		.INIT('h1)
	) name15351 (
		_w15881_,
		_w15882_,
		_w15883_
	);
	LUT2 #(
		.INIT('h8)
	) name15352 (
		_w15880_,
		_w15883_,
		_w15884_
	);
	LUT2 #(
		.INIT('h1)
	) name15353 (
		_w15880_,
		_w15883_,
		_w15885_
	);
	LUT2 #(
		.INIT('h1)
	) name15354 (
		_w15884_,
		_w15885_,
		_w15886_
	);
	LUT2 #(
		.INIT('h4)
	) name15355 (
		ld_pad,
		_w15886_,
		_w15887_
	);
	LUT2 #(
		.INIT('h1)
	) name15356 (
		_w15702_,
		_w15887_,
		_w15888_
	);
	LUT2 #(
		.INIT('h4)
	) name15357 (
		\key[51]_pad ,
		ld_pad,
		_w15889_
	);
	LUT2 #(
		.INIT('h1)
	) name15358 (
		_w15756_,
		_w15860_,
		_w15890_
	);
	LUT2 #(
		.INIT('h2)
	) name15359 (
		_w15757_,
		_w15890_,
		_w15891_
	);
	LUT2 #(
		.INIT('h8)
	) name15360 (
		\u0_w_reg[3][11]/P0001 ,
		_w15867_,
		_w15892_
	);
	LUT2 #(
		.INIT('h2)
	) name15361 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w15893_
	);
	LUT2 #(
		.INIT('h2)
	) name15362 (
		\u0_w_reg[3][15]/P0001 ,
		_w15756_,
		_w15894_
	);
	LUT2 #(
		.INIT('h8)
	) name15363 (
		_w15893_,
		_w15894_,
		_w15895_
	);
	LUT2 #(
		.INIT('h4)
	) name15364 (
		\u0_w_reg[3][11]/P0001 ,
		_w15778_,
		_w15896_
	);
	LUT2 #(
		.INIT('h4)
	) name15365 (
		\u0_w_reg[3][13]/P0001 ,
		_w15896_,
		_w15897_
	);
	LUT2 #(
		.INIT('h1)
	) name15366 (
		\u0_w_reg[3][9]/P0001 ,
		_w15891_,
		_w15898_
	);
	LUT2 #(
		.INIT('h1)
	) name15367 (
		_w15895_,
		_w15897_,
		_w15899_
	);
	LUT2 #(
		.INIT('h8)
	) name15368 (
		_w15898_,
		_w15899_,
		_w15900_
	);
	LUT2 #(
		.INIT('h4)
	) name15369 (
		_w15892_,
		_w15900_,
		_w15901_
	);
	LUT2 #(
		.INIT('h8)
	) name15370 (
		_w15713_,
		_w15751_,
		_w15902_
	);
	LUT2 #(
		.INIT('h4)
	) name15371 (
		\u0_w_reg[3][15]/P0001 ,
		_w15902_,
		_w15903_
	);
	LUT2 #(
		.INIT('h1)
	) name15372 (
		_w15823_,
		_w15903_,
		_w15904_
	);
	LUT2 #(
		.INIT('h2)
	) name15373 (
		\u0_w_reg[3][10]/P0001 ,
		_w15904_,
		_w15905_
	);
	LUT2 #(
		.INIT('h8)
	) name15374 (
		\u0_w_reg[3][15]/P0001 ,
		_w15735_,
		_w15906_
	);
	LUT2 #(
		.INIT('h1)
	) name15375 (
		_w15896_,
		_w15906_,
		_w15907_
	);
	LUT2 #(
		.INIT('h2)
	) name15376 (
		_w15713_,
		_w15907_,
		_w15908_
	);
	LUT2 #(
		.INIT('h4)
	) name15377 (
		\u0_w_reg[3][10]/P0001 ,
		_w15779_,
		_w15909_
	);
	LUT2 #(
		.INIT('h2)
	) name15378 (
		\u0_w_reg[3][9]/P0001 ,
		_w15744_,
		_w15910_
	);
	LUT2 #(
		.INIT('h4)
	) name15379 (
		_w15909_,
		_w15910_,
		_w15911_
	);
	LUT2 #(
		.INIT('h4)
	) name15380 (
		_w15908_,
		_w15911_,
		_w15912_
	);
	LUT2 #(
		.INIT('h4)
	) name15381 (
		_w15905_,
		_w15912_,
		_w15913_
	);
	LUT2 #(
		.INIT('h1)
	) name15382 (
		_w15901_,
		_w15913_,
		_w15914_
	);
	LUT2 #(
		.INIT('h4)
	) name15383 (
		\u0_w_reg[3][12]/P0001 ,
		_w15714_,
		_w15915_
	);
	LUT2 #(
		.INIT('h4)
	) name15384 (
		\u0_w_reg[3][13]/P0001 ,
		_w15915_,
		_w15916_
	);
	LUT2 #(
		.INIT('h1)
	) name15385 (
		_w15805_,
		_w15916_,
		_w15917_
	);
	LUT2 #(
		.INIT('h2)
	) name15386 (
		\u0_w_reg[3][10]/P0001 ,
		_w15917_,
		_w15918_
	);
	LUT2 #(
		.INIT('h8)
	) name15387 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w15919_
	);
	LUT2 #(
		.INIT('h8)
	) name15388 (
		_w15757_,
		_w15919_,
		_w15920_
	);
	LUT2 #(
		.INIT('h1)
	) name15389 (
		_w15706_,
		_w15920_,
		_w15921_
	);
	LUT2 #(
		.INIT('h1)
	) name15390 (
		\u0_w_reg[3][10]/P0001 ,
		_w15921_,
		_w15922_
	);
	LUT2 #(
		.INIT('h1)
	) name15391 (
		_w15711_,
		_w15918_,
		_w15923_
	);
	LUT2 #(
		.INIT('h4)
	) name15392 (
		_w15922_,
		_w15923_,
		_w15924_
	);
	LUT2 #(
		.INIT('h4)
	) name15393 (
		_w15914_,
		_w15924_,
		_w15925_
	);
	LUT2 #(
		.INIT('h1)
	) name15394 (
		\u0_w_reg[3][8]/P0001 ,
		_w15925_,
		_w15926_
	);
	LUT2 #(
		.INIT('h4)
	) name15395 (
		_w15720_,
		_w15745_,
		_w15927_
	);
	LUT2 #(
		.INIT('h2)
	) name15396 (
		\u0_w_reg[3][10]/P0001 ,
		_w15927_,
		_w15928_
	);
	LUT2 #(
		.INIT('h8)
	) name15397 (
		\u0_w_reg[3][13]/P0001 ,
		_w15709_,
		_w15929_
	);
	LUT2 #(
		.INIT('h8)
	) name15398 (
		\u0_w_reg[3][14]/P0001 ,
		_w15929_,
		_w15930_
	);
	LUT2 #(
		.INIT('h8)
	) name15399 (
		_w15838_,
		_w15849_,
		_w15931_
	);
	LUT2 #(
		.INIT('h8)
	) name15400 (
		\u0_w_reg[3][11]/P0001 ,
		_w15802_,
		_w15932_
	);
	LUT2 #(
		.INIT('h1)
	) name15401 (
		_w15853_,
		_w15930_,
		_w15933_
	);
	LUT2 #(
		.INIT('h1)
	) name15402 (
		_w15931_,
		_w15932_,
		_w15934_
	);
	LUT2 #(
		.INIT('h8)
	) name15403 (
		_w15933_,
		_w15934_,
		_w15935_
	);
	LUT2 #(
		.INIT('h4)
	) name15404 (
		_w15872_,
		_w15935_,
		_w15936_
	);
	LUT2 #(
		.INIT('h4)
	) name15405 (
		_w15928_,
		_w15936_,
		_w15937_
	);
	LUT2 #(
		.INIT('h1)
	) name15406 (
		\u0_w_reg[3][9]/P0001 ,
		_w15937_,
		_w15938_
	);
	LUT2 #(
		.INIT('h8)
	) name15407 (
		_w15814_,
		_w15919_,
		_w15939_
	);
	LUT2 #(
		.INIT('h1)
	) name15408 (
		_w15817_,
		_w15939_,
		_w15940_
	);
	LUT2 #(
		.INIT('h8)
	) name15409 (
		_w15751_,
		_w15780_,
		_w15941_
	);
	LUT2 #(
		.INIT('h4)
	) name15410 (
		\u0_w_reg[3][11]/P0001 ,
		_w15725_,
		_w15942_
	);
	LUT2 #(
		.INIT('h4)
	) name15411 (
		\u0_w_reg[3][13]/P0001 ,
		_w15736_,
		_w15943_
	);
	LUT2 #(
		.INIT('h1)
	) name15412 (
		\u0_w_reg[3][10]/P0001 ,
		_w15942_,
		_w15944_
	);
	LUT2 #(
		.INIT('h4)
	) name15413 (
		_w15943_,
		_w15944_,
		_w15945_
	);
	LUT2 #(
		.INIT('h8)
	) name15414 (
		\u0_w_reg[3][12]/P0001 ,
		_w15814_,
		_w15946_
	);
	LUT2 #(
		.INIT('h4)
	) name15415 (
		_w15714_,
		_w15773_,
		_w15947_
	);
	LUT2 #(
		.INIT('h2)
	) name15416 (
		\u0_w_reg[3][10]/P0001 ,
		_w15946_,
		_w15948_
	);
	LUT2 #(
		.INIT('h4)
	) name15417 (
		_w15947_,
		_w15948_,
		_w15949_
	);
	LUT2 #(
		.INIT('h1)
	) name15418 (
		_w15945_,
		_w15949_,
		_w15950_
	);
	LUT2 #(
		.INIT('h2)
	) name15419 (
		_w15940_,
		_w15941_,
		_w15951_
	);
	LUT2 #(
		.INIT('h4)
	) name15420 (
		_w15950_,
		_w15951_,
		_w15952_
	);
	LUT2 #(
		.INIT('h2)
	) name15421 (
		\u0_w_reg[3][9]/P0001 ,
		_w15952_,
		_w15953_
	);
	LUT2 #(
		.INIT('h8)
	) name15422 (
		_w15780_,
		_w15919_,
		_w15954_
	);
	LUT2 #(
		.INIT('h1)
	) name15423 (
		_w15897_,
		_w15954_,
		_w15955_
	);
	LUT2 #(
		.INIT('h1)
	) name15424 (
		\u0_w_reg[3][10]/P0001 ,
		_w15955_,
		_w15956_
	);
	LUT2 #(
		.INIT('h8)
	) name15425 (
		_w15713_,
		_w15724_,
		_w15957_
	);
	LUT2 #(
		.INIT('h4)
	) name15426 (
		\u0_w_reg[3][15]/P0001 ,
		_w15957_,
		_w15958_
	);
	LUT2 #(
		.INIT('h4)
	) name15427 (
		\u0_w_reg[3][11]/P0001 ,
		_w15867_,
		_w15959_
	);
	LUT2 #(
		.INIT('h8)
	) name15428 (
		_w15735_,
		_w15742_,
		_w15960_
	);
	LUT2 #(
		.INIT('h1)
	) name15429 (
		_w15802_,
		_w15826_,
		_w15961_
	);
	LUT2 #(
		.INIT('h4)
	) name15430 (
		_w15960_,
		_w15961_,
		_w15962_
	);
	LUT2 #(
		.INIT('h2)
	) name15431 (
		\u0_w_reg[3][10]/P0001 ,
		_w15962_,
		_w15963_
	);
	LUT2 #(
		.INIT('h1)
	) name15432 (
		_w15958_,
		_w15959_,
		_w15964_
	);
	LUT2 #(
		.INIT('h4)
	) name15433 (
		_w15956_,
		_w15964_,
		_w15965_
	);
	LUT2 #(
		.INIT('h4)
	) name15434 (
		_w15963_,
		_w15965_,
		_w15966_
	);
	LUT2 #(
		.INIT('h4)
	) name15435 (
		_w15953_,
		_w15966_,
		_w15967_
	);
	LUT2 #(
		.INIT('h4)
	) name15436 (
		_w15938_,
		_w15967_,
		_w15968_
	);
	LUT2 #(
		.INIT('h2)
	) name15437 (
		\u0_w_reg[3][8]/P0001 ,
		_w15968_,
		_w15969_
	);
	LUT2 #(
		.INIT('h8)
	) name15438 (
		_w15724_,
		_w15786_,
		_w15970_
	);
	LUT2 #(
		.INIT('h4)
	) name15439 (
		\u0_w_reg[3][13]/P0001 ,
		_w15970_,
		_w15971_
	);
	LUT2 #(
		.INIT('h1)
	) name15440 (
		_w15932_,
		_w15971_,
		_w15972_
	);
	LUT2 #(
		.INIT('h2)
	) name15441 (
		\u0_w_reg[3][10]/P0001 ,
		_w15972_,
		_w15973_
	);
	LUT2 #(
		.INIT('h2)
	) name15442 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w15974_
	);
	LUT2 #(
		.INIT('h4)
	) name15443 (
		\u0_w_reg[3][11]/P0001 ,
		_w15974_,
		_w15975_
	);
	LUT2 #(
		.INIT('h8)
	) name15444 (
		_w15708_,
		_w15822_,
		_w15976_
	);
	LUT2 #(
		.INIT('h1)
	) name15445 (
		_w15758_,
		_w15976_,
		_w15977_
	);
	LUT2 #(
		.INIT('h2)
	) name15446 (
		_w15975_,
		_w15977_,
		_w15978_
	);
	LUT2 #(
		.INIT('h1)
	) name15447 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w15979_
	);
	LUT2 #(
		.INIT('h8)
	) name15448 (
		_w15778_,
		_w15979_,
		_w15980_
	);
	LUT2 #(
		.INIT('h1)
	) name15449 (
		_w15812_,
		_w15980_,
		_w15981_
	);
	LUT2 #(
		.INIT('h2)
	) name15450 (
		_w15919_,
		_w15981_,
		_w15982_
	);
	LUT2 #(
		.INIT('h8)
	) name15451 (
		\u0_w_reg[3][12]/P0001 ,
		_w15756_,
		_w15983_
	);
	LUT2 #(
		.INIT('h1)
	) name15452 (
		_w15771_,
		_w15779_,
		_w15984_
	);
	LUT2 #(
		.INIT('h4)
	) name15453 (
		_w15983_,
		_w15984_,
		_w15985_
	);
	LUT2 #(
		.INIT('h2)
	) name15454 (
		_w15847_,
		_w15985_,
		_w15986_
	);
	LUT2 #(
		.INIT('h2)
	) name15455 (
		_w15940_,
		_w15957_,
		_w15987_
	);
	LUT2 #(
		.INIT('h2)
	) name15456 (
		\u0_w_reg[3][10]/P0001 ,
		_w15987_,
		_w15988_
	);
	LUT2 #(
		.INIT('h8)
	) name15457 (
		_w15756_,
		_w15778_,
		_w15989_
	);
	LUT2 #(
		.INIT('h8)
	) name15458 (
		_w15849_,
		_w15989_,
		_w15990_
	);
	LUT2 #(
		.INIT('h1)
	) name15459 (
		_w15986_,
		_w15990_,
		_w15991_
	);
	LUT2 #(
		.INIT('h4)
	) name15460 (
		_w15988_,
		_w15991_,
		_w15992_
	);
	LUT2 #(
		.INIT('h2)
	) name15461 (
		\u0_w_reg[3][9]/P0001 ,
		_w15992_,
		_w15993_
	);
	LUT2 #(
		.INIT('h1)
	) name15462 (
		_w15978_,
		_w15982_,
		_w15994_
	);
	LUT2 #(
		.INIT('h4)
	) name15463 (
		_w15973_,
		_w15994_,
		_w15995_
	);
	LUT2 #(
		.INIT('h4)
	) name15464 (
		_w15993_,
		_w15995_,
		_w15996_
	);
	LUT2 #(
		.INIT('h4)
	) name15465 (
		_w15926_,
		_w15996_,
		_w15997_
	);
	LUT2 #(
		.INIT('h4)
	) name15466 (
		_w15969_,
		_w15997_,
		_w15998_
	);
	LUT2 #(
		.INIT('h2)
	) name15467 (
		\u0_w_reg[0][19]/P0001 ,
		_w15998_,
		_w15999_
	);
	LUT2 #(
		.INIT('h4)
	) name15468 (
		\u0_w_reg[0][19]/P0001 ,
		_w15998_,
		_w16000_
	);
	LUT2 #(
		.INIT('h1)
	) name15469 (
		_w15999_,
		_w16000_,
		_w16001_
	);
	LUT2 #(
		.INIT('h2)
	) name15470 (
		\u0_w_reg[1][19]/P0001 ,
		\u0_w_reg[2][19]/P0001 ,
		_w16002_
	);
	LUT2 #(
		.INIT('h4)
	) name15471 (
		\u0_w_reg[1][19]/P0001 ,
		\u0_w_reg[2][19]/P0001 ,
		_w16003_
	);
	LUT2 #(
		.INIT('h1)
	) name15472 (
		_w16002_,
		_w16003_,
		_w16004_
	);
	LUT2 #(
		.INIT('h8)
	) name15473 (
		_w16001_,
		_w16004_,
		_w16005_
	);
	LUT2 #(
		.INIT('h1)
	) name15474 (
		_w16001_,
		_w16004_,
		_w16006_
	);
	LUT2 #(
		.INIT('h1)
	) name15475 (
		_w16005_,
		_w16006_,
		_w16007_
	);
	LUT2 #(
		.INIT('h4)
	) name15476 (
		ld_pad,
		_w16007_,
		_w16008_
	);
	LUT2 #(
		.INIT('h1)
	) name15477 (
		_w15889_,
		_w16008_,
		_w16009_
	);
	LUT2 #(
		.INIT('h4)
	) name15478 (
		\key[37]_pad ,
		ld_pad,
		_w16010_
	);
	LUT2 #(
		.INIT('h8)
	) name15479 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w16011_
	);
	LUT2 #(
		.INIT('h2)
	) name15480 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w16012_
	);
	LUT2 #(
		.INIT('h8)
	) name15481 (
		_w16011_,
		_w16012_,
		_w16013_
	);
	LUT2 #(
		.INIT('h4)
	) name15482 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w16014_
	);
	LUT2 #(
		.INIT('h8)
	) name15483 (
		_w16012_,
		_w16014_,
		_w16015_
	);
	LUT2 #(
		.INIT('h1)
	) name15484 (
		_w16013_,
		_w16015_,
		_w16016_
	);
	LUT2 #(
		.INIT('h2)
	) name15485 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w16017_
	);
	LUT2 #(
		.INIT('h4)
	) name15486 (
		\u0_w_reg[3][28]/P0001 ,
		_w16017_,
		_w16018_
	);
	LUT2 #(
		.INIT('h4)
	) name15487 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w16019_
	);
	LUT2 #(
		.INIT('h8)
	) name15488 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w16020_
	);
	LUT2 #(
		.INIT('h8)
	) name15489 (
		_w16019_,
		_w16020_,
		_w16021_
	);
	LUT2 #(
		.INIT('h1)
	) name15490 (
		_w16018_,
		_w16021_,
		_w16022_
	);
	LUT2 #(
		.INIT('h8)
	) name15491 (
		_w16016_,
		_w16022_,
		_w16023_
	);
	LUT2 #(
		.INIT('h1)
	) name15492 (
		\u0_w_reg[3][26]/P0001 ,
		_w16023_,
		_w16024_
	);
	LUT2 #(
		.INIT('h2)
	) name15493 (
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w16025_
	);
	LUT2 #(
		.INIT('h4)
	) name15494 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		_w16026_
	);
	LUT2 #(
		.INIT('h8)
	) name15495 (
		_w16025_,
		_w16026_,
		_w16027_
	);
	LUT2 #(
		.INIT('h8)
	) name15496 (
		\u0_w_reg[3][27]/P0001 ,
		_w16027_,
		_w16028_
	);
	LUT2 #(
		.INIT('h2)
	) name15497 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		_w16029_
	);
	LUT2 #(
		.INIT('h1)
	) name15498 (
		\u0_w_reg[3][29]/P0001 ,
		_w16014_,
		_w16030_
	);
	LUT2 #(
		.INIT('h4)
	) name15499 (
		_w16020_,
		_w16030_,
		_w16031_
	);
	LUT2 #(
		.INIT('h2)
	) name15500 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w16032_
	);
	LUT2 #(
		.INIT('h8)
	) name15501 (
		\u0_w_reg[3][29]/P0001 ,
		_w16032_,
		_w16033_
	);
	LUT2 #(
		.INIT('h1)
	) name15502 (
		_w16031_,
		_w16033_,
		_w16034_
	);
	LUT2 #(
		.INIT('h2)
	) name15503 (
		_w16029_,
		_w16034_,
		_w16035_
	);
	LUT2 #(
		.INIT('h2)
	) name15504 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w16036_
	);
	LUT2 #(
		.INIT('h8)
	) name15505 (
		\u0_w_reg[3][31]/P0001 ,
		_w16011_,
		_w16037_
	);
	LUT2 #(
		.INIT('h8)
	) name15506 (
		\u0_w_reg[3][28]/P0001 ,
		_w16037_,
		_w16038_
	);
	LUT2 #(
		.INIT('h1)
	) name15507 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w16039_
	);
	LUT2 #(
		.INIT('h8)
	) name15508 (
		_w16019_,
		_w16039_,
		_w16040_
	);
	LUT2 #(
		.INIT('h1)
	) name15509 (
		_w16038_,
		_w16040_,
		_w16041_
	);
	LUT2 #(
		.INIT('h2)
	) name15510 (
		_w16036_,
		_w16041_,
		_w16042_
	);
	LUT2 #(
		.INIT('h4)
	) name15511 (
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w16043_
	);
	LUT2 #(
		.INIT('h8)
	) name15512 (
		_w16032_,
		_w16043_,
		_w16044_
	);
	LUT2 #(
		.INIT('h8)
	) name15513 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w16045_
	);
	LUT2 #(
		.INIT('h4)
	) name15514 (
		\u0_w_reg[3][30]/P0001 ,
		_w16045_,
		_w16046_
	);
	LUT2 #(
		.INIT('h8)
	) name15515 (
		_w16017_,
		_w16046_,
		_w16047_
	);
	LUT2 #(
		.INIT('h4)
	) name15516 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w16048_
	);
	LUT2 #(
		.INIT('h8)
	) name15517 (
		\u0_w_reg[3][29]/P0001 ,
		_w16043_,
		_w16049_
	);
	LUT2 #(
		.INIT('h8)
	) name15518 (
		_w16048_,
		_w16049_,
		_w16050_
	);
	LUT2 #(
		.INIT('h1)
	) name15519 (
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w16051_
	);
	LUT2 #(
		.INIT('h4)
	) name15520 (
		\u0_w_reg[3][29]/P0001 ,
		_w16051_,
		_w16052_
	);
	LUT2 #(
		.INIT('h8)
	) name15521 (
		_w16048_,
		_w16052_,
		_w16053_
	);
	LUT2 #(
		.INIT('h1)
	) name15522 (
		_w16044_,
		_w16047_,
		_w16054_
	);
	LUT2 #(
		.INIT('h1)
	) name15523 (
		_w16050_,
		_w16053_,
		_w16055_
	);
	LUT2 #(
		.INIT('h8)
	) name15524 (
		_w16054_,
		_w16055_,
		_w16056_
	);
	LUT2 #(
		.INIT('h2)
	) name15525 (
		\u0_w_reg[3][25]/P0001 ,
		_w16056_,
		_w16057_
	);
	LUT2 #(
		.INIT('h8)
	) name15526 (
		\u0_w_reg[3][29]/P0001 ,
		_w16025_,
		_w16058_
	);
	LUT2 #(
		.INIT('h4)
	) name15527 (
		\u0_w_reg[3][29]/P0001 ,
		_w16043_,
		_w16059_
	);
	LUT2 #(
		.INIT('h8)
	) name15528 (
		\u0_w_reg[3][27]/P0001 ,
		_w16059_,
		_w16060_
	);
	LUT2 #(
		.INIT('h1)
	) name15529 (
		_w16058_,
		_w16060_,
		_w16061_
	);
	LUT2 #(
		.INIT('h1)
	) name15530 (
		\u0_w_reg[3][26]/P0001 ,
		_w16061_,
		_w16062_
	);
	LUT2 #(
		.INIT('h8)
	) name15531 (
		_w16011_,
		_w16048_,
		_w16063_
	);
	LUT2 #(
		.INIT('h8)
	) name15532 (
		\u0_w_reg[3][31]/P0001 ,
		_w16063_,
		_w16064_
	);
	LUT2 #(
		.INIT('h4)
	) name15533 (
		\u0_w_reg[3][29]/P0001 ,
		_w16014_,
		_w16065_
	);
	LUT2 #(
		.INIT('h8)
	) name15534 (
		_w16045_,
		_w16051_,
		_w16066_
	);
	LUT2 #(
		.INIT('h1)
	) name15535 (
		_w16065_,
		_w16066_,
		_w16067_
	);
	LUT2 #(
		.INIT('h2)
	) name15536 (
		\u0_w_reg[3][26]/P0001 ,
		_w16067_,
		_w16068_
	);
	LUT2 #(
		.INIT('h1)
	) name15537 (
		_w16013_,
		_w16064_,
		_w16069_
	);
	LUT2 #(
		.INIT('h4)
	) name15538 (
		_w16068_,
		_w16069_,
		_w16070_
	);
	LUT2 #(
		.INIT('h4)
	) name15539 (
		_w16062_,
		_w16070_,
		_w16071_
	);
	LUT2 #(
		.INIT('h1)
	) name15540 (
		\u0_w_reg[3][25]/P0001 ,
		_w16071_,
		_w16072_
	);
	LUT2 #(
		.INIT('h1)
	) name15541 (
		_w16024_,
		_w16028_,
		_w16073_
	);
	LUT2 #(
		.INIT('h1)
	) name15542 (
		_w16035_,
		_w16042_,
		_w16074_
	);
	LUT2 #(
		.INIT('h8)
	) name15543 (
		_w16073_,
		_w16074_,
		_w16075_
	);
	LUT2 #(
		.INIT('h4)
	) name15544 (
		_w16057_,
		_w16075_,
		_w16076_
	);
	LUT2 #(
		.INIT('h4)
	) name15545 (
		_w16072_,
		_w16076_,
		_w16077_
	);
	LUT2 #(
		.INIT('h2)
	) name15546 (
		\u0_w_reg[3][24]/P0001 ,
		_w16077_,
		_w16078_
	);
	LUT2 #(
		.INIT('h2)
	) name15547 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w16079_
	);
	LUT2 #(
		.INIT('h8)
	) name15548 (
		_w16045_,
		_w16079_,
		_w16080_
	);
	LUT2 #(
		.INIT('h4)
	) name15549 (
		\u0_w_reg[3][29]/P0001 ,
		_w16025_,
		_w16081_
	);
	LUT2 #(
		.INIT('h1)
	) name15550 (
		_w16037_,
		_w16059_,
		_w16082_
	);
	LUT2 #(
		.INIT('h4)
	) name15551 (
		_w16081_,
		_w16082_,
		_w16083_
	);
	LUT2 #(
		.INIT('h2)
	) name15552 (
		_w16048_,
		_w16083_,
		_w16084_
	);
	LUT2 #(
		.INIT('h1)
	) name15553 (
		_w16080_,
		_w16084_,
		_w16085_
	);
	LUT2 #(
		.INIT('h2)
	) name15554 (
		\u0_w_reg[3][26]/P0001 ,
		_w16085_,
		_w16086_
	);
	LUT2 #(
		.INIT('h1)
	) name15555 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w16087_
	);
	LUT2 #(
		.INIT('h8)
	) name15556 (
		_w16051_,
		_w16087_,
		_w16088_
	);
	LUT2 #(
		.INIT('h1)
	) name15557 (
		_w16086_,
		_w16088_,
		_w16089_
	);
	LUT2 #(
		.INIT('h1)
	) name15558 (
		\u0_w_reg[3][25]/P0001 ,
		_w16089_,
		_w16090_
	);
	LUT2 #(
		.INIT('h8)
	) name15559 (
		_w16020_,
		_w16079_,
		_w16091_
	);
	LUT2 #(
		.INIT('h4)
	) name15560 (
		\u0_w_reg[3][26]/P0001 ,
		_w16091_,
		_w16092_
	);
	LUT2 #(
		.INIT('h4)
	) name15561 (
		\u0_w_reg[3][28]/P0001 ,
		_w16012_,
		_w16093_
	);
	LUT2 #(
		.INIT('h1)
	) name15562 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w16094_
	);
	LUT2 #(
		.INIT('h8)
	) name15563 (
		_w16093_,
		_w16094_,
		_w16095_
	);
	LUT2 #(
		.INIT('h1)
	) name15564 (
		_w16092_,
		_w16095_,
		_w16096_
	);
	LUT2 #(
		.INIT('h2)
	) name15565 (
		\u0_w_reg[3][25]/P0001 ,
		_w16096_,
		_w16097_
	);
	LUT2 #(
		.INIT('h8)
	) name15566 (
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w16098_
	);
	LUT2 #(
		.INIT('h4)
	) name15567 (
		\u0_w_reg[3][29]/P0001 ,
		_w16098_,
		_w16099_
	);
	LUT2 #(
		.INIT('h4)
	) name15568 (
		\u0_w_reg[3][27]/P0001 ,
		_w16099_,
		_w16100_
	);
	LUT2 #(
		.INIT('h4)
	) name15569 (
		\u0_w_reg[3][26]/P0001 ,
		_w16100_,
		_w16101_
	);
	LUT2 #(
		.INIT('h8)
	) name15570 (
		_w16017_,
		_w16045_,
		_w16102_
	);
	LUT2 #(
		.INIT('h2)
	) name15571 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w16103_
	);
	LUT2 #(
		.INIT('h8)
	) name15572 (
		_w16102_,
		_w16103_,
		_w16104_
	);
	LUT2 #(
		.INIT('h2)
	) name15573 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w16105_
	);
	LUT2 #(
		.INIT('h8)
	) name15574 (
		_w16036_,
		_w16105_,
		_w16106_
	);
	LUT2 #(
		.INIT('h8)
	) name15575 (
		\u0_w_reg[3][25]/P0001 ,
		_w16011_,
		_w16107_
	);
	LUT2 #(
		.INIT('h8)
	) name15576 (
		_w16106_,
		_w16107_,
		_w16108_
	);
	LUT2 #(
		.INIT('h1)
	) name15577 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		_w16109_
	);
	LUT2 #(
		.INIT('h8)
	) name15578 (
		_w16011_,
		_w16045_,
		_w16110_
	);
	LUT2 #(
		.INIT('h4)
	) name15579 (
		\u0_w_reg[3][31]/P0001 ,
		_w16110_,
		_w16111_
	);
	LUT2 #(
		.INIT('h8)
	) name15580 (
		\u0_w_reg[3][29]/P0001 ,
		_w16087_,
		_w16112_
	);
	LUT2 #(
		.INIT('h8)
	) name15581 (
		\u0_w_reg[3][31]/P0001 ,
		_w16112_,
		_w16113_
	);
	LUT2 #(
		.INIT('h1)
	) name15582 (
		_w16021_,
		_w16111_,
		_w16114_
	);
	LUT2 #(
		.INIT('h4)
	) name15583 (
		_w16113_,
		_w16114_,
		_w16115_
	);
	LUT2 #(
		.INIT('h2)
	) name15584 (
		_w16109_,
		_w16115_,
		_w16116_
	);
	LUT2 #(
		.INIT('h4)
	) name15585 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w16117_
	);
	LUT2 #(
		.INIT('h8)
	) name15586 (
		_w16026_,
		_w16051_,
		_w16118_
	);
	LUT2 #(
		.INIT('h8)
	) name15587 (
		_w16117_,
		_w16118_,
		_w16119_
	);
	LUT2 #(
		.INIT('h8)
	) name15588 (
		_w16039_,
		_w16094_,
		_w16120_
	);
	LUT2 #(
		.INIT('h4)
	) name15589 (
		\u0_w_reg[3][28]/P0001 ,
		_w16094_,
		_w16121_
	);
	LUT2 #(
		.INIT('h8)
	) name15590 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w16122_
	);
	LUT2 #(
		.INIT('h8)
	) name15591 (
		_w16121_,
		_w16122_,
		_w16123_
	);
	LUT2 #(
		.INIT('h8)
	) name15592 (
		_w16043_,
		_w16048_,
		_w16124_
	);
	LUT2 #(
		.INIT('h4)
	) name15593 (
		\u0_w_reg[3][27]/P0001 ,
		_w16051_,
		_w16125_
	);
	LUT2 #(
		.INIT('h8)
	) name15594 (
		\u0_w_reg[3][26]/P0001 ,
		_w16125_,
		_w16126_
	);
	LUT2 #(
		.INIT('h1)
	) name15595 (
		_w16124_,
		_w16126_,
		_w16127_
	);
	LUT2 #(
		.INIT('h1)
	) name15596 (
		\u0_w_reg[3][29]/P0001 ,
		_w16127_,
		_w16128_
	);
	LUT2 #(
		.INIT('h4)
	) name15597 (
		\u0_w_reg[3][27]/P0001 ,
		_w16037_,
		_w16129_
	);
	LUT2 #(
		.INIT('h4)
	) name15598 (
		\u0_w_reg[3][28]/P0001 ,
		_w16129_,
		_w16130_
	);
	LUT2 #(
		.INIT('h1)
	) name15599 (
		\u0_w_reg[3][25]/P0001 ,
		_w16123_,
		_w16131_
	);
	LUT2 #(
		.INIT('h4)
	) name15600 (
		_w16130_,
		_w16131_,
		_w16132_
	);
	LUT2 #(
		.INIT('h4)
	) name15601 (
		_w16128_,
		_w16132_,
		_w16133_
	);
	LUT2 #(
		.INIT('h8)
	) name15602 (
		_w16048_,
		_w16079_,
		_w16134_
	);
	LUT2 #(
		.INIT('h1)
	) name15603 (
		_w16043_,
		_w16087_,
		_w16135_
	);
	LUT2 #(
		.INIT('h1)
	) name15604 (
		\u0_w_reg[3][27]/P0001 ,
		_w16025_,
		_w16136_
	);
	LUT2 #(
		.INIT('h1)
	) name15605 (
		_w16135_,
		_w16136_,
		_w16137_
	);
	LUT2 #(
		.INIT('h1)
	) name15606 (
		_w16134_,
		_w16137_,
		_w16138_
	);
	LUT2 #(
		.INIT('h1)
	) name15607 (
		\u0_w_reg[3][26]/P0001 ,
		_w16138_,
		_w16139_
	);
	LUT2 #(
		.INIT('h4)
	) name15608 (
		\u0_w_reg[3][27]/P0001 ,
		_w16025_,
		_w16140_
	);
	LUT2 #(
		.INIT('h8)
	) name15609 (
		_w16026_,
		_w16140_,
		_w16141_
	);
	LUT2 #(
		.INIT('h8)
	) name15610 (
		\u0_w_reg[3][26]/P0001 ,
		_w16011_,
		_w16142_
	);
	LUT2 #(
		.INIT('h8)
	) name15611 (
		_w16105_,
		_w16142_,
		_w16143_
	);
	LUT2 #(
		.INIT('h8)
	) name15612 (
		_w16012_,
		_w16094_,
		_w16144_
	);
	LUT2 #(
		.INIT('h8)
	) name15613 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w16145_
	);
	LUT2 #(
		.INIT('h8)
	) name15614 (
		\u0_w_reg[3][27]/P0001 ,
		_w16145_,
		_w16146_
	);
	LUT2 #(
		.INIT('h1)
	) name15615 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w16147_
	);
	LUT2 #(
		.INIT('h2)
	) name15616 (
		_w16146_,
		_w16147_,
		_w16148_
	);
	LUT2 #(
		.INIT('h2)
	) name15617 (
		\u0_w_reg[3][25]/P0001 ,
		_w16100_,
		_w16149_
	);
	LUT2 #(
		.INIT('h8)
	) name15618 (
		_w16026_,
		_w16043_,
		_w16150_
	);
	LUT2 #(
		.INIT('h1)
	) name15619 (
		_w16144_,
		_w16150_,
		_w16151_
	);
	LUT2 #(
		.INIT('h4)
	) name15620 (
		_w16141_,
		_w16151_,
		_w16152_
	);
	LUT2 #(
		.INIT('h1)
	) name15621 (
		_w16143_,
		_w16148_,
		_w16153_
	);
	LUT2 #(
		.INIT('h8)
	) name15622 (
		_w16152_,
		_w16153_,
		_w16154_
	);
	LUT2 #(
		.INIT('h8)
	) name15623 (
		_w16149_,
		_w16154_,
		_w16155_
	);
	LUT2 #(
		.INIT('h4)
	) name15624 (
		_w16139_,
		_w16155_,
		_w16156_
	);
	LUT2 #(
		.INIT('h1)
	) name15625 (
		_w16133_,
		_w16156_,
		_w16157_
	);
	LUT2 #(
		.INIT('h8)
	) name15626 (
		\u0_w_reg[3][31]/P0001 ,
		_w16045_,
		_w16158_
	);
	LUT2 #(
		.INIT('h8)
	) name15627 (
		\u0_w_reg[3][29]/P0001 ,
		_w16158_,
		_w16159_
	);
	LUT2 #(
		.INIT('h8)
	) name15628 (
		\u0_w_reg[3][28]/P0001 ,
		_w16019_,
		_w16160_
	);
	LUT2 #(
		.INIT('h4)
	) name15629 (
		\u0_w_reg[3][31]/P0001 ,
		_w16160_,
		_w16161_
	);
	LUT2 #(
		.INIT('h4)
	) name15630 (
		\u0_w_reg[3][27]/P0001 ,
		_w16161_,
		_w16162_
	);
	LUT2 #(
		.INIT('h4)
	) name15631 (
		\u0_w_reg[3][28]/P0001 ,
		_w16051_,
		_w16163_
	);
	LUT2 #(
		.INIT('h2)
	) name15632 (
		\u0_w_reg[3][26]/P0001 ,
		_w16163_,
		_w16164_
	);
	LUT2 #(
		.INIT('h4)
	) name15633 (
		\u0_w_reg[3][29]/P0001 ,
		_w16093_,
		_w16165_
	);
	LUT2 #(
		.INIT('h4)
	) name15634 (
		_w16159_,
		_w16164_,
		_w16166_
	);
	LUT2 #(
		.INIT('h4)
	) name15635 (
		_w16165_,
		_w16166_,
		_w16167_
	);
	LUT2 #(
		.INIT('h4)
	) name15636 (
		_w16162_,
		_w16167_,
		_w16168_
	);
	LUT2 #(
		.INIT('h4)
	) name15637 (
		\u0_w_reg[3][29]/P0001 ,
		_w16105_,
		_w16169_
	);
	LUT2 #(
		.INIT('h8)
	) name15638 (
		\u0_w_reg[3][27]/P0001 ,
		_w16169_,
		_w16170_
	);
	LUT2 #(
		.INIT('h4)
	) name15639 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w16171_
	);
	LUT2 #(
		.INIT('h8)
	) name15640 (
		_w16014_,
		_w16171_,
		_w16172_
	);
	LUT2 #(
		.INIT('h1)
	) name15641 (
		_w16170_,
		_w16172_,
		_w16173_
	);
	LUT2 #(
		.INIT('h1)
	) name15642 (
		\u0_w_reg[3][26]/P0001 ,
		_w16091_,
		_w16174_
	);
	LUT2 #(
		.INIT('h8)
	) name15643 (
		_w16173_,
		_w16174_,
		_w16175_
	);
	LUT2 #(
		.INIT('h1)
	) name15644 (
		_w16168_,
		_w16175_,
		_w16176_
	);
	LUT2 #(
		.INIT('h1)
	) name15645 (
		_w16120_,
		_w16176_,
		_w16177_
	);
	LUT2 #(
		.INIT('h4)
	) name15646 (
		_w16157_,
		_w16177_,
		_w16178_
	);
	LUT2 #(
		.INIT('h1)
	) name15647 (
		\u0_w_reg[3][24]/P0001 ,
		_w16178_,
		_w16179_
	);
	LUT2 #(
		.INIT('h1)
	) name15648 (
		_w16104_,
		_w16108_,
		_w16180_
	);
	LUT2 #(
		.INIT('h4)
	) name15649 (
		_w16119_,
		_w16180_,
		_w16181_
	);
	LUT2 #(
		.INIT('h4)
	) name15650 (
		_w16101_,
		_w16181_,
		_w16182_
	);
	LUT2 #(
		.INIT('h4)
	) name15651 (
		_w16097_,
		_w16182_,
		_w16183_
	);
	LUT2 #(
		.INIT('h4)
	) name15652 (
		_w16116_,
		_w16183_,
		_w16184_
	);
	LUT2 #(
		.INIT('h4)
	) name15653 (
		_w16090_,
		_w16184_,
		_w16185_
	);
	LUT2 #(
		.INIT('h4)
	) name15654 (
		_w16078_,
		_w16185_,
		_w16186_
	);
	LUT2 #(
		.INIT('h4)
	) name15655 (
		_w16179_,
		_w16186_,
		_w16187_
	);
	LUT2 #(
		.INIT('h2)
	) name15656 (
		\u0_w_reg[0][5]/P0001 ,
		_w16187_,
		_w16188_
	);
	LUT2 #(
		.INIT('h4)
	) name15657 (
		\u0_w_reg[0][5]/P0001 ,
		_w16187_,
		_w16189_
	);
	LUT2 #(
		.INIT('h1)
	) name15658 (
		_w16188_,
		_w16189_,
		_w16190_
	);
	LUT2 #(
		.INIT('h2)
	) name15659 (
		\u0_w_reg[1][5]/P0001 ,
		\u0_w_reg[2][5]/P0001 ,
		_w16191_
	);
	LUT2 #(
		.INIT('h4)
	) name15660 (
		\u0_w_reg[1][5]/P0001 ,
		\u0_w_reg[2][5]/P0001 ,
		_w16192_
	);
	LUT2 #(
		.INIT('h1)
	) name15661 (
		_w16191_,
		_w16192_,
		_w16193_
	);
	LUT2 #(
		.INIT('h8)
	) name15662 (
		_w16190_,
		_w16193_,
		_w16194_
	);
	LUT2 #(
		.INIT('h1)
	) name15663 (
		_w16190_,
		_w16193_,
		_w16195_
	);
	LUT2 #(
		.INIT('h1)
	) name15664 (
		_w16194_,
		_w16195_,
		_w16196_
	);
	LUT2 #(
		.INIT('h4)
	) name15665 (
		ld_pad,
		_w16196_,
		_w16197_
	);
	LUT2 #(
		.INIT('h1)
	) name15666 (
		_w16010_,
		_w16197_,
		_w16198_
	);
	LUT2 #(
		.INIT('h2)
	) name15667 (
		\u0_w_reg[0][10]/P0001 ,
		_w15068_,
		_w16199_
	);
	LUT2 #(
		.INIT('h4)
	) name15668 (
		\u0_w_reg[0][10]/P0001 ,
		_w15068_,
		_w16200_
	);
	LUT2 #(
		.INIT('h1)
	) name15669 (
		_w16199_,
		_w16200_,
		_w16201_
	);
	LUT2 #(
		.INIT('h8)
	) name15670 (
		_w13752_,
		_w16201_,
		_w16202_
	);
	LUT2 #(
		.INIT('h1)
	) name15671 (
		_w13752_,
		_w16201_,
		_w16203_
	);
	LUT2 #(
		.INIT('h1)
	) name15672 (
		_w16202_,
		_w16203_,
		_w16204_
	);
	LUT2 #(
		.INIT('h8)
	) name15673 (
		_w13835_,
		_w14804_,
		_w16205_
	);
	LUT2 #(
		.INIT('h1)
	) name15674 (
		_w13835_,
		_w14804_,
		_w16206_
	);
	LUT2 #(
		.INIT('h1)
	) name15675 (
		_w16205_,
		_w16206_,
		_w16207_
	);
	LUT2 #(
		.INIT('h1)
	) name15676 (
		_w16204_,
		_w16207_,
		_w16208_
	);
	LUT2 #(
		.INIT('h8)
	) name15677 (
		_w16204_,
		_w16207_,
		_w16209_
	);
	LUT2 #(
		.INIT('h1)
	) name15678 (
		\ld_r_reg/P0001 ,
		_w16208_,
		_w16210_
	);
	LUT2 #(
		.INIT('h4)
	) name15679 (
		_w16209_,
		_w16210_,
		_w16211_
	);
	LUT2 #(
		.INIT('h2)
	) name15680 (
		\text_in_r_reg[106]/P0001 ,
		\u0_w_reg[0][10]/P0001 ,
		_w16212_
	);
	LUT2 #(
		.INIT('h4)
	) name15681 (
		\text_in_r_reg[106]/P0001 ,
		\u0_w_reg[0][10]/P0001 ,
		_w16213_
	);
	LUT2 #(
		.INIT('h2)
	) name15682 (
		\ld_r_reg/P0001 ,
		_w16212_,
		_w16214_
	);
	LUT2 #(
		.INIT('h4)
	) name15683 (
		_w16213_,
		_w16214_,
		_w16215_
	);
	LUT2 #(
		.INIT('h1)
	) name15684 (
		_w16211_,
		_w16215_,
		_w16216_
	);
	LUT2 #(
		.INIT('h8)
	) name15685 (
		\u0_w_reg[3][19]/P0001 ,
		_w15531_,
		_w16217_
	);
	LUT2 #(
		.INIT('h1)
	) name15686 (
		_w15516_,
		_w15543_,
		_w16218_
	);
	LUT2 #(
		.INIT('h4)
	) name15687 (
		_w16217_,
		_w16218_,
		_w16219_
	);
	LUT2 #(
		.INIT('h2)
	) name15688 (
		\u0_w_reg[3][18]/P0001 ,
		_w16219_,
		_w16220_
	);
	LUT2 #(
		.INIT('h8)
	) name15689 (
		_w15529_,
		_w15638_,
		_w16221_
	);
	LUT2 #(
		.INIT('h8)
	) name15690 (
		_w15562_,
		_w15601_,
		_w16222_
	);
	LUT2 #(
		.INIT('h1)
	) name15691 (
		_w15580_,
		_w15637_,
		_w16223_
	);
	LUT2 #(
		.INIT('h4)
	) name15692 (
		_w15661_,
		_w16223_,
		_w16224_
	);
	LUT2 #(
		.INIT('h1)
	) name15693 (
		_w16221_,
		_w16222_,
		_w16225_
	);
	LUT2 #(
		.INIT('h8)
	) name15694 (
		_w16224_,
		_w16225_,
		_w16226_
	);
	LUT2 #(
		.INIT('h4)
	) name15695 (
		_w16220_,
		_w16226_,
		_w16227_
	);
	LUT2 #(
		.INIT('h1)
	) name15696 (
		\u0_w_reg[3][17]/P0001 ,
		_w16227_,
		_w16228_
	);
	LUT2 #(
		.INIT('h8)
	) name15697 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w16229_
	);
	LUT2 #(
		.INIT('h8)
	) name15698 (
		_w15601_,
		_w16229_,
		_w16230_
	);
	LUT2 #(
		.INIT('h1)
	) name15699 (
		_w15628_,
		_w16230_,
		_w16231_
	);
	LUT2 #(
		.INIT('h4)
	) name15700 (
		\u0_w_reg[3][18]/P0001 ,
		_w15557_,
		_w16232_
	);
	LUT2 #(
		.INIT('h8)
	) name15701 (
		_w15503_,
		_w15648_,
		_w16233_
	);
	LUT2 #(
		.INIT('h1)
	) name15702 (
		_w15527_,
		_w16233_,
		_w16234_
	);
	LUT2 #(
		.INIT('h8)
	) name15703 (
		_w16231_,
		_w16234_,
		_w16235_
	);
	LUT2 #(
		.INIT('h4)
	) name15704 (
		_w16232_,
		_w16235_,
		_w16236_
	);
	LUT2 #(
		.INIT('h2)
	) name15705 (
		\u0_w_reg[3][17]/P0001 ,
		_w16236_,
		_w16237_
	);
	LUT2 #(
		.INIT('h8)
	) name15706 (
		_w15503_,
		_w15505_,
		_w16238_
	);
	LUT2 #(
		.INIT('h4)
	) name15707 (
		\u0_w_reg[3][18]/P0001 ,
		_w15527_,
		_w16239_
	);
	LUT2 #(
		.INIT('h4)
	) name15708 (
		\u0_w_reg[3][22]/P0001 ,
		_w16239_,
		_w16240_
	);
	LUT2 #(
		.INIT('h8)
	) name15709 (
		_w15506_,
		_w15601_,
		_w16241_
	);
	LUT2 #(
		.INIT('h8)
	) name15710 (
		_w15526_,
		_w16229_,
		_w16242_
	);
	LUT2 #(
		.INIT('h1)
	) name15711 (
		_w16241_,
		_w16242_,
		_w16243_
	);
	LUT2 #(
		.INIT('h1)
	) name15712 (
		\u0_w_reg[3][18]/P0001 ,
		_w16243_,
		_w16244_
	);
	LUT2 #(
		.INIT('h4)
	) name15713 (
		_w15537_,
		_w15559_,
		_w16245_
	);
	LUT2 #(
		.INIT('h1)
	) name15714 (
		_w15602_,
		_w16245_,
		_w16246_
	);
	LUT2 #(
		.INIT('h2)
	) name15715 (
		\u0_w_reg[3][17]/P0001 ,
		_w16246_,
		_w16247_
	);
	LUT2 #(
		.INIT('h8)
	) name15716 (
		\u0_w_reg[3][23]/P0001 ,
		_w15521_,
		_w16248_
	);
	LUT2 #(
		.INIT('h4)
	) name15717 (
		\u0_w_reg[3][22]/P0001 ,
		_w16248_,
		_w16249_
	);
	LUT2 #(
		.INIT('h1)
	) name15718 (
		_w15603_,
		_w15618_,
		_w16250_
	);
	LUT2 #(
		.INIT('h4)
	) name15719 (
		_w16249_,
		_w16250_,
		_w16251_
	);
	LUT2 #(
		.INIT('h4)
	) name15720 (
		_w16247_,
		_w16251_,
		_w16252_
	);
	LUT2 #(
		.INIT('h2)
	) name15721 (
		\u0_w_reg[3][18]/P0001 ,
		_w16252_,
		_w16253_
	);
	LUT2 #(
		.INIT('h1)
	) name15722 (
		_w16238_,
		_w16240_,
		_w16254_
	);
	LUT2 #(
		.INIT('h4)
	) name15723 (
		_w16244_,
		_w16254_,
		_w16255_
	);
	LUT2 #(
		.INIT('h4)
	) name15724 (
		_w16237_,
		_w16255_,
		_w16256_
	);
	LUT2 #(
		.INIT('h4)
	) name15725 (
		_w16228_,
		_w16256_,
		_w16257_
	);
	LUT2 #(
		.INIT('h4)
	) name15726 (
		_w16253_,
		_w16257_,
		_w16258_
	);
	LUT2 #(
		.INIT('h2)
	) name15727 (
		\u0_w_reg[3][16]/P0001 ,
		_w16258_,
		_w16259_
	);
	LUT2 #(
		.INIT('h2)
	) name15728 (
		\u0_w_reg[3][18]/P0001 ,
		_w16231_,
		_w16260_
	);
	LUT2 #(
		.INIT('h8)
	) name15729 (
		\u0_w_reg[3][20]/P0001 ,
		_w15549_,
		_w16261_
	);
	LUT2 #(
		.INIT('h4)
	) name15730 (
		\u0_w_reg[3][20]/P0001 ,
		_w15503_,
		_w16262_
	);
	LUT2 #(
		.INIT('h1)
	) name15731 (
		_w16261_,
		_w16262_,
		_w16263_
	);
	LUT2 #(
		.INIT('h4)
	) name15732 (
		_w15583_,
		_w16263_,
		_w16264_
	);
	LUT2 #(
		.INIT('h2)
	) name15733 (
		_w15648_,
		_w16264_,
		_w16265_
	);
	LUT2 #(
		.INIT('h4)
	) name15734 (
		\u0_w_reg[3][20]/P0001 ,
		_w15608_,
		_w16266_
	);
	LUT2 #(
		.INIT('h8)
	) name15735 (
		_w15512_,
		_w16266_,
		_w16267_
	);
	LUT2 #(
		.INIT('h4)
	) name15736 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w16268_
	);
	LUT2 #(
		.INIT('h8)
	) name15737 (
		_w15549_,
		_w16268_,
		_w16269_
	);
	LUT2 #(
		.INIT('h8)
	) name15738 (
		_w15529_,
		_w16269_,
		_w16270_
	);
	LUT2 #(
		.INIT('h1)
	) name15739 (
		_w16267_,
		_w16270_,
		_w16271_
	);
	LUT2 #(
		.INIT('h4)
	) name15740 (
		_w16260_,
		_w16271_,
		_w16272_
	);
	LUT2 #(
		.INIT('h4)
	) name15741 (
		_w16265_,
		_w16272_,
		_w16273_
	);
	LUT2 #(
		.INIT('h2)
	) name15742 (
		\u0_w_reg[3][17]/P0001 ,
		_w16273_,
		_w16274_
	);
	LUT2 #(
		.INIT('h8)
	) name15743 (
		_w15603_,
		_w15608_,
		_w16275_
	);
	LUT2 #(
		.INIT('h8)
	) name15744 (
		\u0_w_reg[3][18]/P0001 ,
		_w16230_,
		_w16276_
	);
	LUT2 #(
		.INIT('h4)
	) name15745 (
		\u0_w_reg[3][17]/P0001 ,
		_w15529_,
		_w16277_
	);
	LUT2 #(
		.INIT('h8)
	) name15746 (
		_w15590_,
		_w16277_,
		_w16278_
	);
	LUT2 #(
		.INIT('h1)
	) name15747 (
		_w16276_,
		_w16278_,
		_w16279_
	);
	LUT2 #(
		.INIT('h1)
	) name15748 (
		\u0_w_reg[3][20]/P0001 ,
		_w16279_,
		_w16280_
	);
	LUT2 #(
		.INIT('h4)
	) name15749 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		_w16281_
	);
	LUT2 #(
		.INIT('h4)
	) name15750 (
		\u0_w_reg[3][19]/P0001 ,
		_w16281_,
		_w16282_
	);
	LUT2 #(
		.INIT('h4)
	) name15751 (
		\u0_w_reg[3][23]/P0001 ,
		_w15519_,
		_w16283_
	);
	LUT2 #(
		.INIT('h8)
	) name15752 (
		_w15549_,
		_w15551_,
		_w16284_
	);
	LUT2 #(
		.INIT('h1)
	) name15753 (
		_w16283_,
		_w16284_,
		_w16285_
	);
	LUT2 #(
		.INIT('h2)
	) name15754 (
		_w16282_,
		_w16285_,
		_w16286_
	);
	LUT2 #(
		.INIT('h8)
	) name15755 (
		_w15503_,
		_w15521_,
		_w16287_
	);
	LUT2 #(
		.INIT('h4)
	) name15756 (
		\u0_w_reg[3][21]/P0001 ,
		_w16287_,
		_w16288_
	);
	LUT2 #(
		.INIT('h8)
	) name15757 (
		\u0_w_reg[3][20]/P0001 ,
		_w16242_,
		_w16289_
	);
	LUT2 #(
		.INIT('h4)
	) name15758 (
		\u0_w_reg[3][18]/P0001 ,
		_w15583_,
		_w16290_
	);
	LUT2 #(
		.INIT('h2)
	) name15759 (
		\u0_w_reg[3][17]/P0001 ,
		_w15607_,
		_w16291_
	);
	LUT2 #(
		.INIT('h1)
	) name15760 (
		_w16217_,
		_w16289_,
		_w16292_
	);
	LUT2 #(
		.INIT('h8)
	) name15761 (
		_w16291_,
		_w16292_,
		_w16293_
	);
	LUT2 #(
		.INIT('h4)
	) name15762 (
		_w16290_,
		_w16293_,
		_w16294_
	);
	LUT2 #(
		.INIT('h8)
	) name15763 (
		\u0_w_reg[3][23]/P0001 ,
		_w15511_,
		_w16295_
	);
	LUT2 #(
		.INIT('h4)
	) name15764 (
		_w15549_,
		_w16295_,
		_w16296_
	);
	LUT2 #(
		.INIT('h2)
	) name15765 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w16297_
	);
	LUT2 #(
		.INIT('h1)
	) name15766 (
		_w15549_,
		_w16297_,
		_w16298_
	);
	LUT2 #(
		.INIT('h2)
	) name15767 (
		_w15551_,
		_w16298_,
		_w16299_
	);
	LUT2 #(
		.INIT('h8)
	) name15768 (
		\u0_w_reg[3][19]/P0001 ,
		_w15629_,
		_w16300_
	);
	LUT2 #(
		.INIT('h1)
	) name15769 (
		\u0_w_reg[3][17]/P0001 ,
		_w16241_,
		_w16301_
	);
	LUT2 #(
		.INIT('h4)
	) name15770 (
		_w16296_,
		_w16301_,
		_w16302_
	);
	LUT2 #(
		.INIT('h4)
	) name15771 (
		_w16299_,
		_w16302_,
		_w16303_
	);
	LUT2 #(
		.INIT('h4)
	) name15772 (
		_w16300_,
		_w16303_,
		_w16304_
	);
	LUT2 #(
		.INIT('h1)
	) name15773 (
		_w16294_,
		_w16304_,
		_w16305_
	);
	LUT2 #(
		.INIT('h1)
	) name15774 (
		_w15528_,
		_w16287_,
		_w16306_
	);
	LUT2 #(
		.INIT('h4)
	) name15775 (
		\u0_w_reg[3][18]/P0001 ,
		_w16306_,
		_w16307_
	);
	LUT2 #(
		.INIT('h8)
	) name15776 (
		\u0_w_reg[3][19]/P0001 ,
		_w15614_,
		_w16308_
	);
	LUT2 #(
		.INIT('h8)
	) name15777 (
		\u0_w_reg[3][22]/P0001 ,
		_w15525_,
		_w16309_
	);
	LUT2 #(
		.INIT('h8)
	) name15778 (
		_w15542_,
		_w16309_,
		_w16310_
	);
	LUT2 #(
		.INIT('h1)
	) name15779 (
		_w15614_,
		_w16310_,
		_w16311_
	);
	LUT2 #(
		.INIT('h2)
	) name15780 (
		\u0_w_reg[3][17]/P0001 ,
		_w16311_,
		_w16312_
	);
	LUT2 #(
		.INIT('h8)
	) name15781 (
		_w15526_,
		_w15539_,
		_w16313_
	);
	LUT2 #(
		.INIT('h2)
	) name15782 (
		\u0_w_reg[3][18]/P0001 ,
		_w16313_,
		_w16314_
	);
	LUT2 #(
		.INIT('h4)
	) name15783 (
		_w16308_,
		_w16314_,
		_w16315_
	);
	LUT2 #(
		.INIT('h4)
	) name15784 (
		_w16312_,
		_w16315_,
		_w16316_
	);
	LUT2 #(
		.INIT('h1)
	) name15785 (
		_w16307_,
		_w16316_,
		_w16317_
	);
	LUT2 #(
		.INIT('h4)
	) name15786 (
		\u0_w_reg[3][21]/P0001 ,
		_w15574_,
		_w16318_
	);
	LUT2 #(
		.INIT('h1)
	) name15787 (
		_w16305_,
		_w16318_,
		_w16319_
	);
	LUT2 #(
		.INIT('h4)
	) name15788 (
		_w16317_,
		_w16319_,
		_w16320_
	);
	LUT2 #(
		.INIT('h1)
	) name15789 (
		\u0_w_reg[3][16]/P0001 ,
		_w16320_,
		_w16321_
	);
	LUT2 #(
		.INIT('h1)
	) name15790 (
		_w16275_,
		_w16288_,
		_w16322_
	);
	LUT2 #(
		.INIT('h4)
	) name15791 (
		_w16280_,
		_w16322_,
		_w16323_
	);
	LUT2 #(
		.INIT('h4)
	) name15792 (
		_w16286_,
		_w16323_,
		_w16324_
	);
	LUT2 #(
		.INIT('h4)
	) name15793 (
		_w16274_,
		_w16324_,
		_w16325_
	);
	LUT2 #(
		.INIT('h4)
	) name15794 (
		_w16259_,
		_w16325_,
		_w16326_
	);
	LUT2 #(
		.INIT('h4)
	) name15795 (
		_w16321_,
		_w16326_,
		_w16327_
	);
	LUT2 #(
		.INIT('h2)
	) name15796 (
		\u0_r0_out_reg[27]/P0001 ,
		\u0_w_reg[0][27]/P0001 ,
		_w16328_
	);
	LUT2 #(
		.INIT('h4)
	) name15797 (
		\u0_r0_out_reg[27]/P0001 ,
		\u0_w_reg[0][27]/P0001 ,
		_w16329_
	);
	LUT2 #(
		.INIT('h1)
	) name15798 (
		_w16328_,
		_w16329_,
		_w16330_
	);
	LUT2 #(
		.INIT('h1)
	) name15799 (
		_w16327_,
		_w16330_,
		_w16331_
	);
	LUT2 #(
		.INIT('h8)
	) name15800 (
		_w16327_,
		_w16330_,
		_w16332_
	);
	LUT2 #(
		.INIT('h1)
	) name15801 (
		ld_pad,
		_w16331_,
		_w16333_
	);
	LUT2 #(
		.INIT('h4)
	) name15802 (
		_w16332_,
		_w16333_,
		_w16334_
	);
	LUT2 #(
		.INIT('h8)
	) name15803 (
		\key[123]_pad ,
		ld_pad,
		_w16335_
	);
	LUT2 #(
		.INIT('h1)
	) name15804 (
		_w16334_,
		_w16335_,
		_w16336_
	);
	LUT2 #(
		.INIT('h4)
	) name15805 (
		\key[91]_pad ,
		ld_pad,
		_w16337_
	);
	LUT2 #(
		.INIT('h2)
	) name15806 (
		\u0_w_reg[1][27]/P0001 ,
		_w16330_,
		_w16338_
	);
	LUT2 #(
		.INIT('h4)
	) name15807 (
		\u0_w_reg[1][27]/P0001 ,
		_w16330_,
		_w16339_
	);
	LUT2 #(
		.INIT('h1)
	) name15808 (
		_w16338_,
		_w16339_,
		_w16340_
	);
	LUT2 #(
		.INIT('h8)
	) name15809 (
		_w16327_,
		_w16340_,
		_w16341_
	);
	LUT2 #(
		.INIT('h1)
	) name15810 (
		_w16327_,
		_w16340_,
		_w16342_
	);
	LUT2 #(
		.INIT('h1)
	) name15811 (
		_w16341_,
		_w16342_,
		_w16343_
	);
	LUT2 #(
		.INIT('h4)
	) name15812 (
		ld_pad,
		_w16343_,
		_w16344_
	);
	LUT2 #(
		.INIT('h1)
	) name15813 (
		_w16337_,
		_w16344_,
		_w16345_
	);
	LUT2 #(
		.INIT('h4)
	) name15814 (
		\key[59]_pad ,
		ld_pad,
		_w16346_
	);
	LUT2 #(
		.INIT('h8)
	) name15815 (
		\u0_w_reg[2][27]/P0001 ,
		_w16343_,
		_w16347_
	);
	LUT2 #(
		.INIT('h1)
	) name15816 (
		\u0_w_reg[2][27]/P0001 ,
		_w16343_,
		_w16348_
	);
	LUT2 #(
		.INIT('h1)
	) name15817 (
		_w16347_,
		_w16348_,
		_w16349_
	);
	LUT2 #(
		.INIT('h4)
	) name15818 (
		ld_pad,
		_w16349_,
		_w16350_
	);
	LUT2 #(
		.INIT('h1)
	) name15819 (
		_w16346_,
		_w16350_,
		_w16351_
	);
	LUT2 #(
		.INIT('h4)
	) name15820 (
		\u0_w_reg[3][27]/P0001 ,
		_w16349_,
		_w16352_
	);
	LUT2 #(
		.INIT('h2)
	) name15821 (
		\u0_w_reg[3][27]/P0001 ,
		_w16349_,
		_w16353_
	);
	LUT2 #(
		.INIT('h1)
	) name15822 (
		ld_pad,
		_w16352_,
		_w16354_
	);
	LUT2 #(
		.INIT('h4)
	) name15823 (
		_w16353_,
		_w16354_,
		_w16355_
	);
	LUT2 #(
		.INIT('h8)
	) name15824 (
		\key[27]_pad ,
		ld_pad,
		_w16356_
	);
	LUT2 #(
		.INIT('h1)
	) name15825 (
		_w16355_,
		_w16356_,
		_w16357_
	);
	LUT2 #(
		.INIT('h4)
	) name15826 (
		\key[35]_pad ,
		ld_pad,
		_w16358_
	);
	LUT2 #(
		.INIT('h4)
	) name15827 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w16359_
	);
	LUT2 #(
		.INIT('h4)
	) name15828 (
		\u0_w_reg[3][27]/P0001 ,
		_w16359_,
		_w16360_
	);
	LUT2 #(
		.INIT('h4)
	) name15829 (
		\u0_w_reg[3][29]/P0001 ,
		_w16360_,
		_w16361_
	);
	LUT2 #(
		.INIT('h8)
	) name15830 (
		\u0_w_reg[3][30]/P0001 ,
		_w16146_,
		_w16362_
	);
	LUT2 #(
		.INIT('h1)
	) name15831 (
		_w16050_,
		_w16362_,
		_w16363_
	);
	LUT2 #(
		.INIT('h1)
	) name15832 (
		\u0_w_reg[3][26]/P0001 ,
		_w16361_,
		_w16364_
	);
	LUT2 #(
		.INIT('h8)
	) name15833 (
		_w16363_,
		_w16364_,
		_w16365_
	);
	LUT2 #(
		.INIT('h8)
	) name15834 (
		_w16020_,
		_w16094_,
		_w16366_
	);
	LUT2 #(
		.INIT('h4)
	) name15835 (
		\u0_w_reg[3][30]/P0001 ,
		_w16158_,
		_w16367_
	);
	LUT2 #(
		.INIT('h2)
	) name15836 (
		\u0_w_reg[3][26]/P0001 ,
		_w16366_,
		_w16368_
	);
	LUT2 #(
		.INIT('h4)
	) name15837 (
		_w16161_,
		_w16368_,
		_w16369_
	);
	LUT2 #(
		.INIT('h4)
	) name15838 (
		_w16367_,
		_w16369_,
		_w16370_
	);
	LUT2 #(
		.INIT('h1)
	) name15839 (
		_w16365_,
		_w16370_,
		_w16371_
	);
	LUT2 #(
		.INIT('h4)
	) name15840 (
		_w16018_,
		_w16061_,
		_w16372_
	);
	LUT2 #(
		.INIT('h2)
	) name15841 (
		\u0_w_reg[3][26]/P0001 ,
		_w16372_,
		_w16373_
	);
	LUT2 #(
		.INIT('h8)
	) name15842 (
		_w16081_,
		_w16117_,
		_w16374_
	);
	LUT2 #(
		.INIT('h8)
	) name15843 (
		\u0_w_reg[3][30]/P0001 ,
		_w16112_,
		_w16375_
	);
	LUT2 #(
		.INIT('h8)
	) name15844 (
		_w16094_,
		_w16158_,
		_w16376_
	);
	LUT2 #(
		.INIT('h1)
	) name15845 (
		\u0_w_reg[3][25]/P0001 ,
		_w16088_,
		_w16377_
	);
	LUT2 #(
		.INIT('h4)
	) name15846 (
		_w16374_,
		_w16377_,
		_w16378_
	);
	LUT2 #(
		.INIT('h1)
	) name15847 (
		_w16375_,
		_w16376_,
		_w16379_
	);
	LUT2 #(
		.INIT('h8)
	) name15848 (
		_w16378_,
		_w16379_,
		_w16380_
	);
	LUT2 #(
		.INIT('h4)
	) name15849 (
		_w16101_,
		_w16380_,
		_w16381_
	);
	LUT2 #(
		.INIT('h4)
	) name15850 (
		_w16373_,
		_w16381_,
		_w16382_
	);
	LUT2 #(
		.INIT('h4)
	) name15851 (
		\u0_w_reg[3][26]/P0001 ,
		_w16052_,
		_w16383_
	);
	LUT2 #(
		.INIT('h2)
	) name15852 (
		\u0_w_reg[3][25]/P0001 ,
		_w16383_,
		_w16384_
	);
	LUT2 #(
		.INIT('h8)
	) name15853 (
		_w16048_,
		_w16145_,
		_w16385_
	);
	LUT2 #(
		.INIT('h1)
	) name15854 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w16386_
	);
	LUT2 #(
		.INIT('h8)
	) name15855 (
		_w16025_,
		_w16386_,
		_w16387_
	);
	LUT2 #(
		.INIT('h8)
	) name15856 (
		\u0_w_reg[3][28]/P0001 ,
		_w16171_,
		_w16388_
	);
	LUT2 #(
		.INIT('h4)
	) name15857 (
		_w16012_,
		_w16079_,
		_w16389_
	);
	LUT2 #(
		.INIT('h1)
	) name15858 (
		_w16388_,
		_w16389_,
		_w16390_
	);
	LUT2 #(
		.INIT('h2)
	) name15859 (
		\u0_w_reg[3][26]/P0001 ,
		_w16390_,
		_w16391_
	);
	LUT2 #(
		.INIT('h8)
	) name15860 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w16392_
	);
	LUT2 #(
		.INIT('h8)
	) name15861 (
		_w16171_,
		_w16392_,
		_w16393_
	);
	LUT2 #(
		.INIT('h1)
	) name15862 (
		_w16091_,
		_w16393_,
		_w16394_
	);
	LUT2 #(
		.INIT('h1)
	) name15863 (
		_w16385_,
		_w16387_,
		_w16395_
	);
	LUT2 #(
		.INIT('h8)
	) name15864 (
		_w16394_,
		_w16395_,
		_w16396_
	);
	LUT2 #(
		.INIT('h8)
	) name15865 (
		_w16384_,
		_w16396_,
		_w16397_
	);
	LUT2 #(
		.INIT('h4)
	) name15866 (
		_w16391_,
		_w16397_,
		_w16398_
	);
	LUT2 #(
		.INIT('h1)
	) name15867 (
		_w16382_,
		_w16398_,
		_w16399_
	);
	LUT2 #(
		.INIT('h1)
	) name15868 (
		_w16028_,
		_w16371_,
		_w16400_
	);
	LUT2 #(
		.INIT('h4)
	) name15869 (
		_w16399_,
		_w16400_,
		_w16401_
	);
	LUT2 #(
		.INIT('h2)
	) name15870 (
		\u0_w_reg[3][24]/P0001 ,
		_w16401_,
		_w16402_
	);
	LUT2 #(
		.INIT('h8)
	) name15871 (
		_w16105_,
		_w16392_,
		_w16403_
	);
	LUT2 #(
		.INIT('h1)
	) name15872 (
		_w16064_,
		_w16403_,
		_w16404_
	);
	LUT2 #(
		.INIT('h1)
	) name15873 (
		\u0_w_reg[3][26]/P0001 ,
		_w16404_,
		_w16405_
	);
	LUT2 #(
		.INIT('h4)
	) name15874 (
		\u0_w_reg[3][29]/P0001 ,
		_w16039_,
		_w16406_
	);
	LUT2 #(
		.INIT('h8)
	) name15875 (
		_w16017_,
		_w16048_,
		_w16407_
	);
	LUT2 #(
		.INIT('h8)
	) name15876 (
		\u0_w_reg[3][30]/P0001 ,
		_w16407_,
		_w16408_
	);
	LUT2 #(
		.INIT('h1)
	) name15877 (
		_w16406_,
		_w16408_,
		_w16409_
	);
	LUT2 #(
		.INIT('h2)
	) name15878 (
		\u0_w_reg[3][26]/P0001 ,
		_w16409_,
		_w16410_
	);
	LUT2 #(
		.INIT('h1)
	) name15879 (
		_w16045_,
		_w16087_,
		_w16411_
	);
	LUT2 #(
		.INIT('h2)
	) name15880 (
		_w16037_,
		_w16411_,
		_w16412_
	);
	LUT2 #(
		.INIT('h4)
	) name15881 (
		\u0_w_reg[3][26]/P0001 ,
		_w16150_,
		_w16413_
	);
	LUT2 #(
		.INIT('h2)
	) name15882 (
		\u0_w_reg[3][25]/P0001 ,
		_w16060_,
		_w16414_
	);
	LUT2 #(
		.INIT('h1)
	) name15883 (
		_w16412_,
		_w16413_,
		_w16415_
	);
	LUT2 #(
		.INIT('h8)
	) name15884 (
		_w16414_,
		_w16415_,
		_w16416_
	);
	LUT2 #(
		.INIT('h4)
	) name15885 (
		_w16410_,
		_w16416_,
		_w16417_
	);
	LUT2 #(
		.INIT('h1)
	) name15886 (
		_w16094_,
		_w16103_,
		_w16418_
	);
	LUT2 #(
		.INIT('h2)
	) name15887 (
		_w16105_,
		_w16418_,
		_w16419_
	);
	LUT2 #(
		.INIT('h8)
	) name15888 (
		\u0_w_reg[3][27]/P0001 ,
		_w16092_,
		_w16420_
	);
	LUT2 #(
		.INIT('h8)
	) name15889 (
		\u0_w_reg[3][31]/P0001 ,
		_w16036_,
		_w16421_
	);
	LUT2 #(
		.INIT('h4)
	) name15890 (
		_w16094_,
		_w16421_,
		_w16422_
	);
	LUT2 #(
		.INIT('h1)
	) name15891 (
		\u0_w_reg[3][25]/P0001 ,
		_w16361_,
		_w16423_
	);
	LUT2 #(
		.INIT('h1)
	) name15892 (
		_w16419_,
		_w16422_,
		_w16424_
	);
	LUT2 #(
		.INIT('h8)
	) name15893 (
		_w16423_,
		_w16424_,
		_w16425_
	);
	LUT2 #(
		.INIT('h4)
	) name15894 (
		_w16420_,
		_w16425_,
		_w16426_
	);
	LUT2 #(
		.INIT('h1)
	) name15895 (
		_w16417_,
		_w16426_,
		_w16427_
	);
	LUT2 #(
		.INIT('h8)
	) name15896 (
		_w16026_,
		_w16098_,
		_w16428_
	);
	LUT2 #(
		.INIT('h1)
	) name15897 (
		_w16165_,
		_w16428_,
		_w16429_
	);
	LUT2 #(
		.INIT('h2)
	) name15898 (
		\u0_w_reg[3][26]/P0001 ,
		_w16429_,
		_w16430_
	);
	LUT2 #(
		.INIT('h4)
	) name15899 (
		\u0_w_reg[3][27]/P0001 ,
		_w16040_,
		_w16431_
	);
	LUT2 #(
		.INIT('h1)
	) name15900 (
		_w16405_,
		_w16431_,
		_w16432_
	);
	LUT2 #(
		.INIT('h4)
	) name15901 (
		_w16430_,
		_w16432_,
		_w16433_
	);
	LUT2 #(
		.INIT('h4)
	) name15902 (
		_w16427_,
		_w16433_,
		_w16434_
	);
	LUT2 #(
		.INIT('h1)
	) name15903 (
		\u0_w_reg[3][24]/P0001 ,
		_w16434_,
		_w16435_
	);
	LUT2 #(
		.INIT('h2)
	) name15904 (
		\u0_w_reg[3][26]/P0001 ,
		_w16394_,
		_w16436_
	);
	LUT2 #(
		.INIT('h8)
	) name15905 (
		_w16032_,
		_w16142_,
		_w16437_
	);
	LUT2 #(
		.INIT('h8)
	) name15906 (
		\u0_w_reg[3][28]/P0001 ,
		_w16094_,
		_w16438_
	);
	LUT2 #(
		.INIT('h4)
	) name15907 (
		\u0_w_reg[3][28]/P0001 ,
		_w16025_,
		_w16439_
	);
	LUT2 #(
		.INIT('h1)
	) name15908 (
		_w16150_,
		_w16438_,
		_w16440_
	);
	LUT2 #(
		.INIT('h4)
	) name15909 (
		_w16439_,
		_w16440_,
		_w16441_
	);
	LUT2 #(
		.INIT('h2)
	) name15910 (
		_w16386_,
		_w16441_,
		_w16442_
	);
	LUT2 #(
		.INIT('h8)
	) name15911 (
		_w16094_,
		_w16359_,
		_w16443_
	);
	LUT2 #(
		.INIT('h8)
	) name15912 (
		_w16117_,
		_w16443_,
		_w16444_
	);
	LUT2 #(
		.INIT('h1)
	) name15913 (
		_w16437_,
		_w16444_,
		_w16445_
	);
	LUT2 #(
		.INIT('h4)
	) name15914 (
		_w16436_,
		_w16445_,
		_w16446_
	);
	LUT2 #(
		.INIT('h4)
	) name15915 (
		_w16442_,
		_w16446_,
		_w16447_
	);
	LUT2 #(
		.INIT('h2)
	) name15916 (
		\u0_w_reg[3][25]/P0001 ,
		_w16447_,
		_w16448_
	);
	LUT2 #(
		.INIT('h8)
	) name15917 (
		_w16169_,
		_w16392_,
		_w16449_
	);
	LUT2 #(
		.INIT('h8)
	) name15918 (
		\u0_w_reg[3][26]/P0001 ,
		_w16099_,
		_w16450_
	);
	LUT2 #(
		.INIT('h8)
	) name15919 (
		_w16098_,
		_w16109_,
		_w16451_
	);
	LUT2 #(
		.INIT('h1)
	) name15920 (
		_w16450_,
		_w16451_,
		_w16452_
	);
	LUT2 #(
		.INIT('h2)
	) name15921 (
		_w16032_,
		_w16452_,
		_w16453_
	);
	LUT2 #(
		.INIT('h8)
	) name15922 (
		\u0_w_reg[3][26]/P0001 ,
		_w16376_,
		_w16454_
	);
	LUT2 #(
		.INIT('h1)
	) name15923 (
		_w16053_,
		_w16431_,
		_w16455_
	);
	LUT2 #(
		.INIT('h4)
	) name15924 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		_w16456_
	);
	LUT2 #(
		.INIT('h4)
	) name15925 (
		_w16455_,
		_w16456_,
		_w16457_
	);
	LUT2 #(
		.INIT('h1)
	) name15926 (
		_w16449_,
		_w16454_,
		_w16458_
	);
	LUT2 #(
		.INIT('h4)
	) name15927 (
		_w16453_,
		_w16458_,
		_w16459_
	);
	LUT2 #(
		.INIT('h4)
	) name15928 (
		_w16457_,
		_w16459_,
		_w16460_
	);
	LUT2 #(
		.INIT('h4)
	) name15929 (
		_w16448_,
		_w16460_,
		_w16461_
	);
	LUT2 #(
		.INIT('h4)
	) name15930 (
		_w16435_,
		_w16461_,
		_w16462_
	);
	LUT2 #(
		.INIT('h4)
	) name15931 (
		_w16402_,
		_w16462_,
		_w16463_
	);
	LUT2 #(
		.INIT('h2)
	) name15932 (
		\u0_w_reg[0][3]/P0001 ,
		_w16463_,
		_w16464_
	);
	LUT2 #(
		.INIT('h4)
	) name15933 (
		\u0_w_reg[0][3]/P0001 ,
		_w16463_,
		_w16465_
	);
	LUT2 #(
		.INIT('h1)
	) name15934 (
		_w16464_,
		_w16465_,
		_w16466_
	);
	LUT2 #(
		.INIT('h2)
	) name15935 (
		\u0_w_reg[1][3]/P0001 ,
		\u0_w_reg[2][3]/P0001 ,
		_w16467_
	);
	LUT2 #(
		.INIT('h4)
	) name15936 (
		\u0_w_reg[1][3]/P0001 ,
		\u0_w_reg[2][3]/P0001 ,
		_w16468_
	);
	LUT2 #(
		.INIT('h1)
	) name15937 (
		_w16467_,
		_w16468_,
		_w16469_
	);
	LUT2 #(
		.INIT('h8)
	) name15938 (
		_w16466_,
		_w16469_,
		_w16470_
	);
	LUT2 #(
		.INIT('h1)
	) name15939 (
		_w16466_,
		_w16469_,
		_w16471_
	);
	LUT2 #(
		.INIT('h1)
	) name15940 (
		_w16470_,
		_w16471_,
		_w16472_
	);
	LUT2 #(
		.INIT('h4)
	) name15941 (
		ld_pad,
		_w16472_,
		_w16473_
	);
	LUT2 #(
		.INIT('h1)
	) name15942 (
		_w16358_,
		_w16473_,
		_w16474_
	);
	LUT2 #(
		.INIT('h4)
	) name15943 (
		\key[43]_pad ,
		ld_pad,
		_w16475_
	);
	LUT2 #(
		.INIT('h8)
	) name15944 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w16476_
	);
	LUT2 #(
		.INIT('h4)
	) name15945 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w16477_
	);
	LUT2 #(
		.INIT('h8)
	) name15946 (
		_w16476_,
		_w16477_,
		_w16478_
	);
	LUT2 #(
		.INIT('h4)
	) name15947 (
		\u0_w_reg[3][3]/P0001 ,
		_w16478_,
		_w16479_
	);
	LUT2 #(
		.INIT('h1)
	) name15948 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w16480_
	);
	LUT2 #(
		.INIT('h4)
	) name15949 (
		\u0_w_reg[3][4]/P0001 ,
		_w16480_,
		_w16481_
	);
	LUT2 #(
		.INIT('h4)
	) name15950 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		_w16482_
	);
	LUT2 #(
		.INIT('h2)
	) name15951 (
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w16483_
	);
	LUT2 #(
		.INIT('h8)
	) name15952 (
		_w16482_,
		_w16483_,
		_w16484_
	);
	LUT2 #(
		.INIT('h8)
	) name15953 (
		\u0_w_reg[3][4]/P0001 ,
		_w16484_,
		_w16485_
	);
	LUT2 #(
		.INIT('h1)
	) name15954 (
		_w16481_,
		_w16485_,
		_w16486_
	);
	LUT2 #(
		.INIT('h2)
	) name15955 (
		\u0_w_reg[3][2]/P0001 ,
		_w16486_,
		_w16487_
	);
	LUT2 #(
		.INIT('h2)
	) name15956 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w16488_
	);
	LUT2 #(
		.INIT('h4)
	) name15957 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w16489_
	);
	LUT2 #(
		.INIT('h8)
	) name15958 (
		_w16488_,
		_w16489_,
		_w16490_
	);
	LUT2 #(
		.INIT('h4)
	) name15959 (
		\u0_w_reg[3][2]/P0001 ,
		_w16490_,
		_w16491_
	);
	LUT2 #(
		.INIT('h8)
	) name15960 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w16492_
	);
	LUT2 #(
		.INIT('h1)
	) name15961 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w16493_
	);
	LUT2 #(
		.INIT('h8)
	) name15962 (
		_w16492_,
		_w16493_,
		_w16494_
	);
	LUT2 #(
		.INIT('h8)
	) name15963 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w16495_
	);
	LUT2 #(
		.INIT('h8)
	) name15964 (
		\u0_w_reg[3][4]/P0001 ,
		_w16492_,
		_w16496_
	);
	LUT2 #(
		.INIT('h8)
	) name15965 (
		_w16495_,
		_w16496_,
		_w16497_
	);
	LUT2 #(
		.INIT('h2)
	) name15966 (
		\u0_w_reg[3][1]/P0001 ,
		_w16494_,
		_w16498_
	);
	LUT2 #(
		.INIT('h4)
	) name15967 (
		_w16479_,
		_w16498_,
		_w16499_
	);
	LUT2 #(
		.INIT('h1)
	) name15968 (
		_w16491_,
		_w16497_,
		_w16500_
	);
	LUT2 #(
		.INIT('h8)
	) name15969 (
		_w16499_,
		_w16500_,
		_w16501_
	);
	LUT2 #(
		.INIT('h4)
	) name15970 (
		_w16487_,
		_w16501_,
		_w16502_
	);
	LUT2 #(
		.INIT('h4)
	) name15971 (
		\u0_w_reg[3][5]/P0001 ,
		_w16489_,
		_w16503_
	);
	LUT2 #(
		.INIT('h4)
	) name15972 (
		\u0_w_reg[3][3]/P0001 ,
		_w16503_,
		_w16504_
	);
	LUT2 #(
		.INIT('h2)
	) name15973 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w16505_
	);
	LUT2 #(
		.INIT('h2)
	) name15974 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w16506_
	);
	LUT2 #(
		.INIT('h1)
	) name15975 (
		_w16480_,
		_w16506_,
		_w16507_
	);
	LUT2 #(
		.INIT('h2)
	) name15976 (
		_w16505_,
		_w16507_,
		_w16508_
	);
	LUT2 #(
		.INIT('h4)
	) name15977 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w16509_
	);
	LUT2 #(
		.INIT('h8)
	) name15978 (
		_w16492_,
		_w16509_,
		_w16510_
	);
	LUT2 #(
		.INIT('h8)
	) name15979 (
		_w16488_,
		_w16510_,
		_w16511_
	);
	LUT2 #(
		.INIT('h2)
	) name15980 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w16512_
	);
	LUT2 #(
		.INIT('h2)
	) name15981 (
		\u0_w_reg[3][7]/P0001 ,
		_w16493_,
		_w16513_
	);
	LUT2 #(
		.INIT('h8)
	) name15982 (
		_w16512_,
		_w16513_,
		_w16514_
	);
	LUT2 #(
		.INIT('h1)
	) name15983 (
		\u0_w_reg[3][1]/P0001 ,
		_w16504_,
		_w16515_
	);
	LUT2 #(
		.INIT('h1)
	) name15984 (
		_w16508_,
		_w16511_,
		_w16516_
	);
	LUT2 #(
		.INIT('h4)
	) name15985 (
		_w16514_,
		_w16516_,
		_w16517_
	);
	LUT2 #(
		.INIT('h8)
	) name15986 (
		_w16515_,
		_w16517_,
		_w16518_
	);
	LUT2 #(
		.INIT('h1)
	) name15987 (
		_w16502_,
		_w16518_,
		_w16519_
	);
	LUT2 #(
		.INIT('h1)
	) name15988 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w16520_
	);
	LUT2 #(
		.INIT('h4)
	) name15989 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w16521_
	);
	LUT2 #(
		.INIT('h4)
	) name15990 (
		\u0_w_reg[3][7]/P0001 ,
		_w16521_,
		_w16522_
	);
	LUT2 #(
		.INIT('h8)
	) name15991 (
		_w16520_,
		_w16522_,
		_w16523_
	);
	LUT2 #(
		.INIT('h8)
	) name15992 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w16524_
	);
	LUT2 #(
		.INIT('h8)
	) name15993 (
		_w16481_,
		_w16524_,
		_w16525_
	);
	LUT2 #(
		.INIT('h8)
	) name15994 (
		\u0_w_reg[3][2]/P0001 ,
		_w16476_,
		_w16526_
	);
	LUT2 #(
		.INIT('h8)
	) name15995 (
		_w16477_,
		_w16526_,
		_w16527_
	);
	LUT2 #(
		.INIT('h8)
	) name15996 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w16528_
	);
	LUT2 #(
		.INIT('h8)
	) name15997 (
		_w16482_,
		_w16528_,
		_w16529_
	);
	LUT2 #(
		.INIT('h8)
	) name15998 (
		\u0_w_reg[3][6]/P0001 ,
		_w16529_,
		_w16530_
	);
	LUT2 #(
		.INIT('h2)
	) name15999 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w16531_
	);
	LUT2 #(
		.INIT('h8)
	) name16000 (
		\u0_w_reg[3][4]/P0001 ,
		_w16531_,
		_w16532_
	);
	LUT2 #(
		.INIT('h8)
	) name16001 (
		\u0_w_reg[3][6]/P0001 ,
		_w16532_,
		_w16533_
	);
	LUT2 #(
		.INIT('h1)
	) name16002 (
		_w16530_,
		_w16533_,
		_w16534_
	);
	LUT2 #(
		.INIT('h1)
	) name16003 (
		\u0_w_reg[3][2]/P0001 ,
		_w16534_,
		_w16535_
	);
	LUT2 #(
		.INIT('h1)
	) name16004 (
		\u0_w_reg[3][0]/P0001 ,
		_w16523_,
		_w16536_
	);
	LUT2 #(
		.INIT('h1)
	) name16005 (
		_w16525_,
		_w16527_,
		_w16537_
	);
	LUT2 #(
		.INIT('h8)
	) name16006 (
		_w16536_,
		_w16537_,
		_w16538_
	);
	LUT2 #(
		.INIT('h4)
	) name16007 (
		_w16535_,
		_w16538_,
		_w16539_
	);
	LUT2 #(
		.INIT('h4)
	) name16008 (
		_w16519_,
		_w16539_,
		_w16540_
	);
	LUT2 #(
		.INIT('h8)
	) name16009 (
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w16541_
	);
	LUT2 #(
		.INIT('h4)
	) name16010 (
		\u0_w_reg[3][5]/P0001 ,
		_w16541_,
		_w16542_
	);
	LUT2 #(
		.INIT('h4)
	) name16011 (
		\u0_w_reg[3][3]/P0001 ,
		_w16542_,
		_w16543_
	);
	LUT2 #(
		.INIT('h8)
	) name16012 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w16544_
	);
	LUT2 #(
		.INIT('h8)
	) name16013 (
		_w16480_,
		_w16544_,
		_w16545_
	);
	LUT2 #(
		.INIT('h1)
	) name16014 (
		_w16543_,
		_w16545_,
		_w16546_
	);
	LUT2 #(
		.INIT('h1)
	) name16015 (
		\u0_w_reg[3][2]/P0001 ,
		_w16546_,
		_w16547_
	);
	LUT2 #(
		.INIT('h1)
	) name16016 (
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w16548_
	);
	LUT2 #(
		.INIT('h8)
	) name16017 (
		_w16520_,
		_w16548_,
		_w16549_
	);
	LUT2 #(
		.INIT('h8)
	) name16018 (
		_w16495_,
		_w16506_,
		_w16550_
	);
	LUT2 #(
		.INIT('h2)
	) name16019 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w16551_
	);
	LUT2 #(
		.INIT('h2)
	) name16020 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w16552_
	);
	LUT2 #(
		.INIT('h8)
	) name16021 (
		_w16551_,
		_w16552_,
		_w16553_
	);
	LUT2 #(
		.INIT('h1)
	) name16022 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w16554_
	);
	LUT2 #(
		.INIT('h2)
	) name16023 (
		_w16494_,
		_w16554_,
		_w16555_
	);
	LUT2 #(
		.INIT('h8)
	) name16024 (
		_w16495_,
		_w16520_,
		_w16556_
	);
	LUT2 #(
		.INIT('h1)
	) name16025 (
		_w16549_,
		_w16550_,
		_w16557_
	);
	LUT2 #(
		.INIT('h1)
	) name16026 (
		_w16553_,
		_w16556_,
		_w16558_
	);
	LUT2 #(
		.INIT('h8)
	) name16027 (
		_w16557_,
		_w16558_,
		_w16559_
	);
	LUT2 #(
		.INIT('h4)
	) name16028 (
		_w16555_,
		_w16559_,
		_w16560_
	);
	LUT2 #(
		.INIT('h4)
	) name16029 (
		_w16547_,
		_w16560_,
		_w16561_
	);
	LUT2 #(
		.INIT('h1)
	) name16030 (
		\u0_w_reg[3][1]/P0001 ,
		_w16561_,
		_w16562_
	);
	LUT2 #(
		.INIT('h8)
	) name16031 (
		_w16488_,
		_w16528_,
		_w16563_
	);
	LUT2 #(
		.INIT('h4)
	) name16032 (
		\u0_w_reg[3][3]/P0001 ,
		_w16563_,
		_w16564_
	);
	LUT2 #(
		.INIT('h8)
	) name16033 (
		\u0_w_reg[3][3]/P0001 ,
		_w16476_,
		_w16565_
	);
	LUT2 #(
		.INIT('h8)
	) name16034 (
		\u0_w_reg[3][6]/P0001 ,
		_w16565_,
		_w16566_
	);
	LUT2 #(
		.INIT('h1)
	) name16035 (
		_w16564_,
		_w16566_,
		_w16567_
	);
	LUT2 #(
		.INIT('h1)
	) name16036 (
		\u0_w_reg[3][2]/P0001 ,
		_w16504_,
		_w16568_
	);
	LUT2 #(
		.INIT('h8)
	) name16037 (
		_w16567_,
		_w16568_,
		_w16569_
	);
	LUT2 #(
		.INIT('h4)
	) name16038 (
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w16570_
	);
	LUT2 #(
		.INIT('h8)
	) name16039 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w16571_
	);
	LUT2 #(
		.INIT('h8)
	) name16040 (
		_w16570_,
		_w16571_,
		_w16572_
	);
	LUT2 #(
		.INIT('h8)
	) name16041 (
		\u0_w_reg[3][4]/P0001 ,
		_w16522_,
		_w16573_
	);
	LUT2 #(
		.INIT('h4)
	) name16042 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w16574_
	);
	LUT2 #(
		.INIT('h8)
	) name16043 (
		_w16505_,
		_w16574_,
		_w16575_
	);
	LUT2 #(
		.INIT('h2)
	) name16044 (
		\u0_w_reg[3][2]/P0001 ,
		_w16572_,
		_w16576_
	);
	LUT2 #(
		.INIT('h4)
	) name16045 (
		_w16575_,
		_w16576_,
		_w16577_
	);
	LUT2 #(
		.INIT('h4)
	) name16046 (
		_w16573_,
		_w16577_,
		_w16578_
	);
	LUT2 #(
		.INIT('h1)
	) name16047 (
		_w16569_,
		_w16578_,
		_w16579_
	);
	LUT2 #(
		.INIT('h2)
	) name16048 (
		\u0_w_reg[3][4]/P0001 ,
		_w16544_,
		_w16580_
	);
	LUT2 #(
		.INIT('h8)
	) name16049 (
		_w16476_,
		_w16580_,
		_w16581_
	);
	LUT2 #(
		.INIT('h8)
	) name16050 (
		\u0_w_reg[3][4]/P0001 ,
		_w16574_,
		_w16582_
	);
	LUT2 #(
		.INIT('h2)
	) name16051 (
		_w16488_,
		_w16531_,
		_w16583_
	);
	LUT2 #(
		.INIT('h1)
	) name16052 (
		_w16582_,
		_w16583_,
		_w16584_
	);
	LUT2 #(
		.INIT('h2)
	) name16053 (
		\u0_w_reg[3][2]/P0001 ,
		_w16584_,
		_w16585_
	);
	LUT2 #(
		.INIT('h1)
	) name16054 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w16586_
	);
	LUT2 #(
		.INIT('h8)
	) name16055 (
		_w16493_,
		_w16586_,
		_w16587_
	);
	LUT2 #(
		.INIT('h1)
	) name16056 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w16588_
	);
	LUT2 #(
		.INIT('h8)
	) name16057 (
		_w16483_,
		_w16588_,
		_w16589_
	);
	LUT2 #(
		.INIT('h8)
	) name16058 (
		_w16544_,
		_w16574_,
		_w16590_
	);
	LUT2 #(
		.INIT('h1)
	) name16059 (
		_w16587_,
		_w16589_,
		_w16591_
	);
	LUT2 #(
		.INIT('h4)
	) name16060 (
		_w16590_,
		_w16591_,
		_w16592_
	);
	LUT2 #(
		.INIT('h4)
	) name16061 (
		_w16581_,
		_w16592_,
		_w16593_
	);
	LUT2 #(
		.INIT('h4)
	) name16062 (
		_w16585_,
		_w16593_,
		_w16594_
	);
	LUT2 #(
		.INIT('h2)
	) name16063 (
		\u0_w_reg[3][1]/P0001 ,
		_w16594_,
		_w16595_
	);
	LUT2 #(
		.INIT('h4)
	) name16064 (
		\u0_w_reg[3][4]/P0001 ,
		_w16551_,
		_w16596_
	);
	LUT2 #(
		.INIT('h8)
	) name16065 (
		_w16544_,
		_w16596_,
		_w16597_
	);
	LUT2 #(
		.INIT('h2)
	) name16066 (
		\u0_w_reg[3][0]/P0001 ,
		_w16597_,
		_w16598_
	);
	LUT2 #(
		.INIT('h4)
	) name16067 (
		_w16579_,
		_w16598_,
		_w16599_
	);
	LUT2 #(
		.INIT('h4)
	) name16068 (
		_w16562_,
		_w16599_,
		_w16600_
	);
	LUT2 #(
		.INIT('h4)
	) name16069 (
		_w16595_,
		_w16600_,
		_w16601_
	);
	LUT2 #(
		.INIT('h1)
	) name16070 (
		_w16540_,
		_w16601_,
		_w16602_
	);
	LUT2 #(
		.INIT('h1)
	) name16071 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		_w16603_
	);
	LUT2 #(
		.INIT('h8)
	) name16072 (
		_w16489_,
		_w16544_,
		_w16604_
	);
	LUT2 #(
		.INIT('h8)
	) name16073 (
		_w16603_,
		_w16604_,
		_w16605_
	);
	LUT2 #(
		.INIT('h8)
	) name16074 (
		_w16494_,
		_w16554_,
		_w16606_
	);
	LUT2 #(
		.INIT('h4)
	) name16075 (
		\u0_w_reg[3][4]/P0001 ,
		_w16483_,
		_w16607_
	);
	LUT2 #(
		.INIT('h8)
	) name16076 (
		\u0_w_reg[3][4]/P0001 ,
		_w16493_,
		_w16608_
	);
	LUT2 #(
		.INIT('h1)
	) name16077 (
		_w16490_,
		_w16607_,
		_w16609_
	);
	LUT2 #(
		.INIT('h4)
	) name16078 (
		_w16608_,
		_w16609_,
		_w16610_
	);
	LUT2 #(
		.INIT('h2)
	) name16079 (
		_w16588_,
		_w16610_,
		_w16611_
	);
	LUT2 #(
		.INIT('h2)
	) name16080 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w16612_
	);
	LUT2 #(
		.INIT('h8)
	) name16081 (
		_w16495_,
		_w16612_,
		_w16613_
	);
	LUT2 #(
		.INIT('h1)
	) name16082 (
		_w16563_,
		_w16613_,
		_w16614_
	);
	LUT2 #(
		.INIT('h2)
	) name16083 (
		\u0_w_reg[3][2]/P0001 ,
		_w16614_,
		_w16615_
	);
	LUT2 #(
		.INIT('h8)
	) name16084 (
		_w16524_,
		_w16542_,
		_w16616_
	);
	LUT2 #(
		.INIT('h1)
	) name16085 (
		_w16606_,
		_w16616_,
		_w16617_
	);
	LUT2 #(
		.INIT('h4)
	) name16086 (
		_w16615_,
		_w16617_,
		_w16618_
	);
	LUT2 #(
		.INIT('h4)
	) name16087 (
		_w16611_,
		_w16618_,
		_w16619_
	);
	LUT2 #(
		.INIT('h2)
	) name16088 (
		\u0_w_reg[3][1]/P0001 ,
		_w16619_,
		_w16620_
	);
	LUT2 #(
		.INIT('h4)
	) name16089 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		_w16621_
	);
	LUT2 #(
		.INIT('h4)
	) name16090 (
		\u0_w_reg[3][3]/P0001 ,
		_w16548_,
		_w16622_
	);
	LUT2 #(
		.INIT('h4)
	) name16091 (
		\u0_w_reg[3][5]/P0001 ,
		_w16622_,
		_w16623_
	);
	LUT2 #(
		.INIT('h8)
	) name16092 (
		\u0_w_reg[3][4]/P0001 ,
		_w16623_,
		_w16624_
	);
	LUT2 #(
		.INIT('h1)
	) name16093 (
		_w16523_,
		_w16624_,
		_w16625_
	);
	LUT2 #(
		.INIT('h2)
	) name16094 (
		_w16621_,
		_w16625_,
		_w16626_
	);
	LUT2 #(
		.INIT('h8)
	) name16095 (
		_w16477_,
		_w16574_,
		_w16627_
	);
	LUT2 #(
		.INIT('h1)
	) name16096 (
		_w16575_,
		_w16627_,
		_w16628_
	);
	LUT2 #(
		.INIT('h2)
	) name16097 (
		_w16524_,
		_w16628_,
		_w16629_
	);
	LUT2 #(
		.INIT('h4)
	) name16098 (
		\u0_w_reg[3][5]/P0001 ,
		_w16532_,
		_w16630_
	);
	LUT2 #(
		.INIT('h8)
	) name16099 (
		\u0_w_reg[3][6]/P0001 ,
		_w16630_,
		_w16631_
	);
	LUT2 #(
		.INIT('h1)
	) name16100 (
		_w16605_,
		_w16629_,
		_w16632_
	);
	LUT2 #(
		.INIT('h4)
	) name16101 (
		_w16631_,
		_w16632_,
		_w16633_
	);
	LUT2 #(
		.INIT('h4)
	) name16102 (
		_w16626_,
		_w16633_,
		_w16634_
	);
	LUT2 #(
		.INIT('h4)
	) name16103 (
		_w16620_,
		_w16634_,
		_w16635_
	);
	LUT2 #(
		.INIT('h4)
	) name16104 (
		_w16602_,
		_w16635_,
		_w16636_
	);
	LUT2 #(
		.INIT('h2)
	) name16105 (
		\u0_w_reg[0][11]/P0001 ,
		_w16636_,
		_w16637_
	);
	LUT2 #(
		.INIT('h4)
	) name16106 (
		\u0_w_reg[0][11]/P0001 ,
		_w16636_,
		_w16638_
	);
	LUT2 #(
		.INIT('h1)
	) name16107 (
		_w16637_,
		_w16638_,
		_w16639_
	);
	LUT2 #(
		.INIT('h2)
	) name16108 (
		\u0_w_reg[1][11]/P0001 ,
		\u0_w_reg[2][11]/P0001 ,
		_w16640_
	);
	LUT2 #(
		.INIT('h4)
	) name16109 (
		\u0_w_reg[1][11]/P0001 ,
		\u0_w_reg[2][11]/P0001 ,
		_w16641_
	);
	LUT2 #(
		.INIT('h1)
	) name16110 (
		_w16640_,
		_w16641_,
		_w16642_
	);
	LUT2 #(
		.INIT('h8)
	) name16111 (
		_w16639_,
		_w16642_,
		_w16643_
	);
	LUT2 #(
		.INIT('h1)
	) name16112 (
		_w16639_,
		_w16642_,
		_w16644_
	);
	LUT2 #(
		.INIT('h1)
	) name16113 (
		_w16643_,
		_w16644_,
		_w16645_
	);
	LUT2 #(
		.INIT('h4)
	) name16114 (
		ld_pad,
		_w16645_,
		_w16646_
	);
	LUT2 #(
		.INIT('h1)
	) name16115 (
		_w16475_,
		_w16646_,
		_w16647_
	);
	LUT2 #(
		.INIT('h4)
	) name16116 (
		\key[44]_pad ,
		ld_pad,
		_w16648_
	);
	LUT2 #(
		.INIT('h4)
	) name16117 (
		\u0_w_reg[3][4]/P0001 ,
		_w16476_,
		_w16649_
	);
	LUT2 #(
		.INIT('h8)
	) name16118 (
		_w16548_,
		_w16571_,
		_w16650_
	);
	LUT2 #(
		.INIT('h1)
	) name16119 (
		_w16649_,
		_w16650_,
		_w16651_
	);
	LUT2 #(
		.INIT('h1)
	) name16120 (
		\u0_w_reg[3][2]/P0001 ,
		_w16651_,
		_w16652_
	);
	LUT2 #(
		.INIT('h1)
	) name16121 (
		\u0_w_reg[3][5]/P0001 ,
		_w16477_,
		_w16653_
	);
	LUT2 #(
		.INIT('h2)
	) name16122 (
		_w16492_,
		_w16653_,
		_w16654_
	);
	LUT2 #(
		.INIT('h1)
	) name16123 (
		_w16652_,
		_w16654_,
		_w16655_
	);
	LUT2 #(
		.INIT('h1)
	) name16124 (
		\u0_w_reg[3][1]/P0001 ,
		_w16655_,
		_w16656_
	);
	LUT2 #(
		.INIT('h8)
	) name16125 (
		_w16483_,
		_w16612_,
		_w16657_
	);
	LUT2 #(
		.INIT('h1)
	) name16126 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w16658_
	);
	LUT2 #(
		.INIT('h8)
	) name16127 (
		_w16493_,
		_w16658_,
		_w16659_
	);
	LUT2 #(
		.INIT('h4)
	) name16128 (
		\u0_w_reg[3][3]/P0001 ,
		_w16659_,
		_w16660_
	);
	LUT2 #(
		.INIT('h1)
	) name16129 (
		_w16590_,
		_w16657_,
		_w16661_
	);
	LUT2 #(
		.INIT('h4)
	) name16130 (
		_w16660_,
		_w16661_,
		_w16662_
	);
	LUT2 #(
		.INIT('h1)
	) name16131 (
		\u0_w_reg[3][2]/P0001 ,
		_w16662_,
		_w16663_
	);
	LUT2 #(
		.INIT('h4)
	) name16132 (
		\u0_w_reg[3][4]/P0001 ,
		_w16524_,
		_w16664_
	);
	LUT2 #(
		.INIT('h4)
	) name16133 (
		\u0_w_reg[3][6]/P0001 ,
		_w16664_,
		_w16665_
	);
	LUT2 #(
		.INIT('h4)
	) name16134 (
		\u0_w_reg[3][1]/P0001 ,
		_w16563_,
		_w16666_
	);
	LUT2 #(
		.INIT('h4)
	) name16135 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w16667_
	);
	LUT2 #(
		.INIT('h4)
	) name16136 (
		\u0_w_reg[3][7]/P0001 ,
		_w16667_,
		_w16668_
	);
	LUT2 #(
		.INIT('h1)
	) name16137 (
		_w16494_,
		_w16668_,
		_w16669_
	);
	LUT2 #(
		.INIT('h4)
	) name16138 (
		_w16666_,
		_w16669_,
		_w16670_
	);
	LUT2 #(
		.INIT('h2)
	) name16139 (
		\u0_w_reg[3][2]/P0001 ,
		_w16670_,
		_w16671_
	);
	LUT2 #(
		.INIT('h1)
	) name16140 (
		_w16575_,
		_w16607_,
		_w16672_
	);
	LUT2 #(
		.INIT('h1)
	) name16141 (
		\u0_w_reg[3][2]/P0001 ,
		_w16672_,
		_w16673_
	);
	LUT2 #(
		.INIT('h8)
	) name16142 (
		_w16552_,
		_w16570_,
		_w16674_
	);
	LUT2 #(
		.INIT('h8)
	) name16143 (
		\u0_w_reg[3][3]/P0001 ,
		_w16658_,
		_w16675_
	);
	LUT2 #(
		.INIT('h8)
	) name16144 (
		_w16488_,
		_w16675_,
		_w16676_
	);
	LUT2 #(
		.INIT('h1)
	) name16145 (
		_w16674_,
		_w16676_,
		_w16677_
	);
	LUT2 #(
		.INIT('h4)
	) name16146 (
		_w16624_,
		_w16677_,
		_w16678_
	);
	LUT2 #(
		.INIT('h4)
	) name16147 (
		_w16673_,
		_w16678_,
		_w16679_
	);
	LUT2 #(
		.INIT('h2)
	) name16148 (
		\u0_w_reg[3][1]/P0001 ,
		_w16679_,
		_w16680_
	);
	LUT2 #(
		.INIT('h2)
	) name16149 (
		\u0_w_reg[3][0]/P0001 ,
		_w16527_,
		_w16681_
	);
	LUT2 #(
		.INIT('h4)
	) name16150 (
		_w16665_,
		_w16681_,
		_w16682_
	);
	LUT2 #(
		.INIT('h4)
	) name16151 (
		_w16663_,
		_w16682_,
		_w16683_
	);
	LUT2 #(
		.INIT('h4)
	) name16152 (
		_w16671_,
		_w16683_,
		_w16684_
	);
	LUT2 #(
		.INIT('h4)
	) name16153 (
		_w16656_,
		_w16684_,
		_w16685_
	);
	LUT2 #(
		.INIT('h4)
	) name16154 (
		_w16680_,
		_w16685_,
		_w16686_
	);
	LUT2 #(
		.INIT('h8)
	) name16155 (
		\u0_w_reg[3][4]/P0001 ,
		_w16495_,
		_w16687_
	);
	LUT2 #(
		.INIT('h8)
	) name16156 (
		\u0_w_reg[3][2]/P0001 ,
		_w16687_,
		_w16688_
	);
	LUT2 #(
		.INIT('h2)
	) name16157 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		_w16689_
	);
	LUT2 #(
		.INIT('h1)
	) name16158 (
		_w16612_,
		_w16689_,
		_w16690_
	);
	LUT2 #(
		.INIT('h2)
	) name16159 (
		_w16548_,
		_w16690_,
		_w16691_
	);
	LUT2 #(
		.INIT('h8)
	) name16160 (
		\u0_w_reg[3][5]/P0001 ,
		_w16589_,
		_w16692_
	);
	LUT2 #(
		.INIT('h1)
	) name16161 (
		_w16688_,
		_w16691_,
		_w16693_
	);
	LUT2 #(
		.INIT('h4)
	) name16162 (
		_w16692_,
		_w16693_,
		_w16694_
	);
	LUT2 #(
		.INIT('h1)
	) name16163 (
		\u0_w_reg[3][1]/P0001 ,
		_w16694_,
		_w16695_
	);
	LUT2 #(
		.INIT('h8)
	) name16164 (
		_w16509_,
		_w16542_,
		_w16696_
	);
	LUT2 #(
		.INIT('h8)
	) name16165 (
		_w16488_,
		_w16658_,
		_w16697_
	);
	LUT2 #(
		.INIT('h1)
	) name16166 (
		_w16696_,
		_w16697_,
		_w16698_
	);
	LUT2 #(
		.INIT('h1)
	) name16167 (
		\u0_w_reg[3][3]/P0001 ,
		_w16698_,
		_w16699_
	);
	LUT2 #(
		.INIT('h4)
	) name16168 (
		\u0_w_reg[3][4]/P0001 ,
		_w16521_,
		_w16700_
	);
	LUT2 #(
		.INIT('h8)
	) name16169 (
		_w16493_,
		_w16531_,
		_w16701_
	);
	LUT2 #(
		.INIT('h1)
	) name16170 (
		_w16700_,
		_w16701_,
		_w16702_
	);
	LUT2 #(
		.INIT('h2)
	) name16171 (
		\u0_w_reg[3][2]/P0001 ,
		_w16612_,
		_w16703_
	);
	LUT2 #(
		.INIT('h4)
	) name16172 (
		_w16702_,
		_w16703_,
		_w16704_
	);
	LUT2 #(
		.INIT('h8)
	) name16173 (
		_w16489_,
		_w16493_,
		_w16705_
	);
	LUT2 #(
		.INIT('h8)
	) name16174 (
		\u0_w_reg[3][5]/P0001 ,
		_w16570_,
		_w16706_
	);
	LUT2 #(
		.INIT('h4)
	) name16175 (
		_w16612_,
		_w16706_,
		_w16707_
	);
	LUT2 #(
		.INIT('h1)
	) name16176 (
		_w16705_,
		_w16707_,
		_w16708_
	);
	LUT2 #(
		.INIT('h1)
	) name16177 (
		\u0_w_reg[3][2]/P0001 ,
		_w16708_,
		_w16709_
	);
	LUT2 #(
		.INIT('h8)
	) name16178 (
		_w16512_,
		_w16582_,
		_w16710_
	);
	LUT2 #(
		.INIT('h1)
	) name16179 (
		_w16533_,
		_w16550_,
		_w16711_
	);
	LUT2 #(
		.INIT('h4)
	) name16180 (
		_w16710_,
		_w16711_,
		_w16712_
	);
	LUT2 #(
		.INIT('h4)
	) name16181 (
		_w16709_,
		_w16712_,
		_w16713_
	);
	LUT2 #(
		.INIT('h2)
	) name16182 (
		\u0_w_reg[3][1]/P0001 ,
		_w16713_,
		_w16714_
	);
	LUT2 #(
		.INIT('h1)
	) name16183 (
		\u0_w_reg[3][0]/P0001 ,
		_w16704_,
		_w16715_
	);
	LUT2 #(
		.INIT('h4)
	) name16184 (
		_w16699_,
		_w16715_,
		_w16716_
	);
	LUT2 #(
		.INIT('h4)
	) name16185 (
		_w16695_,
		_w16716_,
		_w16717_
	);
	LUT2 #(
		.INIT('h4)
	) name16186 (
		_w16714_,
		_w16717_,
		_w16718_
	);
	LUT2 #(
		.INIT('h1)
	) name16187 (
		_w16686_,
		_w16718_,
		_w16719_
	);
	LUT2 #(
		.INIT('h8)
	) name16188 (
		_w16522_,
		_w16554_,
		_w16720_
	);
	LUT2 #(
		.INIT('h1)
	) name16189 (
		_w16688_,
		_w16720_,
		_w16721_
	);
	LUT2 #(
		.INIT('h2)
	) name16190 (
		\u0_w_reg[3][3]/P0001 ,
		_w16721_,
		_w16722_
	);
	LUT2 #(
		.INIT('h8)
	) name16191 (
		_w16544_,
		_w16649_,
		_w16723_
	);
	LUT2 #(
		.INIT('h1)
	) name16192 (
		\u0_w_reg[3][2]/P0001 ,
		_w16723_,
		_w16724_
	);
	LUT2 #(
		.INIT('h4)
	) name16193 (
		\u0_w_reg[3][3]/P0001 ,
		_w16521_,
		_w16725_
	);
	LUT2 #(
		.INIT('h4)
	) name16194 (
		_w16658_,
		_w16725_,
		_w16726_
	);
	LUT2 #(
		.INIT('h2)
	) name16195 (
		_w16724_,
		_w16726_,
		_w16727_
	);
	LUT2 #(
		.INIT('h8)
	) name16196 (
		_w16544_,
		_w16551_,
		_w16728_
	);
	LUT2 #(
		.INIT('h8)
	) name16197 (
		_w16488_,
		_w16612_,
		_w16729_
	);
	LUT2 #(
		.INIT('h4)
	) name16198 (
		\u0_w_reg[3][3]/P0001 ,
		_w16705_,
		_w16730_
	);
	LUT2 #(
		.INIT('h2)
	) name16199 (
		\u0_w_reg[3][2]/P0001 ,
		_w16730_,
		_w16731_
	);
	LUT2 #(
		.INIT('h8)
	) name16200 (
		_w16492_,
		_w16608_,
		_w16732_
	);
	LUT2 #(
		.INIT('h1)
	) name16201 (
		_w16728_,
		_w16729_,
		_w16733_
	);
	LUT2 #(
		.INIT('h4)
	) name16202 (
		_w16732_,
		_w16733_,
		_w16734_
	);
	LUT2 #(
		.INIT('h8)
	) name16203 (
		_w16731_,
		_w16734_,
		_w16735_
	);
	LUT2 #(
		.INIT('h1)
	) name16204 (
		_w16727_,
		_w16735_,
		_w16736_
	);
	LUT2 #(
		.INIT('h8)
	) name16205 (
		_w16495_,
		_w16532_,
		_w16737_
	);
	LUT2 #(
		.INIT('h2)
	) name16206 (
		_w16482_,
		_w16509_,
		_w16738_
	);
	LUT2 #(
		.INIT('h8)
	) name16207 (
		_w16548_,
		_w16738_,
		_w16739_
	);
	LUT2 #(
		.INIT('h1)
	) name16208 (
		\u0_w_reg[3][1]/P0001 ,
		_w16737_,
		_w16740_
	);
	LUT2 #(
		.INIT('h4)
	) name16209 (
		_w16739_,
		_w16740_,
		_w16741_
	);
	LUT2 #(
		.INIT('h4)
	) name16210 (
		_w16736_,
		_w16741_,
		_w16742_
	);
	LUT2 #(
		.INIT('h4)
	) name16211 (
		\u0_w_reg[3][5]/P0001 ,
		_w16612_,
		_w16743_
	);
	LUT2 #(
		.INIT('h8)
	) name16212 (
		_w16570_,
		_w16743_,
		_w16744_
	);
	LUT2 #(
		.INIT('h8)
	) name16213 (
		_w16483_,
		_w16512_,
		_w16745_
	);
	LUT2 #(
		.INIT('h1)
	) name16214 (
		_w16590_,
		_w16745_,
		_w16746_
	);
	LUT2 #(
		.INIT('h2)
	) name16215 (
		\u0_w_reg[3][4]/P0001 ,
		_w16746_,
		_w16747_
	);
	LUT2 #(
		.INIT('h2)
	) name16216 (
		\u0_w_reg[3][3]/P0001 ,
		_w16548_,
		_w16748_
	);
	LUT2 #(
		.INIT('h1)
	) name16217 (
		_w16549_,
		_w16748_,
		_w16749_
	);
	LUT2 #(
		.INIT('h1)
	) name16218 (
		\u0_w_reg[3][5]/P0001 ,
		_w16749_,
		_w16750_
	);
	LUT2 #(
		.INIT('h1)
	) name16219 (
		_w16479_,
		_w16750_,
		_w16751_
	);
	LUT2 #(
		.INIT('h1)
	) name16220 (
		\u0_w_reg[3][2]/P0001 ,
		_w16751_,
		_w16752_
	);
	LUT2 #(
		.INIT('h8)
	) name16221 (
		\u0_w_reg[3][5]/P0001 ,
		_w16548_,
		_w16753_
	);
	LUT2 #(
		.INIT('h8)
	) name16222 (
		_w16524_,
		_w16753_,
		_w16754_
	);
	LUT2 #(
		.INIT('h2)
	) name16223 (
		\u0_w_reg[3][1]/P0001 ,
		_w16744_,
		_w16755_
	);
	LUT2 #(
		.INIT('h4)
	) name16224 (
		_w16754_,
		_w16755_,
		_w16756_
	);
	LUT2 #(
		.INIT('h4)
	) name16225 (
		_w16747_,
		_w16756_,
		_w16757_
	);
	LUT2 #(
		.INIT('h4)
	) name16226 (
		_w16752_,
		_w16757_,
		_w16758_
	);
	LUT2 #(
		.INIT('h1)
	) name16227 (
		_w16742_,
		_w16758_,
		_w16759_
	);
	LUT2 #(
		.INIT('h1)
	) name16228 (
		_w16722_,
		_w16759_,
		_w16760_
	);
	LUT2 #(
		.INIT('h4)
	) name16229 (
		_w16719_,
		_w16760_,
		_w16761_
	);
	LUT2 #(
		.INIT('h2)
	) name16230 (
		\u0_w_reg[0][12]/P0001 ,
		_w16761_,
		_w16762_
	);
	LUT2 #(
		.INIT('h4)
	) name16231 (
		\u0_w_reg[0][12]/P0001 ,
		_w16761_,
		_w16763_
	);
	LUT2 #(
		.INIT('h1)
	) name16232 (
		_w16762_,
		_w16763_,
		_w16764_
	);
	LUT2 #(
		.INIT('h2)
	) name16233 (
		\u0_w_reg[1][12]/P0001 ,
		\u0_w_reg[2][12]/P0001 ,
		_w16765_
	);
	LUT2 #(
		.INIT('h4)
	) name16234 (
		\u0_w_reg[1][12]/P0001 ,
		\u0_w_reg[2][12]/P0001 ,
		_w16766_
	);
	LUT2 #(
		.INIT('h1)
	) name16235 (
		_w16765_,
		_w16766_,
		_w16767_
	);
	LUT2 #(
		.INIT('h8)
	) name16236 (
		_w16764_,
		_w16767_,
		_w16768_
	);
	LUT2 #(
		.INIT('h1)
	) name16237 (
		_w16764_,
		_w16767_,
		_w16769_
	);
	LUT2 #(
		.INIT('h1)
	) name16238 (
		_w16768_,
		_w16769_,
		_w16770_
	);
	LUT2 #(
		.INIT('h4)
	) name16239 (
		ld_pad,
		_w16770_,
		_w16771_
	);
	LUT2 #(
		.INIT('h1)
	) name16240 (
		_w16648_,
		_w16771_,
		_w16772_
	);
	LUT2 #(
		.INIT('h8)
	) name16241 (
		\key[120]_pad ,
		ld_pad,
		_w16773_
	);
	LUT2 #(
		.INIT('h8)
	) name16242 (
		\u0_w_reg[3][21]/P0001 ,
		_w15520_,
		_w16774_
	);
	LUT2 #(
		.INIT('h1)
	) name16243 (
		_w15518_,
		_w16774_,
		_w16775_
	);
	LUT2 #(
		.INIT('h2)
	) name16244 (
		_w16266_,
		_w16775_,
		_w16776_
	);
	LUT2 #(
		.INIT('h8)
	) name16245 (
		\u0_w_reg[3][18]/P0001 ,
		_w15516_,
		_w16777_
	);
	LUT2 #(
		.INIT('h8)
	) name16246 (
		\u0_w_reg[3][19]/P0001 ,
		_w16777_,
		_w16778_
	);
	LUT2 #(
		.INIT('h8)
	) name16247 (
		\u0_w_reg[3][20]/P0001 ,
		_w16229_,
		_w16779_
	);
	LUT2 #(
		.INIT('h1)
	) name16248 (
		_w15660_,
		_w16779_,
		_w16780_
	);
	LUT2 #(
		.INIT('h2)
	) name16249 (
		\u0_w_reg[3][23]/P0001 ,
		_w16780_,
		_w16781_
	);
	LUT2 #(
		.INIT('h2)
	) name16250 (
		_w15520_,
		_w15521_,
		_w16782_
	);
	LUT2 #(
		.INIT('h2)
	) name16251 (
		\u0_w_reg[3][17]/P0001 ,
		_w16782_,
		_w16783_
	);
	LUT2 #(
		.INIT('h4)
	) name16252 (
		_w16778_,
		_w16783_,
		_w16784_
	);
	LUT2 #(
		.INIT('h4)
	) name16253 (
		_w16781_,
		_w16784_,
		_w16785_
	);
	LUT2 #(
		.INIT('h1)
	) name16254 (
		_w16283_,
		_w16313_,
		_w16786_
	);
	LUT2 #(
		.INIT('h1)
	) name16255 (
		\u0_w_reg[3][19]/P0001 ,
		_w16786_,
		_w16787_
	);
	LUT2 #(
		.INIT('h2)
	) name16256 (
		_w15526_,
		_w16229_,
		_w16788_
	);
	LUT2 #(
		.INIT('h2)
	) name16257 (
		\u0_w_reg[3][18]/P0001 ,
		_w16788_,
		_w16789_
	);
	LUT2 #(
		.INIT('h1)
	) name16258 (
		\u0_w_reg[3][18]/P0001 ,
		_w15522_,
		_w16790_
	);
	LUT2 #(
		.INIT('h1)
	) name16259 (
		_w16789_,
		_w16790_,
		_w16791_
	);
	LUT2 #(
		.INIT('h1)
	) name16260 (
		\u0_w_reg[3][17]/P0001 ,
		_w16791_,
		_w16792_
	);
	LUT2 #(
		.INIT('h4)
	) name16261 (
		_w16787_,
		_w16792_,
		_w16793_
	);
	LUT2 #(
		.INIT('h1)
	) name16262 (
		_w16785_,
		_w16793_,
		_w16794_
	);
	LUT2 #(
		.INIT('h8)
	) name16263 (
		_w15506_,
		_w15549_,
		_w16795_
	);
	LUT2 #(
		.INIT('h1)
	) name16264 (
		_w16242_,
		_w16795_,
		_w16796_
	);
	LUT2 #(
		.INIT('h4)
	) name16265 (
		_w15561_,
		_w16796_,
		_w16797_
	);
	LUT2 #(
		.INIT('h1)
	) name16266 (
		\u0_w_reg[3][18]/P0001 ,
		_w16797_,
		_w16798_
	);
	LUT2 #(
		.INIT('h1)
	) name16267 (
		_w16776_,
		_w16798_,
		_w16799_
	);
	LUT2 #(
		.INIT('h4)
	) name16268 (
		_w16794_,
		_w16799_,
		_w16800_
	);
	LUT2 #(
		.INIT('h1)
	) name16269 (
		\u0_w_reg[3][16]/P0001 ,
		_w16800_,
		_w16801_
	);
	LUT2 #(
		.INIT('h4)
	) name16270 (
		\u0_w_reg[3][20]/P0001 ,
		_w15587_,
		_w16802_
	);
	LUT2 #(
		.INIT('h1)
	) name16271 (
		_w15563_,
		_w16802_,
		_w16803_
	);
	LUT2 #(
		.INIT('h2)
	) name16272 (
		\u0_w_reg[3][18]/P0001 ,
		_w16269_,
		_w16804_
	);
	LUT2 #(
		.INIT('h4)
	) name16273 (
		_w15561_,
		_w16804_,
		_w16805_
	);
	LUT2 #(
		.INIT('h8)
	) name16274 (
		_w16803_,
		_w16805_,
		_w16806_
	);
	LUT2 #(
		.INIT('h8)
	) name16275 (
		_w15525_,
		_w15542_,
		_w16807_
	);
	LUT2 #(
		.INIT('h1)
	) name16276 (
		_w15518_,
		_w15613_,
		_w16808_
	);
	LUT2 #(
		.INIT('h2)
	) name16277 (
		\u0_w_reg[3][19]/P0001 ,
		_w16808_,
		_w16809_
	);
	LUT2 #(
		.INIT('h1)
	) name16278 (
		\u0_w_reg[3][18]/P0001 ,
		_w16807_,
		_w16810_
	);
	LUT2 #(
		.INIT('h4)
	) name16279 (
		_w15514_,
		_w16810_,
		_w16811_
	);
	LUT2 #(
		.INIT('h4)
	) name16280 (
		_w16809_,
		_w16811_,
		_w16812_
	);
	LUT2 #(
		.INIT('h1)
	) name16281 (
		_w16806_,
		_w16812_,
		_w16813_
	);
	LUT2 #(
		.INIT('h4)
	) name16282 (
		\u0_w_reg[3][19]/P0001 ,
		_w15516_,
		_w16814_
	);
	LUT2 #(
		.INIT('h8)
	) name16283 (
		_w15530_,
		_w15662_,
		_w16815_
	);
	LUT2 #(
		.INIT('h1)
	) name16284 (
		_w15545_,
		_w15585_,
		_w16816_
	);
	LUT2 #(
		.INIT('h2)
	) name16285 (
		\u0_w_reg[3][18]/P0001 ,
		_w16816_,
		_w16817_
	);
	LUT2 #(
		.INIT('h1)
	) name16286 (
		_w15543_,
		_w15600_,
		_w16818_
	);
	LUT2 #(
		.INIT('h1)
	) name16287 (
		\u0_w_reg[3][19]/P0001 ,
		_w16818_,
		_w16819_
	);
	LUT2 #(
		.INIT('h8)
	) name16288 (
		_w15530_,
		_w15660_,
		_w16820_
	);
	LUT2 #(
		.INIT('h8)
	) name16289 (
		\u0_w_reg[3][20]/P0001 ,
		_w16820_,
		_w16821_
	);
	LUT2 #(
		.INIT('h1)
	) name16290 (
		\u0_w_reg[3][17]/P0001 ,
		_w15556_,
		_w16822_
	);
	LUT2 #(
		.INIT('h4)
	) name16291 (
		_w15662_,
		_w16822_,
		_w16823_
	);
	LUT2 #(
		.INIT('h4)
	) name16292 (
		_w16817_,
		_w16823_,
		_w16824_
	);
	LUT2 #(
		.INIT('h4)
	) name16293 (
		_w16821_,
		_w16824_,
		_w16825_
	);
	LUT2 #(
		.INIT('h4)
	) name16294 (
		_w16819_,
		_w16825_,
		_w16826_
	);
	LUT2 #(
		.INIT('h4)
	) name16295 (
		\u0_w_reg[3][18]/P0001 ,
		_w15512_,
		_w16827_
	);
	LUT2 #(
		.INIT('h2)
	) name16296 (
		\u0_w_reg[3][17]/P0001 ,
		_w15618_,
		_w16828_
	);
	LUT2 #(
		.INIT('h4)
	) name16297 (
		_w16827_,
		_w16828_,
		_w16829_
	);
	LUT2 #(
		.INIT('h4)
	) name16298 (
		_w16232_,
		_w16829_,
		_w16830_
	);
	LUT2 #(
		.INIT('h1)
	) name16299 (
		_w16826_,
		_w16830_,
		_w16831_
	);
	LUT2 #(
		.INIT('h1)
	) name16300 (
		_w16814_,
		_w16815_,
		_w16832_
	);
	LUT2 #(
		.INIT('h4)
	) name16301 (
		_w16813_,
		_w16832_,
		_w16833_
	);
	LUT2 #(
		.INIT('h4)
	) name16302 (
		_w16831_,
		_w16833_,
		_w16834_
	);
	LUT2 #(
		.INIT('h2)
	) name16303 (
		\u0_w_reg[3][16]/P0001 ,
		_w16834_,
		_w16835_
	);
	LUT2 #(
		.INIT('h8)
	) name16304 (
		_w15529_,
		_w15544_,
		_w16836_
	);
	LUT2 #(
		.INIT('h8)
	) name16305 (
		_w15507_,
		_w15542_,
		_w16837_
	);
	LUT2 #(
		.INIT('h1)
	) name16306 (
		_w16836_,
		_w16837_,
		_w16838_
	);
	LUT2 #(
		.INIT('h2)
	) name16307 (
		\u0_w_reg[3][22]/P0001 ,
		_w16838_,
		_w16839_
	);
	LUT2 #(
		.INIT('h8)
	) name16308 (
		\u0_w_reg[3][20]/P0001 ,
		_w15518_,
		_w16840_
	);
	LUT2 #(
		.INIT('h8)
	) name16309 (
		_w15511_,
		_w16840_,
		_w16841_
	);
	LUT2 #(
		.INIT('h1)
	) name16310 (
		_w15657_,
		_w16795_,
		_w16842_
	);
	LUT2 #(
		.INIT('h4)
	) name16311 (
		_w16841_,
		_w16842_,
		_w16843_
	);
	LUT2 #(
		.INIT('h1)
	) name16312 (
		\u0_w_reg[3][23]/P0001 ,
		_w16843_,
		_w16844_
	);
	LUT2 #(
		.INIT('h8)
	) name16313 (
		_w15531_,
		_w15608_,
		_w16845_
	);
	LUT2 #(
		.INIT('h2)
	) name16314 (
		\u0_w_reg[3][17]/P0001 ,
		_w16239_,
		_w16846_
	);
	LUT2 #(
		.INIT('h4)
	) name16315 (
		_w16845_,
		_w16846_,
		_w16847_
	);
	LUT2 #(
		.INIT('h4)
	) name16316 (
		_w16844_,
		_w16847_,
		_w16848_
	);
	LUT2 #(
		.INIT('h1)
	) name16317 (
		_w15512_,
		_w15531_,
		_w16849_
	);
	LUT2 #(
		.INIT('h2)
	) name16318 (
		_w15507_,
		_w16849_,
		_w16850_
	);
	LUT2 #(
		.INIT('h8)
	) name16319 (
		_w15512_,
		_w15613_,
		_w16851_
	);
	LUT2 #(
		.INIT('h8)
	) name16320 (
		_w15529_,
		_w16851_,
		_w16852_
	);
	LUT2 #(
		.INIT('h8)
	) name16321 (
		_w15559_,
		_w15613_,
		_w16853_
	);
	LUT2 #(
		.INIT('h8)
	) name16322 (
		\u0_w_reg[3][20]/P0001 ,
		_w15503_,
		_w16854_
	);
	LUT2 #(
		.INIT('h1)
	) name16323 (
		_w15638_,
		_w16853_,
		_w16855_
	);
	LUT2 #(
		.INIT('h4)
	) name16324 (
		_w16854_,
		_w16855_,
		_w16856_
	);
	LUT2 #(
		.INIT('h2)
	) name16325 (
		_w15648_,
		_w16856_,
		_w16857_
	);
	LUT2 #(
		.INIT('h1)
	) name16326 (
		\u0_w_reg[3][17]/P0001 ,
		_w15656_,
		_w16858_
	);
	LUT2 #(
		.INIT('h4)
	) name16327 (
		_w16852_,
		_w16858_,
		_w16859_
	);
	LUT2 #(
		.INIT('h4)
	) name16328 (
		_w16850_,
		_w16859_,
		_w16860_
	);
	LUT2 #(
		.INIT('h4)
	) name16329 (
		_w16857_,
		_w16860_,
		_w16861_
	);
	LUT2 #(
		.INIT('h1)
	) name16330 (
		_w16848_,
		_w16861_,
		_w16862_
	);
	LUT2 #(
		.INIT('h1)
	) name16331 (
		_w16839_,
		_w16862_,
		_w16863_
	);
	LUT2 #(
		.INIT('h4)
	) name16332 (
		_w16801_,
		_w16863_,
		_w16864_
	);
	LUT2 #(
		.INIT('h4)
	) name16333 (
		_w16835_,
		_w16864_,
		_w16865_
	);
	LUT2 #(
		.INIT('h2)
	) name16334 (
		\u0_r0_out_reg[24]/P0001 ,
		\u0_w_reg[0][24]/P0001 ,
		_w16866_
	);
	LUT2 #(
		.INIT('h4)
	) name16335 (
		\u0_r0_out_reg[24]/P0001 ,
		\u0_w_reg[0][24]/P0001 ,
		_w16867_
	);
	LUT2 #(
		.INIT('h1)
	) name16336 (
		_w16866_,
		_w16867_,
		_w16868_
	);
	LUT2 #(
		.INIT('h1)
	) name16337 (
		_w16865_,
		_w16868_,
		_w16869_
	);
	LUT2 #(
		.INIT('h8)
	) name16338 (
		_w16865_,
		_w16868_,
		_w16870_
	);
	LUT2 #(
		.INIT('h1)
	) name16339 (
		_w16869_,
		_w16870_,
		_w16871_
	);
	LUT2 #(
		.INIT('h4)
	) name16340 (
		ld_pad,
		_w16871_,
		_w16872_
	);
	LUT2 #(
		.INIT('h1)
	) name16341 (
		_w16773_,
		_w16872_,
		_w16873_
	);
	LUT2 #(
		.INIT('h1)
	) name16342 (
		_w15625_,
		_w16289_,
		_w16874_
	);
	LUT2 #(
		.INIT('h4)
	) name16343 (
		\u0_w_reg[3][19]/P0001 ,
		_w15530_,
		_w16875_
	);
	LUT2 #(
		.INIT('h8)
	) name16344 (
		\u0_w_reg[3][20]/P0001 ,
		_w16875_,
		_w16876_
	);
	LUT2 #(
		.INIT('h2)
	) name16345 (
		_w16874_,
		_w16876_,
		_w16877_
	);
	LUT2 #(
		.INIT('h1)
	) name16346 (
		\u0_w_reg[3][18]/P0001 ,
		_w16877_,
		_w16878_
	);
	LUT2 #(
		.INIT('h1)
	) name16347 (
		_w15592_,
		_w16878_,
		_w16879_
	);
	LUT2 #(
		.INIT('h2)
	) name16348 (
		\u0_w_reg[3][17]/P0001 ,
		_w16879_,
		_w16880_
	);
	LUT2 #(
		.INIT('h1)
	) name16349 (
		_w15549_,
		_w16313_,
		_w16881_
	);
	LUT2 #(
		.INIT('h2)
	) name16350 (
		_w15608_,
		_w16881_,
		_w16882_
	);
	LUT2 #(
		.INIT('h4)
	) name16351 (
		_w15525_,
		_w15549_,
		_w16883_
	);
	LUT2 #(
		.INIT('h4)
	) name16352 (
		_w15613_,
		_w16883_,
		_w16884_
	);
	LUT2 #(
		.INIT('h8)
	) name16353 (
		_w15648_,
		_w16774_,
		_w16885_
	);
	LUT2 #(
		.INIT('h8)
	) name16354 (
		\u0_w_reg[3][18]/P0001 ,
		_w15527_,
		_w16886_
	);
	LUT2 #(
		.INIT('h1)
	) name16355 (
		_w15650_,
		_w16853_,
		_w16887_
	);
	LUT2 #(
		.INIT('h4)
	) name16356 (
		_w16249_,
		_w16887_,
		_w16888_
	);
	LUT2 #(
		.INIT('h1)
	) name16357 (
		\u0_w_reg[3][18]/P0001 ,
		_w16888_,
		_w16889_
	);
	LUT2 #(
		.INIT('h1)
	) name16358 (
		_w16884_,
		_w16885_,
		_w16890_
	);
	LUT2 #(
		.INIT('h4)
	) name16359 (
		_w16886_,
		_w16890_,
		_w16891_
	);
	LUT2 #(
		.INIT('h4)
	) name16360 (
		_w16882_,
		_w16891_,
		_w16892_
	);
	LUT2 #(
		.INIT('h4)
	) name16361 (
		_w16889_,
		_w16892_,
		_w16893_
	);
	LUT2 #(
		.INIT('h1)
	) name16362 (
		\u0_w_reg[3][17]/P0001 ,
		_w16893_,
		_w16894_
	);
	LUT2 #(
		.INIT('h8)
	) name16363 (
		_w15518_,
		_w16266_,
		_w16895_
	);
	LUT2 #(
		.INIT('h2)
	) name16364 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w16896_
	);
	LUT2 #(
		.INIT('h8)
	) name16365 (
		_w16895_,
		_w16896_,
		_w16897_
	);
	LUT2 #(
		.INIT('h1)
	) name16366 (
		_w15601_,
		_w16774_,
		_w16898_
	);
	LUT2 #(
		.INIT('h2)
	) name16367 (
		_w15507_,
		_w16898_,
		_w16899_
	);
	LUT2 #(
		.INIT('h1)
	) name16368 (
		_w15506_,
		_w16840_,
		_w16900_
	);
	LUT2 #(
		.INIT('h8)
	) name16369 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		_w16901_
	);
	LUT2 #(
		.INIT('h8)
	) name16370 (
		\u0_w_reg[3][23]/P0001 ,
		_w16901_,
		_w16902_
	);
	LUT2 #(
		.INIT('h4)
	) name16371 (
		_w16900_,
		_w16902_,
		_w16903_
	);
	LUT2 #(
		.INIT('h1)
	) name16372 (
		_w15606_,
		_w15618_,
		_w16904_
	);
	LUT2 #(
		.INIT('h4)
	) name16373 (
		_w15655_,
		_w16904_,
		_w16905_
	);
	LUT2 #(
		.INIT('h2)
	) name16374 (
		_w15608_,
		_w16905_,
		_w16906_
	);
	LUT2 #(
		.INIT('h1)
	) name16375 (
		_w15531_,
		_w16774_,
		_w16907_
	);
	LUT2 #(
		.INIT('h2)
	) name16376 (
		_w15506_,
		_w16907_,
		_w16908_
	);
	LUT2 #(
		.INIT('h8)
	) name16377 (
		_w15511_,
		_w15516_,
		_w16909_
	);
	LUT2 #(
		.INIT('h2)
	) name16378 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		_w16910_
	);
	LUT2 #(
		.INIT('h1)
	) name16379 (
		_w16261_,
		_w16309_,
		_w16911_
	);
	LUT2 #(
		.INIT('h2)
	) name16380 (
		_w16910_,
		_w16911_,
		_w16912_
	);
	LUT2 #(
		.INIT('h1)
	) name16381 (
		\u0_w_reg[3][21]/P0001 ,
		_w15588_,
		_w16913_
	);
	LUT2 #(
		.INIT('h2)
	) name16382 (
		_w15520_,
		_w16913_,
		_w16914_
	);
	LUT2 #(
		.INIT('h1)
	) name16383 (
		_w15543_,
		_w16914_,
		_w16915_
	);
	LUT2 #(
		.INIT('h1)
	) name16384 (
		\u0_w_reg[3][19]/P0001 ,
		_w16915_,
		_w16916_
	);
	LUT2 #(
		.INIT('h8)
	) name16385 (
		_w15503_,
		_w15511_,
		_w16917_
	);
	LUT2 #(
		.INIT('h8)
	) name16386 (
		_w16268_,
		_w16297_,
		_w16918_
	);
	LUT2 #(
		.INIT('h8)
	) name16387 (
		_w15504_,
		_w15590_,
		_w16919_
	);
	LUT2 #(
		.INIT('h1)
	) name16388 (
		\u0_w_reg[3][17]/P0001 ,
		_w16917_,
		_w16920_
	);
	LUT2 #(
		.INIT('h1)
	) name16389 (
		_w16918_,
		_w16919_,
		_w16921_
	);
	LUT2 #(
		.INIT('h8)
	) name16390 (
		_w16920_,
		_w16921_,
		_w16922_
	);
	LUT2 #(
		.INIT('h1)
	) name16391 (
		_w15647_,
		_w16777_,
		_w16923_
	);
	LUT2 #(
		.INIT('h8)
	) name16392 (
		_w16922_,
		_w16923_,
		_w16924_
	);
	LUT2 #(
		.INIT('h4)
	) name16393 (
		_w16916_,
		_w16924_,
		_w16925_
	);
	LUT2 #(
		.INIT('h8)
	) name16394 (
		_w15613_,
		_w16297_,
		_w16926_
	);
	LUT2 #(
		.INIT('h2)
	) name16395 (
		\u0_w_reg[3][17]/P0001 ,
		_w16926_,
		_w16927_
	);
	LUT2 #(
		.INIT('h4)
	) name16396 (
		_w16852_,
		_w16927_,
		_w16928_
	);
	LUT2 #(
		.INIT('h1)
	) name16397 (
		_w16925_,
		_w16928_,
		_w16929_
	);
	LUT2 #(
		.INIT('h2)
	) name16398 (
		\u0_w_reg[3][16]/P0001 ,
		_w16909_,
		_w16930_
	);
	LUT2 #(
		.INIT('h4)
	) name16399 (
		_w16908_,
		_w16930_,
		_w16931_
	);
	LUT2 #(
		.INIT('h4)
	) name16400 (
		_w16912_,
		_w16931_,
		_w16932_
	);
	LUT2 #(
		.INIT('h4)
	) name16401 (
		_w16906_,
		_w16932_,
		_w16933_
	);
	LUT2 #(
		.INIT('h4)
	) name16402 (
		_w16929_,
		_w16933_,
		_w16934_
	);
	LUT2 #(
		.INIT('h8)
	) name16403 (
		_w15529_,
		_w15542_,
		_w16935_
	);
	LUT2 #(
		.INIT('h1)
	) name16404 (
		\u0_w_reg[3][17]/P0001 ,
		_w15527_,
		_w16936_
	);
	LUT2 #(
		.INIT('h4)
	) name16405 (
		_w16935_,
		_w16936_,
		_w16937_
	);
	LUT2 #(
		.INIT('h1)
	) name16406 (
		_w15613_,
		_w16229_,
		_w16938_
	);
	LUT2 #(
		.INIT('h1)
	) name16407 (
		\u0_w_reg[3][18]/P0001 ,
		_w15542_,
		_w16939_
	);
	LUT2 #(
		.INIT('h4)
	) name16408 (
		_w16938_,
		_w16939_,
		_w16940_
	);
	LUT2 #(
		.INIT('h4)
	) name16409 (
		\u0_w_reg[3][19]/P0001 ,
		_w15520_,
		_w16941_
	);
	LUT2 #(
		.INIT('h1)
	) name16410 (
		_w15540_,
		_w16941_,
		_w16942_
	);
	LUT2 #(
		.INIT('h2)
	) name16411 (
		\u0_w_reg[3][18]/P0001 ,
		_w16942_,
		_w16943_
	);
	LUT2 #(
		.INIT('h8)
	) name16412 (
		\u0_w_reg[3][21]/P0001 ,
		_w15575_,
		_w16944_
	);
	LUT2 #(
		.INIT('h2)
	) name16413 (
		\u0_w_reg[3][17]/P0001 ,
		_w16944_,
		_w16945_
	);
	LUT2 #(
		.INIT('h1)
	) name16414 (
		_w16940_,
		_w16943_,
		_w16946_
	);
	LUT2 #(
		.INIT('h8)
	) name16415 (
		_w16945_,
		_w16946_,
		_w16947_
	);
	LUT2 #(
		.INIT('h1)
	) name16416 (
		_w16937_,
		_w16947_,
		_w16948_
	);
	LUT2 #(
		.INIT('h8)
	) name16417 (
		_w15602_,
		_w15608_,
		_w16949_
	);
	LUT2 #(
		.INIT('h8)
	) name16418 (
		\u0_w_reg[3][22]/P0001 ,
		_w16949_,
		_w16950_
	);
	LUT2 #(
		.INIT('h1)
	) name16419 (
		\u0_w_reg[3][16]/P0001 ,
		_w15628_,
		_w16951_
	);
	LUT2 #(
		.INIT('h4)
	) name16420 (
		_w15659_,
		_w16951_,
		_w16952_
	);
	LUT2 #(
		.INIT('h4)
	) name16421 (
		_w16950_,
		_w16952_,
		_w16953_
	);
	LUT2 #(
		.INIT('h4)
	) name16422 (
		_w16948_,
		_w16953_,
		_w16954_
	);
	LUT2 #(
		.INIT('h1)
	) name16423 (
		_w16934_,
		_w16954_,
		_w16955_
	);
	LUT2 #(
		.INIT('h1)
	) name16424 (
		_w16270_,
		_w16897_,
		_w16956_
	);
	LUT2 #(
		.INIT('h1)
	) name16425 (
		_w16899_,
		_w16903_,
		_w16957_
	);
	LUT2 #(
		.INIT('h8)
	) name16426 (
		_w16956_,
		_w16957_,
		_w16958_
	);
	LUT2 #(
		.INIT('h4)
	) name16427 (
		_w16880_,
		_w16958_,
		_w16959_
	);
	LUT2 #(
		.INIT('h4)
	) name16428 (
		_w16894_,
		_w16959_,
		_w16960_
	);
	LUT2 #(
		.INIT('h4)
	) name16429 (
		_w16955_,
		_w16960_,
		_w16961_
	);
	LUT2 #(
		.INIT('h2)
	) name16430 (
		\u0_w_reg[0][26]/P0001 ,
		_w16961_,
		_w16962_
	);
	LUT2 #(
		.INIT('h4)
	) name16431 (
		\u0_w_reg[0][26]/P0001 ,
		_w16961_,
		_w16963_
	);
	LUT2 #(
		.INIT('h1)
	) name16432 (
		_w16962_,
		_w16963_,
		_w16964_
	);
	LUT2 #(
		.INIT('h1)
	) name16433 (
		\u0_r0_out_reg[26]/P0001 ,
		_w16964_,
		_w16965_
	);
	LUT2 #(
		.INIT('h8)
	) name16434 (
		\u0_r0_out_reg[26]/P0001 ,
		_w16964_,
		_w16966_
	);
	LUT2 #(
		.INIT('h1)
	) name16435 (
		ld_pad,
		_w16965_,
		_w16967_
	);
	LUT2 #(
		.INIT('h4)
	) name16436 (
		_w16966_,
		_w16967_,
		_w16968_
	);
	LUT2 #(
		.INIT('h8)
	) name16437 (
		\key[122]_pad ,
		ld_pad,
		_w16969_
	);
	LUT2 #(
		.INIT('h1)
	) name16438 (
		_w16968_,
		_w16969_,
		_w16970_
	);
	LUT2 #(
		.INIT('h4)
	) name16439 (
		_w15539_,
		_w15660_,
		_w16971_
	);
	LUT2 #(
		.INIT('h4)
	) name16440 (
		\u0_w_reg[3][20]/P0001 ,
		_w15592_,
		_w16972_
	);
	LUT2 #(
		.INIT('h1)
	) name16441 (
		_w15583_,
		_w16854_,
		_w16973_
	);
	LUT2 #(
		.INIT('h4)
	) name16442 (
		_w16972_,
		_w16973_,
		_w16974_
	);
	LUT2 #(
		.INIT('h2)
	) name16443 (
		\u0_w_reg[3][18]/P0001 ,
		_w16974_,
		_w16975_
	);
	LUT2 #(
		.INIT('h2)
	) name16444 (
		_w16803_,
		_w16971_,
		_w16976_
	);
	LUT2 #(
		.INIT('h4)
	) name16445 (
		_w16975_,
		_w16976_,
		_w16977_
	);
	LUT2 #(
		.INIT('h2)
	) name16446 (
		\u0_w_reg[3][17]/P0001 ,
		_w16977_,
		_w16978_
	);
	LUT2 #(
		.INIT('h1)
	) name16447 (
		_w15576_,
		_w16851_,
		_w16979_
	);
	LUT2 #(
		.INIT('h1)
	) name16448 (
		\u0_w_reg[3][18]/P0001 ,
		_w16979_,
		_w16980_
	);
	LUT2 #(
		.INIT('h1)
	) name16449 (
		_w15630_,
		_w16217_,
		_w16981_
	);
	LUT2 #(
		.INIT('h8)
	) name16450 (
		_w16306_,
		_w16981_,
		_w16982_
	);
	LUT2 #(
		.INIT('h2)
	) name16451 (
		\u0_w_reg[3][18]/P0001 ,
		_w16982_,
		_w16983_
	);
	LUT2 #(
		.INIT('h1)
	) name16452 (
		_w15638_,
		_w16248_,
		_w16984_
	);
	LUT2 #(
		.INIT('h2)
	) name16453 (
		\u0_w_reg[3][18]/P0001 ,
		_w16984_,
		_w16985_
	);
	LUT2 #(
		.INIT('h1)
	) name16454 (
		_w15628_,
		_w16885_,
		_w16986_
	);
	LUT2 #(
		.INIT('h4)
	) name16455 (
		_w16985_,
		_w16986_,
		_w16987_
	);
	LUT2 #(
		.INIT('h4)
	) name16456 (
		_w15627_,
		_w16987_,
		_w16988_
	);
	LUT2 #(
		.INIT('h1)
	) name16457 (
		\u0_w_reg[3][17]/P0001 ,
		_w16988_,
		_w16989_
	);
	LUT2 #(
		.INIT('h1)
	) name16458 (
		_w16980_,
		_w16983_,
		_w16990_
	);
	LUT2 #(
		.INIT('h4)
	) name16459 (
		_w16989_,
		_w16990_,
		_w16991_
	);
	LUT2 #(
		.INIT('h4)
	) name16460 (
		_w16978_,
		_w16991_,
		_w16992_
	);
	LUT2 #(
		.INIT('h2)
	) name16461 (
		\u0_w_reg[3][16]/P0001 ,
		_w16992_,
		_w16993_
	);
	LUT2 #(
		.INIT('h4)
	) name16462 (
		\u0_w_reg[3][19]/P0001 ,
		_w16261_,
		_w16994_
	);
	LUT2 #(
		.INIT('h4)
	) name16463 (
		_w15520_,
		_w15662_,
		_w16995_
	);
	LUT2 #(
		.INIT('h1)
	) name16464 (
		_w16230_,
		_w16310_,
		_w16996_
	);
	LUT2 #(
		.INIT('h1)
	) name16465 (
		_w16994_,
		_w16995_,
		_w16997_
	);
	LUT2 #(
		.INIT('h8)
	) name16466 (
		_w16996_,
		_w16997_,
		_w16998_
	);
	LUT2 #(
		.INIT('h1)
	) name16467 (
		\u0_w_reg[3][18]/P0001 ,
		_w16998_,
		_w16999_
	);
	LUT2 #(
		.INIT('h4)
	) name16468 (
		\u0_w_reg[3][20]/P0001 ,
		_w16875_,
		_w17000_
	);
	LUT2 #(
		.INIT('h1)
	) name16469 (
		_w15504_,
		_w16309_,
		_w17001_
	);
	LUT2 #(
		.INIT('h2)
	) name16470 (
		_w15601_,
		_w17001_,
		_w17002_
	);
	LUT2 #(
		.INIT('h8)
	) name16471 (
		_w15608_,
		_w16774_,
		_w17003_
	);
	LUT2 #(
		.INIT('h1)
	) name16472 (
		\u0_w_reg[3][17]/P0001 ,
		_w16836_,
		_w17004_
	);
	LUT2 #(
		.INIT('h4)
	) name16473 (
		_w16851_,
		_w17004_,
		_w17005_
	);
	LUT2 #(
		.INIT('h1)
	) name16474 (
		_w17000_,
		_w17003_,
		_w17006_
	);
	LUT2 #(
		.INIT('h8)
	) name16475 (
		_w17005_,
		_w17006_,
		_w17007_
	);
	LUT2 #(
		.INIT('h4)
	) name16476 (
		_w17002_,
		_w17007_,
		_w17008_
	);
	LUT2 #(
		.INIT('h2)
	) name16477 (
		_w15511_,
		_w15616_,
		_w17009_
	);
	LUT2 #(
		.INIT('h4)
	) name16478 (
		\u0_w_reg[3][18]/P0001 ,
		_w15630_,
		_w17010_
	);
	LUT2 #(
		.INIT('h2)
	) name16479 (
		\u0_w_reg[3][17]/P0001 ,
		_w15650_,
		_w17011_
	);
	LUT2 #(
		.INIT('h4)
	) name16480 (
		_w17010_,
		_w17011_,
		_w17012_
	);
	LUT2 #(
		.INIT('h4)
	) name16481 (
		_w17009_,
		_w17012_,
		_w17013_
	);
	LUT2 #(
		.INIT('h1)
	) name16482 (
		_w17008_,
		_w17013_,
		_w17014_
	);
	LUT2 #(
		.INIT('h1)
	) name16483 (
		_w16999_,
		_w17014_,
		_w17015_
	);
	LUT2 #(
		.INIT('h1)
	) name16484 (
		\u0_w_reg[3][16]/P0001 ,
		_w17015_,
		_w17016_
	);
	LUT2 #(
		.INIT('h8)
	) name16485 (
		_w15520_,
		_w16266_,
		_w17017_
	);
	LUT2 #(
		.INIT('h4)
	) name16486 (
		\u0_w_reg[3][18]/P0001 ,
		_w15618_,
		_w17018_
	);
	LUT2 #(
		.INIT('h8)
	) name16487 (
		\u0_w_reg[3][18]/P0001 ,
		_w16313_,
		_w17019_
	);
	LUT2 #(
		.INIT('h8)
	) name16488 (
		\u0_w_reg[3][21]/P0001 ,
		_w15530_,
		_w17020_
	);
	LUT2 #(
		.INIT('h8)
	) name16489 (
		_w15529_,
		_w17020_,
		_w17021_
	);
	LUT2 #(
		.INIT('h1)
	) name16490 (
		_w15580_,
		_w15629_,
		_w17022_
	);
	LUT2 #(
		.INIT('h1)
	) name16491 (
		_w16249_,
		_w17017_,
		_w17023_
	);
	LUT2 #(
		.INIT('h1)
	) name16492 (
		_w17018_,
		_w17019_,
		_w17024_
	);
	LUT2 #(
		.INIT('h4)
	) name16493 (
		_w17021_,
		_w17024_,
		_w17025_
	);
	LUT2 #(
		.INIT('h8)
	) name16494 (
		_w17022_,
		_w17023_,
		_w17026_
	);
	LUT2 #(
		.INIT('h8)
	) name16495 (
		_w17025_,
		_w17026_,
		_w17027_
	);
	LUT2 #(
		.INIT('h1)
	) name16496 (
		\u0_w_reg[3][17]/P0001 ,
		_w17027_,
		_w17028_
	);
	LUT2 #(
		.INIT('h8)
	) name16497 (
		\u0_w_reg[3][17]/P0001 ,
		_w15659_,
		_w17029_
	);
	LUT2 #(
		.INIT('h1)
	) name16498 (
		_w15600_,
		_w15630_,
		_w17030_
	);
	LUT2 #(
		.INIT('h1)
	) name16499 (
		\u0_w_reg[3][19]/P0001 ,
		_w17030_,
		_w17031_
	);
	LUT2 #(
		.INIT('h8)
	) name16500 (
		_w15525_,
		_w15591_,
		_w17032_
	);
	LUT2 #(
		.INIT('h1)
	) name16501 (
		_w16795_,
		_w17032_,
		_w17033_
	);
	LUT2 #(
		.INIT('h1)
	) name16502 (
		\u0_w_reg[3][16]/P0001 ,
		_w17033_,
		_w17034_
	);
	LUT2 #(
		.INIT('h8)
	) name16503 (
		_w15504_,
		_w17020_,
		_w17035_
	);
	LUT2 #(
		.INIT('h1)
	) name16504 (
		_w15637_,
		_w16284_,
		_w17036_
	);
	LUT2 #(
		.INIT('h4)
	) name16505 (
		_w17035_,
		_w17036_,
		_w17037_
	);
	LUT2 #(
		.INIT('h2)
	) name16506 (
		\u0_w_reg[3][17]/P0001 ,
		_w17037_,
		_w17038_
	);
	LUT2 #(
		.INIT('h1)
	) name16507 (
		_w16288_,
		_w17034_,
		_w17039_
	);
	LUT2 #(
		.INIT('h4)
	) name16508 (
		_w17038_,
		_w17039_,
		_w17040_
	);
	LUT2 #(
		.INIT('h2)
	) name16509 (
		\u0_w_reg[3][18]/P0001 ,
		_w17040_,
		_w17041_
	);
	LUT2 #(
		.INIT('h1)
	) name16510 (
		_w16300_,
		_w17029_,
		_w17042_
	);
	LUT2 #(
		.INIT('h4)
	) name16511 (
		_w17031_,
		_w17042_,
		_w17043_
	);
	LUT2 #(
		.INIT('h4)
	) name16512 (
		_w17028_,
		_w17043_,
		_w17044_
	);
	LUT2 #(
		.INIT('h4)
	) name16513 (
		_w17041_,
		_w17044_,
		_w17045_
	);
	LUT2 #(
		.INIT('h4)
	) name16514 (
		_w17016_,
		_w17045_,
		_w17046_
	);
	LUT2 #(
		.INIT('h4)
	) name16515 (
		_w16993_,
		_w17046_,
		_w17047_
	);
	LUT2 #(
		.INIT('h2)
	) name16516 (
		\u0_r0_out_reg[30]/P0001 ,
		_w17047_,
		_w17048_
	);
	LUT2 #(
		.INIT('h4)
	) name16517 (
		\u0_r0_out_reg[30]/P0001 ,
		_w17047_,
		_w17049_
	);
	LUT2 #(
		.INIT('h1)
	) name16518 (
		_w17048_,
		_w17049_,
		_w17050_
	);
	LUT2 #(
		.INIT('h1)
	) name16519 (
		\u0_w_reg[0][30]/P0001 ,
		_w17050_,
		_w17051_
	);
	LUT2 #(
		.INIT('h8)
	) name16520 (
		\u0_w_reg[0][30]/P0001 ,
		_w17050_,
		_w17052_
	);
	LUT2 #(
		.INIT('h1)
	) name16521 (
		ld_pad,
		_w17051_,
		_w17053_
	);
	LUT2 #(
		.INIT('h4)
	) name16522 (
		_w17052_,
		_w17053_,
		_w17054_
	);
	LUT2 #(
		.INIT('h8)
	) name16523 (
		\key[126]_pad ,
		ld_pad,
		_w17055_
	);
	LUT2 #(
		.INIT('h1)
	) name16524 (
		_w17054_,
		_w17055_,
		_w17056_
	);
	LUT2 #(
		.INIT('h1)
	) name16525 (
		_w15543_,
		_w15606_,
		_w17057_
	);
	LUT2 #(
		.INIT('h2)
	) name16526 (
		_w15648_,
		_w17057_,
		_w17058_
	);
	LUT2 #(
		.INIT('h8)
	) name16527 (
		_w15518_,
		_w15537_,
		_w17059_
	);
	LUT2 #(
		.INIT('h1)
	) name16528 (
		_w15562_,
		_w17059_,
		_w17060_
	);
	LUT2 #(
		.INIT('h1)
	) name16529 (
		\u0_w_reg[3][18]/P0001 ,
		_w17060_,
		_w17061_
	);
	LUT2 #(
		.INIT('h1)
	) name16530 (
		_w16841_,
		_w17032_,
		_w17062_
	);
	LUT2 #(
		.INIT('h8)
	) name16531 (
		_w16945_,
		_w17062_,
		_w17063_
	);
	LUT2 #(
		.INIT('h4)
	) name16532 (
		_w17061_,
		_w17063_,
		_w17064_
	);
	LUT2 #(
		.INIT('h1)
	) name16533 (
		\u0_w_reg[3][17]/P0001 ,
		_w15600_,
		_w17065_
	);
	LUT2 #(
		.INIT('h1)
	) name16534 (
		_w16802_,
		_w16949_,
		_w17066_
	);
	LUT2 #(
		.INIT('h8)
	) name16535 (
		_w17065_,
		_w17066_,
		_w17067_
	);
	LUT2 #(
		.INIT('h1)
	) name16536 (
		_w17064_,
		_w17067_,
		_w17068_
	);
	LUT2 #(
		.INIT('h1)
	) name16537 (
		_w15663_,
		_w16289_,
		_w17069_
	);
	LUT2 #(
		.INIT('h2)
	) name16538 (
		\u0_w_reg[3][18]/P0001 ,
		_w17069_,
		_w17070_
	);
	LUT2 #(
		.INIT('h4)
	) name16539 (
		\u0_w_reg[3][17]/P0001 ,
		_w16268_,
		_w17071_
	);
	LUT2 #(
		.INIT('h1)
	) name16540 (
		_w16284_,
		_w17071_,
		_w17072_
	);
	LUT2 #(
		.INIT('h1)
	) name16541 (
		\u0_w_reg[3][18]/P0001 ,
		_w17072_,
		_w17073_
	);
	LUT2 #(
		.INIT('h1)
	) name16542 (
		_w15651_,
		_w15656_,
		_w17074_
	);
	LUT2 #(
		.INIT('h1)
	) name16543 (
		_w17058_,
		_w17073_,
		_w17075_
	);
	LUT2 #(
		.INIT('h8)
	) name16544 (
		_w17074_,
		_w17075_,
		_w17076_
	);
	LUT2 #(
		.INIT('h4)
	) name16545 (
		_w17070_,
		_w17076_,
		_w17077_
	);
	LUT2 #(
		.INIT('h4)
	) name16546 (
		_w17068_,
		_w17077_,
		_w17078_
	);
	LUT2 #(
		.INIT('h1)
	) name16547 (
		\u0_w_reg[3][16]/P0001 ,
		_w17078_,
		_w17079_
	);
	LUT2 #(
		.INIT('h4)
	) name16548 (
		\u0_w_reg[3][21]/P0001 ,
		_w15522_,
		_w17080_
	);
	LUT2 #(
		.INIT('h1)
	) name16549 (
		_w15581_,
		_w17080_,
		_w17081_
	);
	LUT2 #(
		.INIT('h1)
	) name16550 (
		\u0_w_reg[3][18]/P0001 ,
		_w17081_,
		_w17082_
	);
	LUT2 #(
		.INIT('h8)
	) name16551 (
		_w15518_,
		_w16248_,
		_w17083_
	);
	LUT2 #(
		.INIT('h8)
	) name16552 (
		\u0_w_reg[3][21]/P0001 ,
		_w16309_,
		_w17084_
	);
	LUT2 #(
		.INIT('h1)
	) name16553 (
		_w15584_,
		_w17083_,
		_w17085_
	);
	LUT2 #(
		.INIT('h4)
	) name16554 (
		_w17084_,
		_w17085_,
		_w17086_
	);
	LUT2 #(
		.INIT('h2)
	) name16555 (
		_w16281_,
		_w17086_,
		_w17087_
	);
	LUT2 #(
		.INIT('h8)
	) name16556 (
		\u0_w_reg[3][20]/P0001 ,
		_w16233_,
		_w17088_
	);
	LUT2 #(
		.INIT('h8)
	) name16557 (
		\u0_w_reg[3][20]/P0001 ,
		_w15559_,
		_w17089_
	);
	LUT2 #(
		.INIT('h8)
	) name16558 (
		\u0_w_reg[3][23]/P0001 ,
		_w15539_,
		_w17090_
	);
	LUT2 #(
		.INIT('h1)
	) name16559 (
		_w17089_,
		_w17090_,
		_w17091_
	);
	LUT2 #(
		.INIT('h2)
	) name16560 (
		_w15511_,
		_w17091_,
		_w17092_
	);
	LUT2 #(
		.INIT('h1)
	) name16561 (
		_w15586_,
		_w16807_,
		_w17093_
	);
	LUT2 #(
		.INIT('h1)
	) name16562 (
		_w16895_,
		_w17088_,
		_w17094_
	);
	LUT2 #(
		.INIT('h8)
	) name16563 (
		_w17093_,
		_w17094_,
		_w17095_
	);
	LUT2 #(
		.INIT('h4)
	) name16564 (
		_w17092_,
		_w17095_,
		_w17096_
	);
	LUT2 #(
		.INIT('h1)
	) name16565 (
		_w15525_,
		_w15648_,
		_w17097_
	);
	LUT2 #(
		.INIT('h2)
	) name16566 (
		\u0_w_reg[3][22]/P0001 ,
		_w17097_,
		_w17098_
	);
	LUT2 #(
		.INIT('h1)
	) name16567 (
		_w16827_,
		_w17098_,
		_w17099_
	);
	LUT2 #(
		.INIT('h1)
	) name16568 (
		\u0_w_reg[3][23]/P0001 ,
		_w17099_,
		_w17100_
	);
	LUT2 #(
		.INIT('h8)
	) name16569 (
		\u0_w_reg[3][23]/P0001 ,
		_w15508_,
		_w17101_
	);
	LUT2 #(
		.INIT('h1)
	) name16570 (
		_w15513_,
		_w16261_,
		_w17102_
	);
	LUT2 #(
		.INIT('h4)
	) name16571 (
		_w16854_,
		_w17102_,
		_w17103_
	);
	LUT2 #(
		.INIT('h1)
	) name16572 (
		\u0_w_reg[3][18]/P0001 ,
		_w17103_,
		_w17104_
	);
	LUT2 #(
		.INIT('h1)
	) name16573 (
		_w15657_,
		_w17101_,
		_w17105_
	);
	LUT2 #(
		.INIT('h4)
	) name16574 (
		_w17100_,
		_w17105_,
		_w17106_
	);
	LUT2 #(
		.INIT('h4)
	) name16575 (
		_w17104_,
		_w17106_,
		_w17107_
	);
	LUT2 #(
		.INIT('h8)
	) name16576 (
		_w17096_,
		_w17107_,
		_w17108_
	);
	LUT2 #(
		.INIT('h2)
	) name16577 (
		\u0_w_reg[3][16]/P0001 ,
		_w17108_,
		_w17109_
	);
	LUT2 #(
		.INIT('h4)
	) name16578 (
		\u0_w_reg[3][20]/P0001 ,
		_w15601_,
		_w17110_
	);
	LUT2 #(
		.INIT('h8)
	) name16579 (
		_w15529_,
		_w17110_,
		_w17111_
	);
	LUT2 #(
		.INIT('h2)
	) name16580 (
		_w16936_,
		_w17111_,
		_w17112_
	);
	LUT2 #(
		.INIT('h4)
	) name16581 (
		_w17058_,
		_w17112_,
		_w17113_
	);
	LUT2 #(
		.INIT('h4)
	) name16582 (
		_w17109_,
		_w17113_,
		_w17114_
	);
	LUT2 #(
		.INIT('h1)
	) name16583 (
		_w15539_,
		_w16261_,
		_w17115_
	);
	LUT2 #(
		.INIT('h8)
	) name16584 (
		\u0_w_reg[3][19]/P0001 ,
		_w15503_,
		_w17116_
	);
	LUT2 #(
		.INIT('h1)
	) name16585 (
		_w16941_,
		_w17116_,
		_w17117_
	);
	LUT2 #(
		.INIT('h8)
	) name16586 (
		_w17115_,
		_w17117_,
		_w17118_
	);
	LUT2 #(
		.INIT('h2)
	) name16587 (
		\u0_w_reg[3][18]/P0001 ,
		_w17118_,
		_w17119_
	);
	LUT2 #(
		.INIT('h1)
	) name16588 (
		_w16820_,
		_w17083_,
		_w17120_
	);
	LUT2 #(
		.INIT('h4)
	) name16589 (
		_w17119_,
		_w17120_,
		_w17121_
	);
	LUT2 #(
		.INIT('h8)
	) name16590 (
		_w17096_,
		_w17121_,
		_w17122_
	);
	LUT2 #(
		.INIT('h2)
	) name16591 (
		\u0_w_reg[3][16]/P0001 ,
		_w17122_,
		_w17123_
	);
	LUT2 #(
		.INIT('h2)
	) name16592 (
		_w15559_,
		_w16268_,
		_w17124_
	);
	LUT2 #(
		.INIT('h2)
	) name16593 (
		_w16786_,
		_w17124_,
		_w17125_
	);
	LUT2 #(
		.INIT('h2)
	) name16594 (
		\u0_w_reg[3][19]/P0001 ,
		_w17125_,
		_w17126_
	);
	LUT2 #(
		.INIT('h1)
	) name16595 (
		\u0_w_reg[3][18]/P0001 ,
		_w17126_,
		_w17127_
	);
	LUT2 #(
		.INIT('h2)
	) name16596 (
		\u0_w_reg[3][23]/P0001 ,
		_w17115_,
		_w17128_
	);
	LUT2 #(
		.INIT('h1)
	) name16597 (
		_w16853_,
		_w17128_,
		_w17129_
	);
	LUT2 #(
		.INIT('h1)
	) name16598 (
		\u0_w_reg[3][19]/P0001 ,
		_w17129_,
		_w17130_
	);
	LUT2 #(
		.INIT('h2)
	) name16599 (
		\u0_w_reg[3][18]/P0001 ,
		_w15538_,
		_w17131_
	);
	LUT2 #(
		.INIT('h4)
	) name16600 (
		_w15625_,
		_w17131_,
		_w17132_
	);
	LUT2 #(
		.INIT('h4)
	) name16601 (
		_w17130_,
		_w17132_,
		_w17133_
	);
	LUT2 #(
		.INIT('h1)
	) name16602 (
		_w17127_,
		_w17133_,
		_w17134_
	);
	LUT2 #(
		.INIT('h2)
	) name16603 (
		\u0_w_reg[3][17]/P0001 ,
		_w17123_,
		_w17135_
	);
	LUT2 #(
		.INIT('h4)
	) name16604 (
		_w17134_,
		_w17135_,
		_w17136_
	);
	LUT2 #(
		.INIT('h1)
	) name16605 (
		_w17114_,
		_w17136_,
		_w17137_
	);
	LUT2 #(
		.INIT('h1)
	) name16606 (
		_w17082_,
		_w17087_,
		_w17138_
	);
	LUT2 #(
		.INIT('h4)
	) name16607 (
		_w17079_,
		_w17138_,
		_w17139_
	);
	LUT2 #(
		.INIT('h4)
	) name16608 (
		_w17137_,
		_w17139_,
		_w17140_
	);
	LUT2 #(
		.INIT('h2)
	) name16609 (
		\u0_w_reg[0][31]/P0001 ,
		_w17140_,
		_w17141_
	);
	LUT2 #(
		.INIT('h4)
	) name16610 (
		\u0_w_reg[0][31]/P0001 ,
		_w17140_,
		_w17142_
	);
	LUT2 #(
		.INIT('h1)
	) name16611 (
		_w17141_,
		_w17142_,
		_w17143_
	);
	LUT2 #(
		.INIT('h1)
	) name16612 (
		\u0_r0_out_reg[31]/P0001 ,
		_w17143_,
		_w17144_
	);
	LUT2 #(
		.INIT('h8)
	) name16613 (
		\u0_r0_out_reg[31]/P0001 ,
		_w17143_,
		_w17145_
	);
	LUT2 #(
		.INIT('h1)
	) name16614 (
		ld_pad,
		_w17144_,
		_w17146_
	);
	LUT2 #(
		.INIT('h4)
	) name16615 (
		_w17145_,
		_w17146_,
		_w17147_
	);
	LUT2 #(
		.INIT('h8)
	) name16616 (
		\key[127]_pad ,
		ld_pad,
		_w17148_
	);
	LUT2 #(
		.INIT('h1)
	) name16617 (
		_w17147_,
		_w17148_,
		_w17149_
	);
	LUT2 #(
		.INIT('h2)
	) name16618 (
		\u0_r0_out_reg[26]/P0001 ,
		\u0_w_reg[1][26]/P0001 ,
		_w17150_
	);
	LUT2 #(
		.INIT('h4)
	) name16619 (
		\u0_r0_out_reg[26]/P0001 ,
		\u0_w_reg[1][26]/P0001 ,
		_w17151_
	);
	LUT2 #(
		.INIT('h1)
	) name16620 (
		_w17150_,
		_w17151_,
		_w17152_
	);
	LUT2 #(
		.INIT('h4)
	) name16621 (
		_w16964_,
		_w17152_,
		_w17153_
	);
	LUT2 #(
		.INIT('h2)
	) name16622 (
		_w16964_,
		_w17152_,
		_w17154_
	);
	LUT2 #(
		.INIT('h1)
	) name16623 (
		ld_pad,
		_w17153_,
		_w17155_
	);
	LUT2 #(
		.INIT('h4)
	) name16624 (
		_w17154_,
		_w17155_,
		_w17156_
	);
	LUT2 #(
		.INIT('h8)
	) name16625 (
		\key[90]_pad ,
		ld_pad,
		_w17157_
	);
	LUT2 #(
		.INIT('h1)
	) name16626 (
		_w17156_,
		_w17157_,
		_w17158_
	);
	LUT2 #(
		.INIT('h2)
	) name16627 (
		\u0_w_reg[0][30]/P0001 ,
		\u0_w_reg[1][30]/P0001 ,
		_w17159_
	);
	LUT2 #(
		.INIT('h4)
	) name16628 (
		\u0_w_reg[0][30]/P0001 ,
		\u0_w_reg[1][30]/P0001 ,
		_w17160_
	);
	LUT2 #(
		.INIT('h1)
	) name16629 (
		_w17159_,
		_w17160_,
		_w17161_
	);
	LUT2 #(
		.INIT('h4)
	) name16630 (
		_w17050_,
		_w17161_,
		_w17162_
	);
	LUT2 #(
		.INIT('h2)
	) name16631 (
		_w17050_,
		_w17161_,
		_w17163_
	);
	LUT2 #(
		.INIT('h1)
	) name16632 (
		ld_pad,
		_w17162_,
		_w17164_
	);
	LUT2 #(
		.INIT('h4)
	) name16633 (
		_w17163_,
		_w17164_,
		_w17165_
	);
	LUT2 #(
		.INIT('h8)
	) name16634 (
		\key[94]_pad ,
		ld_pad,
		_w17166_
	);
	LUT2 #(
		.INIT('h1)
	) name16635 (
		_w17165_,
		_w17166_,
		_w17167_
	);
	LUT2 #(
		.INIT('h2)
	) name16636 (
		\u0_r0_out_reg[31]/P0001 ,
		\u0_w_reg[1][31]/P0001 ,
		_w17168_
	);
	LUT2 #(
		.INIT('h4)
	) name16637 (
		\u0_r0_out_reg[31]/P0001 ,
		\u0_w_reg[1][31]/P0001 ,
		_w17169_
	);
	LUT2 #(
		.INIT('h1)
	) name16638 (
		_w17168_,
		_w17169_,
		_w17170_
	);
	LUT2 #(
		.INIT('h4)
	) name16639 (
		_w17143_,
		_w17170_,
		_w17171_
	);
	LUT2 #(
		.INIT('h2)
	) name16640 (
		_w17143_,
		_w17170_,
		_w17172_
	);
	LUT2 #(
		.INIT('h1)
	) name16641 (
		ld_pad,
		_w17171_,
		_w17173_
	);
	LUT2 #(
		.INIT('h4)
	) name16642 (
		_w17172_,
		_w17173_,
		_w17174_
	);
	LUT2 #(
		.INIT('h8)
	) name16643 (
		\key[95]_pad ,
		ld_pad,
		_w17175_
	);
	LUT2 #(
		.INIT('h1)
	) name16644 (
		_w17174_,
		_w17175_,
		_w17176_
	);
	LUT2 #(
		.INIT('h8)
	) name16645 (
		\key[56]_pad ,
		ld_pad,
		_w17177_
	);
	LUT2 #(
		.INIT('h2)
	) name16646 (
		\u0_w_reg[1][24]/P0002 ,
		\u0_w_reg[2][24]/P0001 ,
		_w17178_
	);
	LUT2 #(
		.INIT('h4)
	) name16647 (
		\u0_w_reg[1][24]/P0002 ,
		\u0_w_reg[2][24]/P0001 ,
		_w17179_
	);
	LUT2 #(
		.INIT('h1)
	) name16648 (
		_w17178_,
		_w17179_,
		_w17180_
	);
	LUT2 #(
		.INIT('h4)
	) name16649 (
		_w16868_,
		_w17180_,
		_w17181_
	);
	LUT2 #(
		.INIT('h2)
	) name16650 (
		_w16868_,
		_w17180_,
		_w17182_
	);
	LUT2 #(
		.INIT('h1)
	) name16651 (
		_w17181_,
		_w17182_,
		_w17183_
	);
	LUT2 #(
		.INIT('h8)
	) name16652 (
		_w16865_,
		_w17183_,
		_w17184_
	);
	LUT2 #(
		.INIT('h1)
	) name16653 (
		_w16865_,
		_w17183_,
		_w17185_
	);
	LUT2 #(
		.INIT('h1)
	) name16654 (
		ld_pad,
		_w17184_,
		_w17186_
	);
	LUT2 #(
		.INIT('h4)
	) name16655 (
		_w17185_,
		_w17186_,
		_w17187_
	);
	LUT2 #(
		.INIT('h1)
	) name16656 (
		_w17177_,
		_w17187_,
		_w17188_
	);
	LUT2 #(
		.INIT('h4)
	) name16657 (
		\key[58]_pad ,
		ld_pad,
		_w17189_
	);
	LUT2 #(
		.INIT('h8)
	) name16658 (
		\u0_w_reg[2][26]/P0001 ,
		_w17152_,
		_w17190_
	);
	LUT2 #(
		.INIT('h1)
	) name16659 (
		\u0_w_reg[2][26]/P0001 ,
		_w17152_,
		_w17191_
	);
	LUT2 #(
		.INIT('h1)
	) name16660 (
		_w17190_,
		_w17191_,
		_w17192_
	);
	LUT2 #(
		.INIT('h8)
	) name16661 (
		_w16964_,
		_w17192_,
		_w17193_
	);
	LUT2 #(
		.INIT('h1)
	) name16662 (
		_w16964_,
		_w17192_,
		_w17194_
	);
	LUT2 #(
		.INIT('h1)
	) name16663 (
		_w17193_,
		_w17194_,
		_w17195_
	);
	LUT2 #(
		.INIT('h4)
	) name16664 (
		ld_pad,
		_w17195_,
		_w17196_
	);
	LUT2 #(
		.INIT('h1)
	) name16665 (
		_w17189_,
		_w17196_,
		_w17197_
	);
	LUT2 #(
		.INIT('h4)
	) name16666 (
		\key[62]_pad ,
		ld_pad,
		_w17198_
	);
	LUT2 #(
		.INIT('h8)
	) name16667 (
		\u0_w_reg[2][30]/P0001 ,
		_w17161_,
		_w17199_
	);
	LUT2 #(
		.INIT('h1)
	) name16668 (
		\u0_w_reg[2][30]/P0001 ,
		_w17161_,
		_w17200_
	);
	LUT2 #(
		.INIT('h1)
	) name16669 (
		_w17199_,
		_w17200_,
		_w17201_
	);
	LUT2 #(
		.INIT('h8)
	) name16670 (
		_w17050_,
		_w17201_,
		_w17202_
	);
	LUT2 #(
		.INIT('h1)
	) name16671 (
		_w17050_,
		_w17201_,
		_w17203_
	);
	LUT2 #(
		.INIT('h1)
	) name16672 (
		_w17202_,
		_w17203_,
		_w17204_
	);
	LUT2 #(
		.INIT('h4)
	) name16673 (
		ld_pad,
		_w17204_,
		_w17205_
	);
	LUT2 #(
		.INIT('h1)
	) name16674 (
		_w17198_,
		_w17205_,
		_w17206_
	);
	LUT2 #(
		.INIT('h4)
	) name16675 (
		\key[63]_pad ,
		ld_pad,
		_w17207_
	);
	LUT2 #(
		.INIT('h8)
	) name16676 (
		\u0_w_reg[2][31]/P0001 ,
		_w17170_,
		_w17208_
	);
	LUT2 #(
		.INIT('h1)
	) name16677 (
		\u0_w_reg[2][31]/P0001 ,
		_w17170_,
		_w17209_
	);
	LUT2 #(
		.INIT('h1)
	) name16678 (
		_w17208_,
		_w17209_,
		_w17210_
	);
	LUT2 #(
		.INIT('h8)
	) name16679 (
		_w17143_,
		_w17210_,
		_w17211_
	);
	LUT2 #(
		.INIT('h1)
	) name16680 (
		_w17143_,
		_w17210_,
		_w17212_
	);
	LUT2 #(
		.INIT('h1)
	) name16681 (
		_w17211_,
		_w17212_,
		_w17213_
	);
	LUT2 #(
		.INIT('h4)
	) name16682 (
		ld_pad,
		_w17213_,
		_w17214_
	);
	LUT2 #(
		.INIT('h1)
	) name16683 (
		_w17207_,
		_w17214_,
		_w17215_
	);
	LUT2 #(
		.INIT('h8)
	) name16684 (
		\key[24]_pad ,
		ld_pad,
		_w17216_
	);
	LUT2 #(
		.INIT('h1)
	) name16685 (
		\u0_w_reg[3][24]/P0001 ,
		_w16871_,
		_w17217_
	);
	LUT2 #(
		.INIT('h8)
	) name16686 (
		\u0_w_reg[3][24]/P0001 ,
		_w16871_,
		_w17218_
	);
	LUT2 #(
		.INIT('h1)
	) name16687 (
		_w17217_,
		_w17218_,
		_w17219_
	);
	LUT2 #(
		.INIT('h2)
	) name16688 (
		_w17180_,
		_w17219_,
		_w17220_
	);
	LUT2 #(
		.INIT('h4)
	) name16689 (
		_w17180_,
		_w17219_,
		_w17221_
	);
	LUT2 #(
		.INIT('h1)
	) name16690 (
		ld_pad,
		_w17220_,
		_w17222_
	);
	LUT2 #(
		.INIT('h4)
	) name16691 (
		_w17221_,
		_w17222_,
		_w17223_
	);
	LUT2 #(
		.INIT('h1)
	) name16692 (
		_w17216_,
		_w17223_,
		_w17224_
	);
	LUT2 #(
		.INIT('h4)
	) name16693 (
		\u0_w_reg[3][26]/P0001 ,
		_w17195_,
		_w17225_
	);
	LUT2 #(
		.INIT('h2)
	) name16694 (
		\u0_w_reg[3][26]/P0001 ,
		_w17195_,
		_w17226_
	);
	LUT2 #(
		.INIT('h1)
	) name16695 (
		ld_pad,
		_w17225_,
		_w17227_
	);
	LUT2 #(
		.INIT('h4)
	) name16696 (
		_w17226_,
		_w17227_,
		_w17228_
	);
	LUT2 #(
		.INIT('h8)
	) name16697 (
		\key[26]_pad ,
		ld_pad,
		_w17229_
	);
	LUT2 #(
		.INIT('h1)
	) name16698 (
		_w17228_,
		_w17229_,
		_w17230_
	);
	LUT2 #(
		.INIT('h4)
	) name16699 (
		\u0_w_reg[3][30]/P0001 ,
		_w17204_,
		_w17231_
	);
	LUT2 #(
		.INIT('h2)
	) name16700 (
		\u0_w_reg[3][30]/P0001 ,
		_w17204_,
		_w17232_
	);
	LUT2 #(
		.INIT('h1)
	) name16701 (
		ld_pad,
		_w17231_,
		_w17233_
	);
	LUT2 #(
		.INIT('h4)
	) name16702 (
		_w17232_,
		_w17233_,
		_w17234_
	);
	LUT2 #(
		.INIT('h8)
	) name16703 (
		\key[30]_pad ,
		ld_pad,
		_w17235_
	);
	LUT2 #(
		.INIT('h1)
	) name16704 (
		_w17234_,
		_w17235_,
		_w17236_
	);
	LUT2 #(
		.INIT('h4)
	) name16705 (
		\u0_w_reg[3][31]/P0001 ,
		_w17213_,
		_w17237_
	);
	LUT2 #(
		.INIT('h2)
	) name16706 (
		\u0_w_reg[3][31]/P0001 ,
		_w17213_,
		_w17238_
	);
	LUT2 #(
		.INIT('h1)
	) name16707 (
		ld_pad,
		_w17237_,
		_w17239_
	);
	LUT2 #(
		.INIT('h4)
	) name16708 (
		_w17238_,
		_w17239_,
		_w17240_
	);
	LUT2 #(
		.INIT('h8)
	) name16709 (
		\key[31]_pad ,
		ld_pad,
		_w17241_
	);
	LUT2 #(
		.INIT('h1)
	) name16710 (
		_w17240_,
		_w17241_,
		_w17242_
	);
	LUT2 #(
		.INIT('h4)
	) name16711 (
		ld_pad,
		_w15880_,
		_w17243_
	);
	LUT2 #(
		.INIT('h8)
	) name16712 (
		\key[117]_pad ,
		ld_pad,
		_w17244_
	);
	LUT2 #(
		.INIT('h1)
	) name16713 (
		_w17243_,
		_w17244_,
		_w17245_
	);
	LUT2 #(
		.INIT('h1)
	) name16714 (
		\u0_w_reg[1][21]/P0001 ,
		_w15880_,
		_w17246_
	);
	LUT2 #(
		.INIT('h8)
	) name16715 (
		\u0_w_reg[1][21]/P0001 ,
		_w15880_,
		_w17247_
	);
	LUT2 #(
		.INIT('h1)
	) name16716 (
		ld_pad,
		_w17246_,
		_w17248_
	);
	LUT2 #(
		.INIT('h4)
	) name16717 (
		_w17247_,
		_w17248_,
		_w17249_
	);
	LUT2 #(
		.INIT('h8)
	) name16718 (
		\key[85]_pad ,
		ld_pad,
		_w17250_
	);
	LUT2 #(
		.INIT('h1)
	) name16719 (
		_w17249_,
		_w17250_,
		_w17251_
	);
	LUT2 #(
		.INIT('h4)
	) name16720 (
		\u0_w_reg[3][21]/P0001 ,
		_w15886_,
		_w17252_
	);
	LUT2 #(
		.INIT('h2)
	) name16721 (
		\u0_w_reg[3][21]/P0001 ,
		_w15886_,
		_w17253_
	);
	LUT2 #(
		.INIT('h1)
	) name16722 (
		ld_pad,
		_w17252_,
		_w17254_
	);
	LUT2 #(
		.INIT('h4)
	) name16723 (
		_w17253_,
		_w17254_,
		_w17255_
	);
	LUT2 #(
		.INIT('h8)
	) name16724 (
		\key[21]_pad ,
		ld_pad,
		_w17256_
	);
	LUT2 #(
		.INIT('h1)
	) name16725 (
		_w17255_,
		_w17256_,
		_w17257_
	);
	LUT2 #(
		.INIT('h4)
	) name16726 (
		\key[39]_pad ,
		ld_pad,
		_w17258_
	);
	LUT2 #(
		.INIT('h8)
	) name16727 (
		\u0_w_reg[3][30]/P0001 ,
		_w16105_,
		_w17259_
	);
	LUT2 #(
		.INIT('h8)
	) name16728 (
		_w16386_,
		_w17259_,
		_w17260_
	);
	LUT2 #(
		.INIT('h4)
	) name16729 (
		\u0_w_reg[3][28]/P0001 ,
		_w16122_,
		_w17261_
	);
	LUT2 #(
		.INIT('h8)
	) name16730 (
		_w16019_,
		_w17261_,
		_w17262_
	);
	LUT2 #(
		.INIT('h2)
	) name16731 (
		\u0_w_reg[3][28]/P0001 ,
		_w16079_,
		_w17263_
	);
	LUT2 #(
		.INIT('h1)
	) name16732 (
		\u0_w_reg[3][28]/P0001 ,
		_w16098_,
		_w17264_
	);
	LUT2 #(
		.INIT('h2)
	) name16733 (
		_w16036_,
		_w17263_,
		_w17265_
	);
	LUT2 #(
		.INIT('h4)
	) name16734 (
		_w17264_,
		_w17265_,
		_w17266_
	);
	LUT2 #(
		.INIT('h1)
	) name16735 (
		_w16143_,
		_w16407_,
		_w17267_
	);
	LUT2 #(
		.INIT('h1)
	) name16736 (
		_w17260_,
		_w17262_,
		_w17268_
	);
	LUT2 #(
		.INIT('h8)
	) name16737 (
		_w17267_,
		_w17268_,
		_w17269_
	);
	LUT2 #(
		.INIT('h4)
	) name16738 (
		_w17266_,
		_w17269_,
		_w17270_
	);
	LUT2 #(
		.INIT('h8)
	) name16739 (
		\u0_w_reg[3][28]/P0001 ,
		_w16140_,
		_w17271_
	);
	LUT2 #(
		.INIT('h4)
	) name16740 (
		_w16099_,
		_w17263_,
		_w17272_
	);
	LUT2 #(
		.INIT('h1)
	) name16741 (
		_w16058_,
		_w16140_,
		_w17273_
	);
	LUT2 #(
		.INIT('h4)
	) name16742 (
		_w17272_,
		_w17273_,
		_w17274_
	);
	LUT2 #(
		.INIT('h1)
	) name16743 (
		\u0_w_reg[3][26]/P0001 ,
		_w17274_,
		_w17275_
	);
	LUT2 #(
		.INIT('h8)
	) name16744 (
		_w16032_,
		_w16079_,
		_w17276_
	);
	LUT2 #(
		.INIT('h4)
	) name16745 (
		\u0_w_reg[3][28]/P0001 ,
		_w16171_,
		_w17277_
	);
	LUT2 #(
		.INIT('h8)
	) name16746 (
		_w16036_,
		_w17277_,
		_w17278_
	);
	LUT2 #(
		.INIT('h1)
	) name16747 (
		_w17271_,
		_w17276_,
		_w17279_
	);
	LUT2 #(
		.INIT('h4)
	) name16748 (
		_w17278_,
		_w17279_,
		_w17280_
	);
	LUT2 #(
		.INIT('h4)
	) name16749 (
		_w17275_,
		_w17280_,
		_w17281_
	);
	LUT2 #(
		.INIT('h8)
	) name16750 (
		_w17270_,
		_w17281_,
		_w17282_
	);
	LUT2 #(
		.INIT('h2)
	) name16751 (
		\u0_w_reg[3][24]/P0001 ,
		_w17282_,
		_w17283_
	);
	LUT2 #(
		.INIT('h8)
	) name16752 (
		_w16117_,
		_w17277_,
		_w17284_
	);
	LUT2 #(
		.INIT('h8)
	) name16753 (
		_w16017_,
		_w16087_,
		_w17285_
	);
	LUT2 #(
		.INIT('h1)
	) name16754 (
		_w16129_,
		_w17285_,
		_w17286_
	);
	LUT2 #(
		.INIT('h4)
	) name16755 (
		\u0_w_reg[3][29]/P0001 ,
		_w16066_,
		_w17287_
	);
	LUT2 #(
		.INIT('h1)
	) name16756 (
		\u0_w_reg[3][26]/P0001 ,
		_w16141_,
		_w17288_
	);
	LUT2 #(
		.INIT('h4)
	) name16757 (
		_w17287_,
		_w17288_,
		_w17289_
	);
	LUT2 #(
		.INIT('h8)
	) name16758 (
		_w17286_,
		_w17289_,
		_w17290_
	);
	LUT2 #(
		.INIT('h8)
	) name16759 (
		_w16388_,
		_w16392_,
		_w17291_
	);
	LUT2 #(
		.INIT('h2)
	) name16760 (
		\u0_w_reg[3][26]/P0001 ,
		_w16063_,
		_w17292_
	);
	LUT2 #(
		.INIT('h4)
	) name16761 (
		_w16144_,
		_w17292_,
		_w17293_
	);
	LUT2 #(
		.INIT('h4)
	) name16762 (
		_w17291_,
		_w17293_,
		_w17294_
	);
	LUT2 #(
		.INIT('h1)
	) name16763 (
		_w17290_,
		_w17294_,
		_w17295_
	);
	LUT2 #(
		.INIT('h1)
	) name16764 (
		\u0_w_reg[3][25]/P0001 ,
		_w16385_,
		_w17296_
	);
	LUT2 #(
		.INIT('h4)
	) name16765 (
		_w17284_,
		_w17296_,
		_w17297_
	);
	LUT2 #(
		.INIT('h4)
	) name16766 (
		_w17295_,
		_w17297_,
		_w17298_
	);
	LUT2 #(
		.INIT('h4)
	) name16767 (
		_w17283_,
		_w17298_,
		_w17299_
	);
	LUT2 #(
		.INIT('h1)
	) name16768 (
		_w16014_,
		_w16438_,
		_w17300_
	);
	LUT2 #(
		.INIT('h8)
	) name16769 (
		\u0_w_reg[3][27]/P0001 ,
		_w16025_,
		_w17301_
	);
	LUT2 #(
		.INIT('h1)
	) name16770 (
		_w16125_,
		_w17301_,
		_w17302_
	);
	LUT2 #(
		.INIT('h8)
	) name16771 (
		_w17300_,
		_w17302_,
		_w17303_
	);
	LUT2 #(
		.INIT('h2)
	) name16772 (
		\u0_w_reg[3][26]/P0001 ,
		_w17303_,
		_w17304_
	);
	LUT2 #(
		.INIT('h8)
	) name16773 (
		_w16171_,
		_w16386_,
		_w17305_
	);
	LUT2 #(
		.INIT('h4)
	) name16774 (
		\u0_w_reg[3][30]/P0001 ,
		_w17305_,
		_w17306_
	);
	LUT2 #(
		.INIT('h1)
	) name16775 (
		_w17291_,
		_w17306_,
		_w17307_
	);
	LUT2 #(
		.INIT('h4)
	) name16776 (
		_w17304_,
		_w17307_,
		_w17308_
	);
	LUT2 #(
		.INIT('h8)
	) name16777 (
		_w17270_,
		_w17308_,
		_w17309_
	);
	LUT2 #(
		.INIT('h2)
	) name16778 (
		\u0_w_reg[3][24]/P0001 ,
		_w17309_,
		_w17310_
	);
	LUT2 #(
		.INIT('h2)
	) name16779 (
		\u0_w_reg[3][31]/P0001 ,
		_w17300_,
		_w17311_
	);
	LUT2 #(
		.INIT('h1)
	) name16780 (
		_w16118_,
		_w17311_,
		_w17312_
	);
	LUT2 #(
		.INIT('h1)
	) name16781 (
		\u0_w_reg[3][27]/P0001 ,
		_w17312_,
		_w17313_
	);
	LUT2 #(
		.INIT('h2)
	) name16782 (
		\u0_w_reg[3][26]/P0001 ,
		_w16013_,
		_w17314_
	);
	LUT2 #(
		.INIT('h4)
	) name16783 (
		_w16172_,
		_w17314_,
		_w17315_
	);
	LUT2 #(
		.INIT('h4)
	) name16784 (
		_w17313_,
		_w17315_,
		_w17316_
	);
	LUT2 #(
		.INIT('h1)
	) name16785 (
		_w16040_,
		_w16428_,
		_w17317_
	);
	LUT2 #(
		.INIT('h8)
	) name16786 (
		\u0_w_reg[3][29]/P0001 ,
		_w16051_,
		_w17318_
	);
	LUT2 #(
		.INIT('h2)
	) name16787 (
		_w17317_,
		_w17318_,
		_w17319_
	);
	LUT2 #(
		.INIT('h2)
	) name16788 (
		\u0_w_reg[3][27]/P0001 ,
		_w17319_,
		_w17320_
	);
	LUT2 #(
		.INIT('h4)
	) name16789 (
		_w16080_,
		_w17289_,
		_w17321_
	);
	LUT2 #(
		.INIT('h4)
	) name16790 (
		_w17320_,
		_w17321_,
		_w17322_
	);
	LUT2 #(
		.INIT('h1)
	) name16791 (
		_w17316_,
		_w17322_,
		_w17323_
	);
	LUT2 #(
		.INIT('h2)
	) name16792 (
		\u0_w_reg[3][25]/P0001 ,
		_w17310_,
		_w17324_
	);
	LUT2 #(
		.INIT('h4)
	) name16793 (
		_w17323_,
		_w17324_,
		_w17325_
	);
	LUT2 #(
		.INIT('h1)
	) name16794 (
		_w17299_,
		_w17325_,
		_w17326_
	);
	LUT2 #(
		.INIT('h8)
	) name16795 (
		\u0_w_reg[3][28]/P0001 ,
		_w16100_,
		_w17327_
	);
	LUT2 #(
		.INIT('h8)
	) name16796 (
		_w16012_,
		_w16019_,
		_w17328_
	);
	LUT2 #(
		.INIT('h1)
	) name16797 (
		_w16046_,
		_w17328_,
		_w17329_
	);
	LUT2 #(
		.INIT('h1)
	) name16798 (
		\u0_w_reg[3][26]/P0001 ,
		_w17329_,
		_w17330_
	);
	LUT2 #(
		.INIT('h4)
	) name16799 (
		\u0_w_reg[3][30]/P0001 ,
		_w16146_,
		_w17331_
	);
	LUT2 #(
		.INIT('h8)
	) name16800 (
		_w16036_,
		_w16160_,
		_w17332_
	);
	LUT2 #(
		.INIT('h2)
	) name16801 (
		\u0_w_reg[3][25]/P0001 ,
		_w17331_,
		_w17333_
	);
	LUT2 #(
		.INIT('h4)
	) name16802 (
		_w17332_,
		_w17333_,
		_w17334_
	);
	LUT2 #(
		.INIT('h1)
	) name16803 (
		_w17327_,
		_w17330_,
		_w17335_
	);
	LUT2 #(
		.INIT('h8)
	) name16804 (
		_w17334_,
		_w17335_,
		_w17336_
	);
	LUT2 #(
		.INIT('h4)
	) name16805 (
		\u0_w_reg[3][28]/P0001 ,
		_w16146_,
		_w17337_
	);
	LUT2 #(
		.INIT('h8)
	) name16806 (
		_w16122_,
		_w16388_,
		_w17338_
	);
	LUT2 #(
		.INIT('h8)
	) name16807 (
		\u0_w_reg[3][26]/P0001 ,
		_w16052_,
		_w17339_
	);
	LUT2 #(
		.INIT('h1)
	) name16808 (
		\u0_w_reg[3][25]/P0001 ,
		_w17337_,
		_w17340_
	);
	LUT2 #(
		.INIT('h1)
	) name16809 (
		_w17338_,
		_w17339_,
		_w17341_
	);
	LUT2 #(
		.INIT('h8)
	) name16810 (
		_w17340_,
		_w17341_,
		_w17342_
	);
	LUT2 #(
		.INIT('h1)
	) name16811 (
		_w17336_,
		_w17342_,
		_w17343_
	);
	LUT2 #(
		.INIT('h4)
	) name16812 (
		\u0_w_reg[3][31]/P0001 ,
		_w16123_,
		_w17344_
	);
	LUT2 #(
		.INIT('h8)
	) name16813 (
		_w16094_,
		_w16105_,
		_w17345_
	);
	LUT2 #(
		.INIT('h1)
	) name16814 (
		\u0_w_reg[3][26]/P0001 ,
		_w16111_,
		_w17346_
	);
	LUT2 #(
		.INIT('h4)
	) name16815 (
		\u0_w_reg[3][25]/P0001 ,
		_w16359_,
		_w17347_
	);
	LUT2 #(
		.INIT('h1)
	) name16816 (
		_w17345_,
		_w17347_,
		_w17348_
	);
	LUT2 #(
		.INIT('h8)
	) name16817 (
		_w17286_,
		_w17348_,
		_w17349_
	);
	LUT2 #(
		.INIT('h8)
	) name16818 (
		_w17346_,
		_w17349_,
		_w17350_
	);
	LUT2 #(
		.INIT('h8)
	) name16819 (
		_w16011_,
		_w16158_,
		_w17351_
	);
	LUT2 #(
		.INIT('h2)
	) name16820 (
		\u0_w_reg[3][26]/P0001 ,
		_w16047_,
		_w17352_
	);
	LUT2 #(
		.INIT('h4)
	) name16821 (
		_w17351_,
		_w17352_,
		_w17353_
	);
	LUT2 #(
		.INIT('h1)
	) name16822 (
		_w17350_,
		_w17353_,
		_w17354_
	);
	LUT2 #(
		.INIT('h1)
	) name16823 (
		_w17343_,
		_w17344_,
		_w17355_
	);
	LUT2 #(
		.INIT('h4)
	) name16824 (
		_w17354_,
		_w17355_,
		_w17356_
	);
	LUT2 #(
		.INIT('h1)
	) name16825 (
		\u0_w_reg[3][24]/P0001 ,
		_w17356_,
		_w17357_
	);
	LUT2 #(
		.INIT('h1)
	) name16826 (
		_w17326_,
		_w17357_,
		_w17358_
	);
	LUT2 #(
		.INIT('h2)
	) name16827 (
		\u0_w_reg[0][7]/P0001 ,
		_w17358_,
		_w17359_
	);
	LUT2 #(
		.INIT('h4)
	) name16828 (
		\u0_w_reg[0][7]/P0001 ,
		_w17358_,
		_w17360_
	);
	LUT2 #(
		.INIT('h1)
	) name16829 (
		_w17359_,
		_w17360_,
		_w17361_
	);
	LUT2 #(
		.INIT('h2)
	) name16830 (
		\u0_w_reg[1][7]/P0001 ,
		\u0_w_reg[2][7]/P0001 ,
		_w17362_
	);
	LUT2 #(
		.INIT('h4)
	) name16831 (
		\u0_w_reg[1][7]/P0001 ,
		\u0_w_reg[2][7]/P0001 ,
		_w17363_
	);
	LUT2 #(
		.INIT('h1)
	) name16832 (
		_w17362_,
		_w17363_,
		_w17364_
	);
	LUT2 #(
		.INIT('h8)
	) name16833 (
		_w17361_,
		_w17364_,
		_w17365_
	);
	LUT2 #(
		.INIT('h1)
	) name16834 (
		_w17361_,
		_w17364_,
		_w17366_
	);
	LUT2 #(
		.INIT('h1)
	) name16835 (
		_w17365_,
		_w17366_,
		_w17367_
	);
	LUT2 #(
		.INIT('h4)
	) name16836 (
		ld_pad,
		_w17367_,
		_w17368_
	);
	LUT2 #(
		.INIT('h1)
	) name16837 (
		_w17258_,
		_w17368_,
		_w17369_
	);
	LUT2 #(
		.INIT('h4)
	) name16838 (
		ld_pad,
		_w16001_,
		_w17370_
	);
	LUT2 #(
		.INIT('h8)
	) name16839 (
		\key[115]_pad ,
		ld_pad,
		_w17371_
	);
	LUT2 #(
		.INIT('h1)
	) name16840 (
		_w17370_,
		_w17371_,
		_w17372_
	);
	LUT2 #(
		.INIT('h1)
	) name16841 (
		\u0_w_reg[1][19]/P0001 ,
		_w16001_,
		_w17373_
	);
	LUT2 #(
		.INIT('h8)
	) name16842 (
		\u0_w_reg[1][19]/P0001 ,
		_w16001_,
		_w17374_
	);
	LUT2 #(
		.INIT('h1)
	) name16843 (
		ld_pad,
		_w17373_,
		_w17375_
	);
	LUT2 #(
		.INIT('h4)
	) name16844 (
		_w17374_,
		_w17375_,
		_w17376_
	);
	LUT2 #(
		.INIT('h8)
	) name16845 (
		\key[83]_pad ,
		ld_pad,
		_w17377_
	);
	LUT2 #(
		.INIT('h1)
	) name16846 (
		_w17376_,
		_w17377_,
		_w17378_
	);
	LUT2 #(
		.INIT('h4)
	) name16847 (
		\u0_w_reg[3][19]/P0001 ,
		_w16007_,
		_w17379_
	);
	LUT2 #(
		.INIT('h2)
	) name16848 (
		\u0_w_reg[3][19]/P0001 ,
		_w16007_,
		_w17380_
	);
	LUT2 #(
		.INIT('h1)
	) name16849 (
		ld_pad,
		_w17379_,
		_w17381_
	);
	LUT2 #(
		.INIT('h4)
	) name16850 (
		_w17380_,
		_w17381_,
		_w17382_
	);
	LUT2 #(
		.INIT('h8)
	) name16851 (
		\key[19]_pad ,
		ld_pad,
		_w17383_
	);
	LUT2 #(
		.INIT('h1)
	) name16852 (
		_w17382_,
		_w17383_,
		_w17384_
	);
	LUT2 #(
		.INIT('h4)
	) name16853 (
		ld_pad,
		_w16190_,
		_w17385_
	);
	LUT2 #(
		.INIT('h8)
	) name16854 (
		\key[101]_pad ,
		ld_pad,
		_w17386_
	);
	LUT2 #(
		.INIT('h1)
	) name16855 (
		_w17385_,
		_w17386_,
		_w17387_
	);
	LUT2 #(
		.INIT('h1)
	) name16856 (
		\u0_w_reg[1][5]/P0001 ,
		_w16190_,
		_w17388_
	);
	LUT2 #(
		.INIT('h8)
	) name16857 (
		\u0_w_reg[1][5]/P0001 ,
		_w16190_,
		_w17389_
	);
	LUT2 #(
		.INIT('h1)
	) name16858 (
		ld_pad,
		_w17388_,
		_w17390_
	);
	LUT2 #(
		.INIT('h4)
	) name16859 (
		_w17389_,
		_w17390_,
		_w17391_
	);
	LUT2 #(
		.INIT('h8)
	) name16860 (
		\key[69]_pad ,
		ld_pad,
		_w17392_
	);
	LUT2 #(
		.INIT('h1)
	) name16861 (
		_w17391_,
		_w17392_,
		_w17393_
	);
	LUT2 #(
		.INIT('h4)
	) name16862 (
		\u0_w_reg[3][5]/P0001 ,
		_w16196_,
		_w17394_
	);
	LUT2 #(
		.INIT('h2)
	) name16863 (
		\u0_w_reg[3][5]/P0001 ,
		_w16196_,
		_w17395_
	);
	LUT2 #(
		.INIT('h1)
	) name16864 (
		ld_pad,
		_w17394_,
		_w17396_
	);
	LUT2 #(
		.INIT('h4)
	) name16865 (
		_w17395_,
		_w17396_,
		_w17397_
	);
	LUT2 #(
		.INIT('h8)
	) name16866 (
		\key[5]_pad ,
		ld_pad,
		_w17398_
	);
	LUT2 #(
		.INIT('h1)
	) name16867 (
		_w17397_,
		_w17398_,
		_w17399_
	);
	LUT2 #(
		.INIT('h4)
	) name16868 (
		\key[32]_pad ,
		ld_pad,
		_w17400_
	);
	LUT2 #(
		.INIT('h4)
	) name16869 (
		\u0_w_reg[3][29]/P0001 ,
		_w16032_,
		_w17401_
	);
	LUT2 #(
		.INIT('h4)
	) name16870 (
		\u0_w_reg[3][27]/P0001 ,
		_w16052_,
		_w17402_
	);
	LUT2 #(
		.INIT('h8)
	) name16871 (
		\u0_w_reg[3][29]/P0001 ,
		_w17259_,
		_w17403_
	);
	LUT2 #(
		.INIT('h1)
	) name16872 (
		_w17402_,
		_w17403_,
		_w17404_
	);
	LUT2 #(
		.INIT('h2)
	) name16873 (
		\u0_w_reg[3][26]/P0001 ,
		_w17404_,
		_w17405_
	);
	LUT2 #(
		.INIT('h1)
	) name16874 (
		_w16450_,
		_w17306_,
		_w17406_
	);
	LUT2 #(
		.INIT('h2)
	) name16875 (
		\u0_w_reg[3][28]/P0001 ,
		_w17406_,
		_w17407_
	);
	LUT2 #(
		.INIT('h1)
	) name16876 (
		\u0_w_reg[3][25]/P0001 ,
		_w17285_,
		_w17408_
	);
	LUT2 #(
		.INIT('h1)
	) name16877 (
		_w16044_,
		_w17401_,
		_w17409_
	);
	LUT2 #(
		.INIT('h8)
	) name16878 (
		_w17408_,
		_w17409_,
		_w17410_
	);
	LUT2 #(
		.INIT('h4)
	) name16879 (
		_w17405_,
		_w17410_,
		_w17411_
	);
	LUT2 #(
		.INIT('h4)
	) name16880 (
		_w17407_,
		_w17411_,
		_w17412_
	);
	LUT2 #(
		.INIT('h4)
	) name16881 (
		\u0_w_reg[3][26]/P0001 ,
		_w16011_,
		_w17413_
	);
	LUT2 #(
		.INIT('h1)
	) name16882 (
		_w16161_,
		_w17413_,
		_w17414_
	);
	LUT2 #(
		.INIT('h8)
	) name16883 (
		_w16384_,
		_w17414_,
		_w17415_
	);
	LUT2 #(
		.INIT('h1)
	) name16884 (
		_w17412_,
		_w17415_,
		_w17416_
	);
	LUT2 #(
		.INIT('h4)
	) name16885 (
		\u0_w_reg[3][28]/P0001 ,
		_w16060_,
		_w17417_
	);
	LUT2 #(
		.INIT('h1)
	) name16886 (
		_w16047_,
		_w17337_,
		_w17418_
	);
	LUT2 #(
		.INIT('h2)
	) name16887 (
		\u0_w_reg[3][26]/P0001 ,
		_w16443_,
		_w17419_
	);
	LUT2 #(
		.INIT('h4)
	) name16888 (
		_w16050_,
		_w17419_,
		_w17420_
	);
	LUT2 #(
		.INIT('h8)
	) name16889 (
		_w17418_,
		_w17420_,
		_w17421_
	);
	LUT2 #(
		.INIT('h8)
	) name16890 (
		\u0_w_reg[3][27]/P0001 ,
		_w16019_,
		_w17422_
	);
	LUT2 #(
		.INIT('h1)
	) name16891 (
		\u0_w_reg[3][26]/P0001 ,
		_w17422_,
		_w17423_
	);
	LUT2 #(
		.INIT('h1)
	) name16892 (
		_w16093_,
		_w16407_,
		_w17424_
	);
	LUT2 #(
		.INIT('h4)
	) name16893 (
		_w16038_,
		_w17424_,
		_w17425_
	);
	LUT2 #(
		.INIT('h8)
	) name16894 (
		_w17423_,
		_w17425_,
		_w17426_
	);
	LUT2 #(
		.INIT('h1)
	) name16895 (
		_w17421_,
		_w17426_,
		_w17427_
	);
	LUT2 #(
		.INIT('h4)
	) name16896 (
		\u0_w_reg[3][27]/P0001 ,
		_w16058_,
		_w17428_
	);
	LUT2 #(
		.INIT('h2)
	) name16897 (
		\u0_w_reg[3][24]/P0001 ,
		_w17428_,
		_w17429_
	);
	LUT2 #(
		.INIT('h4)
	) name16898 (
		_w17417_,
		_w17429_,
		_w17430_
	);
	LUT2 #(
		.INIT('h4)
	) name16899 (
		_w17427_,
		_w17430_,
		_w17431_
	);
	LUT2 #(
		.INIT('h4)
	) name16900 (
		_w17416_,
		_w17431_,
		_w17432_
	);
	LUT2 #(
		.INIT('h1)
	) name16901 (
		_w16019_,
		_w17318_,
		_w17433_
	);
	LUT2 #(
		.INIT('h2)
	) name16902 (
		_w17261_,
		_w17433_,
		_w17434_
	);
	LUT2 #(
		.INIT('h8)
	) name16903 (
		\u0_w_reg[3][26]/P0001 ,
		_w16145_,
		_w17435_
	);
	LUT2 #(
		.INIT('h4)
	) name16904 (
		_w16392_,
		_w17435_,
		_w17436_
	);
	LUT2 #(
		.INIT('h1)
	) name16905 (
		\u0_w_reg[3][27]/P0001 ,
		_w17317_,
		_w17437_
	);
	LUT2 #(
		.INIT('h4)
	) name16906 (
		\u0_w_reg[3][26]/P0001 ,
		_w16066_,
		_w17438_
	);
	LUT2 #(
		.INIT('h1)
	) name16907 (
		\u0_w_reg[3][25]/P0001 ,
		_w17436_,
		_w17439_
	);
	LUT2 #(
		.INIT('h4)
	) name16908 (
		_w17438_,
		_w17439_,
		_w17440_
	);
	LUT2 #(
		.INIT('h4)
	) name16909 (
		_w17437_,
		_w17440_,
		_w17441_
	);
	LUT2 #(
		.INIT('h8)
	) name16910 (
		_w16012_,
		_w16142_,
		_w17442_
	);
	LUT2 #(
		.INIT('h8)
	) name16911 (
		_w16020_,
		_w16392_,
		_w17443_
	);
	LUT2 #(
		.INIT('h4)
	) name16912 (
		_w16045_,
		_w16051_,
		_w17444_
	);
	LUT2 #(
		.INIT('h2)
	) name16913 (
		\u0_w_reg[3][25]/P0001 ,
		_w17305_,
		_w17445_
	);
	LUT2 #(
		.INIT('h1)
	) name16914 (
		_w17443_,
		_w17444_,
		_w17446_
	);
	LUT2 #(
		.INIT('h8)
	) name16915 (
		_w17445_,
		_w17446_,
		_w17447_
	);
	LUT2 #(
		.INIT('h4)
	) name16916 (
		_w17442_,
		_w17447_,
		_w17448_
	);
	LUT2 #(
		.INIT('h1)
	) name16917 (
		_w17441_,
		_w17448_,
		_w17449_
	);
	LUT2 #(
		.INIT('h8)
	) name16918 (
		_w16087_,
		_w16094_,
		_w17450_
	);
	LUT2 #(
		.INIT('h2)
	) name16919 (
		_w16363_,
		_w17450_,
		_w17451_
	);
	LUT2 #(
		.INIT('h1)
	) name16920 (
		\u0_w_reg[3][26]/P0001 ,
		_w17451_,
		_w17452_
	);
	LUT2 #(
		.INIT('h1)
	) name16921 (
		\u0_w_reg[3][24]/P0001 ,
		_w17434_,
		_w17453_
	);
	LUT2 #(
		.INIT('h4)
	) name16922 (
		_w17452_,
		_w17453_,
		_w17454_
	);
	LUT2 #(
		.INIT('h4)
	) name16923 (
		_w17449_,
		_w17454_,
		_w17455_
	);
	LUT2 #(
		.INIT('h1)
	) name16924 (
		_w17432_,
		_w17455_,
		_w17456_
	);
	LUT2 #(
		.INIT('h8)
	) name16925 (
		_w16020_,
		_w16117_,
		_w17457_
	);
	LUT2 #(
		.INIT('h8)
	) name16926 (
		_w16018_,
		_w16036_,
		_w17458_
	);
	LUT2 #(
		.INIT('h1)
	) name16927 (
		_w17457_,
		_w17458_,
		_w17459_
	);
	LUT2 #(
		.INIT('h2)
	) name16928 (
		\u0_w_reg[3][30]/P0001 ,
		_w17459_,
		_w17460_
	);
	LUT2 #(
		.INIT('h1)
	) name16929 (
		_w16060_,
		_w16162_,
		_w17461_
	);
	LUT2 #(
		.INIT('h2)
	) name16930 (
		\u0_w_reg[3][26]/P0001 ,
		_w17461_,
		_w17462_
	);
	LUT2 #(
		.INIT('h4)
	) name16931 (
		\u0_w_reg[3][31]/P0001 ,
		_w17450_,
		_w17463_
	);
	LUT2 #(
		.INIT('h8)
	) name16932 (
		\u0_w_reg[3][27]/P0001 ,
		_w16118_,
		_w17464_
	);
	LUT2 #(
		.INIT('h4)
	) name16933 (
		\u0_w_reg[3][26]/P0001 ,
		_w16385_,
		_w17465_
	);
	LUT2 #(
		.INIT('h1)
	) name16934 (
		_w17463_,
		_w17464_,
		_w17466_
	);
	LUT2 #(
		.INIT('h4)
	) name16935 (
		_w17465_,
		_w17466_,
		_w17467_
	);
	LUT2 #(
		.INIT('h4)
	) name16936 (
		_w17462_,
		_w17467_,
		_w17468_
	);
	LUT2 #(
		.INIT('h2)
	) name16937 (
		\u0_w_reg[3][25]/P0001 ,
		_w17468_,
		_w17469_
	);
	LUT2 #(
		.INIT('h8)
	) name16938 (
		\u0_w_reg[3][26]/P0001 ,
		_w16087_,
		_w17470_
	);
	LUT2 #(
		.INIT('h1)
	) name16939 (
		_w16011_,
		_w16059_,
		_w17471_
	);
	LUT2 #(
		.INIT('h2)
	) name16940 (
		_w17470_,
		_w17471_,
		_w17472_
	);
	LUT2 #(
		.INIT('h4)
	) name16941 (
		_w16026_,
		_w16140_,
		_w17473_
	);
	LUT2 #(
		.INIT('h8)
	) name16942 (
		_w16051_,
		_w16112_,
		_w17474_
	);
	LUT2 #(
		.INIT('h1)
	) name16943 (
		_w16028_,
		_w17473_,
		_w17475_
	);
	LUT2 #(
		.INIT('h4)
	) name16944 (
		_w17474_,
		_w17475_,
		_w17476_
	);
	LUT2 #(
		.INIT('h1)
	) name16945 (
		\u0_w_reg[3][26]/P0001 ,
		_w17476_,
		_w17477_
	);
	LUT2 #(
		.INIT('h1)
	) name16946 (
		_w16104_,
		_w17472_,
		_w17478_
	);
	LUT2 #(
		.INIT('h4)
	) name16947 (
		_w17477_,
		_w17478_,
		_w17479_
	);
	LUT2 #(
		.INIT('h1)
	) name16948 (
		\u0_w_reg[3][25]/P0001 ,
		_w17479_,
		_w17480_
	);
	LUT2 #(
		.INIT('h1)
	) name16949 (
		_w17460_,
		_w17469_,
		_w17481_
	);
	LUT2 #(
		.INIT('h4)
	) name16950 (
		_w17480_,
		_w17481_,
		_w17482_
	);
	LUT2 #(
		.INIT('h4)
	) name16951 (
		_w17456_,
		_w17482_,
		_w17483_
	);
	LUT2 #(
		.INIT('h2)
	) name16952 (
		\u0_w_reg[0][0]/P0001 ,
		_w17483_,
		_w17484_
	);
	LUT2 #(
		.INIT('h4)
	) name16953 (
		\u0_w_reg[0][0]/P0001 ,
		_w17483_,
		_w17485_
	);
	LUT2 #(
		.INIT('h1)
	) name16954 (
		_w17484_,
		_w17485_,
		_w17486_
	);
	LUT2 #(
		.INIT('h2)
	) name16955 (
		\u0_w_reg[1][0]/P0001 ,
		\u0_w_reg[2][0]/P0001 ,
		_w17487_
	);
	LUT2 #(
		.INIT('h4)
	) name16956 (
		\u0_w_reg[1][0]/P0001 ,
		\u0_w_reg[2][0]/P0001 ,
		_w17488_
	);
	LUT2 #(
		.INIT('h1)
	) name16957 (
		_w17487_,
		_w17488_,
		_w17489_
	);
	LUT2 #(
		.INIT('h8)
	) name16958 (
		_w17486_,
		_w17489_,
		_w17490_
	);
	LUT2 #(
		.INIT('h1)
	) name16959 (
		_w17486_,
		_w17489_,
		_w17491_
	);
	LUT2 #(
		.INIT('h1)
	) name16960 (
		_w17490_,
		_w17491_,
		_w17492_
	);
	LUT2 #(
		.INIT('h4)
	) name16961 (
		ld_pad,
		_w17492_,
		_w17493_
	);
	LUT2 #(
		.INIT('h1)
	) name16962 (
		_w17400_,
		_w17493_,
		_w17494_
	);
	LUT2 #(
		.INIT('h4)
	) name16963 (
		\key[42]_pad ,
		ld_pad,
		_w17495_
	);
	LUT2 #(
		.INIT('h8)
	) name16964 (
		\u0_w_reg[3][5]/P0001 ,
		_w16745_,
		_w17496_
	);
	LUT2 #(
		.INIT('h2)
	) name16965 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		_w17497_
	);
	LUT2 #(
		.INIT('h4)
	) name16966 (
		_w16488_,
		_w17497_,
		_w17498_
	);
	LUT2 #(
		.INIT('h8)
	) name16967 (
		_w16580_,
		_w17498_,
		_w17499_
	);
	LUT2 #(
		.INIT('h8)
	) name16968 (
		_w16505_,
		_w16551_,
		_w17500_
	);
	LUT2 #(
		.INIT('h8)
	) name16969 (
		\u0_w_reg[3][5]/P0001 ,
		_w16541_,
		_w17501_
	);
	LUT2 #(
		.INIT('h1)
	) name16970 (
		_w17500_,
		_w17501_,
		_w17502_
	);
	LUT2 #(
		.INIT('h4)
	) name16971 (
		_w16573_,
		_w17502_,
		_w17503_
	);
	LUT2 #(
		.INIT('h2)
	) name16972 (
		_w16524_,
		_w17503_,
		_w17504_
	);
	LUT2 #(
		.INIT('h8)
	) name16973 (
		_w16520_,
		_w16551_,
		_w17505_
	);
	LUT2 #(
		.INIT('h4)
	) name16974 (
		\u0_w_reg[3][6]/P0001 ,
		_w17505_,
		_w17506_
	);
	LUT2 #(
		.INIT('h1)
	) name16975 (
		\u0_w_reg[3][5]/P0001 ,
		_w16554_,
		_w17507_
	);
	LUT2 #(
		.INIT('h2)
	) name16976 (
		_w16622_,
		_w17507_,
		_w17508_
	);
	LUT2 #(
		.INIT('h1)
	) name16977 (
		\u0_w_reg[3][1]/P0001 ,
		_w16550_,
		_w17509_
	);
	LUT2 #(
		.INIT('h1)
	) name16978 (
		_w16604_,
		_w16674_,
		_w17510_
	);
	LUT2 #(
		.INIT('h1)
	) name16979 (
		_w16745_,
		_w17505_,
		_w17511_
	);
	LUT2 #(
		.INIT('h8)
	) name16980 (
		_w17510_,
		_w17511_,
		_w17512_
	);
	LUT2 #(
		.INIT('h4)
	) name16981 (
		_w16696_,
		_w17509_,
		_w17513_
	);
	LUT2 #(
		.INIT('h4)
	) name16982 (
		_w17508_,
		_w17513_,
		_w17514_
	);
	LUT2 #(
		.INIT('h8)
	) name16983 (
		_w17512_,
		_w17514_,
		_w17515_
	);
	LUT2 #(
		.INIT('h4)
	) name16984 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w17516_
	);
	LUT2 #(
		.INIT('h8)
	) name16985 (
		_w16495_,
		_w16658_,
		_w17517_
	);
	LUT2 #(
		.INIT('h8)
	) name16986 (
		_w17516_,
		_w17517_,
		_w17518_
	);
	LUT2 #(
		.INIT('h4)
	) name16987 (
		\u0_w_reg[3][4]/P0001 ,
		_w16548_,
		_w17519_
	);
	LUT2 #(
		.INIT('h8)
	) name16988 (
		\u0_w_reg[3][2]/P0001 ,
		_w17519_,
		_w17520_
	);
	LUT2 #(
		.INIT('h2)
	) name16989 (
		\u0_w_reg[3][1]/P0001 ,
		_w17518_,
		_w17521_
	);
	LUT2 #(
		.INIT('h4)
	) name16990 (
		_w17520_,
		_w17521_,
		_w17522_
	);
	LUT2 #(
		.INIT('h1)
	) name16991 (
		_w17515_,
		_w17522_,
		_w17523_
	);
	LUT2 #(
		.INIT('h2)
	) name16992 (
		\u0_w_reg[3][0]/P0001 ,
		_w16730_,
		_w17524_
	);
	LUT2 #(
		.INIT('h1)
	) name16993 (
		_w17496_,
		_w17499_,
		_w17525_
	);
	LUT2 #(
		.INIT('h4)
	) name16994 (
		_w17506_,
		_w17525_,
		_w17526_
	);
	LUT2 #(
		.INIT('h8)
	) name16995 (
		_w17524_,
		_w17526_,
		_w17527_
	);
	LUT2 #(
		.INIT('h4)
	) name16996 (
		_w17504_,
		_w17527_,
		_w17528_
	);
	LUT2 #(
		.INIT('h4)
	) name16997 (
		_w17523_,
		_w17528_,
		_w17529_
	);
	LUT2 #(
		.INIT('h8)
	) name16998 (
		_w16488_,
		_w16492_,
		_w17530_
	);
	LUT2 #(
		.INIT('h2)
	) name16999 (
		\u0_w_reg[3][1]/P0001 ,
		_w17530_,
		_w17531_
	);
	LUT2 #(
		.INIT('h8)
	) name17000 (
		\u0_w_reg[3][3]/P0001 ,
		_w16541_,
		_w17532_
	);
	LUT2 #(
		.INIT('h8)
	) name17001 (
		\u0_w_reg[3][3]/P0001 ,
		_w16521_,
		_w17533_
	);
	LUT2 #(
		.INIT('h1)
	) name17002 (
		\u0_w_reg[3][2]/P0001 ,
		_w17533_,
		_w17534_
	);
	LUT2 #(
		.INIT('h1)
	) name17003 (
		_w16481_,
		_w17532_,
		_w17535_
	);
	LUT2 #(
		.INIT('h8)
	) name17004 (
		_w17534_,
		_w17535_,
		_w17536_
	);
	LUT2 #(
		.INIT('h2)
	) name17005 (
		\u0_w_reg[3][2]/P0001 ,
		_w16622_,
		_w17537_
	);
	LUT2 #(
		.INIT('h4)
	) name17006 (
		_w16657_,
		_w17537_,
		_w17538_
	);
	LUT2 #(
		.INIT('h1)
	) name17007 (
		_w17536_,
		_w17538_,
		_w17539_
	);
	LUT2 #(
		.INIT('h2)
	) name17008 (
		_w17531_,
		_w17539_,
		_w17540_
	);
	LUT2 #(
		.INIT('h8)
	) name17009 (
		_w16551_,
		_w17516_,
		_w17541_
	);
	LUT2 #(
		.INIT('h1)
	) name17010 (
		\u0_w_reg[3][1]/P0001 ,
		_w16529_,
		_w17542_
	);
	LUT2 #(
		.INIT('h4)
	) name17011 (
		_w17541_,
		_w17542_,
		_w17543_
	);
	LUT2 #(
		.INIT('h1)
	) name17012 (
		_w17540_,
		_w17543_,
		_w17544_
	);
	LUT2 #(
		.INIT('h8)
	) name17013 (
		\u0_w_reg[3][4]/P0001 ,
		_w16616_,
		_w17545_
	);
	LUT2 #(
		.INIT('h8)
	) name17014 (
		_w16586_,
		_w16729_,
		_w17546_
	);
	LUT2 #(
		.INIT('h1)
	) name17015 (
		\u0_w_reg[3][0]/P0001 ,
		_w16563_,
		_w17547_
	);
	LUT2 #(
		.INIT('h4)
	) name17016 (
		_w17546_,
		_w17547_,
		_w17548_
	);
	LUT2 #(
		.INIT('h4)
	) name17017 (
		_w17545_,
		_w17548_,
		_w17549_
	);
	LUT2 #(
		.INIT('h4)
	) name17018 (
		_w17544_,
		_w17549_,
		_w17550_
	);
	LUT2 #(
		.INIT('h1)
	) name17019 (
		_w17529_,
		_w17550_,
		_w17551_
	);
	LUT2 #(
		.INIT('h1)
	) name17020 (
		_w16572_,
		_w16697_,
		_w17552_
	);
	LUT2 #(
		.INIT('h4)
	) name17021 (
		_w16737_,
		_w17552_,
		_w17553_
	);
	LUT2 #(
		.INIT('h1)
	) name17022 (
		\u0_w_reg[3][2]/P0001 ,
		_w17553_,
		_w17554_
	);
	LUT2 #(
		.INIT('h1)
	) name17023 (
		_w16478_,
		_w16493_,
		_w17555_
	);
	LUT2 #(
		.INIT('h2)
	) name17024 (
		_w16524_,
		_w17555_,
		_w17556_
	);
	LUT2 #(
		.INIT('h2)
	) name17025 (
		_w16493_,
		_w16658_,
		_w17557_
	);
	LUT2 #(
		.INIT('h4)
	) name17026 (
		_w16667_,
		_w17557_,
		_w17558_
	);
	LUT2 #(
		.INIT('h8)
	) name17027 (
		_w16588_,
		_w16753_,
		_w17559_
	);
	LUT2 #(
		.INIT('h8)
	) name17028 (
		_w16526_,
		_w16667_,
		_w17560_
	);
	LUT2 #(
		.INIT('h1)
	) name17029 (
		\u0_w_reg[3][1]/P0001 ,
		_w17558_,
		_w17561_
	);
	LUT2 #(
		.INIT('h1)
	) name17030 (
		_w17559_,
		_w17560_,
		_w17562_
	);
	LUT2 #(
		.INIT('h8)
	) name17031 (
		_w17561_,
		_w17562_,
		_w17563_
	);
	LUT2 #(
		.INIT('h4)
	) name17032 (
		_w17556_,
		_w17563_,
		_w17564_
	);
	LUT2 #(
		.INIT('h4)
	) name17033 (
		_w17554_,
		_w17564_,
		_w17565_
	);
	LUT2 #(
		.INIT('h8)
	) name17034 (
		\u0_w_reg[3][4]/P0001 ,
		_w16521_,
		_w17566_
	);
	LUT2 #(
		.INIT('h1)
	) name17035 (
		_w16520_,
		_w17566_,
		_w17567_
	);
	LUT2 #(
		.INIT('h2)
	) name17036 (
		\u0_w_reg[3][7]/P0001 ,
		_w17567_,
		_w17568_
	);
	LUT2 #(
		.INIT('h8)
	) name17037 (
		_w16658_,
		_w17533_,
		_w17569_
	);
	LUT2 #(
		.INIT('h1)
	) name17038 (
		_w17568_,
		_w17569_,
		_w17570_
	);
	LUT2 #(
		.INIT('h2)
	) name17039 (
		\u0_w_reg[3][2]/P0001 ,
		_w17570_,
		_w17571_
	);
	LUT2 #(
		.INIT('h1)
	) name17040 (
		_w16497_,
		_w16627_,
		_w17572_
	);
	LUT2 #(
		.INIT('h8)
	) name17041 (
		_w16570_,
		_w16667_,
		_w17573_
	);
	LUT2 #(
		.INIT('h2)
	) name17042 (
		_w17572_,
		_w17573_,
		_w17574_
	);
	LUT2 #(
		.INIT('h1)
	) name17043 (
		\u0_w_reg[3][2]/P0001 ,
		_w17574_,
		_w17575_
	);
	LUT2 #(
		.INIT('h2)
	) name17044 (
		\u0_w_reg[3][1]/P0001 ,
		_w16543_,
		_w17576_
	);
	LUT2 #(
		.INIT('h4)
	) name17045 (
		_w17571_,
		_w17576_,
		_w17577_
	);
	LUT2 #(
		.INIT('h4)
	) name17046 (
		_w17575_,
		_w17577_,
		_w17578_
	);
	LUT2 #(
		.INIT('h1)
	) name17047 (
		_w17565_,
		_w17578_,
		_w17579_
	);
	LUT2 #(
		.INIT('h1)
	) name17048 (
		_w16574_,
		_w16753_,
		_w17580_
	);
	LUT2 #(
		.INIT('h8)
	) name17049 (
		\u0_w_reg[3][2]/P0001 ,
		_w16520_,
		_w17581_
	);
	LUT2 #(
		.INIT('h4)
	) name17050 (
		_w17580_,
		_w17581_,
		_w17582_
	);
	LUT2 #(
		.INIT('h1)
	) name17051 (
		_w16606_,
		_w17582_,
		_w17583_
	);
	LUT2 #(
		.INIT('h4)
	) name17052 (
		_w17551_,
		_w17583_,
		_w17584_
	);
	LUT2 #(
		.INIT('h4)
	) name17053 (
		_w17579_,
		_w17584_,
		_w17585_
	);
	LUT2 #(
		.INIT('h2)
	) name17054 (
		\u0_w_reg[0][10]/P0001 ,
		_w17585_,
		_w17586_
	);
	LUT2 #(
		.INIT('h4)
	) name17055 (
		\u0_w_reg[0][10]/P0001 ,
		_w17585_,
		_w17587_
	);
	LUT2 #(
		.INIT('h1)
	) name17056 (
		_w17586_,
		_w17587_,
		_w17588_
	);
	LUT2 #(
		.INIT('h2)
	) name17057 (
		\u0_w_reg[1][10]/P0001 ,
		\u0_w_reg[2][10]/P0001 ,
		_w17589_
	);
	LUT2 #(
		.INIT('h4)
	) name17058 (
		\u0_w_reg[1][10]/P0001 ,
		\u0_w_reg[2][10]/P0001 ,
		_w17590_
	);
	LUT2 #(
		.INIT('h1)
	) name17059 (
		_w17589_,
		_w17590_,
		_w17591_
	);
	LUT2 #(
		.INIT('h8)
	) name17060 (
		_w17588_,
		_w17591_,
		_w17592_
	);
	LUT2 #(
		.INIT('h1)
	) name17061 (
		_w17588_,
		_w17591_,
		_w17593_
	);
	LUT2 #(
		.INIT('h1)
	) name17062 (
		_w17592_,
		_w17593_,
		_w17594_
	);
	LUT2 #(
		.INIT('h4)
	) name17063 (
		ld_pad,
		_w17594_,
		_w17595_
	);
	LUT2 #(
		.INIT('h1)
	) name17064 (
		_w17495_,
		_w17595_,
		_w17596_
	);
	LUT2 #(
		.INIT('h4)
	) name17065 (
		\key[48]_pad ,
		ld_pad,
		_w17597_
	);
	LUT2 #(
		.INIT('h8)
	) name17066 (
		\u0_w_reg[3][13]/P0001 ,
		_w15736_,
		_w17598_
	);
	LUT2 #(
		.INIT('h1)
	) name17067 (
		_w15708_,
		_w17598_,
		_w17599_
	);
	LUT2 #(
		.INIT('h2)
	) name17068 (
		_w15800_,
		_w17599_,
		_w17600_
	);
	LUT2 #(
		.INIT('h1)
	) name17069 (
		_w15805_,
		_w15976_,
		_w17601_
	);
	LUT2 #(
		.INIT('h1)
	) name17070 (
		\u0_w_reg[3][11]/P0001 ,
		_w17601_,
		_w17602_
	);
	LUT2 #(
		.INIT('h4)
	) name17071 (
		\u0_w_reg[3][10]/P0001 ,
		_w15737_,
		_w17603_
	);
	LUT2 #(
		.INIT('h8)
	) name17072 (
		\u0_w_reg[3][10]/P0001 ,
		_w15780_,
		_w17604_
	);
	LUT2 #(
		.INIT('h4)
	) name17073 (
		_w15919_,
		_w17604_,
		_w17605_
	);
	LUT2 #(
		.INIT('h1)
	) name17074 (
		\u0_w_reg[3][9]/P0001 ,
		_w17603_,
		_w17606_
	);
	LUT2 #(
		.INIT('h4)
	) name17075 (
		_w17605_,
		_w17606_,
		_w17607_
	);
	LUT2 #(
		.INIT('h4)
	) name17076 (
		_w17602_,
		_w17607_,
		_w17608_
	);
	LUT2 #(
		.INIT('h4)
	) name17077 (
		\u0_w_reg[3][11]/P0001 ,
		_w15736_,
		_w17609_
	);
	LUT2 #(
		.INIT('h8)
	) name17078 (
		_w15814_,
		_w15847_,
		_w17610_
	);
	LUT2 #(
		.INIT('h4)
	) name17079 (
		\u0_w_reg[3][15]/P0001 ,
		_w15791_,
		_w17611_
	);
	LUT2 #(
		.INIT('h1)
	) name17080 (
		_w15704_,
		_w17611_,
		_w17612_
	);
	LUT2 #(
		.INIT('h2)
	) name17081 (
		\u0_w_reg[3][11]/P0001 ,
		_w17612_,
		_w17613_
	);
	LUT2 #(
		.INIT('h2)
	) name17082 (
		\u0_w_reg[3][9]/P0001 ,
		_w15820_,
		_w17614_
	);
	LUT2 #(
		.INIT('h1)
	) name17083 (
		_w17609_,
		_w17610_,
		_w17615_
	);
	LUT2 #(
		.INIT('h8)
	) name17084 (
		_w17614_,
		_w17615_,
		_w17616_
	);
	LUT2 #(
		.INIT('h4)
	) name17085 (
		_w17613_,
		_w17616_,
		_w17617_
	);
	LUT2 #(
		.INIT('h1)
	) name17086 (
		_w17608_,
		_w17617_,
		_w17618_
	);
	LUT2 #(
		.INIT('h8)
	) name17087 (
		_w15709_,
		_w15756_,
		_w17619_
	);
	LUT2 #(
		.INIT('h1)
	) name17088 (
		_w15954_,
		_w17619_,
		_w17620_
	);
	LUT2 #(
		.INIT('h4)
	) name17089 (
		_w15753_,
		_w17620_,
		_w17621_
	);
	LUT2 #(
		.INIT('h1)
	) name17090 (
		\u0_w_reg[3][10]/P0001 ,
		_w17621_,
		_w17622_
	);
	LUT2 #(
		.INIT('h1)
	) name17091 (
		\u0_w_reg[3][8]/P0001 ,
		_w17600_,
		_w17623_
	);
	LUT2 #(
		.INIT('h4)
	) name17092 (
		_w17622_,
		_w17623_,
		_w17624_
	);
	LUT2 #(
		.INIT('h4)
	) name17093 (
		_w17618_,
		_w17624_,
		_w17625_
	);
	LUT2 #(
		.INIT('h1)
	) name17094 (
		_w15704_,
		_w17609_,
		_w17626_
	);
	LUT2 #(
		.INIT('h1)
	) name17095 (
		\u0_w_reg[3][13]/P0001 ,
		_w17626_,
		_w17627_
	);
	LUT2 #(
		.INIT('h1)
	) name17096 (
		_w15851_,
		_w17627_,
		_w17628_
	);
	LUT2 #(
		.INIT('h2)
	) name17097 (
		\u0_w_reg[3][10]/P0001 ,
		_w17628_,
		_w17629_
	);
	LUT2 #(
		.INIT('h8)
	) name17098 (
		_w15709_,
		_w15719_,
		_w17630_
	);
	LUT2 #(
		.INIT('h2)
	) name17099 (
		\u0_w_reg[3][13]/P0001 ,
		_w15742_,
		_w17631_
	);
	LUT2 #(
		.INIT('h2)
	) name17100 (
		_w15724_,
		_w17631_,
		_w17632_
	);
	LUT2 #(
		.INIT('h8)
	) name17101 (
		_w15802_,
		_w15847_,
		_w17633_
	);
	LUT2 #(
		.INIT('h1)
	) name17102 (
		_w17630_,
		_w17632_,
		_w17634_
	);
	LUT2 #(
		.INIT('h4)
	) name17103 (
		_w17633_,
		_w17634_,
		_w17635_
	);
	LUT2 #(
		.INIT('h4)
	) name17104 (
		_w17629_,
		_w17635_,
		_w17636_
	);
	LUT2 #(
		.INIT('h1)
	) name17105 (
		\u0_w_reg[3][9]/P0001 ,
		_w17636_,
		_w17637_
	);
	LUT2 #(
		.INIT('h8)
	) name17106 (
		_w15724_,
		_w15780_,
		_w17638_
	);
	LUT2 #(
		.INIT('h1)
	) name17107 (
		_w15755_,
		_w17638_,
		_w17639_
	);
	LUT2 #(
		.INIT('h2)
	) name17108 (
		\u0_w_reg[3][10]/P0001 ,
		_w15989_,
		_w17640_
	);
	LUT2 #(
		.INIT('h4)
	) name17109 (
		_w15753_,
		_w17640_,
		_w17641_
	);
	LUT2 #(
		.INIT('h8)
	) name17110 (
		_w17639_,
		_w17641_,
		_w17642_
	);
	LUT2 #(
		.INIT('h8)
	) name17111 (
		_w15719_,
		_w15751_,
		_w17643_
	);
	LUT2 #(
		.INIT('h8)
	) name17112 (
		\u0_w_reg[3][11]/P0001 ,
		_w15708_,
		_w17644_
	);
	LUT2 #(
		.INIT('h1)
	) name17113 (
		\u0_w_reg[3][10]/P0001 ,
		_w17644_,
		_w17645_
	);
	LUT2 #(
		.INIT('h1)
	) name17114 (
		_w15915_,
		_w17643_,
		_w17646_
	);
	LUT2 #(
		.INIT('h4)
	) name17115 (
		_w15705_,
		_w17646_,
		_w17647_
	);
	LUT2 #(
		.INIT('h8)
	) name17116 (
		_w17645_,
		_w17647_,
		_w17648_
	);
	LUT2 #(
		.INIT('h1)
	) name17117 (
		_w17642_,
		_w17648_,
		_w17649_
	);
	LUT2 #(
		.INIT('h1)
	) name17118 (
		\u0_w_reg[3][13]/P0001 ,
		_w15736_,
		_w17650_
	);
	LUT2 #(
		.INIT('h1)
	) name17119 (
		\u0_w_reg[3][10]/P0001 ,
		_w15773_,
		_w17651_
	);
	LUT2 #(
		.INIT('h4)
	) name17120 (
		_w17650_,
		_w17651_,
		_w17652_
	);
	LUT2 #(
		.INIT('h1)
	) name17121 (
		_w15826_,
		_w17652_,
		_w17653_
	);
	LUT2 #(
		.INIT('h2)
	) name17122 (
		\u0_w_reg[3][9]/P0001 ,
		_w17653_,
		_w17654_
	);
	LUT2 #(
		.INIT('h8)
	) name17123 (
		_w15724_,
		_w15814_,
		_w17655_
	);
	LUT2 #(
		.INIT('h4)
	) name17124 (
		\u0_w_reg[3][14]/P0001 ,
		_w17655_,
		_w17656_
	);
	LUT2 #(
		.INIT('h2)
	) name17125 (
		\u0_w_reg[3][8]/P0001 ,
		_w15784_,
		_w17657_
	);
	LUT2 #(
		.INIT('h4)
	) name17126 (
		_w17656_,
		_w17657_,
		_w17658_
	);
	LUT2 #(
		.INIT('h4)
	) name17127 (
		_w17654_,
		_w17658_,
		_w17659_
	);
	LUT2 #(
		.INIT('h4)
	) name17128 (
		_w17649_,
		_w17659_,
		_w17660_
	);
	LUT2 #(
		.INIT('h4)
	) name17129 (
		_w17637_,
		_w17660_,
		_w17661_
	);
	LUT2 #(
		.INIT('h1)
	) name17130 (
		_w17625_,
		_w17661_,
		_w17662_
	);
	LUT2 #(
		.INIT('h8)
	) name17131 (
		_w15720_,
		_w15893_,
		_w17663_
	);
	LUT2 #(
		.INIT('h8)
	) name17132 (
		_w15703_,
		_w15849_,
		_w17664_
	);
	LUT2 #(
		.INIT('h1)
	) name17133 (
		_w17663_,
		_w17664_,
		_w17665_
	);
	LUT2 #(
		.INIT('h2)
	) name17134 (
		\u0_w_reg[3][14]/P0001 ,
		_w17665_,
		_w17666_
	);
	LUT2 #(
		.INIT('h8)
	) name17135 (
		_w15713_,
		_w15822_,
		_w17667_
	);
	LUT2 #(
		.INIT('h8)
	) name17136 (
		_w15849_,
		_w17667_,
		_w17668_
	);
	LUT2 #(
		.INIT('h8)
	) name17137 (
		_w15756_,
		_w15896_,
		_w17669_
	);
	LUT2 #(
		.INIT('h1)
	) name17138 (
		_w15930_,
		_w17669_,
		_w17670_
	);
	LUT2 #(
		.INIT('h2)
	) name17139 (
		\u0_w_reg[3][10]/P0001 ,
		_w17670_,
		_w17671_
	);
	LUT2 #(
		.INIT('h8)
	) name17140 (
		_w15773_,
		_w15822_,
		_w17672_
	);
	LUT2 #(
		.INIT('h1)
	) name17141 (
		_w15838_,
		_w15850_,
		_w17673_
	);
	LUT2 #(
		.INIT('h4)
	) name17142 (
		_w17672_,
		_w17673_,
		_w17674_
	);
	LUT2 #(
		.INIT('h2)
	) name17143 (
		_w15847_,
		_w17674_,
		_w17675_
	);
	LUT2 #(
		.INIT('h1)
	) name17144 (
		\u0_w_reg[3][9]/P0001 ,
		_w15861_,
		_w17676_
	);
	LUT2 #(
		.INIT('h4)
	) name17145 (
		_w17668_,
		_w17676_,
		_w17677_
	);
	LUT2 #(
		.INIT('h4)
	) name17146 (
		_w17671_,
		_w17677_,
		_w17678_
	);
	LUT2 #(
		.INIT('h4)
	) name17147 (
		_w17675_,
		_w17678_,
		_w17679_
	);
	LUT2 #(
		.INIT('h4)
	) name17148 (
		\u0_w_reg[3][10]/P0001 ,
		_w15941_,
		_w17680_
	);
	LUT2 #(
		.INIT('h8)
	) name17149 (
		_w15743_,
		_w15803_,
		_w17681_
	);
	LUT2 #(
		.INIT('h8)
	) name17150 (
		_w15724_,
		_w15773_,
		_w17682_
	);
	LUT2 #(
		.INIT('h8)
	) name17151 (
		\u0_w_reg[3][12]/P0001 ,
		_w15708_,
		_w17683_
	);
	LUT2 #(
		.INIT('h8)
	) name17152 (
		_w15893_,
		_w17683_,
		_w17684_
	);
	LUT2 #(
		.INIT('h1)
	) name17153 (
		_w17619_,
		_w17682_,
		_w17685_
	);
	LUT2 #(
		.INIT('h4)
	) name17154 (
		_w17684_,
		_w17685_,
		_w17686_
	);
	LUT2 #(
		.INIT('h1)
	) name17155 (
		\u0_w_reg[3][15]/P0001 ,
		_w17686_,
		_w17687_
	);
	LUT2 #(
		.INIT('h2)
	) name17156 (
		\u0_w_reg[3][9]/P0001 ,
		_w17680_,
		_w17688_
	);
	LUT2 #(
		.INIT('h4)
	) name17157 (
		_w17681_,
		_w17688_,
		_w17689_
	);
	LUT2 #(
		.INIT('h4)
	) name17158 (
		_w17687_,
		_w17689_,
		_w17690_
	);
	LUT2 #(
		.INIT('h1)
	) name17159 (
		_w17679_,
		_w17690_,
		_w17691_
	);
	LUT2 #(
		.INIT('h1)
	) name17160 (
		_w17666_,
		_w17691_,
		_w17692_
	);
	LUT2 #(
		.INIT('h4)
	) name17161 (
		_w17662_,
		_w17692_,
		_w17693_
	);
	LUT2 #(
		.INIT('h2)
	) name17162 (
		\u0_w_reg[0][16]/P0001 ,
		_w17693_,
		_w17694_
	);
	LUT2 #(
		.INIT('h4)
	) name17163 (
		\u0_w_reg[0][16]/P0001 ,
		_w17693_,
		_w17695_
	);
	LUT2 #(
		.INIT('h1)
	) name17164 (
		_w17694_,
		_w17695_,
		_w17696_
	);
	LUT2 #(
		.INIT('h2)
	) name17165 (
		\u0_w_reg[1][16]/P0001 ,
		\u0_w_reg[2][16]/P0001 ,
		_w17697_
	);
	LUT2 #(
		.INIT('h4)
	) name17166 (
		\u0_w_reg[1][16]/P0001 ,
		\u0_w_reg[2][16]/P0001 ,
		_w17698_
	);
	LUT2 #(
		.INIT('h1)
	) name17167 (
		_w17697_,
		_w17698_,
		_w17699_
	);
	LUT2 #(
		.INIT('h8)
	) name17168 (
		_w17696_,
		_w17699_,
		_w17700_
	);
	LUT2 #(
		.INIT('h1)
	) name17169 (
		_w17696_,
		_w17699_,
		_w17701_
	);
	LUT2 #(
		.INIT('h1)
	) name17170 (
		_w17700_,
		_w17701_,
		_w17702_
	);
	LUT2 #(
		.INIT('h4)
	) name17171 (
		ld_pad,
		_w17702_,
		_w17703_
	);
	LUT2 #(
		.INIT('h1)
	) name17172 (
		_w17597_,
		_w17703_,
		_w17704_
	);
	LUT2 #(
		.INIT('h4)
	) name17173 (
		\key[50]_pad ,
		ld_pad,
		_w17705_
	);
	LUT2 #(
		.INIT('h1)
	) name17174 (
		_w15814_,
		_w17598_,
		_w17706_
	);
	LUT2 #(
		.INIT('h2)
	) name17175 (
		_w15709_,
		_w17706_,
		_w17707_
	);
	LUT2 #(
		.INIT('h1)
	) name17176 (
		_w15703_,
		_w15915_,
		_w17708_
	);
	LUT2 #(
		.INIT('h2)
	) name17177 (
		_w15708_,
		_w17708_,
		_w17709_
	);
	LUT2 #(
		.INIT('h1)
	) name17178 (
		_w15896_,
		_w17707_,
		_w17710_
	);
	LUT2 #(
		.INIT('h4)
	) name17179 (
		_w17709_,
		_w17710_,
		_w17711_
	);
	LUT2 #(
		.INIT('h2)
	) name17180 (
		\u0_w_reg[3][10]/P0001 ,
		_w17711_,
		_w17712_
	);
	LUT2 #(
		.INIT('h2)
	) name17181 (
		\u0_w_reg[3][9]/P0001 ,
		_w17712_,
		_w17713_
	);
	LUT2 #(
		.INIT('h1)
	) name17182 (
		_w15756_,
		_w15805_,
		_w17714_
	);
	LUT2 #(
		.INIT('h2)
	) name17183 (
		\u0_w_reg[3][11]/P0001 ,
		_w17714_,
		_w17715_
	);
	LUT2 #(
		.INIT('h4)
	) name17184 (
		_w15941_,
		_w15974_,
		_w17716_
	);
	LUT2 #(
		.INIT('h4)
	) name17185 (
		_w17707_,
		_w17716_,
		_w17717_
	);
	LUT2 #(
		.INIT('h4)
	) name17186 (
		_w17715_,
		_w17717_,
		_w17718_
	);
	LUT2 #(
		.INIT('h8)
	) name17187 (
		\u0_w_reg[3][13]/P0001 ,
		_w17609_,
		_w17719_
	);
	LUT2 #(
		.INIT('h1)
	) name17188 (
		\u0_w_reg[3][10]/P0001 ,
		_w17719_,
		_w17720_
	);
	LUT2 #(
		.INIT('h8)
	) name17189 (
		_w15713_,
		_w15735_,
		_w17721_
	);
	LUT2 #(
		.INIT('h4)
	) name17190 (
		\u0_w_reg[3][15]/P0001 ,
		_w17721_,
		_w17722_
	);
	LUT2 #(
		.INIT('h1)
	) name17191 (
		_w15960_,
		_w17672_,
		_w17723_
	);
	LUT2 #(
		.INIT('h4)
	) name17192 (
		_w17722_,
		_w17723_,
		_w17724_
	);
	LUT2 #(
		.INIT('h8)
	) name17193 (
		_w17720_,
		_w17724_,
		_w17725_
	);
	LUT2 #(
		.INIT('h1)
	) name17194 (
		_w17718_,
		_w17725_,
		_w17726_
	);
	LUT2 #(
		.INIT('h4)
	) name17195 (
		_w15751_,
		_w15756_,
		_w17727_
	);
	LUT2 #(
		.INIT('h4)
	) name17196 (
		_w15822_,
		_w17727_,
		_w17728_
	);
	LUT2 #(
		.INIT('h1)
	) name17197 (
		_w17726_,
		_w17728_,
		_w17729_
	);
	LUT2 #(
		.INIT('h1)
	) name17198 (
		_w17713_,
		_w17729_,
		_w17730_
	);
	LUT2 #(
		.INIT('h8)
	) name17199 (
		\u0_w_reg[3][15]/P0001 ,
		_w17721_,
		_w17731_
	);
	LUT2 #(
		.INIT('h1)
	) name17200 (
		_w15815_,
		_w17731_,
		_w17732_
	);
	LUT2 #(
		.INIT('h4)
	) name17201 (
		_w15752_,
		_w17732_,
		_w17733_
	);
	LUT2 #(
		.INIT('h1)
	) name17202 (
		\u0_w_reg[3][10]/P0001 ,
		_w17733_,
		_w17734_
	);
	LUT2 #(
		.INIT('h1)
	) name17203 (
		_w15788_,
		_w17734_,
		_w17735_
	);
	LUT2 #(
		.INIT('h2)
	) name17204 (
		\u0_w_reg[3][9]/P0001 ,
		_w17735_,
		_w17736_
	);
	LUT2 #(
		.INIT('h8)
	) name17205 (
		\u0_w_reg[3][12]/P0001 ,
		_w15773_,
		_w17737_
	);
	LUT2 #(
		.INIT('h4)
	) name17206 (
		\u0_w_reg[3][15]/P0001 ,
		_w17737_,
		_w17738_
	);
	LUT2 #(
		.INIT('h1)
	) name17207 (
		_w15826_,
		_w15840_,
		_w17739_
	);
	LUT2 #(
		.INIT('h4)
	) name17208 (
		_w17738_,
		_w17739_,
		_w17740_
	);
	LUT2 #(
		.INIT('h2)
	) name17209 (
		_w15799_,
		_w17740_,
		_w17741_
	);
	LUT2 #(
		.INIT('h8)
	) name17210 (
		_w15778_,
		_w15860_,
		_w17742_
	);
	LUT2 #(
		.INIT('h8)
	) name17211 (
		_w15725_,
		_w15893_,
		_w17743_
	);
	LUT2 #(
		.INIT('h1)
	) name17212 (
		\u0_w_reg[3][13]/P0001 ,
		_w15782_,
		_w17744_
	);
	LUT2 #(
		.INIT('h2)
	) name17213 (
		_w17609_,
		_w17744_,
		_w17745_
	);
	LUT2 #(
		.INIT('h1)
	) name17214 (
		\u0_w_reg[3][9]/P0001 ,
		_w15970_,
		_w17746_
	);
	LUT2 #(
		.INIT('h1)
	) name17215 (
		_w17630_,
		_w17742_,
		_w17747_
	);
	LUT2 #(
		.INIT('h4)
	) name17216 (
		_w17743_,
		_w17747_,
		_w17748_
	);
	LUT2 #(
		.INIT('h1)
	) name17217 (
		_w15731_,
		_w17611_,
		_w17749_
	);
	LUT2 #(
		.INIT('h4)
	) name17218 (
		_w17745_,
		_w17746_,
		_w17750_
	);
	LUT2 #(
		.INIT('h8)
	) name17219 (
		_w17749_,
		_w17750_,
		_w17751_
	);
	LUT2 #(
		.INIT('h8)
	) name17220 (
		_w17748_,
		_w17751_,
		_w17752_
	);
	LUT2 #(
		.INIT('h8)
	) name17221 (
		_w15822_,
		_w15860_,
		_w17753_
	);
	LUT2 #(
		.INIT('h2)
	) name17222 (
		\u0_w_reg[3][9]/P0001 ,
		_w17753_,
		_w17754_
	);
	LUT2 #(
		.INIT('h4)
	) name17223 (
		_w17668_,
		_w17754_,
		_w17755_
	);
	LUT2 #(
		.INIT('h1)
	) name17224 (
		_w17752_,
		_w17755_,
		_w17756_
	);
	LUT2 #(
		.INIT('h8)
	) name17225 (
		\u0_w_reg[3][10]/P0001 ,
		_w15784_,
		_w17757_
	);
	LUT2 #(
		.INIT('h8)
	) name17226 (
		_w15736_,
		_w15929_,
		_w17758_
	);
	LUT2 #(
		.INIT('h2)
	) name17227 (
		\u0_w_reg[3][12]/P0001 ,
		_w15919_,
		_w17759_
	);
	LUT2 #(
		.INIT('h2)
	) name17228 (
		_w15726_,
		_w15773_,
		_w17760_
	);
	LUT2 #(
		.INIT('h8)
	) name17229 (
		_w17759_,
		_w17760_,
		_w17761_
	);
	LUT2 #(
		.INIT('h2)
	) name17230 (
		\u0_w_reg[3][8]/P0001 ,
		_w17669_,
		_w17762_
	);
	LUT2 #(
		.INIT('h1)
	) name17231 (
		_w17758_,
		_w17761_,
		_w17763_
	);
	LUT2 #(
		.INIT('h8)
	) name17232 (
		_w17762_,
		_w17763_,
		_w17764_
	);
	LUT2 #(
		.INIT('h4)
	) name17233 (
		_w17757_,
		_w17764_,
		_w17765_
	);
	LUT2 #(
		.INIT('h4)
	) name17234 (
		_w17741_,
		_w17765_,
		_w17766_
	);
	LUT2 #(
		.INIT('h4)
	) name17235 (
		_w17756_,
		_w17766_,
		_w17767_
	);
	LUT2 #(
		.INIT('h8)
	) name17236 (
		_w15719_,
		_w15849_,
		_w17768_
	);
	LUT2 #(
		.INIT('h1)
	) name17237 (
		\u0_w_reg[3][9]/P0001 ,
		_w15941_,
		_w17769_
	);
	LUT2 #(
		.INIT('h4)
	) name17238 (
		_w17768_,
		_w17769_,
		_w17770_
	);
	LUT2 #(
		.INIT('h4)
	) name17239 (
		\u0_w_reg[3][14]/P0001 ,
		_w15781_,
		_w17771_
	);
	LUT2 #(
		.INIT('h8)
	) name17240 (
		\u0_w_reg[3][11]/P0001 ,
		_w15786_,
		_w17772_
	);
	LUT2 #(
		.INIT('h1)
	) name17241 (
		_w15823_,
		_w17772_,
		_w17773_
	);
	LUT2 #(
		.INIT('h8)
	) name17242 (
		_w17645_,
		_w17773_,
		_w17774_
	);
	LUT2 #(
		.INIT('h2)
	) name17243 (
		\u0_w_reg[3][10]/P0001 ,
		_w15717_,
		_w17775_
	);
	LUT2 #(
		.INIT('h4)
	) name17244 (
		_w17609_,
		_w17775_,
		_w17776_
	);
	LUT2 #(
		.INIT('h1)
	) name17245 (
		_w17774_,
		_w17776_,
		_w17777_
	);
	LUT2 #(
		.INIT('h2)
	) name17246 (
		\u0_w_reg[3][9]/P0001 ,
		_w17771_,
		_w17778_
	);
	LUT2 #(
		.INIT('h4)
	) name17247 (
		_w17777_,
		_w17778_,
		_w17779_
	);
	LUT2 #(
		.INIT('h1)
	) name17248 (
		_w17770_,
		_w17779_,
		_w17780_
	);
	LUT2 #(
		.INIT('h8)
	) name17249 (
		_w15708_,
		_w15906_,
		_w17781_
	);
	LUT2 #(
		.INIT('h8)
	) name17250 (
		\u0_w_reg[3][10]/P0001 ,
		_w17781_,
		_w17782_
	);
	LUT2 #(
		.INIT('h1)
	) name17251 (
		\u0_w_reg[3][8]/P0001 ,
		_w15817_,
		_w17783_
	);
	LUT2 #(
		.INIT('h4)
	) name17252 (
		_w15864_,
		_w17783_,
		_w17784_
	);
	LUT2 #(
		.INIT('h4)
	) name17253 (
		_w17782_,
		_w17784_,
		_w17785_
	);
	LUT2 #(
		.INIT('h4)
	) name17254 (
		_w17780_,
		_w17785_,
		_w17786_
	);
	LUT2 #(
		.INIT('h1)
	) name17255 (
		_w17767_,
		_w17786_,
		_w17787_
	);
	LUT2 #(
		.INIT('h1)
	) name17256 (
		_w15990_,
		_w17736_,
		_w17788_
	);
	LUT2 #(
		.INIT('h4)
	) name17257 (
		_w17730_,
		_w17788_,
		_w17789_
	);
	LUT2 #(
		.INIT('h4)
	) name17258 (
		_w17787_,
		_w17789_,
		_w17790_
	);
	LUT2 #(
		.INIT('h2)
	) name17259 (
		\u0_w_reg[0][18]/P0001 ,
		_w17790_,
		_w17791_
	);
	LUT2 #(
		.INIT('h4)
	) name17260 (
		\u0_w_reg[0][18]/P0001 ,
		_w17790_,
		_w17792_
	);
	LUT2 #(
		.INIT('h1)
	) name17261 (
		_w17791_,
		_w17792_,
		_w17793_
	);
	LUT2 #(
		.INIT('h2)
	) name17262 (
		\u0_w_reg[1][18]/P0001 ,
		\u0_w_reg[2][18]/P0001 ,
		_w17794_
	);
	LUT2 #(
		.INIT('h4)
	) name17263 (
		\u0_w_reg[1][18]/P0001 ,
		\u0_w_reg[2][18]/P0001 ,
		_w17795_
	);
	LUT2 #(
		.INIT('h1)
	) name17264 (
		_w17794_,
		_w17795_,
		_w17796_
	);
	LUT2 #(
		.INIT('h8)
	) name17265 (
		_w17793_,
		_w17796_,
		_w17797_
	);
	LUT2 #(
		.INIT('h1)
	) name17266 (
		_w17793_,
		_w17796_,
		_w17798_
	);
	LUT2 #(
		.INIT('h1)
	) name17267 (
		_w17797_,
		_w17798_,
		_w17799_
	);
	LUT2 #(
		.INIT('h4)
	) name17268 (
		ld_pad,
		_w17799_,
		_w17800_
	);
	LUT2 #(
		.INIT('h1)
	) name17269 (
		_w17705_,
		_w17800_,
		_w17801_
	);
	LUT2 #(
		.INIT('h2)
	) name17270 (
		\u0_w_reg[3][26]/P0001 ,
		_w17273_,
		_w17802_
	);
	LUT2 #(
		.INIT('h8)
	) name17271 (
		_w16103_,
		_w16359_,
		_w17803_
	);
	LUT2 #(
		.INIT('h8)
	) name17272 (
		_w16359_,
		_w16392_,
		_w17804_
	);
	LUT2 #(
		.INIT('h4)
	) name17273 (
		\u0_w_reg[3][27]/P0001 ,
		_w16079_,
		_w17805_
	);
	LUT2 #(
		.INIT('h4)
	) name17274 (
		\u0_w_reg[3][31]/P0001 ,
		_w17805_,
		_w17806_
	);
	LUT2 #(
		.INIT('h4)
	) name17275 (
		\u0_w_reg[3][26]/P0001 ,
		_w16021_,
		_w17807_
	);
	LUT2 #(
		.INIT('h8)
	) name17276 (
		_w16125_,
		_w16147_,
		_w17808_
	);
	LUT2 #(
		.INIT('h1)
	) name17277 (
		_w17803_,
		_w17804_,
		_w17809_
	);
	LUT2 #(
		.INIT('h8)
	) name17278 (
		_w17408_,
		_w17809_,
		_w17810_
	);
	LUT2 #(
		.INIT('h1)
	) name17279 (
		_w17806_,
		_w17807_,
		_w17811_
	);
	LUT2 #(
		.INIT('h4)
	) name17280 (
		_w17808_,
		_w17811_,
		_w17812_
	);
	LUT2 #(
		.INIT('h4)
	) name17281 (
		_w17802_,
		_w17810_,
		_w17813_
	);
	LUT2 #(
		.INIT('h8)
	) name17282 (
		_w17812_,
		_w17813_,
		_w17814_
	);
	LUT2 #(
		.INIT('h1)
	) name17283 (
		\u0_w_reg[3][26]/P0001 ,
		_w16027_,
		_w17815_
	);
	LUT2 #(
		.INIT('h1)
	) name17284 (
		_w16164_,
		_w16386_,
		_w17816_
	);
	LUT2 #(
		.INIT('h4)
	) name17285 (
		_w17815_,
		_w17816_,
		_w17817_
	);
	LUT2 #(
		.INIT('h2)
	) name17286 (
		\u0_w_reg[3][25]/P0001 ,
		_w17817_,
		_w17818_
	);
	LUT2 #(
		.INIT('h1)
	) name17287 (
		_w17814_,
		_w17818_,
		_w17819_
	);
	LUT2 #(
		.INIT('h8)
	) name17288 (
		\u0_w_reg[3][28]/P0001 ,
		_w17318_,
		_w17820_
	);
	LUT2 #(
		.INIT('h1)
	) name17289 (
		_w16037_,
		_w16161_,
		_w17821_
	);
	LUT2 #(
		.INIT('h4)
	) name17290 (
		_w17820_,
		_w17821_,
		_w17822_
	);
	LUT2 #(
		.INIT('h2)
	) name17291 (
		_w16122_,
		_w17822_,
		_w17823_
	);
	LUT2 #(
		.INIT('h8)
	) name17292 (
		_w16036_,
		_w16058_,
		_w17824_
	);
	LUT2 #(
		.INIT('h4)
	) name17293 (
		\u0_w_reg[3][30]/P0001 ,
		_w16360_,
		_w17825_
	);
	LUT2 #(
		.INIT('h4)
	) name17294 (
		\u0_w_reg[3][29]/P0001 ,
		_w17825_,
		_w17826_
	);
	LUT2 #(
		.INIT('h2)
	) name17295 (
		_w16029_,
		_w16392_,
		_w17827_
	);
	LUT2 #(
		.INIT('h8)
	) name17296 (
		_w17263_,
		_w17827_,
		_w17828_
	);
	LUT2 #(
		.INIT('h2)
	) name17297 (
		\u0_w_reg[3][24]/P0001 ,
		_w17474_,
		_w17829_
	);
	LUT2 #(
		.INIT('h1)
	) name17298 (
		_w17824_,
		_w17828_,
		_w17830_
	);
	LUT2 #(
		.INIT('h8)
	) name17299 (
		_w17829_,
		_w17830_,
		_w17831_
	);
	LUT2 #(
		.INIT('h4)
	) name17300 (
		_w17826_,
		_w17831_,
		_w17832_
	);
	LUT2 #(
		.INIT('h4)
	) name17301 (
		_w17823_,
		_w17832_,
		_w17833_
	);
	LUT2 #(
		.INIT('h4)
	) name17302 (
		_w17819_,
		_w17833_,
		_w17834_
	);
	LUT2 #(
		.INIT('h8)
	) name17303 (
		\u0_w_reg[3][27]/P0001 ,
		_w16098_,
		_w17835_
	);
	LUT2 #(
		.INIT('h1)
	) name17304 (
		_w16406_,
		_w17835_,
		_w17836_
	);
	LUT2 #(
		.INIT('h8)
	) name17305 (
		_w17423_,
		_w17836_,
		_w17837_
	);
	LUT2 #(
		.INIT('h2)
	) name17306 (
		\u0_w_reg[3][26]/P0001 ,
		_w16015_,
		_w17838_
	);
	LUT2 #(
		.INIT('h4)
	) name17307 (
		_w16125_,
		_w17838_,
		_w17839_
	);
	LUT2 #(
		.INIT('h1)
	) name17308 (
		_w17837_,
		_w17839_,
		_w17840_
	);
	LUT2 #(
		.INIT('h1)
	) name17309 (
		_w17331_,
		_w17840_,
		_w17841_
	);
	LUT2 #(
		.INIT('h2)
	) name17310 (
		\u0_w_reg[3][25]/P0001 ,
		_w17841_,
		_w17842_
	);
	LUT2 #(
		.INIT('h8)
	) name17311 (
		_w16045_,
		_w16450_,
		_w17843_
	);
	LUT2 #(
		.INIT('h8)
	) name17312 (
		_w16017_,
		_w16117_,
		_w17844_
	);
	LUT2 #(
		.INIT('h1)
	) name17313 (
		_w16385_,
		_w17844_,
		_w17845_
	);
	LUT2 #(
		.INIT('h1)
	) name17314 (
		\u0_w_reg[3][25]/P0001 ,
		_w17845_,
		_w17846_
	);
	LUT2 #(
		.INIT('h1)
	) name17315 (
		\u0_w_reg[3][24]/P0001 ,
		_w16091_,
		_w17847_
	);
	LUT2 #(
		.INIT('h4)
	) name17316 (
		_w16119_,
		_w17847_,
		_w17848_
	);
	LUT2 #(
		.INIT('h4)
	) name17317 (
		_w17843_,
		_w17848_,
		_w17849_
	);
	LUT2 #(
		.INIT('h4)
	) name17318 (
		_w17846_,
		_w17849_,
		_w17850_
	);
	LUT2 #(
		.INIT('h4)
	) name17319 (
		_w17842_,
		_w17850_,
		_w17851_
	);
	LUT2 #(
		.INIT('h1)
	) name17320 (
		_w17834_,
		_w17851_,
		_w17852_
	);
	LUT2 #(
		.INIT('h1)
	) name17321 (
		_w16172_,
		_w17351_,
		_w17853_
	);
	LUT2 #(
		.INIT('h4)
	) name17322 (
		_w16124_,
		_w17853_,
		_w17854_
	);
	LUT2 #(
		.INIT('h1)
	) name17323 (
		\u0_w_reg[3][26]/P0001 ,
		_w17854_,
		_w17855_
	);
	LUT2 #(
		.INIT('h2)
	) name17324 (
		_w16149_,
		_w17855_,
		_w17856_
	);
	LUT2 #(
		.INIT('h1)
	) name17325 (
		_w16118_,
		_w16367_,
		_w17857_
	);
	LUT2 #(
		.INIT('h8)
	) name17326 (
		_w17346_,
		_w17857_,
		_w17858_
	);
	LUT2 #(
		.INIT('h1)
	) name17327 (
		_w16094_,
		_w16428_,
		_w17859_
	);
	LUT2 #(
		.INIT('h2)
	) name17328 (
		\u0_w_reg[3][27]/P0001 ,
		_w17859_,
		_w17860_
	);
	LUT2 #(
		.INIT('h2)
	) name17329 (
		\u0_w_reg[3][26]/P0001 ,
		_w16385_,
		_w17861_
	);
	LUT2 #(
		.INIT('h4)
	) name17330 (
		_w17860_,
		_w17861_,
		_w17862_
	);
	LUT2 #(
		.INIT('h1)
	) name17331 (
		_w17858_,
		_w17862_,
		_w17863_
	);
	LUT2 #(
		.INIT('h8)
	) name17332 (
		_w16386_,
		_w17318_,
		_w17864_
	);
	LUT2 #(
		.INIT('h1)
	) name17333 (
		\u0_w_reg[3][25]/P0001 ,
		_w17864_,
		_w17865_
	);
	LUT2 #(
		.INIT('h4)
	) name17334 (
		_w16048_,
		_w16094_,
		_w17866_
	);
	LUT2 #(
		.INIT('h4)
	) name17335 (
		_w16039_,
		_w17866_,
		_w17867_
	);
	LUT2 #(
		.INIT('h2)
	) name17336 (
		_w17865_,
		_w17867_,
		_w17868_
	);
	LUT2 #(
		.INIT('h4)
	) name17337 (
		_w17863_,
		_w17868_,
		_w17869_
	);
	LUT2 #(
		.INIT('h1)
	) name17338 (
		_w17856_,
		_w17869_,
		_w17870_
	);
	LUT2 #(
		.INIT('h8)
	) name17339 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		_w17871_
	);
	LUT2 #(
		.INIT('h1)
	) name17340 (
		_w16021_,
		_w16360_,
		_w17872_
	);
	LUT2 #(
		.INIT('h2)
	) name17341 (
		_w17871_,
		_w17872_,
		_w17873_
	);
	LUT2 #(
		.INIT('h8)
	) name17342 (
		\u0_w_reg[3][25]/P0001 ,
		_w16122_,
		_w17874_
	);
	LUT2 #(
		.INIT('h8)
	) name17343 (
		_w16040_,
		_w17874_,
		_w17875_
	);
	LUT2 #(
		.INIT('h1)
	) name17344 (
		_w16171_,
		_w17318_,
		_w17876_
	);
	LUT2 #(
		.INIT('h2)
	) name17345 (
		_w17470_,
		_w17876_,
		_w17877_
	);
	LUT2 #(
		.INIT('h1)
	) name17346 (
		_w16444_,
		_w17875_,
		_w17878_
	);
	LUT2 #(
		.INIT('h4)
	) name17347 (
		_w17873_,
		_w17878_,
		_w17879_
	);
	LUT2 #(
		.INIT('h4)
	) name17348 (
		_w17877_,
		_w17879_,
		_w17880_
	);
	LUT2 #(
		.INIT('h4)
	) name17349 (
		_w17870_,
		_w17880_,
		_w17881_
	);
	LUT2 #(
		.INIT('h4)
	) name17350 (
		_w17852_,
		_w17881_,
		_w17882_
	);
	LUT2 #(
		.INIT('h2)
	) name17351 (
		\u0_w_reg[0][2]/P0001 ,
		_w17882_,
		_w17883_
	);
	LUT2 #(
		.INIT('h4)
	) name17352 (
		\u0_w_reg[0][2]/P0001 ,
		_w17882_,
		_w17884_
	);
	LUT2 #(
		.INIT('h1)
	) name17353 (
		_w17883_,
		_w17884_,
		_w17885_
	);
	LUT2 #(
		.INIT('h8)
	) name17354 (
		\u0_w_reg[1][2]/P0001 ,
		_w17885_,
		_w17886_
	);
	LUT2 #(
		.INIT('h1)
	) name17355 (
		\u0_w_reg[1][2]/P0001 ,
		_w17885_,
		_w17887_
	);
	LUT2 #(
		.INIT('h1)
	) name17356 (
		_w17886_,
		_w17887_,
		_w17888_
	);
	LUT2 #(
		.INIT('h8)
	) name17357 (
		\u0_w_reg[2][2]/P0001 ,
		_w17888_,
		_w17889_
	);
	LUT2 #(
		.INIT('h1)
	) name17358 (
		\u0_w_reg[2][2]/P0001 ,
		_w17888_,
		_w17890_
	);
	LUT2 #(
		.INIT('h1)
	) name17359 (
		_w17889_,
		_w17890_,
		_w17891_
	);
	LUT2 #(
		.INIT('h4)
	) name17360 (
		ld_pad,
		_w17891_,
		_w17892_
	);
	LUT2 #(
		.INIT('h8)
	) name17361 (
		\key[34]_pad ,
		ld_pad,
		_w17893_
	);
	LUT2 #(
		.INIT('h1)
	) name17362 (
		_w17892_,
		_w17893_,
		_w17894_
	);
	LUT2 #(
		.INIT('h4)
	) name17363 (
		\key[46]_pad ,
		ld_pad,
		_w17895_
	);
	LUT2 #(
		.INIT('h8)
	) name17364 (
		_w16493_,
		_w16520_,
		_w17896_
	);
	LUT2 #(
		.INIT('h8)
	) name17365 (
		_w16542_,
		_w16667_,
		_w17897_
	);
	LUT2 #(
		.INIT('h2)
	) name17366 (
		\u0_w_reg[3][2]/P0001 ,
		_w17897_,
		_w17898_
	);
	LUT2 #(
		.INIT('h4)
	) name17367 (
		_w17896_,
		_w17898_,
		_w17899_
	);
	LUT2 #(
		.INIT('h4)
	) name17368 (
		\u0_w_reg[3][3]/P0001 ,
		_w16608_,
		_w17900_
	);
	LUT2 #(
		.INIT('h4)
	) name17369 (
		_w16548_,
		_w16743_,
		_w17901_
	);
	LUT2 #(
		.INIT('h1)
	) name17370 (
		\u0_w_reg[3][2]/P0001 ,
		_w16590_,
		_w17902_
	);
	LUT2 #(
		.INIT('h4)
	) name17371 (
		_w16485_,
		_w17902_,
		_w17903_
	);
	LUT2 #(
		.INIT('h1)
	) name17372 (
		_w17900_,
		_w17901_,
		_w17904_
	);
	LUT2 #(
		.INIT('h8)
	) name17373 (
		_w17903_,
		_w17904_,
		_w17905_
	);
	LUT2 #(
		.INIT('h1)
	) name17374 (
		_w17899_,
		_w17905_,
		_w17906_
	);
	LUT2 #(
		.INIT('h8)
	) name17375 (
		\u0_w_reg[3][7]/P0001 ,
		_w16743_,
		_w17907_
	);
	LUT2 #(
		.INIT('h8)
	) name17376 (
		_w16520_,
		_w16570_,
		_w17908_
	);
	LUT2 #(
		.INIT('h1)
	) name17377 (
		\u0_w_reg[3][1]/P0001 ,
		_w16510_,
		_w17909_
	);
	LUT2 #(
		.INIT('h1)
	) name17378 (
		_w17517_,
		_w17908_,
		_w17910_
	);
	LUT2 #(
		.INIT('h8)
	) name17379 (
		_w17909_,
		_w17910_,
		_w17911_
	);
	LUT2 #(
		.INIT('h1)
	) name17380 (
		_w16754_,
		_w17897_,
		_w17912_
	);
	LUT2 #(
		.INIT('h4)
	) name17381 (
		_w17907_,
		_w17912_,
		_w17913_
	);
	LUT2 #(
		.INIT('h8)
	) name17382 (
		_w17911_,
		_w17913_,
		_w17914_
	);
	LUT2 #(
		.INIT('h8)
	) name17383 (
		\u0_w_reg[3][4]/P0001 ,
		_w16476_,
		_w17915_
	);
	LUT2 #(
		.INIT('h1)
	) name17384 (
		_w16481_,
		_w17915_,
		_w17916_
	);
	LUT2 #(
		.INIT('h1)
	) name17385 (
		\u0_w_reg[3][2]/P0001 ,
		_w16659_,
		_w17917_
	);
	LUT2 #(
		.INIT('h1)
	) name17386 (
		_w16524_,
		_w17916_,
		_w17918_
	);
	LUT2 #(
		.INIT('h4)
	) name17387 (
		_w17917_,
		_w17918_,
		_w17919_
	);
	LUT2 #(
		.INIT('h2)
	) name17388 (
		\u0_w_reg[3][1]/P0001 ,
		_w16737_,
		_w17920_
	);
	LUT2 #(
		.INIT('h4)
	) name17389 (
		_w17919_,
		_w17920_,
		_w17921_
	);
	LUT2 #(
		.INIT('h1)
	) name17390 (
		_w17914_,
		_w17921_,
		_w17922_
	);
	LUT2 #(
		.INIT('h1)
	) name17391 (
		_w17906_,
		_w17922_,
		_w17923_
	);
	LUT2 #(
		.INIT('h1)
	) name17392 (
		\u0_w_reg[3][0]/P0001 ,
		_w17923_,
		_w17924_
	);
	LUT2 #(
		.INIT('h1)
	) name17393 (
		_w16622_,
		_w17530_,
		_w17925_
	);
	LUT2 #(
		.INIT('h1)
	) name17394 (
		\u0_w_reg[3][4]/P0001 ,
		_w17925_,
		_w17926_
	);
	LUT2 #(
		.INIT('h4)
	) name17395 (
		\u0_w_reg[3][7]/P0001 ,
		_w16608_,
		_w17927_
	);
	LUT2 #(
		.INIT('h1)
	) name17396 (
		_w17926_,
		_w17927_,
		_w17928_
	);
	LUT2 #(
		.INIT('h2)
	) name17397 (
		\u0_w_reg[3][2]/P0001 ,
		_w17928_,
		_w17929_
	);
	LUT2 #(
		.INIT('h1)
	) name17398 (
		_w17546_,
		_w17929_,
		_w17930_
	);
	LUT2 #(
		.INIT('h2)
	) name17399 (
		\u0_w_reg[3][1]/P0001 ,
		_w17930_,
		_w17931_
	);
	LUT2 #(
		.INIT('h8)
	) name17400 (
		_w16548_,
		_w16664_,
		_w17932_
	);
	LUT2 #(
		.INIT('h1)
	) name17401 (
		_w16573_,
		_w17530_,
		_w17933_
	);
	LUT2 #(
		.INIT('h1)
	) name17402 (
		\u0_w_reg[3][2]/P0001 ,
		_w17933_,
		_w17934_
	);
	LUT2 #(
		.INIT('h4)
	) name17403 (
		\u0_w_reg[3][2]/P0001 ,
		_w16563_,
		_w17935_
	);
	LUT2 #(
		.INIT('h1)
	) name17404 (
		_w16556_,
		_w16572_,
		_w17936_
	);
	LUT2 #(
		.INIT('h4)
	) name17405 (
		_w16527_,
		_w17936_,
		_w17937_
	);
	LUT2 #(
		.INIT('h1)
	) name17406 (
		_w17932_,
		_w17935_,
		_w17938_
	);
	LUT2 #(
		.INIT('h8)
	) name17407 (
		_w17937_,
		_w17938_,
		_w17939_
	);
	LUT2 #(
		.INIT('h4)
	) name17408 (
		_w17934_,
		_w17939_,
		_w17940_
	);
	LUT2 #(
		.INIT('h1)
	) name17409 (
		\u0_w_reg[3][1]/P0001 ,
		_w17940_,
		_w17941_
	);
	LUT2 #(
		.INIT('h1)
	) name17410 (
		_w16623_,
		_w16631_,
		_w17942_
	);
	LUT2 #(
		.INIT('h1)
	) name17411 (
		_w16509_,
		_w17942_,
		_w17943_
	);
	LUT2 #(
		.INIT('h1)
	) name17412 (
		_w16627_,
		_w16630_,
		_w17944_
	);
	LUT2 #(
		.INIT('h1)
	) name17413 (
		\u0_w_reg[3][2]/P0001 ,
		_w17944_,
		_w17945_
	);
	LUT2 #(
		.INIT('h1)
	) name17414 (
		_w16496_,
		_w16522_,
		_w17946_
	);
	LUT2 #(
		.INIT('h2)
	) name17415 (
		\u0_w_reg[3][2]/P0001 ,
		_w17946_,
		_w17947_
	);
	LUT2 #(
		.INIT('h1)
	) name17416 (
		_w16563_,
		_w17559_,
		_w17948_
	);
	LUT2 #(
		.INIT('h4)
	) name17417 (
		_w17947_,
		_w17948_,
		_w17949_
	);
	LUT2 #(
		.INIT('h4)
	) name17418 (
		_w17945_,
		_w17949_,
		_w17950_
	);
	LUT2 #(
		.INIT('h1)
	) name17419 (
		\u0_w_reg[3][1]/P0001 ,
		_w17950_,
		_w17951_
	);
	LUT2 #(
		.INIT('h8)
	) name17420 (
		\u0_w_reg[3][4]/P0001 ,
		_w16488_,
		_w17952_
	);
	LUT2 #(
		.INIT('h8)
	) name17421 (
		_w16588_,
		_w17952_,
		_w17953_
	);
	LUT2 #(
		.INIT('h1)
	) name17422 (
		_w16494_,
		_w16659_,
		_w17954_
	);
	LUT2 #(
		.INIT('h8)
	) name17423 (
		_w16534_,
		_w17954_,
		_w17955_
	);
	LUT2 #(
		.INIT('h2)
	) name17424 (
		\u0_w_reg[3][2]/P0001 ,
		_w17955_,
		_w17956_
	);
	LUT2 #(
		.INIT('h8)
	) name17425 (
		_w16588_,
		_w16653_,
		_w17957_
	);
	LUT2 #(
		.INIT('h8)
	) name17426 (
		_w16476_,
		_w16612_,
		_w17958_
	);
	LUT2 #(
		.INIT('h8)
	) name17427 (
		_w16488_,
		_w16532_,
		_w17959_
	);
	LUT2 #(
		.INIT('h4)
	) name17428 (
		\u0_w_reg[3][3]/P0001 ,
		_w16627_,
		_w17960_
	);
	LUT2 #(
		.INIT('h8)
	) name17429 (
		\u0_w_reg[3][4]/P0001 ,
		_w16483_,
		_w17961_
	);
	LUT2 #(
		.INIT('h1)
	) name17430 (
		_w16490_,
		_w17961_,
		_w17962_
	);
	LUT2 #(
		.INIT('h4)
	) name17431 (
		_w17960_,
		_w17962_,
		_w17963_
	);
	LUT2 #(
		.INIT('h2)
	) name17432 (
		\u0_w_reg[3][2]/P0001 ,
		_w17963_,
		_w17964_
	);
	LUT2 #(
		.INIT('h1)
	) name17433 (
		_w17957_,
		_w17958_,
		_w17965_
	);
	LUT2 #(
		.INIT('h4)
	) name17434 (
		_w17959_,
		_w17965_,
		_w17966_
	);
	LUT2 #(
		.INIT('h4)
	) name17435 (
		_w17964_,
		_w17966_,
		_w17967_
	);
	LUT2 #(
		.INIT('h2)
	) name17436 (
		\u0_w_reg[3][1]/P0001 ,
		_w17967_,
		_w17968_
	);
	LUT2 #(
		.INIT('h4)
	) name17437 (
		\u0_w_reg[3][2]/P0001 ,
		_w16495_,
		_w17969_
	);
	LUT2 #(
		.INIT('h8)
	) name17438 (
		_w16658_,
		_w17969_,
		_w17970_
	);
	LUT2 #(
		.INIT('h1)
	) name17439 (
		_w17953_,
		_w17970_,
		_w17971_
	);
	LUT2 #(
		.INIT('h4)
	) name17440 (
		_w17956_,
		_w17971_,
		_w17972_
	);
	LUT2 #(
		.INIT('h4)
	) name17441 (
		_w17951_,
		_w17972_,
		_w17973_
	);
	LUT2 #(
		.INIT('h4)
	) name17442 (
		_w17968_,
		_w17973_,
		_w17974_
	);
	LUT2 #(
		.INIT('h2)
	) name17443 (
		\u0_w_reg[3][0]/P0001 ,
		_w17974_,
		_w17975_
	);
	LUT2 #(
		.INIT('h1)
	) name17444 (
		_w16511_,
		_w17943_,
		_w17976_
	);
	LUT2 #(
		.INIT('h4)
	) name17445 (
		_w17941_,
		_w17976_,
		_w17977_
	);
	LUT2 #(
		.INIT('h4)
	) name17446 (
		_w17931_,
		_w17977_,
		_w17978_
	);
	LUT2 #(
		.INIT('h4)
	) name17447 (
		_w17924_,
		_w17978_,
		_w17979_
	);
	LUT2 #(
		.INIT('h4)
	) name17448 (
		_w17975_,
		_w17979_,
		_w17980_
	);
	LUT2 #(
		.INIT('h2)
	) name17449 (
		\u0_w_reg[0][14]/P0001 ,
		_w17980_,
		_w17981_
	);
	LUT2 #(
		.INIT('h4)
	) name17450 (
		\u0_w_reg[0][14]/P0001 ,
		_w17980_,
		_w17982_
	);
	LUT2 #(
		.INIT('h1)
	) name17451 (
		_w17981_,
		_w17982_,
		_w17983_
	);
	LUT2 #(
		.INIT('h2)
	) name17452 (
		\u0_w_reg[1][14]/P0001 ,
		\u0_w_reg[2][14]/P0001 ,
		_w17984_
	);
	LUT2 #(
		.INIT('h4)
	) name17453 (
		\u0_w_reg[1][14]/P0001 ,
		\u0_w_reg[2][14]/P0001 ,
		_w17985_
	);
	LUT2 #(
		.INIT('h1)
	) name17454 (
		_w17984_,
		_w17985_,
		_w17986_
	);
	LUT2 #(
		.INIT('h8)
	) name17455 (
		_w17983_,
		_w17986_,
		_w17987_
	);
	LUT2 #(
		.INIT('h1)
	) name17456 (
		_w17983_,
		_w17986_,
		_w17988_
	);
	LUT2 #(
		.INIT('h1)
	) name17457 (
		_w17987_,
		_w17988_,
		_w17989_
	);
	LUT2 #(
		.INIT('h4)
	) name17458 (
		ld_pad,
		_w17989_,
		_w17990_
	);
	LUT2 #(
		.INIT('h1)
	) name17459 (
		_w17895_,
		_w17990_,
		_w17991_
	);
	LUT2 #(
		.INIT('h4)
	) name17460 (
		\key[54]_pad ,
		ld_pad,
		_w17992_
	);
	LUT2 #(
		.INIT('h2)
	) name17461 (
		\u0_w_reg[3][10]/P0001 ,
		_w15838_,
		_w17993_
	);
	LUT2 #(
		.INIT('h4)
	) name17462 (
		_w15906_,
		_w17993_,
		_w17994_
	);
	LUT2 #(
		.INIT('h1)
	) name17463 (
		_w17720_,
		_w17994_,
		_w17995_
	);
	LUT2 #(
		.INIT('h1)
	) name17464 (
		\u0_w_reg[3][10]/P0001 ,
		_w15816_,
		_w17996_
	);
	LUT2 #(
		.INIT('h1)
	) name17465 (
		\u0_w_reg[3][9]/P0001 ,
		_w15817_,
		_w17997_
	);
	LUT2 #(
		.INIT('h4)
	) name17466 (
		_w17995_,
		_w17997_,
		_w17998_
	);
	LUT2 #(
		.INIT('h4)
	) name17467 (
		_w17996_,
		_w17998_,
		_w17999_
	);
	LUT2 #(
		.INIT('h8)
	) name17468 (
		\u0_w_reg[3][15]/P0001 ,
		_w15710_,
		_w18000_
	);
	LUT2 #(
		.INIT('h1)
	) name17469 (
		_w15779_,
		_w15850_,
		_w18001_
	);
	LUT2 #(
		.INIT('h4)
	) name17470 (
		_w18000_,
		_w18001_,
		_w18002_
	);
	LUT2 #(
		.INIT('h2)
	) name17471 (
		\u0_w_reg[3][10]/P0001 ,
		_w18002_,
		_w18003_
	);
	LUT2 #(
		.INIT('h8)
	) name17472 (
		_w15732_,
		_w15847_,
		_w18004_
	);
	LUT2 #(
		.INIT('h2)
	) name17473 (
		\u0_w_reg[3][9]/P0001 ,
		_w18004_,
		_w18005_
	);
	LUT2 #(
		.INIT('h8)
	) name17474 (
		_w17639_,
		_w18005_,
		_w18006_
	);
	LUT2 #(
		.INIT('h4)
	) name17475 (
		_w18003_,
		_w18006_,
		_w18007_
	);
	LUT2 #(
		.INIT('h1)
	) name17476 (
		_w17999_,
		_w18007_,
		_w18008_
	);
	LUT2 #(
		.INIT('h1)
	) name17477 (
		_w15832_,
		_w15920_,
		_w18009_
	);
	LUT2 #(
		.INIT('h4)
	) name17478 (
		_w15744_,
		_w18009_,
		_w18010_
	);
	LUT2 #(
		.INIT('h8)
	) name17479 (
		_w15707_,
		_w18010_,
		_w18011_
	);
	LUT2 #(
		.INIT('h1)
	) name17480 (
		\u0_w_reg[3][10]/P0001 ,
		_w15774_,
		_w18012_
	);
	LUT2 #(
		.INIT('h4)
	) name17481 (
		_w17667_,
		_w18012_,
		_w18013_
	);
	LUT2 #(
		.INIT('h1)
	) name17482 (
		_w18011_,
		_w18013_,
		_w18014_
	);
	LUT2 #(
		.INIT('h1)
	) name17483 (
		_w18008_,
		_w18014_,
		_w18015_
	);
	LUT2 #(
		.INIT('h2)
	) name17484 (
		\u0_w_reg[3][8]/P0001 ,
		_w18015_,
		_w18016_
	);
	LUT2 #(
		.INIT('h8)
	) name17485 (
		_w15751_,
		_w15787_,
		_w18017_
	);
	LUT2 #(
		.INIT('h1)
	) name17486 (
		_w17619_,
		_w18017_,
		_w18018_
	);
	LUT2 #(
		.INIT('h2)
	) name17487 (
		\u0_w_reg[3][10]/P0001 ,
		_w18018_,
		_w18019_
	);
	LUT2 #(
		.INIT('h1)
	) name17488 (
		_w15741_,
		_w15756_,
		_w18020_
	);
	LUT2 #(
		.INIT('h2)
	) name17489 (
		_w15751_,
		_w18020_,
		_w18021_
	);
	LUT2 #(
		.INIT('h8)
	) name17490 (
		_w15724_,
		_w17650_,
		_w18022_
	);
	LUT2 #(
		.INIT('h1)
	) name17491 (
		_w15939_,
		_w18022_,
		_w18023_
	);
	LUT2 #(
		.INIT('h4)
	) name17492 (
		_w18021_,
		_w18023_,
		_w18024_
	);
	LUT2 #(
		.INIT('h1)
	) name17493 (
		\u0_w_reg[3][10]/P0001 ,
		_w18024_,
		_w18025_
	);
	LUT2 #(
		.INIT('h8)
	) name17494 (
		_w15799_,
		_w17598_,
		_w18026_
	);
	LUT2 #(
		.INIT('h8)
	) name17495 (
		_w15709_,
		_w15742_,
		_w18027_
	);
	LUT2 #(
		.INIT('h1)
	) name17496 (
		\u0_w_reg[3][9]/P0001 ,
		_w17655_,
		_w18028_
	);
	LUT2 #(
		.INIT('h1)
	) name17497 (
		_w17664_,
		_w17667_,
		_w18029_
	);
	LUT2 #(
		.INIT('h4)
	) name17498 (
		_w18027_,
		_w18029_,
		_w18030_
	);
	LUT2 #(
		.INIT('h4)
	) name17499 (
		_w18017_,
		_w18028_,
		_w18031_
	);
	LUT2 #(
		.INIT('h4)
	) name17500 (
		_w18026_,
		_w18031_,
		_w18032_
	);
	LUT2 #(
		.INIT('h8)
	) name17501 (
		_w18030_,
		_w18032_,
		_w18033_
	);
	LUT2 #(
		.INIT('h4)
	) name17502 (
		_w15824_,
		_w15893_,
		_w18034_
	);
	LUT2 #(
		.INIT('h4)
	) name17503 (
		\u0_w_reg[3][10]/P0001 ,
		_w15832_,
		_w18035_
	);
	LUT2 #(
		.INIT('h2)
	) name17504 (
		\u0_w_reg[3][9]/P0001 ,
		_w17722_,
		_w18036_
	);
	LUT2 #(
		.INIT('h4)
	) name17505 (
		_w18035_,
		_w18036_,
		_w18037_
	);
	LUT2 #(
		.INIT('h4)
	) name17506 (
		_w18034_,
		_w18037_,
		_w18038_
	);
	LUT2 #(
		.INIT('h1)
	) name17507 (
		_w18033_,
		_w18038_,
		_w18039_
	);
	LUT2 #(
		.INIT('h1)
	) name17508 (
		_w18019_,
		_w18025_,
		_w18040_
	);
	LUT2 #(
		.INIT('h4)
	) name17509 (
		_w18039_,
		_w18040_,
		_w18041_
	);
	LUT2 #(
		.INIT('h1)
	) name17510 (
		\u0_w_reg[3][8]/P0001 ,
		_w18041_,
		_w18042_
	);
	LUT2 #(
		.INIT('h2)
	) name17511 (
		\u0_w_reg[3][10]/P0001 ,
		_w15805_,
		_w18043_
	);
	LUT2 #(
		.INIT('h4)
	) name17512 (
		_w15865_,
		_w18043_,
		_w18044_
	);
	LUT2 #(
		.INIT('h2)
	) name17513 (
		_w15818_,
		_w15826_,
		_w18045_
	);
	LUT2 #(
		.INIT('h4)
	) name17514 (
		_w17771_,
		_w18045_,
		_w18046_
	);
	LUT2 #(
		.INIT('h1)
	) name17515 (
		_w18044_,
		_w18046_,
		_w18047_
	);
	LUT2 #(
		.INIT('h1)
	) name17516 (
		_w15930_,
		_w15960_,
		_w18048_
	);
	LUT2 #(
		.INIT('h4)
	) name17517 (
		_w18047_,
		_w18048_,
		_w18049_
	);
	LUT2 #(
		.INIT('h1)
	) name17518 (
		\u0_w_reg[3][9]/P0001 ,
		_w18049_,
		_w18050_
	);
	LUT2 #(
		.INIT('h4)
	) name17519 (
		\u0_w_reg[3][15]/P0001 ,
		_w17619_,
		_w18051_
	);
	LUT2 #(
		.INIT('h1)
	) name17520 (
		_w15920_,
		_w17609_,
		_w18052_
	);
	LUT2 #(
		.INIT('h2)
	) name17521 (
		_w15803_,
		_w18052_,
		_w18053_
	);
	LUT2 #(
		.INIT('h8)
	) name17522 (
		_w15726_,
		_w15863_,
		_w18054_
	);
	LUT2 #(
		.INIT('h8)
	) name17523 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w18055_
	);
	LUT2 #(
		.INIT('h1)
	) name17524 (
		_w17609_,
		_w17771_,
		_w18056_
	);
	LUT2 #(
		.INIT('h1)
	) name17525 (
		\u0_w_reg[3][12]/P0001 ,
		_w18056_,
		_w18057_
	);
	LUT2 #(
		.INIT('h1)
	) name17526 (
		_w15758_,
		_w18057_,
		_w18058_
	);
	LUT2 #(
		.INIT('h2)
	) name17527 (
		_w18055_,
		_w18058_,
		_w18059_
	);
	LUT2 #(
		.INIT('h1)
	) name17528 (
		_w15892_,
		_w18051_,
		_w18060_
	);
	LUT2 #(
		.INIT('h1)
	) name17529 (
		_w18053_,
		_w18054_,
		_w18061_
	);
	LUT2 #(
		.INIT('h8)
	) name17530 (
		_w18060_,
		_w18061_,
		_w18062_
	);
	LUT2 #(
		.INIT('h4)
	) name17531 (
		_w18059_,
		_w18062_,
		_w18063_
	);
	LUT2 #(
		.INIT('h4)
	) name17532 (
		_w18050_,
		_w18063_,
		_w18064_
	);
	LUT2 #(
		.INIT('h4)
	) name17533 (
		_w18042_,
		_w18064_,
		_w18065_
	);
	LUT2 #(
		.INIT('h4)
	) name17534 (
		_w18016_,
		_w18065_,
		_w18066_
	);
	LUT2 #(
		.INIT('h2)
	) name17535 (
		\u0_w_reg[0][22]/P0001 ,
		_w18066_,
		_w18067_
	);
	LUT2 #(
		.INIT('h4)
	) name17536 (
		\u0_w_reg[0][22]/P0001 ,
		_w18066_,
		_w18068_
	);
	LUT2 #(
		.INIT('h1)
	) name17537 (
		_w18067_,
		_w18068_,
		_w18069_
	);
	LUT2 #(
		.INIT('h2)
	) name17538 (
		\u0_w_reg[1][22]/P0001 ,
		\u0_w_reg[2][22]/P0001 ,
		_w18070_
	);
	LUT2 #(
		.INIT('h4)
	) name17539 (
		\u0_w_reg[1][22]/P0001 ,
		\u0_w_reg[2][22]/P0001 ,
		_w18071_
	);
	LUT2 #(
		.INIT('h1)
	) name17540 (
		_w18070_,
		_w18071_,
		_w18072_
	);
	LUT2 #(
		.INIT('h8)
	) name17541 (
		_w18069_,
		_w18072_,
		_w18073_
	);
	LUT2 #(
		.INIT('h1)
	) name17542 (
		_w18069_,
		_w18072_,
		_w18074_
	);
	LUT2 #(
		.INIT('h1)
	) name17543 (
		_w18073_,
		_w18074_,
		_w18075_
	);
	LUT2 #(
		.INIT('h4)
	) name17544 (
		ld_pad,
		_w18075_,
		_w18076_
	);
	LUT2 #(
		.INIT('h1)
	) name17545 (
		_w17992_,
		_w18076_,
		_w18077_
	);
	LUT2 #(
		.INIT('h4)
	) name17546 (
		\key[38]_pad ,
		ld_pad,
		_w18078_
	);
	LUT2 #(
		.INIT('h8)
	) name17547 (
		_w16030_,
		_w16386_,
		_w18079_
	);
	LUT2 #(
		.INIT('h2)
	) name17548 (
		\u0_w_reg[3][25]/P0001 ,
		_w18079_,
		_w18080_
	);
	LUT2 #(
		.INIT('h8)
	) name17549 (
		_w17418_,
		_w18080_,
		_w18081_
	);
	LUT2 #(
		.INIT('h8)
	) name17550 (
		_w16019_,
		_w16360_,
		_w18082_
	);
	LUT2 #(
		.INIT('h1)
	) name17551 (
		_w16150_,
		_w17259_,
		_w18083_
	);
	LUT2 #(
		.INIT('h4)
	) name17552 (
		_w18082_,
		_w18083_,
		_w18084_
	);
	LUT2 #(
		.INIT('h8)
	) name17553 (
		_w18081_,
		_w18084_,
		_w18085_
	);
	LUT2 #(
		.INIT('h4)
	) name17554 (
		_w16091_,
		_w17865_,
		_w18086_
	);
	LUT2 #(
		.INIT('h1)
	) name17555 (
		_w16081_,
		_w16158_,
		_w18087_
	);
	LUT2 #(
		.INIT('h8)
	) name17556 (
		_w18086_,
		_w18087_,
		_w18088_
	);
	LUT2 #(
		.INIT('h1)
	) name17557 (
		_w18085_,
		_w18088_,
		_w18089_
	);
	LUT2 #(
		.INIT('h2)
	) name17558 (
		\u0_w_reg[3][26]/P0001 ,
		_w16060_,
		_w18090_
	);
	LUT2 #(
		.INIT('h4)
	) name17559 (
		_w16120_,
		_w16404_,
		_w18091_
	);
	LUT2 #(
		.INIT('h8)
	) name17560 (
		_w18090_,
		_w18091_,
		_w18092_
	);
	LUT2 #(
		.INIT('h4)
	) name17561 (
		_w18089_,
		_w18092_,
		_w18093_
	);
	LUT2 #(
		.INIT('h8)
	) name17562 (
		_w16173_,
		_w18086_,
		_w18094_
	);
	LUT2 #(
		.INIT('h1)
	) name17563 (
		_w18081_,
		_w18094_,
		_w18095_
	);
	LUT2 #(
		.INIT('h4)
	) name17564 (
		_w16134_,
		_w17815_,
		_w18096_
	);
	LUT2 #(
		.INIT('h4)
	) name17565 (
		_w18095_,
		_w18096_,
		_w18097_
	);
	LUT2 #(
		.INIT('h2)
	) name17566 (
		\u0_w_reg[3][24]/P0001 ,
		_w18093_,
		_w18098_
	);
	LUT2 #(
		.INIT('h4)
	) name17567 (
		_w18097_,
		_w18098_,
		_w18099_
	);
	LUT2 #(
		.INIT('h4)
	) name17568 (
		_w16051_,
		_w17401_,
		_w18100_
	);
	LUT2 #(
		.INIT('h1)
	) name17569 (
		\u0_w_reg[3][26]/P0001 ,
		_w16393_,
		_w18101_
	);
	LUT2 #(
		.INIT('h4)
	) name17570 (
		\u0_w_reg[3][27]/P0001 ,
		_w16438_,
		_w18102_
	);
	LUT2 #(
		.INIT('h1)
	) name17571 (
		_w16408_,
		_w18100_,
		_w18103_
	);
	LUT2 #(
		.INIT('h2)
	) name17572 (
		_w18101_,
		_w18102_,
		_w18104_
	);
	LUT2 #(
		.INIT('h8)
	) name17573 (
		_w18103_,
		_w18104_,
		_w18105_
	);
	LUT2 #(
		.INIT('h2)
	) name17574 (
		\u0_w_reg[3][26]/P0001 ,
		_w17450_,
		_w18106_
	);
	LUT2 #(
		.INIT('h4)
	) name17575 (
		_w17327_,
		_w18106_,
		_w18107_
	);
	LUT2 #(
		.INIT('h1)
	) name17576 (
		_w18105_,
		_w18107_,
		_w18108_
	);
	LUT2 #(
		.INIT('h8)
	) name17577 (
		\u0_w_reg[3][31]/P0001 ,
		_w17401_,
		_w18109_
	);
	LUT2 #(
		.INIT('h8)
	) name17578 (
		_w16122_,
		_w17318_,
		_w18110_
	);
	LUT2 #(
		.INIT('h1)
	) name17579 (
		\u0_w_reg[3][25]/P0001 ,
		_w16027_,
		_w18111_
	);
	LUT2 #(
		.INIT('h4)
	) name17580 (
		_w17457_,
		_w18111_,
		_w18112_
	);
	LUT2 #(
		.INIT('h1)
	) name17581 (
		_w17825_,
		_w18109_,
		_w18113_
	);
	LUT2 #(
		.INIT('h4)
	) name17582 (
		_w18110_,
		_w18113_,
		_w18114_
	);
	LUT2 #(
		.INIT('h4)
	) name17583 (
		_w17327_,
		_w18112_,
		_w18115_
	);
	LUT2 #(
		.INIT('h8)
	) name17584 (
		_w18114_,
		_w18115_,
		_w18116_
	);
	LUT2 #(
		.INIT('h4)
	) name17585 (
		\u0_w_reg[3][26]/P0001 ,
		_w16120_,
		_w18117_
	);
	LUT2 #(
		.INIT('h8)
	) name17586 (
		\u0_w_reg[3][28]/P0001 ,
		_w16145_,
		_w18118_
	);
	LUT2 #(
		.INIT('h1)
	) name17587 (
		_w16406_,
		_w18118_,
		_w18119_
	);
	LUT2 #(
		.INIT('h2)
	) name17588 (
		_w16036_,
		_w18119_,
		_w18120_
	);
	LUT2 #(
		.INIT('h2)
	) name17589 (
		\u0_w_reg[3][25]/P0001 ,
		_w16111_,
		_w18121_
	);
	LUT2 #(
		.INIT('h4)
	) name17590 (
		_w18117_,
		_w18121_,
		_w18122_
	);
	LUT2 #(
		.INIT('h4)
	) name17591 (
		_w18120_,
		_w18122_,
		_w18123_
	);
	LUT2 #(
		.INIT('h1)
	) name17592 (
		_w18116_,
		_w18123_,
		_w18124_
	);
	LUT2 #(
		.INIT('h1)
	) name17593 (
		_w18108_,
		_w18124_,
		_w18125_
	);
	LUT2 #(
		.INIT('h1)
	) name17594 (
		\u0_w_reg[3][24]/P0001 ,
		_w18125_,
		_w18126_
	);
	LUT2 #(
		.INIT('h1)
	) name17595 (
		\u0_w_reg[3][26]/P0001 ,
		_w16161_,
		_w18127_
	);
	LUT2 #(
		.INIT('h1)
	) name17596 (
		_w16091_,
		_w17331_,
		_w18128_
	);
	LUT2 #(
		.INIT('h8)
	) name17597 (
		_w18127_,
		_w18128_,
		_w18129_
	);
	LUT2 #(
		.INIT('h8)
	) name17598 (
		_w16032_,
		_w16051_,
		_w18130_
	);
	LUT2 #(
		.INIT('h2)
	) name17599 (
		\u0_w_reg[3][26]/P0001 ,
		_w16428_,
		_w18131_
	);
	LUT2 #(
		.INIT('h4)
	) name17600 (
		_w18130_,
		_w18131_,
		_w18132_
	);
	LUT2 #(
		.INIT('h1)
	) name17601 (
		_w18129_,
		_w18132_,
		_w18133_
	);
	LUT2 #(
		.INIT('h1)
	) name17602 (
		_w16367_,
		_w16375_,
		_w18134_
	);
	LUT2 #(
		.INIT('h4)
	) name17603 (
		_w18133_,
		_w18134_,
		_w18135_
	);
	LUT2 #(
		.INIT('h1)
	) name17604 (
		\u0_w_reg[3][25]/P0001 ,
		_w18135_,
		_w18136_
	);
	LUT2 #(
		.INIT('h1)
	) name17605 (
		_w16449_,
		_w17402_,
		_w18137_
	);
	LUT2 #(
		.INIT('h2)
	) name17606 (
		\u0_w_reg[3][26]/P0001 ,
		_w18137_,
		_w18138_
	);
	LUT2 #(
		.INIT('h8)
	) name17607 (
		\u0_w_reg[3][25]/P0001 ,
		_w16119_,
		_w18139_
	);
	LUT2 #(
		.INIT('h1)
	) name17608 (
		_w16169_,
		_w17337_,
		_w18140_
	);
	LUT2 #(
		.INIT('h1)
	) name17609 (
		\u0_w_reg[3][30]/P0001 ,
		_w18140_,
		_w18141_
	);
	LUT2 #(
		.INIT('h1)
	) name17610 (
		_w16088_,
		_w18141_,
		_w18142_
	);
	LUT2 #(
		.INIT('h2)
	) name17611 (
		_w17871_,
		_w18142_,
		_w18143_
	);
	LUT2 #(
		.INIT('h1)
	) name17612 (
		_w16420_,
		_w17463_,
		_w18144_
	);
	LUT2 #(
		.INIT('h4)
	) name17613 (
		_w18139_,
		_w18144_,
		_w18145_
	);
	LUT2 #(
		.INIT('h4)
	) name17614 (
		_w18138_,
		_w18145_,
		_w18146_
	);
	LUT2 #(
		.INIT('h4)
	) name17615 (
		_w18143_,
		_w18146_,
		_w18147_
	);
	LUT2 #(
		.INIT('h4)
	) name17616 (
		_w18136_,
		_w18147_,
		_w18148_
	);
	LUT2 #(
		.INIT('h4)
	) name17617 (
		_w18126_,
		_w18148_,
		_w18149_
	);
	LUT2 #(
		.INIT('h4)
	) name17618 (
		_w18099_,
		_w18149_,
		_w18150_
	);
	LUT2 #(
		.INIT('h2)
	) name17619 (
		\u0_w_reg[0][6]/P0001 ,
		_w18150_,
		_w18151_
	);
	LUT2 #(
		.INIT('h4)
	) name17620 (
		\u0_w_reg[0][6]/P0001 ,
		_w18150_,
		_w18152_
	);
	LUT2 #(
		.INIT('h1)
	) name17621 (
		_w18151_,
		_w18152_,
		_w18153_
	);
	LUT2 #(
		.INIT('h2)
	) name17622 (
		\u0_w_reg[1][6]/P0001 ,
		\u0_w_reg[2][6]/P0001 ,
		_w18154_
	);
	LUT2 #(
		.INIT('h4)
	) name17623 (
		\u0_w_reg[1][6]/P0001 ,
		\u0_w_reg[2][6]/P0001 ,
		_w18155_
	);
	LUT2 #(
		.INIT('h1)
	) name17624 (
		_w18154_,
		_w18155_,
		_w18156_
	);
	LUT2 #(
		.INIT('h8)
	) name17625 (
		_w18153_,
		_w18156_,
		_w18157_
	);
	LUT2 #(
		.INIT('h1)
	) name17626 (
		_w18153_,
		_w18156_,
		_w18158_
	);
	LUT2 #(
		.INIT('h1)
	) name17627 (
		_w18157_,
		_w18158_,
		_w18159_
	);
	LUT2 #(
		.INIT('h4)
	) name17628 (
		ld_pad,
		_w18159_,
		_w18160_
	);
	LUT2 #(
		.INIT('h1)
	) name17629 (
		_w18078_,
		_w18160_,
		_w18161_
	);
	LUT2 #(
		.INIT('h4)
	) name17630 (
		\key[45]_pad ,
		ld_pad,
		_w18162_
	);
	LUT2 #(
		.INIT('h8)
	) name17631 (
		\u0_w_reg[3][4]/P0001 ,
		_w16480_,
		_w18163_
	);
	LUT2 #(
		.INIT('h1)
	) name17632 (
		\u0_w_reg[3][4]/P0001 ,
		_w16482_,
		_w18164_
	);
	LUT2 #(
		.INIT('h4)
	) name17633 (
		_w16521_,
		_w18164_,
		_w18165_
	);
	LUT2 #(
		.INIT('h1)
	) name17634 (
		_w18163_,
		_w18165_,
		_w18166_
	);
	LUT2 #(
		.INIT('h2)
	) name17635 (
		\u0_w_reg[3][1]/P0001 ,
		_w18166_,
		_w18167_
	);
	LUT2 #(
		.INIT('h1)
	) name17636 (
		_w16657_,
		_w16728_,
		_w18168_
	);
	LUT2 #(
		.INIT('h1)
	) name17637 (
		\u0_w_reg[3][2]/P0001 ,
		_w16596_,
		_w18169_
	);
	LUT2 #(
		.INIT('h8)
	) name17638 (
		_w18168_,
		_w18169_,
		_w18170_
	);
	LUT2 #(
		.INIT('h4)
	) name17639 (
		_w18167_,
		_w18170_,
		_w18171_
	);
	LUT2 #(
		.INIT('h2)
	) name17640 (
		\u0_w_reg[3][2]/P0001 ,
		_w16523_,
		_w18172_
	);
	LUT2 #(
		.INIT('h4)
	) name17641 (
		_w16530_,
		_w18172_,
		_w18173_
	);
	LUT2 #(
		.INIT('h1)
	) name17642 (
		_w18171_,
		_w18173_,
		_w18174_
	);
	LUT2 #(
		.INIT('h8)
	) name17643 (
		_w16570_,
		_w16612_,
		_w18175_
	);
	LUT2 #(
		.INIT('h1)
	) name17644 (
		_w16564_,
		_w17959_,
		_w18176_
	);
	LUT2 #(
		.INIT('h2)
	) name17645 (
		\u0_w_reg[3][1]/P0001 ,
		_w18175_,
		_w18177_
	);
	LUT2 #(
		.INIT('h4)
	) name17646 (
		_w16624_,
		_w18177_,
		_w18178_
	);
	LUT2 #(
		.INIT('h8)
	) name17647 (
		_w18176_,
		_w18178_,
		_w18179_
	);
	LUT2 #(
		.INIT('h8)
	) name17648 (
		_w16495_,
		_w16586_,
		_w18180_
	);
	LUT2 #(
		.INIT('h1)
	) name17649 (
		\u0_w_reg[3][1]/P0001 ,
		_w18180_,
		_w18181_
	);
	LUT2 #(
		.INIT('h1)
	) name17650 (
		_w16650_,
		_w16700_,
		_w18182_
	);
	LUT2 #(
		.INIT('h2)
	) name17651 (
		\u0_w_reg[3][2]/P0001 ,
		_w18182_,
		_w18183_
	);
	LUT2 #(
		.INIT('h4)
	) name17652 (
		\u0_w_reg[3][2]/P0001 ,
		_w16494_,
		_w18184_
	);
	LUT2 #(
		.INIT('h1)
	) name17653 (
		_w16530_,
		_w16728_,
		_w18185_
	);
	LUT2 #(
		.INIT('h2)
	) name17654 (
		_w18181_,
		_w18184_,
		_w18186_
	);
	LUT2 #(
		.INIT('h8)
	) name17655 (
		_w18185_,
		_w18186_,
		_w18187_
	);
	LUT2 #(
		.INIT('h4)
	) name17656 (
		_w18183_,
		_w18187_,
		_w18188_
	);
	LUT2 #(
		.INIT('h1)
	) name17657 (
		_w18179_,
		_w18188_,
		_w18189_
	);
	LUT2 #(
		.INIT('h1)
	) name17658 (
		_w16597_,
		_w16696_,
		_w18190_
	);
	LUT2 #(
		.INIT('h4)
	) name17659 (
		_w18174_,
		_w18190_,
		_w18191_
	);
	LUT2 #(
		.INIT('h4)
	) name17660 (
		_w18189_,
		_w18191_,
		_w18192_
	);
	LUT2 #(
		.INIT('h2)
	) name17661 (
		\u0_w_reg[3][0]/P0001 ,
		_w18192_,
		_w18193_
	);
	LUT2 #(
		.INIT('h8)
	) name17662 (
		\u0_w_reg[3][3]/P0001 ,
		_w16570_,
		_w18194_
	);
	LUT2 #(
		.INIT('h1)
	) name17663 (
		_w16607_,
		_w17952_,
		_w18195_
	);
	LUT2 #(
		.INIT('h1)
	) name17664 (
		\u0_w_reg[3][3]/P0001 ,
		_w18195_,
		_w18196_
	);
	LUT2 #(
		.INIT('h1)
	) name17665 (
		_w18194_,
		_w18196_,
		_w18197_
	);
	LUT2 #(
		.INIT('h1)
	) name17666 (
		\u0_w_reg[3][2]/P0001 ,
		_w18197_,
		_w18198_
	);
	LUT2 #(
		.INIT('h1)
	) name17667 (
		_w16556_,
		_w16688_,
		_w18199_
	);
	LUT2 #(
		.INIT('h1)
	) name17668 (
		\u0_w_reg[3][7]/P0001 ,
		_w18199_,
		_w18200_
	);
	LUT2 #(
		.INIT('h4)
	) name17669 (
		_w16554_,
		_w16565_,
		_w18201_
	);
	LUT2 #(
		.INIT('h1)
	) name17670 (
		_w16490_,
		_w16701_,
		_w18202_
	);
	LUT2 #(
		.INIT('h4)
	) name17671 (
		_w16543_,
		_w18202_,
		_w18203_
	);
	LUT2 #(
		.INIT('h4)
	) name17672 (
		_w18201_,
		_w18203_,
		_w18204_
	);
	LUT2 #(
		.INIT('h4)
	) name17673 (
		_w18200_,
		_w18204_,
		_w18205_
	);
	LUT2 #(
		.INIT('h4)
	) name17674 (
		_w18198_,
		_w18205_,
		_w18206_
	);
	LUT2 #(
		.INIT('h2)
	) name17675 (
		\u0_w_reg[3][1]/P0001 ,
		_w18206_,
		_w18207_
	);
	LUT2 #(
		.INIT('h1)
	) name17676 (
		_w16665_,
		_w17573_,
		_w18208_
	);
	LUT2 #(
		.INIT('h1)
	) name17677 (
		\u0_w_reg[3][5]/P0001 ,
		_w18208_,
		_w18209_
	);
	LUT2 #(
		.INIT('h8)
	) name17678 (
		\u0_w_reg[3][2]/P0001 ,
		_w16623_,
		_w18210_
	);
	LUT2 #(
		.INIT('h1)
	) name17679 (
		_w16479_,
		_w18210_,
		_w18211_
	);
	LUT2 #(
		.INIT('h4)
	) name17680 (
		_w18209_,
		_w18211_,
		_w18212_
	);
	LUT2 #(
		.INIT('h1)
	) name17681 (
		\u0_w_reg[3][1]/P0001 ,
		_w18212_,
		_w18213_
	);
	LUT2 #(
		.INIT('h2)
	) name17682 (
		\u0_w_reg[3][3]/P0001 ,
		_w17916_,
		_w18214_
	);
	LUT2 #(
		.INIT('h8)
	) name17683 (
		_w16521_,
		_w16668_,
		_w18215_
	);
	LUT2 #(
		.INIT('h1)
	) name17684 (
		_w17519_,
		_w18215_,
		_w18216_
	);
	LUT2 #(
		.INIT('h4)
	) name17685 (
		_w18214_,
		_w18216_,
		_w18217_
	);
	LUT2 #(
		.INIT('h2)
	) name17686 (
		\u0_w_reg[3][2]/P0001 ,
		_w18217_,
		_w18218_
	);
	LUT2 #(
		.INIT('h1)
	) name17687 (
		_w16659_,
		_w17935_,
		_w18219_
	);
	LUT2 #(
		.INIT('h4)
	) name17688 (
		_w17945_,
		_w18219_,
		_w18220_
	);
	LUT2 #(
		.INIT('h4)
	) name17689 (
		_w18218_,
		_w18220_,
		_w18221_
	);
	LUT2 #(
		.INIT('h4)
	) name17690 (
		_w18213_,
		_w18221_,
		_w18222_
	);
	LUT2 #(
		.INIT('h4)
	) name17691 (
		_w18207_,
		_w18222_,
		_w18223_
	);
	LUT2 #(
		.INIT('h1)
	) name17692 (
		\u0_w_reg[3][0]/P0001 ,
		_w18223_,
		_w18224_
	);
	LUT2 #(
		.INIT('h8)
	) name17693 (
		\u0_w_reg[3][3]/P0001 ,
		_w17952_,
		_w18225_
	);
	LUT2 #(
		.INIT('h4)
	) name17694 (
		\u0_w_reg[3][5]/P0001 ,
		_w16570_,
		_w18226_
	);
	LUT2 #(
		.INIT('h1)
	) name17695 (
		_w16522_,
		_w17501_,
		_w18227_
	);
	LUT2 #(
		.INIT('h4)
	) name17696 (
		_w18226_,
		_w18227_,
		_w18228_
	);
	LUT2 #(
		.INIT('h2)
	) name17697 (
		_w16667_,
		_w18228_,
		_w18229_
	);
	LUT2 #(
		.INIT('h1)
	) name17698 (
		_w18225_,
		_w18229_,
		_w18230_
	);
	LUT2 #(
		.INIT('h2)
	) name17699 (
		\u0_w_reg[3][2]/P0001 ,
		_w18230_,
		_w18231_
	);
	LUT2 #(
		.INIT('h8)
	) name17700 (
		_w16588_,
		_w16649_,
		_w18232_
	);
	LUT2 #(
		.INIT('h8)
	) name17701 (
		_w16509_,
		_w16728_,
		_w18233_
	);
	LUT2 #(
		.INIT('h1)
	) name17702 (
		_w16549_,
		_w16696_,
		_w18234_
	);
	LUT2 #(
		.INIT('h1)
	) name17703 (
		_w18232_,
		_w18233_,
		_w18235_
	);
	LUT2 #(
		.INIT('h8)
	) name17704 (
		_w18234_,
		_w18235_,
		_w18236_
	);
	LUT2 #(
		.INIT('h4)
	) name17705 (
		_w18231_,
		_w18236_,
		_w18237_
	);
	LUT2 #(
		.INIT('h1)
	) name17706 (
		\u0_w_reg[3][1]/P0001 ,
		_w18237_,
		_w18238_
	);
	LUT2 #(
		.INIT('h1)
	) name17707 (
		_w16543_,
		_w16676_,
		_w18239_
	);
	LUT2 #(
		.INIT('h1)
	) name17708 (
		\u0_w_reg[3][2]/P0001 ,
		_w18239_,
		_w18240_
	);
	LUT2 #(
		.INIT('h8)
	) name17709 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		_w18241_
	);
	LUT2 #(
		.INIT('h8)
	) name17710 (
		_w16485_,
		_w18241_,
		_w18242_
	);
	LUT2 #(
		.INIT('h8)
	) name17711 (
		\u0_w_reg[3][3]/P0001 ,
		_w16659_,
		_w18243_
	);
	LUT2 #(
		.INIT('h1)
	) name17712 (
		_w17935_,
		_w18243_,
		_w18244_
	);
	LUT2 #(
		.INIT('h2)
	) name17713 (
		\u0_w_reg[3][1]/P0001 ,
		_w18244_,
		_w18245_
	);
	LUT2 #(
		.INIT('h8)
	) name17714 (
		_w16506_,
		_w18225_,
		_w18246_
	);
	LUT2 #(
		.INIT('h1)
	) name17715 (
		_w18242_,
		_w18246_,
		_w18247_
	);
	LUT2 #(
		.INIT('h4)
	) name17716 (
		_w18240_,
		_w18247_,
		_w18248_
	);
	LUT2 #(
		.INIT('h4)
	) name17717 (
		_w18245_,
		_w18248_,
		_w18249_
	);
	LUT2 #(
		.INIT('h4)
	) name17718 (
		_w18238_,
		_w18249_,
		_w18250_
	);
	LUT2 #(
		.INIT('h4)
	) name17719 (
		_w18193_,
		_w18250_,
		_w18251_
	);
	LUT2 #(
		.INIT('h4)
	) name17720 (
		_w18224_,
		_w18251_,
		_w18252_
	);
	LUT2 #(
		.INIT('h2)
	) name17721 (
		\u0_w_reg[0][13]/P0001 ,
		_w18252_,
		_w18253_
	);
	LUT2 #(
		.INIT('h4)
	) name17722 (
		\u0_w_reg[0][13]/P0001 ,
		_w18252_,
		_w18254_
	);
	LUT2 #(
		.INIT('h1)
	) name17723 (
		_w18253_,
		_w18254_,
		_w18255_
	);
	LUT2 #(
		.INIT('h2)
	) name17724 (
		\u0_w_reg[1][13]/P0001 ,
		\u0_w_reg[2][13]/P0001 ,
		_w18256_
	);
	LUT2 #(
		.INIT('h4)
	) name17725 (
		\u0_w_reg[1][13]/P0001 ,
		\u0_w_reg[2][13]/P0001 ,
		_w18257_
	);
	LUT2 #(
		.INIT('h1)
	) name17726 (
		_w18256_,
		_w18257_,
		_w18258_
	);
	LUT2 #(
		.INIT('h8)
	) name17727 (
		_w18255_,
		_w18258_,
		_w18259_
	);
	LUT2 #(
		.INIT('h1)
	) name17728 (
		_w18255_,
		_w18258_,
		_w18260_
	);
	LUT2 #(
		.INIT('h1)
	) name17729 (
		_w18259_,
		_w18260_,
		_w18261_
	);
	LUT2 #(
		.INIT('h4)
	) name17730 (
		ld_pad,
		_w18261_,
		_w18262_
	);
	LUT2 #(
		.INIT('h1)
	) name17731 (
		_w18162_,
		_w18262_,
		_w18263_
	);
	LUT2 #(
		.INIT('h8)
	) name17732 (
		_w16512_,
		_w17566_,
		_w18264_
	);
	LUT2 #(
		.INIT('h1)
	) name17733 (
		_w16505_,
		_w16522_,
		_w18265_
	);
	LUT2 #(
		.INIT('h2)
	) name17734 (
		_w17516_,
		_w18265_,
		_w18266_
	);
	LUT2 #(
		.INIT('h2)
	) name17735 (
		_w17531_,
		_w17897_,
		_w18267_
	);
	LUT2 #(
		.INIT('h4)
	) name17736 (
		_w18264_,
		_w18267_,
		_w18268_
	);
	LUT2 #(
		.INIT('h4)
	) name17737 (
		_w18266_,
		_w18268_,
		_w18269_
	);
	LUT2 #(
		.INIT('h8)
	) name17738 (
		_w16493_,
		_w16506_,
		_w18270_
	);
	LUT2 #(
		.INIT('h8)
	) name17739 (
		_w16524_,
		_w16582_,
		_w18271_
	);
	LUT2 #(
		.INIT('h1)
	) name17740 (
		\u0_w_reg[3][1]/P0001 ,
		_w17958_,
		_w18272_
	);
	LUT2 #(
		.INIT('h4)
	) name17741 (
		_w18270_,
		_w18272_,
		_w18273_
	);
	LUT2 #(
		.INIT('h4)
	) name17742 (
		_w18271_,
		_w18273_,
		_w18274_
	);
	LUT2 #(
		.INIT('h1)
	) name17743 (
		_w18269_,
		_w18274_,
		_w18275_
	);
	LUT2 #(
		.INIT('h1)
	) name17744 (
		_w16596_,
		_w17501_,
		_w18276_
	);
	LUT2 #(
		.INIT('h2)
	) name17745 (
		_w16588_,
		_w18276_,
		_w18277_
	);
	LUT2 #(
		.INIT('h8)
	) name17746 (
		_w16489_,
		_w16603_,
		_w18278_
	);
	LUT2 #(
		.INIT('h8)
	) name17747 (
		_w16495_,
		_w16528_,
		_w18279_
	);
	LUT2 #(
		.INIT('h1)
	) name17748 (
		_w16659_,
		_w18279_,
		_w18280_
	);
	LUT2 #(
		.INIT('h2)
	) name17749 (
		_w16524_,
		_w18280_,
		_w18281_
	);
	LUT2 #(
		.INIT('h8)
	) name17750 (
		\u0_w_reg[3][4]/P0001 ,
		_w16587_,
		_w18282_
	);
	LUT2 #(
		.INIT('h1)
	) name17751 (
		\u0_w_reg[3][0]/P0001 ,
		_w18278_,
		_w18283_
	);
	LUT2 #(
		.INIT('h4)
	) name17752 (
		_w18233_,
		_w18283_,
		_w18284_
	);
	LUT2 #(
		.INIT('h4)
	) name17753 (
		_w18282_,
		_w18284_,
		_w18285_
	);
	LUT2 #(
		.INIT('h1)
	) name17754 (
		_w18246_,
		_w18277_,
		_w18286_
	);
	LUT2 #(
		.INIT('h4)
	) name17755 (
		_w18281_,
		_w18286_,
		_w18287_
	);
	LUT2 #(
		.INIT('h8)
	) name17756 (
		_w18285_,
		_w18287_,
		_w18288_
	);
	LUT2 #(
		.INIT('h4)
	) name17757 (
		_w18275_,
		_w18288_,
		_w18289_
	);
	LUT2 #(
		.INIT('h2)
	) name17758 (
		\u0_w_reg[3][2]/P0001 ,
		_w16504_,
		_w18290_
	);
	LUT2 #(
		.INIT('h1)
	) name17759 (
		\u0_w_reg[3][2]/P0001 ,
		_w16608_,
		_w18291_
	);
	LUT2 #(
		.INIT('h1)
	) name17760 (
		_w16687_,
		_w17961_,
		_w18292_
	);
	LUT2 #(
		.INIT('h8)
	) name17761 (
		_w18291_,
		_w18292_,
		_w18293_
	);
	LUT2 #(
		.INIT('h1)
	) name17762 (
		_w18290_,
		_w18293_,
		_w18294_
	);
	LUT2 #(
		.INIT('h4)
	) name17763 (
		\u0_w_reg[3][3]/P0001 ,
		_w16483_,
		_w18295_
	);
	LUT2 #(
		.INIT('h4)
	) name17764 (
		_w16552_,
		_w18295_,
		_w18296_
	);
	LUT2 #(
		.INIT('h4)
	) name17765 (
		_w16729_,
		_w18181_,
		_w18297_
	);
	LUT2 #(
		.INIT('h4)
	) name17766 (
		_w18296_,
		_w18297_,
		_w18298_
	);
	LUT2 #(
		.INIT('h4)
	) name17767 (
		_w18294_,
		_w18298_,
		_w18299_
	);
	LUT2 #(
		.INIT('h8)
	) name17768 (
		\u0_w_reg[3][3]/P0001 ,
		_w16483_,
		_w18300_
	);
	LUT2 #(
		.INIT('h1)
	) name17769 (
		_w16477_,
		_w16608_,
		_w18301_
	);
	LUT2 #(
		.INIT('h1)
	) name17770 (
		_w16622_,
		_w18300_,
		_w18302_
	);
	LUT2 #(
		.INIT('h8)
	) name17771 (
		_w18301_,
		_w18302_,
		_w18303_
	);
	LUT2 #(
		.INIT('h2)
	) name17772 (
		\u0_w_reg[3][2]/P0001 ,
		_w18303_,
		_w18304_
	);
	LUT2 #(
		.INIT('h8)
	) name17773 (
		_w16588_,
		_w18226_,
		_w18305_
	);
	LUT2 #(
		.INIT('h8)
	) name17774 (
		_w16496_,
		_w16521_,
		_w18306_
	);
	LUT2 #(
		.INIT('h2)
	) name17775 (
		\u0_w_reg[3][1]/P0001 ,
		_w18305_,
		_w18307_
	);
	LUT2 #(
		.INIT('h4)
	) name17776 (
		_w18306_,
		_w18307_,
		_w18308_
	);
	LUT2 #(
		.INIT('h4)
	) name17777 (
		_w18304_,
		_w18308_,
		_w18309_
	);
	LUT2 #(
		.INIT('h1)
	) name17778 (
		_w18299_,
		_w18309_,
		_w18310_
	);
	LUT2 #(
		.INIT('h1)
	) name17779 (
		_w16550_,
		_w16589_,
		_w18311_
	);
	LUT2 #(
		.INIT('h2)
	) name17780 (
		\u0_w_reg[3][4]/P0001 ,
		_w18311_,
		_w18312_
	);
	LUT2 #(
		.INIT('h8)
	) name17781 (
		_w16524_,
		_w16700_,
		_w18313_
	);
	LUT2 #(
		.INIT('h4)
	) name17782 (
		\u0_w_reg[3][4]/P0001 ,
		_w16541_,
		_w18314_
	);
	LUT2 #(
		.INIT('h1)
	) name17783 (
		_w17952_,
		_w18314_,
		_w18315_
	);
	LUT2 #(
		.INIT('h2)
	) name17784 (
		_w16512_,
		_w18315_,
		_w18316_
	);
	LUT2 #(
		.INIT('h8)
	) name17785 (
		\u0_w_reg[3][5]/P0001 ,
		_w16668_,
		_w18317_
	);
	LUT2 #(
		.INIT('h2)
	) name17786 (
		\u0_w_reg[3][0]/P0001 ,
		_w18313_,
		_w18318_
	);
	LUT2 #(
		.INIT('h4)
	) name17787 (
		_w18317_,
		_w18318_,
		_w18319_
	);
	LUT2 #(
		.INIT('h1)
	) name17788 (
		_w18312_,
		_w18316_,
		_w18320_
	);
	LUT2 #(
		.INIT('h8)
	) name17789 (
		_w18319_,
		_w18320_,
		_w18321_
	);
	LUT2 #(
		.INIT('h4)
	) name17790 (
		_w18310_,
		_w18321_,
		_w18322_
	);
	LUT2 #(
		.INIT('h1)
	) name17791 (
		_w18289_,
		_w18322_,
		_w18323_
	);
	LUT2 #(
		.INIT('h8)
	) name17792 (
		_w16521_,
		_w16658_,
		_w18324_
	);
	LUT2 #(
		.INIT('h1)
	) name17793 (
		_w16478_,
		_w18324_,
		_w18325_
	);
	LUT2 #(
		.INIT('h2)
	) name17794 (
		_w16488_,
		_w16489_,
		_w18326_
	);
	LUT2 #(
		.INIT('h2)
	) name17795 (
		_w18325_,
		_w18326_,
		_w18327_
	);
	LUT2 #(
		.INIT('h2)
	) name17796 (
		\u0_w_reg[3][3]/P0001 ,
		_w18327_,
		_w18328_
	);
	LUT2 #(
		.INIT('h1)
	) name17797 (
		\u0_w_reg[3][2]/P0001 ,
		_w18328_,
		_w18329_
	);
	LUT2 #(
		.INIT('h1)
	) name17798 (
		_w16575_,
		_w16697_,
		_w18330_
	);
	LUT2 #(
		.INIT('h4)
	) name17799 (
		_w18314_,
		_w18330_,
		_w18331_
	);
	LUT2 #(
		.INIT('h1)
	) name17800 (
		\u0_w_reg[3][3]/P0001 ,
		_w18331_,
		_w18332_
	);
	LUT2 #(
		.INIT('h2)
	) name17801 (
		\u0_w_reg[3][2]/P0001 ,
		_w16627_,
		_w18333_
	);
	LUT2 #(
		.INIT('h4)
	) name17802 (
		_w16728_,
		_w18333_,
		_w18334_
	);
	LUT2 #(
		.INIT('h4)
	) name17803 (
		_w18332_,
		_w18334_,
		_w18335_
	);
	LUT2 #(
		.INIT('h2)
	) name17804 (
		\u0_w_reg[3][1]/P0001 ,
		_w18329_,
		_w18336_
	);
	LUT2 #(
		.INIT('h4)
	) name17805 (
		_w18335_,
		_w18336_,
		_w18337_
	);
	LUT2 #(
		.INIT('h4)
	) name17806 (
		\u0_w_reg[3][2]/P0001 ,
		_w17907_,
		_w18338_
	);
	LUT2 #(
		.INIT('h1)
	) name17807 (
		_w16529_,
		_w18277_,
		_w18339_
	);
	LUT2 #(
		.INIT('h4)
	) name17808 (
		_w18338_,
		_w18339_,
		_w18340_
	);
	LUT2 #(
		.INIT('h1)
	) name17809 (
		\u0_w_reg[3][1]/P0001 ,
		_w18340_,
		_w18341_
	);
	LUT2 #(
		.INIT('h8)
	) name17810 (
		_w17516_,
		_w17927_,
		_w18342_
	);
	LUT2 #(
		.INIT('h8)
	) name17811 (
		_w16621_,
		_w16687_,
		_w18343_
	);
	LUT2 #(
		.INIT('h1)
	) name17812 (
		_w17970_,
		_w18343_,
		_w18344_
	);
	LUT2 #(
		.INIT('h1)
	) name17813 (
		\u0_w_reg[3][3]/P0001 ,
		_w18344_,
		_w18345_
	);
	LUT2 #(
		.INIT('h1)
	) name17814 (
		_w16701_,
		_w18306_,
		_w18346_
	);
	LUT2 #(
		.INIT('h2)
	) name17815 (
		_w16621_,
		_w18346_,
		_w18347_
	);
	LUT2 #(
		.INIT('h1)
	) name17816 (
		_w18342_,
		_w18345_,
		_w18348_
	);
	LUT2 #(
		.INIT('h4)
	) name17817 (
		_w18347_,
		_w18348_,
		_w18349_
	);
	LUT2 #(
		.INIT('h4)
	) name17818 (
		_w18341_,
		_w18349_,
		_w18350_
	);
	LUT2 #(
		.INIT('h4)
	) name17819 (
		_w18337_,
		_w18350_,
		_w18351_
	);
	LUT2 #(
		.INIT('h4)
	) name17820 (
		_w18323_,
		_w18351_,
		_w18352_
	);
	LUT2 #(
		.INIT('h2)
	) name17821 (
		\u0_w_reg[0][15]/P0001 ,
		_w18352_,
		_w18353_
	);
	LUT2 #(
		.INIT('h4)
	) name17822 (
		\u0_w_reg[0][15]/P0001 ,
		_w18352_,
		_w18354_
	);
	LUT2 #(
		.INIT('h1)
	) name17823 (
		_w18353_,
		_w18354_,
		_w18355_
	);
	LUT2 #(
		.INIT('h8)
	) name17824 (
		\u0_w_reg[1][15]/P0001 ,
		_w18355_,
		_w18356_
	);
	LUT2 #(
		.INIT('h1)
	) name17825 (
		\u0_w_reg[1][15]/P0001 ,
		_w18355_,
		_w18357_
	);
	LUT2 #(
		.INIT('h1)
	) name17826 (
		_w18356_,
		_w18357_,
		_w18358_
	);
	LUT2 #(
		.INIT('h8)
	) name17827 (
		\u0_w_reg[2][15]/P0001 ,
		_w18358_,
		_w18359_
	);
	LUT2 #(
		.INIT('h1)
	) name17828 (
		\u0_w_reg[2][15]/P0001 ,
		_w18358_,
		_w18360_
	);
	LUT2 #(
		.INIT('h1)
	) name17829 (
		_w18359_,
		_w18360_,
		_w18361_
	);
	LUT2 #(
		.INIT('h4)
	) name17830 (
		ld_pad,
		_w18361_,
		_w18362_
	);
	LUT2 #(
		.INIT('h8)
	) name17831 (
		\key[47]_pad ,
		ld_pad,
		_w18363_
	);
	LUT2 #(
		.INIT('h1)
	) name17832 (
		_w18362_,
		_w18363_,
		_w18364_
	);
	LUT2 #(
		.INIT('h4)
	) name17833 (
		\key[40]_pad ,
		ld_pad,
		_w18365_
	);
	LUT2 #(
		.INIT('h4)
	) name17834 (
		\u0_w_reg[3][3]/P0001 ,
		_w17517_,
		_w18366_
	);
	LUT2 #(
		.INIT('h1)
	) name17835 (
		_w16494_,
		_w18215_,
		_w18367_
	);
	LUT2 #(
		.INIT('h4)
	) name17836 (
		_w18366_,
		_w18367_,
		_w18368_
	);
	LUT2 #(
		.INIT('h2)
	) name17837 (
		\u0_w_reg[3][2]/P0001 ,
		_w18368_,
		_w18369_
	);
	LUT2 #(
		.INIT('h4)
	) name17838 (
		\u0_w_reg[3][2]/P0001 ,
		_w16529_,
		_w18370_
	);
	LUT2 #(
		.INIT('h2)
	) name17839 (
		\u0_w_reg[3][1]/P0001 ,
		_w16660_,
		_w18371_
	);
	LUT2 #(
		.INIT('h1)
	) name17840 (
		_w16676_,
		_w18370_,
		_w18372_
	);
	LUT2 #(
		.INIT('h8)
	) name17841 (
		_w18371_,
		_w18372_,
		_w18373_
	);
	LUT2 #(
		.INIT('h4)
	) name17842 (
		_w18369_,
		_w18373_,
		_w18374_
	);
	LUT2 #(
		.INIT('h1)
	) name17843 (
		_w16556_,
		_w17959_,
		_w18375_
	);
	LUT2 #(
		.INIT('h8)
	) name17844 (
		_w16731_,
		_w18375_,
		_w18376_
	);
	LUT2 #(
		.INIT('h1)
	) name17845 (
		_w16522_,
		_w17961_,
		_w18377_
	);
	LUT2 #(
		.INIT('h1)
	) name17846 (
		\u0_w_reg[3][3]/P0001 ,
		_w18377_,
		_w18378_
	);
	LUT2 #(
		.INIT('h1)
	) name17847 (
		\u0_w_reg[3][2]/P0001 ,
		_w17506_,
		_w18379_
	);
	LUT2 #(
		.INIT('h4)
	) name17848 (
		_w18378_,
		_w18379_,
		_w18380_
	);
	LUT2 #(
		.INIT('h1)
	) name17849 (
		_w18376_,
		_w18380_,
		_w18381_
	);
	LUT2 #(
		.INIT('h1)
	) name17850 (
		\u0_w_reg[3][1]/P0001 ,
		_w17518_,
		_w18382_
	);
	LUT2 #(
		.INIT('h4)
	) name17851 (
		_w18381_,
		_w18382_,
		_w18383_
	);
	LUT2 #(
		.INIT('h1)
	) name17852 (
		_w18374_,
		_w18383_,
		_w18384_
	);
	LUT2 #(
		.INIT('h8)
	) name17853 (
		_w16509_,
		_w17532_,
		_w18385_
	);
	LUT2 #(
		.INIT('h2)
	) name17854 (
		_w16567_,
		_w17896_,
		_w18386_
	);
	LUT2 #(
		.INIT('h1)
	) name17855 (
		\u0_w_reg[3][2]/P0001 ,
		_w18386_,
		_w18387_
	);
	LUT2 #(
		.INIT('h1)
	) name17856 (
		_w16521_,
		_w16753_,
		_w18388_
	);
	LUT2 #(
		.INIT('h2)
	) name17857 (
		_w16664_,
		_w18388_,
		_w18389_
	);
	LUT2 #(
		.INIT('h4)
	) name17858 (
		\u0_w_reg[3][2]/P0001 ,
		_w16650_,
		_w18390_
	);
	LUT2 #(
		.INIT('h1)
	) name17859 (
		\u0_w_reg[3][3]/P0001 ,
		_w18325_,
		_w18391_
	);
	LUT2 #(
		.INIT('h2)
	) name17860 (
		_w16526_,
		_w16544_,
		_w18392_
	);
	LUT2 #(
		.INIT('h1)
	) name17861 (
		\u0_w_reg[3][1]/P0001 ,
		_w18390_,
		_w18393_
	);
	LUT2 #(
		.INIT('h4)
	) name17862 (
		_w18392_,
		_w18393_,
		_w18394_
	);
	LUT2 #(
		.INIT('h4)
	) name17863 (
		_w18391_,
		_w18394_,
		_w18395_
	);
	LUT2 #(
		.INIT('h8)
	) name17864 (
		\u0_w_reg[3][4]/P0001 ,
		_w16541_,
		_w18396_
	);
	LUT2 #(
		.INIT('h1)
	) name17865 (
		_w16550_,
		_w18396_,
		_w18397_
	);
	LUT2 #(
		.INIT('h2)
	) name17866 (
		\u0_w_reg[3][3]/P0001 ,
		_w18397_,
		_w18398_
	);
	LUT2 #(
		.INIT('h8)
	) name17867 (
		_w16574_,
		_w16588_,
		_w18399_
	);
	LUT2 #(
		.INIT('h2)
	) name17868 (
		\u0_w_reg[3][1]/P0001 ,
		_w16622_,
		_w18400_
	);
	LUT2 #(
		.INIT('h1)
	) name17869 (
		_w17519_,
		_w18399_,
		_w18401_
	);
	LUT2 #(
		.INIT('h8)
	) name17870 (
		_w18400_,
		_w18401_,
		_w18402_
	);
	LUT2 #(
		.INIT('h4)
	) name17871 (
		_w18398_,
		_w18402_,
		_w18403_
	);
	LUT2 #(
		.INIT('h1)
	) name17872 (
		_w18395_,
		_w18403_,
		_w18404_
	);
	LUT2 #(
		.INIT('h1)
	) name17873 (
		\u0_w_reg[3][0]/P0001 ,
		_w18389_,
		_w18405_
	);
	LUT2 #(
		.INIT('h4)
	) name17874 (
		_w18387_,
		_w18405_,
		_w18406_
	);
	LUT2 #(
		.INIT('h4)
	) name17875 (
		_w18404_,
		_w18406_,
		_w18407_
	);
	LUT2 #(
		.INIT('h1)
	) name17876 (
		_w16675_,
		_w18279_,
		_w18408_
	);
	LUT2 #(
		.INIT('h8)
	) name17877 (
		_w17534_,
		_w18408_,
		_w18409_
	);
	LUT2 #(
		.INIT('h4)
	) name17878 (
		_w18317_,
		_w18409_,
		_w18410_
	);
	LUT2 #(
		.INIT('h2)
	) name17879 (
		\u0_w_reg[3][2]/P0001 ,
		_w16705_,
		_w18411_
	);
	LUT2 #(
		.INIT('h4)
	) name17880 (
		_w17958_,
		_w18411_,
		_w18412_
	);
	LUT2 #(
		.INIT('h8)
	) name17881 (
		_w18176_,
		_w18412_,
		_w18413_
	);
	LUT2 #(
		.INIT('h1)
	) name17882 (
		_w18410_,
		_w18413_,
		_w18414_
	);
	LUT2 #(
		.INIT('h1)
	) name17883 (
		_w16622_,
		_w18396_,
		_w18415_
	);
	LUT2 #(
		.INIT('h2)
	) name17884 (
		_w16689_,
		_w18415_,
		_w18416_
	);
	LUT2 #(
		.INIT('h1)
	) name17885 (
		_w16550_,
		_w18305_,
		_w18417_
	);
	LUT2 #(
		.INIT('h2)
	) name17886 (
		\u0_w_reg[3][4]/P0001 ,
		_w18417_,
		_w18418_
	);
	LUT2 #(
		.INIT('h1)
	) name17887 (
		\u0_w_reg[3][1]/P0001 ,
		_w16743_,
		_w18419_
	);
	LUT2 #(
		.INIT('h1)
	) name17888 (
		_w17505_,
		_w18175_,
		_w18420_
	);
	LUT2 #(
		.INIT('h8)
	) name17889 (
		_w18419_,
		_w18420_,
		_w18421_
	);
	LUT2 #(
		.INIT('h4)
	) name17890 (
		_w18416_,
		_w18421_,
		_w18422_
	);
	LUT2 #(
		.INIT('h4)
	) name17891 (
		_w18418_,
		_w18422_,
		_w18423_
	);
	LUT2 #(
		.INIT('h2)
	) name17892 (
		\u0_w_reg[3][1]/P0001 ,
		_w16587_,
		_w18424_
	);
	LUT2 #(
		.INIT('h4)
	) name17893 (
		_w17969_,
		_w18424_,
		_w18425_
	);
	LUT2 #(
		.INIT('h4)
	) name17894 (
		_w16573_,
		_w18425_,
		_w18426_
	);
	LUT2 #(
		.INIT('h1)
	) name17895 (
		_w18423_,
		_w18426_,
		_w18427_
	);
	LUT2 #(
		.INIT('h2)
	) name17896 (
		\u0_w_reg[3][0]/P0001 ,
		_w16484_,
		_w18428_
	);
	LUT2 #(
		.INIT('h4)
	) name17897 (
		_w16744_,
		_w18428_,
		_w18429_
	);
	LUT2 #(
		.INIT('h4)
	) name17898 (
		_w18414_,
		_w18429_,
		_w18430_
	);
	LUT2 #(
		.INIT('h4)
	) name17899 (
		_w18427_,
		_w18430_,
		_w18431_
	);
	LUT2 #(
		.INIT('h1)
	) name17900 (
		_w18407_,
		_w18431_,
		_w18432_
	);
	LUT2 #(
		.INIT('h1)
	) name17901 (
		_w18384_,
		_w18385_,
		_w18433_
	);
	LUT2 #(
		.INIT('h4)
	) name17902 (
		_w18432_,
		_w18433_,
		_w18434_
	);
	LUT2 #(
		.INIT('h2)
	) name17903 (
		\u0_w_reg[0][8]/P0001 ,
		_w18434_,
		_w18435_
	);
	LUT2 #(
		.INIT('h4)
	) name17904 (
		\u0_w_reg[0][8]/P0001 ,
		_w18434_,
		_w18436_
	);
	LUT2 #(
		.INIT('h1)
	) name17905 (
		_w18435_,
		_w18436_,
		_w18437_
	);
	LUT2 #(
		.INIT('h2)
	) name17906 (
		\u0_w_reg[1][8]/P0001 ,
		\u0_w_reg[2][8]/P0001 ,
		_w18438_
	);
	LUT2 #(
		.INIT('h4)
	) name17907 (
		\u0_w_reg[1][8]/P0001 ,
		\u0_w_reg[2][8]/P0001 ,
		_w18439_
	);
	LUT2 #(
		.INIT('h1)
	) name17908 (
		_w18438_,
		_w18439_,
		_w18440_
	);
	LUT2 #(
		.INIT('h8)
	) name17909 (
		_w18437_,
		_w18440_,
		_w18441_
	);
	LUT2 #(
		.INIT('h1)
	) name17910 (
		_w18437_,
		_w18440_,
		_w18442_
	);
	LUT2 #(
		.INIT('h1)
	) name17911 (
		_w18441_,
		_w18442_,
		_w18443_
	);
	LUT2 #(
		.INIT('h4)
	) name17912 (
		ld_pad,
		_w18443_,
		_w18444_
	);
	LUT2 #(
		.INIT('h1)
	) name17913 (
		_w18365_,
		_w18444_,
		_w18445_
	);
	LUT2 #(
		.INIT('h4)
	) name17914 (
		_w15588_,
		_w15592_,
		_w18446_
	);
	LUT2 #(
		.INIT('h8)
	) name17915 (
		\u0_w_reg[3][19]/P0001 ,
		_w15590_,
		_w18447_
	);
	LUT2 #(
		.INIT('h1)
	) name17916 (
		_w16840_,
		_w17110_,
		_w18448_
	);
	LUT2 #(
		.INIT('h4)
	) name17917 (
		_w18447_,
		_w18448_,
		_w18449_
	);
	LUT2 #(
		.INIT('h2)
	) name17918 (
		\u0_w_reg[3][18]/P0001 ,
		_w18449_,
		_w18450_
	);
	LUT2 #(
		.INIT('h2)
	) name17919 (
		_w16874_,
		_w18450_,
		_w18451_
	);
	LUT2 #(
		.INIT('h2)
	) name17920 (
		\u0_w_reg[3][17]/P0001 ,
		_w18451_,
		_w18452_
	);
	LUT2 #(
		.INIT('h8)
	) name17921 (
		_w15529_,
		_w15530_,
		_w18453_
	);
	LUT2 #(
		.INIT('h8)
	) name17922 (
		_w15560_,
		_w16268_,
		_w18454_
	);
	LUT2 #(
		.INIT('h1)
	) name17923 (
		_w15530_,
		_w15542_,
		_w18455_
	);
	LUT2 #(
		.INIT('h2)
	) name17924 (
		_w15521_,
		_w18455_,
		_w18456_
	);
	LUT2 #(
		.INIT('h1)
	) name17925 (
		_w18453_,
		_w18454_,
		_w18457_
	);
	LUT2 #(
		.INIT('h4)
	) name17926 (
		_w18456_,
		_w18457_,
		_w18458_
	);
	LUT2 #(
		.INIT('h1)
	) name17927 (
		\u0_w_reg[3][17]/P0001 ,
		_w18458_,
		_w18459_
	);
	LUT2 #(
		.INIT('h1)
	) name17928 (
		_w16814_,
		_w16944_,
		_w18460_
	);
	LUT2 #(
		.INIT('h1)
	) name17929 (
		\u0_w_reg[3][18]/P0001 ,
		_w18460_,
		_w18461_
	);
	LUT2 #(
		.INIT('h2)
	) name17930 (
		_w16283_,
		_w16901_,
		_w18462_
	);
	LUT2 #(
		.INIT('h4)
	) name17931 (
		_w15608_,
		_w15655_,
		_w18463_
	);
	LUT2 #(
		.INIT('h1)
	) name17932 (
		_w18446_,
		_w18463_,
		_w18464_
	);
	LUT2 #(
		.INIT('h4)
	) name17933 (
		_w18462_,
		_w18464_,
		_w18465_
	);
	LUT2 #(
		.INIT('h4)
	) name17934 (
		_w18461_,
		_w18465_,
		_w18466_
	);
	LUT2 #(
		.INIT('h4)
	) name17935 (
		_w18459_,
		_w18466_,
		_w18467_
	);
	LUT2 #(
		.INIT('h4)
	) name17936 (
		_w18452_,
		_w18467_,
		_w18468_
	);
	LUT2 #(
		.INIT('h2)
	) name17937 (
		\u0_w_reg[3][16]/P0001 ,
		_w18468_,
		_w18469_
	);
	LUT2 #(
		.INIT('h8)
	) name17938 (
		\u0_w_reg[3][19]/P0001 ,
		_w16840_,
		_w18470_
	);
	LUT2 #(
		.INIT('h1)
	) name17939 (
		_w15550_,
		_w16875_,
		_w18471_
	);
	LUT2 #(
		.INIT('h4)
	) name17940 (
		_w18470_,
		_w18471_,
		_w18472_
	);
	LUT2 #(
		.INIT('h1)
	) name17941 (
		\u0_w_reg[3][18]/P0001 ,
		_w18472_,
		_w18473_
	);
	LUT2 #(
		.INIT('h4)
	) name17942 (
		\u0_w_reg[3][19]/P0001 ,
		_w15606_,
		_w18474_
	);
	LUT2 #(
		.INIT('h1)
	) name17943 (
		_w15615_,
		_w18474_,
		_w18475_
	);
	LUT2 #(
		.INIT('h2)
	) name17944 (
		\u0_w_reg[3][18]/P0001 ,
		_w18475_,
		_w18476_
	);
	LUT2 #(
		.INIT('h2)
	) name17945 (
		\u0_w_reg[3][17]/P0001 ,
		_w15584_,
		_w18477_
	);
	LUT2 #(
		.INIT('h8)
	) name17946 (
		_w15541_,
		_w18477_,
		_w18478_
	);
	LUT2 #(
		.INIT('h4)
	) name17947 (
		_w18473_,
		_w18478_,
		_w18479_
	);
	LUT2 #(
		.INIT('h4)
	) name17948 (
		_w18476_,
		_w18479_,
		_w18480_
	);
	LUT2 #(
		.INIT('h4)
	) name17949 (
		\u0_w_reg[3][20]/P0001 ,
		_w16242_,
		_w18481_
	);
	LUT2 #(
		.INIT('h8)
	) name17950 (
		_w15660_,
		_w17090_,
		_w18482_
	);
	LUT2 #(
		.INIT('h1)
	) name17951 (
		\u0_w_reg[3][17]/P0001 ,
		_w16276_,
		_w18483_
	);
	LUT2 #(
		.INIT('h1)
	) name17952 (
		_w16288_,
		_w16909_,
		_w18484_
	);
	LUT2 #(
		.INIT('h1)
	) name17953 (
		_w17018_,
		_w18481_,
		_w18485_
	);
	LUT2 #(
		.INIT('h4)
	) name17954 (
		_w18482_,
		_w18485_,
		_w18486_
	);
	LUT2 #(
		.INIT('h8)
	) name17955 (
		_w18483_,
		_w18484_,
		_w18487_
	);
	LUT2 #(
		.INIT('h8)
	) name17956 (
		_w18486_,
		_w18487_,
		_w18488_
	);
	LUT2 #(
		.INIT('h1)
	) name17957 (
		_w18480_,
		_w18488_,
		_w18489_
	);
	LUT2 #(
		.INIT('h8)
	) name17958 (
		_w15529_,
		_w16313_,
		_w18490_
	);
	LUT2 #(
		.INIT('h1)
	) name17959 (
		_w15557_,
		_w15613_,
		_w18491_
	);
	LUT2 #(
		.INIT('h2)
	) name17960 (
		_w15511_,
		_w18491_,
		_w18492_
	);
	LUT2 #(
		.INIT('h1)
	) name17961 (
		_w15637_,
		_w15656_,
		_w18493_
	);
	LUT2 #(
		.INIT('h4)
	) name17962 (
		_w18490_,
		_w18493_,
		_w18494_
	);
	LUT2 #(
		.INIT('h1)
	) name17963 (
		_w16240_,
		_w18492_,
		_w18495_
	);
	LUT2 #(
		.INIT('h8)
	) name17964 (
		_w18494_,
		_w18495_,
		_w18496_
	);
	LUT2 #(
		.INIT('h4)
	) name17965 (
		_w18489_,
		_w18496_,
		_w18497_
	);
	LUT2 #(
		.INIT('h1)
	) name17966 (
		\u0_w_reg[3][16]/P0001 ,
		_w18497_,
		_w18498_
	);
	LUT2 #(
		.INIT('h1)
	) name17967 (
		_w15513_,
		_w15625_,
		_w18499_
	);
	LUT2 #(
		.INIT('h2)
	) name17968 (
		\u0_w_reg[3][19]/P0001 ,
		_w18499_,
		_w18500_
	);
	LUT2 #(
		.INIT('h1)
	) name17969 (
		_w17032_,
		_w18500_,
		_w18501_
	);
	LUT2 #(
		.INIT('h2)
	) name17970 (
		_w16901_,
		_w18501_,
		_w18502_
	);
	LUT2 #(
		.INIT('h1)
	) name17971 (
		_w15603_,
		_w15630_,
		_w18503_
	);
	LUT2 #(
		.INIT('h2)
	) name17972 (
		_w15608_,
		_w18503_,
		_w18504_
	);
	LUT2 #(
		.INIT('h1)
	) name17973 (
		_w15531_,
		_w15620_,
		_w18505_
	);
	LUT2 #(
		.INIT('h4)
	) name17974 (
		_w15514_,
		_w18505_,
		_w18506_
	);
	LUT2 #(
		.INIT('h2)
	) name17975 (
		_w16282_,
		_w18506_,
		_w18507_
	);
	LUT2 #(
		.INIT('h1)
	) name17976 (
		_w15560_,
		_w15630_,
		_w18508_
	);
	LUT2 #(
		.INIT('h1)
	) name17977 (
		_w15544_,
		_w18508_,
		_w18509_
	);
	LUT2 #(
		.INIT('h1)
	) name17978 (
		_w15584_,
		_w16851_,
		_w18510_
	);
	LUT2 #(
		.INIT('h4)
	) name17979 (
		_w18509_,
		_w18510_,
		_w18511_
	);
	LUT2 #(
		.INIT('h2)
	) name17980 (
		_w16910_,
		_w18511_,
		_w18512_
	);
	LUT2 #(
		.INIT('h1)
	) name17981 (
		_w15558_,
		_w17059_,
		_w18513_
	);
	LUT2 #(
		.INIT('h4)
	) name17982 (
		_w16802_,
		_w18513_,
		_w18514_
	);
	LUT2 #(
		.INIT('h1)
	) name17983 (
		\u0_w_reg[3][18]/P0001 ,
		_w18514_,
		_w18515_
	);
	LUT2 #(
		.INIT('h1)
	) name17984 (
		_w15563_,
		_w16222_,
		_w18516_
	);
	LUT2 #(
		.INIT('h4)
	) name17985 (
		_w18515_,
		_w18516_,
		_w18517_
	);
	LUT2 #(
		.INIT('h1)
	) name17986 (
		\u0_w_reg[3][17]/P0001 ,
		_w18517_,
		_w18518_
	);
	LUT2 #(
		.INIT('h1)
	) name17987 (
		_w18504_,
		_w18507_,
		_w18519_
	);
	LUT2 #(
		.INIT('h4)
	) name17988 (
		_w18502_,
		_w18519_,
		_w18520_
	);
	LUT2 #(
		.INIT('h4)
	) name17989 (
		_w18512_,
		_w18520_,
		_w18521_
	);
	LUT2 #(
		.INIT('h4)
	) name17990 (
		_w18518_,
		_w18521_,
		_w18522_
	);
	LUT2 #(
		.INIT('h4)
	) name17991 (
		_w18469_,
		_w18522_,
		_w18523_
	);
	LUT2 #(
		.INIT('h4)
	) name17992 (
		_w18498_,
		_w18523_,
		_w18524_
	);
	LUT2 #(
		.INIT('h2)
	) name17993 (
		\u0_w_reg[0][25]/P0001 ,
		_w18524_,
		_w18525_
	);
	LUT2 #(
		.INIT('h4)
	) name17994 (
		\u0_w_reg[0][25]/P0001 ,
		_w18524_,
		_w18526_
	);
	LUT2 #(
		.INIT('h1)
	) name17995 (
		_w18525_,
		_w18526_,
		_w18527_
	);
	LUT2 #(
		.INIT('h1)
	) name17996 (
		\u0_r0_out_reg[25]/P0001 ,
		_w18527_,
		_w18528_
	);
	LUT2 #(
		.INIT('h8)
	) name17997 (
		\u0_r0_out_reg[25]/P0001 ,
		_w18527_,
		_w18529_
	);
	LUT2 #(
		.INIT('h1)
	) name17998 (
		ld_pad,
		_w18528_,
		_w18530_
	);
	LUT2 #(
		.INIT('h4)
	) name17999 (
		_w18529_,
		_w18530_,
		_w18531_
	);
	LUT2 #(
		.INIT('h8)
	) name18000 (
		\key[121]_pad ,
		ld_pad,
		_w18532_
	);
	LUT2 #(
		.INIT('h1)
	) name18001 (
		_w18531_,
		_w18532_,
		_w18533_
	);
	LUT2 #(
		.INIT('h2)
	) name18002 (
		\u0_r0_out_reg[25]/P0001 ,
		\u0_w_reg[1][25]/P0001 ,
		_w18534_
	);
	LUT2 #(
		.INIT('h4)
	) name18003 (
		\u0_r0_out_reg[25]/P0001 ,
		\u0_w_reg[1][25]/P0001 ,
		_w18535_
	);
	LUT2 #(
		.INIT('h1)
	) name18004 (
		_w18534_,
		_w18535_,
		_w18536_
	);
	LUT2 #(
		.INIT('h4)
	) name18005 (
		_w18527_,
		_w18536_,
		_w18537_
	);
	LUT2 #(
		.INIT('h2)
	) name18006 (
		_w18527_,
		_w18536_,
		_w18538_
	);
	LUT2 #(
		.INIT('h1)
	) name18007 (
		ld_pad,
		_w18537_,
		_w18539_
	);
	LUT2 #(
		.INIT('h4)
	) name18008 (
		_w18538_,
		_w18539_,
		_w18540_
	);
	LUT2 #(
		.INIT('h8)
	) name18009 (
		\key[89]_pad ,
		ld_pad,
		_w18541_
	);
	LUT2 #(
		.INIT('h1)
	) name18010 (
		_w18540_,
		_w18541_,
		_w18542_
	);
	LUT2 #(
		.INIT('h4)
	) name18011 (
		\key[57]_pad ,
		ld_pad,
		_w18543_
	);
	LUT2 #(
		.INIT('h8)
	) name18012 (
		\u0_w_reg[2][25]/P0001 ,
		_w18536_,
		_w18544_
	);
	LUT2 #(
		.INIT('h1)
	) name18013 (
		\u0_w_reg[2][25]/P0001 ,
		_w18536_,
		_w18545_
	);
	LUT2 #(
		.INIT('h1)
	) name18014 (
		_w18544_,
		_w18545_,
		_w18546_
	);
	LUT2 #(
		.INIT('h8)
	) name18015 (
		_w18527_,
		_w18546_,
		_w18547_
	);
	LUT2 #(
		.INIT('h1)
	) name18016 (
		_w18527_,
		_w18546_,
		_w18548_
	);
	LUT2 #(
		.INIT('h1)
	) name18017 (
		_w18547_,
		_w18548_,
		_w18549_
	);
	LUT2 #(
		.INIT('h4)
	) name18018 (
		ld_pad,
		_w18549_,
		_w18550_
	);
	LUT2 #(
		.INIT('h1)
	) name18019 (
		_w18543_,
		_w18550_,
		_w18551_
	);
	LUT2 #(
		.INIT('h4)
	) name18020 (
		\u0_w_reg[3][25]/P0001 ,
		_w18549_,
		_w18552_
	);
	LUT2 #(
		.INIT('h2)
	) name18021 (
		\u0_w_reg[3][25]/P0001 ,
		_w18549_,
		_w18553_
	);
	LUT2 #(
		.INIT('h1)
	) name18022 (
		ld_pad,
		_w18552_,
		_w18554_
	);
	LUT2 #(
		.INIT('h4)
	) name18023 (
		_w18553_,
		_w18554_,
		_w18555_
	);
	LUT2 #(
		.INIT('h8)
	) name18024 (
		\key[25]_pad ,
		ld_pad,
		_w18556_
	);
	LUT2 #(
		.INIT('h1)
	) name18025 (
		_w18555_,
		_w18556_,
		_w18557_
	);
	LUT2 #(
		.INIT('h4)
	) name18026 (
		\u0_w_reg[3][15]/P0001 ,
		_w17644_,
		_w18558_
	);
	LUT2 #(
		.INIT('h1)
	) name18027 (
		_w15754_,
		_w18558_,
		_w18559_
	);
	LUT2 #(
		.INIT('h1)
	) name18028 (
		\u0_w_reg[3][10]/P0001 ,
		_w18559_,
		_w18560_
	);
	LUT2 #(
		.INIT('h1)
	) name18029 (
		_w17684_,
		_w17771_,
		_w18561_
	);
	LUT2 #(
		.INIT('h4)
	) name18030 (
		_w18017_,
		_w18561_,
		_w18562_
	);
	LUT2 #(
		.INIT('h4)
	) name18031 (
		_w18560_,
		_w18562_,
		_w18563_
	);
	LUT2 #(
		.INIT('h2)
	) name18032 (
		\u0_w_reg[3][9]/P0001 ,
		_w18563_,
		_w18564_
	);
	LUT2 #(
		.INIT('h8)
	) name18033 (
		_w15799_,
		_w15946_,
		_w18565_
	);
	LUT2 #(
		.INIT('h1)
	) name18034 (
		_w15804_,
		_w17638_,
		_w18566_
	);
	LUT2 #(
		.INIT('h4)
	) name18035 (
		_w18565_,
		_w18566_,
		_w18567_
	);
	LUT2 #(
		.INIT('h1)
	) name18036 (
		\u0_w_reg[3][9]/P0001 ,
		_w18567_,
		_w18568_
	);
	LUT2 #(
		.INIT('h1)
	) name18037 (
		_w15758_,
		_w17722_,
		_w18569_
	);
	LUT2 #(
		.INIT('h1)
	) name18038 (
		\u0_w_reg[3][10]/P0001 ,
		_w18569_,
		_w18570_
	);
	LUT2 #(
		.INIT('h8)
	) name18039 (
		\u0_w_reg[3][10]/P0001 ,
		_w17731_,
		_w18571_
	);
	LUT2 #(
		.INIT('h4)
	) name18040 (
		_w15757_,
		_w15847_,
		_w18572_
	);
	LUT2 #(
		.INIT('h8)
	) name18041 (
		_w17631_,
		_w18572_,
		_w18573_
	);
	LUT2 #(
		.INIT('h8)
	) name18042 (
		_w15803_,
		_w15865_,
		_w18574_
	);
	LUT2 #(
		.INIT('h1)
	) name18043 (
		\u0_w_reg[3][8]/P0001 ,
		_w15980_,
		_w18575_
	);
	LUT2 #(
		.INIT('h4)
	) name18044 (
		_w15861_,
		_w18575_,
		_w18576_
	);
	LUT2 #(
		.INIT('h1)
	) name18045 (
		_w18573_,
		_w18574_,
		_w18577_
	);
	LUT2 #(
		.INIT('h8)
	) name18046 (
		_w18576_,
		_w18577_,
		_w18578_
	);
	LUT2 #(
		.INIT('h4)
	) name18047 (
		_w18571_,
		_w18578_,
		_w18579_
	);
	LUT2 #(
		.INIT('h1)
	) name18048 (
		_w18568_,
		_w18570_,
		_w18580_
	);
	LUT2 #(
		.INIT('h8)
	) name18049 (
		_w18579_,
		_w18580_,
		_w18581_
	);
	LUT2 #(
		.INIT('h4)
	) name18050 (
		_w18564_,
		_w18581_,
		_w18582_
	);
	LUT2 #(
		.INIT('h4)
	) name18051 (
		_w15787_,
		_w17651_,
		_w18583_
	);
	LUT2 #(
		.INIT('h1)
	) name18052 (
		_w15942_,
		_w18583_,
		_w18584_
	);
	LUT2 #(
		.INIT('h2)
	) name18053 (
		\u0_w_reg[3][12]/P0001 ,
		_w18584_,
		_w18585_
	);
	LUT2 #(
		.INIT('h4)
	) name18054 (
		\u0_w_reg[3][10]/P0001 ,
		_w15741_,
		_w18586_
	);
	LUT2 #(
		.INIT('h8)
	) name18055 (
		_w15803_,
		_w15896_,
		_w18587_
	);
	LUT2 #(
		.INIT('h8)
	) name18056 (
		_w15725_,
		_w15847_,
		_w18588_
	);
	LUT2 #(
		.INIT('h1)
	) name18057 (
		\u0_w_reg[3][9]/P0001 ,
		_w17682_,
		_w18589_
	);
	LUT2 #(
		.INIT('h4)
	) name18058 (
		_w18588_,
		_w18589_,
		_w18590_
	);
	LUT2 #(
		.INIT('h1)
	) name18059 (
		_w18586_,
		_w18587_,
		_w18591_
	);
	LUT2 #(
		.INIT('h8)
	) name18060 (
		_w18590_,
		_w18591_,
		_w18592_
	);
	LUT2 #(
		.INIT('h4)
	) name18061 (
		_w18585_,
		_w18592_,
		_w18593_
	);
	LUT2 #(
		.INIT('h8)
	) name18062 (
		\u0_w_reg[3][11]/P0001 ,
		_w15725_,
		_w18594_
	);
	LUT2 #(
		.INIT('h1)
	) name18063 (
		_w15716_,
		_w15983_,
		_w18595_
	);
	LUT2 #(
		.INIT('h1)
	) name18064 (
		_w17609_,
		_w18594_,
		_w18596_
	);
	LUT2 #(
		.INIT('h8)
	) name18065 (
		_w18595_,
		_w18596_,
		_w18597_
	);
	LUT2 #(
		.INIT('h2)
	) name18066 (
		\u0_w_reg[3][10]/P0001 ,
		_w18597_,
		_w18598_
	);
	LUT2 #(
		.INIT('h2)
	) name18067 (
		\u0_w_reg[3][9]/P0001 ,
		_w17781_,
		_w18599_
	);
	LUT2 #(
		.INIT('h4)
	) name18068 (
		\u0_w_reg[3][14]/P0001 ,
		_w17610_,
		_w18600_
	);
	LUT2 #(
		.INIT('h2)
	) name18069 (
		_w18599_,
		_w18600_,
		_w18601_
	);
	LUT2 #(
		.INIT('h4)
	) name18070 (
		_w18598_,
		_w18601_,
		_w18602_
	);
	LUT2 #(
		.INIT('h1)
	) name18071 (
		_w18593_,
		_w18602_,
		_w18603_
	);
	LUT2 #(
		.INIT('h8)
	) name18072 (
		\u0_w_reg[3][12]/P0001 ,
		_w18588_,
		_w18604_
	);
	LUT2 #(
		.INIT('h8)
	) name18073 (
		\u0_w_reg[3][15]/P0001 ,
		_w15716_,
		_w18605_
	);
	LUT2 #(
		.INIT('h1)
	) name18074 (
		_w17737_,
		_w18605_,
		_w18606_
	);
	LUT2 #(
		.INIT('h2)
	) name18075 (
		_w15893_,
		_w18606_,
		_w18607_
	);
	LUT2 #(
		.INIT('h8)
	) name18076 (
		_w15738_,
		_w15799_,
		_w18608_
	);
	LUT2 #(
		.INIT('h2)
	) name18077 (
		\u0_w_reg[3][8]/P0001 ,
		_w17643_,
		_w18609_
	);
	LUT2 #(
		.INIT('h4)
	) name18078 (
		_w15792_,
		_w18609_,
		_w18610_
	);
	LUT2 #(
		.INIT('h1)
	) name18079 (
		_w18604_,
		_w18608_,
		_w18611_
	);
	LUT2 #(
		.INIT('h8)
	) name18080 (
		_w18610_,
		_w18611_,
		_w18612_
	);
	LUT2 #(
		.INIT('h4)
	) name18081 (
		_w18607_,
		_w18612_,
		_w18613_
	);
	LUT2 #(
		.INIT('h4)
	) name18082 (
		_w18603_,
		_w18613_,
		_w18614_
	);
	LUT2 #(
		.INIT('h1)
	) name18083 (
		_w18582_,
		_w18614_,
		_w18615_
	);
	LUT2 #(
		.INIT('h4)
	) name18084 (
		_w17598_,
		_w17601_,
		_w18616_
	);
	LUT2 #(
		.INIT('h2)
	) name18085 (
		\u0_w_reg[3][11]/P0001 ,
		_w18616_,
		_w18617_
	);
	LUT2 #(
		.INIT('h1)
	) name18086 (
		\u0_w_reg[3][10]/P0001 ,
		_w15837_,
		_w18618_
	);
	LUT2 #(
		.INIT('h4)
	) name18087 (
		_w18617_,
		_w18618_,
		_w18619_
	);
	LUT2 #(
		.INIT('h1)
	) name18088 (
		_w15802_,
		_w17672_,
		_w18620_
	);
	LUT2 #(
		.INIT('h4)
	) name18089 (
		_w18605_,
		_w18620_,
		_w18621_
	);
	LUT2 #(
		.INIT('h1)
	) name18090 (
		\u0_w_reg[3][11]/P0001 ,
		_w18621_,
		_w18622_
	);
	LUT2 #(
		.INIT('h2)
	) name18091 (
		\u0_w_reg[3][10]/P0001 ,
		_w15715_,
		_w18623_
	);
	LUT2 #(
		.INIT('h4)
	) name18092 (
		_w15815_,
		_w18623_,
		_w18624_
	);
	LUT2 #(
		.INIT('h4)
	) name18093 (
		_w18622_,
		_w18624_,
		_w18625_
	);
	LUT2 #(
		.INIT('h2)
	) name18094 (
		\u0_w_reg[3][9]/P0001 ,
		_w18619_,
		_w18626_
	);
	LUT2 #(
		.INIT('h4)
	) name18095 (
		_w18625_,
		_w18626_,
		_w18627_
	);
	LUT2 #(
		.INIT('h8)
	) name18096 (
		_w15735_,
		_w15943_,
		_w18628_
	);
	LUT2 #(
		.INIT('h1)
	) name18097 (
		_w15785_,
		_w18628_,
		_w18629_
	);
	LUT2 #(
		.INIT('h1)
	) name18098 (
		\u0_w_reg[3][10]/P0001 ,
		_w18629_,
		_w18630_
	);
	LUT2 #(
		.INIT('h1)
	) name18099 (
		_w15789_,
		_w15902_,
		_w18631_
	);
	LUT2 #(
		.INIT('h4)
	) name18100 (
		_w17781_,
		_w18631_,
		_w18632_
	);
	LUT2 #(
		.INIT('h2)
	) name18101 (
		_w15974_,
		_w18632_,
		_w18633_
	);
	LUT2 #(
		.INIT('h4)
	) name18102 (
		\u0_w_reg[3][12]/P0001 ,
		_w15814_,
		_w18634_
	);
	LUT2 #(
		.INIT('h8)
	) name18103 (
		_w15849_,
		_w18634_,
		_w18635_
	);
	LUT2 #(
		.INIT('h1)
	) name18104 (
		_w15941_,
		_w18573_,
		_w18636_
	);
	LUT2 #(
		.INIT('h4)
	) name18105 (
		_w18635_,
		_w18636_,
		_w18637_
	);
	LUT2 #(
		.INIT('h1)
	) name18106 (
		\u0_w_reg[3][9]/P0001 ,
		_w18637_,
		_w18638_
	);
	LUT2 #(
		.INIT('h1)
	) name18107 (
		_w18630_,
		_w18633_,
		_w18639_
	);
	LUT2 #(
		.INIT('h4)
	) name18108 (
		_w18638_,
		_w18639_,
		_w18640_
	);
	LUT2 #(
		.INIT('h4)
	) name18109 (
		_w18627_,
		_w18640_,
		_w18641_
	);
	LUT2 #(
		.INIT('h4)
	) name18110 (
		_w18615_,
		_w18641_,
		_w18642_
	);
	LUT2 #(
		.INIT('h2)
	) name18111 (
		\u0_w_reg[0][23]/P0001 ,
		_w18642_,
		_w18643_
	);
	LUT2 #(
		.INIT('h4)
	) name18112 (
		\u0_w_reg[0][23]/P0001 ,
		_w18642_,
		_w18644_
	);
	LUT2 #(
		.INIT('h1)
	) name18113 (
		_w18643_,
		_w18644_,
		_w18645_
	);
	LUT2 #(
		.INIT('h8)
	) name18114 (
		\u0_w_reg[1][23]/P0001 ,
		_w18645_,
		_w18646_
	);
	LUT2 #(
		.INIT('h1)
	) name18115 (
		\u0_w_reg[1][23]/P0001 ,
		_w18645_,
		_w18647_
	);
	LUT2 #(
		.INIT('h1)
	) name18116 (
		_w18646_,
		_w18647_,
		_w18648_
	);
	LUT2 #(
		.INIT('h8)
	) name18117 (
		\u0_w_reg[2][23]/P0001 ,
		_w18648_,
		_w18649_
	);
	LUT2 #(
		.INIT('h1)
	) name18118 (
		\u0_w_reg[2][23]/P0001 ,
		_w18648_,
		_w18650_
	);
	LUT2 #(
		.INIT('h1)
	) name18119 (
		_w18649_,
		_w18650_,
		_w18651_
	);
	LUT2 #(
		.INIT('h4)
	) name18120 (
		ld_pad,
		_w18651_,
		_w18652_
	);
	LUT2 #(
		.INIT('h8)
	) name18121 (
		\key[55]_pad ,
		ld_pad,
		_w18653_
	);
	LUT2 #(
		.INIT('h1)
	) name18122 (
		_w18652_,
		_w18653_,
		_w18654_
	);
	LUT2 #(
		.INIT('h4)
	) name18123 (
		ld_pad,
		_w16466_,
		_w18655_
	);
	LUT2 #(
		.INIT('h8)
	) name18124 (
		\key[99]_pad ,
		ld_pad,
		_w18656_
	);
	LUT2 #(
		.INIT('h1)
	) name18125 (
		_w18655_,
		_w18656_,
		_w18657_
	);
	LUT2 #(
		.INIT('h1)
	) name18126 (
		\u0_w_reg[1][3]/P0001 ,
		_w16466_,
		_w18658_
	);
	LUT2 #(
		.INIT('h8)
	) name18127 (
		\u0_w_reg[1][3]/P0001 ,
		_w16466_,
		_w18659_
	);
	LUT2 #(
		.INIT('h1)
	) name18128 (
		ld_pad,
		_w18658_,
		_w18660_
	);
	LUT2 #(
		.INIT('h4)
	) name18129 (
		_w18659_,
		_w18660_,
		_w18661_
	);
	LUT2 #(
		.INIT('h8)
	) name18130 (
		\key[67]_pad ,
		ld_pad,
		_w18662_
	);
	LUT2 #(
		.INIT('h1)
	) name18131 (
		_w18661_,
		_w18662_,
		_w18663_
	);
	LUT2 #(
		.INIT('h4)
	) name18132 (
		\u0_w_reg[3][3]/P0001 ,
		_w16472_,
		_w18664_
	);
	LUT2 #(
		.INIT('h2)
	) name18133 (
		\u0_w_reg[3][3]/P0001 ,
		_w16472_,
		_w18665_
	);
	LUT2 #(
		.INIT('h1)
	) name18134 (
		ld_pad,
		_w18664_,
		_w18666_
	);
	LUT2 #(
		.INIT('h4)
	) name18135 (
		_w18665_,
		_w18666_,
		_w18667_
	);
	LUT2 #(
		.INIT('h8)
	) name18136 (
		\key[3]_pad ,
		ld_pad,
		_w18668_
	);
	LUT2 #(
		.INIT('h1)
	) name18137 (
		_w18667_,
		_w18668_,
		_w18669_
	);
	LUT2 #(
		.INIT('h4)
	) name18138 (
		ld_pad,
		_w16639_,
		_w18670_
	);
	LUT2 #(
		.INIT('h8)
	) name18139 (
		\key[107]_pad ,
		ld_pad,
		_w18671_
	);
	LUT2 #(
		.INIT('h1)
	) name18140 (
		_w18670_,
		_w18671_,
		_w18672_
	);
	LUT2 #(
		.INIT('h1)
	) name18141 (
		\u0_w_reg[1][11]/P0001 ,
		_w16639_,
		_w18673_
	);
	LUT2 #(
		.INIT('h8)
	) name18142 (
		\u0_w_reg[1][11]/P0001 ,
		_w16639_,
		_w18674_
	);
	LUT2 #(
		.INIT('h1)
	) name18143 (
		ld_pad,
		_w18673_,
		_w18675_
	);
	LUT2 #(
		.INIT('h4)
	) name18144 (
		_w18674_,
		_w18675_,
		_w18676_
	);
	LUT2 #(
		.INIT('h8)
	) name18145 (
		\key[75]_pad ,
		ld_pad,
		_w18677_
	);
	LUT2 #(
		.INIT('h1)
	) name18146 (
		_w18676_,
		_w18677_,
		_w18678_
	);
	LUT2 #(
		.INIT('h4)
	) name18147 (
		\u0_w_reg[3][11]/P0001 ,
		_w16645_,
		_w18679_
	);
	LUT2 #(
		.INIT('h2)
	) name18148 (
		\u0_w_reg[3][11]/P0001 ,
		_w16645_,
		_w18680_
	);
	LUT2 #(
		.INIT('h1)
	) name18149 (
		ld_pad,
		_w18679_,
		_w18681_
	);
	LUT2 #(
		.INIT('h4)
	) name18150 (
		_w18680_,
		_w18681_,
		_w18682_
	);
	LUT2 #(
		.INIT('h8)
	) name18151 (
		\key[11]_pad ,
		ld_pad,
		_w18683_
	);
	LUT2 #(
		.INIT('h1)
	) name18152 (
		_w18682_,
		_w18683_,
		_w18684_
	);
	LUT2 #(
		.INIT('h4)
	) name18153 (
		\key[49]_pad ,
		ld_pad,
		_w18685_
	);
	LUT2 #(
		.INIT('h2)
	) name18154 (
		_w15732_,
		_w17759_,
		_w18686_
	);
	LUT2 #(
		.INIT('h4)
	) name18155 (
		\u0_w_reg[3][11]/P0001 ,
		_w15742_,
		_w18687_
	);
	LUT2 #(
		.INIT('h1)
	) name18156 (
		\u0_w_reg[3][10]/P0001 ,
		_w18687_,
		_w18688_
	);
	LUT2 #(
		.INIT('h4)
	) name18157 (
		_w18686_,
		_w18688_,
		_w18689_
	);
	LUT2 #(
		.INIT('h4)
	) name18158 (
		\u0_w_reg[3][11]/P0001 ,
		_w15840_,
		_w18690_
	);
	LUT2 #(
		.INIT('h2)
	) name18159 (
		\u0_w_reg[3][10]/P0001 ,
		_w15821_,
		_w18691_
	);
	LUT2 #(
		.INIT('h4)
	) name18160 (
		_w18690_,
		_w18691_,
		_w18692_
	);
	LUT2 #(
		.INIT('h1)
	) name18161 (
		_w18689_,
		_w18692_,
		_w18693_
	);
	LUT2 #(
		.INIT('h8)
	) name18162 (
		_w15718_,
		_w15790_,
		_w18694_
	);
	LUT2 #(
		.INIT('h4)
	) name18163 (
		_w18693_,
		_w18694_,
		_w18695_
	);
	LUT2 #(
		.INIT('h1)
	) name18164 (
		_w15812_,
		_w15846_,
		_w18696_
	);
	LUT2 #(
		.INIT('h2)
	) name18165 (
		_w15919_,
		_w18696_,
		_w18697_
	);
	LUT2 #(
		.INIT('h1)
	) name18166 (
		_w15757_,
		_w15896_,
		_w18698_
	);
	LUT2 #(
		.INIT('h2)
	) name18167 (
		_w15730_,
		_w18698_,
		_w18699_
	);
	LUT2 #(
		.INIT('h8)
	) name18168 (
		_w15787_,
		_w15799_,
		_w18700_
	);
	LUT2 #(
		.INIT('h1)
	) name18169 (
		\u0_w_reg[3][9]/P0001 ,
		_w18700_,
		_w18701_
	);
	LUT2 #(
		.INIT('h4)
	) name18170 (
		_w17757_,
		_w18701_,
		_w18702_
	);
	LUT2 #(
		.INIT('h1)
	) name18171 (
		_w18697_,
		_w18699_,
		_w18703_
	);
	LUT2 #(
		.INIT('h8)
	) name18172 (
		_w18702_,
		_w18703_,
		_w18704_
	);
	LUT2 #(
		.INIT('h1)
	) name18173 (
		_w18695_,
		_w18704_,
		_w18705_
	);
	LUT2 #(
		.INIT('h1)
	) name18174 (
		_w15822_,
		_w15943_,
		_w18706_
	);
	LUT2 #(
		.INIT('h2)
	) name18175 (
		_w15893_,
		_w18706_,
		_w18707_
	);
	LUT2 #(
		.INIT('h8)
	) name18176 (
		_w15805_,
		_w15849_,
		_w18708_
	);
	LUT2 #(
		.INIT('h1)
	) name18177 (
		_w15853_,
		_w15861_,
		_w18709_
	);
	LUT2 #(
		.INIT('h4)
	) name18178 (
		_w18708_,
		_w18709_,
		_w18710_
	);
	LUT2 #(
		.INIT('h1)
	) name18179 (
		_w15959_,
		_w18707_,
		_w18711_
	);
	LUT2 #(
		.INIT('h8)
	) name18180 (
		_w18710_,
		_w18711_,
		_w18712_
	);
	LUT2 #(
		.INIT('h4)
	) name18181 (
		_w18705_,
		_w18712_,
		_w18713_
	);
	LUT2 #(
		.INIT('h1)
	) name18182 (
		\u0_w_reg[3][8]/P0001 ,
		_w18713_,
		_w18714_
	);
	LUT2 #(
		.INIT('h1)
	) name18183 (
		_w15865_,
		_w15960_,
		_w18715_
	);
	LUT2 #(
		.INIT('h2)
	) name18184 (
		_w15803_,
		_w18715_,
		_w18716_
	);
	LUT2 #(
		.INIT('h1)
	) name18185 (
		_w15820_,
		_w15839_,
		_w18717_
	);
	LUT2 #(
		.INIT('h4)
	) name18186 (
		_w15705_,
		_w18717_,
		_w18718_
	);
	LUT2 #(
		.INIT('h2)
	) name18187 (
		_w15975_,
		_w18718_,
		_w18719_
	);
	LUT2 #(
		.INIT('h1)
	) name18188 (
		_w15823_,
		_w15929_,
		_w18720_
	);
	LUT2 #(
		.INIT('h1)
	) name18189 (
		\u0_w_reg[3][14]/P0001 ,
		_w18720_,
		_w18721_
	);
	LUT2 #(
		.INIT('h1)
	) name18190 (
		_w15789_,
		_w17667_,
		_w18722_
	);
	LUT2 #(
		.INIT('h4)
	) name18191 (
		_w17719_,
		_w18722_,
		_w18723_
	);
	LUT2 #(
		.INIT('h4)
	) name18192 (
		_w18721_,
		_w18723_,
		_w18724_
	);
	LUT2 #(
		.INIT('h2)
	) name18193 (
		_w15726_,
		_w18724_,
		_w18725_
	);
	LUT2 #(
		.INIT('h1)
	) name18194 (
		_w15971_,
		_w17721_,
		_w18726_
	);
	LUT2 #(
		.INIT('h4)
	) name18195 (
		_w18017_,
		_w18726_,
		_w18727_
	);
	LUT2 #(
		.INIT('h2)
	) name18196 (
		_w18055_,
		_w18727_,
		_w18728_
	);
	LUT2 #(
		.INIT('h1)
	) name18197 (
		_w15759_,
		_w17638_,
		_w18729_
	);
	LUT2 #(
		.INIT('h4)
	) name18198 (
		_w18558_,
		_w18729_,
		_w18730_
	);
	LUT2 #(
		.INIT('h1)
	) name18199 (
		\u0_w_reg[3][10]/P0001 ,
		_w18730_,
		_w18731_
	);
	LUT2 #(
		.INIT('h1)
	) name18200 (
		_w15755_,
		_w15932_,
		_w18732_
	);
	LUT2 #(
		.INIT('h4)
	) name18201 (
		_w18731_,
		_w18732_,
		_w18733_
	);
	LUT2 #(
		.INIT('h1)
	) name18202 (
		\u0_w_reg[3][9]/P0001 ,
		_w18733_,
		_w18734_
	);
	LUT2 #(
		.INIT('h1)
	) name18203 (
		_w17683_,
		_w17772_,
		_w18735_
	);
	LUT2 #(
		.INIT('h4)
	) name18204 (
		_w18634_,
		_w18735_,
		_w18736_
	);
	LUT2 #(
		.INIT('h2)
	) name18205 (
		\u0_w_reg[3][10]/P0001 ,
		_w18736_,
		_w18737_
	);
	LUT2 #(
		.INIT('h2)
	) name18206 (
		_w17732_,
		_w18737_,
		_w18738_
	);
	LUT2 #(
		.INIT('h2)
	) name18207 (
		\u0_w_reg[3][9]/P0001 ,
		_w18738_,
		_w18739_
	);
	LUT2 #(
		.INIT('h1)
	) name18208 (
		_w15742_,
		_w15859_,
		_w18740_
	);
	LUT2 #(
		.INIT('h1)
	) name18209 (
		_w15735_,
		_w15849_,
		_w18741_
	);
	LUT2 #(
		.INIT('h4)
	) name18210 (
		_w15929_,
		_w18741_,
		_w18742_
	);
	LUT2 #(
		.INIT('h1)
	) name18211 (
		_w18740_,
		_w18742_,
		_w18743_
	);
	LUT2 #(
		.INIT('h1)
	) name18212 (
		_w15976_,
		_w18743_,
		_w18744_
	);
	LUT2 #(
		.INIT('h1)
	) name18213 (
		\u0_w_reg[3][9]/P0001 ,
		_w18744_,
		_w18745_
	);
	LUT2 #(
		.INIT('h4)
	) name18214 (
		_w15782_,
		_w15787_,
		_w18746_
	);
	LUT2 #(
		.INIT('h1)
	) name18215 (
		_w17738_,
		_w18746_,
		_w18747_
	);
	LUT2 #(
		.INIT('h1)
	) name18216 (
		\u0_w_reg[3][11]/P0001 ,
		_w18747_,
		_w18748_
	);
	LUT2 #(
		.INIT('h1)
	) name18217 (
		_w15784_,
		_w15976_,
		_w18749_
	);
	LUT2 #(
		.INIT('h1)
	) name18218 (
		_w17738_,
		_w17771_,
		_w18750_
	);
	LUT2 #(
		.INIT('h8)
	) name18219 (
		_w18749_,
		_w18750_,
		_w18751_
	);
	LUT2 #(
		.INIT('h1)
	) name18220 (
		\u0_w_reg[3][10]/P0001 ,
		_w18751_,
		_w18752_
	);
	LUT2 #(
		.INIT('h1)
	) name18221 (
		_w18745_,
		_w18748_,
		_w18753_
	);
	LUT2 #(
		.INIT('h4)
	) name18222 (
		_w18752_,
		_w18753_,
		_w18754_
	);
	LUT2 #(
		.INIT('h4)
	) name18223 (
		_w18739_,
		_w18754_,
		_w18755_
	);
	LUT2 #(
		.INIT('h2)
	) name18224 (
		\u0_w_reg[3][8]/P0001 ,
		_w18755_,
		_w18756_
	);
	LUT2 #(
		.INIT('h1)
	) name18225 (
		_w18716_,
		_w18719_,
		_w18757_
	);
	LUT2 #(
		.INIT('h4)
	) name18226 (
		_w18725_,
		_w18757_,
		_w18758_
	);
	LUT2 #(
		.INIT('h4)
	) name18227 (
		_w18728_,
		_w18758_,
		_w18759_
	);
	LUT2 #(
		.INIT('h4)
	) name18228 (
		_w18734_,
		_w18759_,
		_w18760_
	);
	LUT2 #(
		.INIT('h4)
	) name18229 (
		_w18714_,
		_w18760_,
		_w18761_
	);
	LUT2 #(
		.INIT('h4)
	) name18230 (
		_w18756_,
		_w18761_,
		_w18762_
	);
	LUT2 #(
		.INIT('h2)
	) name18231 (
		\u0_w_reg[0][17]/P0001 ,
		_w18762_,
		_w18763_
	);
	LUT2 #(
		.INIT('h4)
	) name18232 (
		\u0_w_reg[0][17]/P0001 ,
		_w18762_,
		_w18764_
	);
	LUT2 #(
		.INIT('h1)
	) name18233 (
		_w18763_,
		_w18764_,
		_w18765_
	);
	LUT2 #(
		.INIT('h2)
	) name18234 (
		\u0_w_reg[1][17]/P0001 ,
		\u0_w_reg[2][17]/P0001 ,
		_w18766_
	);
	LUT2 #(
		.INIT('h4)
	) name18235 (
		\u0_w_reg[1][17]/P0001 ,
		\u0_w_reg[2][17]/P0001 ,
		_w18767_
	);
	LUT2 #(
		.INIT('h1)
	) name18236 (
		_w18766_,
		_w18767_,
		_w18768_
	);
	LUT2 #(
		.INIT('h8)
	) name18237 (
		_w18765_,
		_w18768_,
		_w18769_
	);
	LUT2 #(
		.INIT('h1)
	) name18238 (
		_w18765_,
		_w18768_,
		_w18770_
	);
	LUT2 #(
		.INIT('h1)
	) name18239 (
		_w18769_,
		_w18770_,
		_w18771_
	);
	LUT2 #(
		.INIT('h4)
	) name18240 (
		ld_pad,
		_w18771_,
		_w18772_
	);
	LUT2 #(
		.INIT('h1)
	) name18241 (
		_w18685_,
		_w18772_,
		_w18773_
	);
	LUT2 #(
		.INIT('h4)
	) name18242 (
		\key[33]_pad ,
		ld_pad,
		_w18774_
	);
	LUT2 #(
		.INIT('h1)
	) name18243 (
		_w16160_,
		_w17277_,
		_w18775_
	);
	LUT2 #(
		.INIT('h4)
	) name18244 (
		_w17835_,
		_w18775_,
		_w18776_
	);
	LUT2 #(
		.INIT('h2)
	) name18245 (
		\u0_w_reg[3][26]/P0001 ,
		_w18776_,
		_w18777_
	);
	LUT2 #(
		.INIT('h2)
	) name18246 (
		_w17853_,
		_w18777_,
		_w18778_
	);
	LUT2 #(
		.INIT('h2)
	) name18247 (
		\u0_w_reg[3][25]/P0001 ,
		_w18778_,
		_w18779_
	);
	LUT2 #(
		.INIT('h1)
	) name18248 (
		_w16043_,
		_w16102_,
		_w18780_
	);
	LUT2 #(
		.INIT('h1)
	) name18249 (
		_w16045_,
		_w16117_,
		_w18781_
	);
	LUT2 #(
		.INIT('h4)
	) name18250 (
		_w16112_,
		_w18781_,
		_w18782_
	);
	LUT2 #(
		.INIT('h1)
	) name18251 (
		_w18780_,
		_w18782_,
		_w18783_
	);
	LUT2 #(
		.INIT('h1)
	) name18252 (
		_w16040_,
		_w18783_,
		_w18784_
	);
	LUT2 #(
		.INIT('h1)
	) name18253 (
		\u0_w_reg[3][25]/P0001 ,
		_w18784_,
		_w18785_
	);
	LUT2 #(
		.INIT('h2)
	) name18254 (
		_w16099_,
		_w16147_,
		_w18786_
	);
	LUT2 #(
		.INIT('h1)
	) name18255 (
		_w17820_,
		_w18786_,
		_w18787_
	);
	LUT2 #(
		.INIT('h1)
	) name18256 (
		\u0_w_reg[3][27]/P0001 ,
		_w18787_,
		_w18788_
	);
	LUT2 #(
		.INIT('h1)
	) name18257 (
		_w16040_,
		_w17331_,
		_w18789_
	);
	LUT2 #(
		.INIT('h1)
	) name18258 (
		_w17428_,
		_w17820_,
		_w18790_
	);
	LUT2 #(
		.INIT('h8)
	) name18259 (
		_w18789_,
		_w18790_,
		_w18791_
	);
	LUT2 #(
		.INIT('h1)
	) name18260 (
		\u0_w_reg[3][26]/P0001 ,
		_w18791_,
		_w18792_
	);
	LUT2 #(
		.INIT('h1)
	) name18261 (
		_w18785_,
		_w18788_,
		_w18793_
	);
	LUT2 #(
		.INIT('h4)
	) name18262 (
		_w18792_,
		_w18793_,
		_w18794_
	);
	LUT2 #(
		.INIT('h4)
	) name18263 (
		_w18779_,
		_w18794_,
		_w18795_
	);
	LUT2 #(
		.INIT('h2)
	) name18264 (
		\u0_w_reg[3][24]/P0001 ,
		_w18795_,
		_w18796_
	);
	LUT2 #(
		.INIT('h2)
	) name18265 (
		\u0_w_reg[3][26]/P0001 ,
		_w16393_,
		_w18797_
	);
	LUT2 #(
		.INIT('h4)
	) name18266 (
		_w18082_,
		_w18127_,
		_w18798_
	);
	LUT2 #(
		.INIT('h1)
	) name18267 (
		_w18797_,
		_w18798_,
		_w18799_
	);
	LUT2 #(
		.INIT('h8)
	) name18268 (
		_w16033_,
		_w16098_,
		_w18800_
	);
	LUT2 #(
		.INIT('h1)
	) name18269 (
		\u0_w_reg[3][25]/P0001 ,
		_w16449_,
		_w18801_
	);
	LUT2 #(
		.INIT('h1)
	) name18270 (
		_w17824_,
		_w18800_,
		_w18802_
	);
	LUT2 #(
		.INIT('h8)
	) name18271 (
		_w18801_,
		_w18802_,
		_w18803_
	);
	LUT2 #(
		.INIT('h4)
	) name18272 (
		_w18799_,
		_w18803_,
		_w18804_
	);
	LUT2 #(
		.INIT('h1)
	) name18273 (
		_w16129_,
		_w18118_,
		_w18805_
	);
	LUT2 #(
		.INIT('h2)
	) name18274 (
		\u0_w_reg[3][26]/P0001 ,
		_w18805_,
		_w18806_
	);
	LUT2 #(
		.INIT('h4)
	) name18275 (
		\u0_w_reg[3][27]/P0001 ,
		_w16043_,
		_w18807_
	);
	LUT2 #(
		.INIT('h8)
	) name18276 (
		\u0_w_reg[3][28]/P0001 ,
		_w17422_,
		_w18808_
	);
	LUT2 #(
		.INIT('h1)
	) name18277 (
		_w16121_,
		_w18807_,
		_w18809_
	);
	LUT2 #(
		.INIT('h4)
	) name18278 (
		_w18808_,
		_w18809_,
		_w18810_
	);
	LUT2 #(
		.INIT('h1)
	) name18279 (
		\u0_w_reg[3][26]/P0001 ,
		_w18810_,
		_w18811_
	);
	LUT2 #(
		.INIT('h2)
	) name18280 (
		\u0_w_reg[3][25]/P0001 ,
		_w16144_,
		_w18812_
	);
	LUT2 #(
		.INIT('h8)
	) name18281 (
		_w16016_,
		_w18812_,
		_w18813_
	);
	LUT2 #(
		.INIT('h4)
	) name18282 (
		_w18806_,
		_w18813_,
		_w18814_
	);
	LUT2 #(
		.INIT('h4)
	) name18283 (
		_w18811_,
		_w18814_,
		_w18815_
	);
	LUT2 #(
		.INIT('h1)
	) name18284 (
		_w18804_,
		_w18815_,
		_w18816_
	);
	LUT2 #(
		.INIT('h8)
	) name18285 (
		_w16091_,
		_w16386_,
		_w18817_
	);
	LUT2 #(
		.INIT('h1)
	) name18286 (
		_w16039_,
		_w16052_,
		_w18818_
	);
	LUT2 #(
		.INIT('h2)
	) name18287 (
		_w16036_,
		_w18818_,
		_w18819_
	);
	LUT2 #(
		.INIT('h8)
	) name18288 (
		_w16117_,
		_w16428_,
		_w18820_
	);
	LUT2 #(
		.INIT('h1)
	) name18289 (
		_w16088_,
		_w16104_,
		_w18821_
	);
	LUT2 #(
		.INIT('h1)
	) name18290 (
		_w18817_,
		_w18820_,
		_w18822_
	);
	LUT2 #(
		.INIT('h8)
	) name18291 (
		_w18821_,
		_w18822_,
		_w18823_
	);
	LUT2 #(
		.INIT('h4)
	) name18292 (
		_w18819_,
		_w18823_,
		_w18824_
	);
	LUT2 #(
		.INIT('h4)
	) name18293 (
		_w18816_,
		_w18824_,
		_w18825_
	);
	LUT2 #(
		.INIT('h1)
	) name18294 (
		\u0_w_reg[3][24]/P0001 ,
		_w18825_,
		_w18826_
	);
	LUT2 #(
		.INIT('h4)
	) name18295 (
		_w16020_,
		_w17805_,
		_w18827_
	);
	LUT2 #(
		.INIT('h4)
	) name18296 (
		\u0_w_reg[3][31]/P0001 ,
		_w17866_,
		_w18828_
	);
	LUT2 #(
		.INIT('h1)
	) name18297 (
		_w16027_,
		_w18827_,
		_w18829_
	);
	LUT2 #(
		.INIT('h4)
	) name18298 (
		_w18828_,
		_w18829_,
		_w18830_
	);
	LUT2 #(
		.INIT('h2)
	) name18299 (
		_w16029_,
		_w18830_,
		_w18831_
	);
	LUT2 #(
		.INIT('h8)
	) name18300 (
		_w16099_,
		_w16411_,
		_w18832_
	);
	LUT2 #(
		.INIT('h1)
	) name18301 (
		_w16110_,
		_w18832_,
		_w18833_
	);
	LUT2 #(
		.INIT('h2)
	) name18302 (
		_w17871_,
		_w18833_,
		_w18834_
	);
	LUT2 #(
		.INIT('h1)
	) name18303 (
		_w16059_,
		_w16163_,
		_w18835_
	);
	LUT2 #(
		.INIT('h4)
	) name18304 (
		_w16038_,
		_w18835_,
		_w18836_
	);
	LUT2 #(
		.INIT('h4)
	) name18305 (
		\u0_w_reg[3][25]/P0001 ,
		_w16036_,
		_w18837_
	);
	LUT2 #(
		.INIT('h4)
	) name18306 (
		_w18836_,
		_w18837_,
		_w18838_
	);
	LUT2 #(
		.INIT('h1)
	) name18307 (
		_w16053_,
		_w17328_,
		_w18839_
	);
	LUT2 #(
		.INIT('h4)
	) name18308 (
		_w17337_,
		_w18839_,
		_w18840_
	);
	LUT2 #(
		.INIT('h1)
	) name18309 (
		\u0_w_reg[3][26]/P0001 ,
		_w18840_,
		_w18841_
	);
	LUT2 #(
		.INIT('h1)
	) name18310 (
		_w16047_,
		_w16376_,
		_w18842_
	);
	LUT2 #(
		.INIT('h4)
	) name18311 (
		_w18841_,
		_w18842_,
		_w18843_
	);
	LUT2 #(
		.INIT('h1)
	) name18312 (
		\u0_w_reg[3][25]/P0001 ,
		_w18843_,
		_w18844_
	);
	LUT2 #(
		.INIT('h1)
	) name18313 (
		_w16454_,
		_w17344_,
		_w18845_
	);
	LUT2 #(
		.INIT('h4)
	) name18314 (
		_w18834_,
		_w18845_,
		_w18846_
	);
	LUT2 #(
		.INIT('h4)
	) name18315 (
		_w18838_,
		_w18846_,
		_w18847_
	);
	LUT2 #(
		.INIT('h4)
	) name18316 (
		_w18831_,
		_w18847_,
		_w18848_
	);
	LUT2 #(
		.INIT('h4)
	) name18317 (
		_w18844_,
		_w18848_,
		_w18849_
	);
	LUT2 #(
		.INIT('h4)
	) name18318 (
		_w18796_,
		_w18849_,
		_w18850_
	);
	LUT2 #(
		.INIT('h4)
	) name18319 (
		_w18826_,
		_w18850_,
		_w18851_
	);
	LUT2 #(
		.INIT('h2)
	) name18320 (
		\u0_w_reg[0][1]/P0001 ,
		_w18851_,
		_w18852_
	);
	LUT2 #(
		.INIT('h4)
	) name18321 (
		\u0_w_reg[0][1]/P0001 ,
		_w18851_,
		_w18853_
	);
	LUT2 #(
		.INIT('h1)
	) name18322 (
		_w18852_,
		_w18853_,
		_w18854_
	);
	LUT2 #(
		.INIT('h2)
	) name18323 (
		\u0_w_reg[1][1]/P0001 ,
		\u0_w_reg[2][1]/P0001 ,
		_w18855_
	);
	LUT2 #(
		.INIT('h4)
	) name18324 (
		\u0_w_reg[1][1]/P0001 ,
		\u0_w_reg[2][1]/P0001 ,
		_w18856_
	);
	LUT2 #(
		.INIT('h1)
	) name18325 (
		_w18855_,
		_w18856_,
		_w18857_
	);
	LUT2 #(
		.INIT('h8)
	) name18326 (
		_w18854_,
		_w18857_,
		_w18858_
	);
	LUT2 #(
		.INIT('h1)
	) name18327 (
		_w18854_,
		_w18857_,
		_w18859_
	);
	LUT2 #(
		.INIT('h1)
	) name18328 (
		_w18858_,
		_w18859_,
		_w18860_
	);
	LUT2 #(
		.INIT('h4)
	) name18329 (
		ld_pad,
		_w18860_,
		_w18861_
	);
	LUT2 #(
		.INIT('h1)
	) name18330 (
		_w18774_,
		_w18861_,
		_w18862_
	);
	LUT2 #(
		.INIT('h4)
	) name18331 (
		\key[41]_pad ,
		ld_pad,
		_w18863_
	);
	LUT2 #(
		.INIT('h1)
	) name18332 (
		_w16503_,
		_w17532_,
		_w18864_
	);
	LUT2 #(
		.INIT('h4)
	) name18333 (
		_w17566_,
		_w18864_,
		_w18865_
	);
	LUT2 #(
		.INIT('h2)
	) name18334 (
		\u0_w_reg[3][2]/P0001 ,
		_w18865_,
		_w18866_
	);
	LUT2 #(
		.INIT('h2)
	) name18335 (
		_w17572_,
		_w18866_,
		_w18867_
	);
	LUT2 #(
		.INIT('h2)
	) name18336 (
		\u0_w_reg[3][1]/P0001 ,
		_w18867_,
		_w18868_
	);
	LUT2 #(
		.INIT('h2)
	) name18337 (
		_w16542_,
		_w16554_,
		_w18869_
	);
	LUT2 #(
		.INIT('h1)
	) name18338 (
		_w17500_,
		_w18869_,
		_w18870_
	);
	LUT2 #(
		.INIT('h1)
	) name18339 (
		\u0_w_reg[3][3]/P0001 ,
		_w18870_,
		_w18871_
	);
	LUT2 #(
		.INIT('h1)
	) name18340 (
		_w16484_,
		_w17500_,
		_w18872_
	);
	LUT2 #(
		.INIT('h1)
	) name18341 (
		_w17530_,
		_w18324_,
		_w18873_
	);
	LUT2 #(
		.INIT('h8)
	) name18342 (
		_w18872_,
		_w18873_,
		_w18874_
	);
	LUT2 #(
		.INIT('h1)
	) name18343 (
		\u0_w_reg[3][2]/P0001 ,
		_w18874_,
		_w18875_
	);
	LUT2 #(
		.INIT('h4)
	) name18344 (
		_w16552_,
		_w18194_,
		_w18876_
	);
	LUT2 #(
		.INIT('h1)
	) name18345 (
		_w16532_,
		_w17908_,
		_w18877_
	);
	LUT2 #(
		.INIT('h2)
	) name18346 (
		\u0_w_reg[3][5]/P0001 ,
		_w18877_,
		_w18878_
	);
	LUT2 #(
		.INIT('h1)
	) name18347 (
		_w18324_,
		_w18876_,
		_w18879_
	);
	LUT2 #(
		.INIT('h4)
	) name18348 (
		_w18878_,
		_w18879_,
		_w18880_
	);
	LUT2 #(
		.INIT('h1)
	) name18349 (
		\u0_w_reg[3][1]/P0001 ,
		_w18880_,
		_w18881_
	);
	LUT2 #(
		.INIT('h1)
	) name18350 (
		_w18871_,
		_w18875_,
		_w18882_
	);
	LUT2 #(
		.INIT('h4)
	) name18351 (
		_w18881_,
		_w18882_,
		_w18883_
	);
	LUT2 #(
		.INIT('h4)
	) name18352 (
		_w18868_,
		_w18883_,
		_w18884_
	);
	LUT2 #(
		.INIT('h2)
	) name18353 (
		\u0_w_reg[3][0]/P0001 ,
		_w18884_,
		_w18885_
	);
	LUT2 #(
		.INIT('h4)
	) name18354 (
		_w16512_,
		_w16573_,
		_w18886_
	);
	LUT2 #(
		.INIT('h8)
	) name18355 (
		_w16588_,
		_w16627_,
		_w18887_
	);
	LUT2 #(
		.INIT('h1)
	) name18356 (
		\u0_w_reg[3][1]/P0001 ,
		_w16616_,
		_w18888_
	);
	LUT2 #(
		.INIT('h1)
	) name18357 (
		_w16723_,
		_w17496_,
		_w18889_
	);
	LUT2 #(
		.INIT('h4)
	) name18358 (
		_w18887_,
		_w18889_,
		_w18890_
	);
	LUT2 #(
		.INIT('h4)
	) name18359 (
		_w18886_,
		_w18888_,
		_w18891_
	);
	LUT2 #(
		.INIT('h8)
	) name18360 (
		_w18890_,
		_w18891_,
		_w18892_
	);
	LUT2 #(
		.INIT('h4)
	) name18361 (
		\u0_w_reg[3][3]/P0001 ,
		_w16570_,
		_w18893_
	);
	LUT2 #(
		.INIT('h4)
	) name18362 (
		_w16580_,
		_w16653_,
		_w18894_
	);
	LUT2 #(
		.INIT('h1)
	) name18363 (
		_w18893_,
		_w18894_,
		_w18895_
	);
	LUT2 #(
		.INIT('h1)
	) name18364 (
		\u0_w_reg[3][2]/P0001 ,
		_w18895_,
		_w18896_
	);
	LUT2 #(
		.INIT('h8)
	) name18365 (
		_w16482_,
		_w16541_,
		_w18897_
	);
	LUT2 #(
		.INIT('h1)
	) name18366 (
		_w17915_,
		_w18897_,
		_w18898_
	);
	LUT2 #(
		.INIT('h2)
	) name18367 (
		\u0_w_reg[3][2]/P0001 ,
		_w18898_,
		_w18899_
	);
	LUT2 #(
		.INIT('h2)
	) name18368 (
		\u0_w_reg[3][1]/P0001 ,
		_w16701_,
		_w18900_
	);
	LUT2 #(
		.INIT('h8)
	) name18369 (
		_w18168_,
		_w18900_,
		_w18901_
	);
	LUT2 #(
		.INIT('h4)
	) name18370 (
		_w18899_,
		_w18901_,
		_w18902_
	);
	LUT2 #(
		.INIT('h4)
	) name18371 (
		_w18896_,
		_w18902_,
		_w18903_
	);
	LUT2 #(
		.INIT('h1)
	) name18372 (
		_w18892_,
		_w18903_,
		_w18904_
	);
	LUT2 #(
		.INIT('h4)
	) name18373 (
		\u0_w_reg[3][3]/P0001 ,
		_w17935_,
		_w18905_
	);
	LUT2 #(
		.INIT('h2)
	) name18374 (
		\u0_w_reg[3][2]/P0001 ,
		_w17959_,
		_w18906_
	);
	LUT2 #(
		.INIT('h1)
	) name18375 (
		_w16724_,
		_w18906_,
		_w18907_
	);
	LUT2 #(
		.INIT('h1)
	) name18376 (
		_w16506_,
		_w16548_,
		_w18908_
	);
	LUT2 #(
		.INIT('h2)
	) name18377 (
		_w16520_,
		_w18908_,
		_w18909_
	);
	LUT2 #(
		.INIT('h1)
	) name18378 (
		_w18210_,
		_w18909_,
		_w18910_
	);
	LUT2 #(
		.INIT('h4)
	) name18379 (
		_w18905_,
		_w18910_,
		_w18911_
	);
	LUT2 #(
		.INIT('h4)
	) name18380 (
		_w18907_,
		_w18911_,
		_w18912_
	);
	LUT2 #(
		.INIT('h4)
	) name18381 (
		_w18904_,
		_w18912_,
		_w18913_
	);
	LUT2 #(
		.INIT('h1)
	) name18382 (
		\u0_w_reg[3][0]/P0001 ,
		_w18913_,
		_w18914_
	);
	LUT2 #(
		.INIT('h1)
	) name18383 (
		_w16545_,
		_w17958_,
		_w18915_
	);
	LUT2 #(
		.INIT('h4)
	) name18384 (
		_w16624_,
		_w18915_,
		_w18916_
	);
	LUT2 #(
		.INIT('h1)
	) name18385 (
		\u0_w_reg[3][2]/P0001 ,
		_w18916_,
		_w18917_
	);
	LUT2 #(
		.INIT('h1)
	) name18386 (
		_w16732_,
		_w17959_,
		_w18918_
	);
	LUT2 #(
		.INIT('h4)
	) name18387 (
		_w18917_,
		_w18918_,
		_w18919_
	);
	LUT2 #(
		.INIT('h1)
	) name18388 (
		\u0_w_reg[3][1]/P0001 ,
		_w18919_,
		_w18920_
	);
	LUT2 #(
		.INIT('h1)
	) name18389 (
		_w16525_,
		_w18271_,
		_w18921_
	);
	LUT2 #(
		.INIT('h1)
	) name18390 (
		\u0_w_reg[3][6]/P0001 ,
		_w18921_,
		_w18922_
	);
	LUT2 #(
		.INIT('h1)
	) name18391 (
		_w17519_,
		_w18226_,
		_w18923_
	);
	LUT2 #(
		.INIT('h4)
	) name18392 (
		_w18279_,
		_w18923_,
		_w18924_
	);
	LUT2 #(
		.INIT('h4)
	) name18393 (
		\u0_w_reg[3][3]/P0001 ,
		_w16621_,
		_w18925_
	);
	LUT2 #(
		.INIT('h4)
	) name18394 (
		_w18924_,
		_w18925_,
		_w18926_
	);
	LUT2 #(
		.INIT('h1)
	) name18395 (
		_w16627_,
		_w16687_,
		_w18927_
	);
	LUT2 #(
		.INIT('h2)
	) name18396 (
		\u0_w_reg[3][3]/P0001 ,
		_w18927_,
		_w18928_
	);
	LUT2 #(
		.INIT('h2)
	) name18397 (
		_w17898_,
		_w18928_,
		_w18929_
	);
	LUT2 #(
		.INIT('h1)
	) name18398 (
		_w16481_,
		_w16482_,
		_w18930_
	);
	LUT2 #(
		.INIT('h1)
	) name18399 (
		\u0_w_reg[3][6]/P0001 ,
		_w16528_,
		_w18931_
	);
	LUT2 #(
		.INIT('h4)
	) name18400 (
		_w18930_,
		_w18931_,
		_w18932_
	);
	LUT2 #(
		.INIT('h1)
	) name18401 (
		\u0_w_reg[3][2]/P0001 ,
		_w16701_,
		_w18933_
	);
	LUT2 #(
		.INIT('h4)
	) name18402 (
		_w17517_,
		_w18933_,
		_w18934_
	);
	LUT2 #(
		.INIT('h4)
	) name18403 (
		_w18932_,
		_w18934_,
		_w18935_
	);
	LUT2 #(
		.INIT('h2)
	) name18404 (
		\u0_w_reg[3][1]/P0001 ,
		_w18929_,
		_w18936_
	);
	LUT2 #(
		.INIT('h4)
	) name18405 (
		_w18935_,
		_w18936_,
		_w18937_
	);
	LUT2 #(
		.INIT('h1)
	) name18406 (
		_w18922_,
		_w18926_,
		_w18938_
	);
	LUT2 #(
		.INIT('h4)
	) name18407 (
		_w18937_,
		_w18938_,
		_w18939_
	);
	LUT2 #(
		.INIT('h4)
	) name18408 (
		_w18920_,
		_w18939_,
		_w18940_
	);
	LUT2 #(
		.INIT('h4)
	) name18409 (
		_w18885_,
		_w18940_,
		_w18941_
	);
	LUT2 #(
		.INIT('h4)
	) name18410 (
		_w18914_,
		_w18941_,
		_w18942_
	);
	LUT2 #(
		.INIT('h2)
	) name18411 (
		\u0_w_reg[0][9]/P0001 ,
		_w18942_,
		_w18943_
	);
	LUT2 #(
		.INIT('h4)
	) name18412 (
		\u0_w_reg[0][9]/P0001 ,
		_w18942_,
		_w18944_
	);
	LUT2 #(
		.INIT('h1)
	) name18413 (
		_w18943_,
		_w18944_,
		_w18945_
	);
	LUT2 #(
		.INIT('h2)
	) name18414 (
		\u0_w_reg[1][9]/P0001 ,
		\u0_w_reg[2][9]/P0001 ,
		_w18946_
	);
	LUT2 #(
		.INIT('h4)
	) name18415 (
		\u0_w_reg[1][9]/P0001 ,
		\u0_w_reg[2][9]/P0001 ,
		_w18947_
	);
	LUT2 #(
		.INIT('h1)
	) name18416 (
		_w18946_,
		_w18947_,
		_w18948_
	);
	LUT2 #(
		.INIT('h8)
	) name18417 (
		_w18945_,
		_w18948_,
		_w18949_
	);
	LUT2 #(
		.INIT('h1)
	) name18418 (
		_w18945_,
		_w18948_,
		_w18950_
	);
	LUT2 #(
		.INIT('h1)
	) name18419 (
		_w18949_,
		_w18950_,
		_w18951_
	);
	LUT2 #(
		.INIT('h4)
	) name18420 (
		ld_pad,
		_w18951_,
		_w18952_
	);
	LUT2 #(
		.INIT('h1)
	) name18421 (
		_w18863_,
		_w18952_,
		_w18953_
	);
	LUT2 #(
		.INIT('h4)
	) name18422 (
		ld_pad,
		_w16764_,
		_w18954_
	);
	LUT2 #(
		.INIT('h8)
	) name18423 (
		\key[108]_pad ,
		ld_pad,
		_w18955_
	);
	LUT2 #(
		.INIT('h1)
	) name18424 (
		_w18954_,
		_w18955_,
		_w18956_
	);
	LUT2 #(
		.INIT('h1)
	) name18425 (
		\u0_w_reg[1][12]/P0001 ,
		_w16764_,
		_w18957_
	);
	LUT2 #(
		.INIT('h8)
	) name18426 (
		\u0_w_reg[1][12]/P0001 ,
		_w16764_,
		_w18958_
	);
	LUT2 #(
		.INIT('h1)
	) name18427 (
		ld_pad,
		_w18957_,
		_w18959_
	);
	LUT2 #(
		.INIT('h4)
	) name18428 (
		_w18958_,
		_w18959_,
		_w18960_
	);
	LUT2 #(
		.INIT('h8)
	) name18429 (
		\key[76]_pad ,
		ld_pad,
		_w18961_
	);
	LUT2 #(
		.INIT('h1)
	) name18430 (
		_w18960_,
		_w18961_,
		_w18962_
	);
	LUT2 #(
		.INIT('h1)
	) name18431 (
		_w15717_,
		_w15939_,
		_w18963_
	);
	LUT2 #(
		.INIT('h4)
	) name18432 (
		_w18051_,
		_w18963_,
		_w18964_
	);
	LUT2 #(
		.INIT('h1)
	) name18433 (
		\u0_w_reg[3][10]/P0001 ,
		_w18964_,
		_w18965_
	);
	LUT2 #(
		.INIT('h8)
	) name18434 (
		_w15817_,
		_w15974_,
		_w18966_
	);
	LUT2 #(
		.INIT('h4)
	) name18435 (
		\u0_w_reg[3][15]/P0001 ,
		_w15751_,
		_w18967_
	);
	LUT2 #(
		.INIT('h1)
	) name18436 (
		_w15805_,
		_w15862_,
		_w18968_
	);
	LUT2 #(
		.INIT('h4)
	) name18437 (
		_w18967_,
		_w18968_,
		_w18969_
	);
	LUT2 #(
		.INIT('h2)
	) name18438 (
		\u0_w_reg[3][10]/P0001 ,
		_w18969_,
		_w18970_
	);
	LUT2 #(
		.INIT('h1)
	) name18439 (
		_w15771_,
		_w15802_,
		_w18971_
	);
	LUT2 #(
		.INIT('h1)
	) name18440 (
		\u0_w_reg[3][10]/P0001 ,
		_w18971_,
		_w18972_
	);
	LUT2 #(
		.INIT('h1)
	) name18441 (
		_w15863_,
		_w17742_,
		_w18973_
	);
	LUT2 #(
		.INIT('h8)
	) name18442 (
		_w15760_,
		_w18973_,
		_w18974_
	);
	LUT2 #(
		.INIT('h4)
	) name18443 (
		_w18972_,
		_w18974_,
		_w18975_
	);
	LUT2 #(
		.INIT('h1)
	) name18444 (
		_w15737_,
		_w15846_,
		_w18976_
	);
	LUT2 #(
		.INIT('h1)
	) name18445 (
		\u0_w_reg[3][10]/P0001 ,
		_w18976_,
		_w18977_
	);
	LUT2 #(
		.INIT('h4)
	) name18446 (
		_w15781_,
		_w17746_,
		_w18978_
	);
	LUT2 #(
		.INIT('h4)
	) name18447 (
		_w18977_,
		_w18978_,
		_w18979_
	);
	LUT2 #(
		.INIT('h1)
	) name18448 (
		_w18975_,
		_w18979_,
		_w18980_
	);
	LUT2 #(
		.INIT('h2)
	) name18449 (
		\u0_w_reg[3][8]/P0001 ,
		_w17681_,
		_w18981_
	);
	LUT2 #(
		.INIT('h4)
	) name18450 (
		_w18966_,
		_w18981_,
		_w18982_
	);
	LUT2 #(
		.INIT('h4)
	) name18451 (
		_w18965_,
		_w18982_,
		_w18983_
	);
	LUT2 #(
		.INIT('h4)
	) name18452 (
		_w18970_,
		_w18983_,
		_w18984_
	);
	LUT2 #(
		.INIT('h4)
	) name18453 (
		_w18980_,
		_w18984_,
		_w18985_
	);
	LUT2 #(
		.INIT('h2)
	) name18454 (
		\u0_w_reg[3][13]/P0001 ,
		_w15724_,
		_w18986_
	);
	LUT2 #(
		.INIT('h8)
	) name18455 (
		_w15742_,
		_w18986_,
		_w18987_
	);
	LUT2 #(
		.INIT('h1)
	) name18456 (
		_w15989_,
		_w18987_,
		_w18988_
	);
	LUT2 #(
		.INIT('h1)
	) name18457 (
		\u0_w_reg[3][10]/P0001 ,
		_w18988_,
		_w18989_
	);
	LUT2 #(
		.INIT('h8)
	) name18458 (
		_w15893_,
		_w15946_,
		_w18990_
	);
	LUT2 #(
		.INIT('h2)
	) name18459 (
		\u0_w_reg[3][9]/P0001 ,
		_w15920_,
		_w18991_
	);
	LUT2 #(
		.INIT('h4)
	) name18460 (
		_w17611_,
		_w18991_,
		_w18992_
	);
	LUT2 #(
		.INIT('h4)
	) name18461 (
		_w18990_,
		_w18992_,
		_w18993_
	);
	LUT2 #(
		.INIT('h4)
	) name18462 (
		_w18989_,
		_w18993_,
		_w18994_
	);
	LUT2 #(
		.INIT('h8)
	) name18463 (
		_w15741_,
		_w15847_,
		_w18995_
	);
	LUT2 #(
		.INIT('h8)
	) name18464 (
		\u0_w_reg[3][12]/P0001 ,
		_w15791_,
		_w18996_
	);
	LUT2 #(
		.INIT('h1)
	) name18465 (
		\u0_w_reg[3][9]/P0001 ,
		_w15804_,
		_w18997_
	);
	LUT2 #(
		.INIT('h4)
	) name18466 (
		_w15865_,
		_w18997_,
		_w18998_
	);
	LUT2 #(
		.INIT('h1)
	) name18467 (
		_w18995_,
		_w18996_,
		_w18999_
	);
	LUT2 #(
		.INIT('h8)
	) name18468 (
		_w18998_,
		_w18999_,
		_w19000_
	);
	LUT2 #(
		.INIT('h1)
	) name18469 (
		_w18994_,
		_w19000_,
		_w19001_
	);
	LUT2 #(
		.INIT('h1)
	) name18470 (
		_w15731_,
		_w17672_,
		_w19002_
	);
	LUT2 #(
		.INIT('h1)
	) name18471 (
		\u0_w_reg[3][11]/P0001 ,
		_w19002_,
		_w19003_
	);
	LUT2 #(
		.INIT('h1)
	) name18472 (
		_w15710_,
		_w18628_,
		_w19004_
	);
	LUT2 #(
		.INIT('h2)
	) name18473 (
		\u0_w_reg[3][10]/P0001 ,
		_w19004_,
		_w19005_
	);
	LUT2 #(
		.INIT('h1)
	) name18474 (
		\u0_w_reg[3][8]/P0001 ,
		_w19003_,
		_w19006_
	);
	LUT2 #(
		.INIT('h4)
	) name18475 (
		_w19005_,
		_w19006_,
		_w19007_
	);
	LUT2 #(
		.INIT('h4)
	) name18476 (
		_w19001_,
		_w19007_,
		_w19008_
	);
	LUT2 #(
		.INIT('h1)
	) name18477 (
		_w18985_,
		_w19008_,
		_w19009_
	);
	LUT2 #(
		.INIT('h4)
	) name18478 (
		\u0_w_reg[3][10]/P0001 ,
		_w15976_,
		_w19010_
	);
	LUT2 #(
		.INIT('h1)
	) name18479 (
		_w18996_,
		_w19010_,
		_w19011_
	);
	LUT2 #(
		.INIT('h2)
	) name18480 (
		\u0_w_reg[3][11]/P0001 ,
		_w19011_,
		_w19012_
	);
	LUT2 #(
		.INIT('h2)
	) name18481 (
		_w15756_,
		_w15907_,
		_w19013_
	);
	LUT2 #(
		.INIT('h1)
	) name18482 (
		_w15715_,
		_w17682_,
		_w19014_
	);
	LUT2 #(
		.INIT('h4)
	) name18483 (
		_w17719_,
		_w19014_,
		_w19015_
	);
	LUT2 #(
		.INIT('h4)
	) name18484 (
		_w19013_,
		_w19015_,
		_w19016_
	);
	LUT2 #(
		.INIT('h2)
	) name18485 (
		\u0_w_reg[3][10]/P0001 ,
		_w19016_,
		_w19017_
	);
	LUT2 #(
		.INIT('h2)
	) name18486 (
		_w15708_,
		_w15822_,
		_w19018_
	);
	LUT2 #(
		.INIT('h8)
	) name18487 (
		_w15847_,
		_w19018_,
		_w19019_
	);
	LUT2 #(
		.INIT('h1)
	) name18488 (
		\u0_w_reg[3][9]/P0001 ,
		_w17722_,
		_w19020_
	);
	LUT2 #(
		.INIT('h1)
	) name18489 (
		_w17758_,
		_w18708_,
		_w19021_
	);
	LUT2 #(
		.INIT('h4)
	) name18490 (
		_w19019_,
		_w19021_,
		_w19022_
	);
	LUT2 #(
		.INIT('h8)
	) name18491 (
		_w19020_,
		_w19022_,
		_w19023_
	);
	LUT2 #(
		.INIT('h4)
	) name18492 (
		_w19017_,
		_w19023_,
		_w19024_
	);
	LUT2 #(
		.INIT('h1)
	) name18493 (
		_w15805_,
		_w15832_,
		_w19025_
	);
	LUT2 #(
		.INIT('h2)
	) name18494 (
		_w15847_,
		_w19025_,
		_w19026_
	);
	LUT2 #(
		.INIT('h8)
	) name18495 (
		\u0_w_reg[3][12]/P0001 ,
		_w17743_,
		_w19027_
	);
	LUT2 #(
		.INIT('h8)
	) name18496 (
		_w15849_,
		_w17650_,
		_w19028_
	);
	LUT2 #(
		.INIT('h1)
	) name18497 (
		_w17656_,
		_w18026_,
		_w19029_
	);
	LUT2 #(
		.INIT('h1)
	) name18498 (
		_w19027_,
		_w19028_,
		_w19030_
	);
	LUT2 #(
		.INIT('h8)
	) name18499 (
		_w19029_,
		_w19030_,
		_w19031_
	);
	LUT2 #(
		.INIT('h2)
	) name18500 (
		_w18599_,
		_w19026_,
		_w19032_
	);
	LUT2 #(
		.INIT('h8)
	) name18501 (
		_w19031_,
		_w19032_,
		_w19033_
	);
	LUT2 #(
		.INIT('h1)
	) name18502 (
		_w19024_,
		_w19033_,
		_w19034_
	);
	LUT2 #(
		.INIT('h1)
	) name18503 (
		_w19012_,
		_w19034_,
		_w19035_
	);
	LUT2 #(
		.INIT('h4)
	) name18504 (
		_w19009_,
		_w19035_,
		_w19036_
	);
	LUT2 #(
		.INIT('h2)
	) name18505 (
		\u0_w_reg[0][20]/P0001 ,
		_w19036_,
		_w19037_
	);
	LUT2 #(
		.INIT('h4)
	) name18506 (
		\u0_w_reg[0][20]/P0001 ,
		_w19036_,
		_w19038_
	);
	LUT2 #(
		.INIT('h1)
	) name18507 (
		_w19037_,
		_w19038_,
		_w19039_
	);
	LUT2 #(
		.INIT('h8)
	) name18508 (
		\u0_w_reg[1][20]/P0001 ,
		_w19039_,
		_w19040_
	);
	LUT2 #(
		.INIT('h1)
	) name18509 (
		\u0_w_reg[1][20]/P0001 ,
		_w19039_,
		_w19041_
	);
	LUT2 #(
		.INIT('h1)
	) name18510 (
		_w19040_,
		_w19041_,
		_w19042_
	);
	LUT2 #(
		.INIT('h8)
	) name18511 (
		\u0_w_reg[2][20]/P0001 ,
		_w19042_,
		_w19043_
	);
	LUT2 #(
		.INIT('h1)
	) name18512 (
		\u0_w_reg[2][20]/P0001 ,
		_w19042_,
		_w19044_
	);
	LUT2 #(
		.INIT('h1)
	) name18513 (
		_w19043_,
		_w19044_,
		_w19045_
	);
	LUT2 #(
		.INIT('h4)
	) name18514 (
		ld_pad,
		_w19045_,
		_w19046_
	);
	LUT2 #(
		.INIT('h8)
	) name18515 (
		\key[52]_pad ,
		ld_pad,
		_w19047_
	);
	LUT2 #(
		.INIT('h1)
	) name18516 (
		_w19046_,
		_w19047_,
		_w19048_
	);
	LUT2 #(
		.INIT('h4)
	) name18517 (
		\key[36]_pad ,
		ld_pad,
		_w19049_
	);
	LUT2 #(
		.INIT('h1)
	) name18518 (
		_w16118_,
		_w17807_,
		_w19050_
	);
	LUT2 #(
		.INIT('h1)
	) name18519 (
		\u0_w_reg[3][27]/P0001 ,
		_w19050_,
		_w19051_
	);
	LUT2 #(
		.INIT('h8)
	) name18520 (
		_w16019_,
		_w16087_,
		_w19052_
	);
	LUT2 #(
		.INIT('h1)
	) name18521 (
		_w17287_,
		_w19052_,
		_w19053_
	);
	LUT2 #(
		.INIT('h2)
	) name18522 (
		\u0_w_reg[3][26]/P0001 ,
		_w19053_,
		_w19054_
	);
	LUT2 #(
		.INIT('h8)
	) name18523 (
		\u0_w_reg[3][28]/P0001 ,
		_w16142_,
		_w19055_
	);
	LUT2 #(
		.INIT('h4)
	) name18524 (
		\u0_w_reg[3][26]/P0001 ,
		_w17428_,
		_w19056_
	);
	LUT2 #(
		.INIT('h1)
	) name18525 (
		_w17339_,
		_w18130_,
		_w19057_
	);
	LUT2 #(
		.INIT('h4)
	) name18526 (
		_w19055_,
		_w19057_,
		_w19058_
	);
	LUT2 #(
		.INIT('h4)
	) name18527 (
		_w19056_,
		_w19058_,
		_w19059_
	);
	LUT2 #(
		.INIT('h1)
	) name18528 (
		\u0_w_reg[3][25]/P0001 ,
		_w19059_,
		_w19060_
	);
	LUT2 #(
		.INIT('h8)
	) name18529 (
		_w16036_,
		_w16388_,
		_w19061_
	);
	LUT2 #(
		.INIT('h8)
	) name18530 (
		\u0_w_reg[3][26]/P0001 ,
		_w16058_,
		_w19062_
	);
	LUT2 #(
		.INIT('h4)
	) name18531 (
		_w16032_,
		_w16049_,
		_w19063_
	);
	LUT2 #(
		.INIT('h1)
	) name18532 (
		_w16443_,
		_w19063_,
		_w19064_
	);
	LUT2 #(
		.INIT('h1)
	) name18533 (
		\u0_w_reg[3][26]/P0001 ,
		_w19064_,
		_w19065_
	);
	LUT2 #(
		.INIT('h1)
	) name18534 (
		_w16403_,
		_w19061_,
		_w19066_
	);
	LUT2 #(
		.INIT('h4)
	) name18535 (
		_w19062_,
		_w19066_,
		_w19067_
	);
	LUT2 #(
		.INIT('h4)
	) name18536 (
		_w19065_,
		_w19067_,
		_w19068_
	);
	LUT2 #(
		.INIT('h2)
	) name18537 (
		\u0_w_reg[3][25]/P0001 ,
		_w19068_,
		_w19069_
	);
	LUT2 #(
		.INIT('h1)
	) name18538 (
		_w19051_,
		_w19054_,
		_w19070_
	);
	LUT2 #(
		.INIT('h4)
	) name18539 (
		_w19060_,
		_w19070_,
		_w19071_
	);
	LUT2 #(
		.INIT('h4)
	) name18540 (
		_w19069_,
		_w19071_,
		_w19072_
	);
	LUT2 #(
		.INIT('h1)
	) name18541 (
		\u0_w_reg[3][24]/P0001 ,
		_w19072_,
		_w19073_
	);
	LUT2 #(
		.INIT('h1)
	) name18542 (
		_w16013_,
		_w17276_,
		_w19074_
	);
	LUT2 #(
		.INIT('h4)
	) name18543 (
		_w16376_,
		_w19074_,
		_w19075_
	);
	LUT2 #(
		.INIT('h4)
	) name18544 (
		_w17806_,
		_w19075_,
		_w19076_
	);
	LUT2 #(
		.INIT('h4)
	) name18545 (
		_w17826_,
		_w19076_,
		_w19077_
	);
	LUT2 #(
		.INIT('h2)
	) name18546 (
		\u0_w_reg[3][26]/P0001 ,
		_w19077_,
		_w19078_
	);
	LUT2 #(
		.INIT('h2)
	) name18547 (
		_w16019_,
		_w16039_,
		_w19079_
	);
	LUT2 #(
		.INIT('h8)
	) name18548 (
		_w16386_,
		_w19079_,
		_w19080_
	);
	LUT2 #(
		.INIT('h1)
	) name18549 (
		_w16111_,
		_w17474_,
		_w19081_
	);
	LUT2 #(
		.INIT('h1)
	) name18550 (
		_w18820_,
		_w19080_,
		_w19082_
	);
	LUT2 #(
		.INIT('h8)
	) name18551 (
		_w19081_,
		_w19082_,
		_w19083_
	);
	LUT2 #(
		.INIT('h4)
	) name18552 (
		_w19078_,
		_w19083_,
		_w19084_
	);
	LUT2 #(
		.INIT('h1)
	) name18553 (
		\u0_w_reg[3][25]/P0001 ,
		_w19084_,
		_w19085_
	);
	LUT2 #(
		.INIT('h8)
	) name18554 (
		_w16036_,
		_w17259_,
		_w19086_
	);
	LUT2 #(
		.INIT('h1)
	) name18555 (
		_w16120_,
		_w16428_,
		_w19087_
	);
	LUT2 #(
		.INIT('h2)
	) name18556 (
		_w16386_,
		_w19087_,
		_w19088_
	);
	LUT2 #(
		.INIT('h4)
	) name18557 (
		_w16051_,
		_w16117_,
		_w19089_
	);
	LUT2 #(
		.INIT('h1)
	) name18558 (
		_w16044_,
		_w17443_,
		_w19090_
	);
	LUT2 #(
		.INIT('h4)
	) name18559 (
		_w19089_,
		_w19090_,
		_w19091_
	);
	LUT2 #(
		.INIT('h1)
	) name18560 (
		\u0_w_reg[3][29]/P0001 ,
		_w19091_,
		_w19092_
	);
	LUT2 #(
		.INIT('h1)
	) name18561 (
		_w18110_,
		_w19086_,
		_w19093_
	);
	LUT2 #(
		.INIT('h4)
	) name18562 (
		_w19088_,
		_w19093_,
		_w19094_
	);
	LUT2 #(
		.INIT('h4)
	) name18563 (
		_w19092_,
		_w19094_,
		_w19095_
	);
	LUT2 #(
		.INIT('h2)
	) name18564 (
		\u0_w_reg[3][25]/P0001 ,
		_w19095_,
		_w19096_
	);
	LUT2 #(
		.INIT('h4)
	) name18565 (
		\u0_w_reg[3][26]/P0001 ,
		_w16040_,
		_w19097_
	);
	LUT2 #(
		.INIT('h1)
	) name18566 (
		_w19055_,
		_w19097_,
		_w19098_
	);
	LUT2 #(
		.INIT('h2)
	) name18567 (
		\u0_w_reg[3][27]/P0001 ,
		_w19098_,
		_w19099_
	);
	LUT2 #(
		.INIT('h8)
	) name18568 (
		_w16032_,
		_w16103_,
		_w19100_
	);
	LUT2 #(
		.INIT('h4)
	) name18569 (
		\u0_w_reg[3][25]/P0001 ,
		_w16091_,
		_w19101_
	);
	LUT2 #(
		.INIT('h1)
	) name18570 (
		_w16428_,
		_w19101_,
		_w19102_
	);
	LUT2 #(
		.INIT('h8)
	) name18571 (
		_w18090_,
		_w19102_,
		_w19103_
	);
	LUT2 #(
		.INIT('h1)
	) name18572 (
		_w16015_,
		_w17463_,
		_w19104_
	);
	LUT2 #(
		.INIT('h8)
	) name18573 (
		_w18101_,
		_w19104_,
		_w19105_
	);
	LUT2 #(
		.INIT('h1)
	) name18574 (
		_w19103_,
		_w19105_,
		_w19106_
	);
	LUT2 #(
		.INIT('h8)
	) name18575 (
		\u0_w_reg[3][31]/P0001 ,
		_w16026_,
		_w19107_
	);
	LUT2 #(
		.INIT('h1)
	) name18576 (
		_w16066_,
		_w19107_,
		_w19108_
	);
	LUT2 #(
		.INIT('h1)
	) name18577 (
		\u0_w_reg[3][26]/P0001 ,
		_w19108_,
		_w19109_
	);
	LUT2 #(
		.INIT('h1)
	) name18578 (
		\u0_w_reg[3][25]/P0001 ,
		_w16146_,
		_w19110_
	);
	LUT2 #(
		.INIT('h4)
	) name18579 (
		_w17804_,
		_w19110_,
		_w19111_
	);
	LUT2 #(
		.INIT('h4)
	) name18580 (
		_w19109_,
		_w19111_,
		_w19112_
	);
	LUT2 #(
		.INIT('h1)
	) name18581 (
		_w16366_,
		_w16439_,
		_w19113_
	);
	LUT2 #(
		.INIT('h1)
	) name18582 (
		\u0_w_reg[3][26]/P0001 ,
		_w19113_,
		_w19114_
	);
	LUT2 #(
		.INIT('h2)
	) name18583 (
		\u0_w_reg[3][25]/P0001 ,
		_w17803_,
		_w19115_
	);
	LUT2 #(
		.INIT('h4)
	) name18584 (
		_w16053_,
		_w19115_,
		_w19116_
	);
	LUT2 #(
		.INIT('h4)
	) name18585 (
		_w17464_,
		_w19116_,
		_w19117_
	);
	LUT2 #(
		.INIT('h4)
	) name18586 (
		_w19114_,
		_w19117_,
		_w19118_
	);
	LUT2 #(
		.INIT('h1)
	) name18587 (
		_w19112_,
		_w19118_,
		_w19119_
	);
	LUT2 #(
		.INIT('h1)
	) name18588 (
		_w16106_,
		_w19100_,
		_w19120_
	);
	LUT2 #(
		.INIT('h4)
	) name18589 (
		_w19106_,
		_w19120_,
		_w19121_
	);
	LUT2 #(
		.INIT('h4)
	) name18590 (
		_w19119_,
		_w19121_,
		_w19122_
	);
	LUT2 #(
		.INIT('h2)
	) name18591 (
		\u0_w_reg[3][24]/P0001 ,
		_w19122_,
		_w19123_
	);
	LUT2 #(
		.INIT('h1)
	) name18592 (
		_w19096_,
		_w19099_,
		_w19124_
	);
	LUT2 #(
		.INIT('h4)
	) name18593 (
		_w19085_,
		_w19124_,
		_w19125_
	);
	LUT2 #(
		.INIT('h4)
	) name18594 (
		_w19123_,
		_w19125_,
		_w19126_
	);
	LUT2 #(
		.INIT('h4)
	) name18595 (
		_w19073_,
		_w19126_,
		_w19127_
	);
	LUT2 #(
		.INIT('h2)
	) name18596 (
		\u0_w_reg[0][4]/P0001 ,
		_w19127_,
		_w19128_
	);
	LUT2 #(
		.INIT('h4)
	) name18597 (
		\u0_w_reg[0][4]/P0001 ,
		_w19127_,
		_w19129_
	);
	LUT2 #(
		.INIT('h1)
	) name18598 (
		_w19128_,
		_w19129_,
		_w19130_
	);
	LUT2 #(
		.INIT('h2)
	) name18599 (
		\u0_w_reg[1][4]/P0001 ,
		\u0_w_reg[2][4]/P0001 ,
		_w19131_
	);
	LUT2 #(
		.INIT('h4)
	) name18600 (
		\u0_w_reg[1][4]/P0001 ,
		\u0_w_reg[2][4]/P0001 ,
		_w19132_
	);
	LUT2 #(
		.INIT('h1)
	) name18601 (
		_w19131_,
		_w19132_,
		_w19133_
	);
	LUT2 #(
		.INIT('h8)
	) name18602 (
		_w19130_,
		_w19133_,
		_w19134_
	);
	LUT2 #(
		.INIT('h1)
	) name18603 (
		_w19130_,
		_w19133_,
		_w19135_
	);
	LUT2 #(
		.INIT('h1)
	) name18604 (
		_w19134_,
		_w19135_,
		_w19136_
	);
	LUT2 #(
		.INIT('h4)
	) name18605 (
		ld_pad,
		_w19136_,
		_w19137_
	);
	LUT2 #(
		.INIT('h1)
	) name18606 (
		_w19049_,
		_w19137_,
		_w19138_
	);
	LUT2 #(
		.INIT('h4)
	) name18607 (
		\u0_w_reg[3][12]/P0001 ,
		_w16770_,
		_w19139_
	);
	LUT2 #(
		.INIT('h2)
	) name18608 (
		\u0_w_reg[3][12]/P0001 ,
		_w16770_,
		_w19140_
	);
	LUT2 #(
		.INIT('h1)
	) name18609 (
		ld_pad,
		_w19139_,
		_w19141_
	);
	LUT2 #(
		.INIT('h4)
	) name18610 (
		_w19140_,
		_w19141_,
		_w19142_
	);
	LUT2 #(
		.INIT('h8)
	) name18611 (
		\key[12]_pad ,
		ld_pad,
		_w19143_
	);
	LUT2 #(
		.INIT('h1)
	) name18612 (
		_w19142_,
		_w19143_,
		_w19144_
	);
	LUT2 #(
		.INIT('h1)
	) name18613 (
		_w15637_,
		_w18447_,
		_w19145_
	);
	LUT2 #(
		.INIT('h1)
	) name18614 (
		\u0_w_reg[3][21]/P0001 ,
		_w19145_,
		_w19146_
	);
	LUT2 #(
		.INIT('h1)
	) name18615 (
		_w15540_,
		_w19146_,
		_w19147_
	);
	LUT2 #(
		.INIT('h1)
	) name18616 (
		\u0_w_reg[3][18]/P0001 ,
		_w19147_,
		_w19148_
	);
	LUT2 #(
		.INIT('h8)
	) name18617 (
		_w15628_,
		_w16281_,
		_w19149_
	);
	LUT2 #(
		.INIT('h8)
	) name18618 (
		_w15504_,
		_w16297_,
		_w19150_
	);
	LUT2 #(
		.INIT('h8)
	) name18619 (
		_w15511_,
		_w15551_,
		_w19151_
	);
	LUT2 #(
		.INIT('h1)
	) name18620 (
		_w15522_,
		_w15582_,
		_w19152_
	);
	LUT2 #(
		.INIT('h1)
	) name18621 (
		\u0_w_reg[3][18]/P0001 ,
		_w19152_,
		_w19153_
	);
	LUT2 #(
		.INIT('h1)
	) name18622 (
		_w15587_,
		_w16919_,
		_w19154_
	);
	LUT2 #(
		.INIT('h4)
	) name18623 (
		_w19153_,
		_w19154_,
		_w19155_
	);
	LUT2 #(
		.INIT('h1)
	) name18624 (
		\u0_w_reg[3][17]/P0001 ,
		_w19155_,
		_w19156_
	);
	LUT2 #(
		.INIT('h1)
	) name18625 (
		_w15603_,
		_w16262_,
		_w19157_
	);
	LUT2 #(
		.INIT('h1)
	) name18626 (
		\u0_w_reg[3][18]/P0001 ,
		_w19157_,
		_w19158_
	);
	LUT2 #(
		.INIT('h1)
	) name18627 (
		_w15558_,
		_w16918_,
		_w19159_
	);
	LUT2 #(
		.INIT('h4)
	) name18628 (
		_w15658_,
		_w19159_,
		_w19160_
	);
	LUT2 #(
		.INIT('h4)
	) name18629 (
		_w19158_,
		_w19160_,
		_w19161_
	);
	LUT2 #(
		.INIT('h2)
	) name18630 (
		\u0_w_reg[3][17]/P0001 ,
		_w19161_,
		_w19162_
	);
	LUT2 #(
		.INIT('h1)
	) name18631 (
		_w19150_,
		_w19151_,
		_w19163_
	);
	LUT2 #(
		.INIT('h4)
	) name18632 (
		_w16845_,
		_w19163_,
		_w19164_
	);
	LUT2 #(
		.INIT('h1)
	) name18633 (
		_w17019_,
		_w19149_,
		_w19165_
	);
	LUT2 #(
		.INIT('h8)
	) name18634 (
		_w19164_,
		_w19165_,
		_w19166_
	);
	LUT2 #(
		.INIT('h4)
	) name18635 (
		_w19148_,
		_w19166_,
		_w19167_
	);
	LUT2 #(
		.INIT('h4)
	) name18636 (
		_w19156_,
		_w19167_,
		_w19168_
	);
	LUT2 #(
		.INIT('h4)
	) name18637 (
		_w19162_,
		_w19168_,
		_w19169_
	);
	LUT2 #(
		.INIT('h2)
	) name18638 (
		\u0_w_reg[3][16]/P0001 ,
		_w19169_,
		_w19170_
	);
	LUT2 #(
		.INIT('h1)
	) name18639 (
		_w16269_,
		_w16774_,
		_w19171_
	);
	LUT2 #(
		.INIT('h1)
	) name18640 (
		\u0_w_reg[3][19]/P0001 ,
		_w19171_,
		_w19172_
	);
	LUT2 #(
		.INIT('h1)
	) name18641 (
		_w15538_,
		_w15657_,
		_w19173_
	);
	LUT2 #(
		.INIT('h4)
	) name18642 (
		_w16222_,
		_w19173_,
		_w19174_
	);
	LUT2 #(
		.INIT('h4)
	) name18643 (
		_w19172_,
		_w19174_,
		_w19175_
	);
	LUT2 #(
		.INIT('h2)
	) name18644 (
		\u0_w_reg[3][18]/P0001 ,
		_w19175_,
		_w19176_
	);
	LUT2 #(
		.INIT('h8)
	) name18645 (
		\u0_w_reg[3][21]/P0001 ,
		_w15637_,
		_w19177_
	);
	LUT2 #(
		.INIT('h2)
	) name18646 (
		\u0_w_reg[3][22]/P0001 ,
		_w15613_,
		_w19178_
	);
	LUT2 #(
		.INIT('h8)
	) name18647 (
		_w15660_,
		_w19178_,
		_w19179_
	);
	LUT2 #(
		.INIT('h1)
	) name18648 (
		_w15650_,
		_w18490_,
		_w19180_
	);
	LUT2 #(
		.INIT('h1)
	) name18649 (
		_w19177_,
		_w19179_,
		_w19181_
	);
	LUT2 #(
		.INIT('h8)
	) name18650 (
		_w19180_,
		_w19181_,
		_w19182_
	);
	LUT2 #(
		.INIT('h4)
	) name18651 (
		_w19176_,
		_w19182_,
		_w19183_
	);
	LUT2 #(
		.INIT('h1)
	) name18652 (
		\u0_w_reg[3][17]/P0001 ,
		_w19183_,
		_w19184_
	);
	LUT2 #(
		.INIT('h4)
	) name18653 (
		_w15504_,
		_w17020_,
		_w19185_
	);
	LUT2 #(
		.INIT('h1)
	) name18654 (
		_w16269_,
		_w19185_,
		_w19186_
	);
	LUT2 #(
		.INIT('h1)
	) name18655 (
		\u0_w_reg[3][18]/P0001 ,
		_w19186_,
		_w19187_
	);
	LUT2 #(
		.INIT('h8)
	) name18656 (
		_w15511_,
		_w15602_,
		_w19188_
	);
	LUT2 #(
		.INIT('h2)
	) name18657 (
		\u0_w_reg[3][17]/P0001 ,
		_w16287_,
		_w19189_
	);
	LUT2 #(
		.INIT('h4)
	) name18658 (
		_w16777_,
		_w19189_,
		_w19190_
	);
	LUT2 #(
		.INIT('h4)
	) name18659 (
		_w19188_,
		_w19190_,
		_w19191_
	);
	LUT2 #(
		.INIT('h4)
	) name18660 (
		_w19187_,
		_w19191_,
		_w19192_
	);
	LUT2 #(
		.INIT('h8)
	) name18661 (
		\u0_w_reg[3][18]/P0001 ,
		_w15513_,
		_w19193_
	);
	LUT2 #(
		.INIT('h8)
	) name18662 (
		_w15504_,
		_w15520_,
		_w19194_
	);
	LUT2 #(
		.INIT('h4)
	) name18663 (
		\u0_w_reg[3][18]/P0001 ,
		_w16814_,
		_w19195_
	);
	LUT2 #(
		.INIT('h1)
	) name18664 (
		_w19193_,
		_w19194_,
		_w19196_
	);
	LUT2 #(
		.INIT('h8)
	) name18665 (
		_w17065_,
		_w19196_,
		_w19197_
	);
	LUT2 #(
		.INIT('h4)
	) name18666 (
		_w19195_,
		_w19197_,
		_w19198_
	);
	LUT2 #(
		.INIT('h1)
	) name18667 (
		_w19192_,
		_w19198_,
		_w19199_
	);
	LUT2 #(
		.INIT('h4)
	) name18668 (
		\u0_w_reg[3][19]/P0001 ,
		_w15519_,
		_w19200_
	);
	LUT2 #(
		.INIT('h1)
	) name18669 (
		_w17080_,
		_w19200_,
		_w19201_
	);
	LUT2 #(
		.INIT('h2)
	) name18670 (
		\u0_w_reg[3][18]/P0001 ,
		_w19201_,
		_w19202_
	);
	LUT2 #(
		.INIT('h1)
	) name18671 (
		_w15647_,
		_w16853_,
		_w19203_
	);
	LUT2 #(
		.INIT('h1)
	) name18672 (
		\u0_w_reg[3][19]/P0001 ,
		_w19203_,
		_w19204_
	);
	LUT2 #(
		.INIT('h1)
	) name18673 (
		_w19202_,
		_w19204_,
		_w19205_
	);
	LUT2 #(
		.INIT('h4)
	) name18674 (
		_w19199_,
		_w19205_,
		_w19206_
	);
	LUT2 #(
		.INIT('h1)
	) name18675 (
		\u0_w_reg[3][16]/P0001 ,
		_w19206_,
		_w19207_
	);
	LUT2 #(
		.INIT('h4)
	) name18676 (
		\u0_w_reg[3][18]/P0001 ,
		_w16283_,
		_w19208_
	);
	LUT2 #(
		.INIT('h1)
	) name18677 (
		_w19193_,
		_w19208_,
		_w19209_
	);
	LUT2 #(
		.INIT('h2)
	) name18678 (
		\u0_w_reg[3][19]/P0001 ,
		_w19209_,
		_w19210_
	);
	LUT2 #(
		.INIT('h8)
	) name18679 (
		\u0_w_reg[3][20]/P0001 ,
		_w16917_,
		_w19211_
	);
	LUT2 #(
		.INIT('h4)
	) name18680 (
		_w15520_,
		_w15529_,
		_w19212_
	);
	LUT2 #(
		.INIT('h1)
	) name18681 (
		_w15556_,
		_w19212_,
		_w19213_
	);
	LUT2 #(
		.INIT('h1)
	) name18682 (
		\u0_w_reg[3][21]/P0001 ,
		_w19213_,
		_w19214_
	);
	LUT2 #(
		.INIT('h1)
	) name18683 (
		_w15630_,
		_w16313_,
		_w19215_
	);
	LUT2 #(
		.INIT('h2)
	) name18684 (
		_w15648_,
		_w19215_,
		_w19216_
	);
	LUT2 #(
		.INIT('h1)
	) name18685 (
		_w17003_,
		_w17083_,
		_w19217_
	);
	LUT2 #(
		.INIT('h4)
	) name18686 (
		_w19211_,
		_w19217_,
		_w19218_
	);
	LUT2 #(
		.INIT('h1)
	) name18687 (
		_w19214_,
		_w19216_,
		_w19219_
	);
	LUT2 #(
		.INIT('h8)
	) name18688 (
		_w19218_,
		_w19219_,
		_w19220_
	);
	LUT2 #(
		.INIT('h2)
	) name18689 (
		\u0_w_reg[3][17]/P0001 ,
		_w19220_,
		_w19221_
	);
	LUT2 #(
		.INIT('h1)
	) name18690 (
		_w19210_,
		_w19221_,
		_w19222_
	);
	LUT2 #(
		.INIT('h4)
	) name18691 (
		_w19184_,
		_w19222_,
		_w19223_
	);
	LUT2 #(
		.INIT('h4)
	) name18692 (
		_w19207_,
		_w19223_,
		_w19224_
	);
	LUT2 #(
		.INIT('h4)
	) name18693 (
		_w19170_,
		_w19224_,
		_w19225_
	);
	LUT2 #(
		.INIT('h4)
	) name18694 (
		\u0_r0_out_reg[28]/P0001 ,
		_w19225_,
		_w19226_
	);
	LUT2 #(
		.INIT('h2)
	) name18695 (
		\u0_r0_out_reg[28]/P0001 ,
		_w19225_,
		_w19227_
	);
	LUT2 #(
		.INIT('h1)
	) name18696 (
		_w19226_,
		_w19227_,
		_w19228_
	);
	LUT2 #(
		.INIT('h8)
	) name18697 (
		\u0_w_reg[0][28]/P0001 ,
		_w19228_,
		_w19229_
	);
	LUT2 #(
		.INIT('h1)
	) name18698 (
		\u0_w_reg[0][28]/P0001 ,
		_w19228_,
		_w19230_
	);
	LUT2 #(
		.INIT('h1)
	) name18699 (
		_w19229_,
		_w19230_,
		_w19231_
	);
	LUT2 #(
		.INIT('h4)
	) name18700 (
		ld_pad,
		_w19231_,
		_w19232_
	);
	LUT2 #(
		.INIT('h8)
	) name18701 (
		\key[124]_pad ,
		ld_pad,
		_w19233_
	);
	LUT2 #(
		.INIT('h1)
	) name18702 (
		_w19232_,
		_w19233_,
		_w19234_
	);
	LUT2 #(
		.INIT('h1)
	) name18703 (
		\u0_w_reg[1][28]/P0001 ,
		_w19231_,
		_w19235_
	);
	LUT2 #(
		.INIT('h8)
	) name18704 (
		\u0_w_reg[1][28]/P0001 ,
		_w19231_,
		_w19236_
	);
	LUT2 #(
		.INIT('h1)
	) name18705 (
		ld_pad,
		_w19235_,
		_w19237_
	);
	LUT2 #(
		.INIT('h4)
	) name18706 (
		_w19236_,
		_w19237_,
		_w19238_
	);
	LUT2 #(
		.INIT('h8)
	) name18707 (
		\key[92]_pad ,
		ld_pad,
		_w19239_
	);
	LUT2 #(
		.INIT('h1)
	) name18708 (
		_w19238_,
		_w19239_,
		_w19240_
	);
	LUT2 #(
		.INIT('h2)
	) name18709 (
		\u0_w_reg[0][28]/P0001 ,
		\u0_w_reg[2][28]/P0001 ,
		_w19241_
	);
	LUT2 #(
		.INIT('h4)
	) name18710 (
		\u0_w_reg[0][28]/P0001 ,
		\u0_w_reg[2][28]/P0001 ,
		_w19242_
	);
	LUT2 #(
		.INIT('h1)
	) name18711 (
		_w19241_,
		_w19242_,
		_w19243_
	);
	LUT2 #(
		.INIT('h8)
	) name18712 (
		_w19228_,
		_w19243_,
		_w19244_
	);
	LUT2 #(
		.INIT('h1)
	) name18713 (
		_w19228_,
		_w19243_,
		_w19245_
	);
	LUT2 #(
		.INIT('h1)
	) name18714 (
		_w19244_,
		_w19245_,
		_w19246_
	);
	LUT2 #(
		.INIT('h4)
	) name18715 (
		\u0_w_reg[1][28]/P0001 ,
		_w19246_,
		_w19247_
	);
	LUT2 #(
		.INIT('h2)
	) name18716 (
		\u0_w_reg[1][28]/P0001 ,
		_w19246_,
		_w19248_
	);
	LUT2 #(
		.INIT('h1)
	) name18717 (
		ld_pad,
		_w19247_,
		_w19249_
	);
	LUT2 #(
		.INIT('h4)
	) name18718 (
		_w19248_,
		_w19249_,
		_w19250_
	);
	LUT2 #(
		.INIT('h8)
	) name18719 (
		\key[60]_pad ,
		ld_pad,
		_w19251_
	);
	LUT2 #(
		.INIT('h1)
	) name18720 (
		_w19250_,
		_w19251_,
		_w19252_
	);
	LUT2 #(
		.INIT('h8)
	) name18721 (
		\key[28]_pad ,
		ld_pad,
		_w19253_
	);
	LUT2 #(
		.INIT('h2)
	) name18722 (
		\u0_w_reg[1][28]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w19254_
	);
	LUT2 #(
		.INIT('h4)
	) name18723 (
		\u0_w_reg[1][28]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w19255_
	);
	LUT2 #(
		.INIT('h1)
	) name18724 (
		_w19254_,
		_w19255_,
		_w19256_
	);
	LUT2 #(
		.INIT('h8)
	) name18725 (
		_w19246_,
		_w19256_,
		_w19257_
	);
	LUT2 #(
		.INIT('h1)
	) name18726 (
		_w19246_,
		_w19256_,
		_w19258_
	);
	LUT2 #(
		.INIT('h1)
	) name18727 (
		ld_pad,
		_w19257_,
		_w19259_
	);
	LUT2 #(
		.INIT('h4)
	) name18728 (
		_w19258_,
		_w19259_,
		_w19260_
	);
	LUT2 #(
		.INIT('h1)
	) name18729 (
		_w19253_,
		_w19260_,
		_w19261_
	);
	LUT2 #(
		.INIT('h4)
	) name18730 (
		ld_pad,
		_w17361_,
		_w19262_
	);
	LUT2 #(
		.INIT('h8)
	) name18731 (
		\key[103]_pad ,
		ld_pad,
		_w19263_
	);
	LUT2 #(
		.INIT('h1)
	) name18732 (
		_w19262_,
		_w19263_,
		_w19264_
	);
	LUT2 #(
		.INIT('h1)
	) name18733 (
		\u0_w_reg[1][7]/P0001 ,
		_w17361_,
		_w19265_
	);
	LUT2 #(
		.INIT('h8)
	) name18734 (
		\u0_w_reg[1][7]/P0001 ,
		_w17361_,
		_w19266_
	);
	LUT2 #(
		.INIT('h1)
	) name18735 (
		ld_pad,
		_w19265_,
		_w19267_
	);
	LUT2 #(
		.INIT('h4)
	) name18736 (
		_w19266_,
		_w19267_,
		_w19268_
	);
	LUT2 #(
		.INIT('h8)
	) name18737 (
		\key[71]_pad ,
		ld_pad,
		_w19269_
	);
	LUT2 #(
		.INIT('h1)
	) name18738 (
		_w19268_,
		_w19269_,
		_w19270_
	);
	LUT2 #(
		.INIT('h4)
	) name18739 (
		\u0_w_reg[3][7]/P0001 ,
		_w17367_,
		_w19271_
	);
	LUT2 #(
		.INIT('h2)
	) name18740 (
		\u0_w_reg[3][7]/P0001 ,
		_w17367_,
		_w19272_
	);
	LUT2 #(
		.INIT('h1)
	) name18741 (
		ld_pad,
		_w19271_,
		_w19273_
	);
	LUT2 #(
		.INIT('h4)
	) name18742 (
		_w19272_,
		_w19273_,
		_w19274_
	);
	LUT2 #(
		.INIT('h8)
	) name18743 (
		\key[7]_pad ,
		ld_pad,
		_w19275_
	);
	LUT2 #(
		.INIT('h1)
	) name18744 (
		_w19274_,
		_w19275_,
		_w19276_
	);
	LUT2 #(
		.INIT('h4)
	) name18745 (
		ld_pad,
		_w17486_,
		_w19277_
	);
	LUT2 #(
		.INIT('h8)
	) name18746 (
		\key[96]_pad ,
		ld_pad,
		_w19278_
	);
	LUT2 #(
		.INIT('h1)
	) name18747 (
		_w19277_,
		_w19278_,
		_w19279_
	);
	LUT2 #(
		.INIT('h4)
	) name18748 (
		ld_pad,
		_w17588_,
		_w19280_
	);
	LUT2 #(
		.INIT('h8)
	) name18749 (
		\key[106]_pad ,
		ld_pad,
		_w19281_
	);
	LUT2 #(
		.INIT('h1)
	) name18750 (
		_w19280_,
		_w19281_,
		_w19282_
	);
	LUT2 #(
		.INIT('h4)
	) name18751 (
		ld_pad,
		_w17696_,
		_w19283_
	);
	LUT2 #(
		.INIT('h8)
	) name18752 (
		\key[112]_pad ,
		ld_pad,
		_w19284_
	);
	LUT2 #(
		.INIT('h1)
	) name18753 (
		_w19283_,
		_w19284_,
		_w19285_
	);
	LUT2 #(
		.INIT('h4)
	) name18754 (
		ld_pad,
		_w17793_,
		_w19286_
	);
	LUT2 #(
		.INIT('h8)
	) name18755 (
		\key[114]_pad ,
		ld_pad,
		_w19287_
	);
	LUT2 #(
		.INIT('h1)
	) name18756 (
		_w19286_,
		_w19287_,
		_w19288_
	);
	LUT2 #(
		.INIT('h4)
	) name18757 (
		ld_pad,
		_w17885_,
		_w19289_
	);
	LUT2 #(
		.INIT('h8)
	) name18758 (
		\key[98]_pad ,
		ld_pad,
		_w19290_
	);
	LUT2 #(
		.INIT('h1)
	) name18759 (
		_w19289_,
		_w19290_,
		_w19291_
	);
	LUT2 #(
		.INIT('h1)
	) name18760 (
		\u0_w_reg[1][0]/P0001 ,
		_w17486_,
		_w19292_
	);
	LUT2 #(
		.INIT('h8)
	) name18761 (
		\u0_w_reg[1][0]/P0001 ,
		_w17486_,
		_w19293_
	);
	LUT2 #(
		.INIT('h1)
	) name18762 (
		ld_pad,
		_w19292_,
		_w19294_
	);
	LUT2 #(
		.INIT('h4)
	) name18763 (
		_w19293_,
		_w19294_,
		_w19295_
	);
	LUT2 #(
		.INIT('h8)
	) name18764 (
		\key[64]_pad ,
		ld_pad,
		_w19296_
	);
	LUT2 #(
		.INIT('h1)
	) name18765 (
		_w19295_,
		_w19296_,
		_w19297_
	);
	LUT2 #(
		.INIT('h1)
	) name18766 (
		\u0_w_reg[1][10]/P0001 ,
		_w17588_,
		_w19298_
	);
	LUT2 #(
		.INIT('h8)
	) name18767 (
		\u0_w_reg[1][10]/P0001 ,
		_w17588_,
		_w19299_
	);
	LUT2 #(
		.INIT('h1)
	) name18768 (
		ld_pad,
		_w19298_,
		_w19300_
	);
	LUT2 #(
		.INIT('h4)
	) name18769 (
		_w19299_,
		_w19300_,
		_w19301_
	);
	LUT2 #(
		.INIT('h8)
	) name18770 (
		\key[74]_pad ,
		ld_pad,
		_w19302_
	);
	LUT2 #(
		.INIT('h1)
	) name18771 (
		_w19301_,
		_w19302_,
		_w19303_
	);
	LUT2 #(
		.INIT('h1)
	) name18772 (
		\u0_w_reg[1][16]/P0001 ,
		_w17696_,
		_w19304_
	);
	LUT2 #(
		.INIT('h8)
	) name18773 (
		\u0_w_reg[1][16]/P0001 ,
		_w17696_,
		_w19305_
	);
	LUT2 #(
		.INIT('h1)
	) name18774 (
		ld_pad,
		_w19304_,
		_w19306_
	);
	LUT2 #(
		.INIT('h4)
	) name18775 (
		_w19305_,
		_w19306_,
		_w19307_
	);
	LUT2 #(
		.INIT('h8)
	) name18776 (
		\key[80]_pad ,
		ld_pad,
		_w19308_
	);
	LUT2 #(
		.INIT('h1)
	) name18777 (
		_w19307_,
		_w19308_,
		_w19309_
	);
	LUT2 #(
		.INIT('h1)
	) name18778 (
		\u0_w_reg[1][18]/P0001 ,
		_w17793_,
		_w19310_
	);
	LUT2 #(
		.INIT('h8)
	) name18779 (
		\u0_w_reg[1][18]/P0001 ,
		_w17793_,
		_w19311_
	);
	LUT2 #(
		.INIT('h1)
	) name18780 (
		ld_pad,
		_w19310_,
		_w19312_
	);
	LUT2 #(
		.INIT('h4)
	) name18781 (
		_w19311_,
		_w19312_,
		_w19313_
	);
	LUT2 #(
		.INIT('h8)
	) name18782 (
		\key[82]_pad ,
		ld_pad,
		_w19314_
	);
	LUT2 #(
		.INIT('h1)
	) name18783 (
		_w19313_,
		_w19314_,
		_w19315_
	);
	LUT2 #(
		.INIT('h4)
	) name18784 (
		ld_pad,
		_w17888_,
		_w19316_
	);
	LUT2 #(
		.INIT('h8)
	) name18785 (
		\key[66]_pad ,
		ld_pad,
		_w19317_
	);
	LUT2 #(
		.INIT('h1)
	) name18786 (
		_w19316_,
		_w19317_,
		_w19318_
	);
	LUT2 #(
		.INIT('h4)
	) name18787 (
		\u0_w_reg[3][0]/P0001 ,
		_w17492_,
		_w19319_
	);
	LUT2 #(
		.INIT('h2)
	) name18788 (
		\u0_w_reg[3][0]/P0001 ,
		_w17492_,
		_w19320_
	);
	LUT2 #(
		.INIT('h1)
	) name18789 (
		ld_pad,
		_w19319_,
		_w19321_
	);
	LUT2 #(
		.INIT('h4)
	) name18790 (
		_w19320_,
		_w19321_,
		_w19322_
	);
	LUT2 #(
		.INIT('h8)
	) name18791 (
		\key[0]_pad ,
		ld_pad,
		_w19323_
	);
	LUT2 #(
		.INIT('h1)
	) name18792 (
		_w19322_,
		_w19323_,
		_w19324_
	);
	LUT2 #(
		.INIT('h4)
	) name18793 (
		\u0_w_reg[3][10]/P0001 ,
		_w17594_,
		_w19325_
	);
	LUT2 #(
		.INIT('h2)
	) name18794 (
		\u0_w_reg[3][10]/P0001 ,
		_w17594_,
		_w19326_
	);
	LUT2 #(
		.INIT('h1)
	) name18795 (
		ld_pad,
		_w19325_,
		_w19327_
	);
	LUT2 #(
		.INIT('h4)
	) name18796 (
		_w19326_,
		_w19327_,
		_w19328_
	);
	LUT2 #(
		.INIT('h8)
	) name18797 (
		\key[10]_pad ,
		ld_pad,
		_w19329_
	);
	LUT2 #(
		.INIT('h1)
	) name18798 (
		_w19328_,
		_w19329_,
		_w19330_
	);
	LUT2 #(
		.INIT('h4)
	) name18799 (
		\u0_w_reg[3][16]/P0001 ,
		_w17702_,
		_w19331_
	);
	LUT2 #(
		.INIT('h2)
	) name18800 (
		\u0_w_reg[3][16]/P0001 ,
		_w17702_,
		_w19332_
	);
	LUT2 #(
		.INIT('h1)
	) name18801 (
		ld_pad,
		_w19331_,
		_w19333_
	);
	LUT2 #(
		.INIT('h4)
	) name18802 (
		_w19332_,
		_w19333_,
		_w19334_
	);
	LUT2 #(
		.INIT('h8)
	) name18803 (
		\key[16]_pad ,
		ld_pad,
		_w19335_
	);
	LUT2 #(
		.INIT('h1)
	) name18804 (
		_w19334_,
		_w19335_,
		_w19336_
	);
	LUT2 #(
		.INIT('h4)
	) name18805 (
		\u0_w_reg[3][18]/P0001 ,
		_w17799_,
		_w19337_
	);
	LUT2 #(
		.INIT('h2)
	) name18806 (
		\u0_w_reg[3][18]/P0001 ,
		_w17799_,
		_w19338_
	);
	LUT2 #(
		.INIT('h1)
	) name18807 (
		ld_pad,
		_w19337_,
		_w19339_
	);
	LUT2 #(
		.INIT('h4)
	) name18808 (
		_w19338_,
		_w19339_,
		_w19340_
	);
	LUT2 #(
		.INIT('h8)
	) name18809 (
		\key[18]_pad ,
		ld_pad,
		_w19341_
	);
	LUT2 #(
		.INIT('h1)
	) name18810 (
		_w19340_,
		_w19341_,
		_w19342_
	);
	LUT2 #(
		.INIT('h1)
	) name18811 (
		\u0_w_reg[3][2]/P0001 ,
		_w17891_,
		_w19343_
	);
	LUT2 #(
		.INIT('h8)
	) name18812 (
		\u0_w_reg[3][2]/P0001 ,
		_w17891_,
		_w19344_
	);
	LUT2 #(
		.INIT('h1)
	) name18813 (
		ld_pad,
		_w19343_,
		_w19345_
	);
	LUT2 #(
		.INIT('h4)
	) name18814 (
		_w19344_,
		_w19345_,
		_w19346_
	);
	LUT2 #(
		.INIT('h8)
	) name18815 (
		\key[2]_pad ,
		ld_pad,
		_w19347_
	);
	LUT2 #(
		.INIT('h1)
	) name18816 (
		_w19346_,
		_w19347_,
		_w19348_
	);
	LUT2 #(
		.INIT('h1)
	) name18817 (
		\u0_w_reg[0][5]/P0001 ,
		_w12580_,
		_w19349_
	);
	LUT2 #(
		.INIT('h8)
	) name18818 (
		\u0_w_reg[0][5]/P0001 ,
		_w12580_,
		_w19350_
	);
	LUT2 #(
		.INIT('h1)
	) name18819 (
		_w19349_,
		_w19350_,
		_w19351_
	);
	LUT2 #(
		.INIT('h4)
	) name18820 (
		ld_pad,
		_w17983_,
		_w19352_
	);
	LUT2 #(
		.INIT('h8)
	) name18821 (
		\key[110]_pad ,
		ld_pad,
		_w19353_
	);
	LUT2 #(
		.INIT('h1)
	) name18822 (
		_w19352_,
		_w19353_,
		_w19354_
	);
	LUT2 #(
		.INIT('h4)
	) name18823 (
		ld_pad,
		_w18069_,
		_w19355_
	);
	LUT2 #(
		.INIT('h8)
	) name18824 (
		\key[118]_pad ,
		ld_pad,
		_w19356_
	);
	LUT2 #(
		.INIT('h1)
	) name18825 (
		_w19355_,
		_w19356_,
		_w19357_
	);
	LUT2 #(
		.INIT('h4)
	) name18826 (
		ld_pad,
		_w18153_,
		_w19358_
	);
	LUT2 #(
		.INIT('h8)
	) name18827 (
		\key[102]_pad ,
		ld_pad,
		_w19359_
	);
	LUT2 #(
		.INIT('h1)
	) name18828 (
		_w19358_,
		_w19359_,
		_w19360_
	);
	LUT2 #(
		.INIT('h1)
	) name18829 (
		\u0_w_reg[1][14]/P0001 ,
		_w17983_,
		_w19361_
	);
	LUT2 #(
		.INIT('h8)
	) name18830 (
		\u0_w_reg[1][14]/P0001 ,
		_w17983_,
		_w19362_
	);
	LUT2 #(
		.INIT('h1)
	) name18831 (
		ld_pad,
		_w19361_,
		_w19363_
	);
	LUT2 #(
		.INIT('h4)
	) name18832 (
		_w19362_,
		_w19363_,
		_w19364_
	);
	LUT2 #(
		.INIT('h8)
	) name18833 (
		\key[78]_pad ,
		ld_pad,
		_w19365_
	);
	LUT2 #(
		.INIT('h1)
	) name18834 (
		_w19364_,
		_w19365_,
		_w19366_
	);
	LUT2 #(
		.INIT('h1)
	) name18835 (
		\u0_w_reg[1][22]/P0001 ,
		_w18069_,
		_w19367_
	);
	LUT2 #(
		.INIT('h8)
	) name18836 (
		\u0_w_reg[1][22]/P0001 ,
		_w18069_,
		_w19368_
	);
	LUT2 #(
		.INIT('h1)
	) name18837 (
		ld_pad,
		_w19367_,
		_w19369_
	);
	LUT2 #(
		.INIT('h4)
	) name18838 (
		_w19368_,
		_w19369_,
		_w19370_
	);
	LUT2 #(
		.INIT('h8)
	) name18839 (
		\key[86]_pad ,
		ld_pad,
		_w19371_
	);
	LUT2 #(
		.INIT('h1)
	) name18840 (
		_w19370_,
		_w19371_,
		_w19372_
	);
	LUT2 #(
		.INIT('h1)
	) name18841 (
		\u0_w_reg[1][6]/P0001 ,
		_w18153_,
		_w19373_
	);
	LUT2 #(
		.INIT('h8)
	) name18842 (
		\u0_w_reg[1][6]/P0001 ,
		_w18153_,
		_w19374_
	);
	LUT2 #(
		.INIT('h1)
	) name18843 (
		ld_pad,
		_w19373_,
		_w19375_
	);
	LUT2 #(
		.INIT('h4)
	) name18844 (
		_w19374_,
		_w19375_,
		_w19376_
	);
	LUT2 #(
		.INIT('h8)
	) name18845 (
		\key[70]_pad ,
		ld_pad,
		_w19377_
	);
	LUT2 #(
		.INIT('h1)
	) name18846 (
		_w19376_,
		_w19377_,
		_w19378_
	);
	LUT2 #(
		.INIT('h4)
	) name18847 (
		\u0_w_reg[3][14]/P0001 ,
		_w17989_,
		_w19379_
	);
	LUT2 #(
		.INIT('h2)
	) name18848 (
		\u0_w_reg[3][14]/P0001 ,
		_w17989_,
		_w19380_
	);
	LUT2 #(
		.INIT('h1)
	) name18849 (
		ld_pad,
		_w19379_,
		_w19381_
	);
	LUT2 #(
		.INIT('h4)
	) name18850 (
		_w19380_,
		_w19381_,
		_w19382_
	);
	LUT2 #(
		.INIT('h8)
	) name18851 (
		\key[14]_pad ,
		ld_pad,
		_w19383_
	);
	LUT2 #(
		.INIT('h1)
	) name18852 (
		_w19382_,
		_w19383_,
		_w19384_
	);
	LUT2 #(
		.INIT('h4)
	) name18853 (
		\u0_w_reg[3][22]/P0001 ,
		_w18075_,
		_w19385_
	);
	LUT2 #(
		.INIT('h2)
	) name18854 (
		\u0_w_reg[3][22]/P0001 ,
		_w18075_,
		_w19386_
	);
	LUT2 #(
		.INIT('h1)
	) name18855 (
		ld_pad,
		_w19385_,
		_w19387_
	);
	LUT2 #(
		.INIT('h4)
	) name18856 (
		_w19386_,
		_w19387_,
		_w19388_
	);
	LUT2 #(
		.INIT('h8)
	) name18857 (
		\key[22]_pad ,
		ld_pad,
		_w19389_
	);
	LUT2 #(
		.INIT('h1)
	) name18858 (
		_w19388_,
		_w19389_,
		_w19390_
	);
	LUT2 #(
		.INIT('h4)
	) name18859 (
		\u0_w_reg[3][6]/P0001 ,
		_w18159_,
		_w19391_
	);
	LUT2 #(
		.INIT('h2)
	) name18860 (
		\u0_w_reg[3][6]/P0001 ,
		_w18159_,
		_w19392_
	);
	LUT2 #(
		.INIT('h1)
	) name18861 (
		ld_pad,
		_w19391_,
		_w19393_
	);
	LUT2 #(
		.INIT('h4)
	) name18862 (
		_w19392_,
		_w19393_,
		_w19394_
	);
	LUT2 #(
		.INIT('h8)
	) name18863 (
		\key[6]_pad ,
		ld_pad,
		_w19395_
	);
	LUT2 #(
		.INIT('h1)
	) name18864 (
		_w19394_,
		_w19395_,
		_w19396_
	);
	LUT2 #(
		.INIT('h4)
	) name18865 (
		ld_pad,
		_w18255_,
		_w19397_
	);
	LUT2 #(
		.INIT('h8)
	) name18866 (
		\key[109]_pad ,
		ld_pad,
		_w19398_
	);
	LUT2 #(
		.INIT('h1)
	) name18867 (
		_w19397_,
		_w19398_,
		_w19399_
	);
	LUT2 #(
		.INIT('h4)
	) name18868 (
		ld_pad,
		_w18355_,
		_w19400_
	);
	LUT2 #(
		.INIT('h8)
	) name18869 (
		\key[111]_pad ,
		ld_pad,
		_w19401_
	);
	LUT2 #(
		.INIT('h1)
	) name18870 (
		_w19400_,
		_w19401_,
		_w19402_
	);
	LUT2 #(
		.INIT('h4)
	) name18871 (
		ld_pad,
		_w18437_,
		_w19403_
	);
	LUT2 #(
		.INIT('h8)
	) name18872 (
		\key[104]_pad ,
		ld_pad,
		_w19404_
	);
	LUT2 #(
		.INIT('h1)
	) name18873 (
		_w19403_,
		_w19404_,
		_w19405_
	);
	LUT2 #(
		.INIT('h1)
	) name18874 (
		\u0_w_reg[1][13]/P0001 ,
		_w18255_,
		_w19406_
	);
	LUT2 #(
		.INIT('h8)
	) name18875 (
		\u0_w_reg[1][13]/P0001 ,
		_w18255_,
		_w19407_
	);
	LUT2 #(
		.INIT('h1)
	) name18876 (
		ld_pad,
		_w19406_,
		_w19408_
	);
	LUT2 #(
		.INIT('h4)
	) name18877 (
		_w19407_,
		_w19408_,
		_w19409_
	);
	LUT2 #(
		.INIT('h8)
	) name18878 (
		\key[77]_pad ,
		ld_pad,
		_w19410_
	);
	LUT2 #(
		.INIT('h1)
	) name18879 (
		_w19409_,
		_w19410_,
		_w19411_
	);
	LUT2 #(
		.INIT('h4)
	) name18880 (
		ld_pad,
		_w18358_,
		_w19412_
	);
	LUT2 #(
		.INIT('h8)
	) name18881 (
		\key[79]_pad ,
		ld_pad,
		_w19413_
	);
	LUT2 #(
		.INIT('h1)
	) name18882 (
		_w19412_,
		_w19413_,
		_w19414_
	);
	LUT2 #(
		.INIT('h1)
	) name18883 (
		\u0_w_reg[1][8]/P0001 ,
		_w18437_,
		_w19415_
	);
	LUT2 #(
		.INIT('h8)
	) name18884 (
		\u0_w_reg[1][8]/P0001 ,
		_w18437_,
		_w19416_
	);
	LUT2 #(
		.INIT('h1)
	) name18885 (
		ld_pad,
		_w19415_,
		_w19417_
	);
	LUT2 #(
		.INIT('h4)
	) name18886 (
		_w19416_,
		_w19417_,
		_w19418_
	);
	LUT2 #(
		.INIT('h8)
	) name18887 (
		\key[72]_pad ,
		ld_pad,
		_w19419_
	);
	LUT2 #(
		.INIT('h1)
	) name18888 (
		_w19418_,
		_w19419_,
		_w19420_
	);
	LUT2 #(
		.INIT('h4)
	) name18889 (
		\u0_w_reg[3][13]/P0001 ,
		_w18261_,
		_w19421_
	);
	LUT2 #(
		.INIT('h2)
	) name18890 (
		\u0_w_reg[3][13]/P0001 ,
		_w18261_,
		_w19422_
	);
	LUT2 #(
		.INIT('h1)
	) name18891 (
		ld_pad,
		_w19421_,
		_w19423_
	);
	LUT2 #(
		.INIT('h4)
	) name18892 (
		_w19422_,
		_w19423_,
		_w19424_
	);
	LUT2 #(
		.INIT('h8)
	) name18893 (
		\key[13]_pad ,
		ld_pad,
		_w19425_
	);
	LUT2 #(
		.INIT('h1)
	) name18894 (
		_w19424_,
		_w19425_,
		_w19426_
	);
	LUT2 #(
		.INIT('h1)
	) name18895 (
		\u0_w_reg[3][15]/P0001 ,
		_w18361_,
		_w19427_
	);
	LUT2 #(
		.INIT('h8)
	) name18896 (
		\u0_w_reg[3][15]/P0001 ,
		_w18361_,
		_w19428_
	);
	LUT2 #(
		.INIT('h1)
	) name18897 (
		ld_pad,
		_w19427_,
		_w19429_
	);
	LUT2 #(
		.INIT('h4)
	) name18898 (
		_w19428_,
		_w19429_,
		_w19430_
	);
	LUT2 #(
		.INIT('h8)
	) name18899 (
		\key[15]_pad ,
		ld_pad,
		_w19431_
	);
	LUT2 #(
		.INIT('h1)
	) name18900 (
		_w19430_,
		_w19431_,
		_w19432_
	);
	LUT2 #(
		.INIT('h4)
	) name18901 (
		\u0_w_reg[3][8]/P0001 ,
		_w18443_,
		_w19433_
	);
	LUT2 #(
		.INIT('h2)
	) name18902 (
		\u0_w_reg[3][8]/P0001 ,
		_w18443_,
		_w19434_
	);
	LUT2 #(
		.INIT('h1)
	) name18903 (
		ld_pad,
		_w19433_,
		_w19435_
	);
	LUT2 #(
		.INIT('h4)
	) name18904 (
		_w19434_,
		_w19435_,
		_w19436_
	);
	LUT2 #(
		.INIT('h8)
	) name18905 (
		\key[8]_pad ,
		ld_pad,
		_w19437_
	);
	LUT2 #(
		.INIT('h1)
	) name18906 (
		_w19436_,
		_w19437_,
		_w19438_
	);
	LUT2 #(
		.INIT('h1)
	) name18907 (
		\u0_w_reg[0][29]/P0001 ,
		_w12714_,
		_w19439_
	);
	LUT2 #(
		.INIT('h8)
	) name18908 (
		\u0_w_reg[0][29]/P0001 ,
		_w12714_,
		_w19440_
	);
	LUT2 #(
		.INIT('h1)
	) name18909 (
		_w19439_,
		_w19440_,
		_w19441_
	);
	LUT2 #(
		.INIT('h1)
	) name18910 (
		\u0_w_reg[3][29]/P0001 ,
		_w1479_,
		_w19442_
	);
	LUT2 #(
		.INIT('h8)
	) name18911 (
		\u0_w_reg[3][29]/P0001 ,
		_w1479_,
		_w19443_
	);
	LUT2 #(
		.INIT('h1)
	) name18912 (
		_w19442_,
		_w19443_,
		_w19444_
	);
	LUT2 #(
		.INIT('h1)
	) name18913 (
		\u0_w_reg[2][29]/P0001 ,
		_w1142_,
		_w19445_
	);
	LUT2 #(
		.INIT('h8)
	) name18914 (
		\u0_w_reg[2][29]/P0001 ,
		_w1142_,
		_w19446_
	);
	LUT2 #(
		.INIT('h1)
	) name18915 (
		_w19445_,
		_w19446_,
		_w19447_
	);
	LUT2 #(
		.INIT('h1)
	) name18916 (
		\u0_w_reg[1][29]/P0002 ,
		_w9289_,
		_w19448_
	);
	LUT2 #(
		.INIT('h8)
	) name18917 (
		\u0_w_reg[1][29]/P0002 ,
		_w9289_,
		_w19449_
	);
	LUT2 #(
		.INIT('h1)
	) name18918 (
		_w19448_,
		_w19449_,
		_w19450_
	);
	LUT2 #(
		.INIT('h4)
	) name18919 (
		ld_pad,
		_w18645_,
		_w19451_
	);
	LUT2 #(
		.INIT('h8)
	) name18920 (
		\key[119]_pad ,
		ld_pad,
		_w19452_
	);
	LUT2 #(
		.INIT('h1)
	) name18921 (
		_w19451_,
		_w19452_,
		_w19453_
	);
	LUT2 #(
		.INIT('h4)
	) name18922 (
		ld_pad,
		_w18648_,
		_w19454_
	);
	LUT2 #(
		.INIT('h8)
	) name18923 (
		\key[87]_pad ,
		ld_pad,
		_w19455_
	);
	LUT2 #(
		.INIT('h1)
	) name18924 (
		_w19454_,
		_w19455_,
		_w19456_
	);
	LUT2 #(
		.INIT('h1)
	) name18925 (
		\u0_w_reg[3][23]/P0001 ,
		_w18651_,
		_w19457_
	);
	LUT2 #(
		.INIT('h8)
	) name18926 (
		\u0_w_reg[3][23]/P0001 ,
		_w18651_,
		_w19458_
	);
	LUT2 #(
		.INIT('h1)
	) name18927 (
		ld_pad,
		_w19457_,
		_w19459_
	);
	LUT2 #(
		.INIT('h4)
	) name18928 (
		_w19458_,
		_w19459_,
		_w19460_
	);
	LUT2 #(
		.INIT('h8)
	) name18929 (
		\key[23]_pad ,
		ld_pad,
		_w19461_
	);
	LUT2 #(
		.INIT('h1)
	) name18930 (
		_w19460_,
		_w19461_,
		_w19462_
	);
	LUT2 #(
		.INIT('h1)
	) name18931 (
		\u0_w_reg[3][8]/P0001 ,
		_w3592_,
		_w19463_
	);
	LUT2 #(
		.INIT('h8)
	) name18932 (
		\u0_w_reg[3][8]/P0001 ,
		_w3592_,
		_w19464_
	);
	LUT2 #(
		.INIT('h1)
	) name18933 (
		_w19463_,
		_w19464_,
		_w19465_
	);
	LUT2 #(
		.INIT('h1)
	) name18934 (
		\u0_w_reg[0][11]/P0001 ,
		_w14567_,
		_w19466_
	);
	LUT2 #(
		.INIT('h8)
	) name18935 (
		\u0_w_reg[0][11]/P0001 ,
		_w14567_,
		_w19467_
	);
	LUT2 #(
		.INIT('h1)
	) name18936 (
		_w19466_,
		_w19467_,
		_w19468_
	);
	LUT2 #(
		.INIT('h1)
	) name18937 (
		\u0_w_reg[3][11]/P0001 ,
		_w4059_,
		_w19469_
	);
	LUT2 #(
		.INIT('h8)
	) name18938 (
		\u0_w_reg[3][11]/P0001 ,
		_w4059_,
		_w19470_
	);
	LUT2 #(
		.INIT('h1)
	) name18939 (
		_w19469_,
		_w19470_,
		_w19471_
	);
	LUT2 #(
		.INIT('h1)
	) name18940 (
		\u0_w_reg[2][11]/P0001 ,
		_w7206_,
		_w19472_
	);
	LUT2 #(
		.INIT('h8)
	) name18941 (
		\u0_w_reg[2][11]/P0001 ,
		_w7206_,
		_w19473_
	);
	LUT2 #(
		.INIT('h1)
	) name18942 (
		_w19472_,
		_w19473_,
		_w19474_
	);
	LUT2 #(
		.INIT('h1)
	) name18943 (
		\u0_w_reg[1][11]/P0001 ,
		_w10775_,
		_w19475_
	);
	LUT2 #(
		.INIT('h8)
	) name18944 (
		\u0_w_reg[1][11]/P0001 ,
		_w10775_,
		_w19476_
	);
	LUT2 #(
		.INIT('h1)
	) name18945 (
		_w19475_,
		_w19476_,
		_w19477_
	);
	LUT2 #(
		.INIT('h1)
	) name18946 (
		\u0_w_reg[0][12]/P0001 ,
		_w12827_,
		_w19478_
	);
	LUT2 #(
		.INIT('h8)
	) name18947 (
		\u0_w_reg[0][12]/P0001 ,
		_w12827_,
		_w19479_
	);
	LUT2 #(
		.INIT('h1)
	) name18948 (
		_w19478_,
		_w19479_,
		_w19480_
	);
	LUT2 #(
		.INIT('h1)
	) name18949 (
		\u0_w_reg[2][12]/P0001 ,
		_w6055_,
		_w19481_
	);
	LUT2 #(
		.INIT('h8)
	) name18950 (
		\u0_w_reg[2][12]/P0001 ,
		_w6055_,
		_w19482_
	);
	LUT2 #(
		.INIT('h1)
	) name18951 (
		_w19481_,
		_w19482_,
		_w19483_
	);
	LUT2 #(
		.INIT('h1)
	) name18952 (
		\u0_w_reg[1][12]/P0001 ,
		_w9516_,
		_w19484_
	);
	LUT2 #(
		.INIT('h8)
	) name18953 (
		\u0_w_reg[1][12]/P0001 ,
		_w9516_,
		_w19485_
	);
	LUT2 #(
		.INIT('h1)
	) name18954 (
		_w19484_,
		_w19485_,
		_w19486_
	);
	LUT2 #(
		.INIT('h1)
	) name18955 (
		\u0_w_reg[0][8]/P0001 ,
		_w13379_,
		_w19487_
	);
	LUT2 #(
		.INIT('h8)
	) name18956 (
		\u0_w_reg[0][8]/P0001 ,
		_w13379_,
		_w19488_
	);
	LUT2 #(
		.INIT('h1)
	) name18957 (
		_w19487_,
		_w19488_,
		_w19489_
	);
	LUT2 #(
		.INIT('h1)
	) name18958 (
		\u0_w_reg[0][24]/P0001 ,
		_w14316_,
		_w19490_
	);
	LUT2 #(
		.INIT('h8)
	) name18959 (
		\u0_w_reg[0][24]/P0001 ,
		_w14316_,
		_w19491_
	);
	LUT2 #(
		.INIT('h1)
	) name18960 (
		_w19490_,
		_w19491_,
		_w19492_
	);
	LUT2 #(
		.INIT('h1)
	) name18961 (
		\u0_w_reg[0][27]/P0001 ,
		_w14970_,
		_w19493_
	);
	LUT2 #(
		.INIT('h8)
	) name18962 (
		\u0_w_reg[0][27]/P0001 ,
		_w14970_,
		_w19494_
	);
	LUT2 #(
		.INIT('h1)
	) name18963 (
		_w19493_,
		_w19494_,
		_w19495_
	);
	LUT2 #(
		.INIT('h1)
	) name18964 (
		\u0_w_reg[3][24]/P0001 ,
		_w4161_,
		_w19496_
	);
	LUT2 #(
		.INIT('h8)
	) name18965 (
		\u0_w_reg[3][24]/P0001 ,
		_w4161_,
		_w19497_
	);
	LUT2 #(
		.INIT('h1)
	) name18966 (
		_w19496_,
		_w19497_,
		_w19498_
	);
	LUT2 #(
		.INIT('h1)
	) name18967 (
		\u0_w_reg[3][27]/P0001 ,
		_w3888_,
		_w19499_
	);
	LUT2 #(
		.INIT('h8)
	) name18968 (
		\u0_w_reg[3][27]/P0001 ,
		_w3888_,
		_w19500_
	);
	LUT2 #(
		.INIT('h1)
	) name18969 (
		_w19499_,
		_w19500_,
		_w19501_
	);
	LUT2 #(
		.INIT('h1)
	) name18970 (
		\u0_w_reg[2][8]/P0001 ,
		_w6927_,
		_w19502_
	);
	LUT2 #(
		.INIT('h8)
	) name18971 (
		\u0_w_reg[2][8]/P0001 ,
		_w6927_,
		_w19503_
	);
	LUT2 #(
		.INIT('h1)
	) name18972 (
		_w19502_,
		_w19503_,
		_w19504_
	);
	LUT2 #(
		.INIT('h1)
	) name18973 (
		\u0_w_reg[2][24]/P0001 ,
		_w6472_,
		_w19505_
	);
	LUT2 #(
		.INIT('h8)
	) name18974 (
		\u0_w_reg[2][24]/P0001 ,
		_w6472_,
		_w19506_
	);
	LUT2 #(
		.INIT('h1)
	) name18975 (
		_w19505_,
		_w19506_,
		_w19507_
	);
	LUT2 #(
		.INIT('h1)
	) name18976 (
		\u0_w_reg[2][27]/P0001 ,
		_w7040_,
		_w19508_
	);
	LUT2 #(
		.INIT('h8)
	) name18977 (
		\u0_w_reg[2][27]/P0001 ,
		_w7040_,
		_w19509_
	);
	LUT2 #(
		.INIT('h1)
	) name18978 (
		_w19508_,
		_w19509_,
		_w19510_
	);
	LUT2 #(
		.INIT('h1)
	) name18979 (
		\u0_w_reg[1][8]/P0001 ,
		_w11073_,
		_w19511_
	);
	LUT2 #(
		.INIT('h8)
	) name18980 (
		\u0_w_reg[1][8]/P0001 ,
		_w11073_,
		_w19512_
	);
	LUT2 #(
		.INIT('h1)
	) name18981 (
		_w19511_,
		_w19512_,
		_w19513_
	);
	LUT2 #(
		.INIT('h1)
	) name18982 (
		\u0_w_reg[1][24]/P0002 ,
		_w10248_,
		_w19514_
	);
	LUT2 #(
		.INIT('h8)
	) name18983 (
		\u0_w_reg[1][24]/P0002 ,
		_w10248_,
		_w19515_
	);
	LUT2 #(
		.INIT('h1)
	) name18984 (
		_w19514_,
		_w19515_,
		_w19516_
	);
	LUT2 #(
		.INIT('h1)
	) name18985 (
		\u0_w_reg[1][27]/P0001 ,
		_w10602_,
		_w19517_
	);
	LUT2 #(
		.INIT('h8)
	) name18986 (
		\u0_w_reg[1][27]/P0001 ,
		_w10602_,
		_w19518_
	);
	LUT2 #(
		.INIT('h1)
	) name18987 (
		_w19517_,
		_w19518_,
		_w19519_
	);
	LUT2 #(
		.INIT('h4)
	) name18988 (
		ld_pad,
		_w18765_,
		_w19520_
	);
	LUT2 #(
		.INIT('h8)
	) name18989 (
		\key[113]_pad ,
		ld_pad,
		_w19521_
	);
	LUT2 #(
		.INIT('h1)
	) name18990 (
		_w19520_,
		_w19521_,
		_w19522_
	);
	LUT2 #(
		.INIT('h4)
	) name18991 (
		ld_pad,
		_w18854_,
		_w19523_
	);
	LUT2 #(
		.INIT('h8)
	) name18992 (
		\key[97]_pad ,
		ld_pad,
		_w19524_
	);
	LUT2 #(
		.INIT('h1)
	) name18993 (
		_w19523_,
		_w19524_,
		_w19525_
	);
	LUT2 #(
		.INIT('h4)
	) name18994 (
		ld_pad,
		_w18945_,
		_w19526_
	);
	LUT2 #(
		.INIT('h8)
	) name18995 (
		\key[105]_pad ,
		ld_pad,
		_w19527_
	);
	LUT2 #(
		.INIT('h1)
	) name18996 (
		_w19526_,
		_w19527_,
		_w19528_
	);
	LUT2 #(
		.INIT('h1)
	) name18997 (
		\u0_w_reg[1][17]/P0001 ,
		_w18765_,
		_w19529_
	);
	LUT2 #(
		.INIT('h8)
	) name18998 (
		\u0_w_reg[1][17]/P0001 ,
		_w18765_,
		_w19530_
	);
	LUT2 #(
		.INIT('h1)
	) name18999 (
		ld_pad,
		_w19529_,
		_w19531_
	);
	LUT2 #(
		.INIT('h4)
	) name19000 (
		_w19530_,
		_w19531_,
		_w19532_
	);
	LUT2 #(
		.INIT('h8)
	) name19001 (
		\key[81]_pad ,
		ld_pad,
		_w19533_
	);
	LUT2 #(
		.INIT('h1)
	) name19002 (
		_w19532_,
		_w19533_,
		_w19534_
	);
	LUT2 #(
		.INIT('h1)
	) name19003 (
		\u0_w_reg[1][1]/P0001 ,
		_w18854_,
		_w19535_
	);
	LUT2 #(
		.INIT('h8)
	) name19004 (
		\u0_w_reg[1][1]/P0001 ,
		_w18854_,
		_w19536_
	);
	LUT2 #(
		.INIT('h1)
	) name19005 (
		ld_pad,
		_w19535_,
		_w19537_
	);
	LUT2 #(
		.INIT('h4)
	) name19006 (
		_w19536_,
		_w19537_,
		_w19538_
	);
	LUT2 #(
		.INIT('h8)
	) name19007 (
		\key[65]_pad ,
		ld_pad,
		_w19539_
	);
	LUT2 #(
		.INIT('h1)
	) name19008 (
		_w19538_,
		_w19539_,
		_w19540_
	);
	LUT2 #(
		.INIT('h1)
	) name19009 (
		\u0_w_reg[1][9]/P0001 ,
		_w18945_,
		_w19541_
	);
	LUT2 #(
		.INIT('h8)
	) name19010 (
		\u0_w_reg[1][9]/P0001 ,
		_w18945_,
		_w19542_
	);
	LUT2 #(
		.INIT('h1)
	) name19011 (
		ld_pad,
		_w19541_,
		_w19543_
	);
	LUT2 #(
		.INIT('h4)
	) name19012 (
		_w19542_,
		_w19543_,
		_w19544_
	);
	LUT2 #(
		.INIT('h8)
	) name19013 (
		\key[73]_pad ,
		ld_pad,
		_w19545_
	);
	LUT2 #(
		.INIT('h1)
	) name19014 (
		_w19544_,
		_w19545_,
		_w19546_
	);
	LUT2 #(
		.INIT('h4)
	) name19015 (
		\u0_w_reg[3][17]/P0001 ,
		_w18771_,
		_w19547_
	);
	LUT2 #(
		.INIT('h2)
	) name19016 (
		\u0_w_reg[3][17]/P0001 ,
		_w18771_,
		_w19548_
	);
	LUT2 #(
		.INIT('h1)
	) name19017 (
		ld_pad,
		_w19547_,
		_w19549_
	);
	LUT2 #(
		.INIT('h4)
	) name19018 (
		_w19548_,
		_w19549_,
		_w19550_
	);
	LUT2 #(
		.INIT('h8)
	) name19019 (
		\key[17]_pad ,
		ld_pad,
		_w19551_
	);
	LUT2 #(
		.INIT('h1)
	) name19020 (
		_w19550_,
		_w19551_,
		_w19552_
	);
	LUT2 #(
		.INIT('h4)
	) name19021 (
		\u0_w_reg[3][1]/P0001 ,
		_w18860_,
		_w19553_
	);
	LUT2 #(
		.INIT('h2)
	) name19022 (
		\u0_w_reg[3][1]/P0001 ,
		_w18860_,
		_w19554_
	);
	LUT2 #(
		.INIT('h1)
	) name19023 (
		ld_pad,
		_w19553_,
		_w19555_
	);
	LUT2 #(
		.INIT('h4)
	) name19024 (
		_w19554_,
		_w19555_,
		_w19556_
	);
	LUT2 #(
		.INIT('h8)
	) name19025 (
		\key[1]_pad ,
		ld_pad,
		_w19557_
	);
	LUT2 #(
		.INIT('h1)
	) name19026 (
		_w19556_,
		_w19557_,
		_w19558_
	);
	LUT2 #(
		.INIT('h4)
	) name19027 (
		\u0_w_reg[3][9]/P0001 ,
		_w18951_,
		_w19559_
	);
	LUT2 #(
		.INIT('h2)
	) name19028 (
		\u0_w_reg[3][9]/P0001 ,
		_w18951_,
		_w19560_
	);
	LUT2 #(
		.INIT('h1)
	) name19029 (
		ld_pad,
		_w19559_,
		_w19561_
	);
	LUT2 #(
		.INIT('h4)
	) name19030 (
		_w19560_,
		_w19561_,
		_w19562_
	);
	LUT2 #(
		.INIT('h8)
	) name19031 (
		\key[9]_pad ,
		ld_pad,
		_w19563_
	);
	LUT2 #(
		.INIT('h1)
	) name19032 (
		_w19562_,
		_w19563_,
		_w19564_
	);
	LUT2 #(
		.INIT('h1)
	) name19033 (
		\u0_w_reg[0][19]/P0001 ,
		_w14491_,
		_w19565_
	);
	LUT2 #(
		.INIT('h8)
	) name19034 (
		\u0_w_reg[0][19]/P0001 ,
		_w14491_,
		_w19566_
	);
	LUT2 #(
		.INIT('h1)
	) name19035 (
		_w19565_,
		_w19566_,
		_w19567_
	);
	LUT2 #(
		.INIT('h1)
	) name19036 (
		\u0_w_reg[3][19]/P0001 ,
		_w3966_,
		_w19568_
	);
	LUT2 #(
		.INIT('h8)
	) name19037 (
		\u0_w_reg[3][19]/P0001 ,
		_w3966_,
		_w19569_
	);
	LUT2 #(
		.INIT('h1)
	) name19038 (
		_w19568_,
		_w19569_,
		_w19570_
	);
	LUT2 #(
		.INIT('h1)
	) name19039 (
		\u0_w_reg[2][19]/P0001 ,
		_w7115_,
		_w19571_
	);
	LUT2 #(
		.INIT('h8)
	) name19040 (
		\u0_w_reg[2][19]/P0001 ,
		_w7115_,
		_w19572_
	);
	LUT2 #(
		.INIT('h1)
	) name19041 (
		_w19571_,
		_w19572_,
		_w19573_
	);
	LUT2 #(
		.INIT('h1)
	) name19042 (
		\u0_w_reg[1][19]/P0001 ,
		_w10682_,
		_w19574_
	);
	LUT2 #(
		.INIT('h8)
	) name19043 (
		\u0_w_reg[1][19]/P0001 ,
		_w10682_,
		_w19575_
	);
	LUT2 #(
		.INIT('h1)
	) name19044 (
		_w19574_,
		_w19575_,
		_w19576_
	);
	LUT2 #(
		.INIT('h1)
	) name19045 (
		\u0_w_reg[0][9]/P0001 ,
		_w13835_,
		_w19577_
	);
	LUT2 #(
		.INIT('h8)
	) name19046 (
		\u0_w_reg[0][9]/P0001 ,
		_w13835_,
		_w19578_
	);
	LUT2 #(
		.INIT('h1)
	) name19047 (
		_w19577_,
		_w19578_,
		_w19579_
	);
	LUT2 #(
		.INIT('h1)
	) name19048 (
		\u0_w_reg[2][9]/P0001 ,
		_w6743_,
		_w19580_
	);
	LUT2 #(
		.INIT('h8)
	) name19049 (
		\u0_w_reg[2][9]/P0001 ,
		_w6743_,
		_w19581_
	);
	LUT2 #(
		.INIT('h1)
	) name19050 (
		_w19580_,
		_w19581_,
		_w19582_
	);
	LUT2 #(
		.INIT('h1)
	) name19051 (
		\u0_w_reg[1][9]/P0001 ,
		_w10508_,
		_w19583_
	);
	LUT2 #(
		.INIT('h8)
	) name19052 (
		\u0_w_reg[1][9]/P0001 ,
		_w10508_,
		_w19584_
	);
	LUT2 #(
		.INIT('h1)
	) name19053 (
		_w19583_,
		_w19584_,
		_w19585_
	);
	LUT2 #(
		.INIT('h1)
	) name19054 (
		\u0_w_reg[0][13]/P0001 ,
		_w12405_,
		_w19586_
	);
	LUT2 #(
		.INIT('h8)
	) name19055 (
		\u0_w_reg[0][13]/P0001 ,
		_w12405_,
		_w19587_
	);
	LUT2 #(
		.INIT('h1)
	) name19056 (
		_w19586_,
		_w19587_,
		_w19588_
	);
	LUT2 #(
		.INIT('h1)
	) name19057 (
		\u0_w_reg[0][21]/P0001 ,
		_w12233_,
		_w19589_
	);
	LUT2 #(
		.INIT('h8)
	) name19058 (
		\u0_w_reg[0][21]/P0001 ,
		_w12233_,
		_w19590_
	);
	LUT2 #(
		.INIT('h1)
	) name19059 (
		_w19589_,
		_w19590_,
		_w19591_
	);
	LUT2 #(
		.INIT('h1)
	) name19060 (
		\u0_w_reg[3][13]/P0001 ,
		_w2939_,
		_w19592_
	);
	LUT2 #(
		.INIT('h8)
	) name19061 (
		\u0_w_reg[3][13]/P0001 ,
		_w2939_,
		_w19593_
	);
	LUT2 #(
		.INIT('h1)
	) name19062 (
		_w19592_,
		_w19593_,
		_w19594_
	);
	LUT2 #(
		.INIT('h1)
	) name19063 (
		\u0_w_reg[3][21]/P0001 ,
		_w2835_,
		_w19595_
	);
	LUT2 #(
		.INIT('h8)
	) name19064 (
		\u0_w_reg[3][21]/P0001 ,
		_w2835_,
		_w19596_
	);
	LUT2 #(
		.INIT('h1)
	) name19065 (
		_w19595_,
		_w19596_,
		_w19597_
	);
	LUT2 #(
		.INIT('h1)
	) name19066 (
		\u0_w_reg[2][13]/P0001 ,
		_w5931_,
		_w19598_
	);
	LUT2 #(
		.INIT('h8)
	) name19067 (
		\u0_w_reg[2][13]/P0001 ,
		_w5931_,
		_w19599_
	);
	LUT2 #(
		.INIT('h1)
	) name19068 (
		_w19598_,
		_w19599_,
		_w19600_
	);
	LUT2 #(
		.INIT('h1)
	) name19069 (
		\u0_w_reg[2][21]/P0001 ,
		_w973_,
		_w19601_
	);
	LUT2 #(
		.INIT('h8)
	) name19070 (
		\u0_w_reg[2][21]/P0001 ,
		_w973_,
		_w19602_
	);
	LUT2 #(
		.INIT('h1)
	) name19071 (
		_w19601_,
		_w19602_,
		_w19603_
	);
	LUT2 #(
		.INIT('h1)
	) name19072 (
		\u0_w_reg[1][13]/P0001 ,
		_w8678_,
		_w19604_
	);
	LUT2 #(
		.INIT('h8)
	) name19073 (
		\u0_w_reg[1][13]/P0001 ,
		_w8678_,
		_w19605_
	);
	LUT2 #(
		.INIT('h1)
	) name19074 (
		_w19604_,
		_w19605_,
		_w19606_
	);
	LUT2 #(
		.INIT('h1)
	) name19075 (
		\u0_w_reg[1][21]/P0001 ,
		_w8507_,
		_w19607_
	);
	LUT2 #(
		.INIT('h8)
	) name19076 (
		\u0_w_reg[1][21]/P0001 ,
		_w8507_,
		_w19608_
	);
	LUT2 #(
		.INIT('h1)
	) name19077 (
		_w19607_,
		_w19608_,
		_w19609_
	);
	LUT2 #(
		.INIT('h4)
	) name19078 (
		ld_pad,
		_w19039_,
		_w19610_
	);
	LUT2 #(
		.INIT('h8)
	) name19079 (
		\key[116]_pad ,
		ld_pad,
		_w19611_
	);
	LUT2 #(
		.INIT('h1)
	) name19080 (
		_w19610_,
		_w19611_,
		_w19612_
	);
	LUT2 #(
		.INIT('h4)
	) name19081 (
		ld_pad,
		_w19130_,
		_w19613_
	);
	LUT2 #(
		.INIT('h8)
	) name19082 (
		\key[100]_pad ,
		ld_pad,
		_w19614_
	);
	LUT2 #(
		.INIT('h1)
	) name19083 (
		_w19613_,
		_w19614_,
		_w19615_
	);
	LUT2 #(
		.INIT('h4)
	) name19084 (
		ld_pad,
		_w19042_,
		_w19616_
	);
	LUT2 #(
		.INIT('h8)
	) name19085 (
		\key[84]_pad ,
		ld_pad,
		_w19617_
	);
	LUT2 #(
		.INIT('h1)
	) name19086 (
		_w19616_,
		_w19617_,
		_w19618_
	);
	LUT2 #(
		.INIT('h1)
	) name19087 (
		\u0_w_reg[1][4]/P0001 ,
		_w19130_,
		_w19619_
	);
	LUT2 #(
		.INIT('h8)
	) name19088 (
		\u0_w_reg[1][4]/P0001 ,
		_w19130_,
		_w19620_
	);
	LUT2 #(
		.INIT('h1)
	) name19089 (
		ld_pad,
		_w19619_,
		_w19621_
	);
	LUT2 #(
		.INIT('h4)
	) name19090 (
		_w19620_,
		_w19621_,
		_w19622_
	);
	LUT2 #(
		.INIT('h8)
	) name19091 (
		\key[68]_pad ,
		ld_pad,
		_w19623_
	);
	LUT2 #(
		.INIT('h1)
	) name19092 (
		_w19622_,
		_w19623_,
		_w19624_
	);
	LUT2 #(
		.INIT('h1)
	) name19093 (
		\u0_w_reg[3][20]/P0001 ,
		_w19045_,
		_w19625_
	);
	LUT2 #(
		.INIT('h8)
	) name19094 (
		\u0_w_reg[3][20]/P0001 ,
		_w19045_,
		_w19626_
	);
	LUT2 #(
		.INIT('h1)
	) name19095 (
		ld_pad,
		_w19625_,
		_w19627_
	);
	LUT2 #(
		.INIT('h4)
	) name19096 (
		_w19626_,
		_w19627_,
		_w19628_
	);
	LUT2 #(
		.INIT('h8)
	) name19097 (
		\key[20]_pad ,
		ld_pad,
		_w19629_
	);
	LUT2 #(
		.INIT('h1)
	) name19098 (
		_w19628_,
		_w19629_,
		_w19630_
	);
	LUT2 #(
		.INIT('h4)
	) name19099 (
		\u0_w_reg[3][4]/P0001 ,
		_w19136_,
		_w19631_
	);
	LUT2 #(
		.INIT('h2)
	) name19100 (
		\u0_w_reg[3][4]/P0001 ,
		_w19136_,
		_w19632_
	);
	LUT2 #(
		.INIT('h1)
	) name19101 (
		ld_pad,
		_w19631_,
		_w19633_
	);
	LUT2 #(
		.INIT('h4)
	) name19102 (
		_w19632_,
		_w19633_,
		_w19634_
	);
	LUT2 #(
		.INIT('h8)
	) name19103 (
		\key[4]_pad ,
		ld_pad,
		_w19635_
	);
	LUT2 #(
		.INIT('h1)
	) name19104 (
		_w19634_,
		_w19635_,
		_w19636_
	);
	LUT2 #(
		.INIT('h1)
	) name19105 (
		\u0_w_reg[0][3]/P0001 ,
		_w14651_,
		_w19637_
	);
	LUT2 #(
		.INIT('h8)
	) name19106 (
		\u0_w_reg[0][3]/P0001 ,
		_w14651_,
		_w19638_
	);
	LUT2 #(
		.INIT('h1)
	) name19107 (
		_w19637_,
		_w19638_,
		_w19639_
	);
	LUT2 #(
		.INIT('h1)
	) name19108 (
		\u0_w_reg[3][9]/P0001 ,
		_w4248_,
		_w19640_
	);
	LUT2 #(
		.INIT('h8)
	) name19109 (
		\u0_w_reg[3][9]/P0001 ,
		_w4248_,
		_w19641_
	);
	LUT2 #(
		.INIT('h1)
	) name19110 (
		_w19640_,
		_w19641_,
		_w19642_
	);
	LUT2 #(
		.INIT('h1)
	) name19111 (
		\u0_w_reg[0][17]/P0001 ,
		_w14210_,
		_w19643_
	);
	LUT2 #(
		.INIT('h8)
	) name19112 (
		\u0_w_reg[0][17]/P0001 ,
		_w14210_,
		_w19644_
	);
	LUT2 #(
		.INIT('h1)
	) name19113 (
		_w19643_,
		_w19644_,
		_w19645_
	);
	LUT2 #(
		.INIT('h1)
	) name19114 (
		\u0_w_reg[3][17]/P0001 ,
		_w3681_,
		_w19646_
	);
	LUT2 #(
		.INIT('h8)
	) name19115 (
		\u0_w_reg[3][17]/P0001 ,
		_w3681_,
		_w19647_
	);
	LUT2 #(
		.INIT('h1)
	) name19116 (
		_w19646_,
		_w19647_,
		_w19648_
	);
	LUT2 #(
		.INIT('h1)
	) name19117 (
		\u0_w_reg[2][17]/P0001 ,
		_w6304_,
		_w19649_
	);
	LUT2 #(
		.INIT('h8)
	) name19118 (
		\u0_w_reg[2][17]/P0001 ,
		_w6304_,
		_w19650_
	);
	LUT2 #(
		.INIT('h1)
	) name19119 (
		_w19649_,
		_w19650_,
		_w19651_
	);
	LUT2 #(
		.INIT('h1)
	) name19120 (
		\u0_w_reg[1][17]/P0001 ,
		_w10081_,
		_w19652_
	);
	LUT2 #(
		.INIT('h8)
	) name19121 (
		\u0_w_reg[1][17]/P0001 ,
		_w10081_,
		_w19653_
	);
	LUT2 #(
		.INIT('h1)
	) name19122 (
		_w19652_,
		_w19653_,
		_w19654_
	);
	LUT2 #(
		.INIT('h1)
	) name19123 (
		\u0_w_reg[0][4]/P0001 ,
		_w12962_,
		_w19655_
	);
	LUT2 #(
		.INIT('h8)
	) name19124 (
		\u0_w_reg[0][4]/P0001 ,
		_w12962_,
		_w19656_
	);
	LUT2 #(
		.INIT('h1)
	) name19125 (
		_w19655_,
		_w19656_,
		_w19657_
	);
	LUT2 #(
		.INIT('h1)
	) name19126 (
		\u0_w_reg[3][12]/P0001 ,
		_w3069_,
		_w19658_
	);
	LUT2 #(
		.INIT('h8)
	) name19127 (
		\u0_w_reg[3][12]/P0001 ,
		_w3069_,
		_w19659_
	);
	LUT2 #(
		.INIT('h1)
	) name19128 (
		_w19658_,
		_w19659_,
		_w19660_
	);
	LUT2 #(
		.INIT('h1)
	) name19129 (
		\u0_w_reg[0][16]/P0001 ,
		_w13465_,
		_w19661_
	);
	LUT2 #(
		.INIT('h8)
	) name19130 (
		\u0_w_reg[0][16]/P0001 ,
		_w13465_,
		_w19662_
	);
	LUT2 #(
		.INIT('h1)
	) name19131 (
		_w19661_,
		_w19662_,
		_w19663_
	);
	LUT2 #(
		.INIT('h1)
	) name19132 (
		\u0_w_reg[3][16]/P0001 ,
		_w4674_,
		_w19664_
	);
	LUT2 #(
		.INIT('h8)
	) name19133 (
		\u0_w_reg[3][16]/P0001 ,
		_w4674_,
		_w19665_
	);
	LUT2 #(
		.INIT('h1)
	) name19134 (
		_w19664_,
		_w19665_,
		_w19666_
	);
	LUT2 #(
		.INIT('h1)
	) name19135 (
		\u0_w_reg[2][16]/P0001 ,
		_w7408_,
		_w19667_
	);
	LUT2 #(
		.INIT('h8)
	) name19136 (
		\u0_w_reg[2][16]/P0001 ,
		_w7408_,
		_w19668_
	);
	LUT2 #(
		.INIT('h1)
	) name19137 (
		_w19667_,
		_w19668_,
		_w19669_
	);
	LUT2 #(
		.INIT('h1)
	) name19138 (
		\u0_w_reg[1][16]/P0001 ,
		_w10996_,
		_w19670_
	);
	LUT2 #(
		.INIT('h8)
	) name19139 (
		\u0_w_reg[1][16]/P0001 ,
		_w10996_,
		_w19671_
	);
	LUT2 #(
		.INIT('h1)
	) name19140 (
		_w19670_,
		_w19671_,
		_w19672_
	);
	LUT2 #(
		.INIT('h1)
	) name19141 (
		\u0_w_reg[0][1]/P0001 ,
		_w13752_,
		_w19673_
	);
	LUT2 #(
		.INIT('h8)
	) name19142 (
		\u0_w_reg[0][1]/P0001 ,
		_w13752_,
		_w19674_
	);
	LUT2 #(
		.INIT('h1)
	) name19143 (
		_w19673_,
		_w19674_,
		_w19675_
	);
	LUT2 #(
		.INIT('h1)
	) name19144 (
		\u0_w_reg[0][6]/P0001 ,
		_w15289_,
		_w19676_
	);
	LUT2 #(
		.INIT('h8)
	) name19145 (
		\u0_w_reg[0][6]/P0001 ,
		_w15289_,
		_w19677_
	);
	LUT2 #(
		.INIT('h1)
	) name19146 (
		_w19676_,
		_w19677_,
		_w19678_
	);
	LUT2 #(
		.INIT('h1)
	) name19147 (
		\u0_w_reg[0][0]/P0001 ,
		_w14113_,
		_w19679_
	);
	LUT2 #(
		.INIT('h8)
	) name19148 (
		\u0_w_reg[0][0]/P0001 ,
		_w14113_,
		_w19680_
	);
	LUT2 #(
		.INIT('h1)
	) name19149 (
		_w19679_,
		_w19680_,
		_w19681_
	);
	LUT2 #(
		.INIT('h1)
	) name19150 (
		\u0_w_reg[0][10]/P0001 ,
		_w14894_,
		_w19682_
	);
	LUT2 #(
		.INIT('h8)
	) name19151 (
		\u0_w_reg[0][10]/P0001 ,
		_w14894_,
		_w19683_
	);
	LUT2 #(
		.INIT('h1)
	) name19152 (
		_w19682_,
		_w19683_,
		_w19684_
	);
	LUT2 #(
		.INIT('h1)
	) name19153 (
		\u0_w_reg[0][15]/P0001 ,
		_w13922_,
		_w19685_
	);
	LUT2 #(
		.INIT('h8)
	) name19154 (
		\u0_w_reg[0][15]/P0001 ,
		_w13922_,
		_w19686_
	);
	LUT2 #(
		.INIT('h1)
	) name19155 (
		_w19685_,
		_w19686_,
		_w19687_
	);
	LUT2 #(
		.INIT('h1)
	) name19156 (
		\u0_w_reg[0][31]/P0001 ,
		_w14400_,
		_w19688_
	);
	LUT2 #(
		.INIT('h8)
	) name19157 (
		\u0_w_reg[0][31]/P0001 ,
		_w14400_,
		_w19689_
	);
	LUT2 #(
		.INIT('h1)
	) name19158 (
		_w19688_,
		_w19689_,
		_w19690_
	);
	LUT2 #(
		.INIT('h1)
	) name19159 (
		\u0_w_reg[3][31]/P0001 ,
		_w2304_,
		_w19691_
	);
	LUT2 #(
		.INIT('h8)
	) name19160 (
		\u0_w_reg[3][31]/P0001 ,
		_w2304_,
		_w19692_
	);
	LUT2 #(
		.INIT('h1)
	) name19161 (
		_w19691_,
		_w19692_,
		_w19693_
	);
	LUT2 #(
		.INIT('h1)
	) name19162 (
		\u0_w_reg[2][10]/P0001 ,
		_w7655_,
		_w19694_
	);
	LUT2 #(
		.INIT('h8)
	) name19163 (
		\u0_w_reg[2][10]/P0001 ,
		_w7655_,
		_w19695_
	);
	LUT2 #(
		.INIT('h1)
	) name19164 (
		_w19694_,
		_w19695_,
		_w19696_
	);
	LUT2 #(
		.INIT('h1)
	) name19165 (
		\u0_w_reg[2][15]/P0001 ,
		_w5631_,
		_w19697_
	);
	LUT2 #(
		.INIT('h8)
	) name19166 (
		\u0_w_reg[2][15]/P0001 ,
		_w5631_,
		_w19698_
	);
	LUT2 #(
		.INIT('h1)
	) name19167 (
		_w19697_,
		_w19698_,
		_w19699_
	);
	LUT2 #(
		.INIT('h1)
	) name19168 (
		\u0_w_reg[2][31]/P0001 ,
		_w5417_,
		_w19700_
	);
	LUT2 #(
		.INIT('h8)
	) name19169 (
		\u0_w_reg[2][31]/P0001 ,
		_w5417_,
		_w19701_
	);
	LUT2 #(
		.INIT('h1)
	) name19170 (
		_w19700_,
		_w19701_,
		_w19702_
	);
	LUT2 #(
		.INIT('h1)
	) name19171 (
		\u0_w_reg[1][10]/P0001 ,
		_w11384_,
		_w19703_
	);
	LUT2 #(
		.INIT('h8)
	) name19172 (
		\u0_w_reg[1][10]/P0001 ,
		_w11384_,
		_w19704_
	);
	LUT2 #(
		.INIT('h1)
	) name19173 (
		_w19703_,
		_w19704_,
		_w19705_
	);
	LUT2 #(
		.INIT('h1)
	) name19174 (
		\u0_w_reg[1][15]/P0001 ,
		_w9980_,
		_w19706_
	);
	LUT2 #(
		.INIT('h8)
	) name19175 (
		\u0_w_reg[1][15]/P0001 ,
		_w9980_,
		_w19707_
	);
	LUT2 #(
		.INIT('h1)
	) name19176 (
		_w19706_,
		_w19707_,
		_w19708_
	);
	LUT2 #(
		.INIT('h1)
	) name19177 (
		\u0_w_reg[1][31]/P0001 ,
		_w9783_,
		_w19709_
	);
	LUT2 #(
		.INIT('h8)
	) name19178 (
		\u0_w_reg[1][31]/P0001 ,
		_w9783_,
		_w19710_
	);
	LUT2 #(
		.INIT('h1)
	) name19179 (
		_w19709_,
		_w19710_,
		_w19711_
	);
	LUT2 #(
		.INIT('h1)
	) name19180 (
		\u0_w_reg[0][18]/P0001 ,
		_w14729_,
		_w19712_
	);
	LUT2 #(
		.INIT('h8)
	) name19181 (
		\u0_w_reg[0][18]/P0001 ,
		_w14729_,
		_w19713_
	);
	LUT2 #(
		.INIT('h1)
	) name19182 (
		_w19712_,
		_w19713_,
		_w19714_
	);
	LUT2 #(
		.INIT('h1)
	) name19183 (
		\u0_w_reg[3][18]/P0001 ,
		_w4433_,
		_w19715_
	);
	LUT2 #(
		.INIT('h8)
	) name19184 (
		\u0_w_reg[3][18]/P0001 ,
		_w4433_,
		_w19716_
	);
	LUT2 #(
		.INIT('h1)
	) name19185 (
		_w19715_,
		_w19716_,
		_w19717_
	);
	LUT2 #(
		.INIT('h1)
	) name19186 (
		\u0_w_reg[2][18]/P0001 ,
		_w7508_,
		_w19718_
	);
	LUT2 #(
		.INIT('h8)
	) name19187 (
		\u0_w_reg[2][18]/P0001 ,
		_w7508_,
		_w19719_
	);
	LUT2 #(
		.INIT('h1)
	) name19188 (
		_w19718_,
		_w19719_,
		_w19720_
	);
	LUT2 #(
		.INIT('h1)
	) name19189 (
		\u0_w_reg[1][18]/P0001 ,
		_w11240_,
		_w19721_
	);
	LUT2 #(
		.INIT('h8)
	) name19190 (
		\u0_w_reg[1][18]/P0001 ,
		_w11240_,
		_w19722_
	);
	LUT2 #(
		.INIT('h1)
	) name19191 (
		_w19721_,
		_w19722_,
		_w19723_
	);
	LUT2 #(
		.INIT('h1)
	) name19192 (
		\u0_w_reg[0][23]/P0001 ,
		_w13558_,
		_w19724_
	);
	LUT2 #(
		.INIT('h8)
	) name19193 (
		\u0_w_reg[0][23]/P0001 ,
		_w13558_,
		_w19725_
	);
	LUT2 #(
		.INIT('h1)
	) name19194 (
		_w19724_,
		_w19725_,
		_w19726_
	);
	LUT2 #(
		.INIT('h1)
	) name19195 (
		\u0_w_reg[3][15]/P0001 ,
		_w2529_,
		_w19727_
	);
	LUT2 #(
		.INIT('h8)
	) name19196 (
		\u0_w_reg[3][15]/P0001 ,
		_w2529_,
		_w19728_
	);
	LUT2 #(
		.INIT('h1)
	) name19197 (
		_w19727_,
		_w19728_,
		_w19729_
	);
	LUT2 #(
		.INIT('h1)
	) name19198 (
		\u0_w_reg[3][23]/P0001 ,
		_w2199_,
		_w19730_
	);
	LUT2 #(
		.INIT('h8)
	) name19199 (
		\u0_w_reg[3][23]/P0001 ,
		_w2199_,
		_w19731_
	);
	LUT2 #(
		.INIT('h1)
	) name19200 (
		_w19730_,
		_w19731_,
		_w19732_
	);
	LUT2 #(
		.INIT('h1)
	) name19201 (
		\u0_w_reg[2][23]/P0001 ,
		_w5516_,
		_w19733_
	);
	LUT2 #(
		.INIT('h8)
	) name19202 (
		\u0_w_reg[2][23]/P0001 ,
		_w5516_,
		_w19734_
	);
	LUT2 #(
		.INIT('h1)
	) name19203 (
		_w19733_,
		_w19734_,
		_w19735_
	);
	LUT2 #(
		.INIT('h1)
	) name19204 (
		\u0_w_reg[1][23]/P0001 ,
		_w9874_,
		_w19736_
	);
	LUT2 #(
		.INIT('h8)
	) name19205 (
		\u0_w_reg[1][23]/P0001 ,
		_w9874_,
		_w19737_
	);
	LUT2 #(
		.INIT('h1)
	) name19206 (
		_w19736_,
		_w19737_,
		_w19738_
	);
	LUT2 #(
		.INIT('h1)
	) name19207 (
		\u0_w_reg[0][26]/P0001 ,
		_w14801_,
		_w19739_
	);
	LUT2 #(
		.INIT('h8)
	) name19208 (
		\u0_w_reg[0][26]/P0001 ,
		_w14801_,
		_w19740_
	);
	LUT2 #(
		.INIT('h1)
	) name19209 (
		_w19739_,
		_w19740_,
		_w19741_
	);
	LUT2 #(
		.INIT('h1)
	) name19210 (
		\u0_w_reg[3][26]/P0001 ,
		_w4505_,
		_w19742_
	);
	LUT2 #(
		.INIT('h8)
	) name19211 (
		\u0_w_reg[3][26]/P0001 ,
		_w4505_,
		_w19743_
	);
	LUT2 #(
		.INIT('h1)
	) name19212 (
		_w19742_,
		_w19743_,
		_w19744_
	);
	LUT2 #(
		.INIT('h1)
	) name19213 (
		\u0_w_reg[2][26]/P0001 ,
		_w7580_,
		_w19745_
	);
	LUT2 #(
		.INIT('h8)
	) name19214 (
		\u0_w_reg[2][26]/P0001 ,
		_w7580_,
		_w19746_
	);
	LUT2 #(
		.INIT('h1)
	) name19215 (
		_w19745_,
		_w19746_,
		_w19747_
	);
	LUT2 #(
		.INIT('h1)
	) name19216 (
		\u0_w_reg[1][26]/P0001 ,
		_w11312_,
		_w19748_
	);
	LUT2 #(
		.INIT('h8)
	) name19217 (
		\u0_w_reg[1][26]/P0001 ,
		_w11312_,
		_w19749_
	);
	LUT2 #(
		.INIT('h1)
	) name19218 (
		_w19748_,
		_w19749_,
		_w19750_
	);
	LUT2 #(
		.INIT('h1)
	) name19219 (
		\u0_w_reg[0][7]/P0001 ,
		_w14033_,
		_w19751_
	);
	LUT2 #(
		.INIT('h8)
	) name19220 (
		\u0_w_reg[0][7]/P0001 ,
		_w14033_,
		_w19752_
	);
	LUT2 #(
		.INIT('h1)
	) name19221 (
		_w19751_,
		_w19752_,
		_w19753_
	);
	LUT2 #(
		.INIT('h1)
	) name19222 (
		\u0_w_reg[0][30]/P0001 ,
		_w13091_,
		_w19754_
	);
	LUT2 #(
		.INIT('h8)
	) name19223 (
		\u0_w_reg[0][30]/P0001 ,
		_w13091_,
		_w19755_
	);
	LUT2 #(
		.INIT('h1)
	) name19224 (
		_w19754_,
		_w19755_,
		_w19756_
	);
	LUT2 #(
		.INIT('h1)
	) name19225 (
		\u0_w_reg[3][30]/P0001 ,
		_w1581_,
		_w19757_
	);
	LUT2 #(
		.INIT('h8)
	) name19226 (
		\u0_w_reg[3][30]/P0001 ,
		_w1581_,
		_w19758_
	);
	LUT2 #(
		.INIT('h1)
	) name19227 (
		_w19757_,
		_w19758_,
		_w19759_
	);
	LUT2 #(
		.INIT('h1)
	) name19228 (
		\u0_w_reg[2][30]/P0001 ,
		_w5191_,
		_w19760_
	);
	LUT2 #(
		.INIT('h8)
	) name19229 (
		\u0_w_reg[2][30]/P0001 ,
		_w5191_,
		_w19761_
	);
	LUT2 #(
		.INIT('h1)
	) name19230 (
		_w19760_,
		_w19761_,
		_w19762_
	);
	LUT2 #(
		.INIT('h1)
	) name19231 (
		\u0_w_reg[1][30]/P0001 ,
		_w9400_,
		_w19763_
	);
	LUT2 #(
		.INIT('h8)
	) name19232 (
		\u0_w_reg[1][30]/P0001 ,
		_w9400_,
		_w19764_
	);
	LUT2 #(
		.INIT('h1)
	) name19233 (
		_w19763_,
		_w19764_,
		_w19765_
	);
	LUT2 #(
		.INIT('h1)
	) name19234 (
		\u0_w_reg[3][10]/P0001 ,
		_w4578_,
		_w19766_
	);
	LUT2 #(
		.INIT('h8)
	) name19235 (
		\u0_w_reg[3][10]/P0001 ,
		_w4578_,
		_w19767_
	);
	LUT2 #(
		.INIT('h1)
	) name19236 (
		_w19766_,
		_w19767_,
		_w19768_
	);
	LUT2 #(
		.INIT('h1)
	) name19237 (
		\u0_w_reg[0][14]/P0001 ,
		_w13284_,
		_w19769_
	);
	LUT2 #(
		.INIT('h8)
	) name19238 (
		\u0_w_reg[0][14]/P0001 ,
		_w13284_,
		_w19770_
	);
	LUT2 #(
		.INIT('h1)
	) name19239 (
		_w19769_,
		_w19770_,
		_w19771_
	);
	LUT2 #(
		.INIT('h1)
	) name19240 (
		\u0_w_reg[0][22]/P0001 ,
		_w13183_,
		_w19772_
	);
	LUT2 #(
		.INIT('h8)
	) name19241 (
		\u0_w_reg[0][22]/P0001 ,
		_w13183_,
		_w19773_
	);
	LUT2 #(
		.INIT('h1)
	) name19242 (
		_w19772_,
		_w19773_,
		_w19774_
	);
	LUT2 #(
		.INIT('h1)
	) name19243 (
		\u0_w_reg[3][14]/P0001 ,
		_w1908_,
		_w19775_
	);
	LUT2 #(
		.INIT('h8)
	) name19244 (
		\u0_w_reg[3][14]/P0001 ,
		_w1908_,
		_w19776_
	);
	LUT2 #(
		.INIT('h1)
	) name19245 (
		_w19775_,
		_w19776_,
		_w19777_
	);
	LUT2 #(
		.INIT('h1)
	) name19246 (
		\u0_w_reg[3][22]/P0001 ,
		_w1738_,
		_w19778_
	);
	LUT2 #(
		.INIT('h8)
	) name19247 (
		\u0_w_reg[3][22]/P0001 ,
		_w1738_,
		_w19779_
	);
	LUT2 #(
		.INIT('h1)
	) name19248 (
		_w19778_,
		_w19779_,
		_w19780_
	);
	LUT2 #(
		.INIT('h1)
	) name19249 (
		\u0_w_reg[2][14]/P0001 ,
		_w850_,
		_w19781_
	);
	LUT2 #(
		.INIT('h8)
	) name19250 (
		\u0_w_reg[2][14]/P0001 ,
		_w850_,
		_w19782_
	);
	LUT2 #(
		.INIT('h1)
	) name19251 (
		_w19781_,
		_w19782_,
		_w19783_
	);
	LUT2 #(
		.INIT('h1)
	) name19252 (
		\u0_w_reg[2][22]/P0001 ,
		_w689_,
		_w19784_
	);
	LUT2 #(
		.INIT('h8)
	) name19253 (
		\u0_w_reg[2][22]/P0001 ,
		_w689_,
		_w19785_
	);
	LUT2 #(
		.INIT('h1)
	) name19254 (
		_w19784_,
		_w19785_,
		_w19786_
	);
	LUT2 #(
		.INIT('h1)
	) name19255 (
		\u0_w_reg[1][14]/P0001 ,
		_w9169_,
		_w19787_
	);
	LUT2 #(
		.INIT('h8)
	) name19256 (
		\u0_w_reg[1][14]/P0001 ,
		_w9169_,
		_w19788_
	);
	LUT2 #(
		.INIT('h1)
	) name19257 (
		_w19787_,
		_w19788_,
		_w19789_
	);
	LUT2 #(
		.INIT('h1)
	) name19258 (
		\u0_w_reg[1][22]/P0001 ,
		_w9063_,
		_w19790_
	);
	LUT2 #(
		.INIT('h8)
	) name19259 (
		\u0_w_reg[1][22]/P0001 ,
		_w9063_,
		_w19791_
	);
	LUT2 #(
		.INIT('h1)
	) name19260 (
		_w19790_,
		_w19791_,
		_w19792_
	);
	LUT2 #(
		.INIT('h1)
	) name19261 (
		\u0_w_reg[0][2]/P0001 ,
		_w15068_,
		_w19793_
	);
	LUT2 #(
		.INIT('h8)
	) name19262 (
		\u0_w_reg[0][2]/P0001 ,
		_w15068_,
		_w19794_
	);
	LUT2 #(
		.INIT('h1)
	) name19263 (
		_w19793_,
		_w19794_,
		_w19795_
	);
	LUT2 #(
		.INIT('h1)
	) name19264 (
		\u0_w_reg[0][25]/P0001 ,
		_w13649_,
		_w19796_
	);
	LUT2 #(
		.INIT('h8)
	) name19265 (
		\u0_w_reg[0][25]/P0001 ,
		_w13649_,
		_w19797_
	);
	LUT2 #(
		.INIT('h1)
	) name19266 (
		_w19796_,
		_w19797_,
		_w19798_
	);
	LUT2 #(
		.INIT('h1)
	) name19267 (
		\u0_w_reg[3][25]/P0001 ,
		_w3768_,
		_w19799_
	);
	LUT2 #(
		.INIT('h8)
	) name19268 (
		\u0_w_reg[3][25]/P0001 ,
		_w3768_,
		_w19800_
	);
	LUT2 #(
		.INIT('h1)
	) name19269 (
		_w19799_,
		_w19800_,
		_w19801_
	);
	LUT2 #(
		.INIT('h1)
	) name19270 (
		\u0_w_reg[2][25]/P0001 ,
		_w6392_,
		_w19802_
	);
	LUT2 #(
		.INIT('h8)
	) name19271 (
		\u0_w_reg[2][25]/P0001 ,
		_w6392_,
		_w19803_
	);
	LUT2 #(
		.INIT('h1)
	) name19272 (
		_w19802_,
		_w19803_,
		_w19804_
	);
	LUT2 #(
		.INIT('h1)
	) name19273 (
		\u0_w_reg[1][25]/P0001 ,
		_w10167_,
		_w19805_
	);
	LUT2 #(
		.INIT('h8)
	) name19274 (
		\u0_w_reg[1][25]/P0001 ,
		_w10167_,
		_w19806_
	);
	LUT2 #(
		.INIT('h1)
	) name19275 (
		_w19805_,
		_w19806_,
		_w19807_
	);
	LUT2 #(
		.INIT('h1)
	) name19276 (
		\u0_w_reg[0][20]/P0001 ,
		_w11951_,
		_w19808_
	);
	LUT2 #(
		.INIT('h8)
	) name19277 (
		\u0_w_reg[0][20]/P0001 ,
		_w11951_,
		_w19809_
	);
	LUT2 #(
		.INIT('h1)
	) name19278 (
		_w19808_,
		_w19809_,
		_w19810_
	);
	LUT2 #(
		.INIT('h1)
	) name19279 (
		\u0_w_reg[3][20]/P0001 ,
		_w2647_,
		_w19811_
	);
	LUT2 #(
		.INIT('h8)
	) name19280 (
		\u0_w_reg[3][20]/P0001 ,
		_w2647_,
		_w19812_
	);
	LUT2 #(
		.INIT('h1)
	) name19281 (
		_w19811_,
		_w19812_,
		_w19813_
	);
	LUT2 #(
		.INIT('h1)
	) name19282 (
		\u0_w_reg[2][20]/P0001 ,
		_w5737_,
		_w19814_
	);
	LUT2 #(
		.INIT('h8)
	) name19283 (
		\u0_w_reg[2][20]/P0001 ,
		_w5737_,
		_w19815_
	);
	LUT2 #(
		.INIT('h1)
	) name19284 (
		_w19814_,
		_w19815_,
		_w19816_
	);
	LUT2 #(
		.INIT('h1)
	) name19285 (
		\u0_w_reg[1][20]/P0001 ,
		_w8213_,
		_w19817_
	);
	LUT2 #(
		.INIT('h8)
	) name19286 (
		\u0_w_reg[1][20]/P0001 ,
		_w8213_,
		_w19818_
	);
	LUT2 #(
		.INIT('h1)
	) name19287 (
		_w19817_,
		_w19818_,
		_w19819_
	);
	LUT2 #(
		.INIT('h1)
	) name19288 (
		\u0_w_reg[0][28]/P0001 ,
		_w12111_,
		_w19820_
	);
	LUT2 #(
		.INIT('h8)
	) name19289 (
		\u0_w_reg[0][28]/P0001 ,
		_w12111_,
		_w19821_
	);
	LUT2 #(
		.INIT('h1)
	) name19290 (
		_w19820_,
		_w19821_,
		_w19822_
	);
	LUT2 #(
		.INIT('h1)
	) name19291 (
		\u0_w_reg[3][28]/P0001 ,
		_w2736_,
		_w19823_
	);
	LUT2 #(
		.INIT('h8)
	) name19292 (
		\u0_w_reg[3][28]/P0001 ,
		_w2736_,
		_w19824_
	);
	LUT2 #(
		.INIT('h1)
	) name19293 (
		_w19823_,
		_w19824_,
		_w19825_
	);
	LUT2 #(
		.INIT('h1)
	) name19294 (
		\u0_w_reg[2][28]/P0001 ,
		_w5830_,
		_w19826_
	);
	LUT2 #(
		.INIT('h8)
	) name19295 (
		\u0_w_reg[2][28]/P0001 ,
		_w5830_,
		_w19827_
	);
	LUT2 #(
		.INIT('h1)
	) name19296 (
		_w19826_,
		_w19827_,
		_w19828_
	);
	LUT2 #(
		.INIT('h1)
	) name19297 (
		\u0_w_reg[1][28]/P0001 ,
		_w8376_,
		_w19829_
	);
	LUT2 #(
		.INIT('h8)
	) name19298 (
		\u0_w_reg[1][28]/P0001 ,
		_w8376_,
		_w19830_
	);
	LUT2 #(
		.INIT('h1)
	) name19299 (
		_w19829_,
		_w19830_,
		_w19831_
	);
	LUT2 #(
		.INIT('h8)
	) name19300 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		\u0_r0_rcnt_reg[1]/P0001 ,
		_w19832_
	);
	LUT2 #(
		.INIT('h1)
	) name19301 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		\u0_r0_rcnt_reg[1]/P0001 ,
		_w19833_
	);
	LUT2 #(
		.INIT('h1)
	) name19302 (
		_w19832_,
		_w19833_,
		_w19834_
	);
	LUT2 #(
		.INIT('h8)
	) name19303 (
		\u0_r0_rcnt_reg[2]/P0001 ,
		_w19832_,
		_w19835_
	);
	LUT2 #(
		.INIT('h1)
	) name19304 (
		\u0_r0_rcnt_reg[2]/P0001 ,
		_w19832_,
		_w19836_
	);
	LUT2 #(
		.INIT('h1)
	) name19305 (
		_w19835_,
		_w19836_,
		_w19837_
	);
	LUT2 #(
		.INIT('h4)
	) name19306 (
		\u0_r0_rcnt_reg[3]/P0001 ,
		_w19837_,
		_w19838_
	);
	LUT2 #(
		.INIT('h4)
	) name19307 (
		_w19834_,
		_w19838_,
		_w19839_
	);
	LUT2 #(
		.INIT('h2)
	) name19308 (
		\u0_r0_rcnt_reg[3]/P0001 ,
		_w19835_,
		_w19840_
	);
	LUT2 #(
		.INIT('h4)
	) name19309 (
		\u0_r0_rcnt_reg[3]/P0001 ,
		_w19835_,
		_w19841_
	);
	LUT2 #(
		.INIT('h1)
	) name19310 (
		_w19840_,
		_w19841_,
		_w19842_
	);
	LUT2 #(
		.INIT('h1)
	) name19311 (
		_w19834_,
		_w19837_,
		_w19843_
	);
	LUT2 #(
		.INIT('h4)
	) name19312 (
		_w19842_,
		_w19843_,
		_w19844_
	);
	LUT2 #(
		.INIT('h1)
	) name19313 (
		_w19839_,
		_w19844_,
		_w19845_
	);
	LUT2 #(
		.INIT('h1)
	) name19314 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		_w19844_,
		_w19846_
	);
	LUT2 #(
		.INIT('h1)
	) name19315 (
		ld_pad,
		_w19846_,
		_w19847_
	);
	LUT2 #(
		.INIT('h4)
	) name19316 (
		_w19845_,
		_w19847_,
		_w19848_
	);
	LUT2 #(
		.INIT('h2)
	) name19317 (
		_w19834_,
		_w19837_,
		_w19849_
	);
	LUT2 #(
		.INIT('h8)
	) name19318 (
		_w19842_,
		_w19849_,
		_w19850_
	);
	LUT2 #(
		.INIT('h2)
	) name19319 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		_w19850_,
		_w19851_
	);
	LUT2 #(
		.INIT('h2)
	) name19320 (
		_w19847_,
		_w19851_,
		_w19852_
	);
	LUT2 #(
		.INIT('h1)
	) name19321 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		_w19850_,
		_w19853_
	);
	LUT2 #(
		.INIT('h2)
	) name19322 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		_w19844_,
		_w19854_
	);
	LUT2 #(
		.INIT('h1)
	) name19323 (
		ld_pad,
		_w19853_,
		_w19855_
	);
	LUT2 #(
		.INIT('h4)
	) name19324 (
		_w19854_,
		_w19855_,
		_w19856_
	);
	LUT2 #(
		.INIT('h1)
	) name19325 (
		ld_pad,
		\u0_r0_rcnt_reg[0]/P0001 ,
		_w19857_
	);
	LUT2 #(
		.INIT('h4)
	) name19326 (
		_w19845_,
		_w19857_,
		_w19858_
	);
	LUT2 #(
		.INIT('h4)
	) name19327 (
		\u0_r0_rcnt_reg[2]/P0001 ,
		_w19833_,
		_w19859_
	);
	LUT2 #(
		.INIT('h1)
	) name19328 (
		_w19844_,
		_w19859_,
		_w19860_
	);
	LUT2 #(
		.INIT('h1)
	) name19329 (
		ld_pad,
		_w19860_,
		_w19861_
	);
	LUT2 #(
		.INIT('h4)
	) name19330 (
		ld_pad,
		_w19834_,
		_w19862_
	);
	LUT2 #(
		.INIT('h4)
	) name19331 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		_w19862_,
		_w19863_
	);
	LUT2 #(
		.INIT('h8)
	) name19332 (
		_w19838_,
		_w19863_,
		_w19864_
	);
	LUT2 #(
		.INIT('h8)
	) name19333 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		_w19862_,
		_w19865_
	);
	LUT2 #(
		.INIT('h8)
	) name19334 (
		_w19838_,
		_w19865_,
		_w19866_
	);
	LUT2 #(
		.INIT('h1)
	) name19335 (
		\dcnt_reg[0]/P0001 ,
		\dcnt_reg[1]/P0001 ,
		_w19867_
	);
	LUT2 #(
		.INIT('h4)
	) name19336 (
		\dcnt_reg[2]/P0001 ,
		_w19867_,
		_w19868_
	);
	LUT2 #(
		.INIT('h2)
	) name19337 (
		\dcnt_reg[3]/P0001 ,
		_w19868_,
		_w19869_
	);
	LUT2 #(
		.INIT('h1)
	) name19338 (
		ld_pad,
		_w19869_,
		_w19870_
	);
	LUT2 #(
		.INIT('h2)
	) name19339 (
		rst_pad,
		_w19870_,
		_w19871_
	);
	LUT2 #(
		.INIT('h1)
	) name19340 (
		ld_pad,
		_w19842_,
		_w19872_
	);
	LUT2 #(
		.INIT('h1)
	) name19341 (
		ld_pad,
		_w19835_,
		_w19873_
	);
	LUT2 #(
		.INIT('h2)
	) name19342 (
		\dcnt_reg[2]/P0001 ,
		_w19867_,
		_w19874_
	);
	LUT2 #(
		.INIT('h8)
	) name19343 (
		\dcnt_reg[3]/P0001 ,
		_w19868_,
		_w19875_
	);
	LUT2 #(
		.INIT('h1)
	) name19344 (
		_w19874_,
		_w19875_,
		_w19876_
	);
	LUT2 #(
		.INIT('h4)
	) name19345 (
		ld_pad,
		rst_pad,
		_w19877_
	);
	LUT2 #(
		.INIT('h4)
	) name19346 (
		_w19876_,
		_w19877_,
		_w19878_
	);
	LUT2 #(
		.INIT('h8)
	) name19347 (
		ld_pad,
		rst_pad,
		_w19879_
	);
	LUT2 #(
		.INIT('h1)
	) name19348 (
		\dcnt_reg[2]/P0001 ,
		\dcnt_reg[3]/P0001 ,
		_w19880_
	);
	LUT2 #(
		.INIT('h8)
	) name19349 (
		_w19867_,
		_w19880_,
		_w19881_
	);
	LUT2 #(
		.INIT('h2)
	) name19350 (
		rst_pad,
		_w19881_,
		_w19882_
	);
	LUT2 #(
		.INIT('h4)
	) name19351 (
		\dcnt_reg[0]/P0001 ,
		_w19882_,
		_w19883_
	);
	LUT2 #(
		.INIT('h1)
	) name19352 (
		_w19879_,
		_w19883_,
		_w19884_
	);
	LUT2 #(
		.INIT('h8)
	) name19353 (
		\dcnt_reg[0]/P0001 ,
		\dcnt_reg[1]/P0001 ,
		_w19885_
	);
	LUT2 #(
		.INIT('h1)
	) name19354 (
		_w19867_,
		_w19885_,
		_w19886_
	);
	LUT2 #(
		.INIT('h2)
	) name19355 (
		_w19882_,
		_w19886_,
		_w19887_
	);
	LUT2 #(
		.INIT('h1)
	) name19356 (
		_w19879_,
		_w19887_,
		_w19888_
	);
	LUT2 #(
		.INIT('h4)
	) name19357 (
		ld_pad,
		_w19837_,
		_w19889_
	);
	LUT2 #(
		.INIT('h2)
	) name19358 (
		\dcnt_reg[0]/P0001 ,
		\dcnt_reg[1]/P0001 ,
		_w19890_
	);
	LUT2 #(
		.INIT('h4)
	) name19359 (
		ld_pad,
		_w19890_,
		_w19891_
	);
	LUT2 #(
		.INIT('h8)
	) name19360 (
		_w19880_,
		_w19891_,
		_w19892_
	);
	LUT2 #(
		.INIT('h2)
	) name19361 (
		\u0_w_reg[1][9]/P0001 ,
		_w11155_,
		_w19893_
	);
	LUT2 #(
		.INIT('h4)
	) name19362 (
		\u0_w_reg[1][9]/P0001 ,
		_w11155_,
		_w19894_
	);
	LUT2 #(
		.INIT('h1)
	) name19363 (
		_w19893_,
		_w19894_,
		_w19895_
	);
	LUT2 #(
		.INIT('h8)
	) name19364 (
		_w10433_,
		_w19895_,
		_w19896_
	);
	LUT2 #(
		.INIT('h1)
	) name19365 (
		_w10433_,
		_w19895_,
		_w19897_
	);
	LUT2 #(
		.INIT('h1)
	) name19366 (
		_w19896_,
		_w19897_,
		_w19898_
	);
	LUT2 #(
		.INIT('h8)
	) name19367 (
		_w10170_,
		_w11643_,
		_w19899_
	);
	LUT2 #(
		.INIT('h1)
	) name19368 (
		_w10170_,
		_w11643_,
		_w19900_
	);
	LUT2 #(
		.INIT('h1)
	) name19369 (
		_w19899_,
		_w19900_,
		_w19901_
	);
	LUT2 #(
		.INIT('h1)
	) name19370 (
		_w19898_,
		_w19901_,
		_w19902_
	);
	LUT2 #(
		.INIT('h8)
	) name19371 (
		_w19898_,
		_w19901_,
		_w19903_
	);
	LUT2 #(
		.INIT('h1)
	) name19372 (
		\ld_r_reg/P0001 ,
		_w19902_,
		_w19904_
	);
	LUT2 #(
		.INIT('h4)
	) name19373 (
		_w19903_,
		_w19904_,
		_w19905_
	);
	LUT2 #(
		.INIT('h1)
	) name19374 (
		\text_in_r_reg[73]/P0001 ,
		\u0_w_reg[1][9]/P0001 ,
		_w19906_
	);
	LUT2 #(
		.INIT('h8)
	) name19375 (
		\text_in_r_reg[73]/P0001 ,
		\u0_w_reg[1][9]/P0001 ,
		_w19907_
	);
	LUT2 #(
		.INIT('h2)
	) name19376 (
		\ld_r_reg/P0001 ,
		_w19906_,
		_w19908_
	);
	LUT2 #(
		.INIT('h4)
	) name19377 (
		_w19907_,
		_w19908_,
		_w19909_
	);
	LUT2 #(
		.INIT('h1)
	) name19378 (
		_w19905_,
		_w19909_,
		_w19910_
	);
	LUT2 #(
		.INIT('h2)
	) name19379 (
		\u0_w_reg[0][0]/P0001 ,
		_w14033_,
		_w19911_
	);
	LUT2 #(
		.INIT('h4)
	) name19380 (
		\u0_w_reg[0][0]/P0001 ,
		_w14033_,
		_w19912_
	);
	LUT2 #(
		.INIT('h1)
	) name19381 (
		_w19911_,
		_w19912_,
		_w19913_
	);
	LUT2 #(
		.INIT('h4)
	) name19382 (
		_w13468_,
		_w14403_,
		_w19914_
	);
	LUT2 #(
		.INIT('h2)
	) name19383 (
		_w13468_,
		_w14403_,
		_w19915_
	);
	LUT2 #(
		.INIT('h1)
	) name19384 (
		_w19914_,
		_w19915_,
		_w19916_
	);
	LUT2 #(
		.INIT('h1)
	) name19385 (
		_w19913_,
		_w19916_,
		_w19917_
	);
	LUT2 #(
		.INIT('h8)
	) name19386 (
		_w19913_,
		_w19916_,
		_w19918_
	);
	LUT2 #(
		.INIT('h1)
	) name19387 (
		\ld_r_reg/P0001 ,
		_w19917_,
		_w19919_
	);
	LUT2 #(
		.INIT('h4)
	) name19388 (
		_w19918_,
		_w19919_,
		_w19920_
	);
	LUT2 #(
		.INIT('h2)
	) name19389 (
		\text_in_r_reg[96]/P0001 ,
		\u0_w_reg[0][0]/P0001 ,
		_w19921_
	);
	LUT2 #(
		.INIT('h4)
	) name19390 (
		\text_in_r_reg[96]/P0001 ,
		\u0_w_reg[0][0]/P0001 ,
		_w19922_
	);
	LUT2 #(
		.INIT('h2)
	) name19391 (
		\ld_r_reg/P0001 ,
		_w19921_,
		_w19923_
	);
	LUT2 #(
		.INIT('h4)
	) name19392 (
		_w19922_,
		_w19923_,
		_w19924_
	);
	LUT2 #(
		.INIT('h1)
	) name19393 (
		_w19920_,
		_w19924_,
		_w19925_
	);
	LUT2 #(
		.INIT('h2)
	) name19394 (
		\u0_w_reg[1][0]/P0001 ,
		_w10430_,
		_w19926_
	);
	LUT2 #(
		.INIT('h4)
	) name19395 (
		\u0_w_reg[1][0]/P0001 ,
		_w10430_,
		_w19927_
	);
	LUT2 #(
		.INIT('h1)
	) name19396 (
		_w19926_,
		_w19927_,
		_w19928_
	);
	LUT2 #(
		.INIT('h8)
	) name19397 (
		_w10251_,
		_w11700_,
		_w19929_
	);
	LUT2 #(
		.INIT('h1)
	) name19398 (
		_w10251_,
		_w11700_,
		_w19930_
	);
	LUT2 #(
		.INIT('h1)
	) name19399 (
		_w19929_,
		_w19930_,
		_w19931_
	);
	LUT2 #(
		.INIT('h1)
	) name19400 (
		_w19928_,
		_w19931_,
		_w19932_
	);
	LUT2 #(
		.INIT('h8)
	) name19401 (
		_w19928_,
		_w19931_,
		_w19933_
	);
	LUT2 #(
		.INIT('h1)
	) name19402 (
		\ld_r_reg/P0001 ,
		_w19932_,
		_w19934_
	);
	LUT2 #(
		.INIT('h4)
	) name19403 (
		_w19933_,
		_w19934_,
		_w19935_
	);
	LUT2 #(
		.INIT('h2)
	) name19404 (
		\text_in_r_reg[64]/P0001 ,
		\u0_w_reg[1][0]/P0001 ,
		_w19936_
	);
	LUT2 #(
		.INIT('h4)
	) name19405 (
		\text_in_r_reg[64]/P0001 ,
		\u0_w_reg[1][0]/P0001 ,
		_w19937_
	);
	LUT2 #(
		.INIT('h2)
	) name19406 (
		\ld_r_reg/P0001 ,
		_w19936_,
		_w19938_
	);
	LUT2 #(
		.INIT('h4)
	) name19407 (
		_w19937_,
		_w19938_,
		_w19939_
	);
	LUT2 #(
		.INIT('h1)
	) name19408 (
		_w19935_,
		_w19939_,
		_w19940_
	);
	LUT2 #(
		.INIT('h2)
	) name19409 (
		\u0_w_reg[2][0]/P0001 ,
		_w6657_,
		_w19941_
	);
	LUT2 #(
		.INIT('h4)
	) name19410 (
		\u0_w_reg[2][0]/P0001 ,
		_w6657_,
		_w19942_
	);
	LUT2 #(
		.INIT('h1)
	) name19411 (
		_w19941_,
		_w19942_,
		_w19943_
	);
	LUT2 #(
		.INIT('h8)
	) name19412 (
		_w6475_,
		_w7931_,
		_w19944_
	);
	LUT2 #(
		.INIT('h1)
	) name19413 (
		_w6475_,
		_w7931_,
		_w19945_
	);
	LUT2 #(
		.INIT('h1)
	) name19414 (
		_w19944_,
		_w19945_,
		_w19946_
	);
	LUT2 #(
		.INIT('h1)
	) name19415 (
		_w19943_,
		_w19946_,
		_w19947_
	);
	LUT2 #(
		.INIT('h8)
	) name19416 (
		_w19943_,
		_w19946_,
		_w19948_
	);
	LUT2 #(
		.INIT('h1)
	) name19417 (
		\ld_r_reg/P0001 ,
		_w19947_,
		_w19949_
	);
	LUT2 #(
		.INIT('h4)
	) name19418 (
		_w19948_,
		_w19949_,
		_w19950_
	);
	LUT2 #(
		.INIT('h2)
	) name19419 (
		\text_in_r_reg[32]/P0001 ,
		\u0_w_reg[2][0]/P0001 ,
		_w19951_
	);
	LUT2 #(
		.INIT('h4)
	) name19420 (
		\text_in_r_reg[32]/P0001 ,
		\u0_w_reg[2][0]/P0001 ,
		_w19952_
	);
	LUT2 #(
		.INIT('h2)
	) name19421 (
		\ld_r_reg/P0001 ,
		_w19951_,
		_w19953_
	);
	LUT2 #(
		.INIT('h4)
	) name19422 (
		_w19952_,
		_w19953_,
		_w19954_
	);
	LUT2 #(
		.INIT('h1)
	) name19423 (
		_w19950_,
		_w19954_,
		_w19955_
	);
	LUT2 #(
		.INIT('h1)
	) name19424 (
		\u0_w_reg[1][24]/P0002 ,
		_w16871_,
		_w19956_
	);
	LUT2 #(
		.INIT('h8)
	) name19425 (
		\u0_w_reg[1][24]/P0002 ,
		_w16871_,
		_w19957_
	);
	LUT2 #(
		.INIT('h1)
	) name19426 (
		ld_pad,
		_w19956_,
		_w19958_
	);
	LUT2 #(
		.INIT('h4)
	) name19427 (
		_w19957_,
		_w19958_,
		_w19959_
	);
	LUT2 #(
		.INIT('h8)
	) name19428 (
		\key[88]_pad ,
		ld_pad,
		_w19960_
	);
	LUT2 #(
		.INIT('h1)
	) name19429 (
		_w19959_,
		_w19960_,
		_w19961_
	);
	LUT2 #(
		.INIT('h4)
	) name19430 (
		_w15677_,
		_w15687_,
		_w19962_
	);
	LUT2 #(
		.INIT('h2)
	) name19431 (
		_w15677_,
		_w15687_,
		_w19963_
	);
	LUT2 #(
		.INIT('h1)
	) name19432 (
		ld_pad,
		_w19962_,
		_w19964_
	);
	LUT2 #(
		.INIT('h4)
	) name19433 (
		_w19963_,
		_w19964_,
		_w19965_
	);
	LUT2 #(
		.INIT('h8)
	) name19434 (
		\key[93]_pad ,
		ld_pad,
		_w19966_
	);
	LUT2 #(
		.INIT('h1)
	) name19435 (
		_w19965_,
		_w19966_,
		_w19967_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g21/_0_  = _w1315_ ;
	assign \g56610/_0_  = _w2092_ ;
	assign \g56611/_0_  = _w2544_ ;
	assign \g56612/_0_  = _w2957_ ;
	assign \g56613/_0_  = _w2978_ ;
	assign \g56614/_0_  = _w3090_ ;
	assign \g56615/_0_  = _w3108_ ;
	assign \g56616/_0_  = _w3220_ ;
	assign \g56617/_0_  = _w3238_ ;
	assign \g56630/_0_  = _w3783_ ;
	assign \g56631/_0_  = _w3801_ ;
	assign \g56632/_0_  = _w3981_ ;
	assign \g56633/_0_  = _w4086_ ;
	assign \g56634/_0_  = _w4263_ ;
	assign \g56635/_0_  = _w4362_ ;
	assign \g56645/_0_  = _w4593_ ;
	assign \g56646/_0_  = _w4689_ ;
	assign \g56647/_0_  = _w4707_ ;
	assign \g56648/_0_  = _w4728_ ;
	assign \g56649/_0_  = _w4746_ ;
	assign \g56650/_0_  = _w4770_ ;
	assign \g56651/_0_  = _w4797_ ;
	assign \g56652/_0_  = _w4884_ ;
	assign \g56666/_0_  = _w4899_ ;
	assign \g56667/_0_  = _w4923_ ;
	assign \g56668/_0_  = _w4938_ ;
	assign \g56669/_0_  = _w4956_ ;
	assign \g56670/_0_  = _w4974_ ;
	assign \g56671/_0_  = _w4992_ ;
	assign \g56672/_0_  = _w5007_ ;
	assign \g56674/_0_  = _w5025_ ;
	assign \g56675/_0_  = _w5040_ ;
	assign \g56704/_0_  = _w5055_ ;
	assign \g56739/_0_  = _w5058_ ;
	assign \g56743/_0_  = _w5061_ ;
	assign \g56763/_0_  = _w5064_ ;
	assign \g56776/_0_  = _w5067_ ;
	assign \g56812/_0_  = _w5070_ ;
	assign \g56818/_0_  = _w5073_ ;
	assign \g56861/_0_  = _w5076_ ;
	assign \g56874/_0_  = _w5079_ ;
	assign \g56919/_0_  = _w5322_ ;
	assign \g56920/_0_  = _w5646_ ;
	assign \g56921/_0_  = _w5949_ ;
	assign \g56923/_0_  = _w5967_ ;
	assign \g56924/_0_  = _w6076_ ;
	assign \g56925/_0_  = _w6195_ ;
	assign \g56926/_0_  = _w6213_ ;
	assign \g56956/_0_  = _w6758_ ;
	assign \g56957/_0_  = _w6942_ ;
	assign \g56958/_0_  = _w6960_ ;
	assign \g56959/_0_  = _w7130_ ;
	assign \g56960/_0_  = _w7233_ ;
	assign \g56961/_0_  = _w7334_ ;
	assign \g56972/_0_  = _w7435_ ;
	assign \g56973/_0_  = _w7670_ ;
	assign \g56974/_0_  = _w7691_ ;
	assign \g56976/_0_  = _w7709_ ;
	assign \g56977/_0_  = _w7733_ ;
	assign \g56978/_0_  = _w7751_ ;
	assign \g56979/_0_  = _w7775_ ;
	assign \g56980/_0_  = _w7871_ ;
	assign \g57008/_0_  = _w7886_ ;
	assign \g57010/_0_  = _w7907_ ;
	assign \g57011/_0_  = _w7925_ ;
	assign \g57012/_0_  = _w7943_ ;
	assign \g57013/_0_  = _w7961_ ;
	assign \g57014/_0_  = _w7979_ ;
	assign \g57015/_0_  = _w7994_ ;
	assign \g57016/_0_  = _w8012_ ;
	assign \g57017/_0_  = _w8030_ ;
	assign \g57086/_0_  = _w8033_ ;
	assign \g57091/_0_  = _w8036_ ;
	assign \g57114/_0_  = _w8039_ ;
	assign \g57129/_0_  = _w8042_ ;
	assign \g57163/_0_  = _w8045_ ;
	assign \g57171/_0_  = _w8048_ ;
	assign \g57204/_0_  = _w8051_ ;
	assign \g57218/_0_  = _w8054_ ;
	assign \g57262/_0_  = _w8868_ ;
	assign \g57263/_0_  = _w9304_ ;
	assign \g57264/_0_  = _w9418_ ;
	assign \g57265/_0_  = _w9537_ ;
	assign \g57266/_0_  = _w9654_ ;
	assign \g57267/_0_  = _w9675_ ;
	assign \g57268/_0_  = _w9693_ ;
	assign \g57269/_0_  = _w9995_ ;
	assign \g57300/_0_  = _w10523_ ;
	assign \g57301/_0_  = _w10697_ ;
	assign \g57302/_0_  = _w10799_ ;
	assign \g57303/_0_  = _w10817_ ;
	assign \g57304/_0_  = _w10919_ ;
	assign \g57316/_0_  = _w11173_ ;
	assign \g57317/_0_  = _w11399_ ;
	assign \g57319/_0_  = _w11420_ ;
	assign \g57320/_0_  = _w11438_ ;
	assign \g57321/_0_  = _w11465_ ;
	assign \g57322/_0_  = _w11486_ ;
	assign \g57323/_0_  = _w11580_ ;
	assign \g57324/_0_  = _w11601_ ;
	assign \g57350/_0_  = _w11619_ ;
	assign \g57353/_0_  = _w11637_ ;
	assign \g57354/_0_  = _w11658_ ;
	assign \g57355/_0_  = _w11676_ ;
	assign \g57356/_0_  = _w11694_ ;
	assign \g57357/_0_  = _w11712_ ;
	assign \g57358/_0_  = _w11730_ ;
	assign \g57359/_0_  = _w11748_ ;
	assign \g57360/_0_  = _w11766_ ;
	assign \g57427/_0_  = _w11769_ ;
	assign \g57432/_0_  = _w11772_ ;
	assign \g57456/_0_  = _w11775_ ;
	assign \g57471/_0_  = _w11778_ ;
	assign \g57506/_0_  = _w11781_ ;
	assign \g57512/_0_  = _w11784_ ;
	assign \g57540/_0_  = _w11787_ ;
	assign \g57547/_0_  = _w11790_ ;
	assign \g57654/_0_  = _w12595_ ;
	assign \g57655/_0_  = _w12848_ ;
	assign \g57656/_0_  = _w12977_ ;
	assign \g57657/_0_  = _w12995_ ;
	assign \g57658/_0_  = _w13299_ ;
	assign \g57676/_0_  = _w13937_ ;
	assign \g57677/_0_  = _w14225_ ;
	assign \g57678/_0_  = _w14415_ ;
	assign \g57679/_0_  = _w14816_ ;
	assign \g57680/_0_  = _w14985_ ;
	assign \g57681/_0_  = _w15083_ ;
	assign \g57682/_0_  = _w15101_ ;
	assign \g57683/_0_  = _w15122_ ;
	assign \g57684/_0_  = _w15143_ ;
	assign \g57685/_0_  = _w15161_ ;
	assign \g57686/_0_  = _w15176_ ;
	assign \g57687/_0_  = _w15194_ ;
	assign \g57688/_0_  = _w15218_ ;
	assign \g57689/_0_  = _w15304_ ;
	assign \g57690/_0_  = _w15322_ ;
	assign \g57691/_0_  = _w15346_ ;
	assign \g57700/_0_  = _w15361_ ;
	assign \g57701/_0_  = _w15379_ ;
	assign \g57702/_0_  = _w15397_ ;
	assign \g57703/_0_  = _w15412_ ;
	assign \g57704/_0_  = _w15433_ ;
	assign \g57705/_0_  = _w15448_ ;
	assign \g57706/_0_  = _w15466_ ;
	assign \g57707/_0_  = _w15484_ ;
	assign \g57708/_0_  = _w15502_ ;
	assign \g57709/_3_  = _w15683_ ;
	assign \g57710/_3_  = _w15695_ ;
	assign \g57711/_0_  = _w15701_ ;
	assign \g57712/_3_  = _w15888_ ;
	assign \g57715/_3_  = _w16009_ ;
	assign \g57716/_3_  = _w16198_ ;
	assign \g57767/_0_  = _w16216_ ;
	assign \g57768/_3_  = _w16336_ ;
	assign \g57769/_3_  = _w16345_ ;
	assign \g57770/_3_  = _w16351_ ;
	assign \g57771/_3_  = _w16357_ ;
	assign \g57777/_3_  = _w16474_ ;
	assign \g57779/_3_  = _w16647_ ;
	assign \g57804/_3_  = _w16772_ ;
	assign \g57805/_3_  = _w16873_ ;
	assign \g57806/_3_  = _w16970_ ;
	assign \g57807/_3_  = _w17056_ ;
	assign \g57808/_3_  = _w17149_ ;
	assign \g57809/_3_  = _w17158_ ;
	assign \g57810/_3_  = _w17167_ ;
	assign \g57811/_3_  = _w17176_ ;
	assign \g57812/_3_  = _w17188_ ;
	assign \g57813/_3_  = _w17197_ ;
	assign \g57814/_3_  = _w17206_ ;
	assign \g57815/_3_  = _w17215_ ;
	assign \g57816/_0_  = _w17224_ ;
	assign \g57817/_3_  = _w17230_ ;
	assign \g57818/_3_  = _w17236_ ;
	assign \g57819/_3_  = _w17242_ ;
	assign \g57822/_3_  = _w17245_ ;
	assign \g57823/_3_  = _w17251_ ;
	assign \g57824/_3_  = _w17257_ ;
	assign \g57830/_3_  = _w17369_ ;
	assign \g57835/_3_  = _w17372_ ;
	assign \g57836/_3_  = _w17378_ ;
	assign \g57837/_3_  = _w17384_ ;
	assign \g57841/_3_  = _w17387_ ;
	assign \g57842/_3_  = _w17393_ ;
	assign \g57843/_3_  = _w17399_ ;
	assign \g57854/_3_  = _w17494_ ;
	assign \g57855/_3_  = _w17596_ ;
	assign \g57856/_3_  = _w17704_ ;
	assign \g57857/_3_  = _w17801_ ;
	assign \g57858/_3_  = _w17894_ ;
	assign \g57859/_3_  = _w17991_ ;
	assign \g57860/_3_  = _w18077_ ;
	assign \g57861/_3_  = _w18161_ ;
	assign \g57871/_3_  = _w18263_ ;
	assign \g57872/_3_  = _w18364_ ;
	assign \g57874/_3_  = _w18445_ ;
	assign \g57968/_3_  = _w18533_ ;
	assign \g57969/_3_  = _w18542_ ;
	assign \g57970/_3_  = _w18551_ ;
	assign \g57971/_3_  = _w18557_ ;
	assign \g57980/_3_  = _w18654_ ;
	assign \g57983/_3_  = _w18657_ ;
	assign \g57984/_3_  = _w18663_ ;
	assign \g57985/_3_  = _w18669_ ;
	assign \g58012/_3_  = _w18672_ ;
	assign \g58013/_3_  = _w18678_ ;
	assign \g58015/_3_  = _w18684_ ;
	assign \g58057/_3_  = _w18773_ ;
	assign \g58058/_3_  = _w18862_ ;
	assign \g58059/_3_  = _w18953_ ;
	assign \g58189/_3_  = _w18956_ ;
	assign \g58190/_3_  = _w18962_ ;
	assign \g58191/_3_  = _w19048_ ;
	assign \g58192/_3_  = _w19138_ ;
	assign \g58193/_3_  = _w19144_ ;
	assign \g58194/_3_  = _w19234_ ;
	assign \g58195/_3_  = _w19240_ ;
	assign \g58196/_3_  = _w19252_ ;
	assign \g58197/_3_  = _w19261_ ;
	assign \g58224/_3_  = _w19264_ ;
	assign \g58226/_3_  = _w19270_ ;
	assign \g58229/_3_  = _w19276_ ;
	assign \g58255/_3_  = _w19279_ ;
	assign \g58256/_3_  = _w19282_ ;
	assign \g58257/_3_  = _w19285_ ;
	assign \g58258/_3_  = _w19288_ ;
	assign \g58259/_3_  = _w19291_ ;
	assign \g58260/_3_  = _w19297_ ;
	assign \g58261/_3_  = _w19303_ ;
	assign \g58262/_3_  = _w19309_ ;
	assign \g58263/_3_  = _w19315_ ;
	assign \g58264/_3_  = _w19318_ ;
	assign \g58265/_3_  = _w19324_ ;
	assign \g58266/_3_  = _w19330_ ;
	assign \g58267/_3_  = _w19336_ ;
	assign \g58268/_3_  = _w19342_ ;
	assign \g58269/_3_  = _w19348_ ;
	assign \g58270/_0_  = _w19351_ ;
	assign \g58271/_3_  = _w19354_ ;
	assign \g58272/_3_  = _w19357_ ;
	assign \g58273/_3_  = _w19360_ ;
	assign \g58274/_3_  = _w19366_ ;
	assign \g58275/_3_  = _w19372_ ;
	assign \g58276/_3_  = _w19378_ ;
	assign \g58277/_3_  = _w19384_ ;
	assign \g58278/_3_  = _w19390_ ;
	assign \g58279/_3_  = _w19396_ ;
	assign \g58285/_3_  = _w19399_ ;
	assign \g58286/_3_  = _w19402_ ;
	assign \g58288/_3_  = _w19405_ ;
	assign \g58289/_3_  = _w19411_ ;
	assign \g58290/_3_  = _w19414_ ;
	assign \g58292/_3_  = _w19420_ ;
	assign \g58294/_3_  = _w19426_ ;
	assign \g58295/_3_  = _w19432_ ;
	assign \g58297/_3_  = _w19438_ ;
	assign \g58330/_0_  = _w19441_ ;
	assign \g58331/_0_  = _w19444_ ;
	assign \g58332/_0_  = _w19447_ ;
	assign \g58333/_0_  = _w19450_ ;
	assign \g58444/_3_  = _w19453_ ;
	assign \g58445/_3_  = _w19456_ ;
	assign \g58446/_3_  = _w19462_ ;
	assign \g58462/_0_  = _w19465_ ;
	assign \g58506/_0_  = _w19468_ ;
	assign \g58507/_0_  = _w19471_ ;
	assign \g58508/_0_  = _w19474_ ;
	assign \g58509/_0_  = _w19477_ ;
	assign \g58531/_0_  = _w19480_ ;
	assign \g58532/_0_  = _w19483_ ;
	assign \g58533/_0_  = _w19486_ ;
	assign \g58550/_0_  = _w19489_ ;
	assign \g58551/_0_  = _w19492_ ;
	assign \g58552/_0_  = _w19495_ ;
	assign \g58553/_0_  = _w19498_ ;
	assign \g58554/_0_  = _w19501_ ;
	assign \g58555/_0_  = _w19504_ ;
	assign \g58556/_0_  = _w19507_ ;
	assign \g58557/_0_  = _w19510_ ;
	assign \g58558/_0_  = _w19513_ ;
	assign \g58559/_0_  = _w19516_ ;
	assign \g58560/_0_  = _w19519_ ;
	assign \g58600/_3_  = _w19522_ ;
	assign \g58601/_3_  = _w19525_ ;
	assign \g58602/_3_  = _w19528_ ;
	assign \g58603/_3_  = _w19534_ ;
	assign \g58604/_3_  = _w19540_ ;
	assign \g58605/_3_  = _w19546_ ;
	assign \g58606/_3_  = _w19552_ ;
	assign \g58607/_3_  = _w19558_ ;
	assign \g58608/_3_  = _w19564_ ;
	assign \g58611/_0_  = _w19567_ ;
	assign \g58612/_0_  = _w19570_ ;
	assign \g58613/_0_  = _w19573_ ;
	assign \g58614/_0_  = _w19576_ ;
	assign \g58617/_0_  = _w19579_ ;
	assign \g58618/_0_  = _w19582_ ;
	assign \g58619/_0_  = _w19585_ ;
	assign \g58634/_0_  = _w19588_ ;
	assign \g58635/_0_  = _w19591_ ;
	assign \g58636/_0_  = _w19594_ ;
	assign \g58637/_0_  = _w19597_ ;
	assign \g58638/_0_  = _w19600_ ;
	assign \g58639/_0_  = _w19603_ ;
	assign \g58640/_0_  = _w19606_ ;
	assign \g58641/_0_  = _w19609_ ;
	assign \g58829/_3_  = _w19612_ ;
	assign \g58830/_3_  = _w19615_ ;
	assign \g58831/_3_  = _w19618_ ;
	assign \g58832/_3_  = _w19624_ ;
	assign \g58833/_3_  = _w19630_ ;
	assign \g58834/_3_  = _w19636_ ;
	assign \g58835/_0_  = _w19639_ ;
	assign \g58844/_0_  = _w19642_ ;
	assign \g58902/_0_  = _w19645_ ;
	assign \g58903/_0_  = _w19648_ ;
	assign \g58904/_0_  = _w19651_ ;
	assign \g58905/_0_  = _w19654_ ;
	assign \g58910/_0_  = _w19657_ ;
	assign \g58913/_0_  = _w19660_ ;
	assign \g58934/_0_  = _w19663_ ;
	assign \g58935/_0_  = _w19666_ ;
	assign \g58936/_0_  = _w19669_ ;
	assign \g58937/_0_  = _w19672_ ;
	assign \g58938/_0_  = _w19675_ ;
	assign \g58970/_0_  = _w19678_ ;
	assign \g58972/_0_  = _w19681_ ;
	assign \g58994/_0_  = _w19684_ ;
	assign \g58995/_0_  = _w19687_ ;
	assign \g58996/_0_  = _w19690_ ;
	assign \g58997/_0_  = _w19693_ ;
	assign \g58998/_0_  = _w19696_ ;
	assign \g58999/_0_  = _w19699_ ;
	assign \g59000/_0_  = _w19702_ ;
	assign \g59002/_0_  = _w19705_ ;
	assign \g59003/_0_  = _w19708_ ;
	assign \g59004/_0_  = _w19711_ ;
	assign \g59254/_0_  = _w19714_ ;
	assign \g59257/_0_  = _w19717_ ;
	assign \g59258/_0_  = _w19720_ ;
	assign \g59259/_0_  = _w19723_ ;
	assign \g59276/_0_  = _w19726_ ;
	assign \g59277/_0_  = _w19729_ ;
	assign \g59278/_0_  = _w19732_ ;
	assign \g59279/_0_  = _w19735_ ;
	assign \g59280/_0_  = _w19738_ ;
	assign \g59291/_0_  = _w19741_ ;
	assign \g59292/_0_  = _w19744_ ;
	assign \g59293/_0_  = _w19747_ ;
	assign \g59294/_0_  = _w19750_ ;
	assign \g59295/_0_  = _w19753_ ;
	assign \g59308/_0_  = _w19756_ ;
	assign \g59309/_0_  = _w19759_ ;
	assign \g59310/_0_  = _w19762_ ;
	assign \g59311/_0_  = _w19765_ ;
	assign \g59330/_0_  = _w19768_ ;
	assign \g59331/_0_  = _w19771_ ;
	assign \g59332/_0_  = _w19774_ ;
	assign \g59333/_0_  = _w19777_ ;
	assign \g59334/_0_  = _w19780_ ;
	assign \g59335/_0_  = _w19783_ ;
	assign \g59336/_0_  = _w19786_ ;
	assign \g59337/_0_  = _w19789_ ;
	assign \g59338/_0_  = _w19792_ ;
	assign \g59339/_0_  = _w19795_ ;
	assign \g59596/_0_  = _w19798_ ;
	assign \g59597/_0_  = _w19801_ ;
	assign \g59598/_0_  = _w19804_ ;
	assign \g59599/_0_  = _w19807_ ;
	assign \g59625/_0_  = _w19810_ ;
	assign \g59626/_0_  = _w19813_ ;
	assign \g59627/_0_  = _w19816_ ;
	assign \g59628/_0_  = _w19819_ ;
	assign \g59837/_0_  = _w19822_ ;
	assign \g59838/_0_  = _w19825_ ;
	assign \g59839/_0_  = _w19828_ ;
	assign \g59840/_0_  = _w19831_ ;
	assign \g60090/_0_  = _w19848_ ;
	assign \g60320/_0_  = _w19852_ ;
	assign \g60321/_0_  = _w19856_ ;
	assign \g60409/_0_  = _w19858_ ;
	assign \g60539/_0_  = _w19861_ ;
	assign \g60860/_0_  = _w19864_ ;
	assign \g60977/_0_  = _w19866_ ;
	assign \g61012/_0_  = _w19871_ ;
	assign \g61185/_0_  = _w19872_ ;
	assign \g61524/_2_  = _w19873_ ;
	assign \g61776/_0_  = _w19878_ ;
	assign \g61895/_0_  = _w19884_ ;
	assign \g61897/_0_  = _w19888_ ;
	assign \g62220/_0_  = _w19889_ ;
	assign \g65958/_0_  = _w19862_ ;
	assign \g72347/_3_  = _w19892_ ;
	assign \g77848/_0_  = _w19857_ ;
	assign \g85056/_0_  = _w19910_ ;
	assign \sa30_reg[0]/_05_  = _w19925_ ;
	assign \sa31_reg[0]/_05_  = _w19940_ ;
	assign \sa32_reg[0]/_05_  = _w19955_ ;
	assign \u0_w_reg[1][24]/_05_  = _w19961_ ;
	assign \u0_w_reg[1][29]/_05_  = _w19967_ ;
endmodule;