module top (\G0_pad , \G10_pad , \G11_pad , \G12_pad , \G13_pad , \G1_pad , \G29_reg/NET0131 , \G2_pad , \G30_reg/NET0131 , \G31_reg/NET0131 , \G32_reg/NET0131 , \G33_reg/NET0131 , \G34_reg/NET0131 , \G35_reg/NET0131 , \G36_reg/NET0131 , \G37_reg/NET0131 , \G38_reg/NET0131 , \G39_reg/NET0131 , \G3_pad , \G40_reg/NET0131 , \G41_reg/NET0131 , \G42_reg/NET0131 , \G43_reg/NET0131 , \G44_reg/NET0131 , \G46_reg/NET0131 , \G4_pad , \G5_pad , \G6_pad , \G7_pad , \G8_pad , \G9_pad , \G532_pad , \G537_pad , \G539_pad , \G542_pad , \G546_pad , \G547_pad , \G548_pad , \G549_pad , \G550_pad , \G551_pad , \G552_pad , \_al_n0 , \_al_n1 , \g1667/_3_ , \g1737/_0_ , \g1744/_0_ , \g1787/_0_ , \g1811/_0_ , \g1830/_0_ , \g1831/_0_ , \g1846/_0_ , \g1852/_0_ , \g1866/_0_ , \g19/_2_ , \g1931/_0_ , \g1945/_0_ , \g2014/_0_ , \g2015/_0_ , \g2643/_0_ , \g2859/_1_ , \g3397/_2_ , \g3546/_0_ , \g3606/_3_ );
	input \G0_pad  ;
	input \G10_pad  ;
	input \G11_pad  ;
	input \G12_pad  ;
	input \G13_pad  ;
	input \G1_pad  ;
	input \G29_reg/NET0131  ;
	input \G2_pad  ;
	input \G30_reg/NET0131  ;
	input \G31_reg/NET0131  ;
	input \G32_reg/NET0131  ;
	input \G33_reg/NET0131  ;
	input \G34_reg/NET0131  ;
	input \G35_reg/NET0131  ;
	input \G36_reg/NET0131  ;
	input \G37_reg/NET0131  ;
	input \G38_reg/NET0131  ;
	input \G39_reg/NET0131  ;
	input \G3_pad  ;
	input \G40_reg/NET0131  ;
	input \G41_reg/NET0131  ;
	input \G42_reg/NET0131  ;
	input \G43_reg/NET0131  ;
	input \G44_reg/NET0131  ;
	input \G46_reg/NET0131  ;
	input \G4_pad  ;
	input \G5_pad  ;
	input \G6_pad  ;
	input \G7_pad  ;
	input \G8_pad  ;
	input \G9_pad  ;
	output \G532_pad  ;
	output \G537_pad  ;
	output \G539_pad  ;
	output \G542_pad  ;
	output \G546_pad  ;
	output \G547_pad  ;
	output \G548_pad  ;
	output \G549_pad  ;
	output \G550_pad  ;
	output \G551_pad  ;
	output \G552_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1667/_3_  ;
	output \g1737/_0_  ;
	output \g1744/_0_  ;
	output \g1787/_0_  ;
	output \g1811/_0_  ;
	output \g1830/_0_  ;
	output \g1831/_0_  ;
	output \g1846/_0_  ;
	output \g1852/_0_  ;
	output \g1866/_0_  ;
	output \g19/_2_  ;
	output \g1931/_0_  ;
	output \g1945/_0_  ;
	output \g2014/_0_  ;
	output \g2015/_0_  ;
	output \g2643/_0_  ;
	output \g2859/_1_  ;
	output \g3397/_2_  ;
	output \g3546/_0_  ;
	output \g3606/_3_  ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\G7_pad ,
		\G8_pad ,
		_w32_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\G30_reg/NET0131 ,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\G11_pad ,
		\G9_pad ,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\G8_pad ,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\G10_pad ,
		\G7_pad ,
		_w36_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		_w35_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		\G10_pad ,
		\G9_pad ,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\G7_pad ,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w33_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		_w37_,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h2)
	) name10 (
		\G32_reg/NET0131 ,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		\G13_pad ,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		\G5_pad ,
		\G6_pad ,
		_w44_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\G3_pad ,
		\G4_pad ,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w44_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\G11_pad ,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\G7_pad ,
		\G8_pad ,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\G8_pad ,
		\G9_pad ,
		_w49_
	);
	LUT2 #(
		.INIT('h2)
	) name18 (
		\G10_pad ,
		\G9_pad ,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		\G10_pad ,
		\G7_pad ,
		_w51_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w48_,
		_w49_,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w50_,
		_w51_,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		_w52_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		\G7_pad ,
		_w38_,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\G8_pad ,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		_w54_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		_w47_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		\G36_reg/NET0131 ,
		\G6_pad ,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		\G4_pad ,
		\G6_pad ,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\G5_pad ,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\G11_pad ,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w54_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		_w59_,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\G3_pad ,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		_w58_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		\G2_pad ,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w43_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\G3_pad ,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		\G1_pad ,
		\G2_pad ,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\G3_pad ,
		\G5_pad ,
		_w71_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		\G4_pad ,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name41 (
		\G2_pad ,
		\G3_pad ,
		_w73_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		\G2_pad ,
		\G3_pad ,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w73_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		_w72_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		\G6_pad ,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		\G4_pad ,
		\G5_pad ,
		_w78_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		\G3_pad ,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w77_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h2)
	) name49 (
		\G1_pad ,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		\G4_pad ,
		\G6_pad ,
		_w82_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		\G5_pad ,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		_w70_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\G1_pad ,
		\G3_pad ,
		_w85_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		\G5_pad ,
		_w60_,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		_w85_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		\G1_pad ,
		\G4_pad ,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		\G5_pad ,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h2)
	) name58 (
		\G1_pad ,
		\G4_pad ,
		_w90_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		\G2_pad ,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		\G6_pad ,
		_w89_,
		_w92_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		_w91_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		_w84_,
		_w87_,
		_w94_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		_w93_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		_w81_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		_w41_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		\G11_pad ,
		\G9_pad ,
		_w98_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		\G10_pad ,
		\G7_pad ,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		\G8_pad ,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		_w98_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		\G7_pad ,
		\G8_pad ,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\G10_pad ,
		_w34_,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		_w102_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w101_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\G3_pad ,
		\G6_pad ,
		_w106_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		\G1_pad ,
		\G4_pad ,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w90_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		_w106_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		_w105_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		\G1_pad ,
		\G3_pad ,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		_w51_,
		_w60_,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		_w35_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		\G8_pad ,
		_w99_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		\G4_pad ,
		\G6_pad ,
		_w115_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		_w98_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		_w114_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		_w113_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h2)
	) name87 (
		_w111_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		_w110_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h2)
	) name89 (
		\G2_pad ,
		\G5_pad ,
		_w121_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		_w120_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		\G10_pad ,
		\G11_pad ,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		_w102_,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		\G9_pad ,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		_w35_,
		_w36_,
		_w126_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w125_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		_w60_,
		_w71_,
		_w128_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		_w127_,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		\G1_pad ,
		\G2_pad ,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w129_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w122_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w97_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		\G13_pad ,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		_w70_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		_w69_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		\G6_pad ,
		_w78_,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w104_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h4)
	) name107 (
		_w136_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name108 (
		\G13_pad ,
		\G43_reg/NET0131 ,
		_w140_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		_w97_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		_w61_,
		_w101_,
		_w142_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		\G36_reg/NET0131 ,
		_w115_,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		_w142_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		\G3_pad ,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		_w68_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		\G4_pad ,
		\G5_pad ,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		\G11_pad ,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\G35_reg/NET0131 ,
		\G3_pad ,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w148_,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w129_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		\G2_pad ,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w67_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		_w43_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		\G13_pad ,
		\G1_pad ,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w133_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w154_,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		\G4_pad ,
		\G5_pad ,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		_w125_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		_w54_,
		_w148_,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w159_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		\G2_pad ,
		_w106_,
		_w162_
	);
	LUT2 #(
		.INIT('h4)
	) name131 (
		_w161_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		_w157_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		_w141_,
		_w146_,
		_w165_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		_w164_,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w139_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		\G12_pad ,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h2)
	) name137 (
		\G12_pad ,
		\G13_pad ,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		\G0_pad ,
		\G3_pad ,
		_w170_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		\G3_pad ,
		\G5_pad ,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		\G4_pad ,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h4)
	) name141 (
		_w170_,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		\G31_reg/NET0131 ,
		\G8_pad ,
		_w174_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		\G10_pad ,
		\G8_pad ,
		_w175_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		\G7_pad ,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h2)
	) name145 (
		\G9_pad ,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h4)
	) name146 (
		\G6_pad ,
		\G7_pad ,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		\G30_reg/NET0131 ,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		\G10_pad ,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		\G9_pad ,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		_w174_,
		_w177_,
		_w182_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		_w181_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		\G11_pad ,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		\G30_reg/NET0131 ,
		\G6_pad ,
		_w185_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		\G31_reg/NET0131 ,
		_w179_,
		_w186_
	);
	LUT2 #(
		.INIT('h2)
	) name155 (
		\G8_pad ,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		\G10_pad ,
		\G8_pad ,
		_w188_
	);
	LUT2 #(
		.INIT('h2)
	) name157 (
		\G9_pad ,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		_w48_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		_w187_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h2)
	) name160 (
		\G11_pad ,
		_w185_,
		_w192_
	);
	LUT2 #(
		.INIT('h4)
	) name161 (
		_w191_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		_w184_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h2)
	) name163 (
		\G46_reg/NET0131 ,
		_w173_,
		_w195_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		_w194_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		_w169_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h2)
	) name166 (
		\G3_pad ,
		\G4_pad ,
		_w198_
	);
	LUT2 #(
		.INIT('h4)
	) name167 (
		\G2_pad ,
		\G5_pad ,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		_w198_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h2)
	) name169 (
		\G1_pad ,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		\G3_pad ,
		\G5_pad ,
		_w202_
	);
	LUT2 #(
		.INIT('h2)
	) name171 (
		\G2_pad ,
		_w85_,
		_w203_
	);
	LUT2 #(
		.INIT('h4)
	) name172 (
		\G2_pad ,
		_w71_,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		_w202_,
		_w203_,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name174 (
		_w204_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h2)
	) name175 (
		\G4_pad ,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		_w201_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h2)
	) name177 (
		\G0_pad ,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		_w197_,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		_w168_,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h4)
	) name180 (
		\G5_pad ,
		_w115_,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		_w123_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		_w61_,
		_w103_,
		_w214_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		_w213_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h2)
	) name184 (
		_w102_,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h4)
	) name185 (
		\G6_pad ,
		_w36_,
		_w217_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		_w35_,
		_w78_,
		_w218_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		_w217_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		_w216_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		\G3_pad ,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		_w46_,
		_w54_,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name191 (
		\G11_pad ,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		_w221_,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		\G12_pad ,
		_w68_,
		_w225_
	);
	LUT2 #(
		.INIT('h4)
	) name194 (
		_w224_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		\G11_pad ,
		\G2_pad ,
		_w227_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\G6_pad ,
		\G9_pad ,
		_w228_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		\G4_pad ,
		_w36_,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		_w228_,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w71_,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h4)
	) name200 (
		\G9_pad ,
		_w99_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		_w106_,
		_w147_,
		_w233_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		_w232_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		_w231_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h2)
	) name204 (
		\G8_pad ,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		_w157_,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h4)
	) name206 (
		\G1_pad ,
		_w134_,
		_w238_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		_w222_,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		_w237_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		\G12_pad ,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h2)
	) name210 (
		_w169_,
		_w196_,
		_w242_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		\G0_pad ,
		\G4_pad ,
		_w243_
	);
	LUT2 #(
		.INIT('h2)
	) name212 (
		\G6_pad ,
		\G9_pad ,
		_w244_
	);
	LUT2 #(
		.INIT('h2)
	) name213 (
		\G11_pad ,
		\G7_pad ,
		_w245_
	);
	LUT2 #(
		.INIT('h2)
	) name214 (
		\G10_pad ,
		\G8_pad ,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		_w202_,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		_w244_,
		_w245_,
		_w248_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		_w247_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		\G11_pad ,
		\G37_reg/NET0131 ,
		_w250_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		_w71_,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		_w100_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		_w249_,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		_w243_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		_w61_,
		_w170_,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		_w126_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w254_,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h2)
	) name226 (
		_w130_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		_w242_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		\G0_pad ,
		_w230_,
		_w260_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		\G38_reg/NET0131 ,
		_w244_,
		_w261_
	);
	LUT2 #(
		.INIT('h1)
	) name230 (
		_w260_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		\G1_pad ,
		\G8_pad ,
		_w263_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		_w71_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		_w262_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		_w259_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		_w241_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h2)
	) name236 (
		_w227_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w226_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h2)
	) name238 (
		_w242_,
		_w258_,
		_w270_
	);
	LUT2 #(
		.INIT('h4)
	) name239 (
		\G12_pad ,
		\G13_pad ,
		_w271_
	);
	LUT2 #(
		.INIT('h4)
	) name240 (
		_w97_,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w132_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h4)
	) name242 (
		\G12_pad ,
		_w43_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name243 (
		_w153_,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w270_,
		_w273_,
		_w276_
	);
	LUT2 #(
		.INIT('h4)
	) name245 (
		_w275_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		\G34_reg/NET0131 ,
		_w36_,
		_w278_
	);
	LUT2 #(
		.INIT('h4)
	) name247 (
		_w49_,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		\G34_reg/NET0131 ,
		\G8_pad ,
		_w280_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		\G6_pad ,
		_w197_,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		_w280_,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		_w39_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h2)
	) name252 (
		\G11_pad ,
		_w48_,
		_w284_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		\G9_pad ,
		_w123_,
		_w285_
	);
	LUT2 #(
		.INIT('h4)
	) name254 (
		_w284_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		\G7_pad ,
		\G9_pad ,
		_w287_
	);
	LUT2 #(
		.INIT('h2)
	) name256 (
		_w188_,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h4)
	) name257 (
		\G8_pad ,
		_w103_,
		_w289_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		_w286_,
		_w288_,
		_w290_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		_w289_,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h2)
	) name260 (
		_w281_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w279_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h4)
	) name262 (
		_w283_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		_w197_,
		_w217_,
		_w295_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		\G8_pad ,
		_w36_,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		\G7_pad ,
		_w188_,
		_w297_
	);
	LUT2 #(
		.INIT('h2)
	) name266 (
		\G34_reg/NET0131 ,
		_w296_,
		_w298_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		_w297_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w295_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h2)
	) name269 (
		\G9_pad ,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		_w34_,
		_w38_,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		\G8_pad ,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h2)
	) name272 (
		_w32_,
		_w50_,
		_w304_
	);
	LUT2 #(
		.INIT('h4)
	) name273 (
		_w123_,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		_w39_,
		_w303_,
		_w306_
	);
	LUT2 #(
		.INIT('h4)
	) name275 (
		_w305_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h2)
	) name276 (
		_w281_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		_w301_,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h4)
	) name278 (
		\G42_reg/NET0131 ,
		_w197_,
		_w310_
	);
	LUT2 #(
		.INIT('h2)
	) name279 (
		\G7_pad ,
		_w50_,
		_w311_
	);
	LUT2 #(
		.INIT('h4)
	) name280 (
		_w189_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		\G11_pad ,
		\G34_reg/NET0131 ,
		_w313_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		_w102_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		_w55_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h4)
	) name284 (
		_w312_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		_w310_,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		_w97_,
		_w271_,
		_w318_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		\G1_pad ,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h4)
	) name288 (
		\G3_pad ,
		_w60_,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w74_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h2)
	) name290 (
		\G5_pad ,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		\G2_pad ,
		\G4_pad ,
		_w323_
	);
	LUT2 #(
		.INIT('h4)
	) name292 (
		\G5_pad ,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h4)
	) name293 (
		\G2_pad ,
		\G6_pad ,
		_w325_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		\G5_pad ,
		\G6_pad ,
		_w326_
	);
	LUT2 #(
		.INIT('h1)
	) name295 (
		_w106_,
		_w325_,
		_w327_
	);
	LUT2 #(
		.INIT('h4)
	) name296 (
		_w326_,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h1)
	) name297 (
		_w71_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		\G4_pad ,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		_w322_,
		_w324_,
		_w331_
	);
	LUT2 #(
		.INIT('h4)
	) name300 (
		_w330_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h2)
	) name301 (
		_w319_,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h2)
	) name302 (
		_w88_,
		_w170_,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		_w197_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		\G13_pad ,
		\G33_reg/NET0131 ,
		_w336_
	);
	LUT2 #(
		.INIT('h8)
	) name305 (
		\G3_pad ,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		\G2_pad ,
		\G5_pad ,
		_w338_
	);
	LUT2 #(
		.INIT('h4)
	) name307 (
		\G12_pad ,
		_w42_,
		_w339_
	);
	LUT2 #(
		.INIT('h4)
	) name308 (
		\G13_pad ,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h4)
	) name309 (
		_w45_,
		_w338_,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name310 (
		_w340_,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		_w337_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h4)
	) name312 (
		_w335_,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h4)
	) name313 (
		_w333_,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h2)
	) name314 (
		\G0_pad ,
		\G29_reg/NET0131 ,
		_w346_
	);
	LUT2 #(
		.INIT('h4)
	) name315 (
		\G0_pad ,
		_w88_,
		_w347_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		\G3_pad ,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w346_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h2)
	) name318 (
		_w197_,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h2)
	) name319 (
		_w71_,
		_w323_,
		_w351_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		_w340_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		\G5_pad ,
		_w88_,
		_w353_
	);
	LUT2 #(
		.INIT('h2)
	) name322 (
		\G2_pad ,
		_w89_,
		_w354_
	);
	LUT2 #(
		.INIT('h4)
	) name323 (
		_w353_,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		_w318_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		_w337_,
		_w352_,
		_w357_
	);
	LUT2 #(
		.INIT('h4)
	) name326 (
		_w350_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h4)
	) name327 (
		_w356_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		_w88_,
		_w170_,
		_w360_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		\G0_pad ,
		\G2_pad ,
		_w361_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		\G1_pad ,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h4)
	) name331 (
		\G4_pad ,
		_w361_,
		_w363_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		\G3_pad ,
		_w362_,
		_w364_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		_w363_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		_w347_,
		_w360_,
		_w366_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		_w365_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h2)
	) name336 (
		_w197_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		\G2_pad ,
		_w85_,
		_w369_
	);
	LUT2 #(
		.INIT('h2)
	) name338 (
		\G4_pad ,
		_w130_,
		_w370_
	);
	LUT2 #(
		.INIT('h4)
	) name339 (
		_w369_,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		_w318_,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		_w368_,
		_w372_,
		_w373_
	);
	LUT2 #(
		.INIT('h2)
	) name342 (
		\G5_pad ,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h4)
	) name343 (
		_w74_,
		_w78_,
		_w375_
	);
	LUT2 #(
		.INIT('h8)
	) name344 (
		_w44_,
		_w74_,
		_w376_
	);
	LUT2 #(
		.INIT('h1)
	) name345 (
		_w320_,
		_w375_,
		_w377_
	);
	LUT2 #(
		.INIT('h4)
	) name346 (
		_w376_,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h2)
	) name347 (
		_w319_,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h8)
	) name348 (
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w380_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		_w340_,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		_w379_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name351 (
		_w374_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h4)
	) name352 (
		\G1_pad ,
		\G5_pad ,
		_w384_
	);
	LUT2 #(
		.INIT('h2)
	) name353 (
		\G4_pad ,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h2)
	) name354 (
		_w203_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h4)
	) name355 (
		\G4_pad ,
		\G5_pad ,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		_w85_,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		_w386_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h2)
	) name358 (
		_w318_,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h2)
	) name359 (
		_w74_,
		_w78_,
		_w391_
	);
	LUT2 #(
		.INIT('h2)
	) name360 (
		\G2_pad ,
		_w147_,
		_w392_
	);
	LUT2 #(
		.INIT('h8)
	) name361 (
		\G5_pad ,
		_w45_,
		_w393_
	);
	LUT2 #(
		.INIT('h2)
	) name362 (
		_w392_,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		_w391_,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h2)
	) name364 (
		_w340_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		_w390_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h2)
	) name366 (
		\G6_pad ,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h4)
	) name367 (
		\G40_reg/NET0131 ,
		_w197_,
		_w399_
	);
	LUT2 #(
		.INIT('h2)
	) name368 (
		_w60_,
		_w338_,
		_w400_
	);
	LUT2 #(
		.INIT('h8)
	) name369 (
		_w319_,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		_w399_,
		_w401_,
		_w402_
	);
	LUT2 #(
		.INIT('h4)
	) name371 (
		_w398_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h8)
	) name372 (
		_w65_,
		_w225_,
		_w404_
	);
	LUT2 #(
		.INIT('h2)
	) name373 (
		\G0_pad ,
		_w198_,
		_w405_
	);
	LUT2 #(
		.INIT('h4)
	) name374 (
		\G0_pad ,
		_w172_,
		_w406_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		\G1_pad ,
		_w405_,
		_w407_
	);
	LUT2 #(
		.INIT('h4)
	) name376 (
		_w406_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		_w72_,
		_w384_,
		_w409_
	);
	LUT2 #(
		.INIT('h2)
	) name378 (
		\G0_pad ,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		_w408_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h2)
	) name380 (
		\G2_pad ,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h8)
	) name381 (
		_w197_,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		_w404_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h2)
	) name383 (
		\G3_pad ,
		_w78_,
		_w415_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		_w338_,
		_w375_,
		_w416_
	);
	LUT2 #(
		.INIT('h4)
	) name385 (
		_w415_,
		_w416_,
		_w417_
	);
	LUT2 #(
		.INIT('h2)
	) name386 (
		\G0_pad ,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		\G1_pad ,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		\G10_pad ,
		\G30_reg/NET0131 ,
		_w420_
	);
	LUT2 #(
		.INIT('h2)
	) name389 (
		\G7_pad ,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h1)
	) name390 (
		\G6_pad ,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h2)
	) name391 (
		_w111_,
		_w387_,
		_w423_
	);
	LUT2 #(
		.INIT('h4)
	) name392 (
		_w78_,
		_w405_,
		_w424_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		_w423_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h8)
	) name394 (
		\G2_pad ,
		_w409_,
		_w426_
	);
	LUT2 #(
		.INIT('h4)
	) name395 (
		_w425_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		_w422_,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h4)
	) name397 (
		_w419_,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		_w318_,
		_w340_,
		_w430_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		\G11_pad ,
		\G7_pad ,
		_w431_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		\G10_pad ,
		\G11_pad ,
		_w432_
	);
	LUT2 #(
		.INIT('h2)
	) name401 (
		\G9_pad ,
		_w431_,
		_w433_
	);
	LUT2 #(
		.INIT('h4)
	) name402 (
		_w432_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		\G31_reg/NET0131 ,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h2)
	) name404 (
		\G6_pad ,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w179_,
		_w436_,
		_w437_
	);
	LUT2 #(
		.INIT('h2)
	) name406 (
		\G8_pad ,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('h4)
	) name407 (
		_w36_,
		_w228_,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name408 (
		\G6_pad ,
		_w188_,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name409 (
		_w48_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		\G9_pad ,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h4)
	) name411 (
		_w38_,
		_w178_,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name412 (
		_w439_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h4)
	) name413 (
		_w442_,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h2)
	) name414 (
		\G11_pad ,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name415 (
		_w86_,
		_w325_,
		_w447_
	);
	LUT2 #(
		.INIT('h4)
	) name416 (
		_w324_,
		_w447_,
		_w448_
	);
	LUT2 #(
		.INIT('h2)
	) name417 (
		\G1_pad ,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h1)
	) name418 (
		_w84_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h2)
	) name419 (
		\G3_pad ,
		_w450_,
		_w451_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		_w126_,
		_w212_,
		_w452_
	);
	LUT2 #(
		.INIT('h8)
	) name421 (
		_w61_,
		_w104_,
		_w453_
	);
	LUT2 #(
		.INIT('h4)
	) name422 (
		\G9_pad ,
		_w326_,
		_w454_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		_w124_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h1)
	) name424 (
		_w452_,
		_w455_,
		_w456_
	);
	LUT2 #(
		.INIT('h4)
	) name425 (
		_w453_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h1)
	) name426 (
		_w124_,
		_w126_,
		_w458_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		\G5_pad ,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h2)
	) name428 (
		_w74_,
		_w83_,
		_w460_
	);
	LUT2 #(
		.INIT('h4)
	) name429 (
		_w128_,
		_w392_,
		_w461_
	);
	LUT2 #(
		.INIT('h1)
	) name430 (
		_w460_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		_w45_,
		_w387_,
		_w463_
	);
	LUT2 #(
		.INIT('h2)
	) name432 (
		_w70_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		_w391_,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		_w99_,
		_w243_,
		_w466_
	);
	LUT2 #(
		.INIT('h2)
	) name435 (
		\G2_pad ,
		_w71_,
		_w467_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		_w204_,
		_w467_,
		_w468_
	);
	LUT2 #(
		.INIT('h2)
	) name437 (
		\G10_pad ,
		_w34_,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name438 (
		_w245_,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h1)
	) name439 (
		\G10_pad ,
		_w98_,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name440 (
		\G6_pad ,
		\G9_pad ,
		_w472_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		_w228_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h1)
	) name442 (
		_w134_,
		_w154_,
		_w474_
	);
	LUT2 #(
		.INIT('h1)
	) name443 (
		\G12_pad ,
		_w474_,
		_w475_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w259_,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		_w55_,
		_w232_,
		_w477_
	);
	LUT2 #(
		.INIT('h2)
	) name446 (
		\G8_pad ,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h8)
	) name447 (
		_w47_,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h1)
	) name448 (
		\G3_pad ,
		\G44_reg/NET0131 ,
		_w480_
	);
	LUT2 #(
		.INIT('h1)
	) name449 (
		_w479_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h2)
	) name450 (
		_w225_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h8)
	) name451 (
		_w54_,
		_w147_,
		_w483_
	);
	LUT2 #(
		.INIT('h4)
	) name452 (
		_w157_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h8)
	) name453 (
		_w238_,
		_w478_,
		_w485_
	);
	LUT2 #(
		.INIT('h1)
	) name454 (
		_w484_,
		_w485_,
		_w486_
	);
	LUT2 #(
		.INIT('h4)
	) name455 (
		\G12_pad ,
		_w106_,
		_w487_
	);
	LUT2 #(
		.INIT('h4)
	) name456 (
		_w486_,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		\G37_reg/NET0131 ,
		\G38_reg/NET0131 ,
		_w489_
	);
	LUT2 #(
		.INIT('h8)
	) name458 (
		_w264_,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		_w259_,
		_w490_,
		_w491_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		_w488_,
		_w491_,
		_w492_
	);
	LUT2 #(
		.INIT('h2)
	) name461 (
		_w227_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name462 (
		_w482_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h2)
	) name463 (
		_w36_,
		_w228_,
		_w495_
	);
	LUT2 #(
		.INIT('h8)
	) name464 (
		_w197_,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('h8)
	) name465 (
		\G34_reg/NET0131 ,
		_w288_,
		_w497_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		_w496_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		_w283_,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h8)
	) name468 (
		_w324_,
		_w339_,
		_w500_
	);
	LUT2 #(
		.INIT('h8)
	) name469 (
		\G0_pad ,
		\G12_pad ,
		_w501_
	);
	LUT2 #(
		.INIT('h8)
	) name470 (
		_w90_,
		_w501_,
		_w502_
	);
	LUT2 #(
		.INIT('h8)
	) name471 (
		_w196_,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		_w500_,
		_w503_,
		_w504_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		\G6_pad ,
		_w54_,
		_w505_
	);
	LUT2 #(
		.INIT('h8)
	) name474 (
		_w114_,
		_w472_,
		_w506_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w505_,
		_w506_,
		_w507_
	);
	assign \G532_pad  = _w211_ ;
	assign \G537_pad  = _w269_ ;
	assign \G539_pad  = _w277_ ;
	assign \G542_pad  = _w294_ ;
	assign \G546_pad  = \G41_reg/NET0131 ;
	assign \G547_pad  = _w309_ ;
	assign \G548_pad  = _w317_ ;
	assign \G549_pad  = _w345_ ;
	assign \G550_pad  = _w359_ ;
	assign \G551_pad  = _w383_ ;
	assign \G552_pad  = _w403_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g1667/_3_  = _w414_ ;
	assign \g1737/_0_  = _w429_ ;
	assign \g1744/_0_  = _w430_ ;
	assign \g1787/_0_  = _w438_ ;
	assign \g1811/_0_  = _w446_ ;
	assign \g1830/_0_  = _w451_ ;
	assign \g1831/_0_  = _w457_ ;
	assign \g1846/_0_  = _w459_ ;
	assign \g1852/_0_  = _w462_ ;
	assign \g1866/_0_  = _w465_ ;
	assign \g19/_2_  = _w466_ ;
	assign \g1931/_0_  = _w468_ ;
	assign \g1945/_0_  = _w470_ ;
	assign \g2014/_0_  = _w471_ ;
	assign \g2015/_0_  = _w473_ ;
	assign \g2643/_0_  = _w476_ ;
	assign \g2859/_1_  = _w494_ ;
	assign \g3397/_2_  = _w499_ ;
	assign \g3546/_0_  = _w504_ ;
	assign \g3606/_3_  = _w507_ ;
endmodule;