module top (\1(0)_pad , \107(12)_pad , \116(13)_pad , \124(14)_pad , \125(15)_pad , \128(16)_pad , \13(1)_pad , \132(17)_pad , \137(18)_pad , \143(19)_pad , \150(20)_pad , \159(21)_pad , \169(22)_pad , \1698(48)_pad , \179(23)_pad , \190(24)_pad , \20(2)_pad , \200(25)_pad , \213(26)_pad , \222(27)_pad , \223(28)_pad , \226(29)_pad , \232(30)_pad , \238(31)_pad , \244(32)_pad , \250(33)_pad , \257(34)_pad , \264(35)_pad , \270(36)_pad , \274(37)_pad , \283(38)_pad , \2897(49)_pad , \294(39)_pad , \303(40)_pad , \311(41)_pad , \317(42)_pad , \322(43)_pad , \326(44)_pad , \329(45)_pad , \33(3)_pad , \330(46)_pad , \343(47)_pad , \41(4)_pad , \45(5)_pad , \50(6)_pad , \58(7)_pad , \68(8)_pad , \77(9)_pad , \87(10)_pad , \97(11)_pad , \2690(1611) , \2709(1587) , \353(405)_pad , \355(399)_pad , \358(1161)_pad , \361(940)_pad , \364(1484)_pad , \367(1585)_pad , \369(1321)_pad , \372(1243)_pad , \381(1626)_pad , \384(1553)_pad , \387(1616)_pad , \390(1603)_pad , \393(1605)_pad , \396(1504)_pad , \399(1428)_pad , \402(1718)_pad , \404(1714) , \407(1657)_pad , \409(1670)_pad , \605(1186) );
	input \1(0)_pad  ;
	input \107(12)_pad  ;
	input \116(13)_pad  ;
	input \124(14)_pad  ;
	input \125(15)_pad  ;
	input \128(16)_pad  ;
	input \13(1)_pad  ;
	input \132(17)_pad  ;
	input \137(18)_pad  ;
	input \143(19)_pad  ;
	input \150(20)_pad  ;
	input \159(21)_pad  ;
	input \169(22)_pad  ;
	input \1698(48)_pad  ;
	input \179(23)_pad  ;
	input \190(24)_pad  ;
	input \20(2)_pad  ;
	input \200(25)_pad  ;
	input \213(26)_pad  ;
	input \222(27)_pad  ;
	input \223(28)_pad  ;
	input \226(29)_pad  ;
	input \232(30)_pad  ;
	input \238(31)_pad  ;
	input \244(32)_pad  ;
	input \250(33)_pad  ;
	input \257(34)_pad  ;
	input \264(35)_pad  ;
	input \270(36)_pad  ;
	input \274(37)_pad  ;
	input \283(38)_pad  ;
	input \2897(49)_pad  ;
	input \294(39)_pad  ;
	input \303(40)_pad  ;
	input \311(41)_pad  ;
	input \317(42)_pad  ;
	input \322(43)_pad  ;
	input \326(44)_pad  ;
	input \329(45)_pad  ;
	input \33(3)_pad  ;
	input \330(46)_pad  ;
	input \343(47)_pad  ;
	input \41(4)_pad  ;
	input \45(5)_pad  ;
	input \50(6)_pad  ;
	input \58(7)_pad  ;
	input \68(8)_pad  ;
	input \77(9)_pad  ;
	input \87(10)_pad  ;
	input \97(11)_pad  ;
	output \2690(1611)  ;
	output \2709(1587)  ;
	output \353(405)_pad  ;
	output \355(399)_pad  ;
	output \358(1161)_pad  ;
	output \361(940)_pad  ;
	output \364(1484)_pad  ;
	output \367(1585)_pad  ;
	output \369(1321)_pad  ;
	output \372(1243)_pad  ;
	output \381(1626)_pad  ;
	output \384(1553)_pad  ;
	output \387(1616)_pad  ;
	output \390(1603)_pad  ;
	output \393(1605)_pad  ;
	output \396(1504)_pad  ;
	output \399(1428)_pad  ;
	output \402(1718)_pad  ;
	output \404(1714)  ;
	output \407(1657)_pad  ;
	output \409(1670)_pad  ;
	output \605(1186)  ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\13(1)_pad ,
		\20(2)_pad ,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\1(0)_pad ,
		\213(26)_pad ,
		_w52_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		_w51_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\1(0)_pad ,
		\13(1)_pad ,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\1(0)_pad ,
		\20(2)_pad ,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\33(3)_pad ,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		_w54_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		\20(2)_pad ,
		\33(3)_pad ,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\68(8)_pad ,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		\58(7)_pad ,
		\68(8)_pad ,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\58(7)_pad ,
		\68(8)_pad ,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		_w60_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		\20(2)_pad ,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\20(2)_pad ,
		\33(3)_pad ,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\159(21)_pad ,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		_w59_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		_w63_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w57_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		\13(1)_pad ,
		\20(2)_pad ,
		_w69_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		\1(0)_pad ,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		\58(7)_pad ,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		\1(0)_pad ,
		\20(2)_pad ,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		_w57_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\58(7)_pad ,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w68_,
		_w71_,
		_w75_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		_w74_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		\33(3)_pad ,
		\41(4)_pad ,
		_w77_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		_w54_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\41(4)_pad ,
		\45(5)_pad ,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		\1(0)_pad ,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w78_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		\232(30)_pad ,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		\274(37)_pad ,
		_w78_,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w80_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		\1698(48)_pad ,
		\33(3)_pad ,
		_w85_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\223(28)_pad ,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h2)
	) name36 (
		\1698(48)_pad ,
		\33(3)_pad ,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\226(29)_pad ,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\33(3)_pad ,
		\87(10)_pad ,
		_w89_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w86_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		_w88_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h2)
	) name41 (
		_w78_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w82_,
		_w84_,
		_w93_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		_w92_,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\169(22)_pad ,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		\179(23)_pad ,
		_w94_,
		_w96_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w76_,
		_w95_,
		_w97_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		_w96_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w53_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		\343(47)_pad ,
		_w53_,
		_w100_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\13(1)_pad ,
		\33(3)_pad ,
		_w101_
	);
	LUT2 #(
		.INIT('h2)
	) name51 (
		_w55_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w70_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		\68(8)_pad ,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		\68(8)_pad ,
		_w73_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		\33(3)_pad ,
		\77(9)_pad ,
		_w106_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		\33(3)_pad ,
		\50(6)_pad ,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		_w106_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		\20(2)_pad ,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		_w57_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		_w104_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		_w105_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		\238(31)_pad ,
		_w81_,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		\226(29)_pad ,
		_w85_,
		_w114_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		\33(3)_pad ,
		\97(11)_pad ,
		_w115_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		\232(30)_pad ,
		_w87_,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w114_,
		_w115_,
		_w117_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		_w116_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		_w78_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		_w84_,
		_w113_,
		_w120_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		_w119_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		\169(22)_pad ,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		\179(23)_pad ,
		_w121_,
		_w123_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w112_,
		_w122_,
		_w124_
	);
	LUT2 #(
		.INIT('h4)
	) name74 (
		_w123_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		\190(24)_pad ,
		_w121_,
		_w126_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		\200(25)_pad ,
		_w121_,
		_w127_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		_w112_,
		_w126_,
		_w128_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		_w127_,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		_w125_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		_w100_,
		_w112_,
		_w131_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		_w130_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		\77(9)_pad ,
		_w70_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\77(9)_pad ,
		_w73_,
		_w134_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		\20(2)_pad ,
		\77(9)_pad ,
		_w135_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\33(3)_pad ,
		\58(7)_pad ,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\20(2)_pad ,
		_w89_,
		_w137_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		_w136_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		_w57_,
		_w135_,
		_w139_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		_w138_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		_w133_,
		_w134_,
		_w141_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		_w140_,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		\244(32)_pad ,
		_w81_,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		\232(30)_pad ,
		_w85_,
		_w144_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		\107(12)_pad ,
		\33(3)_pad ,
		_w145_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		\238(31)_pad ,
		_w87_,
		_w146_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w144_,
		_w145_,
		_w147_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		_w146_,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		_w78_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		_w84_,
		_w143_,
		_w150_
	);
	LUT2 #(
		.INIT('h4)
	) name100 (
		_w149_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		\169(22)_pad ,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		\179(23)_pad ,
		_w151_,
		_w153_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		_w142_,
		_w152_,
		_w154_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		_w153_,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		\238(31)_pad ,
		_w85_,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		\244(32)_pad ,
		_w87_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		\116(13)_pad ,
		\33(3)_pad ,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		_w156_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h4)
	) name109 (
		_w157_,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h2)
	) name110 (
		_w78_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		\1(0)_pad ,
		\45(5)_pad ,
		_w162_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		\250(33)_pad ,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h4)
	) name113 (
		\274(37)_pad ,
		_w162_,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		_w78_,
		_w163_,
		_w165_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		_w164_,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w161_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\179(23)_pad ,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h2)
	) name118 (
		\169(22)_pad ,
		_w167_,
		_w169_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w168_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		\87(10)_pad ,
		_w70_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		\33(3)_pad ,
		_w69_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		\1(0)_pad ,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h2)
	) name123 (
		_w57_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		\87(10)_pad ,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		\107(12)_pad ,
		\87(10)_pad ,
		_w176_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		\97(11)_pad ,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		\20(2)_pad ,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		\68(8)_pad ,
		_w64_,
		_w179_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w115_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		_w178_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w57_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		_w171_,
		_w175_,
		_w183_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		_w182_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		_w170_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		\116(13)_pad ,
		_w70_,
		_w186_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		\116(13)_pad ,
		_w174_,
		_w187_
	);
	LUT2 #(
		.INIT('h4)
	) name137 (
		\116(13)_pad ,
		\20(2)_pad ,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		\283(38)_pad ,
		\33(3)_pad ,
		_w189_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		\33(3)_pad ,
		\97(11)_pad ,
		_w190_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		\20(2)_pad ,
		_w189_,
		_w191_
	);
	LUT2 #(
		.INIT('h4)
	) name141 (
		_w190_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		_w57_,
		_w188_,
		_w193_
	);
	LUT2 #(
		.INIT('h4)
	) name143 (
		_w192_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w186_,
		_w187_,
		_w195_
	);
	LUT2 #(
		.INIT('h4)
	) name145 (
		_w194_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h4)
	) name146 (
		\41(4)_pad ,
		_w162_,
		_w197_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w83_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\264(35)_pad ,
		_w87_,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		\257(34)_pad ,
		_w85_,
		_w200_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		\303(40)_pad ,
		\33(3)_pad ,
		_w201_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w199_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h4)
	) name152 (
		_w200_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h2)
	) name153 (
		_w78_,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		_w78_,
		_w197_,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		\270(36)_pad ,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		_w204_,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h4)
	) name157 (
		_w198_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		\169(22)_pad ,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		\179(23)_pad ,
		_w208_,
		_w210_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		_w209_,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		_w196_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		\107(12)_pad ,
		_w103_,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		\107(12)_pad ,
		_w174_,
		_w214_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		\33(3)_pad ,
		\87(10)_pad ,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w158_,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		\20(2)_pad ,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h4)
	) name167 (
		_w57_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		_w213_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		_w214_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		\264(35)_pad ,
		_w205_,
		_w221_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		\257(34)_pad ,
		_w87_,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		\250(33)_pad ,
		_w85_,
		_w223_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		\294(39)_pad ,
		\33(3)_pad ,
		_w224_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		_w222_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		_w223_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		_w78_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		_w198_,
		_w221_,
		_w228_
	);
	LUT2 #(
		.INIT('h4)
	) name178 (
		_w227_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		\169(22)_pad ,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h4)
	) name180 (
		\179(23)_pad ,
		_w229_,
		_w231_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		_w220_,
		_w230_,
		_w232_
	);
	LUT2 #(
		.INIT('h4)
	) name182 (
		_w231_,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		_w212_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		\190(24)_pad ,
		_w229_,
		_w235_
	);
	LUT2 #(
		.INIT('h2)
	) name185 (
		\200(25)_pad ,
		_w229_,
		_w236_
	);
	LUT2 #(
		.INIT('h2)
	) name186 (
		_w220_,
		_w235_,
		_w237_
	);
	LUT2 #(
		.INIT('h4)
	) name187 (
		_w236_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h8)
	) name188 (
		\257(34)_pad ,
		_w205_,
		_w239_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		\244(32)_pad ,
		_w85_,
		_w240_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		\250(33)_pad ,
		_w87_,
		_w241_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		_w189_,
		_w240_,
		_w242_
	);
	LUT2 #(
		.INIT('h4)
	) name192 (
		_w241_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h2)
	) name193 (
		_w78_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		_w198_,
		_w239_,
		_w245_
	);
	LUT2 #(
		.INIT('h4)
	) name195 (
		_w244_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\190(24)_pad ,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h4)
	) name197 (
		\97(11)_pad ,
		_w70_,
		_w248_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		\97(11)_pad ,
		_w174_,
		_w249_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		\33(3)_pad ,
		\77(9)_pad ,
		_w250_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		\20(2)_pad ,
		_w145_,
		_w251_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		_w250_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		\107(12)_pad ,
		\97(11)_pad ,
		_w253_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		\107(12)_pad ,
		\97(11)_pad ,
		_w254_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		_w253_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\20(2)_pad ,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		_w57_,
		_w252_,
		_w257_
	);
	LUT2 #(
		.INIT('h4)
	) name207 (
		_w256_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		_w248_,
		_w249_,
		_w259_
	);
	LUT2 #(
		.INIT('h4)
	) name209 (
		_w258_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h2)
	) name210 (
		\200(25)_pad ,
		_w246_,
		_w261_
	);
	LUT2 #(
		.INIT('h4)
	) name211 (
		_w247_,
		_w260_,
		_w262_
	);
	LUT2 #(
		.INIT('h4)
	) name212 (
		_w261_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w238_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h4)
	) name214 (
		_w234_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		\169(22)_pad ,
		_w246_,
		_w266_
	);
	LUT2 #(
		.INIT('h4)
	) name216 (
		\179(23)_pad ,
		_w246_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		_w260_,
		_w266_,
		_w268_
	);
	LUT2 #(
		.INIT('h4)
	) name218 (
		_w267_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name219 (
		_w265_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		\190(24)_pad ,
		_w167_,
		_w271_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		\200(25)_pad ,
		_w167_,
		_w272_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		_w184_,
		_w271_,
		_w273_
	);
	LUT2 #(
		.INIT('h4)
	) name223 (
		_w272_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w270_,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w185_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h2)
	) name226 (
		_w100_,
		_w142_,
		_w277_
	);
	LUT2 #(
		.INIT('h2)
	) name227 (
		\200(25)_pad ,
		_w151_,
		_w278_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		\190(24)_pad ,
		_w151_,
		_w279_
	);
	LUT2 #(
		.INIT('h2)
	) name229 (
		_w142_,
		_w278_,
		_w280_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		_w279_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w155_,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h4)
	) name232 (
		_w277_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		_w276_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h1)
	) name234 (
		_w155_,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h2)
	) name235 (
		_w132_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		_w125_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w100_,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h2)
	) name238 (
		_w53_,
		_w76_,
		_w289_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		\190(24)_pad ,
		_w94_,
		_w290_
	);
	LUT2 #(
		.INIT('h2)
	) name240 (
		\200(25)_pad ,
		_w94_,
		_w291_
	);
	LUT2 #(
		.INIT('h2)
	) name241 (
		_w76_,
		_w290_,
		_w292_
	);
	LUT2 #(
		.INIT('h4)
	) name242 (
		_w291_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		_w289_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w98_,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		_w288_,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		_w99_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		\58(7)_pad ,
		_w58_,
		_w298_
	);
	LUT2 #(
		.INIT('h4)
	) name248 (
		\50(6)_pad ,
		_w60_,
		_w299_
	);
	LUT2 #(
		.INIT('h2)
	) name249 (
		\20(2)_pad ,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		\150(20)_pad ,
		_w64_,
		_w301_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		_w298_,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		_w300_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w57_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h4)
	) name254 (
		\50(6)_pad ,
		_w70_,
		_w305_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		\50(6)_pad ,
		_w73_,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		_w304_,
		_w305_,
		_w307_
	);
	LUT2 #(
		.INIT('h4)
	) name257 (
		_w306_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		\226(29)_pad ,
		_w81_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		\222(27)_pad ,
		_w85_,
		_w310_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		\223(28)_pad ,
		_w87_,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w106_,
		_w310_,
		_w312_
	);
	LUT2 #(
		.INIT('h4)
	) name262 (
		_w311_,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		_w78_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		_w84_,
		_w309_,
		_w315_
	);
	LUT2 #(
		.INIT('h4)
	) name265 (
		_w314_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name266 (
		\169(22)_pad ,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		\179(23)_pad ,
		_w316_,
		_w318_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w308_,
		_w317_,
		_w319_
	);
	LUT2 #(
		.INIT('h4)
	) name269 (
		_w318_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		\190(24)_pad ,
		_w316_,
		_w321_
	);
	LUT2 #(
		.INIT('h2)
	) name271 (
		\200(25)_pad ,
		_w316_,
		_w322_
	);
	LUT2 #(
		.INIT('h2)
	) name272 (
		_w308_,
		_w321_,
		_w323_
	);
	LUT2 #(
		.INIT('h4)
	) name273 (
		_w322_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		_w320_,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		_w53_,
		_w308_,
		_w326_
	);
	LUT2 #(
		.INIT('h2)
	) name276 (
		_w325_,
		_w326_,
		_w327_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		_w53_,
		_w320_,
		_w328_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		_w327_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h2)
	) name279 (
		\200(25)_pad ,
		_w208_,
		_w330_
	);
	LUT2 #(
		.INIT('h8)
	) name280 (
		\190(24)_pad ,
		_w208_,
		_w331_
	);
	LUT2 #(
		.INIT('h2)
	) name281 (
		_w196_,
		_w330_,
		_w332_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		_w331_,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		_w212_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		_w185_,
		_w274_,
		_w335_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		_w233_,
		_w269_,
		_w336_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		_w264_,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		_w335_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		_w334_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w100_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		_w207_,
		_w229_,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		_w246_,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		_w168_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		\179(23)_pad ,
		_w167_,
		_w344_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		_w229_,
		_w246_,
		_w345_
	);
	LUT2 #(
		.INIT('h8)
	) name295 (
		_w344_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h4)
	) name296 (
		_w208_,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h2)
	) name297 (
		_w100_,
		_w343_,
		_w348_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		_w347_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h2)
	) name299 (
		\330(46)_pad ,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h4)
	) name300 (
		_w340_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		_w99_,
		_w295_,
		_w352_
	);
	LUT2 #(
		.INIT('h8)
	) name302 (
		_w100_,
		_w155_,
		_w353_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		_w283_,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h8)
	) name304 (
		_w100_,
		_w125_,
		_w355_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		_w132_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		_w354_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name307 (
		_w352_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h8)
	) name308 (
		_w351_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h4)
	) name309 (
		_w329_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h2)
	) name310 (
		_w329_,
		_w359_,
		_w361_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		_w360_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h8)
	) name312 (
		_w297_,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		_w297_,
		_w362_,
		_w364_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		_w363_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h8)
	) name315 (
		\45(5)_pad ,
		_w51_,
		_w366_
	);
	LUT2 #(
		.INIT('h2)
	) name316 (
		\1(0)_pad ,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w365_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h4)
	) name318 (
		\13(1)_pad ,
		_w55_,
		_w369_
	);
	LUT2 #(
		.INIT('h4)
	) name319 (
		\41(4)_pad ,
		_w369_,
		_w370_
	);
	LUT2 #(
		.INIT('h2)
	) name320 (
		_w367_,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h4)
	) name321 (
		\169(22)_pad ,
		\20(2)_pad ,
		_w372_
	);
	LUT2 #(
		.INIT('h2)
	) name322 (
		_w54_,
		_w372_,
		_w373_
	);
	LUT2 #(
		.INIT('h2)
	) name323 (
		\41(4)_pad ,
		\50(6)_pad ,
		_w374_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		\179(23)_pad ,
		\20(2)_pad ,
		_w375_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		\200(25)_pad ,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h8)
	) name326 (
		\190(24)_pad ,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		\125(15)_pad ,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h8)
	) name328 (
		\20(2)_pad ,
		\200(25)_pad ,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name329 (
		_w375_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h4)
	) name330 (
		\190(24)_pad ,
		\20(2)_pad ,
		_w381_
	);
	LUT2 #(
		.INIT('h2)
	) name331 (
		_w380_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		\150(20)_pad ,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		\200(25)_pad ,
		_w375_,
		_w384_
	);
	LUT2 #(
		.INIT('h8)
	) name334 (
		\190(24)_pad ,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h8)
	) name335 (
		\128(16)_pad ,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h8)
	) name336 (
		_w380_,
		_w381_,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		\124(14)_pad ,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h4)
	) name338 (
		\190(24)_pad ,
		_w384_,
		_w389_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		\137(18)_pad ,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h4)
	) name340 (
		\190(24)_pad ,
		_w376_,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		\132(17)_pad ,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		_w375_,
		_w379_,
		_w393_
	);
	LUT2 #(
		.INIT('h8)
	) name343 (
		\190(24)_pad ,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h8)
	) name344 (
		\143(19)_pad ,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h4)
	) name345 (
		\190(24)_pad ,
		_w393_,
		_w396_
	);
	LUT2 #(
		.INIT('h8)
	) name346 (
		\159(21)_pad ,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		\33(3)_pad ,
		\41(4)_pad ,
		_w398_
	);
	LUT2 #(
		.INIT('h4)
	) name348 (
		_w378_,
		_w398_,
		_w399_
	);
	LUT2 #(
		.INIT('h1)
	) name349 (
		_w383_,
		_w386_,
		_w400_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		_w388_,
		_w390_,
		_w401_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		_w392_,
		_w395_,
		_w402_
	);
	LUT2 #(
		.INIT('h4)
	) name352 (
		_w397_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h8)
	) name353 (
		_w400_,
		_w401_,
		_w404_
	);
	LUT2 #(
		.INIT('h8)
	) name354 (
		_w399_,
		_w404_,
		_w405_
	);
	LUT2 #(
		.INIT('h8)
	) name355 (
		_w403_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		\58(7)_pad ,
		_w396_,
		_w407_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		\283(38)_pad ,
		_w387_,
		_w408_
	);
	LUT2 #(
		.INIT('h8)
	) name358 (
		\77(9)_pad ,
		_w394_,
		_w409_
	);
	LUT2 #(
		.INIT('h8)
	) name359 (
		\97(11)_pad ,
		_w391_,
		_w410_
	);
	LUT2 #(
		.INIT('h8)
	) name360 (
		\107(12)_pad ,
		_w385_,
		_w411_
	);
	LUT2 #(
		.INIT('h8)
	) name361 (
		\116(13)_pad ,
		_w377_,
		_w412_
	);
	LUT2 #(
		.INIT('h8)
	) name362 (
		\68(8)_pad ,
		_w382_,
		_w413_
	);
	LUT2 #(
		.INIT('h8)
	) name363 (
		\87(10)_pad ,
		_w389_,
		_w414_
	);
	LUT2 #(
		.INIT('h2)
	) name364 (
		\33(3)_pad ,
		\41(4)_pad ,
		_w415_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w407_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h1)
	) name366 (
		_w408_,
		_w409_,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w410_,
		_w411_,
		_w418_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		_w412_,
		_w413_,
		_w419_
	);
	LUT2 #(
		.INIT('h4)
	) name369 (
		_w414_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h8)
	) name370 (
		_w417_,
		_w418_,
		_w421_
	);
	LUT2 #(
		.INIT('h8)
	) name371 (
		_w416_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h8)
	) name372 (
		_w420_,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h1)
	) name373 (
		_w374_,
		_w406_,
		_w424_
	);
	LUT2 #(
		.INIT('h4)
	) name374 (
		_w423_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		_w373_,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h8)
	) name376 (
		_w101_,
		_w329_,
		_w427_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		_w101_,
		_w373_,
		_w428_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		\50(6)_pad ,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h2)
	) name379 (
		_w371_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h4)
	) name380 (
		_w426_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h4)
	) name381 (
		_w427_,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		_w100_,
		_w276_,
		_w433_
	);
	LUT2 #(
		.INIT('h1)
	) name383 (
		_w351_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		_w98_,
		_w293_,
		_w435_
	);
	LUT2 #(
		.INIT('h8)
	) name385 (
		_w130_,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		_w282_,
		_w325_,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name387 (
		_w436_,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('h4)
	) name388 (
		_w434_,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h4)
	) name389 (
		_w129_,
		_w155_,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name390 (
		_w125_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h1)
	) name391 (
		_w293_,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h1)
	) name392 (
		_w98_,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		_w324_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		_w320_,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h4)
	) name395 (
		_w439_,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h2)
	) name396 (
		_w351_,
		_w354_,
		_w447_
	);
	LUT2 #(
		.INIT('h2)
	) name397 (
		_w356_,
		_w447_,
		_w448_
	);
	LUT2 #(
		.INIT('h8)
	) name398 (
		_w351_,
		_w357_,
		_w449_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		_w448_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		_w100_,
		_w285_,
		_w451_
	);
	LUT2 #(
		.INIT('h4)
	) name401 (
		_w450_,
		_w451_,
		_w452_
	);
	LUT2 #(
		.INIT('h2)
	) name402 (
		_w450_,
		_w451_,
		_w453_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		_w452_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h2)
	) name404 (
		_w446_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w352_,
		_w449_,
		_w456_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		_w359_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h4)
	) name407 (
		_w288_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h2)
	) name408 (
		_w288_,
		_w457_,
		_w459_
	);
	LUT2 #(
		.INIT('h1)
	) name409 (
		_w458_,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('h2)
	) name410 (
		_w455_,
		_w460_,
		_w461_
	);
	LUT2 #(
		.INIT('h2)
	) name411 (
		_w446_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h4)
	) name412 (
		_w365_,
		_w370_,
		_w463_
	);
	LUT2 #(
		.INIT('h4)
	) name413 (
		_w462_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		_w368_,
		_w432_,
		_w465_
	);
	LUT2 #(
		.INIT('h4)
	) name415 (
		_w464_,
		_w465_,
		_w466_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		_w367_,
		_w460_,
		_w467_
	);
	LUT2 #(
		.INIT('h8)
	) name417 (
		\137(18)_pad ,
		_w391_,
		_w468_
	);
	LUT2 #(
		.INIT('h8)
	) name418 (
		\50(6)_pad ,
		_w396_,
		_w469_
	);
	LUT2 #(
		.INIT('h8)
	) name419 (
		\132(17)_pad ,
		_w385_,
		_w470_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		\143(19)_pad ,
		_w389_,
		_w471_
	);
	LUT2 #(
		.INIT('h8)
	) name421 (
		\125(15)_pad ,
		_w387_,
		_w472_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		\150(20)_pad ,
		_w394_,
		_w473_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		\128(16)_pad ,
		_w377_,
		_w474_
	);
	LUT2 #(
		.INIT('h8)
	) name424 (
		\159(21)_pad ,
		_w382_,
		_w475_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		\33(3)_pad ,
		_w468_,
		_w476_
	);
	LUT2 #(
		.INIT('h1)
	) name426 (
		_w469_,
		_w470_,
		_w477_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		_w471_,
		_w472_,
		_w478_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		_w473_,
		_w474_,
		_w479_
	);
	LUT2 #(
		.INIT('h4)
	) name429 (
		_w475_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h8)
	) name430 (
		_w477_,
		_w478_,
		_w481_
	);
	LUT2 #(
		.INIT('h8)
	) name431 (
		_w476_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		_w480_,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h8)
	) name433 (
		\68(8)_pad ,
		_w396_,
		_w484_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		\87(10)_pad ,
		_w394_,
		_w485_
	);
	LUT2 #(
		.INIT('h8)
	) name435 (
		\294(39)_pad ,
		_w387_,
		_w486_
	);
	LUT2 #(
		.INIT('h8)
	) name436 (
		\97(11)_pad ,
		_w389_,
		_w487_
	);
	LUT2 #(
		.INIT('h8)
	) name437 (
		\116(13)_pad ,
		_w385_,
		_w488_
	);
	LUT2 #(
		.INIT('h8)
	) name438 (
		\77(9)_pad ,
		_w382_,
		_w489_
	);
	LUT2 #(
		.INIT('h8)
	) name439 (
		\107(12)_pad ,
		_w391_,
		_w490_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		\283(38)_pad ,
		_w377_,
		_w491_
	);
	LUT2 #(
		.INIT('h2)
	) name441 (
		\33(3)_pad ,
		_w484_,
		_w492_
	);
	LUT2 #(
		.INIT('h1)
	) name442 (
		_w485_,
		_w486_,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name443 (
		_w487_,
		_w488_,
		_w494_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w489_,
		_w490_,
		_w495_
	);
	LUT2 #(
		.INIT('h4)
	) name445 (
		_w491_,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('h8)
	) name446 (
		_w493_,
		_w494_,
		_w497_
	);
	LUT2 #(
		.INIT('h8)
	) name447 (
		_w492_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		_w496_,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h1)
	) name449 (
		_w483_,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h2)
	) name450 (
		_w373_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h2)
	) name451 (
		_w101_,
		_w352_,
		_w502_
	);
	LUT2 #(
		.INIT('h4)
	) name452 (
		\58(7)_pad ,
		_w428_,
		_w503_
	);
	LUT2 #(
		.INIT('h2)
	) name453 (
		_w371_,
		_w503_,
		_w504_
	);
	LUT2 #(
		.INIT('h4)
	) name454 (
		_w501_,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h4)
	) name455 (
		_w502_,
		_w505_,
		_w506_
	);
	LUT2 #(
		.INIT('h4)
	) name456 (
		_w455_,
		_w460_,
		_w507_
	);
	LUT2 #(
		.INIT('h2)
	) name457 (
		_w370_,
		_w461_,
		_w508_
	);
	LUT2 #(
		.INIT('h4)
	) name458 (
		_w507_,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		_w467_,
		_w506_,
		_w510_
	);
	LUT2 #(
		.INIT('h4)
	) name460 (
		_w509_,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		\50(6)_pad ,
		\77(9)_pad ,
		_w512_
	);
	LUT2 #(
		.INIT('h8)
	) name462 (
		_w60_,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h2)
	) name463 (
		\87(10)_pad ,
		_w253_,
		_w514_
	);
	LUT2 #(
		.INIT('h1)
	) name464 (
		\257(34)_pad ,
		\264(35)_pad ,
		_w515_
	);
	LUT2 #(
		.INIT('h8)
	) name465 (
		\257(34)_pad ,
		\264(35)_pad ,
		_w516_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		_w515_,
		_w516_,
		_w517_
	);
	LUT2 #(
		.INIT('h2)
	) name467 (
		\250(33)_pad ,
		\270(36)_pad ,
		_w518_
	);
	LUT2 #(
		.INIT('h4)
	) name468 (
		\250(33)_pad ,
		\270(36)_pad ,
		_w519_
	);
	LUT2 #(
		.INIT('h1)
	) name469 (
		_w518_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h8)
	) name470 (
		_w517_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h1)
	) name471 (
		_w517_,
		_w520_,
		_w522_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		_w521_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h2)
	) name473 (
		\226(29)_pad ,
		\232(30)_pad ,
		_w524_
	);
	LUT2 #(
		.INIT('h4)
	) name474 (
		\226(29)_pad ,
		\232(30)_pad ,
		_w525_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w524_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h2)
	) name476 (
		\238(31)_pad ,
		\244(32)_pad ,
		_w527_
	);
	LUT2 #(
		.INIT('h4)
	) name477 (
		\238(31)_pad ,
		\244(32)_pad ,
		_w528_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		_w527_,
		_w528_,
		_w529_
	);
	LUT2 #(
		.INIT('h8)
	) name479 (
		_w526_,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h1)
	) name480 (
		_w526_,
		_w529_,
		_w531_
	);
	LUT2 #(
		.INIT('h1)
	) name481 (
		_w530_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h8)
	) name482 (
		_w523_,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		_w523_,
		_w532_,
		_w534_
	);
	LUT2 #(
		.INIT('h1)
	) name484 (
		_w533_,
		_w534_,
		_w535_
	);
	LUT2 #(
		.INIT('h8)
	) name485 (
		\232(30)_pad ,
		\58(7)_pad ,
		_w536_
	);
	LUT2 #(
		.INIT('h8)
	) name486 (
		\226(29)_pad ,
		\50(6)_pad ,
		_w537_
	);
	LUT2 #(
		.INIT('h8)
	) name487 (
		\250(33)_pad ,
		\87(10)_pad ,
		_w538_
	);
	LUT2 #(
		.INIT('h8)
	) name488 (
		\244(32)_pad ,
		\77(9)_pad ,
		_w539_
	);
	LUT2 #(
		.INIT('h8)
	) name489 (
		\116(13)_pad ,
		\270(36)_pad ,
		_w540_
	);
	LUT2 #(
		.INIT('h8)
	) name490 (
		\107(12)_pad ,
		\264(35)_pad ,
		_w541_
	);
	LUT2 #(
		.INIT('h8)
	) name491 (
		\238(31)_pad ,
		\68(8)_pad ,
		_w542_
	);
	LUT2 #(
		.INIT('h8)
	) name492 (
		\257(34)_pad ,
		\97(11)_pad ,
		_w543_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		_w536_,
		_w537_,
		_w544_
	);
	LUT2 #(
		.INIT('h1)
	) name494 (
		_w538_,
		_w539_,
		_w545_
	);
	LUT2 #(
		.INIT('h1)
	) name495 (
		_w540_,
		_w541_,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w542_,
		_w543_,
		_w547_
	);
	LUT2 #(
		.INIT('h8)
	) name497 (
		_w546_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		_w544_,
		_w545_,
		_w549_
	);
	LUT2 #(
		.INIT('h8)
	) name499 (
		_w548_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		_w55_,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h2)
	) name501 (
		\50(6)_pad ,
		_w60_,
		_w552_
	);
	LUT2 #(
		.INIT('h8)
	) name502 (
		\1(0)_pad ,
		_w69_,
		_w553_
	);
	LUT2 #(
		.INIT('h8)
	) name503 (
		_w552_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h2)
	) name504 (
		\250(33)_pad ,
		_w515_,
		_w555_
	);
	LUT2 #(
		.INIT('h8)
	) name505 (
		_w369_,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w554_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h4)
	) name507 (
		_w551_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		_w370_,
		_w552_,
		_w559_
	);
	LUT2 #(
		.INIT('h1)
	) name509 (
		\1(0)_pad ,
		_w434_,
		_w560_
	);
	LUT2 #(
		.INIT('h4)
	) name510 (
		\116(13)_pad ,
		_w177_,
		_w561_
	);
	LUT2 #(
		.INIT('h2)
	) name511 (
		\1(0)_pad ,
		_w370_,
		_w562_
	);
	LUT2 #(
		.INIT('h8)
	) name512 (
		_w561_,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h1)
	) name513 (
		_w559_,
		_w563_,
		_w564_
	);
	LUT2 #(
		.INIT('h4)
	) name514 (
		_w560_,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h4)
	) name515 (
		\50(6)_pad ,
		\68(8)_pad ,
		_w566_
	);
	LUT2 #(
		.INIT('h8)
	) name516 (
		\50(6)_pad ,
		\77(9)_pad ,
		_w567_
	);
	LUT2 #(
		.INIT('h8)
	) name517 (
		_w62_,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h1)
	) name518 (
		_w566_,
		_w568_,
		_w569_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		\13(1)_pad ,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h8)
	) name520 (
		\116(13)_pad ,
		_w255_,
		_w571_
	);
	LUT2 #(
		.INIT('h8)
	) name521 (
		_w69_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h1)
	) name522 (
		_w570_,
		_w572_,
		_w573_
	);
	LUT2 #(
		.INIT('h2)
	) name523 (
		\1(0)_pad ,
		_w573_,
		_w574_
	);
	LUT2 #(
		.INIT('h2)
	) name524 (
		\1(0)_pad ,
		_w51_,
		_w575_
	);
	LUT2 #(
		.INIT('h1)
	) name525 (
		_w358_,
		_w438_,
		_w576_
	);
	LUT2 #(
		.INIT('h8)
	) name526 (
		_w358_,
		_w438_,
		_w577_
	);
	LUT2 #(
		.INIT('h2)
	) name527 (
		_w351_,
		_w576_,
		_w578_
	);
	LUT2 #(
		.INIT('h4)
	) name528 (
		_w577_,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h4)
	) name529 (
		_w297_,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h2)
	) name530 (
		_w297_,
		_w579_,
		_w581_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w580_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h8)
	) name532 (
		_w433_,
		_w438_,
		_w583_
	);
	LUT2 #(
		.INIT('h2)
	) name533 (
		_w445_,
		_w583_,
		_w584_
	);
	LUT2 #(
		.INIT('h2)
	) name534 (
		_w582_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h4)
	) name535 (
		_w582_,
		_w584_,
		_w586_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w575_,
		_w585_,
		_w587_
	);
	LUT2 #(
		.INIT('h4)
	) name537 (
		_w586_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		_w574_,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h4)
	) name539 (
		_w276_,
		_w438_,
		_w590_
	);
	LUT2 #(
		.INIT('h2)
	) name540 (
		_w445_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h8)
	) name541 (
		_w339_,
		_w438_,
		_w592_
	);
	LUT2 #(
		.INIT('h1)
	) name542 (
		_w367_,
		_w454_,
		_w593_
	);
	LUT2 #(
		.INIT('h8)
	) name543 (
		\87(10)_pad ,
		_w382_,
		_w594_
	);
	LUT2 #(
		.INIT('h8)
	) name544 (
		\97(11)_pad ,
		_w394_,
		_w595_
	);
	LUT2 #(
		.INIT('h8)
	) name545 (
		\77(9)_pad ,
		_w396_,
		_w596_
	);
	LUT2 #(
		.INIT('h8)
	) name546 (
		\294(39)_pad ,
		_w377_,
		_w597_
	);
	LUT2 #(
		.INIT('h8)
	) name547 (
		\107(12)_pad ,
		_w389_,
		_w598_
	);
	LUT2 #(
		.INIT('h8)
	) name548 (
		\116(13)_pad ,
		_w391_,
		_w599_
	);
	LUT2 #(
		.INIT('h8)
	) name549 (
		\283(38)_pad ,
		_w385_,
		_w600_
	);
	LUT2 #(
		.INIT('h8)
	) name550 (
		\303(40)_pad ,
		_w387_,
		_w601_
	);
	LUT2 #(
		.INIT('h2)
	) name551 (
		\33(3)_pad ,
		_w594_,
		_w602_
	);
	LUT2 #(
		.INIT('h1)
	) name552 (
		_w595_,
		_w596_,
		_w603_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		_w597_,
		_w598_,
		_w604_
	);
	LUT2 #(
		.INIT('h1)
	) name554 (
		_w599_,
		_w600_,
		_w605_
	);
	LUT2 #(
		.INIT('h4)
	) name555 (
		_w601_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h8)
	) name556 (
		_w603_,
		_w604_,
		_w607_
	);
	LUT2 #(
		.INIT('h8)
	) name557 (
		_w602_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h8)
	) name558 (
		_w606_,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('h8)
	) name559 (
		\132(17)_pad ,
		_w377_,
		_w610_
	);
	LUT2 #(
		.INIT('h8)
	) name560 (
		\159(21)_pad ,
		_w394_,
		_w611_
	);
	LUT2 #(
		.INIT('h8)
	) name561 (
		\137(18)_pad ,
		_w385_,
		_w612_
	);
	LUT2 #(
		.INIT('h8)
	) name562 (
		\128(16)_pad ,
		_w387_,
		_w613_
	);
	LUT2 #(
		.INIT('h8)
	) name563 (
		\50(6)_pad ,
		_w382_,
		_w614_
	);
	LUT2 #(
		.INIT('h8)
	) name564 (
		\143(19)_pad ,
		_w391_,
		_w615_
	);
	LUT2 #(
		.INIT('h8)
	) name565 (
		\150(20)_pad ,
		_w389_,
		_w616_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		\33(3)_pad ,
		_w407_,
		_w617_
	);
	LUT2 #(
		.INIT('h1)
	) name567 (
		_w610_,
		_w611_,
		_w618_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		_w612_,
		_w613_,
		_w619_
	);
	LUT2 #(
		.INIT('h1)
	) name569 (
		_w614_,
		_w615_,
		_w620_
	);
	LUT2 #(
		.INIT('h4)
	) name570 (
		_w616_,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h8)
	) name571 (
		_w618_,
		_w619_,
		_w622_
	);
	LUT2 #(
		.INIT('h8)
	) name572 (
		_w617_,
		_w622_,
		_w623_
	);
	LUT2 #(
		.INIT('h8)
	) name573 (
		_w621_,
		_w623_,
		_w624_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		_w609_,
		_w624_,
		_w625_
	);
	LUT2 #(
		.INIT('h2)
	) name575 (
		_w373_,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h8)
	) name576 (
		_w101_,
		_w356_,
		_w627_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		\68(8)_pad ,
		_w428_,
		_w628_
	);
	LUT2 #(
		.INIT('h2)
	) name578 (
		_w371_,
		_w628_,
		_w629_
	);
	LUT2 #(
		.INIT('h4)
	) name579 (
		_w626_,
		_w629_,
		_w630_
	);
	LUT2 #(
		.INIT('h4)
	) name580 (
		_w627_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h4)
	) name581 (
		_w446_,
		_w454_,
		_w632_
	);
	LUT2 #(
		.INIT('h2)
	) name582 (
		_w370_,
		_w455_,
		_w633_
	);
	LUT2 #(
		.INIT('h4)
	) name583 (
		_w632_,
		_w633_,
		_w634_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		_w593_,
		_w631_,
		_w635_
	);
	LUT2 #(
		.INIT('h4)
	) name585 (
		_w634_,
		_w635_,
		_w636_
	);
	LUT2 #(
		.INIT('h4)
	) name586 (
		_w351_,
		_w354_,
		_w637_
	);
	LUT2 #(
		.INIT('h1)
	) name587 (
		_w447_,
		_w637_,
		_w638_
	);
	LUT2 #(
		.INIT('h8)
	) name588 (
		_w433_,
		_w638_,
		_w639_
	);
	LUT2 #(
		.INIT('h1)
	) name589 (
		_w433_,
		_w638_,
		_w640_
	);
	LUT2 #(
		.INIT('h1)
	) name590 (
		_w371_,
		_w639_,
		_w641_
	);
	LUT2 #(
		.INIT('h4)
	) name591 (
		_w640_,
		_w641_,
		_w642_
	);
	LUT2 #(
		.INIT('h8)
	) name592 (
		\97(11)_pad ,
		_w382_,
		_w643_
	);
	LUT2 #(
		.INIT('h8)
	) name593 (
		\107(12)_pad ,
		_w394_,
		_w644_
	);
	LUT2 #(
		.INIT('h8)
	) name594 (
		\87(10)_pad ,
		_w396_,
		_w645_
	);
	LUT2 #(
		.INIT('h8)
	) name595 (
		\303(40)_pad ,
		_w377_,
		_w646_
	);
	LUT2 #(
		.INIT('h8)
	) name596 (
		\116(13)_pad ,
		_w389_,
		_w647_
	);
	LUT2 #(
		.INIT('h8)
	) name597 (
		\283(38)_pad ,
		_w391_,
		_w648_
	);
	LUT2 #(
		.INIT('h8)
	) name598 (
		\294(39)_pad ,
		_w385_,
		_w649_
	);
	LUT2 #(
		.INIT('h8)
	) name599 (
		\311(41)_pad ,
		_w387_,
		_w650_
	);
	LUT2 #(
		.INIT('h2)
	) name600 (
		\33(3)_pad ,
		_w643_,
		_w651_
	);
	LUT2 #(
		.INIT('h1)
	) name601 (
		_w644_,
		_w645_,
		_w652_
	);
	LUT2 #(
		.INIT('h1)
	) name602 (
		_w646_,
		_w647_,
		_w653_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		_w648_,
		_w649_,
		_w654_
	);
	LUT2 #(
		.INIT('h4)
	) name604 (
		_w650_,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h8)
	) name605 (
		_w652_,
		_w653_,
		_w656_
	);
	LUT2 #(
		.INIT('h8)
	) name606 (
		_w651_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h8)
	) name607 (
		_w655_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h8)
	) name608 (
		\137(18)_pad ,
		_w377_,
		_w659_
	);
	LUT2 #(
		.INIT('h8)
	) name609 (
		\50(6)_pad ,
		_w394_,
		_w660_
	);
	LUT2 #(
		.INIT('h8)
	) name610 (
		\143(19)_pad ,
		_w385_,
		_w661_
	);
	LUT2 #(
		.INIT('h8)
	) name611 (
		\132(17)_pad ,
		_w387_,
		_w662_
	);
	LUT2 #(
		.INIT('h8)
	) name612 (
		\58(7)_pad ,
		_w382_,
		_w663_
	);
	LUT2 #(
		.INIT('h8)
	) name613 (
		\150(20)_pad ,
		_w391_,
		_w664_
	);
	LUT2 #(
		.INIT('h8)
	) name614 (
		\159(21)_pad ,
		_w389_,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name615 (
		\33(3)_pad ,
		_w484_,
		_w666_
	);
	LUT2 #(
		.INIT('h1)
	) name616 (
		_w659_,
		_w660_,
		_w667_
	);
	LUT2 #(
		.INIT('h1)
	) name617 (
		_w661_,
		_w662_,
		_w668_
	);
	LUT2 #(
		.INIT('h1)
	) name618 (
		_w663_,
		_w664_,
		_w669_
	);
	LUT2 #(
		.INIT('h4)
	) name619 (
		_w665_,
		_w669_,
		_w670_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		_w667_,
		_w668_,
		_w671_
	);
	LUT2 #(
		.INIT('h8)
	) name621 (
		_w666_,
		_w671_,
		_w672_
	);
	LUT2 #(
		.INIT('h8)
	) name622 (
		_w670_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h1)
	) name623 (
		_w658_,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h2)
	) name624 (
		_w373_,
		_w674_,
		_w675_
	);
	LUT2 #(
		.INIT('h8)
	) name625 (
		_w101_,
		_w354_,
		_w676_
	);
	LUT2 #(
		.INIT('h4)
	) name626 (
		\77(9)_pad ,
		_w428_,
		_w677_
	);
	LUT2 #(
		.INIT('h2)
	) name627 (
		_w371_,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h4)
	) name628 (
		_w675_,
		_w678_,
		_w679_
	);
	LUT2 #(
		.INIT('h4)
	) name629 (
		_w676_,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		_w642_,
		_w680_,
		_w681_
	);
	LUT2 #(
		.INIT('h4)
	) name631 (
		\13(1)_pad ,
		_w64_,
		_w682_
	);
	LUT2 #(
		.INIT('h2)
	) name632 (
		_w100_,
		_w184_,
		_w683_
	);
	LUT2 #(
		.INIT('h2)
	) name633 (
		_w335_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h8)
	) name634 (
		_w100_,
		_w185_,
		_w685_
	);
	LUT2 #(
		.INIT('h1)
	) name635 (
		_w684_,
		_w685_,
		_w686_
	);
	LUT2 #(
		.INIT('h8)
	) name636 (
		_w682_,
		_w686_,
		_w687_
	);
	LUT2 #(
		.INIT('h8)
	) name637 (
		\159(21)_pad ,
		_w391_,
		_w688_
	);
	LUT2 #(
		.INIT('h8)
	) name638 (
		\137(18)_pad ,
		_w387_,
		_w689_
	);
	LUT2 #(
		.INIT('h8)
	) name639 (
		\143(19)_pad ,
		_w377_,
		_w690_
	);
	LUT2 #(
		.INIT('h8)
	) name640 (
		\58(7)_pad ,
		_w394_,
		_w691_
	);
	LUT2 #(
		.INIT('h8)
	) name641 (
		\150(20)_pad ,
		_w385_,
		_w692_
	);
	LUT2 #(
		.INIT('h8)
	) name642 (
		\50(6)_pad ,
		_w389_,
		_w693_
	);
	LUT2 #(
		.INIT('h1)
	) name643 (
		\33(3)_pad ,
		_w413_,
		_w694_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		_w596_,
		_w688_,
		_w695_
	);
	LUT2 #(
		.INIT('h1)
	) name645 (
		_w689_,
		_w690_,
		_w696_
	);
	LUT2 #(
		.INIT('h1)
	) name646 (
		_w691_,
		_w692_,
		_w697_
	);
	LUT2 #(
		.INIT('h4)
	) name647 (
		_w693_,
		_w697_,
		_w698_
	);
	LUT2 #(
		.INIT('h8)
	) name648 (
		_w695_,
		_w696_,
		_w699_
	);
	LUT2 #(
		.INIT('h8)
	) name649 (
		_w694_,
		_w699_,
		_w700_
	);
	LUT2 #(
		.INIT('h8)
	) name650 (
		_w698_,
		_w700_,
		_w701_
	);
	LUT2 #(
		.INIT('h8)
	) name651 (
		\294(39)_pad ,
		_w391_,
		_w702_
	);
	LUT2 #(
		.INIT('h8)
	) name652 (
		\97(11)_pad ,
		_w396_,
		_w703_
	);
	LUT2 #(
		.INIT('h8)
	) name653 (
		\311(41)_pad ,
		_w377_,
		_w704_
	);
	LUT2 #(
		.INIT('h8)
	) name654 (
		\303(40)_pad ,
		_w385_,
		_w705_
	);
	LUT2 #(
		.INIT('h8)
	) name655 (
		\317(42)_pad ,
		_w387_,
		_w706_
	);
	LUT2 #(
		.INIT('h8)
	) name656 (
		\116(13)_pad ,
		_w394_,
		_w707_
	);
	LUT2 #(
		.INIT('h8)
	) name657 (
		\283(38)_pad ,
		_w389_,
		_w708_
	);
	LUT2 #(
		.INIT('h8)
	) name658 (
		\107(12)_pad ,
		_w382_,
		_w709_
	);
	LUT2 #(
		.INIT('h2)
	) name659 (
		\33(3)_pad ,
		_w702_,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name660 (
		_w703_,
		_w704_,
		_w711_
	);
	LUT2 #(
		.INIT('h1)
	) name661 (
		_w705_,
		_w706_,
		_w712_
	);
	LUT2 #(
		.INIT('h1)
	) name662 (
		_w707_,
		_w708_,
		_w713_
	);
	LUT2 #(
		.INIT('h4)
	) name663 (
		_w709_,
		_w713_,
		_w714_
	);
	LUT2 #(
		.INIT('h8)
	) name664 (
		_w711_,
		_w712_,
		_w715_
	);
	LUT2 #(
		.INIT('h8)
	) name665 (
		_w710_,
		_w715_,
		_w716_
	);
	LUT2 #(
		.INIT('h8)
	) name666 (
		_w714_,
		_w716_,
		_w717_
	);
	LUT2 #(
		.INIT('h1)
	) name667 (
		_w701_,
		_w717_,
		_w718_
	);
	LUT2 #(
		.INIT('h2)
	) name668 (
		_w373_,
		_w718_,
		_w719_
	);
	LUT2 #(
		.INIT('h1)
	) name669 (
		_w373_,
		_w682_,
		_w720_
	);
	LUT2 #(
		.INIT('h4)
	) name670 (
		\13(1)_pad ,
		_w56_,
		_w721_
	);
	LUT2 #(
		.INIT('h8)
	) name671 (
		_w523_,
		_w721_,
		_w722_
	);
	LUT2 #(
		.INIT('h2)
	) name672 (
		\87(10)_pad ,
		_w369_,
		_w723_
	);
	LUT2 #(
		.INIT('h2)
	) name673 (
		_w720_,
		_w723_,
		_w724_
	);
	LUT2 #(
		.INIT('h4)
	) name674 (
		_w722_,
		_w724_,
		_w725_
	);
	LUT2 #(
		.INIT('h2)
	) name675 (
		_w371_,
		_w725_,
		_w726_
	);
	LUT2 #(
		.INIT('h4)
	) name676 (
		_w719_,
		_w726_,
		_w727_
	);
	LUT2 #(
		.INIT('h4)
	) name677 (
		_w687_,
		_w727_,
		_w728_
	);
	LUT2 #(
		.INIT('h2)
	) name678 (
		_w100_,
		_w196_,
		_w729_
	);
	LUT2 #(
		.INIT('h2)
	) name679 (
		_w334_,
		_w729_,
		_w730_
	);
	LUT2 #(
		.INIT('h4)
	) name680 (
		_w211_,
		_w729_,
		_w731_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		_w730_,
		_w731_,
		_w732_
	);
	LUT2 #(
		.INIT('h2)
	) name682 (
		\330(46)_pad ,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h4)
	) name683 (
		_w100_,
		_w212_,
		_w734_
	);
	LUT2 #(
		.INIT('h4)
	) name684 (
		_w100_,
		_w233_,
		_w735_
	);
	LUT2 #(
		.INIT('h2)
	) name685 (
		_w100_,
		_w220_,
		_w736_
	);
	LUT2 #(
		.INIT('h1)
	) name686 (
		_w238_,
		_w736_,
		_w737_
	);
	LUT2 #(
		.INIT('h1)
	) name687 (
		_w233_,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h1)
	) name688 (
		_w735_,
		_w738_,
		_w739_
	);
	LUT2 #(
		.INIT('h1)
	) name689 (
		_w734_,
		_w739_,
		_w740_
	);
	LUT2 #(
		.INIT('h1)
	) name690 (
		_w233_,
		_w238_,
		_w741_
	);
	LUT2 #(
		.INIT('h8)
	) name691 (
		_w734_,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h1)
	) name692 (
		_w740_,
		_w742_,
		_w743_
	);
	LUT2 #(
		.INIT('h4)
	) name693 (
		_w733_,
		_w743_,
		_w744_
	);
	LUT2 #(
		.INIT('h2)
	) name694 (
		_w733_,
		_w743_,
		_w745_
	);
	LUT2 #(
		.INIT('h1)
	) name695 (
		_w744_,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h2)
	) name696 (
		_w434_,
		_w746_,
		_w747_
	);
	LUT2 #(
		.INIT('h4)
	) name697 (
		_w100_,
		_w269_,
		_w748_
	);
	LUT2 #(
		.INIT('h2)
	) name698 (
		_w100_,
		_w260_,
		_w749_
	);
	LUT2 #(
		.INIT('h1)
	) name699 (
		_w263_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h1)
	) name700 (
		_w269_,
		_w750_,
		_w751_
	);
	LUT2 #(
		.INIT('h1)
	) name701 (
		_w748_,
		_w751_,
		_w752_
	);
	LUT2 #(
		.INIT('h2)
	) name702 (
		_w733_,
		_w738_,
		_w753_
	);
	LUT2 #(
		.INIT('h1)
	) name703 (
		_w735_,
		_w753_,
		_w754_
	);
	LUT2 #(
		.INIT('h4)
	) name704 (
		_w742_,
		_w754_,
		_w755_
	);
	LUT2 #(
		.INIT('h2)
	) name705 (
		_w742_,
		_w754_,
		_w756_
	);
	LUT2 #(
		.INIT('h1)
	) name706 (
		_w755_,
		_w756_,
		_w757_
	);
	LUT2 #(
		.INIT('h2)
	) name707 (
		_w752_,
		_w757_,
		_w758_
	);
	LUT2 #(
		.INIT('h4)
	) name708 (
		_w752_,
		_w757_,
		_w759_
	);
	LUT2 #(
		.INIT('h1)
	) name709 (
		_w758_,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h2)
	) name710 (
		_w747_,
		_w760_,
		_w761_
	);
	LUT2 #(
		.INIT('h2)
	) name711 (
		_w434_,
		_w761_,
		_w762_
	);
	LUT2 #(
		.INIT('h2)
	) name712 (
		_w370_,
		_w762_,
		_w763_
	);
	LUT2 #(
		.INIT('h2)
	) name713 (
		_w367_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('h4)
	) name714 (
		_w751_,
		_w757_,
		_w765_
	);
	LUT2 #(
		.INIT('h1)
	) name715 (
		_w748_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h1)
	) name716 (
		_w686_,
		_w766_,
		_w767_
	);
	LUT2 #(
		.INIT('h8)
	) name717 (
		_w686_,
		_w766_,
		_w768_
	);
	LUT2 #(
		.INIT('h1)
	) name718 (
		_w767_,
		_w768_,
		_w769_
	);
	LUT2 #(
		.INIT('h4)
	) name719 (
		_w764_,
		_w769_,
		_w770_
	);
	LUT2 #(
		.INIT('h1)
	) name720 (
		_w728_,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('h1)
	) name721 (
		_w367_,
		_w760_,
		_w772_
	);
	LUT2 #(
		.INIT('h2)
	) name722 (
		\97(11)_pad ,
		_w369_,
		_w773_
	);
	LUT2 #(
		.INIT('h1)
	) name723 (
		\116(13)_pad ,
		_w255_,
		_w774_
	);
	LUT2 #(
		.INIT('h1)
	) name724 (
		_w571_,
		_w774_,
		_w775_
	);
	LUT2 #(
		.INIT('h8)
	) name725 (
		\87(10)_pad ,
		_w775_,
		_w776_
	);
	LUT2 #(
		.INIT('h1)
	) name726 (
		\87(10)_pad ,
		_w775_,
		_w777_
	);
	LUT2 #(
		.INIT('h1)
	) name727 (
		_w776_,
		_w777_,
		_w778_
	);
	LUT2 #(
		.INIT('h2)
	) name728 (
		_w721_,
		_w778_,
		_w779_
	);
	LUT2 #(
		.INIT('h2)
	) name729 (
		_w720_,
		_w773_,
		_w780_
	);
	LUT2 #(
		.INIT('h4)
	) name730 (
		_w779_,
		_w780_,
		_w781_
	);
	LUT2 #(
		.INIT('h8)
	) name731 (
		\116(13)_pad ,
		_w382_,
		_w782_
	);
	LUT2 #(
		.INIT('h8)
	) name732 (
		\294(39)_pad ,
		_w389_,
		_w783_
	);
	LUT2 #(
		.INIT('h8)
	) name733 (
		\322(43)_pad ,
		_w387_,
		_w784_
	);
	LUT2 #(
		.INIT('h8)
	) name734 (
		\283(38)_pad ,
		_w394_,
		_w785_
	);
	LUT2 #(
		.INIT('h8)
	) name735 (
		\107(12)_pad ,
		_w396_,
		_w786_
	);
	LUT2 #(
		.INIT('h8)
	) name736 (
		\317(42)_pad ,
		_w377_,
		_w787_
	);
	LUT2 #(
		.INIT('h8)
	) name737 (
		\311(41)_pad ,
		_w385_,
		_w788_
	);
	LUT2 #(
		.INIT('h8)
	) name738 (
		\303(40)_pad ,
		_w391_,
		_w789_
	);
	LUT2 #(
		.INIT('h2)
	) name739 (
		\33(3)_pad ,
		_w782_,
		_w790_
	);
	LUT2 #(
		.INIT('h1)
	) name740 (
		_w783_,
		_w784_,
		_w791_
	);
	LUT2 #(
		.INIT('h1)
	) name741 (
		_w785_,
		_w786_,
		_w792_
	);
	LUT2 #(
		.INIT('h1)
	) name742 (
		_w787_,
		_w788_,
		_w793_
	);
	LUT2 #(
		.INIT('h4)
	) name743 (
		_w789_,
		_w793_,
		_w794_
	);
	LUT2 #(
		.INIT('h8)
	) name744 (
		_w791_,
		_w792_,
		_w795_
	);
	LUT2 #(
		.INIT('h8)
	) name745 (
		_w790_,
		_w795_,
		_w796_
	);
	LUT2 #(
		.INIT('h8)
	) name746 (
		_w794_,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('h8)
	) name747 (
		\50(6)_pad ,
		_w391_,
		_w798_
	);
	LUT2 #(
		.INIT('h8)
	) name748 (
		\143(19)_pad ,
		_w387_,
		_w799_
	);
	LUT2 #(
		.INIT('h8)
	) name749 (
		\150(20)_pad ,
		_w377_,
		_w800_
	);
	LUT2 #(
		.INIT('h8)
	) name750 (
		\68(8)_pad ,
		_w394_,
		_w801_
	);
	LUT2 #(
		.INIT('h8)
	) name751 (
		\159(21)_pad ,
		_w385_,
		_w802_
	);
	LUT2 #(
		.INIT('h8)
	) name752 (
		\58(7)_pad ,
		_w389_,
		_w803_
	);
	LUT2 #(
		.INIT('h1)
	) name753 (
		\33(3)_pad ,
		_w489_,
		_w804_
	);
	LUT2 #(
		.INIT('h1)
	) name754 (
		_w645_,
		_w798_,
		_w805_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		_w799_,
		_w800_,
		_w806_
	);
	LUT2 #(
		.INIT('h1)
	) name756 (
		_w801_,
		_w802_,
		_w807_
	);
	LUT2 #(
		.INIT('h4)
	) name757 (
		_w803_,
		_w807_,
		_w808_
	);
	LUT2 #(
		.INIT('h8)
	) name758 (
		_w805_,
		_w806_,
		_w809_
	);
	LUT2 #(
		.INIT('h8)
	) name759 (
		_w804_,
		_w809_,
		_w810_
	);
	LUT2 #(
		.INIT('h8)
	) name760 (
		_w808_,
		_w810_,
		_w811_
	);
	LUT2 #(
		.INIT('h1)
	) name761 (
		_w797_,
		_w811_,
		_w812_
	);
	LUT2 #(
		.INIT('h2)
	) name762 (
		_w373_,
		_w812_,
		_w813_
	);
	LUT2 #(
		.INIT('h2)
	) name763 (
		_w682_,
		_w752_,
		_w814_
	);
	LUT2 #(
		.INIT('h2)
	) name764 (
		_w371_,
		_w781_,
		_w815_
	);
	LUT2 #(
		.INIT('h4)
	) name765 (
		_w813_,
		_w815_,
		_w816_
	);
	LUT2 #(
		.INIT('h4)
	) name766 (
		_w814_,
		_w816_,
		_w817_
	);
	LUT2 #(
		.INIT('h4)
	) name767 (
		_w747_,
		_w760_,
		_w818_
	);
	LUT2 #(
		.INIT('h2)
	) name768 (
		_w370_,
		_w761_,
		_w819_
	);
	LUT2 #(
		.INIT('h4)
	) name769 (
		_w818_,
		_w819_,
		_w820_
	);
	LUT2 #(
		.INIT('h1)
	) name770 (
		_w772_,
		_w817_,
		_w821_
	);
	LUT2 #(
		.INIT('h4)
	) name771 (
		_w820_,
		_w821_,
		_w822_
	);
	LUT2 #(
		.INIT('h1)
	) name772 (
		_w367_,
		_w746_,
		_w823_
	);
	LUT2 #(
		.INIT('h2)
	) name773 (
		_w682_,
		_w739_,
		_w824_
	);
	LUT2 #(
		.INIT('h1)
	) name774 (
		\107(12)_pad ,
		_w369_,
		_w825_
	);
	LUT2 #(
		.INIT('h4)
	) name775 (
		\33(3)_pad ,
		_w369_,
		_w826_
	);
	LUT2 #(
		.INIT('h4)
	) name776 (
		_w561_,
		_w826_,
		_w827_
	);
	LUT2 #(
		.INIT('h2)
	) name777 (
		\45(5)_pad ,
		_w532_,
		_w828_
	);
	LUT2 #(
		.INIT('h8)
	) name778 (
		\68(8)_pad ,
		\77(9)_pad ,
		_w829_
	);
	LUT2 #(
		.INIT('h1)
	) name779 (
		\45(5)_pad ,
		\50(6)_pad ,
		_w830_
	);
	LUT2 #(
		.INIT('h8)
	) name780 (
		\58(7)_pad ,
		_w830_,
		_w831_
	);
	LUT2 #(
		.INIT('h4)
	) name781 (
		_w829_,
		_w831_,
		_w832_
	);
	LUT2 #(
		.INIT('h8)
	) name782 (
		_w561_,
		_w832_,
		_w833_
	);
	LUT2 #(
		.INIT('h2)
	) name783 (
		_w721_,
		_w833_,
		_w834_
	);
	LUT2 #(
		.INIT('h4)
	) name784 (
		_w828_,
		_w834_,
		_w835_
	);
	LUT2 #(
		.INIT('h1)
	) name785 (
		_w825_,
		_w827_,
		_w836_
	);
	LUT2 #(
		.INIT('h4)
	) name786 (
		_w835_,
		_w836_,
		_w837_
	);
	LUT2 #(
		.INIT('h2)
	) name787 (
		_w720_,
		_w837_,
		_w838_
	);
	LUT2 #(
		.INIT('h8)
	) name788 (
		\150(20)_pad ,
		_w387_,
		_w839_
	);
	LUT2 #(
		.INIT('h8)
	) name789 (
		\50(6)_pad ,
		_w385_,
		_w840_
	);
	LUT2 #(
		.INIT('h8)
	) name790 (
		\68(8)_pad ,
		_w389_,
		_w841_
	);
	LUT2 #(
		.INIT('h8)
	) name791 (
		\58(7)_pad ,
		_w391_,
		_w842_
	);
	LUT2 #(
		.INIT('h8)
	) name792 (
		\159(21)_pad ,
		_w377_,
		_w843_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		\33(3)_pad ,
		_w409_,
		_w844_
	);
	LUT2 #(
		.INIT('h1)
	) name794 (
		_w594_,
		_w703_,
		_w845_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		_w839_,
		_w840_,
		_w846_
	);
	LUT2 #(
		.INIT('h1)
	) name796 (
		_w841_,
		_w842_,
		_w847_
	);
	LUT2 #(
		.INIT('h4)
	) name797 (
		_w843_,
		_w847_,
		_w848_
	);
	LUT2 #(
		.INIT('h8)
	) name798 (
		_w845_,
		_w846_,
		_w849_
	);
	LUT2 #(
		.INIT('h8)
	) name799 (
		_w844_,
		_w849_,
		_w850_
	);
	LUT2 #(
		.INIT('h8)
	) name800 (
		_w848_,
		_w850_,
		_w851_
	);
	LUT2 #(
		.INIT('h8)
	) name801 (
		\303(40)_pad ,
		_w389_,
		_w852_
	);
	LUT2 #(
		.INIT('h8)
	) name802 (
		\116(13)_pad ,
		_w396_,
		_w853_
	);
	LUT2 #(
		.INIT('h8)
	) name803 (
		\317(42)_pad ,
		_w385_,
		_w854_
	);
	LUT2 #(
		.INIT('h8)
	) name804 (
		\326(44)_pad ,
		_w387_,
		_w855_
	);
	LUT2 #(
		.INIT('h8)
	) name805 (
		\283(38)_pad ,
		_w382_,
		_w856_
	);
	LUT2 #(
		.INIT('h8)
	) name806 (
		\294(39)_pad ,
		_w394_,
		_w857_
	);
	LUT2 #(
		.INIT('h8)
	) name807 (
		\322(43)_pad ,
		_w377_,
		_w858_
	);
	LUT2 #(
		.INIT('h8)
	) name808 (
		\311(41)_pad ,
		_w391_,
		_w859_
	);
	LUT2 #(
		.INIT('h2)
	) name809 (
		\33(3)_pad ,
		_w852_,
		_w860_
	);
	LUT2 #(
		.INIT('h1)
	) name810 (
		_w853_,
		_w854_,
		_w861_
	);
	LUT2 #(
		.INIT('h1)
	) name811 (
		_w855_,
		_w856_,
		_w862_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		_w857_,
		_w858_,
		_w863_
	);
	LUT2 #(
		.INIT('h4)
	) name813 (
		_w859_,
		_w863_,
		_w864_
	);
	LUT2 #(
		.INIT('h8)
	) name814 (
		_w861_,
		_w862_,
		_w865_
	);
	LUT2 #(
		.INIT('h8)
	) name815 (
		_w860_,
		_w865_,
		_w866_
	);
	LUT2 #(
		.INIT('h8)
	) name816 (
		_w864_,
		_w866_,
		_w867_
	);
	LUT2 #(
		.INIT('h1)
	) name817 (
		_w851_,
		_w867_,
		_w868_
	);
	LUT2 #(
		.INIT('h2)
	) name818 (
		_w373_,
		_w868_,
		_w869_
	);
	LUT2 #(
		.INIT('h2)
	) name819 (
		_w371_,
		_w838_,
		_w870_
	);
	LUT2 #(
		.INIT('h4)
	) name820 (
		_w869_,
		_w870_,
		_w871_
	);
	LUT2 #(
		.INIT('h4)
	) name821 (
		_w824_,
		_w871_,
		_w872_
	);
	LUT2 #(
		.INIT('h4)
	) name822 (
		_w434_,
		_w746_,
		_w873_
	);
	LUT2 #(
		.INIT('h2)
	) name823 (
		_w370_,
		_w747_,
		_w874_
	);
	LUT2 #(
		.INIT('h4)
	) name824 (
		_w873_,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h1)
	) name825 (
		_w823_,
		_w872_,
		_w876_
	);
	LUT2 #(
		.INIT('h4)
	) name826 (
		_w875_,
		_w876_,
		_w877_
	);
	LUT2 #(
		.INIT('h4)
	) name827 (
		\330(46)_pad ,
		_w732_,
		_w878_
	);
	LUT2 #(
		.INIT('h1)
	) name828 (
		_w371_,
		_w733_,
		_w879_
	);
	LUT2 #(
		.INIT('h4)
	) name829 (
		_w878_,
		_w879_,
		_w880_
	);
	LUT2 #(
		.INIT('h8)
	) name830 (
		_w682_,
		_w732_,
		_w881_
	);
	LUT2 #(
		.INIT('h8)
	) name831 (
		\322(43)_pad ,
		_w385_,
		_w882_
	);
	LUT2 #(
		.INIT('h8)
	) name832 (
		\294(39)_pad ,
		_w382_,
		_w883_
	);
	LUT2 #(
		.INIT('h8)
	) name833 (
		\329(45)_pad ,
		_w387_,
		_w884_
	);
	LUT2 #(
		.INIT('h8)
	) name834 (
		\317(42)_pad ,
		_w391_,
		_w885_
	);
	LUT2 #(
		.INIT('h8)
	) name835 (
		\311(41)_pad ,
		_w389_,
		_w886_
	);
	LUT2 #(
		.INIT('h8)
	) name836 (
		\303(40)_pad ,
		_w394_,
		_w887_
	);
	LUT2 #(
		.INIT('h8)
	) name837 (
		\326(44)_pad ,
		_w377_,
		_w888_
	);
	LUT2 #(
		.INIT('h8)
	) name838 (
		\283(38)_pad ,
		_w396_,
		_w889_
	);
	LUT2 #(
		.INIT('h2)
	) name839 (
		\33(3)_pad ,
		_w882_,
		_w890_
	);
	LUT2 #(
		.INIT('h1)
	) name840 (
		_w883_,
		_w884_,
		_w891_
	);
	LUT2 #(
		.INIT('h1)
	) name841 (
		_w885_,
		_w886_,
		_w892_
	);
	LUT2 #(
		.INIT('h1)
	) name842 (
		_w887_,
		_w888_,
		_w893_
	);
	LUT2 #(
		.INIT('h4)
	) name843 (
		_w889_,
		_w893_,
		_w894_
	);
	LUT2 #(
		.INIT('h8)
	) name844 (
		_w891_,
		_w892_,
		_w895_
	);
	LUT2 #(
		.INIT('h8)
	) name845 (
		_w890_,
		_w895_,
		_w896_
	);
	LUT2 #(
		.INIT('h8)
	) name846 (
		_w894_,
		_w896_,
		_w897_
	);
	LUT2 #(
		.INIT('h8)
	) name847 (
		\159(21)_pad ,
		_w387_,
		_w898_
	);
	LUT2 #(
		.INIT('h8)
	) name848 (
		\68(8)_pad ,
		_w391_,
		_w899_
	);
	LUT2 #(
		.INIT('h8)
	) name849 (
		\58(7)_pad ,
		_w385_,
		_w900_
	);
	LUT2 #(
		.INIT('h8)
	) name850 (
		\77(9)_pad ,
		_w389_,
		_w901_
	);
	LUT2 #(
		.INIT('h8)
	) name851 (
		\50(6)_pad ,
		_w377_,
		_w902_
	);
	LUT2 #(
		.INIT('h1)
	) name852 (
		\33(3)_pad ,
		_w485_,
		_w903_
	);
	LUT2 #(
		.INIT('h1)
	) name853 (
		_w643_,
		_w786_,
		_w904_
	);
	LUT2 #(
		.INIT('h1)
	) name854 (
		_w898_,
		_w899_,
		_w905_
	);
	LUT2 #(
		.INIT('h1)
	) name855 (
		_w900_,
		_w901_,
		_w906_
	);
	LUT2 #(
		.INIT('h4)
	) name856 (
		_w902_,
		_w906_,
		_w907_
	);
	LUT2 #(
		.INIT('h8)
	) name857 (
		_w904_,
		_w905_,
		_w908_
	);
	LUT2 #(
		.INIT('h8)
	) name858 (
		_w903_,
		_w908_,
		_w909_
	);
	LUT2 #(
		.INIT('h8)
	) name859 (
		_w907_,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h1)
	) name860 (
		_w897_,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h2)
	) name861 (
		_w373_,
		_w911_,
		_w912_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		\116(13)_pad ,
		_w369_,
		_w913_
	);
	LUT2 #(
		.INIT('h4)
	) name863 (
		_w514_,
		_w826_,
		_w914_
	);
	LUT2 #(
		.INIT('h4)
	) name864 (
		\45(5)_pad ,
		_w552_,
		_w915_
	);
	LUT2 #(
		.INIT('h1)
	) name865 (
		_w512_,
		_w567_,
		_w916_
	);
	LUT2 #(
		.INIT('h2)
	) name866 (
		_w62_,
		_w916_,
		_w917_
	);
	LUT2 #(
		.INIT('h4)
	) name867 (
		_w62_,
		_w916_,
		_w918_
	);
	LUT2 #(
		.INIT('h1)
	) name868 (
		_w917_,
		_w918_,
		_w919_
	);
	LUT2 #(
		.INIT('h8)
	) name869 (
		\45(5)_pad ,
		_w919_,
		_w920_
	);
	LUT2 #(
		.INIT('h2)
	) name870 (
		_w721_,
		_w915_,
		_w921_
	);
	LUT2 #(
		.INIT('h4)
	) name871 (
		_w920_,
		_w921_,
		_w922_
	);
	LUT2 #(
		.INIT('h1)
	) name872 (
		_w913_,
		_w914_,
		_w923_
	);
	LUT2 #(
		.INIT('h4)
	) name873 (
		_w922_,
		_w923_,
		_w924_
	);
	LUT2 #(
		.INIT('h2)
	) name874 (
		_w720_,
		_w924_,
		_w925_
	);
	LUT2 #(
		.INIT('h2)
	) name875 (
		_w371_,
		_w925_,
		_w926_
	);
	LUT2 #(
		.INIT('h4)
	) name876 (
		_w912_,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h4)
	) name877 (
		_w881_,
		_w927_,
		_w928_
	);
	LUT2 #(
		.INIT('h1)
	) name878 (
		_w880_,
		_w928_,
		_w929_
	);
	LUT2 #(
		.INIT('h1)
	) name879 (
		_w466_,
		_w511_,
		_w930_
	);
	LUT2 #(
		.INIT('h8)
	) name880 (
		_w466_,
		_w511_,
		_w931_
	);
	LUT2 #(
		.INIT('h1)
	) name881 (
		_w930_,
		_w931_,
		_w932_
	);
	LUT2 #(
		.INIT('h2)
	) name882 (
		_w877_,
		_w929_,
		_w933_
	);
	LUT2 #(
		.INIT('h4)
	) name883 (
		_w877_,
		_w929_,
		_w934_
	);
	LUT2 #(
		.INIT('h1)
	) name884 (
		_w933_,
		_w934_,
		_w935_
	);
	LUT2 #(
		.INIT('h8)
	) name885 (
		_w771_,
		_w935_,
		_w936_
	);
	LUT2 #(
		.INIT('h1)
	) name886 (
		_w771_,
		_w935_,
		_w937_
	);
	LUT2 #(
		.INIT('h1)
	) name887 (
		_w936_,
		_w937_,
		_w938_
	);
	LUT2 #(
		.INIT('h4)
	) name888 (
		_w636_,
		_w681_,
		_w939_
	);
	LUT2 #(
		.INIT('h2)
	) name889 (
		_w636_,
		_w681_,
		_w940_
	);
	LUT2 #(
		.INIT('h1)
	) name890 (
		_w939_,
		_w940_,
		_w941_
	);
	LUT2 #(
		.INIT('h2)
	) name891 (
		_w822_,
		_w941_,
		_w942_
	);
	LUT2 #(
		.INIT('h4)
	) name892 (
		_w822_,
		_w941_,
		_w943_
	);
	LUT2 #(
		.INIT('h1)
	) name893 (
		_w942_,
		_w943_,
		_w944_
	);
	LUT2 #(
		.INIT('h8)
	) name894 (
		_w938_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h1)
	) name895 (
		_w938_,
		_w944_,
		_w946_
	);
	LUT2 #(
		.INIT('h1)
	) name896 (
		_w945_,
		_w946_,
		_w947_
	);
	LUT2 #(
		.INIT('h8)
	) name897 (
		_w932_,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h1)
	) name898 (
		_w932_,
		_w947_,
		_w949_
	);
	LUT2 #(
		.INIT('h1)
	) name899 (
		_w948_,
		_w949_,
		_w950_
	);
	LUT2 #(
		.INIT('h2)
	) name900 (
		\213(26)_pad ,
		\343(47)_pad ,
		_w951_
	);
	LUT2 #(
		.INIT('h1)
	) name901 (
		_w932_,
		_w951_,
		_w952_
	);
	LUT2 #(
		.INIT('h4)
	) name902 (
		\2897(49)_pad ,
		_w951_,
		_w953_
	);
	LUT2 #(
		.INIT('h1)
	) name903 (
		_w952_,
		_w953_,
		_w954_
	);
	LUT2 #(
		.INIT('h8)
	) name904 (
		_w947_,
		_w954_,
		_w955_
	);
	LUT2 #(
		.INIT('h1)
	) name905 (
		_w947_,
		_w954_,
		_w956_
	);
	LUT2 #(
		.INIT('h1)
	) name906 (
		_w955_,
		_w956_,
		_w957_
	);
	LUT2 #(
		.INIT('h8)
	) name907 (
		_w681_,
		_w929_,
		_w958_
	);
	LUT2 #(
		.INIT('h8)
	) name908 (
		_w877_,
		_w958_,
		_w959_
	);
	LUT2 #(
		.INIT('h8)
	) name909 (
		_w636_,
		_w959_,
		_w960_
	);
	LUT2 #(
		.INIT('h8)
	) name910 (
		_w822_,
		_w960_,
		_w961_
	);
	LUT2 #(
		.INIT('h8)
	) name911 (
		_w771_,
		_w961_,
		_w962_
	);
	LUT2 #(
		.INIT('h8)
	) name912 (
		_w931_,
		_w962_,
		_w963_
	);
	LUT2 #(
		.INIT('h8)
	) name913 (
		_w931_,
		_w951_,
		_w964_
	);
	LUT2 #(
		.INIT('h2)
	) name914 (
		\213(26)_pad ,
		_w963_,
		_w965_
	);
	LUT2 #(
		.INIT('h4)
	) name915 (
		_w964_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h8)
	) name916 (
		_w778_,
		_w919_,
		_w967_
	);
	LUT2 #(
		.INIT('h1)
	) name917 (
		_w778_,
		_w919_,
		_w968_
	);
	LUT2 #(
		.INIT('h1)
	) name918 (
		_w967_,
		_w968_,
		_w969_
	);
	assign \2690(1611)  = _w466_ ;
	assign \2709(1587)  = _w511_ ;
	assign \353(405)_pad  = _w513_ ;
	assign \355(399)_pad  = _w514_ ;
	assign \358(1161)_pad  = _w535_ ;
	assign \361(940)_pad  = _w558_ ;
	assign \364(1484)_pad  = _w565_ ;
	assign \367(1585)_pad  = _w589_ ;
	assign \369(1321)_pad  = _w591_ ;
	assign \372(1243)_pad  = _w592_ ;
	assign \381(1626)_pad  = _w636_ ;
	assign \384(1553)_pad  = _w681_ ;
	assign \387(1616)_pad  = _w771_ ;
	assign \390(1603)_pad  = _w822_ ;
	assign \393(1605)_pad  = _w877_ ;
	assign \396(1504)_pad  = _w929_ ;
	assign \399(1428)_pad  = _w755_ ;
	assign \402(1718)_pad  = _w950_ ;
	assign \404(1714)  = _w957_ ;
	assign \407(1657)_pad  = _w963_ ;
	assign \409(1670)_pad  = _w966_ ;
	assign \605(1186)  = _w969_ ;
endmodule;