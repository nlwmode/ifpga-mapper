module top (\CarrierSense_Tx2_reg/NET0131 , \Collision_Tx1_reg/NET0131 , \Collision_Tx2_reg/NET0131 , \RstTxPauseRq_reg/NET0131 , \RxAbortRst_reg/NET0131 , \RxAbort_latch_reg/NET0131 , \RxAbort_wb_reg/NET0131 , \RxEnSync_reg/NET0131 , \TPauseRq_reg/NET0131 , \TxPauseRq_sync2_reg/NET0131 , \TxPauseRq_sync3_reg/NET0131 , \WillSendControlFrame_sync2_reg/NET0131 , \WillSendControlFrame_sync3_reg/NET0131 , \WillTransmit_q2_reg/P0001 , \ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131 , \ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131 , \ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131 , \ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131 , \ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131 , \ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131 , \ethreg1_COLLCONF_2_DataOut_reg[0]/NET0131 , \ethreg1_COLLCONF_2_DataOut_reg[1]/NET0131 , \ethreg1_COLLCONF_2_DataOut_reg[2]/NET0131 , \ethreg1_COLLCONF_2_DataOut_reg[3]/NET0131 , \ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131 , \ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131 , \ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131 , \ethreg1_INT_MASK_0_DataOut_reg[0]/NET0131 , \ethreg1_INT_MASK_0_DataOut_reg[1]/NET0131 , \ethreg1_INT_MASK_0_DataOut_reg[2]/NET0131 , \ethreg1_INT_MASK_0_DataOut_reg[3]/NET0131 , \ethreg1_INT_MASK_0_DataOut_reg[4]/NET0131 , \ethreg1_INT_MASK_0_DataOut_reg[5]/NET0131 , \ethreg1_INT_MASK_0_DataOut_reg[6]/NET0131 , \ethreg1_IPGR1_0_DataOut_reg[0]/NET0131 , \ethreg1_IPGR1_0_DataOut_reg[1]/NET0131 , \ethreg1_IPGR1_0_DataOut_reg[2]/NET0131 , \ethreg1_IPGR1_0_DataOut_reg[3]/NET0131 , \ethreg1_IPGR1_0_DataOut_reg[4]/NET0131 , \ethreg1_IPGR1_0_DataOut_reg[5]/NET0131 , \ethreg1_IPGR1_0_DataOut_reg[6]/NET0131 , \ethreg1_IPGR2_0_DataOut_reg[0]/NET0131 , \ethreg1_IPGR2_0_DataOut_reg[1]/NET0131 , \ethreg1_IPGR2_0_DataOut_reg[2]/NET0131 , \ethreg1_IPGR2_0_DataOut_reg[3]/NET0131 , \ethreg1_IPGR2_0_DataOut_reg[4]/NET0131 , \ethreg1_IPGR2_0_DataOut_reg[5]/NET0131 , \ethreg1_IPGR2_0_DataOut_reg[6]/NET0131 , \ethreg1_IPGT_0_DataOut_reg[0]/NET0131 , \ethreg1_IPGT_0_DataOut_reg[1]/NET0131 , \ethreg1_IPGT_0_DataOut_reg[2]/NET0131 , \ethreg1_IPGT_0_DataOut_reg[3]/NET0131 , \ethreg1_IPGT_0_DataOut_reg[4]/NET0131 , \ethreg1_IPGT_0_DataOut_reg[5]/NET0131 , \ethreg1_IPGT_0_DataOut_reg[6]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131 , \ethreg1_MIIADDRESS_0_DataOut_reg[0]/NET0131 , \ethreg1_MIIADDRESS_0_DataOut_reg[1]/NET0131 , \ethreg1_MIIADDRESS_0_DataOut_reg[2]/NET0131 , \ethreg1_MIIADDRESS_0_DataOut_reg[3]/NET0131 , \ethreg1_MIIADDRESS_0_DataOut_reg[4]/NET0131 , \ethreg1_MIIADDRESS_1_DataOut_reg[0]/NET0131 , \ethreg1_MIIADDRESS_1_DataOut_reg[1]/NET0131 , \ethreg1_MIIADDRESS_1_DataOut_reg[2]/NET0131 , \ethreg1_MIIADDRESS_1_DataOut_reg[3]/NET0131 , \ethreg1_MIIADDRESS_1_DataOut_reg[4]/NET0131 , \ethreg1_MIICOMMAND0_DataOut_reg[0]/NET0131 , \ethreg1_MIICOMMAND1_DataOut_reg[0]/NET0131 , \ethreg1_MIICOMMAND2_DataOut_reg[0]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[0]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131 , \ethreg1_MIIMODER_1_DataOut_reg[0]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[0]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[10]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[11]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[12]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[13]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[14]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[15]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[1]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[2]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[3]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[4]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[5]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[6]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[7]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[8]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[9]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[0]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[1]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[2]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[3]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[4]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[5]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[6]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[7]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[0]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[1]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[2]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[3]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[4]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[5]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[6]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[7]/NET0131 , \ethreg1_MODER_0_DataOut_reg[0]/NET0131 , \ethreg1_MODER_0_DataOut_reg[1]/NET0131 , \ethreg1_MODER_0_DataOut_reg[2]/NET0131 , \ethreg1_MODER_0_DataOut_reg[3]/NET0131 , \ethreg1_MODER_0_DataOut_reg[4]/NET0131 , \ethreg1_MODER_0_DataOut_reg[5]/NET0131 , \ethreg1_MODER_0_DataOut_reg[6]/NET0131 , \ethreg1_MODER_0_DataOut_reg[7]/NET0131 , \ethreg1_MODER_1_DataOut_reg[0]/NET0131 , \ethreg1_MODER_1_DataOut_reg[1]/NET0131 , \ethreg1_MODER_1_DataOut_reg[2]/NET0131 , \ethreg1_MODER_1_DataOut_reg[3]/NET0131 , \ethreg1_MODER_1_DataOut_reg[4]/NET0131 , \ethreg1_MODER_1_DataOut_reg[5]/NET0131 , \ethreg1_MODER_1_DataOut_reg[6]/NET0131 , \ethreg1_MODER_1_DataOut_reg[7]/NET0131 , \ethreg1_MODER_2_DataOut_reg[0]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[7]/NET0131 , \ethreg1_ResetRxCIrq_sync2_reg/NET0131 , \ethreg1_ResetRxCIrq_sync3_reg/NET0131 , \ethreg1_ResetTxCIrq_sync2_reg/NET0131 , \ethreg1_SetRxCIrq_reg/NET0131 , \ethreg1_SetRxCIrq_rxclk_reg/NET0131 , \ethreg1_SetRxCIrq_sync2_reg/NET0131 , \ethreg1_SetRxCIrq_sync3_reg/NET0131 , \ethreg1_SetTxCIrq_reg/NET0131 , \ethreg1_SetTxCIrq_sync2_reg/NET0131 , \ethreg1_SetTxCIrq_sync3_reg/NET0131 , \ethreg1_SetTxCIrq_txclk_reg/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[0]/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[1]/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[2]/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[3]/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[4]/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[5]/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[6]/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[7]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[0]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[1]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[2]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[3]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[4]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[5]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[6]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[7]/NET0131 , \ethreg1_TXCTRL_2_DataOut_reg[0]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[0]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[1]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[2]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[3]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[4]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[5]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[6]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131 , \ethreg1_irq_busy_reg/NET0131 , \ethreg1_irq_rxb_reg/NET0131 , \ethreg1_irq_rxc_reg/NET0131 , \ethreg1_irq_rxe_reg/NET0131 , \ethreg1_irq_txb_reg/NET0131 , \ethreg1_irq_txc_reg/NET0131 , \ethreg1_irq_txe_reg/NET0131 , m_wb_ack_i_pad, \m_wb_adr_o[10]_pad , \m_wb_adr_o[11]_pad , \m_wb_adr_o[12]_pad , \m_wb_adr_o[13]_pad , \m_wb_adr_o[14]_pad , \m_wb_adr_o[15]_pad , \m_wb_adr_o[16]_pad , \m_wb_adr_o[17]_pad , \m_wb_adr_o[18]_pad , \m_wb_adr_o[19]_pad , \m_wb_adr_o[20]_pad , \m_wb_adr_o[21]_pad , \m_wb_adr_o[22]_pad , \m_wb_adr_o[23]_pad , \m_wb_adr_o[24]_pad , \m_wb_adr_o[25]_pad , \m_wb_adr_o[26]_pad , \m_wb_adr_o[27]_pad , \m_wb_adr_o[28]_pad , \m_wb_adr_o[29]_pad , \m_wb_adr_o[2]_pad , \m_wb_adr_o[30]_pad , \m_wb_adr_o[31]_pad , \m_wb_adr_o[3]_pad , \m_wb_adr_o[4]_pad , \m_wb_adr_o[5]_pad , \m_wb_adr_o[6]_pad , \m_wb_adr_o[7]_pad , \m_wb_adr_o[8]_pad , \m_wb_adr_o[9]_pad , \m_wb_dat_i[10]_pad , \m_wb_dat_i[11]_pad , \m_wb_dat_i[12]_pad , \m_wb_dat_i[13]_pad , \m_wb_dat_i[14]_pad , \m_wb_dat_i[15]_pad , \m_wb_dat_i[16]_pad , \m_wb_dat_i[17]_pad , \m_wb_dat_i[18]_pad , \m_wb_dat_i[19]_pad , \m_wb_dat_i[1]_pad , \m_wb_dat_i[20]_pad , \m_wb_dat_i[22]_pad , \m_wb_dat_i[23]_pad , \m_wb_dat_i[24]_pad , \m_wb_dat_i[25]_pad , \m_wb_dat_i[26]_pad , \m_wb_dat_i[27]_pad , \m_wb_dat_i[28]_pad , \m_wb_dat_i[29]_pad , \m_wb_dat_i[2]_pad , \m_wb_dat_i[30]_pad , \m_wb_dat_i[31]_pad , \m_wb_dat_i[3]_pad , \m_wb_dat_i[4]_pad , \m_wb_dat_i[5]_pad , \m_wb_dat_i[6]_pad , \m_wb_dat_i[7]_pad , \m_wb_dat_i[8]_pad , m_wb_err_i_pad, \m_wb_sel_o[0]_pad , \m_wb_sel_o[1]_pad , \m_wb_sel_o[2]_pad , \m_wb_sel_o[3]_pad , m_wb_stb_o_pad, m_wb_we_o_pad, \maccontrol1_MuxedAbort_reg/NET0131 , \maccontrol1_MuxedDone_reg/NET0131 , \maccontrol1_TxAbortInLatched_reg/NET0131 , \maccontrol1_TxDoneInLatched_reg/NET0131 , \maccontrol1_TxUsedDataOutDetected_reg/NET0131 , \maccontrol1_receivecontrol1_AddressOK_reg/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[0]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[10]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[11]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[12]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[13]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[14]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[15]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[1]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[2]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[3]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[4]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[5]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[6]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[7]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[8]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[9]/NET0131 , \maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 , \maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 , \maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 , \maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 , \maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131 , \maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131 , \maccontrol1_receivecontrol1_Divider2_reg/NET0131 , \maccontrol1_receivecontrol1_DlyCrcCnt_reg[0]/NET0131 , \maccontrol1_receivecontrol1_DlyCrcCnt_reg[1]/NET0131 , \maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[0]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[10]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[11]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[12]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[13]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[14]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[15]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[1]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[2]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[3]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[4]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[5]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[6]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[7]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[8]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[9]/NET0131 , \maccontrol1_receivecontrol1_OpCodeOK_reg/NET0131 , \maccontrol1_receivecontrol1_PauseTimerEq0_sync2_reg/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[11]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[12]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[14]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[15]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[1]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[5]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[8]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131 , \maccontrol1_receivecontrol1_Pause_reg/NET0131 , \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 , \maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131 , \maccontrol1_receivecontrol1_SlotTimer_reg[0]/NET0131 , \maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131 , \maccontrol1_receivecontrol1_SlotTimer_reg[2]/NET0131 , \maccontrol1_receivecontrol1_SlotTimer_reg[3]/NET0131 , \maccontrol1_receivecontrol1_SlotTimer_reg[4]/NET0131 , \maccontrol1_receivecontrol1_SlotTimer_reg[5]/NET0131 , \maccontrol1_receivecontrol1_TypeLengthOK_reg/NET0131 , \maccontrol1_transmitcontrol1_BlockTxDone_reg/NET0131 , \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 , \maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 , \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 , \maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 , \maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 , \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[0]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[1]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[2]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[3]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[4]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[5]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[6]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[7]/NET0131 , \maccontrol1_transmitcontrol1_ControlEnd_q_reg/P0001 , \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 , \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131 , \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[1]/NET0131 , \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131 , \maccontrol1_transmitcontrol1_SendingCtrlFrm_reg/NET0131 , \maccontrol1_transmitcontrol1_TxCtrlEndFrm_reg/NET0131 , \maccontrol1_transmitcontrol1_TxCtrlStartFrm_q_reg/P0001 , \maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 , \maccontrol1_transmitcontrol1_TxUsedDataIn_q_reg/NET0131 , \maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131 , \macstatus1_CarrierSenseLost_reg/NET0131 , \macstatus1_DeferLatched_reg/NET0131 , \macstatus1_DribbleNibble_reg/NET0131 , \macstatus1_InvalidSymbol_reg/NET0131 , \macstatus1_LatchedCrcError_reg/NET0131 , \macstatus1_LatchedMRxErr_reg/NET0131 , \macstatus1_LateCollLatched_reg/P0002 , \macstatus1_LoadRxStatus_reg/NET0131 , \macstatus1_ReceiveEnd_reg/NET0131 , \macstatus1_ReceivedPacketTooBig_reg/NET0131 , \macstatus1_RetryCntLatched_reg[0]/P0002 , \macstatus1_RetryCntLatched_reg[1]/P0002 , \macstatus1_RetryCntLatched_reg[2]/P0002 , \macstatus1_RetryCntLatched_reg[3]/P0002 , \macstatus1_RetryLimit_reg/P0002 , \macstatus1_RxColWindow_reg/NET0131 , \macstatus1_RxLateCollision_reg/NET0131 , \macstatus1_ShortFrame_reg/NET0131 , mcoll_pad_i_pad, md_pad_i_pad, mdc_pad_o_pad, \miim1_BitCounter_reg[0]/NET0131 , \miim1_BitCounter_reg[1]/NET0131 , \miim1_BitCounter_reg[2]/NET0131 , \miim1_BitCounter_reg[3]/NET0131 , \miim1_BitCounter_reg[4]/NET0131 , \miim1_BitCounter_reg[5]/NET0131 , \miim1_BitCounter_reg[6]/NET0131 , \miim1_EndBusy_reg/NET0131 , \miim1_InProgress_q1_reg/NET0131 , \miim1_InProgress_q2_reg/NET0131 , \miim1_InProgress_q3_reg/NET0131 , \miim1_InProgress_reg/NET0131 , \miim1_LatchByte0_d_reg/NET0131 , \miim1_LatchByte1_d_reg/NET0131 , \miim1_LatchByte_reg[0]/NET0131 , \miim1_LatchByte_reg[1]/NET0131 , \miim1_Nvalid_reg/NET0131 , \miim1_RStatStart_q1_reg/NET0131 , \miim1_RStatStart_q2_reg/NET0131 , \miim1_RStatStart_reg/NET0131 , \miim1_RStat_q2_reg/NET0131 , \miim1_RStat_q3_reg/NET0131 , \miim1_ScanStat_q2_reg/NET0131 , \miim1_SyncStatMdcEn_reg/NET0131 , \miim1_WCtrlDataStart_q1_reg/NET0131 , \miim1_WCtrlDataStart_q2_reg/NET0131 , \miim1_WCtrlDataStart_q_reg/NET0131 , \miim1_WCtrlDataStart_reg/NET0131 , \miim1_WCtrlData_q2_reg/NET0131 , \miim1_WCtrlData_q3_reg/NET0131 , \miim1_WriteOp_reg/NET0131 , \miim1_clkgen_Counter_reg[0]/NET0131 , \miim1_clkgen_Counter_reg[1]/NET0131 , \miim1_clkgen_Counter_reg[2]/NET0131 , \miim1_clkgen_Counter_reg[3]/NET0131 , \miim1_clkgen_Counter_reg[4]/NET0131 , \miim1_clkgen_Counter_reg[5]/NET0131 , \miim1_clkgen_Counter_reg[6]/NET0131 , \miim1_outctrl_Mdo_2d_reg/NET0131 , \miim1_shftrg_LinkFail_reg/NET0131 , \miim1_shftrg_ShiftReg_reg[0]/NET0131 , \miim1_shftrg_ShiftReg_reg[1]/NET0131 , \miim1_shftrg_ShiftReg_reg[2]/NET0131 , \miim1_shftrg_ShiftReg_reg[3]/NET0131 , \miim1_shftrg_ShiftReg_reg[4]/NET0131 , \miim1_shftrg_ShiftReg_reg[5]/NET0131 , \miim1_shftrg_ShiftReg_reg[6]/NET0131 , \miim1_shftrg_ShiftReg_reg[7]/NET0131 , \mrxd_pad_i[0]_pad , \mrxd_pad_i[1]_pad , \mrxd_pad_i[2]_pad , \mrxd_pad_i[3]_pad , mrxdv_pad_i_pad, mrxerr_pad_i_pad, \mtxd_pad_o[0]_pad , \mtxd_pad_o[1]_pad , \mtxd_pad_o[2]_pad , \mtxd_pad_o[3]_pad , mtxen_pad_o_pad, mtxerr_pad_o_pad, \rxethmac1_Broadcast_reg/NET0131 , \rxethmac1_CrcHashGood_reg/P0001 , \rxethmac1_CrcHash_reg[0]/P0001 , \rxethmac1_CrcHash_reg[1]/P0001 , \rxethmac1_CrcHash_reg[2]/P0001 , \rxethmac1_CrcHash_reg[3]/P0001 , \rxethmac1_CrcHash_reg[4]/P0001 , \rxethmac1_CrcHash_reg[5]/P0001 , \rxethmac1_DelayData_reg/NET0131 , \rxethmac1_LatchedByte_reg[0]/NET0131 , \rxethmac1_LatchedByte_reg[1]/NET0131 , \rxethmac1_LatchedByte_reg[2]/NET0131 , \rxethmac1_LatchedByte_reg[3]/NET0131 , \rxethmac1_LatchedByte_reg[4]/NET0131 , \rxethmac1_LatchedByte_reg[5]/NET0131 , \rxethmac1_LatchedByte_reg[6]/NET0131 , \rxethmac1_LatchedByte_reg[7]/NET0131 , \rxethmac1_Multicast_reg/NET0131 , \rxethmac1_RxData_d_reg[0]/NET0131 , \rxethmac1_RxData_d_reg[1]/NET0131 , \rxethmac1_RxData_d_reg[2]/NET0131 , \rxethmac1_RxData_d_reg[3]/NET0131 , \rxethmac1_RxData_d_reg[4]/NET0131 , \rxethmac1_RxData_d_reg[5]/NET0131 , \rxethmac1_RxData_d_reg[6]/NET0131 , \rxethmac1_RxData_d_reg[7]/NET0131 , \rxethmac1_RxData_reg[0]/NET0131 , \rxethmac1_RxData_reg[1]/NET0131 , \rxethmac1_RxData_reg[2]/NET0131 , \rxethmac1_RxData_reg[3]/NET0131 , \rxethmac1_RxData_reg[4]/NET0131 , \rxethmac1_RxData_reg[5]/NET0131 , \rxethmac1_RxData_reg[6]/NET0131 , \rxethmac1_RxData_reg[7]/NET0131 , \rxethmac1_RxEndFrm_d_reg/NET0131 , \rxethmac1_RxEndFrm_reg/NET0131 , \rxethmac1_RxStartFrm_reg/NET0131 , \rxethmac1_RxValid_reg/NET0131 , \rxethmac1_crcrx_Crc_reg[0]/NET0131 , \rxethmac1_crcrx_Crc_reg[10]/NET0131 , \rxethmac1_crcrx_Crc_reg[11]/NET0131 , \rxethmac1_crcrx_Crc_reg[12]/NET0131 , \rxethmac1_crcrx_Crc_reg[13]/NET0131 , \rxethmac1_crcrx_Crc_reg[14]/NET0131 , \rxethmac1_crcrx_Crc_reg[15]/NET0131 , \rxethmac1_crcrx_Crc_reg[16]/NET0131 , \rxethmac1_crcrx_Crc_reg[17]/NET0131 , \rxethmac1_crcrx_Crc_reg[18]/NET0131 , \rxethmac1_crcrx_Crc_reg[19]/NET0131 , \rxethmac1_crcrx_Crc_reg[1]/NET0131 , \rxethmac1_crcrx_Crc_reg[20]/NET0131 , \rxethmac1_crcrx_Crc_reg[21]/NET0131 , \rxethmac1_crcrx_Crc_reg[22]/NET0131 , \rxethmac1_crcrx_Crc_reg[23]/NET0131 , \rxethmac1_crcrx_Crc_reg[24]/NET0131 , \rxethmac1_crcrx_Crc_reg[25]/NET0131 , \rxethmac1_crcrx_Crc_reg[26]/NET0131 , \rxethmac1_crcrx_Crc_reg[27]/NET0131 , \rxethmac1_crcrx_Crc_reg[28]/NET0131 , \rxethmac1_crcrx_Crc_reg[29]/NET0131 , \rxethmac1_crcrx_Crc_reg[2]/NET0131 , \rxethmac1_crcrx_Crc_reg[30]/NET0131 , \rxethmac1_crcrx_Crc_reg[31]/NET0131 , \rxethmac1_crcrx_Crc_reg[3]/NET0131 , \rxethmac1_crcrx_Crc_reg[4]/NET0131 , \rxethmac1_crcrx_Crc_reg[5]/NET0131 , \rxethmac1_crcrx_Crc_reg[6]/NET0131 , \rxethmac1_crcrx_Crc_reg[7]/NET0131 , \rxethmac1_crcrx_Crc_reg[8]/NET0131 , \rxethmac1_crcrx_Crc_reg[9]/NET0131 , \rxethmac1_rxaddrcheck1_AddressMiss_reg/NET0131 , \rxethmac1_rxaddrcheck1_MulticastOK_reg/NET0131 , \rxethmac1_rxaddrcheck1_RxAbort_reg/NET0131 , \rxethmac1_rxaddrcheck1_UnicastOK_reg/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 , \rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 , \rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131 , \rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131 , \rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131 , \rxethmac1_rxcounters1_IFGCounter_reg[0]/NET0131 , \rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131 , \rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131 , \rxethmac1_rxcounters1_IFGCounter_reg[3]/NET0131 , \rxethmac1_rxcounters1_IFGCounter_reg[4]/NET0131 , \rxethmac1_rxstatem1_StateData0_reg/NET0131 , \rxethmac1_rxstatem1_StateData1_reg/NET0131 , \rxethmac1_rxstatem1_StateDrop_reg/NET0131 , \rxethmac1_rxstatem1_StateIdle_reg/NET0131 , \rxethmac1_rxstatem1_StatePreamble_reg/NET0131 , \rxethmac1_rxstatem1_StateSFD_reg/NET0131 , \txethmac1_ColWindow_reg/NET0131 , \txethmac1_PacketFinished_q_reg/NET0131 , \txethmac1_RetryCnt_reg[0]/NET0131 , \txethmac1_RetryCnt_reg[1]/NET0131 , \txethmac1_RetryCnt_reg[2]/NET0131 , \txethmac1_RetryCnt_reg[3]/NET0131 , \txethmac1_StatusLatch_reg/NET0131 , \txethmac1_StopExcessiveDeferOccured_reg/NET0131 , \txethmac1_TxAbort_reg/NET0131 , \txethmac1_TxDone_reg/NET0131 , \txethmac1_TxRetry_reg/NET0131 , \txethmac1_TxUsedData_reg/NET0131 , \txethmac1_random1_RandomLatched_reg[0]/NET0131 , \txethmac1_random1_RandomLatched_reg[1]/NET0131 , \txethmac1_random1_RandomLatched_reg[2]/NET0131 , \txethmac1_random1_RandomLatched_reg[3]/NET0131 , \txethmac1_random1_RandomLatched_reg[4]/NET0131 , \txethmac1_random1_RandomLatched_reg[5]/NET0131 , \txethmac1_random1_RandomLatched_reg[6]/NET0131 , \txethmac1_random1_RandomLatched_reg[7]/NET0131 , \txethmac1_random1_RandomLatched_reg[8]/NET0131 , \txethmac1_random1_RandomLatched_reg[9]/NET0131 , \txethmac1_random1_x_reg[1]/NET0131 , \txethmac1_random1_x_reg[2]/NET0131 , \txethmac1_random1_x_reg[3]/NET0131 , \txethmac1_random1_x_reg[4]/NET0131 , \txethmac1_random1_x_reg[5]/NET0131 , \txethmac1_random1_x_reg[6]/NET0131 , \txethmac1_random1_x_reg[7]/NET0131 , \txethmac1_random1_x_reg[8]/NET0131 , \txethmac1_random1_x_reg[9]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[10]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[11]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[13]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[14]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[15]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[7]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[8]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 , \txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131 , \txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131 , \txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[0]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[10]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[11]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[12]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[13]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[14]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[15]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[1]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[2]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[3]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[4]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[5]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[6]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[7]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[8]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[9]/NET0131 , \txethmac1_txcrc_Crc_reg[0]/NET0131 , \txethmac1_txcrc_Crc_reg[10]/NET0131 , \txethmac1_txcrc_Crc_reg[11]/NET0131 , \txethmac1_txcrc_Crc_reg[12]/NET0131 , \txethmac1_txcrc_Crc_reg[13]/NET0131 , \txethmac1_txcrc_Crc_reg[14]/NET0131 , \txethmac1_txcrc_Crc_reg[15]/NET0131 , \txethmac1_txcrc_Crc_reg[16]/NET0131 , \txethmac1_txcrc_Crc_reg[17]/NET0131 , \txethmac1_txcrc_Crc_reg[18]/NET0131 , \txethmac1_txcrc_Crc_reg[19]/NET0131 , \txethmac1_txcrc_Crc_reg[1]/NET0131 , \txethmac1_txcrc_Crc_reg[20]/NET0131 , \txethmac1_txcrc_Crc_reg[21]/NET0131 , \txethmac1_txcrc_Crc_reg[22]/NET0131 , \txethmac1_txcrc_Crc_reg[23]/NET0131 , \txethmac1_txcrc_Crc_reg[24]/NET0131 , \txethmac1_txcrc_Crc_reg[25]/NET0131 , \txethmac1_txcrc_Crc_reg[26]/NET0131 , \txethmac1_txcrc_Crc_reg[27]/NET0131 , \txethmac1_txcrc_Crc_reg[28]/NET0131 , \txethmac1_txcrc_Crc_reg[29]/NET0131 , \txethmac1_txcrc_Crc_reg[2]/NET0131 , \txethmac1_txcrc_Crc_reg[30]/NET0131 , \txethmac1_txcrc_Crc_reg[31]/NET0131 , \txethmac1_txcrc_Crc_reg[3]/NET0131 , \txethmac1_txcrc_Crc_reg[4]/NET0131 , \txethmac1_txcrc_Crc_reg[5]/NET0131 , \txethmac1_txcrc_Crc_reg[6]/NET0131 , \txethmac1_txcrc_Crc_reg[7]/NET0131 , \txethmac1_txcrc_Crc_reg[8]/NET0131 , \txethmac1_txcrc_Crc_reg[9]/NET0131 , \txethmac1_txstatem1_Rule1_reg/NET0131 , \txethmac1_txstatem1_StateBackOff_reg/NET0131 , \txethmac1_txstatem1_StateData_reg[0]/NET0131 , \txethmac1_txstatem1_StateData_reg[1]/NET0131 , \txethmac1_txstatem1_StateDefer_reg/NET0131 , \txethmac1_txstatem1_StateFCS_reg/NET0131 , \txethmac1_txstatem1_StateIPG_reg/NET0131 , \txethmac1_txstatem1_StateIdle_reg/NET0131 , \txethmac1_txstatem1_StateJam_q_reg/NET0131 , \txethmac1_txstatem1_StateJam_reg/NET0131 , \txethmac1_txstatem1_StatePAD_reg/NET0131 , \txethmac1_txstatem1_StatePreamble_reg/NET0131 , wb_ack_o_pad, \wb_adr_i[10]_pad , \wb_adr_i[11]_pad , \wb_adr_i[2]_pad , \wb_adr_i[3]_pad , \wb_adr_i[4]_pad , \wb_adr_i[5]_pad , \wb_adr_i[6]_pad , \wb_adr_i[7]_pad , \wb_adr_i[8]_pad , \wb_adr_i[9]_pad , wb_cyc_i_pad, \wb_dat_i[0]_pad , \wb_dat_i[10]_pad , \wb_dat_i[11]_pad , \wb_dat_i[12]_pad , \wb_dat_i[13]_pad , \wb_dat_i[14]_pad , \wb_dat_i[15]_pad , \wb_dat_i[16]_pad , \wb_dat_i[17]_pad , \wb_dat_i[18]_pad , \wb_dat_i[19]_pad , \wb_dat_i[1]_pad , \wb_dat_i[20]_pad , \wb_dat_i[21]_pad , \wb_dat_i[22]_pad , \wb_dat_i[23]_pad , \wb_dat_i[24]_pad , \wb_dat_i[25]_pad , \wb_dat_i[26]_pad , \wb_dat_i[27]_pad , \wb_dat_i[28]_pad , \wb_dat_i[29]_pad , \wb_dat_i[2]_pad , \wb_dat_i[30]_pad , \wb_dat_i[31]_pad , \wb_dat_i[3]_pad , \wb_dat_i[4]_pad , \wb_dat_i[5]_pad , \wb_dat_i[6]_pad , \wb_dat_i[7]_pad , \wb_dat_i[8]_pad , \wb_dat_i[9]_pad , wb_err_o_pad, wb_rst_i_pad, \wb_sel_i[0]_pad , \wb_sel_i[1]_pad , \wb_sel_i[2]_pad , \wb_sel_i[3]_pad , wb_stb_i_pad, wb_we_i_pad, \wishbone_BDRead_reg/NET0131 , \wishbone_BDWrite_reg[0]/NET0131 , \wishbone_BDWrite_reg[1]/NET0131 , \wishbone_BDWrite_reg[2]/NET0131 , \wishbone_BDWrite_reg[3]/NET0131 , \wishbone_BlockReadTxDataFromMemory_reg/NET0131 , \wishbone_BlockingIncrementTxPointer_reg/NET0131 , \wishbone_BlockingTxBDRead_reg/NET0131 , \wishbone_BlockingTxStatusWrite_reg/NET0131 , \wishbone_BlockingTxStatusWrite_sync2_reg/NET0131 , \wishbone_BlockingTxStatusWrite_sync3_reg/NET0131 , \wishbone_Busy_IRQ_rck_reg/NET0131 , \wishbone_Busy_IRQ_sync2_reg/P0001 , \wishbone_Busy_IRQ_sync3_reg/P0001 , \wishbone_Busy_IRQ_syncb2_reg/P0001 , \wishbone_Flop_reg/NET0131 , \wishbone_IncrTxPointer_reg/NET0131 , \wishbone_LastByteIn_reg/NET0131 , \wishbone_LastWord_reg/NET0131 , \wishbone_LatchValidBytes_q_reg/NET0131 , \wishbone_LatchValidBytes_reg/NET0131 , \wishbone_LatchedRxLength_reg[0]/NET0131 , \wishbone_LatchedRxLength_reg[10]/NET0131 , \wishbone_LatchedRxLength_reg[11]/NET0131 , \wishbone_LatchedRxLength_reg[12]/NET0131 , \wishbone_LatchedRxLength_reg[13]/NET0131 , \wishbone_LatchedRxLength_reg[14]/NET0131 , \wishbone_LatchedRxLength_reg[15]/NET0131 , \wishbone_LatchedRxLength_reg[1]/NET0131 , \wishbone_LatchedRxLength_reg[2]/NET0131 , \wishbone_LatchedRxLength_reg[3]/NET0131 , \wishbone_LatchedRxLength_reg[4]/NET0131 , \wishbone_LatchedRxLength_reg[5]/NET0131 , \wishbone_LatchedRxLength_reg[6]/NET0131 , \wishbone_LatchedRxLength_reg[7]/NET0131 , \wishbone_LatchedRxLength_reg[8]/NET0131 , \wishbone_LatchedRxLength_reg[9]/NET0131 , \wishbone_LatchedRxStartFrm_reg/NET0131 , \wishbone_LatchedTxLength_reg[0]/NET0131 , \wishbone_LatchedTxLength_reg[10]/NET0131 , \wishbone_LatchedTxLength_reg[11]/NET0131 , \wishbone_LatchedTxLength_reg[12]/NET0131 , \wishbone_LatchedTxLength_reg[13]/NET0131 , \wishbone_LatchedTxLength_reg[14]/NET0131 , \wishbone_LatchedTxLength_reg[15]/NET0131 , \wishbone_LatchedTxLength_reg[1]/NET0131 , \wishbone_LatchedTxLength_reg[2]/NET0131 , \wishbone_LatchedTxLength_reg[3]/NET0131 , \wishbone_LatchedTxLength_reg[4]/NET0131 , \wishbone_LatchedTxLength_reg[5]/NET0131 , \wishbone_LatchedTxLength_reg[6]/NET0131 , \wishbone_LatchedTxLength_reg[7]/NET0131 , \wishbone_LatchedTxLength_reg[8]/NET0131 , \wishbone_LatchedTxLength_reg[9]/NET0131 , \wishbone_MasterWbRX_reg/NET0131 , \wishbone_MasterWbTX_reg/NET0131 , \wishbone_ReadTxDataFromFifo_sync2_reg/NET0131 , \wishbone_ReadTxDataFromFifo_sync3_reg/NET0131 , \wishbone_ReadTxDataFromFifo_syncb2_reg/NET0131 , \wishbone_ReadTxDataFromFifo_syncb3_reg/NET0131 , \wishbone_ReadTxDataFromFifo_tck_reg/NET0131 , \wishbone_ReadTxDataFromMemory_reg/NET0131 , \wishbone_RxAbortLatched_reg/NET0131 , \wishbone_RxAbortSync2_reg/NET0131 , \wishbone_RxAbortSync3_reg/NET0131 , \wishbone_RxAbortSync4_reg/NET0131 , \wishbone_RxAbortSyncb2_reg/NET0131 , \wishbone_RxBDAddress_reg[1]/NET0131 , \wishbone_RxBDAddress_reg[2]/NET0131 , \wishbone_RxBDAddress_reg[3]/NET0131 , \wishbone_RxBDAddress_reg[4]/NET0131 , \wishbone_RxBDAddress_reg[5]/NET0131 , \wishbone_RxBDAddress_reg[6]/NET0131 , \wishbone_RxBDAddress_reg[7]/NET0131 , \wishbone_RxBDRead_reg/NET0131 , \wishbone_RxBDReady_reg/NET0131 , \wishbone_RxB_IRQ_reg/NET0131 , \wishbone_RxByteCnt_reg[0]/NET0131 , \wishbone_RxByteCnt_reg[1]/NET0131 , \wishbone_RxDataLatched1_reg[10]/NET0131 , \wishbone_RxDataLatched1_reg[11]/NET0131 , \wishbone_RxDataLatched1_reg[12]/NET0131 , \wishbone_RxDataLatched1_reg[13]/NET0131 , \wishbone_RxDataLatched1_reg[14]/NET0131 , \wishbone_RxDataLatched1_reg[15]/NET0131 , \wishbone_RxDataLatched1_reg[16]/NET0131 , \wishbone_RxDataLatched1_reg[17]/NET0131 , \wishbone_RxDataLatched1_reg[18]/NET0131 , \wishbone_RxDataLatched1_reg[19]/NET0131 , \wishbone_RxDataLatched1_reg[20]/NET0131 , \wishbone_RxDataLatched1_reg[21]/NET0131 , \wishbone_RxDataLatched1_reg[22]/NET0131 , \wishbone_RxDataLatched1_reg[23]/NET0131 , \wishbone_RxDataLatched1_reg[24]/NET0131 , \wishbone_RxDataLatched1_reg[25]/NET0131 , \wishbone_RxDataLatched1_reg[26]/NET0131 , \wishbone_RxDataLatched1_reg[27]/NET0131 , \wishbone_RxDataLatched1_reg[28]/NET0131 , \wishbone_RxDataLatched1_reg[29]/NET0131 , \wishbone_RxDataLatched1_reg[30]/NET0131 , \wishbone_RxDataLatched1_reg[31]/NET0131 , \wishbone_RxDataLatched1_reg[8]/NET0131 , \wishbone_RxDataLatched1_reg[9]/NET0131 , \wishbone_RxDataLatched2_reg[0]/NET0131 , \wishbone_RxDataLatched2_reg[10]/NET0131 , \wishbone_RxDataLatched2_reg[11]/NET0131 , \wishbone_RxDataLatched2_reg[12]/NET0131 , \wishbone_RxDataLatched2_reg[13]/NET0131 , \wishbone_RxDataLatched2_reg[14]/NET0131 , \wishbone_RxDataLatched2_reg[15]/NET0131 , \wishbone_RxDataLatched2_reg[16]/NET0131 , \wishbone_RxDataLatched2_reg[17]/NET0131 , \wishbone_RxDataLatched2_reg[18]/NET0131 , \wishbone_RxDataLatched2_reg[19]/NET0131 , \wishbone_RxDataLatched2_reg[1]/NET0131 , \wishbone_RxDataLatched2_reg[20]/NET0131 , \wishbone_RxDataLatched2_reg[21]/NET0131 , \wishbone_RxDataLatched2_reg[22]/NET0131 , \wishbone_RxDataLatched2_reg[23]/NET0131 , \wishbone_RxDataLatched2_reg[24]/NET0131 , \wishbone_RxDataLatched2_reg[25]/NET0131 , \wishbone_RxDataLatched2_reg[26]/NET0131 , \wishbone_RxDataLatched2_reg[27]/NET0131 , \wishbone_RxDataLatched2_reg[28]/NET0131 , \wishbone_RxDataLatched2_reg[29]/NET0131 , \wishbone_RxDataLatched2_reg[2]/NET0131 , \wishbone_RxDataLatched2_reg[30]/NET0131 , \wishbone_RxDataLatched2_reg[31]/NET0131 , \wishbone_RxDataLatched2_reg[3]/NET0131 , \wishbone_RxDataLatched2_reg[4]/NET0131 , \wishbone_RxDataLatched2_reg[5]/NET0131 , \wishbone_RxDataLatched2_reg[6]/NET0131 , \wishbone_RxDataLatched2_reg[7]/NET0131 , \wishbone_RxDataLatched2_reg[8]/NET0131 , \wishbone_RxDataLatched2_reg[9]/NET0131 , \wishbone_RxE_IRQ_reg/NET0131 , \wishbone_RxEn_needed_reg/NET0131 , \wishbone_RxEn_q_reg/NET0131 , \wishbone_RxEn_reg/NET0131 , \wishbone_RxEnableWindow_reg/NET0131 , \wishbone_RxOverrun_reg/NET0131 , \wishbone_RxPointerLSB_rst_reg[0]/NET0131 , \wishbone_RxPointerLSB_rst_reg[1]/NET0131 , \wishbone_RxPointerMSB_reg[10]/NET0131 , \wishbone_RxPointerMSB_reg[11]/NET0131 , \wishbone_RxPointerMSB_reg[12]/NET0131 , \wishbone_RxPointerMSB_reg[13]/NET0131 , \wishbone_RxPointerMSB_reg[14]/NET0131 , \wishbone_RxPointerMSB_reg[15]/NET0131 , \wishbone_RxPointerMSB_reg[16]/NET0131 , \wishbone_RxPointerMSB_reg[17]/NET0131 , \wishbone_RxPointerMSB_reg[18]/NET0131 , \wishbone_RxPointerMSB_reg[19]/NET0131 , \wishbone_RxPointerMSB_reg[20]/NET0131 , \wishbone_RxPointerMSB_reg[21]/NET0131 , \wishbone_RxPointerMSB_reg[22]/NET0131 , \wishbone_RxPointerMSB_reg[23]/NET0131 , \wishbone_RxPointerMSB_reg[24]/NET0131 , \wishbone_RxPointerMSB_reg[25]/NET0131 , \wishbone_RxPointerMSB_reg[26]/NET0131 , \wishbone_RxPointerMSB_reg[27]/NET0131 , \wishbone_RxPointerMSB_reg[28]/NET0131 , \wishbone_RxPointerMSB_reg[29]/NET0131 , \wishbone_RxPointerMSB_reg[2]/NET0131 , \wishbone_RxPointerMSB_reg[30]/NET0131 , \wishbone_RxPointerMSB_reg[31]/NET0131 , \wishbone_RxPointerMSB_reg[3]/NET0131 , \wishbone_RxPointerMSB_reg[4]/NET0131 , \wishbone_RxPointerMSB_reg[5]/NET0131 , \wishbone_RxPointerMSB_reg[6]/NET0131 , \wishbone_RxPointerMSB_reg[7]/NET0131 , \wishbone_RxPointerMSB_reg[8]/NET0131 , \wishbone_RxPointerMSB_reg[9]/NET0131 , \wishbone_RxPointerRead_reg/NET0131 , \wishbone_RxReady_reg/NET0131 , \wishbone_RxStatusInLatched_reg[0]/NET0131 , \wishbone_RxStatusInLatched_reg[1]/NET0131 , \wishbone_RxStatusInLatched_reg[2]/NET0131 , \wishbone_RxStatusInLatched_reg[3]/NET0131 , \wishbone_RxStatusInLatched_reg[4]/NET0131 , \wishbone_RxStatusInLatched_reg[5]/NET0131 , \wishbone_RxStatusInLatched_reg[6]/NET0131 , \wishbone_RxStatusInLatched_reg[7]/NET0131 , \wishbone_RxStatusInLatched_reg[8]/NET0131 , \wishbone_RxStatusWriteLatched_reg/NET0131 , \wishbone_RxStatusWriteLatched_sync2_reg/NET0131 , \wishbone_RxStatusWriteLatched_syncb2_reg/NET0131 , \wishbone_RxStatus_reg[13]/NET0131 , \wishbone_RxStatus_reg[14]/NET0131 , \wishbone_RxValidBytes_reg[0]/NET0131 , \wishbone_RxValidBytes_reg[1]/NET0131 , \wishbone_ShiftEndedSync1_reg/NET0131 , \wishbone_ShiftEndedSync2_reg/NET0131 , \wishbone_ShiftEndedSync3_reg/NET0131 , \wishbone_ShiftEndedSync_c1_reg/NET0131 , \wishbone_ShiftEndedSync_c2_reg/NET0131 , \wishbone_ShiftEnded_rck_reg/NET0131 , \wishbone_ShiftEnded_reg/NET0131 , \wishbone_ShiftWillEnd_reg/NET0131 , \wishbone_StartOccured_reg/NET0131 , \wishbone_SyncRxStartFrm_q2_reg/NET0131 , \wishbone_SyncRxStartFrm_q_reg/NET0131 , \wishbone_TxAbortPacketBlocked_reg/NET0131 , \wishbone_TxAbortPacket_NotCleared_reg/NET0131 , \wishbone_TxAbortPacket_reg/NET0131 , \wishbone_TxAbort_q_reg/NET0131 , \wishbone_TxAbort_wb_q_reg/NET0131 , \wishbone_TxAbort_wb_reg/NET0131 , \wishbone_TxBDAddress_reg[1]/NET0131 , \wishbone_TxBDAddress_reg[2]/NET0131 , \wishbone_TxBDAddress_reg[3]/NET0131 , \wishbone_TxBDAddress_reg[4]/NET0131 , \wishbone_TxBDAddress_reg[5]/NET0131 , \wishbone_TxBDAddress_reg[6]/NET0131 , \wishbone_TxBDAddress_reg[7]/NET0131 , \wishbone_TxBDRead_reg/NET0131 , \wishbone_TxBDReady_reg/NET0131 , \wishbone_TxB_IRQ_reg/NET0131 , \wishbone_TxByteCnt_reg[0]/NET0131 , \wishbone_TxByteCnt_reg[1]/NET0131 , \wishbone_TxDataLatched_reg[0]/NET0131 , \wishbone_TxDataLatched_reg[10]/NET0131 , \wishbone_TxDataLatched_reg[11]/NET0131 , \wishbone_TxDataLatched_reg[12]/NET0131 , \wishbone_TxDataLatched_reg[13]/NET0131 , \wishbone_TxDataLatched_reg[14]/NET0131 , \wishbone_TxDataLatched_reg[15]/NET0131 , \wishbone_TxDataLatched_reg[16]/NET0131 , \wishbone_TxDataLatched_reg[17]/NET0131 , \wishbone_TxDataLatched_reg[18]/NET0131 , \wishbone_TxDataLatched_reg[19]/NET0131 , \wishbone_TxDataLatched_reg[1]/NET0131 , \wishbone_TxDataLatched_reg[20]/NET0131 , \wishbone_TxDataLatched_reg[21]/NET0131 , \wishbone_TxDataLatched_reg[22]/NET0131 , \wishbone_TxDataLatched_reg[23]/NET0131 , \wishbone_TxDataLatched_reg[24]/NET0131 , \wishbone_TxDataLatched_reg[25]/NET0131 , \wishbone_TxDataLatched_reg[26]/NET0131 , \wishbone_TxDataLatched_reg[27]/NET0131 , \wishbone_TxDataLatched_reg[28]/NET0131 , \wishbone_TxDataLatched_reg[29]/NET0131 , \wishbone_TxDataLatched_reg[2]/NET0131 , \wishbone_TxDataLatched_reg[30]/NET0131 , \wishbone_TxDataLatched_reg[31]/NET0131 , \wishbone_TxDataLatched_reg[3]/NET0131 , \wishbone_TxDataLatched_reg[4]/NET0131 , \wishbone_TxDataLatched_reg[5]/NET0131 , \wishbone_TxDataLatched_reg[6]/NET0131 , \wishbone_TxDataLatched_reg[7]/NET0131 , \wishbone_TxDataLatched_reg[8]/NET0131 , \wishbone_TxDataLatched_reg[9]/NET0131 , \wishbone_TxData_reg[0]/NET0131 , \wishbone_TxData_reg[1]/NET0131 , \wishbone_TxData_reg[2]/NET0131 , \wishbone_TxData_reg[3]/NET0131 , \wishbone_TxData_reg[4]/NET0131 , \wishbone_TxData_reg[5]/NET0131 , \wishbone_TxData_reg[6]/NET0131 , \wishbone_TxData_reg[7]/NET0131 , \wishbone_TxDonePacketBlocked_reg/NET0131 , \wishbone_TxDonePacket_NotCleared_reg/NET0131 , \wishbone_TxDonePacket_reg/NET0131 , \wishbone_TxDone_wb_q_reg/NET0131 , \wishbone_TxDone_wb_reg/NET0131 , \wishbone_TxE_IRQ_reg/NET0131 , \wishbone_TxEn_needed_reg/NET0131 , \wishbone_TxEn_q_reg/NET0131 , \wishbone_TxEn_reg/NET0131 , \wishbone_TxEndFrm_reg/NET0131 , \wishbone_TxEndFrm_wb_reg/NET0131 , \wishbone_TxLength_reg[0]/NET0131 , \wishbone_TxLength_reg[10]/NET0131 , \wishbone_TxLength_reg[11]/NET0131 , \wishbone_TxLength_reg[12]/NET0131 , \wishbone_TxLength_reg[13]/NET0131 , \wishbone_TxLength_reg[14]/NET0131 , \wishbone_TxLength_reg[15]/NET0131 , \wishbone_TxLength_reg[1]/NET0131 , \wishbone_TxLength_reg[2]/NET0131 , \wishbone_TxLength_reg[3]/NET0131 , \wishbone_TxLength_reg[4]/NET0131 , \wishbone_TxLength_reg[5]/NET0131 , \wishbone_TxLength_reg[6]/NET0131 , \wishbone_TxLength_reg[7]/NET0131 , \wishbone_TxLength_reg[8]/NET0131 , \wishbone_TxLength_reg[9]/NET0131 , \wishbone_TxPointerLSB_reg[0]/NET0131 , \wishbone_TxPointerLSB_reg[1]/NET0131 , \wishbone_TxPointerLSB_rst_reg[0]/NET0131 , \wishbone_TxPointerLSB_rst_reg[1]/NET0131 , \wishbone_TxPointerMSB_reg[10]/NET0131 , \wishbone_TxPointerMSB_reg[11]/NET0131 , \wishbone_TxPointerMSB_reg[12]/NET0131 , \wishbone_TxPointerMSB_reg[13]/NET0131 , \wishbone_TxPointerMSB_reg[14]/NET0131 , \wishbone_TxPointerMSB_reg[15]/NET0131 , \wishbone_TxPointerMSB_reg[16]/NET0131 , \wishbone_TxPointerMSB_reg[17]/NET0131 , \wishbone_TxPointerMSB_reg[18]/NET0131 , \wishbone_TxPointerMSB_reg[19]/NET0131 , \wishbone_TxPointerMSB_reg[20]/NET0131 , \wishbone_TxPointerMSB_reg[21]/NET0131 , \wishbone_TxPointerMSB_reg[22]/NET0131 , \wishbone_TxPointerMSB_reg[23]/NET0131 , \wishbone_TxPointerMSB_reg[24]/NET0131 , \wishbone_TxPointerMSB_reg[25]/NET0131 , \wishbone_TxPointerMSB_reg[26]/NET0131 , \wishbone_TxPointerMSB_reg[27]/NET0131 , \wishbone_TxPointerMSB_reg[28]/NET0131 , \wishbone_TxPointerMSB_reg[29]/NET0131 , \wishbone_TxPointerMSB_reg[2]/NET0131 , \wishbone_TxPointerMSB_reg[30]/NET0131 , \wishbone_TxPointerMSB_reg[31]/NET0131 , \wishbone_TxPointerMSB_reg[3]/NET0131 , \wishbone_TxPointerMSB_reg[4]/NET0131 , \wishbone_TxPointerMSB_reg[5]/NET0131 , \wishbone_TxPointerMSB_reg[6]/NET0131 , \wishbone_TxPointerMSB_reg[7]/NET0131 , \wishbone_TxPointerMSB_reg[8]/NET0131 , \wishbone_TxPointerMSB_reg[9]/NET0131 , \wishbone_TxPointerRead_reg/NET0131 , \wishbone_TxRetryPacketBlocked_reg/NET0131 , \wishbone_TxRetryPacket_NotCleared_reg/NET0131 , \wishbone_TxRetryPacket_reg/NET0131 , \wishbone_TxRetry_q_reg/NET0131 , \wishbone_TxRetry_wb_q_reg/NET0131 , \wishbone_TxRetry_wb_reg/NET0131 , \wishbone_TxStartFrm_reg/NET0131 , \wishbone_TxStartFrm_sync2_reg/NET0131 , \wishbone_TxStartFrm_syncb2_reg/NET0131 , \wishbone_TxStartFrm_wb_reg/NET0131 , \wishbone_TxStatus_reg[11]/NET0131 , \wishbone_TxStatus_reg[12]/NET0131 , \wishbone_TxStatus_reg[13]/NET0131 , \wishbone_TxStatus_reg[14]/NET0131 , \wishbone_TxUnderRun_reg/NET0131 , \wishbone_TxUnderRun_sync1_reg/NET0131 , \wishbone_TxUnderRun_wb_reg/NET0131 , \wishbone_TxUsedData_q_reg/NET0131 , \wishbone_TxValidBytesLatched_reg[0]/NET0131 , \wishbone_TxValidBytesLatched_reg[1]/NET0131 , \wishbone_WB_ACK_O_reg/P0001 , \wishbone_WbEn_q_reg/NET0131 , \wishbone_WbEn_reg/NET0131 , \wishbone_WriteRxDataToFifoSync2_reg/NET0131 , \wishbone_WriteRxDataToFifoSync3_reg/NET0131 , \wishbone_WriteRxDataToFifo_reg/NET0131 , \wishbone_bd_ram_mem0_reg[0][0]/P0001 , \wishbone_bd_ram_mem0_reg[0][1]/P0001 , \wishbone_bd_ram_mem0_reg[0][2]/P0001 , \wishbone_bd_ram_mem0_reg[0][3]/P0001 , \wishbone_bd_ram_mem0_reg[0][4]/P0001 , \wishbone_bd_ram_mem0_reg[0][5]/P0001 , \wishbone_bd_ram_mem0_reg[0][6]/P0001 , \wishbone_bd_ram_mem0_reg[0][7]/P0001 , \wishbone_bd_ram_mem0_reg[100][0]/P0001 , \wishbone_bd_ram_mem0_reg[100][1]/P0001 , \wishbone_bd_ram_mem0_reg[100][2]/P0001 , \wishbone_bd_ram_mem0_reg[100][3]/P0001 , \wishbone_bd_ram_mem0_reg[100][4]/P0001 , \wishbone_bd_ram_mem0_reg[100][5]/P0001 , \wishbone_bd_ram_mem0_reg[100][6]/P0001 , \wishbone_bd_ram_mem0_reg[100][7]/P0001 , \wishbone_bd_ram_mem0_reg[101][0]/P0001 , \wishbone_bd_ram_mem0_reg[101][1]/P0001 , \wishbone_bd_ram_mem0_reg[101][2]/P0001 , \wishbone_bd_ram_mem0_reg[101][3]/P0001 , \wishbone_bd_ram_mem0_reg[101][4]/P0001 , \wishbone_bd_ram_mem0_reg[101][5]/P0001 , \wishbone_bd_ram_mem0_reg[101][6]/P0001 , \wishbone_bd_ram_mem0_reg[101][7]/P0001 , \wishbone_bd_ram_mem0_reg[102][0]/P0001 , \wishbone_bd_ram_mem0_reg[102][1]/P0001 , \wishbone_bd_ram_mem0_reg[102][2]/P0001 , \wishbone_bd_ram_mem0_reg[102][3]/P0001 , \wishbone_bd_ram_mem0_reg[102][4]/P0001 , \wishbone_bd_ram_mem0_reg[102][5]/P0001 , \wishbone_bd_ram_mem0_reg[102][6]/P0001 , \wishbone_bd_ram_mem0_reg[102][7]/P0001 , \wishbone_bd_ram_mem0_reg[103][0]/P0001 , \wishbone_bd_ram_mem0_reg[103][1]/P0001 , \wishbone_bd_ram_mem0_reg[103][2]/P0001 , \wishbone_bd_ram_mem0_reg[103][3]/P0001 , \wishbone_bd_ram_mem0_reg[103][4]/P0001 , \wishbone_bd_ram_mem0_reg[103][5]/P0001 , \wishbone_bd_ram_mem0_reg[103][6]/P0001 , \wishbone_bd_ram_mem0_reg[103][7]/P0001 , \wishbone_bd_ram_mem0_reg[104][0]/P0001 , \wishbone_bd_ram_mem0_reg[104][1]/P0001 , \wishbone_bd_ram_mem0_reg[104][2]/P0001 , \wishbone_bd_ram_mem0_reg[104][3]/P0001 , \wishbone_bd_ram_mem0_reg[104][4]/P0001 , \wishbone_bd_ram_mem0_reg[104][5]/P0001 , \wishbone_bd_ram_mem0_reg[104][6]/P0001 , \wishbone_bd_ram_mem0_reg[104][7]/P0001 , \wishbone_bd_ram_mem0_reg[105][0]/P0001 , \wishbone_bd_ram_mem0_reg[105][1]/P0001 , \wishbone_bd_ram_mem0_reg[105][2]/P0001 , \wishbone_bd_ram_mem0_reg[105][3]/P0001 , \wishbone_bd_ram_mem0_reg[105][4]/P0001 , \wishbone_bd_ram_mem0_reg[105][5]/P0001 , \wishbone_bd_ram_mem0_reg[105][6]/P0001 , \wishbone_bd_ram_mem0_reg[105][7]/P0001 , \wishbone_bd_ram_mem0_reg[106][0]/P0001 , \wishbone_bd_ram_mem0_reg[106][1]/P0001 , \wishbone_bd_ram_mem0_reg[106][2]/P0001 , \wishbone_bd_ram_mem0_reg[106][3]/P0001 , \wishbone_bd_ram_mem0_reg[106][4]/P0001 , \wishbone_bd_ram_mem0_reg[106][5]/P0001 , \wishbone_bd_ram_mem0_reg[106][6]/P0001 , \wishbone_bd_ram_mem0_reg[106][7]/P0001 , \wishbone_bd_ram_mem0_reg[107][0]/P0001 , \wishbone_bd_ram_mem0_reg[107][1]/P0001 , \wishbone_bd_ram_mem0_reg[107][2]/P0001 , \wishbone_bd_ram_mem0_reg[107][3]/P0001 , \wishbone_bd_ram_mem0_reg[107][4]/P0001 , \wishbone_bd_ram_mem0_reg[107][5]/P0001 , \wishbone_bd_ram_mem0_reg[107][6]/P0001 , \wishbone_bd_ram_mem0_reg[107][7]/P0001 , \wishbone_bd_ram_mem0_reg[108][0]/P0001 , \wishbone_bd_ram_mem0_reg[108][1]/P0001 , \wishbone_bd_ram_mem0_reg[108][2]/P0001 , \wishbone_bd_ram_mem0_reg[108][3]/P0001 , \wishbone_bd_ram_mem0_reg[108][4]/P0001 , \wishbone_bd_ram_mem0_reg[108][5]/P0001 , \wishbone_bd_ram_mem0_reg[108][6]/P0001 , \wishbone_bd_ram_mem0_reg[108][7]/P0001 , \wishbone_bd_ram_mem0_reg[109][0]/P0001 , \wishbone_bd_ram_mem0_reg[109][1]/P0001 , \wishbone_bd_ram_mem0_reg[109][2]/P0001 , \wishbone_bd_ram_mem0_reg[109][3]/P0001 , \wishbone_bd_ram_mem0_reg[109][4]/P0001 , \wishbone_bd_ram_mem0_reg[109][5]/P0001 , \wishbone_bd_ram_mem0_reg[109][6]/P0001 , \wishbone_bd_ram_mem0_reg[109][7]/P0001 , \wishbone_bd_ram_mem0_reg[10][0]/P0001 , \wishbone_bd_ram_mem0_reg[10][1]/P0001 , \wishbone_bd_ram_mem0_reg[10][2]/P0001 , \wishbone_bd_ram_mem0_reg[10][3]/P0001 , \wishbone_bd_ram_mem0_reg[10][4]/P0001 , \wishbone_bd_ram_mem0_reg[10][5]/P0001 , \wishbone_bd_ram_mem0_reg[10][6]/P0001 , \wishbone_bd_ram_mem0_reg[10][7]/P0001 , \wishbone_bd_ram_mem0_reg[110][0]/P0001 , \wishbone_bd_ram_mem0_reg[110][1]/P0001 , \wishbone_bd_ram_mem0_reg[110][2]/P0001 , \wishbone_bd_ram_mem0_reg[110][3]/P0001 , \wishbone_bd_ram_mem0_reg[110][4]/P0001 , \wishbone_bd_ram_mem0_reg[110][5]/P0001 , \wishbone_bd_ram_mem0_reg[110][6]/P0001 , \wishbone_bd_ram_mem0_reg[110][7]/P0001 , \wishbone_bd_ram_mem0_reg[111][0]/P0001 , \wishbone_bd_ram_mem0_reg[111][1]/P0001 , \wishbone_bd_ram_mem0_reg[111][2]/P0001 , \wishbone_bd_ram_mem0_reg[111][3]/P0001 , \wishbone_bd_ram_mem0_reg[111][4]/P0001 , \wishbone_bd_ram_mem0_reg[111][5]/P0001 , \wishbone_bd_ram_mem0_reg[111][6]/P0001 , \wishbone_bd_ram_mem0_reg[111][7]/P0001 , \wishbone_bd_ram_mem0_reg[112][0]/P0001 , \wishbone_bd_ram_mem0_reg[112][1]/P0001 , \wishbone_bd_ram_mem0_reg[112][2]/P0001 , \wishbone_bd_ram_mem0_reg[112][3]/P0001 , \wishbone_bd_ram_mem0_reg[112][4]/P0001 , \wishbone_bd_ram_mem0_reg[112][5]/P0001 , \wishbone_bd_ram_mem0_reg[112][6]/P0001 , \wishbone_bd_ram_mem0_reg[112][7]/P0001 , \wishbone_bd_ram_mem0_reg[113][0]/P0001 , \wishbone_bd_ram_mem0_reg[113][1]/P0001 , \wishbone_bd_ram_mem0_reg[113][2]/P0001 , \wishbone_bd_ram_mem0_reg[113][3]/P0001 , \wishbone_bd_ram_mem0_reg[113][4]/P0001 , \wishbone_bd_ram_mem0_reg[113][5]/P0001 , \wishbone_bd_ram_mem0_reg[113][6]/P0001 , \wishbone_bd_ram_mem0_reg[113][7]/P0001 , \wishbone_bd_ram_mem0_reg[114][0]/P0001 , \wishbone_bd_ram_mem0_reg[114][1]/P0001 , \wishbone_bd_ram_mem0_reg[114][2]/P0001 , \wishbone_bd_ram_mem0_reg[114][3]/P0001 , \wishbone_bd_ram_mem0_reg[114][4]/P0001 , \wishbone_bd_ram_mem0_reg[114][5]/P0001 , \wishbone_bd_ram_mem0_reg[114][6]/P0001 , \wishbone_bd_ram_mem0_reg[114][7]/P0001 , \wishbone_bd_ram_mem0_reg[115][0]/P0001 , \wishbone_bd_ram_mem0_reg[115][1]/P0001 , \wishbone_bd_ram_mem0_reg[115][2]/P0001 , \wishbone_bd_ram_mem0_reg[115][3]/P0001 , \wishbone_bd_ram_mem0_reg[115][4]/P0001 , \wishbone_bd_ram_mem0_reg[115][5]/P0001 , \wishbone_bd_ram_mem0_reg[115][6]/P0001 , \wishbone_bd_ram_mem0_reg[115][7]/P0001 , \wishbone_bd_ram_mem0_reg[116][0]/P0001 , \wishbone_bd_ram_mem0_reg[116][1]/P0001 , \wishbone_bd_ram_mem0_reg[116][2]/P0001 , \wishbone_bd_ram_mem0_reg[116][3]/P0001 , \wishbone_bd_ram_mem0_reg[116][4]/P0001 , \wishbone_bd_ram_mem0_reg[116][5]/P0001 , \wishbone_bd_ram_mem0_reg[116][6]/P0001 , \wishbone_bd_ram_mem0_reg[116][7]/P0001 , \wishbone_bd_ram_mem0_reg[117][0]/P0001 , \wishbone_bd_ram_mem0_reg[117][1]/P0001 , \wishbone_bd_ram_mem0_reg[117][2]/P0001 , \wishbone_bd_ram_mem0_reg[117][3]/P0001 , \wishbone_bd_ram_mem0_reg[117][4]/P0001 , \wishbone_bd_ram_mem0_reg[117][5]/P0001 , \wishbone_bd_ram_mem0_reg[117][6]/P0001 , \wishbone_bd_ram_mem0_reg[117][7]/P0001 , \wishbone_bd_ram_mem0_reg[118][0]/P0001 , \wishbone_bd_ram_mem0_reg[118][1]/P0001 , \wishbone_bd_ram_mem0_reg[118][2]/P0001 , \wishbone_bd_ram_mem0_reg[118][3]/P0001 , \wishbone_bd_ram_mem0_reg[118][4]/P0001 , \wishbone_bd_ram_mem0_reg[118][5]/P0001 , \wishbone_bd_ram_mem0_reg[118][6]/P0001 , \wishbone_bd_ram_mem0_reg[118][7]/P0001 , \wishbone_bd_ram_mem0_reg[119][0]/P0001 , \wishbone_bd_ram_mem0_reg[119][1]/P0001 , \wishbone_bd_ram_mem0_reg[119][2]/P0001 , \wishbone_bd_ram_mem0_reg[119][3]/P0001 , \wishbone_bd_ram_mem0_reg[119][4]/P0001 , \wishbone_bd_ram_mem0_reg[119][5]/P0001 , \wishbone_bd_ram_mem0_reg[119][6]/P0001 , \wishbone_bd_ram_mem0_reg[119][7]/P0001 , \wishbone_bd_ram_mem0_reg[11][0]/P0001 , \wishbone_bd_ram_mem0_reg[11][1]/P0001 , \wishbone_bd_ram_mem0_reg[11][2]/P0001 , \wishbone_bd_ram_mem0_reg[11][3]/P0001 , \wishbone_bd_ram_mem0_reg[11][4]/P0001 , \wishbone_bd_ram_mem0_reg[11][5]/P0001 , \wishbone_bd_ram_mem0_reg[11][6]/P0001 , \wishbone_bd_ram_mem0_reg[11][7]/P0001 , \wishbone_bd_ram_mem0_reg[120][0]/P0001 , \wishbone_bd_ram_mem0_reg[120][1]/P0001 , \wishbone_bd_ram_mem0_reg[120][2]/P0001 , \wishbone_bd_ram_mem0_reg[120][3]/P0001 , \wishbone_bd_ram_mem0_reg[120][4]/P0001 , \wishbone_bd_ram_mem0_reg[120][5]/P0001 , \wishbone_bd_ram_mem0_reg[120][6]/P0001 , \wishbone_bd_ram_mem0_reg[120][7]/P0001 , \wishbone_bd_ram_mem0_reg[121][0]/P0001 , \wishbone_bd_ram_mem0_reg[121][1]/P0001 , \wishbone_bd_ram_mem0_reg[121][2]/P0001 , \wishbone_bd_ram_mem0_reg[121][3]/P0001 , \wishbone_bd_ram_mem0_reg[121][4]/P0001 , \wishbone_bd_ram_mem0_reg[121][5]/P0001 , \wishbone_bd_ram_mem0_reg[121][6]/P0001 , \wishbone_bd_ram_mem0_reg[121][7]/P0001 , \wishbone_bd_ram_mem0_reg[122][0]/P0001 , \wishbone_bd_ram_mem0_reg[122][1]/P0001 , \wishbone_bd_ram_mem0_reg[122][2]/P0001 , \wishbone_bd_ram_mem0_reg[122][3]/P0001 , \wishbone_bd_ram_mem0_reg[122][4]/P0001 , \wishbone_bd_ram_mem0_reg[122][5]/P0001 , \wishbone_bd_ram_mem0_reg[122][6]/P0001 , \wishbone_bd_ram_mem0_reg[122][7]/P0001 , \wishbone_bd_ram_mem0_reg[123][0]/P0001 , \wishbone_bd_ram_mem0_reg[123][1]/P0001 , \wishbone_bd_ram_mem0_reg[123][2]/P0001 , \wishbone_bd_ram_mem0_reg[123][3]/P0001 , \wishbone_bd_ram_mem0_reg[123][4]/P0001 , \wishbone_bd_ram_mem0_reg[123][5]/P0001 , \wishbone_bd_ram_mem0_reg[123][6]/P0001 , \wishbone_bd_ram_mem0_reg[123][7]/P0001 , \wishbone_bd_ram_mem0_reg[124][0]/P0001 , \wishbone_bd_ram_mem0_reg[124][1]/P0001 , \wishbone_bd_ram_mem0_reg[124][2]/P0001 , \wishbone_bd_ram_mem0_reg[124][3]/P0001 , \wishbone_bd_ram_mem0_reg[124][4]/P0001 , \wishbone_bd_ram_mem0_reg[124][5]/P0001 , \wishbone_bd_ram_mem0_reg[124][6]/P0001 , \wishbone_bd_ram_mem0_reg[124][7]/P0001 , \wishbone_bd_ram_mem0_reg[125][0]/P0001 , \wishbone_bd_ram_mem0_reg[125][1]/P0001 , \wishbone_bd_ram_mem0_reg[125][2]/P0001 , \wishbone_bd_ram_mem0_reg[125][3]/P0001 , \wishbone_bd_ram_mem0_reg[125][4]/P0001 , \wishbone_bd_ram_mem0_reg[125][5]/P0001 , \wishbone_bd_ram_mem0_reg[125][6]/P0001 , \wishbone_bd_ram_mem0_reg[125][7]/P0001 , \wishbone_bd_ram_mem0_reg[126][0]/P0001 , \wishbone_bd_ram_mem0_reg[126][1]/P0001 , \wishbone_bd_ram_mem0_reg[126][2]/P0001 , \wishbone_bd_ram_mem0_reg[126][3]/P0001 , \wishbone_bd_ram_mem0_reg[126][4]/P0001 , \wishbone_bd_ram_mem0_reg[126][5]/P0001 , \wishbone_bd_ram_mem0_reg[126][6]/P0001 , \wishbone_bd_ram_mem0_reg[126][7]/P0001 , \wishbone_bd_ram_mem0_reg[127][0]/P0001 , \wishbone_bd_ram_mem0_reg[127][1]/P0001 , \wishbone_bd_ram_mem0_reg[127][2]/P0001 , \wishbone_bd_ram_mem0_reg[127][3]/P0001 , \wishbone_bd_ram_mem0_reg[127][4]/P0001 , \wishbone_bd_ram_mem0_reg[127][5]/P0001 , \wishbone_bd_ram_mem0_reg[127][6]/P0001 , \wishbone_bd_ram_mem0_reg[127][7]/P0001 , \wishbone_bd_ram_mem0_reg[128][0]/P0001 , \wishbone_bd_ram_mem0_reg[128][1]/P0001 , \wishbone_bd_ram_mem0_reg[128][2]/P0001 , \wishbone_bd_ram_mem0_reg[128][3]/P0001 , \wishbone_bd_ram_mem0_reg[128][4]/P0001 , \wishbone_bd_ram_mem0_reg[128][5]/P0001 , \wishbone_bd_ram_mem0_reg[128][6]/P0001 , \wishbone_bd_ram_mem0_reg[128][7]/P0001 , \wishbone_bd_ram_mem0_reg[129][0]/P0001 , \wishbone_bd_ram_mem0_reg[129][1]/P0001 , \wishbone_bd_ram_mem0_reg[129][2]/P0001 , \wishbone_bd_ram_mem0_reg[129][3]/P0001 , \wishbone_bd_ram_mem0_reg[129][4]/P0001 , \wishbone_bd_ram_mem0_reg[129][5]/P0001 , \wishbone_bd_ram_mem0_reg[129][6]/P0001 , \wishbone_bd_ram_mem0_reg[129][7]/P0001 , \wishbone_bd_ram_mem0_reg[12][0]/P0001 , \wishbone_bd_ram_mem0_reg[12][1]/P0001 , \wishbone_bd_ram_mem0_reg[12][2]/P0001 , \wishbone_bd_ram_mem0_reg[12][3]/P0001 , \wishbone_bd_ram_mem0_reg[12][4]/P0001 , \wishbone_bd_ram_mem0_reg[12][5]/P0001 , \wishbone_bd_ram_mem0_reg[12][6]/P0001 , \wishbone_bd_ram_mem0_reg[12][7]/P0001 , \wishbone_bd_ram_mem0_reg[130][0]/P0001 , \wishbone_bd_ram_mem0_reg[130][1]/P0001 , \wishbone_bd_ram_mem0_reg[130][2]/P0001 , \wishbone_bd_ram_mem0_reg[130][3]/P0001 , \wishbone_bd_ram_mem0_reg[130][4]/P0001 , \wishbone_bd_ram_mem0_reg[130][5]/P0001 , \wishbone_bd_ram_mem0_reg[130][6]/P0001 , \wishbone_bd_ram_mem0_reg[130][7]/P0001 , \wishbone_bd_ram_mem0_reg[131][0]/P0001 , \wishbone_bd_ram_mem0_reg[131][1]/P0001 , \wishbone_bd_ram_mem0_reg[131][2]/P0001 , \wishbone_bd_ram_mem0_reg[131][3]/P0001 , \wishbone_bd_ram_mem0_reg[131][4]/P0001 , \wishbone_bd_ram_mem0_reg[131][5]/P0001 , \wishbone_bd_ram_mem0_reg[131][6]/P0001 , \wishbone_bd_ram_mem0_reg[131][7]/P0001 , \wishbone_bd_ram_mem0_reg[132][0]/P0001 , \wishbone_bd_ram_mem0_reg[132][1]/P0001 , \wishbone_bd_ram_mem0_reg[132][2]/P0001 , \wishbone_bd_ram_mem0_reg[132][3]/P0001 , \wishbone_bd_ram_mem0_reg[132][4]/P0001 , \wishbone_bd_ram_mem0_reg[132][5]/P0001 , \wishbone_bd_ram_mem0_reg[132][6]/P0001 , \wishbone_bd_ram_mem0_reg[132][7]/P0001 , \wishbone_bd_ram_mem0_reg[133][0]/P0001 , \wishbone_bd_ram_mem0_reg[133][1]/P0001 , \wishbone_bd_ram_mem0_reg[133][2]/P0001 , \wishbone_bd_ram_mem0_reg[133][3]/P0001 , \wishbone_bd_ram_mem0_reg[133][4]/P0001 , \wishbone_bd_ram_mem0_reg[133][5]/P0001 , \wishbone_bd_ram_mem0_reg[133][6]/P0001 , \wishbone_bd_ram_mem0_reg[133][7]/P0001 , \wishbone_bd_ram_mem0_reg[134][0]/P0001 , \wishbone_bd_ram_mem0_reg[134][1]/P0001 , \wishbone_bd_ram_mem0_reg[134][2]/P0001 , \wishbone_bd_ram_mem0_reg[134][3]/P0001 , \wishbone_bd_ram_mem0_reg[134][4]/P0001 , \wishbone_bd_ram_mem0_reg[134][5]/P0001 , \wishbone_bd_ram_mem0_reg[134][6]/P0001 , \wishbone_bd_ram_mem0_reg[134][7]/P0001 , \wishbone_bd_ram_mem0_reg[135][0]/P0001 , \wishbone_bd_ram_mem0_reg[135][1]/P0001 , \wishbone_bd_ram_mem0_reg[135][2]/P0001 , \wishbone_bd_ram_mem0_reg[135][3]/P0001 , \wishbone_bd_ram_mem0_reg[135][4]/P0001 , \wishbone_bd_ram_mem0_reg[135][5]/P0001 , \wishbone_bd_ram_mem0_reg[135][6]/P0001 , \wishbone_bd_ram_mem0_reg[135][7]/P0001 , \wishbone_bd_ram_mem0_reg[136][0]/P0001 , \wishbone_bd_ram_mem0_reg[136][1]/P0001 , \wishbone_bd_ram_mem0_reg[136][2]/P0001 , \wishbone_bd_ram_mem0_reg[136][3]/P0001 , \wishbone_bd_ram_mem0_reg[136][4]/P0001 , \wishbone_bd_ram_mem0_reg[136][5]/P0001 , \wishbone_bd_ram_mem0_reg[136][6]/P0001 , \wishbone_bd_ram_mem0_reg[136][7]/P0001 , \wishbone_bd_ram_mem0_reg[137][0]/P0001 , \wishbone_bd_ram_mem0_reg[137][1]/P0001 , \wishbone_bd_ram_mem0_reg[137][2]/P0001 , \wishbone_bd_ram_mem0_reg[137][3]/P0001 , \wishbone_bd_ram_mem0_reg[137][4]/P0001 , \wishbone_bd_ram_mem0_reg[137][5]/P0001 , \wishbone_bd_ram_mem0_reg[137][6]/P0001 , \wishbone_bd_ram_mem0_reg[137][7]/P0001 , \wishbone_bd_ram_mem0_reg[138][0]/P0001 , \wishbone_bd_ram_mem0_reg[138][1]/P0001 , \wishbone_bd_ram_mem0_reg[138][2]/P0001 , \wishbone_bd_ram_mem0_reg[138][3]/P0001 , \wishbone_bd_ram_mem0_reg[138][4]/P0001 , \wishbone_bd_ram_mem0_reg[138][5]/P0001 , \wishbone_bd_ram_mem0_reg[138][6]/P0001 , \wishbone_bd_ram_mem0_reg[138][7]/P0001 , \wishbone_bd_ram_mem0_reg[139][0]/P0001 , \wishbone_bd_ram_mem0_reg[139][1]/P0001 , \wishbone_bd_ram_mem0_reg[139][2]/P0001 , \wishbone_bd_ram_mem0_reg[139][3]/P0001 , \wishbone_bd_ram_mem0_reg[139][4]/P0001 , \wishbone_bd_ram_mem0_reg[139][5]/P0001 , \wishbone_bd_ram_mem0_reg[139][6]/P0001 , \wishbone_bd_ram_mem0_reg[139][7]/P0001 , \wishbone_bd_ram_mem0_reg[13][0]/P0001 , \wishbone_bd_ram_mem0_reg[13][1]/P0001 , \wishbone_bd_ram_mem0_reg[13][2]/P0001 , \wishbone_bd_ram_mem0_reg[13][3]/P0001 , \wishbone_bd_ram_mem0_reg[13][4]/P0001 , \wishbone_bd_ram_mem0_reg[13][5]/P0001 , \wishbone_bd_ram_mem0_reg[13][6]/P0001 , \wishbone_bd_ram_mem0_reg[13][7]/P0001 , \wishbone_bd_ram_mem0_reg[140][0]/P0001 , \wishbone_bd_ram_mem0_reg[140][1]/P0001 , \wishbone_bd_ram_mem0_reg[140][2]/P0001 , \wishbone_bd_ram_mem0_reg[140][3]/P0001 , \wishbone_bd_ram_mem0_reg[140][4]/P0001 , \wishbone_bd_ram_mem0_reg[140][5]/P0001 , \wishbone_bd_ram_mem0_reg[140][6]/P0001 , \wishbone_bd_ram_mem0_reg[140][7]/P0001 , \wishbone_bd_ram_mem0_reg[141][0]/P0001 , \wishbone_bd_ram_mem0_reg[141][1]/P0001 , \wishbone_bd_ram_mem0_reg[141][2]/P0001 , \wishbone_bd_ram_mem0_reg[141][3]/P0001 , \wishbone_bd_ram_mem0_reg[141][4]/P0001 , \wishbone_bd_ram_mem0_reg[141][5]/P0001 , \wishbone_bd_ram_mem0_reg[141][6]/P0001 , \wishbone_bd_ram_mem0_reg[141][7]/P0001 , \wishbone_bd_ram_mem0_reg[142][0]/P0001 , \wishbone_bd_ram_mem0_reg[142][1]/P0001 , \wishbone_bd_ram_mem0_reg[142][2]/P0001 , \wishbone_bd_ram_mem0_reg[142][3]/P0001 , \wishbone_bd_ram_mem0_reg[142][4]/P0001 , \wishbone_bd_ram_mem0_reg[142][5]/P0001 , \wishbone_bd_ram_mem0_reg[142][6]/P0001 , \wishbone_bd_ram_mem0_reg[142][7]/P0001 , \wishbone_bd_ram_mem0_reg[143][0]/P0001 , \wishbone_bd_ram_mem0_reg[143][1]/P0001 , \wishbone_bd_ram_mem0_reg[143][2]/P0001 , \wishbone_bd_ram_mem0_reg[143][3]/P0001 , \wishbone_bd_ram_mem0_reg[143][4]/P0001 , \wishbone_bd_ram_mem0_reg[143][5]/P0001 , \wishbone_bd_ram_mem0_reg[143][6]/P0001 , \wishbone_bd_ram_mem0_reg[143][7]/P0001 , \wishbone_bd_ram_mem0_reg[144][0]/P0001 , \wishbone_bd_ram_mem0_reg[144][1]/P0001 , \wishbone_bd_ram_mem0_reg[144][2]/P0001 , \wishbone_bd_ram_mem0_reg[144][3]/P0001 , \wishbone_bd_ram_mem0_reg[144][4]/P0001 , \wishbone_bd_ram_mem0_reg[144][5]/P0001 , \wishbone_bd_ram_mem0_reg[144][6]/P0001 , \wishbone_bd_ram_mem0_reg[144][7]/P0001 , \wishbone_bd_ram_mem0_reg[145][0]/P0001 , \wishbone_bd_ram_mem0_reg[145][1]/P0001 , \wishbone_bd_ram_mem0_reg[145][2]/P0001 , \wishbone_bd_ram_mem0_reg[145][3]/P0001 , \wishbone_bd_ram_mem0_reg[145][4]/P0001 , \wishbone_bd_ram_mem0_reg[145][5]/P0001 , \wishbone_bd_ram_mem0_reg[145][6]/P0001 , \wishbone_bd_ram_mem0_reg[145][7]/P0001 , \wishbone_bd_ram_mem0_reg[146][0]/P0001 , \wishbone_bd_ram_mem0_reg[146][1]/P0001 , \wishbone_bd_ram_mem0_reg[146][2]/P0001 , \wishbone_bd_ram_mem0_reg[146][3]/P0001 , \wishbone_bd_ram_mem0_reg[146][4]/P0001 , \wishbone_bd_ram_mem0_reg[146][5]/P0001 , \wishbone_bd_ram_mem0_reg[146][6]/P0001 , \wishbone_bd_ram_mem0_reg[146][7]/P0001 , \wishbone_bd_ram_mem0_reg[147][0]/P0001 , \wishbone_bd_ram_mem0_reg[147][1]/P0001 , \wishbone_bd_ram_mem0_reg[147][2]/P0001 , \wishbone_bd_ram_mem0_reg[147][3]/P0001 , \wishbone_bd_ram_mem0_reg[147][4]/P0001 , \wishbone_bd_ram_mem0_reg[147][5]/P0001 , \wishbone_bd_ram_mem0_reg[147][6]/P0001 , \wishbone_bd_ram_mem0_reg[147][7]/P0001 , \wishbone_bd_ram_mem0_reg[148][0]/P0001 , \wishbone_bd_ram_mem0_reg[148][1]/P0001 , \wishbone_bd_ram_mem0_reg[148][2]/P0001 , \wishbone_bd_ram_mem0_reg[148][3]/P0001 , \wishbone_bd_ram_mem0_reg[148][4]/P0001 , \wishbone_bd_ram_mem0_reg[148][5]/P0001 , \wishbone_bd_ram_mem0_reg[148][6]/P0001 , \wishbone_bd_ram_mem0_reg[148][7]/P0001 , \wishbone_bd_ram_mem0_reg[149][0]/P0001 , \wishbone_bd_ram_mem0_reg[149][1]/P0001 , \wishbone_bd_ram_mem0_reg[149][2]/P0001 , \wishbone_bd_ram_mem0_reg[149][3]/P0001 , \wishbone_bd_ram_mem0_reg[149][4]/P0001 , \wishbone_bd_ram_mem0_reg[149][5]/P0001 , \wishbone_bd_ram_mem0_reg[149][6]/P0001 , \wishbone_bd_ram_mem0_reg[149][7]/P0001 , \wishbone_bd_ram_mem0_reg[14][0]/P0001 , \wishbone_bd_ram_mem0_reg[14][1]/P0001 , \wishbone_bd_ram_mem0_reg[14][2]/P0001 , \wishbone_bd_ram_mem0_reg[14][3]/P0001 , \wishbone_bd_ram_mem0_reg[14][4]/P0001 , \wishbone_bd_ram_mem0_reg[14][5]/P0001 , \wishbone_bd_ram_mem0_reg[14][6]/P0001 , \wishbone_bd_ram_mem0_reg[14][7]/P0001 , \wishbone_bd_ram_mem0_reg[150][0]/P0001 , \wishbone_bd_ram_mem0_reg[150][1]/P0001 , \wishbone_bd_ram_mem0_reg[150][2]/P0001 , \wishbone_bd_ram_mem0_reg[150][3]/P0001 , \wishbone_bd_ram_mem0_reg[150][4]/P0001 , \wishbone_bd_ram_mem0_reg[150][5]/P0001 , \wishbone_bd_ram_mem0_reg[150][6]/P0001 , \wishbone_bd_ram_mem0_reg[150][7]/P0001 , \wishbone_bd_ram_mem0_reg[151][0]/P0001 , \wishbone_bd_ram_mem0_reg[151][1]/P0001 , \wishbone_bd_ram_mem0_reg[151][2]/P0001 , \wishbone_bd_ram_mem0_reg[151][3]/P0001 , \wishbone_bd_ram_mem0_reg[151][4]/P0001 , \wishbone_bd_ram_mem0_reg[151][5]/P0001 , \wishbone_bd_ram_mem0_reg[151][6]/P0001 , \wishbone_bd_ram_mem0_reg[151][7]/P0001 , \wishbone_bd_ram_mem0_reg[152][0]/P0001 , \wishbone_bd_ram_mem0_reg[152][1]/P0001 , \wishbone_bd_ram_mem0_reg[152][2]/P0001 , \wishbone_bd_ram_mem0_reg[152][3]/P0001 , \wishbone_bd_ram_mem0_reg[152][4]/P0001 , \wishbone_bd_ram_mem0_reg[152][5]/P0001 , \wishbone_bd_ram_mem0_reg[152][6]/P0001 , \wishbone_bd_ram_mem0_reg[152][7]/P0001 , \wishbone_bd_ram_mem0_reg[153][0]/P0001 , \wishbone_bd_ram_mem0_reg[153][1]/P0001 , \wishbone_bd_ram_mem0_reg[153][2]/P0001 , \wishbone_bd_ram_mem0_reg[153][3]/P0001 , \wishbone_bd_ram_mem0_reg[153][4]/P0001 , \wishbone_bd_ram_mem0_reg[153][5]/P0001 , \wishbone_bd_ram_mem0_reg[153][6]/P0001 , \wishbone_bd_ram_mem0_reg[153][7]/P0001 , \wishbone_bd_ram_mem0_reg[154][0]/P0001 , \wishbone_bd_ram_mem0_reg[154][1]/P0001 , \wishbone_bd_ram_mem0_reg[154][2]/P0001 , \wishbone_bd_ram_mem0_reg[154][3]/P0001 , \wishbone_bd_ram_mem0_reg[154][4]/P0001 , \wishbone_bd_ram_mem0_reg[154][5]/P0001 , \wishbone_bd_ram_mem0_reg[154][6]/P0001 , \wishbone_bd_ram_mem0_reg[154][7]/P0001 , \wishbone_bd_ram_mem0_reg[155][0]/P0001 , \wishbone_bd_ram_mem0_reg[155][1]/P0001 , \wishbone_bd_ram_mem0_reg[155][2]/P0001 , \wishbone_bd_ram_mem0_reg[155][3]/P0001 , \wishbone_bd_ram_mem0_reg[155][4]/P0001 , \wishbone_bd_ram_mem0_reg[155][5]/P0001 , \wishbone_bd_ram_mem0_reg[155][6]/P0001 , \wishbone_bd_ram_mem0_reg[155][7]/P0001 , \wishbone_bd_ram_mem0_reg[156][0]/P0001 , \wishbone_bd_ram_mem0_reg[156][1]/P0001 , \wishbone_bd_ram_mem0_reg[156][2]/P0001 , \wishbone_bd_ram_mem0_reg[156][3]/P0001 , \wishbone_bd_ram_mem0_reg[156][4]/P0001 , \wishbone_bd_ram_mem0_reg[156][5]/P0001 , \wishbone_bd_ram_mem0_reg[156][6]/P0001 , \wishbone_bd_ram_mem0_reg[156][7]/P0001 , \wishbone_bd_ram_mem0_reg[157][0]/P0001 , \wishbone_bd_ram_mem0_reg[157][1]/P0001 , \wishbone_bd_ram_mem0_reg[157][2]/P0001 , \wishbone_bd_ram_mem0_reg[157][3]/P0001 , \wishbone_bd_ram_mem0_reg[157][4]/P0001 , \wishbone_bd_ram_mem0_reg[157][5]/P0001 , \wishbone_bd_ram_mem0_reg[157][6]/P0001 , \wishbone_bd_ram_mem0_reg[157][7]/P0001 , \wishbone_bd_ram_mem0_reg[158][0]/P0001 , \wishbone_bd_ram_mem0_reg[158][1]/P0001 , \wishbone_bd_ram_mem0_reg[158][2]/P0001 , \wishbone_bd_ram_mem0_reg[158][3]/P0001 , \wishbone_bd_ram_mem0_reg[158][4]/P0001 , \wishbone_bd_ram_mem0_reg[158][5]/P0001 , \wishbone_bd_ram_mem0_reg[158][6]/P0001 , \wishbone_bd_ram_mem0_reg[158][7]/P0001 , \wishbone_bd_ram_mem0_reg[159][0]/P0001 , \wishbone_bd_ram_mem0_reg[159][1]/P0001 , \wishbone_bd_ram_mem0_reg[159][2]/P0001 , \wishbone_bd_ram_mem0_reg[159][3]/P0001 , \wishbone_bd_ram_mem0_reg[159][4]/P0001 , \wishbone_bd_ram_mem0_reg[159][5]/P0001 , \wishbone_bd_ram_mem0_reg[159][6]/P0001 , \wishbone_bd_ram_mem0_reg[159][7]/P0001 , \wishbone_bd_ram_mem0_reg[15][0]/P0001 , \wishbone_bd_ram_mem0_reg[15][1]/P0001 , \wishbone_bd_ram_mem0_reg[15][2]/P0001 , \wishbone_bd_ram_mem0_reg[15][3]/P0001 , \wishbone_bd_ram_mem0_reg[15][4]/P0001 , \wishbone_bd_ram_mem0_reg[15][5]/P0001 , \wishbone_bd_ram_mem0_reg[15][6]/P0001 , \wishbone_bd_ram_mem0_reg[15][7]/P0001 , \wishbone_bd_ram_mem0_reg[160][0]/P0001 , \wishbone_bd_ram_mem0_reg[160][1]/P0001 , \wishbone_bd_ram_mem0_reg[160][2]/P0001 , \wishbone_bd_ram_mem0_reg[160][3]/P0001 , \wishbone_bd_ram_mem0_reg[160][4]/P0001 , \wishbone_bd_ram_mem0_reg[160][5]/P0001 , \wishbone_bd_ram_mem0_reg[160][6]/P0001 , \wishbone_bd_ram_mem0_reg[160][7]/P0001 , \wishbone_bd_ram_mem0_reg[161][0]/P0001 , \wishbone_bd_ram_mem0_reg[161][1]/P0001 , \wishbone_bd_ram_mem0_reg[161][2]/P0001 , \wishbone_bd_ram_mem0_reg[161][3]/P0001 , \wishbone_bd_ram_mem0_reg[161][4]/P0001 , \wishbone_bd_ram_mem0_reg[161][5]/P0001 , \wishbone_bd_ram_mem0_reg[161][6]/P0001 , \wishbone_bd_ram_mem0_reg[161][7]/P0001 , \wishbone_bd_ram_mem0_reg[162][0]/P0001 , \wishbone_bd_ram_mem0_reg[162][1]/P0001 , \wishbone_bd_ram_mem0_reg[162][2]/P0001 , \wishbone_bd_ram_mem0_reg[162][3]/P0001 , \wishbone_bd_ram_mem0_reg[162][4]/P0001 , \wishbone_bd_ram_mem0_reg[162][5]/P0001 , \wishbone_bd_ram_mem0_reg[162][6]/P0001 , \wishbone_bd_ram_mem0_reg[162][7]/P0001 , \wishbone_bd_ram_mem0_reg[163][0]/P0001 , \wishbone_bd_ram_mem0_reg[163][1]/P0001 , \wishbone_bd_ram_mem0_reg[163][2]/P0001 , \wishbone_bd_ram_mem0_reg[163][3]/P0001 , \wishbone_bd_ram_mem0_reg[163][4]/P0001 , \wishbone_bd_ram_mem0_reg[163][5]/P0001 , \wishbone_bd_ram_mem0_reg[163][6]/P0001 , \wishbone_bd_ram_mem0_reg[163][7]/P0001 , \wishbone_bd_ram_mem0_reg[164][0]/P0001 , \wishbone_bd_ram_mem0_reg[164][1]/P0001 , \wishbone_bd_ram_mem0_reg[164][2]/P0001 , \wishbone_bd_ram_mem0_reg[164][3]/P0001 , \wishbone_bd_ram_mem0_reg[164][4]/P0001 , \wishbone_bd_ram_mem0_reg[164][5]/P0001 , \wishbone_bd_ram_mem0_reg[164][6]/P0001 , \wishbone_bd_ram_mem0_reg[164][7]/P0001 , \wishbone_bd_ram_mem0_reg[165][0]/P0001 , \wishbone_bd_ram_mem0_reg[165][1]/P0001 , \wishbone_bd_ram_mem0_reg[165][2]/P0001 , \wishbone_bd_ram_mem0_reg[165][3]/P0001 , \wishbone_bd_ram_mem0_reg[165][4]/P0001 , \wishbone_bd_ram_mem0_reg[165][5]/P0001 , \wishbone_bd_ram_mem0_reg[165][6]/P0001 , \wishbone_bd_ram_mem0_reg[165][7]/P0001 , \wishbone_bd_ram_mem0_reg[166][0]/P0001 , \wishbone_bd_ram_mem0_reg[166][1]/P0001 , \wishbone_bd_ram_mem0_reg[166][2]/P0001 , \wishbone_bd_ram_mem0_reg[166][3]/P0001 , \wishbone_bd_ram_mem0_reg[166][4]/P0001 , \wishbone_bd_ram_mem0_reg[166][5]/P0001 , \wishbone_bd_ram_mem0_reg[166][6]/P0001 , \wishbone_bd_ram_mem0_reg[166][7]/P0001 , \wishbone_bd_ram_mem0_reg[167][0]/P0001 , \wishbone_bd_ram_mem0_reg[167][1]/P0001 , \wishbone_bd_ram_mem0_reg[167][2]/P0001 , \wishbone_bd_ram_mem0_reg[167][3]/P0001 , \wishbone_bd_ram_mem0_reg[167][4]/P0001 , \wishbone_bd_ram_mem0_reg[167][5]/P0001 , \wishbone_bd_ram_mem0_reg[167][6]/P0001 , \wishbone_bd_ram_mem0_reg[167][7]/P0001 , \wishbone_bd_ram_mem0_reg[168][0]/P0001 , \wishbone_bd_ram_mem0_reg[168][1]/P0001 , \wishbone_bd_ram_mem0_reg[168][2]/P0001 , \wishbone_bd_ram_mem0_reg[168][3]/P0001 , \wishbone_bd_ram_mem0_reg[168][4]/P0001 , \wishbone_bd_ram_mem0_reg[168][5]/P0001 , \wishbone_bd_ram_mem0_reg[168][6]/P0001 , \wishbone_bd_ram_mem0_reg[168][7]/P0001 , \wishbone_bd_ram_mem0_reg[169][0]/P0001 , \wishbone_bd_ram_mem0_reg[169][1]/P0001 , \wishbone_bd_ram_mem0_reg[169][2]/P0001 , \wishbone_bd_ram_mem0_reg[169][3]/P0001 , \wishbone_bd_ram_mem0_reg[169][4]/P0001 , \wishbone_bd_ram_mem0_reg[169][5]/P0001 , \wishbone_bd_ram_mem0_reg[169][6]/P0001 , \wishbone_bd_ram_mem0_reg[169][7]/P0001 , \wishbone_bd_ram_mem0_reg[16][0]/P0001 , \wishbone_bd_ram_mem0_reg[16][1]/P0001 , \wishbone_bd_ram_mem0_reg[16][2]/P0001 , \wishbone_bd_ram_mem0_reg[16][3]/P0001 , \wishbone_bd_ram_mem0_reg[16][4]/P0001 , \wishbone_bd_ram_mem0_reg[16][5]/P0001 , \wishbone_bd_ram_mem0_reg[16][6]/P0001 , \wishbone_bd_ram_mem0_reg[16][7]/P0001 , \wishbone_bd_ram_mem0_reg[170][0]/P0001 , \wishbone_bd_ram_mem0_reg[170][1]/P0001 , \wishbone_bd_ram_mem0_reg[170][2]/P0001 , \wishbone_bd_ram_mem0_reg[170][3]/P0001 , \wishbone_bd_ram_mem0_reg[170][4]/P0001 , \wishbone_bd_ram_mem0_reg[170][5]/P0001 , \wishbone_bd_ram_mem0_reg[170][6]/P0001 , \wishbone_bd_ram_mem0_reg[170][7]/P0001 , \wishbone_bd_ram_mem0_reg[171][0]/P0001 , \wishbone_bd_ram_mem0_reg[171][1]/P0001 , \wishbone_bd_ram_mem0_reg[171][2]/P0001 , \wishbone_bd_ram_mem0_reg[171][3]/P0001 , \wishbone_bd_ram_mem0_reg[171][4]/P0001 , \wishbone_bd_ram_mem0_reg[171][5]/P0001 , \wishbone_bd_ram_mem0_reg[171][6]/P0001 , \wishbone_bd_ram_mem0_reg[171][7]/P0001 , \wishbone_bd_ram_mem0_reg[172][0]/P0001 , \wishbone_bd_ram_mem0_reg[172][1]/P0001 , \wishbone_bd_ram_mem0_reg[172][2]/P0001 , \wishbone_bd_ram_mem0_reg[172][3]/P0001 , \wishbone_bd_ram_mem0_reg[172][4]/P0001 , \wishbone_bd_ram_mem0_reg[172][5]/P0001 , \wishbone_bd_ram_mem0_reg[172][6]/P0001 , \wishbone_bd_ram_mem0_reg[172][7]/P0001 , \wishbone_bd_ram_mem0_reg[173][0]/P0001 , \wishbone_bd_ram_mem0_reg[173][1]/P0001 , \wishbone_bd_ram_mem0_reg[173][2]/P0001 , \wishbone_bd_ram_mem0_reg[173][3]/P0001 , \wishbone_bd_ram_mem0_reg[173][4]/P0001 , \wishbone_bd_ram_mem0_reg[173][5]/P0001 , \wishbone_bd_ram_mem0_reg[173][6]/P0001 , \wishbone_bd_ram_mem0_reg[173][7]/P0001 , \wishbone_bd_ram_mem0_reg[174][0]/P0001 , \wishbone_bd_ram_mem0_reg[174][1]/P0001 , \wishbone_bd_ram_mem0_reg[174][2]/P0001 , \wishbone_bd_ram_mem0_reg[174][3]/P0001 , \wishbone_bd_ram_mem0_reg[174][4]/P0001 , \wishbone_bd_ram_mem0_reg[174][5]/P0001 , \wishbone_bd_ram_mem0_reg[174][6]/P0001 , \wishbone_bd_ram_mem0_reg[174][7]/P0001 , \wishbone_bd_ram_mem0_reg[175][0]/P0001 , \wishbone_bd_ram_mem0_reg[175][1]/P0001 , \wishbone_bd_ram_mem0_reg[175][2]/P0001 , \wishbone_bd_ram_mem0_reg[175][3]/P0001 , \wishbone_bd_ram_mem0_reg[175][4]/P0001 , \wishbone_bd_ram_mem0_reg[175][5]/P0001 , \wishbone_bd_ram_mem0_reg[175][6]/P0001 , \wishbone_bd_ram_mem0_reg[175][7]/P0001 , \wishbone_bd_ram_mem0_reg[176][0]/P0001 , \wishbone_bd_ram_mem0_reg[176][1]/P0001 , \wishbone_bd_ram_mem0_reg[176][2]/P0001 , \wishbone_bd_ram_mem0_reg[176][3]/P0001 , \wishbone_bd_ram_mem0_reg[176][4]/P0001 , \wishbone_bd_ram_mem0_reg[176][5]/P0001 , \wishbone_bd_ram_mem0_reg[176][6]/P0001 , \wishbone_bd_ram_mem0_reg[176][7]/P0001 , \wishbone_bd_ram_mem0_reg[177][0]/P0001 , \wishbone_bd_ram_mem0_reg[177][1]/P0001 , \wishbone_bd_ram_mem0_reg[177][2]/P0001 , \wishbone_bd_ram_mem0_reg[177][3]/P0001 , \wishbone_bd_ram_mem0_reg[177][4]/P0001 , \wishbone_bd_ram_mem0_reg[177][5]/P0001 , \wishbone_bd_ram_mem0_reg[177][6]/P0001 , \wishbone_bd_ram_mem0_reg[177][7]/P0001 , \wishbone_bd_ram_mem0_reg[178][0]/P0001 , \wishbone_bd_ram_mem0_reg[178][1]/P0001 , \wishbone_bd_ram_mem0_reg[178][2]/P0001 , \wishbone_bd_ram_mem0_reg[178][3]/P0001 , \wishbone_bd_ram_mem0_reg[178][4]/P0001 , \wishbone_bd_ram_mem0_reg[178][5]/P0001 , \wishbone_bd_ram_mem0_reg[178][6]/P0001 , \wishbone_bd_ram_mem0_reg[178][7]/P0001 , \wishbone_bd_ram_mem0_reg[179][0]/P0001 , \wishbone_bd_ram_mem0_reg[179][1]/P0001 , \wishbone_bd_ram_mem0_reg[179][2]/P0001 , \wishbone_bd_ram_mem0_reg[179][3]/P0001 , \wishbone_bd_ram_mem0_reg[179][4]/P0001 , \wishbone_bd_ram_mem0_reg[179][5]/P0001 , \wishbone_bd_ram_mem0_reg[179][6]/P0001 , \wishbone_bd_ram_mem0_reg[179][7]/P0001 , \wishbone_bd_ram_mem0_reg[17][0]/P0001 , \wishbone_bd_ram_mem0_reg[17][1]/P0001 , \wishbone_bd_ram_mem0_reg[17][2]/P0001 , \wishbone_bd_ram_mem0_reg[17][3]/P0001 , \wishbone_bd_ram_mem0_reg[17][4]/P0001 , \wishbone_bd_ram_mem0_reg[17][5]/P0001 , \wishbone_bd_ram_mem0_reg[17][6]/P0001 , \wishbone_bd_ram_mem0_reg[17][7]/P0001 , \wishbone_bd_ram_mem0_reg[180][0]/P0001 , \wishbone_bd_ram_mem0_reg[180][1]/P0001 , \wishbone_bd_ram_mem0_reg[180][2]/P0001 , \wishbone_bd_ram_mem0_reg[180][3]/P0001 , \wishbone_bd_ram_mem0_reg[180][4]/P0001 , \wishbone_bd_ram_mem0_reg[180][5]/P0001 , \wishbone_bd_ram_mem0_reg[180][6]/P0001 , \wishbone_bd_ram_mem0_reg[180][7]/P0001 , \wishbone_bd_ram_mem0_reg[181][0]/P0001 , \wishbone_bd_ram_mem0_reg[181][1]/P0001 , \wishbone_bd_ram_mem0_reg[181][2]/P0001 , \wishbone_bd_ram_mem0_reg[181][3]/P0001 , \wishbone_bd_ram_mem0_reg[181][4]/P0001 , \wishbone_bd_ram_mem0_reg[181][5]/P0001 , \wishbone_bd_ram_mem0_reg[181][6]/P0001 , \wishbone_bd_ram_mem0_reg[181][7]/P0001 , \wishbone_bd_ram_mem0_reg[182][0]/P0001 , \wishbone_bd_ram_mem0_reg[182][1]/P0001 , \wishbone_bd_ram_mem0_reg[182][2]/P0001 , \wishbone_bd_ram_mem0_reg[182][3]/P0001 , \wishbone_bd_ram_mem0_reg[182][4]/P0001 , \wishbone_bd_ram_mem0_reg[182][5]/P0001 , \wishbone_bd_ram_mem0_reg[182][6]/P0001 , \wishbone_bd_ram_mem0_reg[182][7]/P0001 , \wishbone_bd_ram_mem0_reg[183][0]/P0001 , \wishbone_bd_ram_mem0_reg[183][1]/P0001 , \wishbone_bd_ram_mem0_reg[183][2]/P0001 , \wishbone_bd_ram_mem0_reg[183][3]/P0001 , \wishbone_bd_ram_mem0_reg[183][4]/P0001 , \wishbone_bd_ram_mem0_reg[183][5]/P0001 , \wishbone_bd_ram_mem0_reg[183][6]/P0001 , \wishbone_bd_ram_mem0_reg[183][7]/P0001 , \wishbone_bd_ram_mem0_reg[184][0]/P0001 , \wishbone_bd_ram_mem0_reg[184][1]/P0001 , \wishbone_bd_ram_mem0_reg[184][2]/P0001 , \wishbone_bd_ram_mem0_reg[184][3]/P0001 , \wishbone_bd_ram_mem0_reg[184][4]/P0001 , \wishbone_bd_ram_mem0_reg[184][5]/P0001 , \wishbone_bd_ram_mem0_reg[184][6]/P0001 , \wishbone_bd_ram_mem0_reg[184][7]/P0001 , \wishbone_bd_ram_mem0_reg[185][0]/P0001 , \wishbone_bd_ram_mem0_reg[185][1]/P0001 , \wishbone_bd_ram_mem0_reg[185][2]/P0001 , \wishbone_bd_ram_mem0_reg[185][3]/P0001 , \wishbone_bd_ram_mem0_reg[185][4]/P0001 , \wishbone_bd_ram_mem0_reg[185][5]/P0001 , \wishbone_bd_ram_mem0_reg[185][6]/P0001 , \wishbone_bd_ram_mem0_reg[185][7]/P0001 , \wishbone_bd_ram_mem0_reg[186][0]/P0001 , \wishbone_bd_ram_mem0_reg[186][1]/P0001 , \wishbone_bd_ram_mem0_reg[186][2]/P0001 , \wishbone_bd_ram_mem0_reg[186][3]/P0001 , \wishbone_bd_ram_mem0_reg[186][4]/P0001 , \wishbone_bd_ram_mem0_reg[186][5]/P0001 , \wishbone_bd_ram_mem0_reg[186][6]/P0001 , \wishbone_bd_ram_mem0_reg[186][7]/P0001 , \wishbone_bd_ram_mem0_reg[187][0]/P0001 , \wishbone_bd_ram_mem0_reg[187][1]/P0001 , \wishbone_bd_ram_mem0_reg[187][2]/P0001 , \wishbone_bd_ram_mem0_reg[187][3]/P0001 , \wishbone_bd_ram_mem0_reg[187][4]/P0001 , \wishbone_bd_ram_mem0_reg[187][5]/P0001 , \wishbone_bd_ram_mem0_reg[187][6]/P0001 , \wishbone_bd_ram_mem0_reg[187][7]/P0001 , \wishbone_bd_ram_mem0_reg[188][0]/P0001 , \wishbone_bd_ram_mem0_reg[188][1]/P0001 , \wishbone_bd_ram_mem0_reg[188][2]/P0001 , \wishbone_bd_ram_mem0_reg[188][3]/P0001 , \wishbone_bd_ram_mem0_reg[188][4]/P0001 , \wishbone_bd_ram_mem0_reg[188][5]/P0001 , \wishbone_bd_ram_mem0_reg[188][6]/P0001 , \wishbone_bd_ram_mem0_reg[188][7]/P0001 , \wishbone_bd_ram_mem0_reg[189][0]/P0001 , \wishbone_bd_ram_mem0_reg[189][1]/P0001 , \wishbone_bd_ram_mem0_reg[189][2]/P0001 , \wishbone_bd_ram_mem0_reg[189][3]/P0001 , \wishbone_bd_ram_mem0_reg[189][4]/P0001 , \wishbone_bd_ram_mem0_reg[189][5]/P0001 , \wishbone_bd_ram_mem0_reg[189][6]/P0001 , \wishbone_bd_ram_mem0_reg[189][7]/P0001 , \wishbone_bd_ram_mem0_reg[18][0]/P0001 , \wishbone_bd_ram_mem0_reg[18][1]/P0001 , \wishbone_bd_ram_mem0_reg[18][2]/P0001 , \wishbone_bd_ram_mem0_reg[18][3]/P0001 , \wishbone_bd_ram_mem0_reg[18][4]/P0001 , \wishbone_bd_ram_mem0_reg[18][5]/P0001 , \wishbone_bd_ram_mem0_reg[18][6]/P0001 , \wishbone_bd_ram_mem0_reg[18][7]/P0001 , \wishbone_bd_ram_mem0_reg[190][0]/P0001 , \wishbone_bd_ram_mem0_reg[190][1]/P0001 , \wishbone_bd_ram_mem0_reg[190][2]/P0001 , \wishbone_bd_ram_mem0_reg[190][3]/P0001 , \wishbone_bd_ram_mem0_reg[190][4]/P0001 , \wishbone_bd_ram_mem0_reg[190][5]/P0001 , \wishbone_bd_ram_mem0_reg[190][6]/P0001 , \wishbone_bd_ram_mem0_reg[190][7]/P0001 , \wishbone_bd_ram_mem0_reg[191][0]/P0001 , \wishbone_bd_ram_mem0_reg[191][1]/P0001 , \wishbone_bd_ram_mem0_reg[191][2]/P0001 , \wishbone_bd_ram_mem0_reg[191][3]/P0001 , \wishbone_bd_ram_mem0_reg[191][4]/P0001 , \wishbone_bd_ram_mem0_reg[191][5]/P0001 , \wishbone_bd_ram_mem0_reg[191][6]/P0001 , \wishbone_bd_ram_mem0_reg[191][7]/P0001 , \wishbone_bd_ram_mem0_reg[192][0]/P0001 , \wishbone_bd_ram_mem0_reg[192][1]/P0001 , \wishbone_bd_ram_mem0_reg[192][2]/P0001 , \wishbone_bd_ram_mem0_reg[192][3]/P0001 , \wishbone_bd_ram_mem0_reg[192][4]/P0001 , \wishbone_bd_ram_mem0_reg[192][5]/P0001 , \wishbone_bd_ram_mem0_reg[192][6]/P0001 , \wishbone_bd_ram_mem0_reg[192][7]/P0001 , \wishbone_bd_ram_mem0_reg[193][0]/P0001 , \wishbone_bd_ram_mem0_reg[193][1]/P0001 , \wishbone_bd_ram_mem0_reg[193][2]/P0001 , \wishbone_bd_ram_mem0_reg[193][3]/P0001 , \wishbone_bd_ram_mem0_reg[193][4]/P0001 , \wishbone_bd_ram_mem0_reg[193][5]/P0001 , \wishbone_bd_ram_mem0_reg[193][6]/P0001 , \wishbone_bd_ram_mem0_reg[193][7]/P0001 , \wishbone_bd_ram_mem0_reg[194][0]/P0001 , \wishbone_bd_ram_mem0_reg[194][1]/P0001 , \wishbone_bd_ram_mem0_reg[194][2]/P0001 , \wishbone_bd_ram_mem0_reg[194][3]/P0001 , \wishbone_bd_ram_mem0_reg[194][4]/P0001 , \wishbone_bd_ram_mem0_reg[194][5]/P0001 , \wishbone_bd_ram_mem0_reg[194][6]/P0001 , \wishbone_bd_ram_mem0_reg[194][7]/P0001 , \wishbone_bd_ram_mem0_reg[195][0]/P0001 , \wishbone_bd_ram_mem0_reg[195][1]/P0001 , \wishbone_bd_ram_mem0_reg[195][2]/P0001 , \wishbone_bd_ram_mem0_reg[195][3]/P0001 , \wishbone_bd_ram_mem0_reg[195][4]/P0001 , \wishbone_bd_ram_mem0_reg[195][5]/P0001 , \wishbone_bd_ram_mem0_reg[195][6]/P0001 , \wishbone_bd_ram_mem0_reg[195][7]/P0001 , \wishbone_bd_ram_mem0_reg[196][0]/P0001 , \wishbone_bd_ram_mem0_reg[196][1]/P0001 , \wishbone_bd_ram_mem0_reg[196][2]/P0001 , \wishbone_bd_ram_mem0_reg[196][3]/P0001 , \wishbone_bd_ram_mem0_reg[196][4]/P0001 , \wishbone_bd_ram_mem0_reg[196][5]/P0001 , \wishbone_bd_ram_mem0_reg[196][6]/P0001 , \wishbone_bd_ram_mem0_reg[196][7]/P0001 , \wishbone_bd_ram_mem0_reg[197][0]/P0001 , \wishbone_bd_ram_mem0_reg[197][1]/P0001 , \wishbone_bd_ram_mem0_reg[197][2]/P0001 , \wishbone_bd_ram_mem0_reg[197][3]/P0001 , \wishbone_bd_ram_mem0_reg[197][4]/P0001 , \wishbone_bd_ram_mem0_reg[197][5]/P0001 , \wishbone_bd_ram_mem0_reg[197][6]/P0001 , \wishbone_bd_ram_mem0_reg[197][7]/P0001 , \wishbone_bd_ram_mem0_reg[198][0]/P0001 , \wishbone_bd_ram_mem0_reg[198][1]/P0001 , \wishbone_bd_ram_mem0_reg[198][2]/P0001 , \wishbone_bd_ram_mem0_reg[198][3]/P0001 , \wishbone_bd_ram_mem0_reg[198][4]/P0001 , \wishbone_bd_ram_mem0_reg[198][5]/P0001 , \wishbone_bd_ram_mem0_reg[198][6]/P0001 , \wishbone_bd_ram_mem0_reg[198][7]/P0001 , \wishbone_bd_ram_mem0_reg[199][0]/P0001 , \wishbone_bd_ram_mem0_reg[199][1]/P0001 , \wishbone_bd_ram_mem0_reg[199][2]/P0001 , \wishbone_bd_ram_mem0_reg[199][3]/P0001 , \wishbone_bd_ram_mem0_reg[199][4]/P0001 , \wishbone_bd_ram_mem0_reg[199][5]/P0001 , \wishbone_bd_ram_mem0_reg[199][6]/P0001 , \wishbone_bd_ram_mem0_reg[199][7]/P0001 , \wishbone_bd_ram_mem0_reg[19][0]/P0001 , \wishbone_bd_ram_mem0_reg[19][1]/P0001 , \wishbone_bd_ram_mem0_reg[19][2]/P0001 , \wishbone_bd_ram_mem0_reg[19][3]/P0001 , \wishbone_bd_ram_mem0_reg[19][4]/P0001 , \wishbone_bd_ram_mem0_reg[19][5]/P0001 , \wishbone_bd_ram_mem0_reg[19][6]/P0001 , \wishbone_bd_ram_mem0_reg[19][7]/P0001 , \wishbone_bd_ram_mem0_reg[1][0]/P0001 , \wishbone_bd_ram_mem0_reg[1][1]/P0001 , \wishbone_bd_ram_mem0_reg[1][2]/P0001 , \wishbone_bd_ram_mem0_reg[1][3]/P0001 , \wishbone_bd_ram_mem0_reg[1][4]/P0001 , \wishbone_bd_ram_mem0_reg[1][5]/P0001 , \wishbone_bd_ram_mem0_reg[1][6]/P0001 , \wishbone_bd_ram_mem0_reg[1][7]/P0001 , \wishbone_bd_ram_mem0_reg[200][0]/P0001 , \wishbone_bd_ram_mem0_reg[200][1]/P0001 , \wishbone_bd_ram_mem0_reg[200][2]/P0001 , \wishbone_bd_ram_mem0_reg[200][3]/P0001 , \wishbone_bd_ram_mem0_reg[200][4]/P0001 , \wishbone_bd_ram_mem0_reg[200][5]/P0001 , \wishbone_bd_ram_mem0_reg[200][6]/P0001 , \wishbone_bd_ram_mem0_reg[200][7]/P0001 , \wishbone_bd_ram_mem0_reg[201][0]/P0001 , \wishbone_bd_ram_mem0_reg[201][1]/P0001 , \wishbone_bd_ram_mem0_reg[201][2]/P0001 , \wishbone_bd_ram_mem0_reg[201][3]/P0001 , \wishbone_bd_ram_mem0_reg[201][4]/P0001 , \wishbone_bd_ram_mem0_reg[201][5]/P0001 , \wishbone_bd_ram_mem0_reg[201][6]/P0001 , \wishbone_bd_ram_mem0_reg[201][7]/P0001 , \wishbone_bd_ram_mem0_reg[202][0]/P0001 , \wishbone_bd_ram_mem0_reg[202][1]/P0001 , \wishbone_bd_ram_mem0_reg[202][2]/P0001 , \wishbone_bd_ram_mem0_reg[202][3]/P0001 , \wishbone_bd_ram_mem0_reg[202][4]/P0001 , \wishbone_bd_ram_mem0_reg[202][5]/P0001 , \wishbone_bd_ram_mem0_reg[202][6]/P0001 , \wishbone_bd_ram_mem0_reg[202][7]/P0001 , \wishbone_bd_ram_mem0_reg[203][0]/P0001 , \wishbone_bd_ram_mem0_reg[203][1]/P0001 , \wishbone_bd_ram_mem0_reg[203][2]/P0001 , \wishbone_bd_ram_mem0_reg[203][3]/P0001 , \wishbone_bd_ram_mem0_reg[203][4]/P0001 , \wishbone_bd_ram_mem0_reg[203][5]/P0001 , \wishbone_bd_ram_mem0_reg[203][6]/P0001 , \wishbone_bd_ram_mem0_reg[203][7]/P0001 , \wishbone_bd_ram_mem0_reg[204][0]/P0001 , \wishbone_bd_ram_mem0_reg[204][1]/P0001 , \wishbone_bd_ram_mem0_reg[204][2]/P0001 , \wishbone_bd_ram_mem0_reg[204][3]/P0001 , \wishbone_bd_ram_mem0_reg[204][4]/P0001 , \wishbone_bd_ram_mem0_reg[204][5]/P0001 , \wishbone_bd_ram_mem0_reg[204][6]/P0001 , \wishbone_bd_ram_mem0_reg[204][7]/P0001 , \wishbone_bd_ram_mem0_reg[205][0]/P0001 , \wishbone_bd_ram_mem0_reg[205][1]/P0001 , \wishbone_bd_ram_mem0_reg[205][2]/P0001 , \wishbone_bd_ram_mem0_reg[205][3]/P0001 , \wishbone_bd_ram_mem0_reg[205][4]/P0001 , \wishbone_bd_ram_mem0_reg[205][5]/P0001 , \wishbone_bd_ram_mem0_reg[205][6]/P0001 , \wishbone_bd_ram_mem0_reg[205][7]/P0001 , \wishbone_bd_ram_mem0_reg[206][0]/P0001 , \wishbone_bd_ram_mem0_reg[206][1]/P0001 , \wishbone_bd_ram_mem0_reg[206][2]/P0001 , \wishbone_bd_ram_mem0_reg[206][3]/P0001 , \wishbone_bd_ram_mem0_reg[206][4]/P0001 , \wishbone_bd_ram_mem0_reg[206][5]/P0001 , \wishbone_bd_ram_mem0_reg[206][6]/P0001 , \wishbone_bd_ram_mem0_reg[206][7]/P0001 , \wishbone_bd_ram_mem0_reg[207][0]/P0001 , \wishbone_bd_ram_mem0_reg[207][1]/P0001 , \wishbone_bd_ram_mem0_reg[207][2]/P0001 , \wishbone_bd_ram_mem0_reg[207][3]/P0001 , \wishbone_bd_ram_mem0_reg[207][4]/P0001 , \wishbone_bd_ram_mem0_reg[207][5]/P0001 , \wishbone_bd_ram_mem0_reg[207][6]/P0001 , \wishbone_bd_ram_mem0_reg[207][7]/P0001 , \wishbone_bd_ram_mem0_reg[208][0]/P0001 , \wishbone_bd_ram_mem0_reg[208][1]/P0001 , \wishbone_bd_ram_mem0_reg[208][2]/P0001 , \wishbone_bd_ram_mem0_reg[208][3]/P0001 , \wishbone_bd_ram_mem0_reg[208][4]/P0001 , \wishbone_bd_ram_mem0_reg[208][5]/P0001 , \wishbone_bd_ram_mem0_reg[208][6]/P0001 , \wishbone_bd_ram_mem0_reg[208][7]/P0001 , \wishbone_bd_ram_mem0_reg[209][0]/P0001 , \wishbone_bd_ram_mem0_reg[209][1]/P0001 , \wishbone_bd_ram_mem0_reg[209][2]/P0001 , \wishbone_bd_ram_mem0_reg[209][3]/P0001 , \wishbone_bd_ram_mem0_reg[209][4]/P0001 , \wishbone_bd_ram_mem0_reg[209][5]/P0001 , \wishbone_bd_ram_mem0_reg[209][6]/P0001 , \wishbone_bd_ram_mem0_reg[209][7]/P0001 , \wishbone_bd_ram_mem0_reg[20][0]/P0001 , \wishbone_bd_ram_mem0_reg[20][1]/P0001 , \wishbone_bd_ram_mem0_reg[20][2]/P0001 , \wishbone_bd_ram_mem0_reg[20][3]/P0001 , \wishbone_bd_ram_mem0_reg[20][4]/P0001 , \wishbone_bd_ram_mem0_reg[20][5]/P0001 , \wishbone_bd_ram_mem0_reg[20][6]/P0001 , \wishbone_bd_ram_mem0_reg[20][7]/P0001 , \wishbone_bd_ram_mem0_reg[210][0]/P0001 , \wishbone_bd_ram_mem0_reg[210][1]/P0001 , \wishbone_bd_ram_mem0_reg[210][2]/P0001 , \wishbone_bd_ram_mem0_reg[210][3]/P0001 , \wishbone_bd_ram_mem0_reg[210][4]/P0001 , \wishbone_bd_ram_mem0_reg[210][5]/P0001 , \wishbone_bd_ram_mem0_reg[210][6]/P0001 , \wishbone_bd_ram_mem0_reg[210][7]/P0001 , \wishbone_bd_ram_mem0_reg[211][0]/P0001 , \wishbone_bd_ram_mem0_reg[211][1]/P0001 , \wishbone_bd_ram_mem0_reg[211][2]/P0001 , \wishbone_bd_ram_mem0_reg[211][3]/P0001 , \wishbone_bd_ram_mem0_reg[211][4]/P0001 , \wishbone_bd_ram_mem0_reg[211][5]/P0001 , \wishbone_bd_ram_mem0_reg[211][6]/P0001 , \wishbone_bd_ram_mem0_reg[211][7]/P0001 , \wishbone_bd_ram_mem0_reg[212][0]/P0001 , \wishbone_bd_ram_mem0_reg[212][1]/P0001 , \wishbone_bd_ram_mem0_reg[212][2]/P0001 , \wishbone_bd_ram_mem0_reg[212][3]/P0001 , \wishbone_bd_ram_mem0_reg[212][4]/P0001 , \wishbone_bd_ram_mem0_reg[212][5]/P0001 , \wishbone_bd_ram_mem0_reg[212][6]/P0001 , \wishbone_bd_ram_mem0_reg[212][7]/P0001 , \wishbone_bd_ram_mem0_reg[213][0]/P0001 , \wishbone_bd_ram_mem0_reg[213][1]/P0001 , \wishbone_bd_ram_mem0_reg[213][2]/P0001 , \wishbone_bd_ram_mem0_reg[213][3]/P0001 , \wishbone_bd_ram_mem0_reg[213][4]/P0001 , \wishbone_bd_ram_mem0_reg[213][5]/P0001 , \wishbone_bd_ram_mem0_reg[213][6]/P0001 , \wishbone_bd_ram_mem0_reg[213][7]/P0001 , \wishbone_bd_ram_mem0_reg[214][0]/P0001 , \wishbone_bd_ram_mem0_reg[214][1]/P0001 , \wishbone_bd_ram_mem0_reg[214][2]/P0001 , \wishbone_bd_ram_mem0_reg[214][3]/P0001 , \wishbone_bd_ram_mem0_reg[214][4]/P0001 , \wishbone_bd_ram_mem0_reg[214][5]/P0001 , \wishbone_bd_ram_mem0_reg[214][6]/P0001 , \wishbone_bd_ram_mem0_reg[214][7]/P0001 , \wishbone_bd_ram_mem0_reg[215][0]/P0001 , \wishbone_bd_ram_mem0_reg[215][1]/P0001 , \wishbone_bd_ram_mem0_reg[215][2]/P0001 , \wishbone_bd_ram_mem0_reg[215][3]/P0001 , \wishbone_bd_ram_mem0_reg[215][4]/P0001 , \wishbone_bd_ram_mem0_reg[215][5]/P0001 , \wishbone_bd_ram_mem0_reg[215][6]/P0001 , \wishbone_bd_ram_mem0_reg[215][7]/P0001 , \wishbone_bd_ram_mem0_reg[216][0]/P0001 , \wishbone_bd_ram_mem0_reg[216][1]/P0001 , \wishbone_bd_ram_mem0_reg[216][2]/P0001 , \wishbone_bd_ram_mem0_reg[216][3]/P0001 , \wishbone_bd_ram_mem0_reg[216][4]/P0001 , \wishbone_bd_ram_mem0_reg[216][5]/P0001 , \wishbone_bd_ram_mem0_reg[216][6]/P0001 , \wishbone_bd_ram_mem0_reg[216][7]/P0001 , \wishbone_bd_ram_mem0_reg[217][0]/P0001 , \wishbone_bd_ram_mem0_reg[217][1]/P0001 , \wishbone_bd_ram_mem0_reg[217][2]/P0001 , \wishbone_bd_ram_mem0_reg[217][3]/P0001 , \wishbone_bd_ram_mem0_reg[217][4]/P0001 , \wishbone_bd_ram_mem0_reg[217][5]/P0001 , \wishbone_bd_ram_mem0_reg[217][6]/P0001 , \wishbone_bd_ram_mem0_reg[217][7]/P0001 , \wishbone_bd_ram_mem0_reg[218][0]/P0001 , \wishbone_bd_ram_mem0_reg[218][1]/P0001 , \wishbone_bd_ram_mem0_reg[218][2]/P0001 , \wishbone_bd_ram_mem0_reg[218][3]/P0001 , \wishbone_bd_ram_mem0_reg[218][4]/P0001 , \wishbone_bd_ram_mem0_reg[218][5]/P0001 , \wishbone_bd_ram_mem0_reg[218][6]/P0001 , \wishbone_bd_ram_mem0_reg[218][7]/P0001 , \wishbone_bd_ram_mem0_reg[219][0]/P0001 , \wishbone_bd_ram_mem0_reg[219][1]/P0001 , \wishbone_bd_ram_mem0_reg[219][2]/P0001 , \wishbone_bd_ram_mem0_reg[219][3]/P0001 , \wishbone_bd_ram_mem0_reg[219][4]/P0001 , \wishbone_bd_ram_mem0_reg[219][5]/P0001 , \wishbone_bd_ram_mem0_reg[219][6]/P0001 , \wishbone_bd_ram_mem0_reg[219][7]/P0001 , \wishbone_bd_ram_mem0_reg[21][0]/P0001 , \wishbone_bd_ram_mem0_reg[21][1]/P0001 , \wishbone_bd_ram_mem0_reg[21][2]/P0001 , \wishbone_bd_ram_mem0_reg[21][3]/P0001 , \wishbone_bd_ram_mem0_reg[21][4]/P0001 , \wishbone_bd_ram_mem0_reg[21][5]/P0001 , \wishbone_bd_ram_mem0_reg[21][6]/P0001 , \wishbone_bd_ram_mem0_reg[21][7]/P0001 , \wishbone_bd_ram_mem0_reg[220][0]/P0001 , \wishbone_bd_ram_mem0_reg[220][1]/P0001 , \wishbone_bd_ram_mem0_reg[220][2]/P0001 , \wishbone_bd_ram_mem0_reg[220][3]/P0001 , \wishbone_bd_ram_mem0_reg[220][4]/P0001 , \wishbone_bd_ram_mem0_reg[220][5]/P0001 , \wishbone_bd_ram_mem0_reg[220][6]/P0001 , \wishbone_bd_ram_mem0_reg[220][7]/P0001 , \wishbone_bd_ram_mem0_reg[221][0]/P0001 , \wishbone_bd_ram_mem0_reg[221][1]/P0001 , \wishbone_bd_ram_mem0_reg[221][2]/P0001 , \wishbone_bd_ram_mem0_reg[221][3]/P0001 , \wishbone_bd_ram_mem0_reg[221][4]/P0001 , \wishbone_bd_ram_mem0_reg[221][5]/P0001 , \wishbone_bd_ram_mem0_reg[221][6]/P0001 , \wishbone_bd_ram_mem0_reg[221][7]/P0001 , \wishbone_bd_ram_mem0_reg[222][0]/P0001 , \wishbone_bd_ram_mem0_reg[222][1]/P0001 , \wishbone_bd_ram_mem0_reg[222][2]/P0001 , \wishbone_bd_ram_mem0_reg[222][3]/P0001 , \wishbone_bd_ram_mem0_reg[222][4]/P0001 , \wishbone_bd_ram_mem0_reg[222][5]/P0001 , \wishbone_bd_ram_mem0_reg[222][6]/P0001 , \wishbone_bd_ram_mem0_reg[222][7]/P0001 , \wishbone_bd_ram_mem0_reg[223][0]/P0001 , \wishbone_bd_ram_mem0_reg[223][1]/P0001 , \wishbone_bd_ram_mem0_reg[223][2]/P0001 , \wishbone_bd_ram_mem0_reg[223][3]/P0001 , \wishbone_bd_ram_mem0_reg[223][4]/P0001 , \wishbone_bd_ram_mem0_reg[223][5]/P0001 , \wishbone_bd_ram_mem0_reg[223][6]/P0001 , \wishbone_bd_ram_mem0_reg[223][7]/P0001 , \wishbone_bd_ram_mem0_reg[224][0]/P0001 , \wishbone_bd_ram_mem0_reg[224][1]/P0001 , \wishbone_bd_ram_mem0_reg[224][2]/P0001 , \wishbone_bd_ram_mem0_reg[224][3]/P0001 , \wishbone_bd_ram_mem0_reg[224][4]/P0001 , \wishbone_bd_ram_mem0_reg[224][5]/P0001 , \wishbone_bd_ram_mem0_reg[224][6]/P0001 , \wishbone_bd_ram_mem0_reg[224][7]/P0001 , \wishbone_bd_ram_mem0_reg[225][0]/P0001 , \wishbone_bd_ram_mem0_reg[225][1]/P0001 , \wishbone_bd_ram_mem0_reg[225][2]/P0001 , \wishbone_bd_ram_mem0_reg[225][3]/P0001 , \wishbone_bd_ram_mem0_reg[225][4]/P0001 , \wishbone_bd_ram_mem0_reg[225][5]/P0001 , \wishbone_bd_ram_mem0_reg[225][6]/P0001 , \wishbone_bd_ram_mem0_reg[225][7]/P0001 , \wishbone_bd_ram_mem0_reg[226][0]/P0001 , \wishbone_bd_ram_mem0_reg[226][1]/P0001 , \wishbone_bd_ram_mem0_reg[226][2]/P0001 , \wishbone_bd_ram_mem0_reg[226][3]/P0001 , \wishbone_bd_ram_mem0_reg[226][4]/P0001 , \wishbone_bd_ram_mem0_reg[226][5]/P0001 , \wishbone_bd_ram_mem0_reg[226][6]/P0001 , \wishbone_bd_ram_mem0_reg[226][7]/P0001 , \wishbone_bd_ram_mem0_reg[227][0]/P0001 , \wishbone_bd_ram_mem0_reg[227][1]/P0001 , \wishbone_bd_ram_mem0_reg[227][2]/P0001 , \wishbone_bd_ram_mem0_reg[227][3]/P0001 , \wishbone_bd_ram_mem0_reg[227][4]/P0001 , \wishbone_bd_ram_mem0_reg[227][5]/P0001 , \wishbone_bd_ram_mem0_reg[227][6]/P0001 , \wishbone_bd_ram_mem0_reg[227][7]/P0001 , \wishbone_bd_ram_mem0_reg[228][0]/P0001 , \wishbone_bd_ram_mem0_reg[228][1]/P0001 , \wishbone_bd_ram_mem0_reg[228][2]/P0001 , \wishbone_bd_ram_mem0_reg[228][3]/P0001 , \wishbone_bd_ram_mem0_reg[228][4]/P0001 , \wishbone_bd_ram_mem0_reg[228][5]/P0001 , \wishbone_bd_ram_mem0_reg[228][6]/P0001 , \wishbone_bd_ram_mem0_reg[228][7]/P0001 , \wishbone_bd_ram_mem0_reg[229][0]/P0001 , \wishbone_bd_ram_mem0_reg[229][1]/P0001 , \wishbone_bd_ram_mem0_reg[229][2]/P0001 , \wishbone_bd_ram_mem0_reg[229][3]/P0001 , \wishbone_bd_ram_mem0_reg[229][4]/P0001 , \wishbone_bd_ram_mem0_reg[229][5]/P0001 , \wishbone_bd_ram_mem0_reg[229][6]/P0001 , \wishbone_bd_ram_mem0_reg[229][7]/P0001 , \wishbone_bd_ram_mem0_reg[22][0]/P0001 , \wishbone_bd_ram_mem0_reg[22][1]/P0001 , \wishbone_bd_ram_mem0_reg[22][2]/P0001 , \wishbone_bd_ram_mem0_reg[22][3]/P0001 , \wishbone_bd_ram_mem0_reg[22][4]/P0001 , \wishbone_bd_ram_mem0_reg[22][5]/P0001 , \wishbone_bd_ram_mem0_reg[22][6]/P0001 , \wishbone_bd_ram_mem0_reg[22][7]/P0001 , \wishbone_bd_ram_mem0_reg[230][0]/P0001 , \wishbone_bd_ram_mem0_reg[230][1]/P0001 , \wishbone_bd_ram_mem0_reg[230][2]/P0001 , \wishbone_bd_ram_mem0_reg[230][3]/P0001 , \wishbone_bd_ram_mem0_reg[230][4]/P0001 , \wishbone_bd_ram_mem0_reg[230][5]/P0001 , \wishbone_bd_ram_mem0_reg[230][6]/P0001 , \wishbone_bd_ram_mem0_reg[230][7]/P0001 , \wishbone_bd_ram_mem0_reg[231][0]/P0001 , \wishbone_bd_ram_mem0_reg[231][1]/P0001 , \wishbone_bd_ram_mem0_reg[231][2]/P0001 , \wishbone_bd_ram_mem0_reg[231][3]/P0001 , \wishbone_bd_ram_mem0_reg[231][4]/P0001 , \wishbone_bd_ram_mem0_reg[231][5]/P0001 , \wishbone_bd_ram_mem0_reg[231][6]/P0001 , \wishbone_bd_ram_mem0_reg[231][7]/P0001 , \wishbone_bd_ram_mem0_reg[232][0]/P0001 , \wishbone_bd_ram_mem0_reg[232][1]/P0001 , \wishbone_bd_ram_mem0_reg[232][2]/P0001 , \wishbone_bd_ram_mem0_reg[232][3]/P0001 , \wishbone_bd_ram_mem0_reg[232][4]/P0001 , \wishbone_bd_ram_mem0_reg[232][5]/P0001 , \wishbone_bd_ram_mem0_reg[232][6]/P0001 , \wishbone_bd_ram_mem0_reg[232][7]/P0001 , \wishbone_bd_ram_mem0_reg[233][0]/P0001 , \wishbone_bd_ram_mem0_reg[233][1]/P0001 , \wishbone_bd_ram_mem0_reg[233][2]/P0001 , \wishbone_bd_ram_mem0_reg[233][3]/P0001 , \wishbone_bd_ram_mem0_reg[233][4]/P0001 , \wishbone_bd_ram_mem0_reg[233][5]/P0001 , \wishbone_bd_ram_mem0_reg[233][6]/P0001 , \wishbone_bd_ram_mem0_reg[233][7]/P0001 , \wishbone_bd_ram_mem0_reg[234][0]/P0001 , \wishbone_bd_ram_mem0_reg[234][1]/P0001 , \wishbone_bd_ram_mem0_reg[234][2]/P0001 , \wishbone_bd_ram_mem0_reg[234][3]/P0001 , \wishbone_bd_ram_mem0_reg[234][4]/P0001 , \wishbone_bd_ram_mem0_reg[234][5]/P0001 , \wishbone_bd_ram_mem0_reg[234][6]/P0001 , \wishbone_bd_ram_mem0_reg[234][7]/P0001 , \wishbone_bd_ram_mem0_reg[235][0]/P0001 , \wishbone_bd_ram_mem0_reg[235][1]/P0001 , \wishbone_bd_ram_mem0_reg[235][2]/P0001 , \wishbone_bd_ram_mem0_reg[235][3]/P0001 , \wishbone_bd_ram_mem0_reg[235][4]/P0001 , \wishbone_bd_ram_mem0_reg[235][5]/P0001 , \wishbone_bd_ram_mem0_reg[235][6]/P0001 , \wishbone_bd_ram_mem0_reg[235][7]/P0001 , \wishbone_bd_ram_mem0_reg[236][0]/P0001 , \wishbone_bd_ram_mem0_reg[236][1]/P0001 , \wishbone_bd_ram_mem0_reg[236][2]/P0001 , \wishbone_bd_ram_mem0_reg[236][3]/P0001 , \wishbone_bd_ram_mem0_reg[236][4]/P0001 , \wishbone_bd_ram_mem0_reg[236][5]/P0001 , \wishbone_bd_ram_mem0_reg[236][6]/P0001 , \wishbone_bd_ram_mem0_reg[236][7]/P0001 , \wishbone_bd_ram_mem0_reg[237][0]/P0001 , \wishbone_bd_ram_mem0_reg[237][1]/P0001 , \wishbone_bd_ram_mem0_reg[237][2]/P0001 , \wishbone_bd_ram_mem0_reg[237][3]/P0001 , \wishbone_bd_ram_mem0_reg[237][4]/P0001 , \wishbone_bd_ram_mem0_reg[237][5]/P0001 , \wishbone_bd_ram_mem0_reg[237][6]/P0001 , \wishbone_bd_ram_mem0_reg[237][7]/P0001 , \wishbone_bd_ram_mem0_reg[238][0]/P0001 , \wishbone_bd_ram_mem0_reg[238][1]/P0001 , \wishbone_bd_ram_mem0_reg[238][2]/P0001 , \wishbone_bd_ram_mem0_reg[238][3]/P0001 , \wishbone_bd_ram_mem0_reg[238][4]/P0001 , \wishbone_bd_ram_mem0_reg[238][5]/P0001 , \wishbone_bd_ram_mem0_reg[238][6]/P0001 , \wishbone_bd_ram_mem0_reg[238][7]/P0001 , \wishbone_bd_ram_mem0_reg[239][0]/P0001 , \wishbone_bd_ram_mem0_reg[239][1]/P0001 , \wishbone_bd_ram_mem0_reg[239][2]/P0001 , \wishbone_bd_ram_mem0_reg[239][3]/P0001 , \wishbone_bd_ram_mem0_reg[239][4]/P0001 , \wishbone_bd_ram_mem0_reg[239][5]/P0001 , \wishbone_bd_ram_mem0_reg[239][6]/P0001 , \wishbone_bd_ram_mem0_reg[239][7]/P0001 , \wishbone_bd_ram_mem0_reg[23][0]/P0001 , \wishbone_bd_ram_mem0_reg[23][1]/P0001 , \wishbone_bd_ram_mem0_reg[23][2]/P0001 , \wishbone_bd_ram_mem0_reg[23][3]/P0001 , \wishbone_bd_ram_mem0_reg[23][4]/P0001 , \wishbone_bd_ram_mem0_reg[23][5]/P0001 , \wishbone_bd_ram_mem0_reg[23][6]/P0001 , \wishbone_bd_ram_mem0_reg[23][7]/P0001 , \wishbone_bd_ram_mem0_reg[240][0]/P0001 , \wishbone_bd_ram_mem0_reg[240][1]/P0001 , \wishbone_bd_ram_mem0_reg[240][2]/P0001 , \wishbone_bd_ram_mem0_reg[240][3]/P0001 , \wishbone_bd_ram_mem0_reg[240][4]/P0001 , \wishbone_bd_ram_mem0_reg[240][5]/P0001 , \wishbone_bd_ram_mem0_reg[240][6]/P0001 , \wishbone_bd_ram_mem0_reg[240][7]/P0001 , \wishbone_bd_ram_mem0_reg[241][0]/P0001 , \wishbone_bd_ram_mem0_reg[241][1]/P0001 , \wishbone_bd_ram_mem0_reg[241][2]/P0001 , \wishbone_bd_ram_mem0_reg[241][3]/P0001 , \wishbone_bd_ram_mem0_reg[241][4]/P0001 , \wishbone_bd_ram_mem0_reg[241][5]/P0001 , \wishbone_bd_ram_mem0_reg[241][6]/P0001 , \wishbone_bd_ram_mem0_reg[241][7]/P0001 , \wishbone_bd_ram_mem0_reg[242][0]/P0001 , \wishbone_bd_ram_mem0_reg[242][1]/P0001 , \wishbone_bd_ram_mem0_reg[242][2]/P0001 , \wishbone_bd_ram_mem0_reg[242][3]/P0001 , \wishbone_bd_ram_mem0_reg[242][4]/P0001 , \wishbone_bd_ram_mem0_reg[242][5]/P0001 , \wishbone_bd_ram_mem0_reg[242][6]/P0001 , \wishbone_bd_ram_mem0_reg[242][7]/P0001 , \wishbone_bd_ram_mem0_reg[243][0]/P0001 , \wishbone_bd_ram_mem0_reg[243][1]/P0001 , \wishbone_bd_ram_mem0_reg[243][2]/P0001 , \wishbone_bd_ram_mem0_reg[243][3]/P0001 , \wishbone_bd_ram_mem0_reg[243][4]/P0001 , \wishbone_bd_ram_mem0_reg[243][5]/P0001 , \wishbone_bd_ram_mem0_reg[243][6]/P0001 , \wishbone_bd_ram_mem0_reg[243][7]/P0001 , \wishbone_bd_ram_mem0_reg[244][0]/P0001 , \wishbone_bd_ram_mem0_reg[244][1]/P0001 , \wishbone_bd_ram_mem0_reg[244][2]/P0001 , \wishbone_bd_ram_mem0_reg[244][3]/P0001 , \wishbone_bd_ram_mem0_reg[244][4]/P0001 , \wishbone_bd_ram_mem0_reg[244][5]/P0001 , \wishbone_bd_ram_mem0_reg[244][6]/P0001 , \wishbone_bd_ram_mem0_reg[244][7]/P0001 , \wishbone_bd_ram_mem0_reg[245][0]/P0001 , \wishbone_bd_ram_mem0_reg[245][1]/P0001 , \wishbone_bd_ram_mem0_reg[245][2]/P0001 , \wishbone_bd_ram_mem0_reg[245][3]/P0001 , \wishbone_bd_ram_mem0_reg[245][4]/P0001 , \wishbone_bd_ram_mem0_reg[245][5]/P0001 , \wishbone_bd_ram_mem0_reg[245][6]/P0001 , \wishbone_bd_ram_mem0_reg[245][7]/P0001 , \wishbone_bd_ram_mem0_reg[246][0]/P0001 , \wishbone_bd_ram_mem0_reg[246][1]/P0001 , \wishbone_bd_ram_mem0_reg[246][2]/P0001 , \wishbone_bd_ram_mem0_reg[246][3]/P0001 , \wishbone_bd_ram_mem0_reg[246][4]/P0001 , \wishbone_bd_ram_mem0_reg[246][5]/P0001 , \wishbone_bd_ram_mem0_reg[246][6]/P0001 , \wishbone_bd_ram_mem0_reg[246][7]/P0001 , \wishbone_bd_ram_mem0_reg[247][0]/P0001 , \wishbone_bd_ram_mem0_reg[247][1]/P0001 , \wishbone_bd_ram_mem0_reg[247][2]/P0001 , \wishbone_bd_ram_mem0_reg[247][3]/P0001 , \wishbone_bd_ram_mem0_reg[247][4]/P0001 , \wishbone_bd_ram_mem0_reg[247][5]/P0001 , \wishbone_bd_ram_mem0_reg[247][6]/P0001 , \wishbone_bd_ram_mem0_reg[247][7]/P0001 , \wishbone_bd_ram_mem0_reg[248][0]/P0001 , \wishbone_bd_ram_mem0_reg[248][1]/P0001 , \wishbone_bd_ram_mem0_reg[248][2]/P0001 , \wishbone_bd_ram_mem0_reg[248][3]/P0001 , \wishbone_bd_ram_mem0_reg[248][4]/P0001 , \wishbone_bd_ram_mem0_reg[248][5]/P0001 , \wishbone_bd_ram_mem0_reg[248][6]/P0001 , \wishbone_bd_ram_mem0_reg[248][7]/P0001 , \wishbone_bd_ram_mem0_reg[249][0]/P0001 , \wishbone_bd_ram_mem0_reg[249][1]/P0001 , \wishbone_bd_ram_mem0_reg[249][2]/P0001 , \wishbone_bd_ram_mem0_reg[249][3]/P0001 , \wishbone_bd_ram_mem0_reg[249][4]/P0001 , \wishbone_bd_ram_mem0_reg[249][5]/P0001 , \wishbone_bd_ram_mem0_reg[249][6]/P0001 , \wishbone_bd_ram_mem0_reg[249][7]/P0001 , \wishbone_bd_ram_mem0_reg[24][0]/P0001 , \wishbone_bd_ram_mem0_reg[24][1]/P0001 , \wishbone_bd_ram_mem0_reg[24][2]/P0001 , \wishbone_bd_ram_mem0_reg[24][3]/P0001 , \wishbone_bd_ram_mem0_reg[24][4]/P0001 , \wishbone_bd_ram_mem0_reg[24][5]/P0001 , \wishbone_bd_ram_mem0_reg[24][6]/P0001 , \wishbone_bd_ram_mem0_reg[24][7]/P0001 , \wishbone_bd_ram_mem0_reg[250][0]/P0001 , \wishbone_bd_ram_mem0_reg[250][1]/P0001 , \wishbone_bd_ram_mem0_reg[250][2]/P0001 , \wishbone_bd_ram_mem0_reg[250][3]/P0001 , \wishbone_bd_ram_mem0_reg[250][4]/P0001 , \wishbone_bd_ram_mem0_reg[250][5]/P0001 , \wishbone_bd_ram_mem0_reg[250][6]/P0001 , \wishbone_bd_ram_mem0_reg[250][7]/P0001 , \wishbone_bd_ram_mem0_reg[251][0]/P0001 , \wishbone_bd_ram_mem0_reg[251][1]/P0001 , \wishbone_bd_ram_mem0_reg[251][2]/P0001 , \wishbone_bd_ram_mem0_reg[251][3]/P0001 , \wishbone_bd_ram_mem0_reg[251][4]/P0001 , \wishbone_bd_ram_mem0_reg[251][5]/P0001 , \wishbone_bd_ram_mem0_reg[251][6]/P0001 , \wishbone_bd_ram_mem0_reg[251][7]/P0001 , \wishbone_bd_ram_mem0_reg[252][0]/P0001 , \wishbone_bd_ram_mem0_reg[252][1]/P0001 , \wishbone_bd_ram_mem0_reg[252][2]/P0001 , \wishbone_bd_ram_mem0_reg[252][3]/P0001 , \wishbone_bd_ram_mem0_reg[252][4]/P0001 , \wishbone_bd_ram_mem0_reg[252][5]/P0001 , \wishbone_bd_ram_mem0_reg[252][6]/P0001 , \wishbone_bd_ram_mem0_reg[252][7]/P0001 , \wishbone_bd_ram_mem0_reg[253][0]/P0001 , \wishbone_bd_ram_mem0_reg[253][1]/P0001 , \wishbone_bd_ram_mem0_reg[253][2]/P0001 , \wishbone_bd_ram_mem0_reg[253][3]/P0001 , \wishbone_bd_ram_mem0_reg[253][4]/P0001 , \wishbone_bd_ram_mem0_reg[253][5]/P0001 , \wishbone_bd_ram_mem0_reg[253][6]/P0001 , \wishbone_bd_ram_mem0_reg[253][7]/P0001 , \wishbone_bd_ram_mem0_reg[254][0]/P0001 , \wishbone_bd_ram_mem0_reg[254][1]/P0001 , \wishbone_bd_ram_mem0_reg[254][2]/P0001 , \wishbone_bd_ram_mem0_reg[254][3]/P0001 , \wishbone_bd_ram_mem0_reg[254][4]/P0001 , \wishbone_bd_ram_mem0_reg[254][5]/P0001 , \wishbone_bd_ram_mem0_reg[254][6]/P0001 , \wishbone_bd_ram_mem0_reg[254][7]/P0001 , \wishbone_bd_ram_mem0_reg[255][0]/P0001 , \wishbone_bd_ram_mem0_reg[255][1]/P0001 , \wishbone_bd_ram_mem0_reg[255][2]/P0001 , \wishbone_bd_ram_mem0_reg[255][3]/P0001 , \wishbone_bd_ram_mem0_reg[255][4]/P0001 , \wishbone_bd_ram_mem0_reg[255][5]/P0001 , \wishbone_bd_ram_mem0_reg[255][6]/P0001 , \wishbone_bd_ram_mem0_reg[255][7]/P0001 , \wishbone_bd_ram_mem0_reg[25][0]/P0001 , \wishbone_bd_ram_mem0_reg[25][1]/P0001 , \wishbone_bd_ram_mem0_reg[25][2]/P0001 , \wishbone_bd_ram_mem0_reg[25][3]/P0001 , \wishbone_bd_ram_mem0_reg[25][4]/P0001 , \wishbone_bd_ram_mem0_reg[25][5]/P0001 , \wishbone_bd_ram_mem0_reg[25][6]/P0001 , \wishbone_bd_ram_mem0_reg[25][7]/P0001 , \wishbone_bd_ram_mem0_reg[26][0]/P0001 , \wishbone_bd_ram_mem0_reg[26][1]/P0001 , \wishbone_bd_ram_mem0_reg[26][2]/P0001 , \wishbone_bd_ram_mem0_reg[26][3]/P0001 , \wishbone_bd_ram_mem0_reg[26][4]/P0001 , \wishbone_bd_ram_mem0_reg[26][5]/P0001 , \wishbone_bd_ram_mem0_reg[26][6]/P0001 , \wishbone_bd_ram_mem0_reg[26][7]/P0001 , \wishbone_bd_ram_mem0_reg[27][0]/P0001 , \wishbone_bd_ram_mem0_reg[27][1]/P0001 , \wishbone_bd_ram_mem0_reg[27][2]/P0001 , \wishbone_bd_ram_mem0_reg[27][3]/P0001 , \wishbone_bd_ram_mem0_reg[27][4]/P0001 , \wishbone_bd_ram_mem0_reg[27][5]/P0001 , \wishbone_bd_ram_mem0_reg[27][6]/P0001 , \wishbone_bd_ram_mem0_reg[27][7]/P0001 , \wishbone_bd_ram_mem0_reg[28][0]/P0001 , \wishbone_bd_ram_mem0_reg[28][1]/P0001 , \wishbone_bd_ram_mem0_reg[28][2]/P0001 , \wishbone_bd_ram_mem0_reg[28][3]/P0001 , \wishbone_bd_ram_mem0_reg[28][4]/P0001 , \wishbone_bd_ram_mem0_reg[28][5]/P0001 , \wishbone_bd_ram_mem0_reg[28][6]/P0001 , \wishbone_bd_ram_mem0_reg[28][7]/P0001 , \wishbone_bd_ram_mem0_reg[29][0]/P0001 , \wishbone_bd_ram_mem0_reg[29][1]/P0001 , \wishbone_bd_ram_mem0_reg[29][2]/P0001 , \wishbone_bd_ram_mem0_reg[29][3]/P0001 , \wishbone_bd_ram_mem0_reg[29][4]/P0001 , \wishbone_bd_ram_mem0_reg[29][5]/P0001 , \wishbone_bd_ram_mem0_reg[29][6]/P0001 , \wishbone_bd_ram_mem0_reg[29][7]/P0001 , \wishbone_bd_ram_mem0_reg[2][0]/P0001 , \wishbone_bd_ram_mem0_reg[2][1]/P0001 , \wishbone_bd_ram_mem0_reg[2][2]/P0001 , \wishbone_bd_ram_mem0_reg[2][3]/P0001 , \wishbone_bd_ram_mem0_reg[2][4]/P0001 , \wishbone_bd_ram_mem0_reg[2][5]/P0001 , \wishbone_bd_ram_mem0_reg[2][6]/P0001 , \wishbone_bd_ram_mem0_reg[2][7]/P0001 , \wishbone_bd_ram_mem0_reg[30][0]/P0001 , \wishbone_bd_ram_mem0_reg[30][1]/P0001 , \wishbone_bd_ram_mem0_reg[30][2]/P0001 , \wishbone_bd_ram_mem0_reg[30][3]/P0001 , \wishbone_bd_ram_mem0_reg[30][4]/P0001 , \wishbone_bd_ram_mem0_reg[30][5]/P0001 , \wishbone_bd_ram_mem0_reg[30][6]/P0001 , \wishbone_bd_ram_mem0_reg[30][7]/P0001 , \wishbone_bd_ram_mem0_reg[31][0]/P0001 , \wishbone_bd_ram_mem0_reg[31][1]/P0001 , \wishbone_bd_ram_mem0_reg[31][2]/P0001 , \wishbone_bd_ram_mem0_reg[31][3]/P0001 , \wishbone_bd_ram_mem0_reg[31][4]/P0001 , \wishbone_bd_ram_mem0_reg[31][5]/P0001 , \wishbone_bd_ram_mem0_reg[31][6]/P0001 , \wishbone_bd_ram_mem0_reg[31][7]/P0001 , \wishbone_bd_ram_mem0_reg[32][0]/P0001 , \wishbone_bd_ram_mem0_reg[32][1]/P0001 , \wishbone_bd_ram_mem0_reg[32][2]/P0001 , \wishbone_bd_ram_mem0_reg[32][3]/P0001 , \wishbone_bd_ram_mem0_reg[32][4]/P0001 , \wishbone_bd_ram_mem0_reg[32][5]/P0001 , \wishbone_bd_ram_mem0_reg[32][6]/P0001 , \wishbone_bd_ram_mem0_reg[32][7]/P0001 , \wishbone_bd_ram_mem0_reg[33][0]/P0001 , \wishbone_bd_ram_mem0_reg[33][1]/P0001 , \wishbone_bd_ram_mem0_reg[33][2]/P0001 , \wishbone_bd_ram_mem0_reg[33][3]/P0001 , \wishbone_bd_ram_mem0_reg[33][4]/P0001 , \wishbone_bd_ram_mem0_reg[33][5]/P0001 , \wishbone_bd_ram_mem0_reg[33][6]/P0001 , \wishbone_bd_ram_mem0_reg[33][7]/P0001 , \wishbone_bd_ram_mem0_reg[34][0]/P0001 , \wishbone_bd_ram_mem0_reg[34][1]/P0001 , \wishbone_bd_ram_mem0_reg[34][2]/P0001 , \wishbone_bd_ram_mem0_reg[34][3]/P0001 , \wishbone_bd_ram_mem0_reg[34][4]/P0001 , \wishbone_bd_ram_mem0_reg[34][5]/P0001 , \wishbone_bd_ram_mem0_reg[34][6]/P0001 , \wishbone_bd_ram_mem0_reg[34][7]/P0001 , \wishbone_bd_ram_mem0_reg[35][0]/P0001 , \wishbone_bd_ram_mem0_reg[35][1]/P0001 , \wishbone_bd_ram_mem0_reg[35][2]/P0001 , \wishbone_bd_ram_mem0_reg[35][3]/P0001 , \wishbone_bd_ram_mem0_reg[35][4]/P0001 , \wishbone_bd_ram_mem0_reg[35][5]/P0001 , \wishbone_bd_ram_mem0_reg[35][6]/P0001 , \wishbone_bd_ram_mem0_reg[35][7]/P0001 , \wishbone_bd_ram_mem0_reg[36][0]/P0001 , \wishbone_bd_ram_mem0_reg[36][1]/P0001 , \wishbone_bd_ram_mem0_reg[36][2]/P0001 , \wishbone_bd_ram_mem0_reg[36][3]/P0001 , \wishbone_bd_ram_mem0_reg[36][4]/P0001 , \wishbone_bd_ram_mem0_reg[36][5]/P0001 , \wishbone_bd_ram_mem0_reg[36][6]/P0001 , \wishbone_bd_ram_mem0_reg[36][7]/P0001 , \wishbone_bd_ram_mem0_reg[37][0]/P0001 , \wishbone_bd_ram_mem0_reg[37][1]/P0001 , \wishbone_bd_ram_mem0_reg[37][2]/P0001 , \wishbone_bd_ram_mem0_reg[37][3]/P0001 , \wishbone_bd_ram_mem0_reg[37][4]/P0001 , \wishbone_bd_ram_mem0_reg[37][5]/P0001 , \wishbone_bd_ram_mem0_reg[37][6]/P0001 , \wishbone_bd_ram_mem0_reg[37][7]/P0001 , \wishbone_bd_ram_mem0_reg[38][0]/P0001 , \wishbone_bd_ram_mem0_reg[38][1]/P0001 , \wishbone_bd_ram_mem0_reg[38][2]/P0001 , \wishbone_bd_ram_mem0_reg[38][3]/P0001 , \wishbone_bd_ram_mem0_reg[38][4]/P0001 , \wishbone_bd_ram_mem0_reg[38][5]/P0001 , \wishbone_bd_ram_mem0_reg[38][6]/P0001 , \wishbone_bd_ram_mem0_reg[38][7]/P0001 , \wishbone_bd_ram_mem0_reg[39][0]/P0001 , \wishbone_bd_ram_mem0_reg[39][1]/P0001 , \wishbone_bd_ram_mem0_reg[39][2]/P0001 , \wishbone_bd_ram_mem0_reg[39][3]/P0001 , \wishbone_bd_ram_mem0_reg[39][4]/P0001 , \wishbone_bd_ram_mem0_reg[39][5]/P0001 , \wishbone_bd_ram_mem0_reg[39][6]/P0001 , \wishbone_bd_ram_mem0_reg[39][7]/P0001 , \wishbone_bd_ram_mem0_reg[3][0]/P0001 , \wishbone_bd_ram_mem0_reg[3][1]/P0001 , \wishbone_bd_ram_mem0_reg[3][2]/P0001 , \wishbone_bd_ram_mem0_reg[3][3]/P0001 , \wishbone_bd_ram_mem0_reg[3][4]/P0001 , \wishbone_bd_ram_mem0_reg[3][5]/P0001 , \wishbone_bd_ram_mem0_reg[3][6]/P0001 , \wishbone_bd_ram_mem0_reg[3][7]/P0001 , \wishbone_bd_ram_mem0_reg[40][0]/P0001 , \wishbone_bd_ram_mem0_reg[40][1]/P0001 , \wishbone_bd_ram_mem0_reg[40][2]/P0001 , \wishbone_bd_ram_mem0_reg[40][3]/P0001 , \wishbone_bd_ram_mem0_reg[40][4]/P0001 , \wishbone_bd_ram_mem0_reg[40][5]/P0001 , \wishbone_bd_ram_mem0_reg[40][6]/P0001 , \wishbone_bd_ram_mem0_reg[40][7]/P0001 , \wishbone_bd_ram_mem0_reg[41][0]/P0001 , \wishbone_bd_ram_mem0_reg[41][1]/P0001 , \wishbone_bd_ram_mem0_reg[41][2]/P0001 , \wishbone_bd_ram_mem0_reg[41][3]/P0001 , \wishbone_bd_ram_mem0_reg[41][4]/P0001 , \wishbone_bd_ram_mem0_reg[41][5]/P0001 , \wishbone_bd_ram_mem0_reg[41][6]/P0001 , \wishbone_bd_ram_mem0_reg[41][7]/P0001 , \wishbone_bd_ram_mem0_reg[42][0]/P0001 , \wishbone_bd_ram_mem0_reg[42][1]/P0001 , \wishbone_bd_ram_mem0_reg[42][2]/P0001 , \wishbone_bd_ram_mem0_reg[42][3]/P0001 , \wishbone_bd_ram_mem0_reg[42][4]/P0001 , \wishbone_bd_ram_mem0_reg[42][5]/P0001 , \wishbone_bd_ram_mem0_reg[42][6]/P0001 , \wishbone_bd_ram_mem0_reg[42][7]/P0001 , \wishbone_bd_ram_mem0_reg[43][0]/P0001 , \wishbone_bd_ram_mem0_reg[43][1]/P0001 , \wishbone_bd_ram_mem0_reg[43][2]/P0001 , \wishbone_bd_ram_mem0_reg[43][3]/P0001 , \wishbone_bd_ram_mem0_reg[43][4]/P0001 , \wishbone_bd_ram_mem0_reg[43][5]/P0001 , \wishbone_bd_ram_mem0_reg[43][6]/P0001 , \wishbone_bd_ram_mem0_reg[43][7]/P0001 , \wishbone_bd_ram_mem0_reg[44][0]/P0001 , \wishbone_bd_ram_mem0_reg[44][1]/P0001 , \wishbone_bd_ram_mem0_reg[44][2]/P0001 , \wishbone_bd_ram_mem0_reg[44][3]/P0001 , \wishbone_bd_ram_mem0_reg[44][4]/P0001 , \wishbone_bd_ram_mem0_reg[44][5]/P0001 , \wishbone_bd_ram_mem0_reg[44][6]/P0001 , \wishbone_bd_ram_mem0_reg[44][7]/P0001 , \wishbone_bd_ram_mem0_reg[45][0]/P0001 , \wishbone_bd_ram_mem0_reg[45][1]/P0001 , \wishbone_bd_ram_mem0_reg[45][2]/P0001 , \wishbone_bd_ram_mem0_reg[45][3]/P0001 , \wishbone_bd_ram_mem0_reg[45][4]/P0001 , \wishbone_bd_ram_mem0_reg[45][5]/P0001 , \wishbone_bd_ram_mem0_reg[45][6]/P0001 , \wishbone_bd_ram_mem0_reg[45][7]/P0001 , \wishbone_bd_ram_mem0_reg[46][0]/P0001 , \wishbone_bd_ram_mem0_reg[46][1]/P0001 , \wishbone_bd_ram_mem0_reg[46][2]/P0001 , \wishbone_bd_ram_mem0_reg[46][3]/P0001 , \wishbone_bd_ram_mem0_reg[46][4]/P0001 , \wishbone_bd_ram_mem0_reg[46][5]/P0001 , \wishbone_bd_ram_mem0_reg[46][6]/P0001 , \wishbone_bd_ram_mem0_reg[46][7]/P0001 , \wishbone_bd_ram_mem0_reg[47][0]/P0001 , \wishbone_bd_ram_mem0_reg[47][1]/P0001 , \wishbone_bd_ram_mem0_reg[47][2]/P0001 , \wishbone_bd_ram_mem0_reg[47][3]/P0001 , \wishbone_bd_ram_mem0_reg[47][4]/P0001 , \wishbone_bd_ram_mem0_reg[47][5]/P0001 , \wishbone_bd_ram_mem0_reg[47][6]/P0001 , \wishbone_bd_ram_mem0_reg[47][7]/P0001 , \wishbone_bd_ram_mem0_reg[48][0]/P0001 , \wishbone_bd_ram_mem0_reg[48][1]/P0001 , \wishbone_bd_ram_mem0_reg[48][2]/P0001 , \wishbone_bd_ram_mem0_reg[48][3]/P0001 , \wishbone_bd_ram_mem0_reg[48][4]/P0001 , \wishbone_bd_ram_mem0_reg[48][5]/P0001 , \wishbone_bd_ram_mem0_reg[48][6]/P0001 , \wishbone_bd_ram_mem0_reg[48][7]/P0001 , \wishbone_bd_ram_mem0_reg[49][0]/P0001 , \wishbone_bd_ram_mem0_reg[49][1]/P0001 , \wishbone_bd_ram_mem0_reg[49][2]/P0001 , \wishbone_bd_ram_mem0_reg[49][3]/P0001 , \wishbone_bd_ram_mem0_reg[49][4]/P0001 , \wishbone_bd_ram_mem0_reg[49][5]/P0001 , \wishbone_bd_ram_mem0_reg[49][6]/P0001 , \wishbone_bd_ram_mem0_reg[49][7]/P0001 , \wishbone_bd_ram_mem0_reg[4][0]/P0001 , \wishbone_bd_ram_mem0_reg[4][1]/P0001 , \wishbone_bd_ram_mem0_reg[4][2]/P0001 , \wishbone_bd_ram_mem0_reg[4][3]/P0001 , \wishbone_bd_ram_mem0_reg[4][4]/P0001 , \wishbone_bd_ram_mem0_reg[4][5]/P0001 , \wishbone_bd_ram_mem0_reg[4][6]/P0001 , \wishbone_bd_ram_mem0_reg[4][7]/P0001 , \wishbone_bd_ram_mem0_reg[50][0]/P0001 , \wishbone_bd_ram_mem0_reg[50][1]/P0001 , \wishbone_bd_ram_mem0_reg[50][2]/P0001 , \wishbone_bd_ram_mem0_reg[50][3]/P0001 , \wishbone_bd_ram_mem0_reg[50][4]/P0001 , \wishbone_bd_ram_mem0_reg[50][5]/P0001 , \wishbone_bd_ram_mem0_reg[50][6]/P0001 , \wishbone_bd_ram_mem0_reg[50][7]/P0001 , \wishbone_bd_ram_mem0_reg[51][0]/P0001 , \wishbone_bd_ram_mem0_reg[51][1]/P0001 , \wishbone_bd_ram_mem0_reg[51][2]/P0001 , \wishbone_bd_ram_mem0_reg[51][3]/P0001 , \wishbone_bd_ram_mem0_reg[51][4]/P0001 , \wishbone_bd_ram_mem0_reg[51][5]/P0001 , \wishbone_bd_ram_mem0_reg[51][6]/P0001 , \wishbone_bd_ram_mem0_reg[51][7]/P0001 , \wishbone_bd_ram_mem0_reg[52][0]/P0001 , \wishbone_bd_ram_mem0_reg[52][1]/P0001 , \wishbone_bd_ram_mem0_reg[52][2]/P0001 , \wishbone_bd_ram_mem0_reg[52][3]/P0001 , \wishbone_bd_ram_mem0_reg[52][4]/P0001 , \wishbone_bd_ram_mem0_reg[52][5]/P0001 , \wishbone_bd_ram_mem0_reg[52][6]/P0001 , \wishbone_bd_ram_mem0_reg[52][7]/P0001 , \wishbone_bd_ram_mem0_reg[53][0]/P0001 , \wishbone_bd_ram_mem0_reg[53][1]/P0001 , \wishbone_bd_ram_mem0_reg[53][2]/P0001 , \wishbone_bd_ram_mem0_reg[53][3]/P0001 , \wishbone_bd_ram_mem0_reg[53][4]/P0001 , \wishbone_bd_ram_mem0_reg[53][5]/P0001 , \wishbone_bd_ram_mem0_reg[53][6]/P0001 , \wishbone_bd_ram_mem0_reg[53][7]/P0001 , \wishbone_bd_ram_mem0_reg[54][0]/P0001 , \wishbone_bd_ram_mem0_reg[54][1]/P0001 , \wishbone_bd_ram_mem0_reg[54][2]/P0001 , \wishbone_bd_ram_mem0_reg[54][3]/P0001 , \wishbone_bd_ram_mem0_reg[54][4]/P0001 , \wishbone_bd_ram_mem0_reg[54][5]/P0001 , \wishbone_bd_ram_mem0_reg[54][6]/P0001 , \wishbone_bd_ram_mem0_reg[54][7]/P0001 , \wishbone_bd_ram_mem0_reg[55][0]/P0001 , \wishbone_bd_ram_mem0_reg[55][1]/P0001 , \wishbone_bd_ram_mem0_reg[55][2]/P0001 , \wishbone_bd_ram_mem0_reg[55][3]/P0001 , \wishbone_bd_ram_mem0_reg[55][4]/P0001 , \wishbone_bd_ram_mem0_reg[55][5]/P0001 , \wishbone_bd_ram_mem0_reg[55][6]/P0001 , \wishbone_bd_ram_mem0_reg[55][7]/P0001 , \wishbone_bd_ram_mem0_reg[56][0]/P0001 , \wishbone_bd_ram_mem0_reg[56][1]/P0001 , \wishbone_bd_ram_mem0_reg[56][2]/P0001 , \wishbone_bd_ram_mem0_reg[56][3]/P0001 , \wishbone_bd_ram_mem0_reg[56][4]/P0001 , \wishbone_bd_ram_mem0_reg[56][5]/P0001 , \wishbone_bd_ram_mem0_reg[56][6]/P0001 , \wishbone_bd_ram_mem0_reg[56][7]/P0001 , \wishbone_bd_ram_mem0_reg[57][0]/P0001 , \wishbone_bd_ram_mem0_reg[57][1]/P0001 , \wishbone_bd_ram_mem0_reg[57][2]/P0001 , \wishbone_bd_ram_mem0_reg[57][3]/P0001 , \wishbone_bd_ram_mem0_reg[57][4]/P0001 , \wishbone_bd_ram_mem0_reg[57][5]/P0001 , \wishbone_bd_ram_mem0_reg[57][6]/P0001 , \wishbone_bd_ram_mem0_reg[57][7]/P0001 , \wishbone_bd_ram_mem0_reg[58][0]/P0001 , \wishbone_bd_ram_mem0_reg[58][1]/P0001 , \wishbone_bd_ram_mem0_reg[58][2]/P0001 , \wishbone_bd_ram_mem0_reg[58][3]/P0001 , \wishbone_bd_ram_mem0_reg[58][4]/P0001 , \wishbone_bd_ram_mem0_reg[58][5]/P0001 , \wishbone_bd_ram_mem0_reg[58][6]/P0001 , \wishbone_bd_ram_mem0_reg[58][7]/P0001 , \wishbone_bd_ram_mem0_reg[59][0]/P0001 , \wishbone_bd_ram_mem0_reg[59][1]/P0001 , \wishbone_bd_ram_mem0_reg[59][2]/P0001 , \wishbone_bd_ram_mem0_reg[59][3]/P0001 , \wishbone_bd_ram_mem0_reg[59][4]/P0001 , \wishbone_bd_ram_mem0_reg[59][5]/P0001 , \wishbone_bd_ram_mem0_reg[59][6]/P0001 , \wishbone_bd_ram_mem0_reg[59][7]/P0001 , \wishbone_bd_ram_mem0_reg[5][0]/P0001 , \wishbone_bd_ram_mem0_reg[5][1]/P0001 , \wishbone_bd_ram_mem0_reg[5][2]/P0001 , \wishbone_bd_ram_mem0_reg[5][3]/P0001 , \wishbone_bd_ram_mem0_reg[5][4]/P0001 , \wishbone_bd_ram_mem0_reg[5][5]/P0001 , \wishbone_bd_ram_mem0_reg[5][6]/P0001 , \wishbone_bd_ram_mem0_reg[5][7]/P0001 , \wishbone_bd_ram_mem0_reg[60][0]/P0001 , \wishbone_bd_ram_mem0_reg[60][1]/P0001 , \wishbone_bd_ram_mem0_reg[60][2]/P0001 , \wishbone_bd_ram_mem0_reg[60][3]/P0001 , \wishbone_bd_ram_mem0_reg[60][4]/P0001 , \wishbone_bd_ram_mem0_reg[60][5]/P0001 , \wishbone_bd_ram_mem0_reg[60][6]/P0001 , \wishbone_bd_ram_mem0_reg[60][7]/P0001 , \wishbone_bd_ram_mem0_reg[61][0]/P0001 , \wishbone_bd_ram_mem0_reg[61][1]/P0001 , \wishbone_bd_ram_mem0_reg[61][2]/P0001 , \wishbone_bd_ram_mem0_reg[61][3]/P0001 , \wishbone_bd_ram_mem0_reg[61][4]/P0001 , \wishbone_bd_ram_mem0_reg[61][5]/P0001 , \wishbone_bd_ram_mem0_reg[61][6]/P0001 , \wishbone_bd_ram_mem0_reg[61][7]/P0001 , \wishbone_bd_ram_mem0_reg[62][0]/P0001 , \wishbone_bd_ram_mem0_reg[62][1]/P0001 , \wishbone_bd_ram_mem0_reg[62][2]/P0001 , \wishbone_bd_ram_mem0_reg[62][3]/P0001 , \wishbone_bd_ram_mem0_reg[62][4]/P0001 , \wishbone_bd_ram_mem0_reg[62][5]/P0001 , \wishbone_bd_ram_mem0_reg[62][6]/P0001 , \wishbone_bd_ram_mem0_reg[62][7]/P0001 , \wishbone_bd_ram_mem0_reg[63][0]/P0001 , \wishbone_bd_ram_mem0_reg[63][1]/P0001 , \wishbone_bd_ram_mem0_reg[63][2]/P0001 , \wishbone_bd_ram_mem0_reg[63][3]/P0001 , \wishbone_bd_ram_mem0_reg[63][4]/P0001 , \wishbone_bd_ram_mem0_reg[63][5]/P0001 , \wishbone_bd_ram_mem0_reg[63][6]/P0001 , \wishbone_bd_ram_mem0_reg[63][7]/P0001 , \wishbone_bd_ram_mem0_reg[64][0]/P0001 , \wishbone_bd_ram_mem0_reg[64][1]/P0001 , \wishbone_bd_ram_mem0_reg[64][2]/P0001 , \wishbone_bd_ram_mem0_reg[64][3]/P0001 , \wishbone_bd_ram_mem0_reg[64][4]/P0001 , \wishbone_bd_ram_mem0_reg[64][5]/P0001 , \wishbone_bd_ram_mem0_reg[64][6]/P0001 , \wishbone_bd_ram_mem0_reg[64][7]/P0001 , \wishbone_bd_ram_mem0_reg[65][0]/P0001 , \wishbone_bd_ram_mem0_reg[65][1]/P0001 , \wishbone_bd_ram_mem0_reg[65][2]/P0001 , \wishbone_bd_ram_mem0_reg[65][3]/P0001 , \wishbone_bd_ram_mem0_reg[65][4]/P0001 , \wishbone_bd_ram_mem0_reg[65][5]/P0001 , \wishbone_bd_ram_mem0_reg[65][6]/P0001 , \wishbone_bd_ram_mem0_reg[65][7]/P0001 , \wishbone_bd_ram_mem0_reg[66][0]/P0001 , \wishbone_bd_ram_mem0_reg[66][1]/P0001 , \wishbone_bd_ram_mem0_reg[66][2]/P0001 , \wishbone_bd_ram_mem0_reg[66][3]/P0001 , \wishbone_bd_ram_mem0_reg[66][4]/P0001 , \wishbone_bd_ram_mem0_reg[66][5]/P0001 , \wishbone_bd_ram_mem0_reg[66][6]/P0001 , \wishbone_bd_ram_mem0_reg[66][7]/P0001 , \wishbone_bd_ram_mem0_reg[67][0]/P0001 , \wishbone_bd_ram_mem0_reg[67][1]/P0001 , \wishbone_bd_ram_mem0_reg[67][2]/P0001 , \wishbone_bd_ram_mem0_reg[67][3]/P0001 , \wishbone_bd_ram_mem0_reg[67][4]/P0001 , \wishbone_bd_ram_mem0_reg[67][5]/P0001 , \wishbone_bd_ram_mem0_reg[67][6]/P0001 , \wishbone_bd_ram_mem0_reg[67][7]/P0001 , \wishbone_bd_ram_mem0_reg[68][0]/P0001 , \wishbone_bd_ram_mem0_reg[68][1]/P0001 , \wishbone_bd_ram_mem0_reg[68][2]/P0001 , \wishbone_bd_ram_mem0_reg[68][3]/P0001 , \wishbone_bd_ram_mem0_reg[68][4]/P0001 , \wishbone_bd_ram_mem0_reg[68][5]/P0001 , \wishbone_bd_ram_mem0_reg[68][6]/P0001 , \wishbone_bd_ram_mem0_reg[68][7]/P0001 , \wishbone_bd_ram_mem0_reg[69][0]/P0001 , \wishbone_bd_ram_mem0_reg[69][1]/P0001 , \wishbone_bd_ram_mem0_reg[69][2]/P0001 , \wishbone_bd_ram_mem0_reg[69][3]/P0001 , \wishbone_bd_ram_mem0_reg[69][4]/P0001 , \wishbone_bd_ram_mem0_reg[69][5]/P0001 , \wishbone_bd_ram_mem0_reg[69][6]/P0001 , \wishbone_bd_ram_mem0_reg[69][7]/P0001 , \wishbone_bd_ram_mem0_reg[6][0]/P0001 , \wishbone_bd_ram_mem0_reg[6][1]/P0001 , \wishbone_bd_ram_mem0_reg[6][2]/P0001 , \wishbone_bd_ram_mem0_reg[6][3]/P0001 , \wishbone_bd_ram_mem0_reg[6][4]/P0001 , \wishbone_bd_ram_mem0_reg[6][5]/P0001 , \wishbone_bd_ram_mem0_reg[6][6]/P0001 , \wishbone_bd_ram_mem0_reg[6][7]/P0001 , \wishbone_bd_ram_mem0_reg[70][0]/P0001 , \wishbone_bd_ram_mem0_reg[70][1]/P0001 , \wishbone_bd_ram_mem0_reg[70][2]/P0001 , \wishbone_bd_ram_mem0_reg[70][3]/P0001 , \wishbone_bd_ram_mem0_reg[70][4]/P0001 , \wishbone_bd_ram_mem0_reg[70][5]/P0001 , \wishbone_bd_ram_mem0_reg[70][6]/P0001 , \wishbone_bd_ram_mem0_reg[70][7]/P0001 , \wishbone_bd_ram_mem0_reg[71][0]/P0001 , \wishbone_bd_ram_mem0_reg[71][1]/P0001 , \wishbone_bd_ram_mem0_reg[71][2]/P0001 , \wishbone_bd_ram_mem0_reg[71][3]/P0001 , \wishbone_bd_ram_mem0_reg[71][4]/P0001 , \wishbone_bd_ram_mem0_reg[71][5]/P0001 , \wishbone_bd_ram_mem0_reg[71][6]/P0001 , \wishbone_bd_ram_mem0_reg[71][7]/P0001 , \wishbone_bd_ram_mem0_reg[72][0]/P0001 , \wishbone_bd_ram_mem0_reg[72][1]/P0001 , \wishbone_bd_ram_mem0_reg[72][2]/P0001 , \wishbone_bd_ram_mem0_reg[72][3]/P0001 , \wishbone_bd_ram_mem0_reg[72][4]/P0001 , \wishbone_bd_ram_mem0_reg[72][5]/P0001 , \wishbone_bd_ram_mem0_reg[72][6]/P0001 , \wishbone_bd_ram_mem0_reg[72][7]/P0001 , \wishbone_bd_ram_mem0_reg[73][0]/P0001 , \wishbone_bd_ram_mem0_reg[73][1]/P0001 , \wishbone_bd_ram_mem0_reg[73][2]/P0001 , \wishbone_bd_ram_mem0_reg[73][3]/P0001 , \wishbone_bd_ram_mem0_reg[73][4]/P0001 , \wishbone_bd_ram_mem0_reg[73][5]/P0001 , \wishbone_bd_ram_mem0_reg[73][6]/P0001 , \wishbone_bd_ram_mem0_reg[73][7]/P0001 , \wishbone_bd_ram_mem0_reg[74][0]/P0001 , \wishbone_bd_ram_mem0_reg[74][1]/P0001 , \wishbone_bd_ram_mem0_reg[74][2]/P0001 , \wishbone_bd_ram_mem0_reg[74][3]/P0001 , \wishbone_bd_ram_mem0_reg[74][4]/P0001 , \wishbone_bd_ram_mem0_reg[74][5]/P0001 , \wishbone_bd_ram_mem0_reg[74][6]/P0001 , \wishbone_bd_ram_mem0_reg[74][7]/P0001 , \wishbone_bd_ram_mem0_reg[75][0]/P0001 , \wishbone_bd_ram_mem0_reg[75][1]/P0001 , \wishbone_bd_ram_mem0_reg[75][2]/P0001 , \wishbone_bd_ram_mem0_reg[75][3]/P0001 , \wishbone_bd_ram_mem0_reg[75][4]/P0001 , \wishbone_bd_ram_mem0_reg[75][5]/P0001 , \wishbone_bd_ram_mem0_reg[75][6]/P0001 , \wishbone_bd_ram_mem0_reg[75][7]/P0001 , \wishbone_bd_ram_mem0_reg[76][0]/P0001 , \wishbone_bd_ram_mem0_reg[76][1]/P0001 , \wishbone_bd_ram_mem0_reg[76][2]/P0001 , \wishbone_bd_ram_mem0_reg[76][3]/P0001 , \wishbone_bd_ram_mem0_reg[76][4]/P0001 , \wishbone_bd_ram_mem0_reg[76][5]/P0001 , \wishbone_bd_ram_mem0_reg[76][6]/P0001 , \wishbone_bd_ram_mem0_reg[76][7]/P0001 , \wishbone_bd_ram_mem0_reg[77][0]/P0001 , \wishbone_bd_ram_mem0_reg[77][1]/P0001 , \wishbone_bd_ram_mem0_reg[77][2]/P0001 , \wishbone_bd_ram_mem0_reg[77][3]/P0001 , \wishbone_bd_ram_mem0_reg[77][4]/P0001 , \wishbone_bd_ram_mem0_reg[77][5]/P0001 , \wishbone_bd_ram_mem0_reg[77][6]/P0001 , \wishbone_bd_ram_mem0_reg[77][7]/P0001 , \wishbone_bd_ram_mem0_reg[78][0]/P0001 , \wishbone_bd_ram_mem0_reg[78][1]/P0001 , \wishbone_bd_ram_mem0_reg[78][2]/P0001 , \wishbone_bd_ram_mem0_reg[78][3]/P0001 , \wishbone_bd_ram_mem0_reg[78][4]/P0001 , \wishbone_bd_ram_mem0_reg[78][5]/P0001 , \wishbone_bd_ram_mem0_reg[78][6]/P0001 , \wishbone_bd_ram_mem0_reg[78][7]/P0001 , \wishbone_bd_ram_mem0_reg[79][0]/P0001 , \wishbone_bd_ram_mem0_reg[79][1]/P0001 , \wishbone_bd_ram_mem0_reg[79][2]/P0001 , \wishbone_bd_ram_mem0_reg[79][3]/P0001 , \wishbone_bd_ram_mem0_reg[79][4]/P0001 , \wishbone_bd_ram_mem0_reg[79][5]/P0001 , \wishbone_bd_ram_mem0_reg[79][6]/P0001 , \wishbone_bd_ram_mem0_reg[79][7]/P0001 , \wishbone_bd_ram_mem0_reg[7][0]/P0001 , \wishbone_bd_ram_mem0_reg[7][1]/P0001 , \wishbone_bd_ram_mem0_reg[7][2]/P0001 , \wishbone_bd_ram_mem0_reg[7][3]/P0001 , \wishbone_bd_ram_mem0_reg[7][4]/P0001 , \wishbone_bd_ram_mem0_reg[7][5]/P0001 , \wishbone_bd_ram_mem0_reg[7][6]/P0001 , \wishbone_bd_ram_mem0_reg[7][7]/P0001 , \wishbone_bd_ram_mem0_reg[80][0]/P0001 , \wishbone_bd_ram_mem0_reg[80][1]/P0001 , \wishbone_bd_ram_mem0_reg[80][2]/P0001 , \wishbone_bd_ram_mem0_reg[80][3]/P0001 , \wishbone_bd_ram_mem0_reg[80][4]/P0001 , \wishbone_bd_ram_mem0_reg[80][5]/P0001 , \wishbone_bd_ram_mem0_reg[80][6]/P0001 , \wishbone_bd_ram_mem0_reg[80][7]/P0001 , \wishbone_bd_ram_mem0_reg[81][0]/P0001 , \wishbone_bd_ram_mem0_reg[81][1]/P0001 , \wishbone_bd_ram_mem0_reg[81][2]/P0001 , \wishbone_bd_ram_mem0_reg[81][3]/P0001 , \wishbone_bd_ram_mem0_reg[81][4]/P0001 , \wishbone_bd_ram_mem0_reg[81][5]/P0001 , \wishbone_bd_ram_mem0_reg[81][6]/P0001 , \wishbone_bd_ram_mem0_reg[81][7]/P0001 , \wishbone_bd_ram_mem0_reg[82][0]/P0001 , \wishbone_bd_ram_mem0_reg[82][1]/P0001 , \wishbone_bd_ram_mem0_reg[82][2]/P0001 , \wishbone_bd_ram_mem0_reg[82][3]/P0001 , \wishbone_bd_ram_mem0_reg[82][4]/P0001 , \wishbone_bd_ram_mem0_reg[82][5]/P0001 , \wishbone_bd_ram_mem0_reg[82][6]/P0001 , \wishbone_bd_ram_mem0_reg[82][7]/P0001 , \wishbone_bd_ram_mem0_reg[83][0]/P0001 , \wishbone_bd_ram_mem0_reg[83][1]/P0001 , \wishbone_bd_ram_mem0_reg[83][2]/P0001 , \wishbone_bd_ram_mem0_reg[83][3]/P0001 , \wishbone_bd_ram_mem0_reg[83][4]/P0001 , \wishbone_bd_ram_mem0_reg[83][5]/P0001 , \wishbone_bd_ram_mem0_reg[83][6]/P0001 , \wishbone_bd_ram_mem0_reg[83][7]/P0001 , \wishbone_bd_ram_mem0_reg[84][0]/P0001 , \wishbone_bd_ram_mem0_reg[84][1]/P0001 , \wishbone_bd_ram_mem0_reg[84][2]/P0001 , \wishbone_bd_ram_mem0_reg[84][3]/P0001 , \wishbone_bd_ram_mem0_reg[84][4]/P0001 , \wishbone_bd_ram_mem0_reg[84][5]/P0001 , \wishbone_bd_ram_mem0_reg[84][6]/P0001 , \wishbone_bd_ram_mem0_reg[84][7]/P0001 , \wishbone_bd_ram_mem0_reg[85][0]/P0001 , \wishbone_bd_ram_mem0_reg[85][1]/P0001 , \wishbone_bd_ram_mem0_reg[85][2]/P0001 , \wishbone_bd_ram_mem0_reg[85][3]/P0001 , \wishbone_bd_ram_mem0_reg[85][4]/P0001 , \wishbone_bd_ram_mem0_reg[85][5]/P0001 , \wishbone_bd_ram_mem0_reg[85][6]/P0001 , \wishbone_bd_ram_mem0_reg[85][7]/P0001 , \wishbone_bd_ram_mem0_reg[86][0]/P0001 , \wishbone_bd_ram_mem0_reg[86][1]/P0001 , \wishbone_bd_ram_mem0_reg[86][2]/P0001 , \wishbone_bd_ram_mem0_reg[86][3]/P0001 , \wishbone_bd_ram_mem0_reg[86][4]/P0001 , \wishbone_bd_ram_mem0_reg[86][5]/P0001 , \wishbone_bd_ram_mem0_reg[86][6]/P0001 , \wishbone_bd_ram_mem0_reg[86][7]/P0001 , \wishbone_bd_ram_mem0_reg[87][0]/P0001 , \wishbone_bd_ram_mem0_reg[87][1]/P0001 , \wishbone_bd_ram_mem0_reg[87][2]/P0001 , \wishbone_bd_ram_mem0_reg[87][3]/P0001 , \wishbone_bd_ram_mem0_reg[87][4]/P0001 , \wishbone_bd_ram_mem0_reg[87][5]/P0001 , \wishbone_bd_ram_mem0_reg[87][6]/P0001 , \wishbone_bd_ram_mem0_reg[87][7]/P0001 , \wishbone_bd_ram_mem0_reg[88][0]/P0001 , \wishbone_bd_ram_mem0_reg[88][1]/P0001 , \wishbone_bd_ram_mem0_reg[88][2]/P0001 , \wishbone_bd_ram_mem0_reg[88][3]/P0001 , \wishbone_bd_ram_mem0_reg[88][4]/P0001 , \wishbone_bd_ram_mem0_reg[88][5]/P0001 , \wishbone_bd_ram_mem0_reg[88][6]/P0001 , \wishbone_bd_ram_mem0_reg[88][7]/P0001 , \wishbone_bd_ram_mem0_reg[89][0]/P0001 , \wishbone_bd_ram_mem0_reg[89][1]/P0001 , \wishbone_bd_ram_mem0_reg[89][2]/P0001 , \wishbone_bd_ram_mem0_reg[89][3]/P0001 , \wishbone_bd_ram_mem0_reg[89][4]/P0001 , \wishbone_bd_ram_mem0_reg[89][5]/P0001 , \wishbone_bd_ram_mem0_reg[89][6]/P0001 , \wishbone_bd_ram_mem0_reg[89][7]/P0001 , \wishbone_bd_ram_mem0_reg[8][0]/P0001 , \wishbone_bd_ram_mem0_reg[8][1]/P0001 , \wishbone_bd_ram_mem0_reg[8][2]/P0001 , \wishbone_bd_ram_mem0_reg[8][3]/P0001 , \wishbone_bd_ram_mem0_reg[8][4]/P0001 , \wishbone_bd_ram_mem0_reg[8][5]/P0001 , \wishbone_bd_ram_mem0_reg[8][6]/P0001 , \wishbone_bd_ram_mem0_reg[8][7]/P0001 , \wishbone_bd_ram_mem0_reg[90][0]/P0001 , \wishbone_bd_ram_mem0_reg[90][1]/P0001 , \wishbone_bd_ram_mem0_reg[90][2]/P0001 , \wishbone_bd_ram_mem0_reg[90][3]/P0001 , \wishbone_bd_ram_mem0_reg[90][4]/P0001 , \wishbone_bd_ram_mem0_reg[90][5]/P0001 , \wishbone_bd_ram_mem0_reg[90][6]/P0001 , \wishbone_bd_ram_mem0_reg[90][7]/P0001 , \wishbone_bd_ram_mem0_reg[91][0]/P0001 , \wishbone_bd_ram_mem0_reg[91][1]/P0001 , \wishbone_bd_ram_mem0_reg[91][2]/P0001 , \wishbone_bd_ram_mem0_reg[91][3]/P0001 , \wishbone_bd_ram_mem0_reg[91][4]/P0001 , \wishbone_bd_ram_mem0_reg[91][5]/P0001 , \wishbone_bd_ram_mem0_reg[91][6]/P0001 , \wishbone_bd_ram_mem0_reg[91][7]/P0001 , \wishbone_bd_ram_mem0_reg[92][0]/P0001 , \wishbone_bd_ram_mem0_reg[92][1]/P0001 , \wishbone_bd_ram_mem0_reg[92][2]/P0001 , \wishbone_bd_ram_mem0_reg[92][3]/P0001 , \wishbone_bd_ram_mem0_reg[92][4]/P0001 , \wishbone_bd_ram_mem0_reg[92][5]/P0001 , \wishbone_bd_ram_mem0_reg[92][6]/P0001 , \wishbone_bd_ram_mem0_reg[92][7]/P0001 , \wishbone_bd_ram_mem0_reg[93][0]/P0001 , \wishbone_bd_ram_mem0_reg[93][1]/P0001 , \wishbone_bd_ram_mem0_reg[93][2]/P0001 , \wishbone_bd_ram_mem0_reg[93][3]/P0001 , \wishbone_bd_ram_mem0_reg[93][4]/P0001 , \wishbone_bd_ram_mem0_reg[93][5]/P0001 , \wishbone_bd_ram_mem0_reg[93][6]/P0001 , \wishbone_bd_ram_mem0_reg[93][7]/P0001 , \wishbone_bd_ram_mem0_reg[94][0]/P0001 , \wishbone_bd_ram_mem0_reg[94][1]/P0001 , \wishbone_bd_ram_mem0_reg[94][2]/P0001 , \wishbone_bd_ram_mem0_reg[94][3]/P0001 , \wishbone_bd_ram_mem0_reg[94][4]/P0001 , \wishbone_bd_ram_mem0_reg[94][5]/P0001 , \wishbone_bd_ram_mem0_reg[94][6]/P0001 , \wishbone_bd_ram_mem0_reg[94][7]/P0001 , \wishbone_bd_ram_mem0_reg[95][0]/P0001 , \wishbone_bd_ram_mem0_reg[95][1]/P0001 , \wishbone_bd_ram_mem0_reg[95][2]/P0001 , \wishbone_bd_ram_mem0_reg[95][3]/P0001 , \wishbone_bd_ram_mem0_reg[95][4]/P0001 , \wishbone_bd_ram_mem0_reg[95][5]/P0001 , \wishbone_bd_ram_mem0_reg[95][6]/P0001 , \wishbone_bd_ram_mem0_reg[95][7]/P0001 , \wishbone_bd_ram_mem0_reg[96][0]/P0001 , \wishbone_bd_ram_mem0_reg[96][1]/P0001 , \wishbone_bd_ram_mem0_reg[96][2]/P0001 , \wishbone_bd_ram_mem0_reg[96][3]/P0001 , \wishbone_bd_ram_mem0_reg[96][4]/P0001 , \wishbone_bd_ram_mem0_reg[96][5]/P0001 , \wishbone_bd_ram_mem0_reg[96][6]/P0001 , \wishbone_bd_ram_mem0_reg[96][7]/P0001 , \wishbone_bd_ram_mem0_reg[97][0]/P0001 , \wishbone_bd_ram_mem0_reg[97][1]/P0001 , \wishbone_bd_ram_mem0_reg[97][2]/P0001 , \wishbone_bd_ram_mem0_reg[97][3]/P0001 , \wishbone_bd_ram_mem0_reg[97][4]/P0001 , \wishbone_bd_ram_mem0_reg[97][5]/P0001 , \wishbone_bd_ram_mem0_reg[97][6]/P0001 , \wishbone_bd_ram_mem0_reg[97][7]/P0001 , \wishbone_bd_ram_mem0_reg[98][0]/P0001 , \wishbone_bd_ram_mem0_reg[98][1]/P0001 , \wishbone_bd_ram_mem0_reg[98][2]/P0001 , \wishbone_bd_ram_mem0_reg[98][3]/P0001 , \wishbone_bd_ram_mem0_reg[98][4]/P0001 , \wishbone_bd_ram_mem0_reg[98][5]/P0001 , \wishbone_bd_ram_mem0_reg[98][6]/P0001 , \wishbone_bd_ram_mem0_reg[98][7]/P0001 , \wishbone_bd_ram_mem0_reg[99][0]/P0001 , \wishbone_bd_ram_mem0_reg[99][1]/P0001 , \wishbone_bd_ram_mem0_reg[99][2]/P0001 , \wishbone_bd_ram_mem0_reg[99][3]/P0001 , \wishbone_bd_ram_mem0_reg[99][4]/P0001 , \wishbone_bd_ram_mem0_reg[99][5]/P0001 , \wishbone_bd_ram_mem0_reg[99][6]/P0001 , \wishbone_bd_ram_mem0_reg[99][7]/P0001 , \wishbone_bd_ram_mem0_reg[9][0]/P0001 , \wishbone_bd_ram_mem0_reg[9][1]/P0001 , \wishbone_bd_ram_mem0_reg[9][2]/P0001 , \wishbone_bd_ram_mem0_reg[9][3]/P0001 , \wishbone_bd_ram_mem0_reg[9][4]/P0001 , \wishbone_bd_ram_mem0_reg[9][5]/P0001 , \wishbone_bd_ram_mem0_reg[9][6]/P0001 , \wishbone_bd_ram_mem0_reg[9][7]/P0001 , \wishbone_bd_ram_mem1_reg[0][10]/P0001 , \wishbone_bd_ram_mem1_reg[0][11]/P0001 , \wishbone_bd_ram_mem1_reg[0][12]/P0001 , \wishbone_bd_ram_mem1_reg[0][13]/P0001 , \wishbone_bd_ram_mem1_reg[0][14]/P0001 , \wishbone_bd_ram_mem1_reg[0][15]/P0001 , \wishbone_bd_ram_mem1_reg[0][8]/P0001 , \wishbone_bd_ram_mem1_reg[0][9]/P0001 , \wishbone_bd_ram_mem1_reg[100][10]/P0001 , \wishbone_bd_ram_mem1_reg[100][11]/P0001 , \wishbone_bd_ram_mem1_reg[100][12]/P0001 , \wishbone_bd_ram_mem1_reg[100][13]/P0001 , \wishbone_bd_ram_mem1_reg[100][14]/P0001 , \wishbone_bd_ram_mem1_reg[100][15]/P0001 , \wishbone_bd_ram_mem1_reg[100][8]/P0001 , \wishbone_bd_ram_mem1_reg[100][9]/P0001 , \wishbone_bd_ram_mem1_reg[101][10]/P0001 , \wishbone_bd_ram_mem1_reg[101][11]/P0001 , \wishbone_bd_ram_mem1_reg[101][12]/P0001 , \wishbone_bd_ram_mem1_reg[101][13]/P0001 , \wishbone_bd_ram_mem1_reg[101][14]/P0001 , \wishbone_bd_ram_mem1_reg[101][15]/P0001 , \wishbone_bd_ram_mem1_reg[101][8]/P0001 , \wishbone_bd_ram_mem1_reg[101][9]/P0001 , \wishbone_bd_ram_mem1_reg[102][10]/P0001 , \wishbone_bd_ram_mem1_reg[102][11]/P0001 , \wishbone_bd_ram_mem1_reg[102][12]/P0001 , \wishbone_bd_ram_mem1_reg[102][13]/P0001 , \wishbone_bd_ram_mem1_reg[102][14]/P0001 , \wishbone_bd_ram_mem1_reg[102][15]/P0001 , \wishbone_bd_ram_mem1_reg[102][8]/P0001 , \wishbone_bd_ram_mem1_reg[102][9]/P0001 , \wishbone_bd_ram_mem1_reg[103][10]/P0001 , \wishbone_bd_ram_mem1_reg[103][11]/P0001 , \wishbone_bd_ram_mem1_reg[103][12]/P0001 , \wishbone_bd_ram_mem1_reg[103][13]/P0001 , \wishbone_bd_ram_mem1_reg[103][14]/P0001 , \wishbone_bd_ram_mem1_reg[103][15]/P0001 , \wishbone_bd_ram_mem1_reg[103][8]/P0001 , \wishbone_bd_ram_mem1_reg[103][9]/P0001 , \wishbone_bd_ram_mem1_reg[104][10]/P0001 , \wishbone_bd_ram_mem1_reg[104][11]/P0001 , \wishbone_bd_ram_mem1_reg[104][12]/P0001 , \wishbone_bd_ram_mem1_reg[104][13]/P0001 , \wishbone_bd_ram_mem1_reg[104][14]/P0001 , \wishbone_bd_ram_mem1_reg[104][15]/P0001 , \wishbone_bd_ram_mem1_reg[104][8]/P0001 , \wishbone_bd_ram_mem1_reg[104][9]/P0001 , \wishbone_bd_ram_mem1_reg[105][10]/P0001 , \wishbone_bd_ram_mem1_reg[105][11]/P0001 , \wishbone_bd_ram_mem1_reg[105][12]/P0001 , \wishbone_bd_ram_mem1_reg[105][13]/P0001 , \wishbone_bd_ram_mem1_reg[105][14]/P0001 , \wishbone_bd_ram_mem1_reg[105][15]/P0001 , \wishbone_bd_ram_mem1_reg[105][8]/P0001 , \wishbone_bd_ram_mem1_reg[105][9]/P0001 , \wishbone_bd_ram_mem1_reg[106][10]/P0001 , \wishbone_bd_ram_mem1_reg[106][11]/P0001 , \wishbone_bd_ram_mem1_reg[106][12]/P0001 , \wishbone_bd_ram_mem1_reg[106][13]/P0001 , \wishbone_bd_ram_mem1_reg[106][14]/P0001 , \wishbone_bd_ram_mem1_reg[106][15]/P0001 , \wishbone_bd_ram_mem1_reg[106][8]/P0001 , \wishbone_bd_ram_mem1_reg[106][9]/P0001 , \wishbone_bd_ram_mem1_reg[107][10]/P0001 , \wishbone_bd_ram_mem1_reg[107][11]/P0001 , \wishbone_bd_ram_mem1_reg[107][12]/P0001 , \wishbone_bd_ram_mem1_reg[107][13]/P0001 , \wishbone_bd_ram_mem1_reg[107][14]/P0001 , \wishbone_bd_ram_mem1_reg[107][15]/P0001 , \wishbone_bd_ram_mem1_reg[107][8]/P0001 , \wishbone_bd_ram_mem1_reg[107][9]/P0001 , \wishbone_bd_ram_mem1_reg[108][10]/P0001 , \wishbone_bd_ram_mem1_reg[108][11]/P0001 , \wishbone_bd_ram_mem1_reg[108][12]/P0001 , \wishbone_bd_ram_mem1_reg[108][13]/P0001 , \wishbone_bd_ram_mem1_reg[108][14]/P0001 , \wishbone_bd_ram_mem1_reg[108][15]/P0001 , \wishbone_bd_ram_mem1_reg[108][8]/P0001 , \wishbone_bd_ram_mem1_reg[108][9]/P0001 , \wishbone_bd_ram_mem1_reg[109][10]/P0001 , \wishbone_bd_ram_mem1_reg[109][11]/P0001 , \wishbone_bd_ram_mem1_reg[109][12]/P0001 , \wishbone_bd_ram_mem1_reg[109][13]/P0001 , \wishbone_bd_ram_mem1_reg[109][14]/P0001 , \wishbone_bd_ram_mem1_reg[109][15]/P0001 , \wishbone_bd_ram_mem1_reg[109][8]/P0001 , \wishbone_bd_ram_mem1_reg[109][9]/P0001 , \wishbone_bd_ram_mem1_reg[10][10]/P0001 , \wishbone_bd_ram_mem1_reg[10][11]/P0001 , \wishbone_bd_ram_mem1_reg[10][12]/P0001 , \wishbone_bd_ram_mem1_reg[10][13]/P0001 , \wishbone_bd_ram_mem1_reg[10][14]/P0001 , \wishbone_bd_ram_mem1_reg[10][15]/P0001 , \wishbone_bd_ram_mem1_reg[10][8]/P0001 , \wishbone_bd_ram_mem1_reg[10][9]/P0001 , \wishbone_bd_ram_mem1_reg[110][10]/P0001 , \wishbone_bd_ram_mem1_reg[110][11]/P0001 , \wishbone_bd_ram_mem1_reg[110][12]/P0001 , \wishbone_bd_ram_mem1_reg[110][13]/P0001 , \wishbone_bd_ram_mem1_reg[110][14]/P0001 , \wishbone_bd_ram_mem1_reg[110][15]/P0001 , \wishbone_bd_ram_mem1_reg[110][8]/P0001 , \wishbone_bd_ram_mem1_reg[110][9]/P0001 , \wishbone_bd_ram_mem1_reg[111][10]/P0001 , \wishbone_bd_ram_mem1_reg[111][11]/P0001 , \wishbone_bd_ram_mem1_reg[111][12]/P0001 , \wishbone_bd_ram_mem1_reg[111][13]/P0001 , \wishbone_bd_ram_mem1_reg[111][14]/P0001 , \wishbone_bd_ram_mem1_reg[111][15]/P0001 , \wishbone_bd_ram_mem1_reg[111][8]/P0001 , \wishbone_bd_ram_mem1_reg[111][9]/P0001 , \wishbone_bd_ram_mem1_reg[112][10]/P0001 , \wishbone_bd_ram_mem1_reg[112][11]/P0001 , \wishbone_bd_ram_mem1_reg[112][12]/P0001 , \wishbone_bd_ram_mem1_reg[112][13]/P0001 , \wishbone_bd_ram_mem1_reg[112][14]/P0001 , \wishbone_bd_ram_mem1_reg[112][15]/P0001 , \wishbone_bd_ram_mem1_reg[112][8]/P0001 , \wishbone_bd_ram_mem1_reg[112][9]/P0001 , \wishbone_bd_ram_mem1_reg[113][10]/P0001 , \wishbone_bd_ram_mem1_reg[113][11]/P0001 , \wishbone_bd_ram_mem1_reg[113][12]/P0001 , \wishbone_bd_ram_mem1_reg[113][13]/P0001 , \wishbone_bd_ram_mem1_reg[113][14]/P0001 , \wishbone_bd_ram_mem1_reg[113][15]/P0001 , \wishbone_bd_ram_mem1_reg[113][8]/P0001 , \wishbone_bd_ram_mem1_reg[113][9]/P0001 , \wishbone_bd_ram_mem1_reg[114][10]/P0001 , \wishbone_bd_ram_mem1_reg[114][11]/P0001 , \wishbone_bd_ram_mem1_reg[114][12]/P0001 , \wishbone_bd_ram_mem1_reg[114][13]/P0001 , \wishbone_bd_ram_mem1_reg[114][14]/P0001 , \wishbone_bd_ram_mem1_reg[114][15]/P0001 , \wishbone_bd_ram_mem1_reg[114][8]/P0001 , \wishbone_bd_ram_mem1_reg[114][9]/P0001 , \wishbone_bd_ram_mem1_reg[115][10]/P0001 , \wishbone_bd_ram_mem1_reg[115][11]/P0001 , \wishbone_bd_ram_mem1_reg[115][12]/P0001 , \wishbone_bd_ram_mem1_reg[115][13]/P0001 , \wishbone_bd_ram_mem1_reg[115][14]/P0001 , \wishbone_bd_ram_mem1_reg[115][15]/P0001 , \wishbone_bd_ram_mem1_reg[115][8]/P0001 , \wishbone_bd_ram_mem1_reg[115][9]/P0001 , \wishbone_bd_ram_mem1_reg[116][10]/P0001 , \wishbone_bd_ram_mem1_reg[116][11]/P0001 , \wishbone_bd_ram_mem1_reg[116][12]/P0001 , \wishbone_bd_ram_mem1_reg[116][13]/P0001 , \wishbone_bd_ram_mem1_reg[116][14]/P0001 , \wishbone_bd_ram_mem1_reg[116][15]/P0001 , \wishbone_bd_ram_mem1_reg[116][8]/P0001 , \wishbone_bd_ram_mem1_reg[116][9]/P0001 , \wishbone_bd_ram_mem1_reg[117][10]/P0001 , \wishbone_bd_ram_mem1_reg[117][11]/P0001 , \wishbone_bd_ram_mem1_reg[117][12]/P0001 , \wishbone_bd_ram_mem1_reg[117][13]/P0001 , \wishbone_bd_ram_mem1_reg[117][14]/P0001 , \wishbone_bd_ram_mem1_reg[117][15]/P0001 , \wishbone_bd_ram_mem1_reg[117][8]/P0001 , \wishbone_bd_ram_mem1_reg[117][9]/P0001 , \wishbone_bd_ram_mem1_reg[118][10]/P0001 , \wishbone_bd_ram_mem1_reg[118][11]/P0001 , \wishbone_bd_ram_mem1_reg[118][12]/P0001 , \wishbone_bd_ram_mem1_reg[118][13]/P0001 , \wishbone_bd_ram_mem1_reg[118][14]/P0001 , \wishbone_bd_ram_mem1_reg[118][15]/P0001 , \wishbone_bd_ram_mem1_reg[118][8]/P0001 , \wishbone_bd_ram_mem1_reg[118][9]/P0001 , \wishbone_bd_ram_mem1_reg[119][10]/P0001 , \wishbone_bd_ram_mem1_reg[119][11]/P0001 , \wishbone_bd_ram_mem1_reg[119][12]/P0001 , \wishbone_bd_ram_mem1_reg[119][13]/P0001 , \wishbone_bd_ram_mem1_reg[119][14]/P0001 , \wishbone_bd_ram_mem1_reg[119][15]/P0001 , \wishbone_bd_ram_mem1_reg[119][8]/P0001 , \wishbone_bd_ram_mem1_reg[119][9]/P0001 , \wishbone_bd_ram_mem1_reg[11][10]/P0001 , \wishbone_bd_ram_mem1_reg[11][11]/P0001 , \wishbone_bd_ram_mem1_reg[11][12]/P0001 , \wishbone_bd_ram_mem1_reg[11][13]/P0001 , \wishbone_bd_ram_mem1_reg[11][14]/P0001 , \wishbone_bd_ram_mem1_reg[11][15]/P0001 , \wishbone_bd_ram_mem1_reg[11][8]/P0001 , \wishbone_bd_ram_mem1_reg[11][9]/P0001 , \wishbone_bd_ram_mem1_reg[120][10]/P0001 , \wishbone_bd_ram_mem1_reg[120][11]/P0001 , \wishbone_bd_ram_mem1_reg[120][12]/P0001 , \wishbone_bd_ram_mem1_reg[120][13]/P0001 , \wishbone_bd_ram_mem1_reg[120][14]/P0001 , \wishbone_bd_ram_mem1_reg[120][15]/P0001 , \wishbone_bd_ram_mem1_reg[120][8]/P0001 , \wishbone_bd_ram_mem1_reg[120][9]/P0001 , \wishbone_bd_ram_mem1_reg[121][10]/P0001 , \wishbone_bd_ram_mem1_reg[121][11]/P0001 , \wishbone_bd_ram_mem1_reg[121][12]/P0001 , \wishbone_bd_ram_mem1_reg[121][13]/P0001 , \wishbone_bd_ram_mem1_reg[121][14]/P0001 , \wishbone_bd_ram_mem1_reg[121][15]/P0001 , \wishbone_bd_ram_mem1_reg[121][8]/P0001 , \wishbone_bd_ram_mem1_reg[121][9]/P0001 , \wishbone_bd_ram_mem1_reg[122][10]/P0001 , \wishbone_bd_ram_mem1_reg[122][11]/P0001 , \wishbone_bd_ram_mem1_reg[122][12]/P0001 , \wishbone_bd_ram_mem1_reg[122][13]/P0001 , \wishbone_bd_ram_mem1_reg[122][14]/P0001 , \wishbone_bd_ram_mem1_reg[122][15]/P0001 , \wishbone_bd_ram_mem1_reg[122][8]/P0001 , \wishbone_bd_ram_mem1_reg[122][9]/P0001 , \wishbone_bd_ram_mem1_reg[123][10]/P0001 , \wishbone_bd_ram_mem1_reg[123][11]/P0001 , \wishbone_bd_ram_mem1_reg[123][12]/P0001 , \wishbone_bd_ram_mem1_reg[123][13]/P0001 , \wishbone_bd_ram_mem1_reg[123][14]/P0001 , \wishbone_bd_ram_mem1_reg[123][15]/P0001 , \wishbone_bd_ram_mem1_reg[123][8]/P0001 , \wishbone_bd_ram_mem1_reg[123][9]/P0001 , \wishbone_bd_ram_mem1_reg[124][10]/P0001 , \wishbone_bd_ram_mem1_reg[124][11]/P0001 , \wishbone_bd_ram_mem1_reg[124][12]/P0001 , \wishbone_bd_ram_mem1_reg[124][13]/P0001 , \wishbone_bd_ram_mem1_reg[124][14]/P0001 , \wishbone_bd_ram_mem1_reg[124][15]/P0001 , \wishbone_bd_ram_mem1_reg[124][8]/P0001 , \wishbone_bd_ram_mem1_reg[124][9]/P0001 , \wishbone_bd_ram_mem1_reg[125][10]/P0001 , \wishbone_bd_ram_mem1_reg[125][11]/P0001 , \wishbone_bd_ram_mem1_reg[125][12]/P0001 , \wishbone_bd_ram_mem1_reg[125][13]/P0001 , \wishbone_bd_ram_mem1_reg[125][14]/P0001 , \wishbone_bd_ram_mem1_reg[125][15]/P0001 , \wishbone_bd_ram_mem1_reg[125][8]/P0001 , \wishbone_bd_ram_mem1_reg[125][9]/P0001 , \wishbone_bd_ram_mem1_reg[126][10]/P0001 , \wishbone_bd_ram_mem1_reg[126][11]/P0001 , \wishbone_bd_ram_mem1_reg[126][12]/P0001 , \wishbone_bd_ram_mem1_reg[126][13]/P0001 , \wishbone_bd_ram_mem1_reg[126][14]/P0001 , \wishbone_bd_ram_mem1_reg[126][15]/P0001 , \wishbone_bd_ram_mem1_reg[126][8]/P0001 , \wishbone_bd_ram_mem1_reg[126][9]/P0001 , \wishbone_bd_ram_mem1_reg[127][10]/P0001 , \wishbone_bd_ram_mem1_reg[127][11]/P0001 , \wishbone_bd_ram_mem1_reg[127][12]/P0001 , \wishbone_bd_ram_mem1_reg[127][13]/P0001 , \wishbone_bd_ram_mem1_reg[127][14]/P0001 , \wishbone_bd_ram_mem1_reg[127][15]/P0001 , \wishbone_bd_ram_mem1_reg[127][8]/P0001 , \wishbone_bd_ram_mem1_reg[127][9]/P0001 , \wishbone_bd_ram_mem1_reg[128][10]/P0001 , \wishbone_bd_ram_mem1_reg[128][11]/P0001 , \wishbone_bd_ram_mem1_reg[128][12]/P0001 , \wishbone_bd_ram_mem1_reg[128][13]/P0001 , \wishbone_bd_ram_mem1_reg[128][14]/P0001 , \wishbone_bd_ram_mem1_reg[128][15]/P0001 , \wishbone_bd_ram_mem1_reg[128][8]/P0001 , \wishbone_bd_ram_mem1_reg[128][9]/P0001 , \wishbone_bd_ram_mem1_reg[129][10]/P0001 , \wishbone_bd_ram_mem1_reg[129][11]/P0001 , \wishbone_bd_ram_mem1_reg[129][12]/P0001 , \wishbone_bd_ram_mem1_reg[129][13]/P0001 , \wishbone_bd_ram_mem1_reg[129][14]/P0001 , \wishbone_bd_ram_mem1_reg[129][15]/P0001 , \wishbone_bd_ram_mem1_reg[129][8]/P0001 , \wishbone_bd_ram_mem1_reg[129][9]/P0001 , \wishbone_bd_ram_mem1_reg[12][10]/P0001 , \wishbone_bd_ram_mem1_reg[12][11]/P0001 , \wishbone_bd_ram_mem1_reg[12][12]/P0001 , \wishbone_bd_ram_mem1_reg[12][13]/P0001 , \wishbone_bd_ram_mem1_reg[12][14]/P0001 , \wishbone_bd_ram_mem1_reg[12][15]/P0001 , \wishbone_bd_ram_mem1_reg[12][8]/P0001 , \wishbone_bd_ram_mem1_reg[12][9]/P0001 , \wishbone_bd_ram_mem1_reg[130][10]/P0001 , \wishbone_bd_ram_mem1_reg[130][11]/P0001 , \wishbone_bd_ram_mem1_reg[130][12]/P0001 , \wishbone_bd_ram_mem1_reg[130][13]/P0001 , \wishbone_bd_ram_mem1_reg[130][14]/P0001 , \wishbone_bd_ram_mem1_reg[130][15]/P0001 , \wishbone_bd_ram_mem1_reg[130][8]/P0001 , \wishbone_bd_ram_mem1_reg[130][9]/P0001 , \wishbone_bd_ram_mem1_reg[131][10]/P0001 , \wishbone_bd_ram_mem1_reg[131][11]/P0001 , \wishbone_bd_ram_mem1_reg[131][12]/P0001 , \wishbone_bd_ram_mem1_reg[131][13]/P0001 , \wishbone_bd_ram_mem1_reg[131][14]/P0001 , \wishbone_bd_ram_mem1_reg[131][15]/P0001 , \wishbone_bd_ram_mem1_reg[131][8]/P0001 , \wishbone_bd_ram_mem1_reg[131][9]/P0001 , \wishbone_bd_ram_mem1_reg[132][10]/P0001 , \wishbone_bd_ram_mem1_reg[132][11]/P0001 , \wishbone_bd_ram_mem1_reg[132][12]/P0001 , \wishbone_bd_ram_mem1_reg[132][13]/P0001 , \wishbone_bd_ram_mem1_reg[132][14]/P0001 , \wishbone_bd_ram_mem1_reg[132][15]/P0001 , \wishbone_bd_ram_mem1_reg[132][8]/P0001 , \wishbone_bd_ram_mem1_reg[132][9]/P0001 , \wishbone_bd_ram_mem1_reg[133][10]/P0001 , \wishbone_bd_ram_mem1_reg[133][11]/P0001 , \wishbone_bd_ram_mem1_reg[133][12]/P0001 , \wishbone_bd_ram_mem1_reg[133][13]/P0001 , \wishbone_bd_ram_mem1_reg[133][14]/P0001 , \wishbone_bd_ram_mem1_reg[133][15]/P0001 , \wishbone_bd_ram_mem1_reg[133][8]/P0001 , \wishbone_bd_ram_mem1_reg[133][9]/P0001 , \wishbone_bd_ram_mem1_reg[134][10]/P0001 , \wishbone_bd_ram_mem1_reg[134][11]/P0001 , \wishbone_bd_ram_mem1_reg[134][12]/P0001 , \wishbone_bd_ram_mem1_reg[134][13]/P0001 , \wishbone_bd_ram_mem1_reg[134][14]/P0001 , \wishbone_bd_ram_mem1_reg[134][15]/P0001 , \wishbone_bd_ram_mem1_reg[134][8]/P0001 , \wishbone_bd_ram_mem1_reg[134][9]/P0001 , \wishbone_bd_ram_mem1_reg[135][10]/P0001 , \wishbone_bd_ram_mem1_reg[135][11]/P0001 , \wishbone_bd_ram_mem1_reg[135][12]/P0001 , \wishbone_bd_ram_mem1_reg[135][13]/P0001 , \wishbone_bd_ram_mem1_reg[135][14]/P0001 , \wishbone_bd_ram_mem1_reg[135][15]/P0001 , \wishbone_bd_ram_mem1_reg[135][8]/P0001 , \wishbone_bd_ram_mem1_reg[135][9]/P0001 , \wishbone_bd_ram_mem1_reg[136][10]/P0001 , \wishbone_bd_ram_mem1_reg[136][11]/P0001 , \wishbone_bd_ram_mem1_reg[136][12]/P0001 , \wishbone_bd_ram_mem1_reg[136][13]/P0001 , \wishbone_bd_ram_mem1_reg[136][14]/P0001 , \wishbone_bd_ram_mem1_reg[136][15]/P0001 , \wishbone_bd_ram_mem1_reg[136][8]/P0001 , \wishbone_bd_ram_mem1_reg[136][9]/P0001 , \wishbone_bd_ram_mem1_reg[137][10]/P0001 , \wishbone_bd_ram_mem1_reg[137][11]/P0001 , \wishbone_bd_ram_mem1_reg[137][12]/P0001 , \wishbone_bd_ram_mem1_reg[137][13]/P0001 , \wishbone_bd_ram_mem1_reg[137][14]/P0001 , \wishbone_bd_ram_mem1_reg[137][15]/P0001 , \wishbone_bd_ram_mem1_reg[137][8]/P0001 , \wishbone_bd_ram_mem1_reg[137][9]/P0001 , \wishbone_bd_ram_mem1_reg[138][10]/P0001 , \wishbone_bd_ram_mem1_reg[138][11]/P0001 , \wishbone_bd_ram_mem1_reg[138][12]/P0001 , \wishbone_bd_ram_mem1_reg[138][13]/P0001 , \wishbone_bd_ram_mem1_reg[138][14]/P0001 , \wishbone_bd_ram_mem1_reg[138][15]/P0001 , \wishbone_bd_ram_mem1_reg[138][8]/P0001 , \wishbone_bd_ram_mem1_reg[138][9]/P0001 , \wishbone_bd_ram_mem1_reg[139][10]/P0001 , \wishbone_bd_ram_mem1_reg[139][11]/P0001 , \wishbone_bd_ram_mem1_reg[139][12]/P0001 , \wishbone_bd_ram_mem1_reg[139][13]/P0001 , \wishbone_bd_ram_mem1_reg[139][14]/P0001 , \wishbone_bd_ram_mem1_reg[139][15]/P0001 , \wishbone_bd_ram_mem1_reg[139][8]/P0001 , \wishbone_bd_ram_mem1_reg[139][9]/P0001 , \wishbone_bd_ram_mem1_reg[13][10]/P0001 , \wishbone_bd_ram_mem1_reg[13][11]/P0001 , \wishbone_bd_ram_mem1_reg[13][12]/P0001 , \wishbone_bd_ram_mem1_reg[13][13]/P0001 , \wishbone_bd_ram_mem1_reg[13][14]/P0001 , \wishbone_bd_ram_mem1_reg[13][15]/P0001 , \wishbone_bd_ram_mem1_reg[13][8]/P0001 , \wishbone_bd_ram_mem1_reg[13][9]/P0001 , \wishbone_bd_ram_mem1_reg[140][10]/P0001 , \wishbone_bd_ram_mem1_reg[140][11]/P0001 , \wishbone_bd_ram_mem1_reg[140][12]/P0001 , \wishbone_bd_ram_mem1_reg[140][13]/P0001 , \wishbone_bd_ram_mem1_reg[140][14]/P0001 , \wishbone_bd_ram_mem1_reg[140][15]/P0001 , \wishbone_bd_ram_mem1_reg[140][8]/P0001 , \wishbone_bd_ram_mem1_reg[140][9]/P0001 , \wishbone_bd_ram_mem1_reg[141][10]/P0001 , \wishbone_bd_ram_mem1_reg[141][11]/P0001 , \wishbone_bd_ram_mem1_reg[141][12]/P0001 , \wishbone_bd_ram_mem1_reg[141][13]/P0001 , \wishbone_bd_ram_mem1_reg[141][14]/P0001 , \wishbone_bd_ram_mem1_reg[141][15]/P0001 , \wishbone_bd_ram_mem1_reg[141][8]/P0001 , \wishbone_bd_ram_mem1_reg[141][9]/P0001 , \wishbone_bd_ram_mem1_reg[142][10]/P0001 , \wishbone_bd_ram_mem1_reg[142][11]/P0001 , \wishbone_bd_ram_mem1_reg[142][12]/P0001 , \wishbone_bd_ram_mem1_reg[142][13]/P0001 , \wishbone_bd_ram_mem1_reg[142][14]/P0001 , \wishbone_bd_ram_mem1_reg[142][15]/P0001 , \wishbone_bd_ram_mem1_reg[142][8]/P0001 , \wishbone_bd_ram_mem1_reg[142][9]/P0001 , \wishbone_bd_ram_mem1_reg[143][10]/P0001 , \wishbone_bd_ram_mem1_reg[143][11]/P0001 , \wishbone_bd_ram_mem1_reg[143][12]/P0001 , \wishbone_bd_ram_mem1_reg[143][13]/P0001 , \wishbone_bd_ram_mem1_reg[143][14]/P0001 , \wishbone_bd_ram_mem1_reg[143][15]/P0001 , \wishbone_bd_ram_mem1_reg[143][8]/P0001 , \wishbone_bd_ram_mem1_reg[143][9]/P0001 , \wishbone_bd_ram_mem1_reg[144][10]/P0001 , \wishbone_bd_ram_mem1_reg[144][11]/P0001 , \wishbone_bd_ram_mem1_reg[144][12]/P0001 , \wishbone_bd_ram_mem1_reg[144][13]/P0001 , \wishbone_bd_ram_mem1_reg[144][14]/P0001 , \wishbone_bd_ram_mem1_reg[144][15]/P0001 , \wishbone_bd_ram_mem1_reg[144][8]/P0001 , \wishbone_bd_ram_mem1_reg[144][9]/P0001 , \wishbone_bd_ram_mem1_reg[145][10]/P0001 , \wishbone_bd_ram_mem1_reg[145][11]/P0001 , \wishbone_bd_ram_mem1_reg[145][12]/P0001 , \wishbone_bd_ram_mem1_reg[145][13]/P0001 , \wishbone_bd_ram_mem1_reg[145][14]/P0001 , \wishbone_bd_ram_mem1_reg[145][15]/P0001 , \wishbone_bd_ram_mem1_reg[145][8]/P0001 , \wishbone_bd_ram_mem1_reg[145][9]/P0001 , \wishbone_bd_ram_mem1_reg[146][10]/P0001 , \wishbone_bd_ram_mem1_reg[146][11]/P0001 , \wishbone_bd_ram_mem1_reg[146][12]/P0001 , \wishbone_bd_ram_mem1_reg[146][13]/P0001 , \wishbone_bd_ram_mem1_reg[146][14]/P0001 , \wishbone_bd_ram_mem1_reg[146][15]/P0001 , \wishbone_bd_ram_mem1_reg[146][8]/P0001 , \wishbone_bd_ram_mem1_reg[146][9]/P0001 , \wishbone_bd_ram_mem1_reg[147][10]/P0001 , \wishbone_bd_ram_mem1_reg[147][11]/P0001 , \wishbone_bd_ram_mem1_reg[147][12]/P0001 , \wishbone_bd_ram_mem1_reg[147][13]/P0001 , \wishbone_bd_ram_mem1_reg[147][14]/P0001 , \wishbone_bd_ram_mem1_reg[147][15]/P0001 , \wishbone_bd_ram_mem1_reg[147][8]/P0001 , \wishbone_bd_ram_mem1_reg[147][9]/P0001 , \wishbone_bd_ram_mem1_reg[148][10]/P0001 , \wishbone_bd_ram_mem1_reg[148][11]/P0001 , \wishbone_bd_ram_mem1_reg[148][12]/P0001 , \wishbone_bd_ram_mem1_reg[148][13]/P0001 , \wishbone_bd_ram_mem1_reg[148][14]/P0001 , \wishbone_bd_ram_mem1_reg[148][15]/P0001 , \wishbone_bd_ram_mem1_reg[148][8]/P0001 , \wishbone_bd_ram_mem1_reg[148][9]/P0001 , \wishbone_bd_ram_mem1_reg[149][10]/P0001 , \wishbone_bd_ram_mem1_reg[149][11]/P0001 , \wishbone_bd_ram_mem1_reg[149][12]/P0001 , \wishbone_bd_ram_mem1_reg[149][13]/P0001 , \wishbone_bd_ram_mem1_reg[149][14]/P0001 , \wishbone_bd_ram_mem1_reg[149][15]/P0001 , \wishbone_bd_ram_mem1_reg[149][8]/P0001 , \wishbone_bd_ram_mem1_reg[149][9]/P0001 , \wishbone_bd_ram_mem1_reg[14][10]/P0001 , \wishbone_bd_ram_mem1_reg[14][11]/P0001 , \wishbone_bd_ram_mem1_reg[14][12]/P0001 , \wishbone_bd_ram_mem1_reg[14][13]/P0001 , \wishbone_bd_ram_mem1_reg[14][14]/P0001 , \wishbone_bd_ram_mem1_reg[14][15]/P0001 , \wishbone_bd_ram_mem1_reg[14][8]/P0001 , \wishbone_bd_ram_mem1_reg[14][9]/P0001 , \wishbone_bd_ram_mem1_reg[150][10]/P0001 , \wishbone_bd_ram_mem1_reg[150][11]/P0001 , \wishbone_bd_ram_mem1_reg[150][12]/P0001 , \wishbone_bd_ram_mem1_reg[150][13]/P0001 , \wishbone_bd_ram_mem1_reg[150][14]/P0001 , \wishbone_bd_ram_mem1_reg[150][15]/P0001 , \wishbone_bd_ram_mem1_reg[150][8]/P0001 , \wishbone_bd_ram_mem1_reg[150][9]/P0001 , \wishbone_bd_ram_mem1_reg[151][10]/P0001 , \wishbone_bd_ram_mem1_reg[151][11]/P0001 , \wishbone_bd_ram_mem1_reg[151][12]/P0001 , \wishbone_bd_ram_mem1_reg[151][13]/P0001 , \wishbone_bd_ram_mem1_reg[151][14]/P0001 , \wishbone_bd_ram_mem1_reg[151][15]/P0001 , \wishbone_bd_ram_mem1_reg[151][8]/P0001 , \wishbone_bd_ram_mem1_reg[151][9]/P0001 , \wishbone_bd_ram_mem1_reg[152][10]/P0001 , \wishbone_bd_ram_mem1_reg[152][11]/P0001 , \wishbone_bd_ram_mem1_reg[152][12]/P0001 , \wishbone_bd_ram_mem1_reg[152][13]/P0001 , \wishbone_bd_ram_mem1_reg[152][14]/P0001 , \wishbone_bd_ram_mem1_reg[152][15]/P0001 , \wishbone_bd_ram_mem1_reg[152][8]/P0001 , \wishbone_bd_ram_mem1_reg[152][9]/P0001 , \wishbone_bd_ram_mem1_reg[153][10]/P0001 , \wishbone_bd_ram_mem1_reg[153][11]/P0001 , \wishbone_bd_ram_mem1_reg[153][12]/P0001 , \wishbone_bd_ram_mem1_reg[153][13]/P0001 , \wishbone_bd_ram_mem1_reg[153][14]/P0001 , \wishbone_bd_ram_mem1_reg[153][15]/P0001 , \wishbone_bd_ram_mem1_reg[153][8]/P0001 , \wishbone_bd_ram_mem1_reg[153][9]/P0001 , \wishbone_bd_ram_mem1_reg[154][10]/P0001 , \wishbone_bd_ram_mem1_reg[154][11]/P0001 , \wishbone_bd_ram_mem1_reg[154][12]/P0001 , \wishbone_bd_ram_mem1_reg[154][13]/P0001 , \wishbone_bd_ram_mem1_reg[154][14]/P0001 , \wishbone_bd_ram_mem1_reg[154][15]/P0001 , \wishbone_bd_ram_mem1_reg[154][8]/P0001 , \wishbone_bd_ram_mem1_reg[154][9]/P0001 , \wishbone_bd_ram_mem1_reg[155][10]/P0001 , \wishbone_bd_ram_mem1_reg[155][11]/P0001 , \wishbone_bd_ram_mem1_reg[155][12]/P0001 , \wishbone_bd_ram_mem1_reg[155][13]/P0001 , \wishbone_bd_ram_mem1_reg[155][14]/P0001 , \wishbone_bd_ram_mem1_reg[155][15]/P0001 , \wishbone_bd_ram_mem1_reg[155][8]/P0001 , \wishbone_bd_ram_mem1_reg[155][9]/P0001 , \wishbone_bd_ram_mem1_reg[156][10]/P0001 , \wishbone_bd_ram_mem1_reg[156][11]/P0001 , \wishbone_bd_ram_mem1_reg[156][12]/P0001 , \wishbone_bd_ram_mem1_reg[156][13]/P0001 , \wishbone_bd_ram_mem1_reg[156][14]/P0001 , \wishbone_bd_ram_mem1_reg[156][15]/P0001 , \wishbone_bd_ram_mem1_reg[156][8]/P0001 , \wishbone_bd_ram_mem1_reg[156][9]/P0001 , \wishbone_bd_ram_mem1_reg[157][10]/P0001 , \wishbone_bd_ram_mem1_reg[157][11]/P0001 , \wishbone_bd_ram_mem1_reg[157][12]/P0001 , \wishbone_bd_ram_mem1_reg[157][13]/P0001 , \wishbone_bd_ram_mem1_reg[157][14]/P0001 , \wishbone_bd_ram_mem1_reg[157][15]/P0001 , \wishbone_bd_ram_mem1_reg[157][8]/P0001 , \wishbone_bd_ram_mem1_reg[157][9]/P0001 , \wishbone_bd_ram_mem1_reg[158][10]/P0001 , \wishbone_bd_ram_mem1_reg[158][11]/P0001 , \wishbone_bd_ram_mem1_reg[158][12]/P0001 , \wishbone_bd_ram_mem1_reg[158][13]/P0001 , \wishbone_bd_ram_mem1_reg[158][14]/P0001 , \wishbone_bd_ram_mem1_reg[158][15]/P0001 , \wishbone_bd_ram_mem1_reg[158][8]/P0001 , \wishbone_bd_ram_mem1_reg[158][9]/P0001 , \wishbone_bd_ram_mem1_reg[159][10]/P0001 , \wishbone_bd_ram_mem1_reg[159][11]/P0001 , \wishbone_bd_ram_mem1_reg[159][12]/P0001 , \wishbone_bd_ram_mem1_reg[159][13]/P0001 , \wishbone_bd_ram_mem1_reg[159][14]/P0001 , \wishbone_bd_ram_mem1_reg[159][15]/P0001 , \wishbone_bd_ram_mem1_reg[159][8]/P0001 , \wishbone_bd_ram_mem1_reg[159][9]/P0001 , \wishbone_bd_ram_mem1_reg[15][10]/P0001 , \wishbone_bd_ram_mem1_reg[15][11]/P0001 , \wishbone_bd_ram_mem1_reg[15][12]/P0001 , \wishbone_bd_ram_mem1_reg[15][13]/P0001 , \wishbone_bd_ram_mem1_reg[15][14]/P0001 , \wishbone_bd_ram_mem1_reg[15][15]/P0001 , \wishbone_bd_ram_mem1_reg[15][8]/P0001 , \wishbone_bd_ram_mem1_reg[15][9]/P0001 , \wishbone_bd_ram_mem1_reg[160][10]/P0001 , \wishbone_bd_ram_mem1_reg[160][11]/P0001 , \wishbone_bd_ram_mem1_reg[160][12]/P0001 , \wishbone_bd_ram_mem1_reg[160][13]/P0001 , \wishbone_bd_ram_mem1_reg[160][14]/P0001 , \wishbone_bd_ram_mem1_reg[160][15]/P0001 , \wishbone_bd_ram_mem1_reg[160][8]/P0001 , \wishbone_bd_ram_mem1_reg[160][9]/P0001 , \wishbone_bd_ram_mem1_reg[161][10]/P0001 , \wishbone_bd_ram_mem1_reg[161][11]/P0001 , \wishbone_bd_ram_mem1_reg[161][12]/P0001 , \wishbone_bd_ram_mem1_reg[161][13]/P0001 , \wishbone_bd_ram_mem1_reg[161][14]/P0001 , \wishbone_bd_ram_mem1_reg[161][15]/P0001 , \wishbone_bd_ram_mem1_reg[161][8]/P0001 , \wishbone_bd_ram_mem1_reg[161][9]/P0001 , \wishbone_bd_ram_mem1_reg[162][10]/P0001 , \wishbone_bd_ram_mem1_reg[162][11]/P0001 , \wishbone_bd_ram_mem1_reg[162][12]/P0001 , \wishbone_bd_ram_mem1_reg[162][13]/P0001 , \wishbone_bd_ram_mem1_reg[162][14]/P0001 , \wishbone_bd_ram_mem1_reg[162][15]/P0001 , \wishbone_bd_ram_mem1_reg[162][8]/P0001 , \wishbone_bd_ram_mem1_reg[162][9]/P0001 , \wishbone_bd_ram_mem1_reg[163][10]/P0001 , \wishbone_bd_ram_mem1_reg[163][11]/P0001 , \wishbone_bd_ram_mem1_reg[163][12]/P0001 , \wishbone_bd_ram_mem1_reg[163][13]/P0001 , \wishbone_bd_ram_mem1_reg[163][14]/P0001 , \wishbone_bd_ram_mem1_reg[163][15]/P0001 , \wishbone_bd_ram_mem1_reg[163][8]/P0001 , \wishbone_bd_ram_mem1_reg[163][9]/P0001 , \wishbone_bd_ram_mem1_reg[164][10]/P0001 , \wishbone_bd_ram_mem1_reg[164][11]/P0001 , \wishbone_bd_ram_mem1_reg[164][12]/P0001 , \wishbone_bd_ram_mem1_reg[164][13]/P0001 , \wishbone_bd_ram_mem1_reg[164][14]/P0001 , \wishbone_bd_ram_mem1_reg[164][15]/P0001 , \wishbone_bd_ram_mem1_reg[164][8]/P0001 , \wishbone_bd_ram_mem1_reg[164][9]/P0001 , \wishbone_bd_ram_mem1_reg[165][10]/P0001 , \wishbone_bd_ram_mem1_reg[165][11]/P0001 , \wishbone_bd_ram_mem1_reg[165][12]/P0001 , \wishbone_bd_ram_mem1_reg[165][13]/P0001 , \wishbone_bd_ram_mem1_reg[165][14]/P0001 , \wishbone_bd_ram_mem1_reg[165][15]/P0001 , \wishbone_bd_ram_mem1_reg[165][8]/P0001 , \wishbone_bd_ram_mem1_reg[165][9]/P0001 , \wishbone_bd_ram_mem1_reg[166][10]/P0001 , \wishbone_bd_ram_mem1_reg[166][11]/P0001 , \wishbone_bd_ram_mem1_reg[166][12]/P0001 , \wishbone_bd_ram_mem1_reg[166][13]/P0001 , \wishbone_bd_ram_mem1_reg[166][14]/P0001 , \wishbone_bd_ram_mem1_reg[166][15]/P0001 , \wishbone_bd_ram_mem1_reg[166][8]/P0001 , \wishbone_bd_ram_mem1_reg[166][9]/P0001 , \wishbone_bd_ram_mem1_reg[167][10]/P0001 , \wishbone_bd_ram_mem1_reg[167][11]/P0001 , \wishbone_bd_ram_mem1_reg[167][12]/P0001 , \wishbone_bd_ram_mem1_reg[167][13]/P0001 , \wishbone_bd_ram_mem1_reg[167][14]/P0001 , \wishbone_bd_ram_mem1_reg[167][15]/P0001 , \wishbone_bd_ram_mem1_reg[167][8]/P0001 , \wishbone_bd_ram_mem1_reg[167][9]/P0001 , \wishbone_bd_ram_mem1_reg[168][10]/P0001 , \wishbone_bd_ram_mem1_reg[168][11]/P0001 , \wishbone_bd_ram_mem1_reg[168][12]/P0001 , \wishbone_bd_ram_mem1_reg[168][13]/P0001 , \wishbone_bd_ram_mem1_reg[168][14]/P0001 , \wishbone_bd_ram_mem1_reg[168][15]/P0001 , \wishbone_bd_ram_mem1_reg[168][8]/P0001 , \wishbone_bd_ram_mem1_reg[168][9]/P0001 , \wishbone_bd_ram_mem1_reg[169][10]/P0001 , \wishbone_bd_ram_mem1_reg[169][11]/P0001 , \wishbone_bd_ram_mem1_reg[169][12]/P0001 , \wishbone_bd_ram_mem1_reg[169][13]/P0001 , \wishbone_bd_ram_mem1_reg[169][14]/P0001 , \wishbone_bd_ram_mem1_reg[169][15]/P0001 , \wishbone_bd_ram_mem1_reg[169][8]/P0001 , \wishbone_bd_ram_mem1_reg[169][9]/P0001 , \wishbone_bd_ram_mem1_reg[16][10]/P0001 , \wishbone_bd_ram_mem1_reg[16][11]/P0001 , \wishbone_bd_ram_mem1_reg[16][12]/P0001 , \wishbone_bd_ram_mem1_reg[16][13]/P0001 , \wishbone_bd_ram_mem1_reg[16][14]/P0001 , \wishbone_bd_ram_mem1_reg[16][15]/P0001 , \wishbone_bd_ram_mem1_reg[16][8]/P0001 , \wishbone_bd_ram_mem1_reg[16][9]/P0001 , \wishbone_bd_ram_mem1_reg[170][10]/P0001 , \wishbone_bd_ram_mem1_reg[170][11]/P0001 , \wishbone_bd_ram_mem1_reg[170][12]/P0001 , \wishbone_bd_ram_mem1_reg[170][13]/P0001 , \wishbone_bd_ram_mem1_reg[170][14]/P0001 , \wishbone_bd_ram_mem1_reg[170][15]/P0001 , \wishbone_bd_ram_mem1_reg[170][8]/P0001 , \wishbone_bd_ram_mem1_reg[170][9]/P0001 , \wishbone_bd_ram_mem1_reg[171][10]/P0001 , \wishbone_bd_ram_mem1_reg[171][11]/P0001 , \wishbone_bd_ram_mem1_reg[171][12]/P0001 , \wishbone_bd_ram_mem1_reg[171][13]/P0001 , \wishbone_bd_ram_mem1_reg[171][14]/P0001 , \wishbone_bd_ram_mem1_reg[171][15]/P0001 , \wishbone_bd_ram_mem1_reg[171][8]/P0001 , \wishbone_bd_ram_mem1_reg[171][9]/P0001 , \wishbone_bd_ram_mem1_reg[172][10]/P0001 , \wishbone_bd_ram_mem1_reg[172][11]/P0001 , \wishbone_bd_ram_mem1_reg[172][12]/P0001 , \wishbone_bd_ram_mem1_reg[172][13]/P0001 , \wishbone_bd_ram_mem1_reg[172][14]/P0001 , \wishbone_bd_ram_mem1_reg[172][15]/P0001 , \wishbone_bd_ram_mem1_reg[172][8]/P0001 , \wishbone_bd_ram_mem1_reg[172][9]/P0001 , \wishbone_bd_ram_mem1_reg[173][10]/P0001 , \wishbone_bd_ram_mem1_reg[173][11]/P0001 , \wishbone_bd_ram_mem1_reg[173][12]/P0001 , \wishbone_bd_ram_mem1_reg[173][13]/P0001 , \wishbone_bd_ram_mem1_reg[173][14]/P0001 , \wishbone_bd_ram_mem1_reg[173][15]/P0001 , \wishbone_bd_ram_mem1_reg[173][8]/P0001 , \wishbone_bd_ram_mem1_reg[173][9]/P0001 , \wishbone_bd_ram_mem1_reg[174][10]/P0001 , \wishbone_bd_ram_mem1_reg[174][11]/P0001 , \wishbone_bd_ram_mem1_reg[174][12]/P0001 , \wishbone_bd_ram_mem1_reg[174][13]/P0001 , \wishbone_bd_ram_mem1_reg[174][14]/P0001 , \wishbone_bd_ram_mem1_reg[174][15]/P0001 , \wishbone_bd_ram_mem1_reg[174][8]/P0001 , \wishbone_bd_ram_mem1_reg[174][9]/P0001 , \wishbone_bd_ram_mem1_reg[175][10]/P0001 , \wishbone_bd_ram_mem1_reg[175][11]/P0001 , \wishbone_bd_ram_mem1_reg[175][12]/P0001 , \wishbone_bd_ram_mem1_reg[175][13]/P0001 , \wishbone_bd_ram_mem1_reg[175][14]/P0001 , \wishbone_bd_ram_mem1_reg[175][15]/P0001 , \wishbone_bd_ram_mem1_reg[175][8]/P0001 , \wishbone_bd_ram_mem1_reg[175][9]/P0001 , \wishbone_bd_ram_mem1_reg[176][10]/P0001 , \wishbone_bd_ram_mem1_reg[176][11]/P0001 , \wishbone_bd_ram_mem1_reg[176][12]/P0001 , \wishbone_bd_ram_mem1_reg[176][13]/P0001 , \wishbone_bd_ram_mem1_reg[176][14]/P0001 , \wishbone_bd_ram_mem1_reg[176][15]/P0001 , \wishbone_bd_ram_mem1_reg[176][8]/P0001 , \wishbone_bd_ram_mem1_reg[176][9]/P0001 , \wishbone_bd_ram_mem1_reg[177][10]/P0001 , \wishbone_bd_ram_mem1_reg[177][11]/P0001 , \wishbone_bd_ram_mem1_reg[177][12]/P0001 , \wishbone_bd_ram_mem1_reg[177][13]/P0001 , \wishbone_bd_ram_mem1_reg[177][14]/P0001 , \wishbone_bd_ram_mem1_reg[177][15]/P0001 , \wishbone_bd_ram_mem1_reg[177][8]/P0001 , \wishbone_bd_ram_mem1_reg[177][9]/P0001 , \wishbone_bd_ram_mem1_reg[178][10]/P0001 , \wishbone_bd_ram_mem1_reg[178][11]/P0001 , \wishbone_bd_ram_mem1_reg[178][12]/P0001 , \wishbone_bd_ram_mem1_reg[178][13]/P0001 , \wishbone_bd_ram_mem1_reg[178][14]/P0001 , \wishbone_bd_ram_mem1_reg[178][15]/P0001 , \wishbone_bd_ram_mem1_reg[178][8]/P0001 , \wishbone_bd_ram_mem1_reg[178][9]/P0001 , \wishbone_bd_ram_mem1_reg[179][10]/P0001 , \wishbone_bd_ram_mem1_reg[179][11]/P0001 , \wishbone_bd_ram_mem1_reg[179][12]/P0001 , \wishbone_bd_ram_mem1_reg[179][13]/P0001 , \wishbone_bd_ram_mem1_reg[179][14]/P0001 , \wishbone_bd_ram_mem1_reg[179][15]/P0001 , \wishbone_bd_ram_mem1_reg[179][8]/P0001 , \wishbone_bd_ram_mem1_reg[179][9]/P0001 , \wishbone_bd_ram_mem1_reg[17][10]/P0001 , \wishbone_bd_ram_mem1_reg[17][11]/P0001 , \wishbone_bd_ram_mem1_reg[17][12]/P0001 , \wishbone_bd_ram_mem1_reg[17][13]/P0001 , \wishbone_bd_ram_mem1_reg[17][14]/P0001 , \wishbone_bd_ram_mem1_reg[17][15]/P0001 , \wishbone_bd_ram_mem1_reg[17][8]/P0001 , \wishbone_bd_ram_mem1_reg[17][9]/P0001 , \wishbone_bd_ram_mem1_reg[180][10]/P0001 , \wishbone_bd_ram_mem1_reg[180][11]/P0001 , \wishbone_bd_ram_mem1_reg[180][12]/P0001 , \wishbone_bd_ram_mem1_reg[180][13]/P0001 , \wishbone_bd_ram_mem1_reg[180][14]/P0001 , \wishbone_bd_ram_mem1_reg[180][15]/P0001 , \wishbone_bd_ram_mem1_reg[180][8]/P0001 , \wishbone_bd_ram_mem1_reg[180][9]/P0001 , \wishbone_bd_ram_mem1_reg[181][10]/P0001 , \wishbone_bd_ram_mem1_reg[181][11]/P0001 , \wishbone_bd_ram_mem1_reg[181][12]/P0001 , \wishbone_bd_ram_mem1_reg[181][13]/P0001 , \wishbone_bd_ram_mem1_reg[181][14]/P0001 , \wishbone_bd_ram_mem1_reg[181][15]/P0001 , \wishbone_bd_ram_mem1_reg[181][8]/P0001 , \wishbone_bd_ram_mem1_reg[181][9]/P0001 , \wishbone_bd_ram_mem1_reg[182][10]/P0001 , \wishbone_bd_ram_mem1_reg[182][11]/P0001 , \wishbone_bd_ram_mem1_reg[182][12]/P0001 , \wishbone_bd_ram_mem1_reg[182][13]/P0001 , \wishbone_bd_ram_mem1_reg[182][14]/P0001 , \wishbone_bd_ram_mem1_reg[182][15]/P0001 , \wishbone_bd_ram_mem1_reg[182][8]/P0001 , \wishbone_bd_ram_mem1_reg[182][9]/P0001 , \wishbone_bd_ram_mem1_reg[183][10]/P0001 , \wishbone_bd_ram_mem1_reg[183][11]/P0001 , \wishbone_bd_ram_mem1_reg[183][12]/P0001 , \wishbone_bd_ram_mem1_reg[183][13]/P0001 , \wishbone_bd_ram_mem1_reg[183][14]/P0001 , \wishbone_bd_ram_mem1_reg[183][15]/P0001 , \wishbone_bd_ram_mem1_reg[183][8]/P0001 , \wishbone_bd_ram_mem1_reg[183][9]/P0001 , \wishbone_bd_ram_mem1_reg[184][10]/P0001 , \wishbone_bd_ram_mem1_reg[184][11]/P0001 , \wishbone_bd_ram_mem1_reg[184][12]/P0001 , \wishbone_bd_ram_mem1_reg[184][13]/P0001 , \wishbone_bd_ram_mem1_reg[184][14]/P0001 , \wishbone_bd_ram_mem1_reg[184][15]/P0001 , \wishbone_bd_ram_mem1_reg[184][8]/P0001 , \wishbone_bd_ram_mem1_reg[184][9]/P0001 , \wishbone_bd_ram_mem1_reg[185][10]/P0001 , \wishbone_bd_ram_mem1_reg[185][11]/P0001 , \wishbone_bd_ram_mem1_reg[185][12]/P0001 , \wishbone_bd_ram_mem1_reg[185][13]/P0001 , \wishbone_bd_ram_mem1_reg[185][14]/P0001 , \wishbone_bd_ram_mem1_reg[185][15]/P0001 , \wishbone_bd_ram_mem1_reg[185][8]/P0001 , \wishbone_bd_ram_mem1_reg[185][9]/P0001 , \wishbone_bd_ram_mem1_reg[186][10]/P0001 , \wishbone_bd_ram_mem1_reg[186][11]/P0001 , \wishbone_bd_ram_mem1_reg[186][12]/P0001 , \wishbone_bd_ram_mem1_reg[186][13]/P0001 , \wishbone_bd_ram_mem1_reg[186][14]/P0001 , \wishbone_bd_ram_mem1_reg[186][15]/P0001 , \wishbone_bd_ram_mem1_reg[186][8]/P0001 , \wishbone_bd_ram_mem1_reg[186][9]/P0001 , \wishbone_bd_ram_mem1_reg[187][10]/P0001 , \wishbone_bd_ram_mem1_reg[187][11]/P0001 , \wishbone_bd_ram_mem1_reg[187][12]/P0001 , \wishbone_bd_ram_mem1_reg[187][13]/P0001 , \wishbone_bd_ram_mem1_reg[187][14]/P0001 , \wishbone_bd_ram_mem1_reg[187][15]/P0001 , \wishbone_bd_ram_mem1_reg[187][8]/P0001 , \wishbone_bd_ram_mem1_reg[187][9]/P0001 , \wishbone_bd_ram_mem1_reg[188][10]/P0001 , \wishbone_bd_ram_mem1_reg[188][11]/P0001 , \wishbone_bd_ram_mem1_reg[188][12]/P0001 , \wishbone_bd_ram_mem1_reg[188][13]/P0001 , \wishbone_bd_ram_mem1_reg[188][14]/P0001 , \wishbone_bd_ram_mem1_reg[188][15]/P0001 , \wishbone_bd_ram_mem1_reg[188][8]/P0001 , \wishbone_bd_ram_mem1_reg[188][9]/P0001 , \wishbone_bd_ram_mem1_reg[189][10]/P0001 , \wishbone_bd_ram_mem1_reg[189][11]/P0001 , \wishbone_bd_ram_mem1_reg[189][12]/P0001 , \wishbone_bd_ram_mem1_reg[189][13]/P0001 , \wishbone_bd_ram_mem1_reg[189][14]/P0001 , \wishbone_bd_ram_mem1_reg[189][15]/P0001 , \wishbone_bd_ram_mem1_reg[189][8]/P0001 , \wishbone_bd_ram_mem1_reg[189][9]/P0001 , \wishbone_bd_ram_mem1_reg[18][10]/P0001 , \wishbone_bd_ram_mem1_reg[18][11]/P0001 , \wishbone_bd_ram_mem1_reg[18][12]/P0001 , \wishbone_bd_ram_mem1_reg[18][13]/P0001 , \wishbone_bd_ram_mem1_reg[18][14]/P0001 , \wishbone_bd_ram_mem1_reg[18][15]/P0001 , \wishbone_bd_ram_mem1_reg[18][8]/P0001 , \wishbone_bd_ram_mem1_reg[18][9]/P0001 , \wishbone_bd_ram_mem1_reg[190][10]/P0001 , \wishbone_bd_ram_mem1_reg[190][11]/P0001 , \wishbone_bd_ram_mem1_reg[190][12]/P0001 , \wishbone_bd_ram_mem1_reg[190][13]/P0001 , \wishbone_bd_ram_mem1_reg[190][14]/P0001 , \wishbone_bd_ram_mem1_reg[190][15]/P0001 , \wishbone_bd_ram_mem1_reg[190][8]/P0001 , \wishbone_bd_ram_mem1_reg[190][9]/P0001 , \wishbone_bd_ram_mem1_reg[191][10]/P0001 , \wishbone_bd_ram_mem1_reg[191][11]/P0001 , \wishbone_bd_ram_mem1_reg[191][12]/P0001 , \wishbone_bd_ram_mem1_reg[191][13]/P0001 , \wishbone_bd_ram_mem1_reg[191][14]/P0001 , \wishbone_bd_ram_mem1_reg[191][15]/P0001 , \wishbone_bd_ram_mem1_reg[191][8]/P0001 , \wishbone_bd_ram_mem1_reg[191][9]/P0001 , \wishbone_bd_ram_mem1_reg[192][10]/P0001 , \wishbone_bd_ram_mem1_reg[192][11]/P0001 , \wishbone_bd_ram_mem1_reg[192][12]/P0001 , \wishbone_bd_ram_mem1_reg[192][13]/P0001 , \wishbone_bd_ram_mem1_reg[192][14]/P0001 , \wishbone_bd_ram_mem1_reg[192][15]/P0001 , \wishbone_bd_ram_mem1_reg[192][8]/P0001 , \wishbone_bd_ram_mem1_reg[192][9]/P0001 , \wishbone_bd_ram_mem1_reg[193][10]/P0001 , \wishbone_bd_ram_mem1_reg[193][11]/P0001 , \wishbone_bd_ram_mem1_reg[193][12]/P0001 , \wishbone_bd_ram_mem1_reg[193][13]/P0001 , \wishbone_bd_ram_mem1_reg[193][14]/P0001 , \wishbone_bd_ram_mem1_reg[193][15]/P0001 , \wishbone_bd_ram_mem1_reg[193][8]/P0001 , \wishbone_bd_ram_mem1_reg[193][9]/P0001 , \wishbone_bd_ram_mem1_reg[194][10]/P0001 , \wishbone_bd_ram_mem1_reg[194][11]/P0001 , \wishbone_bd_ram_mem1_reg[194][12]/P0001 , \wishbone_bd_ram_mem1_reg[194][13]/P0001 , \wishbone_bd_ram_mem1_reg[194][14]/P0001 , \wishbone_bd_ram_mem1_reg[194][15]/P0001 , \wishbone_bd_ram_mem1_reg[194][8]/P0001 , \wishbone_bd_ram_mem1_reg[194][9]/P0001 , \wishbone_bd_ram_mem1_reg[195][10]/P0001 , \wishbone_bd_ram_mem1_reg[195][11]/P0001 , \wishbone_bd_ram_mem1_reg[195][12]/P0001 , \wishbone_bd_ram_mem1_reg[195][13]/P0001 , \wishbone_bd_ram_mem1_reg[195][14]/P0001 , \wishbone_bd_ram_mem1_reg[195][15]/P0001 , \wishbone_bd_ram_mem1_reg[195][8]/P0001 , \wishbone_bd_ram_mem1_reg[195][9]/P0001 , \wishbone_bd_ram_mem1_reg[196][10]/P0001 , \wishbone_bd_ram_mem1_reg[196][11]/P0001 , \wishbone_bd_ram_mem1_reg[196][12]/P0001 , \wishbone_bd_ram_mem1_reg[196][13]/P0001 , \wishbone_bd_ram_mem1_reg[196][14]/P0001 , \wishbone_bd_ram_mem1_reg[196][15]/P0001 , \wishbone_bd_ram_mem1_reg[196][8]/P0001 , \wishbone_bd_ram_mem1_reg[196][9]/P0001 , \wishbone_bd_ram_mem1_reg[197][10]/P0001 , \wishbone_bd_ram_mem1_reg[197][11]/P0001 , \wishbone_bd_ram_mem1_reg[197][12]/P0001 , \wishbone_bd_ram_mem1_reg[197][13]/P0001 , \wishbone_bd_ram_mem1_reg[197][14]/P0001 , \wishbone_bd_ram_mem1_reg[197][15]/P0001 , \wishbone_bd_ram_mem1_reg[197][8]/P0001 , \wishbone_bd_ram_mem1_reg[197][9]/P0001 , \wishbone_bd_ram_mem1_reg[198][10]/P0001 , \wishbone_bd_ram_mem1_reg[198][11]/P0001 , \wishbone_bd_ram_mem1_reg[198][12]/P0001 , \wishbone_bd_ram_mem1_reg[198][13]/P0001 , \wishbone_bd_ram_mem1_reg[198][14]/P0001 , \wishbone_bd_ram_mem1_reg[198][15]/P0001 , \wishbone_bd_ram_mem1_reg[198][8]/P0001 , \wishbone_bd_ram_mem1_reg[198][9]/P0001 , \wishbone_bd_ram_mem1_reg[199][10]/P0001 , \wishbone_bd_ram_mem1_reg[199][11]/P0001 , \wishbone_bd_ram_mem1_reg[199][12]/P0001 , \wishbone_bd_ram_mem1_reg[199][13]/P0001 , \wishbone_bd_ram_mem1_reg[199][14]/P0001 , \wishbone_bd_ram_mem1_reg[199][15]/P0001 , \wishbone_bd_ram_mem1_reg[199][8]/P0001 , \wishbone_bd_ram_mem1_reg[199][9]/P0001 , \wishbone_bd_ram_mem1_reg[19][10]/P0001 , \wishbone_bd_ram_mem1_reg[19][11]/P0001 , \wishbone_bd_ram_mem1_reg[19][12]/P0001 , \wishbone_bd_ram_mem1_reg[19][13]/P0001 , \wishbone_bd_ram_mem1_reg[19][14]/P0001 , \wishbone_bd_ram_mem1_reg[19][15]/P0001 , \wishbone_bd_ram_mem1_reg[19][8]/P0001 , \wishbone_bd_ram_mem1_reg[19][9]/P0001 , \wishbone_bd_ram_mem1_reg[1][10]/P0001 , \wishbone_bd_ram_mem1_reg[1][11]/P0001 , \wishbone_bd_ram_mem1_reg[1][12]/P0001 , \wishbone_bd_ram_mem1_reg[1][13]/P0001 , \wishbone_bd_ram_mem1_reg[1][14]/P0001 , \wishbone_bd_ram_mem1_reg[1][15]/P0001 , \wishbone_bd_ram_mem1_reg[1][8]/P0001 , \wishbone_bd_ram_mem1_reg[1][9]/P0001 , \wishbone_bd_ram_mem1_reg[200][10]/P0001 , \wishbone_bd_ram_mem1_reg[200][11]/P0001 , \wishbone_bd_ram_mem1_reg[200][12]/P0001 , \wishbone_bd_ram_mem1_reg[200][13]/P0001 , \wishbone_bd_ram_mem1_reg[200][14]/P0001 , \wishbone_bd_ram_mem1_reg[200][15]/P0001 , \wishbone_bd_ram_mem1_reg[200][8]/P0001 , \wishbone_bd_ram_mem1_reg[200][9]/P0001 , \wishbone_bd_ram_mem1_reg[201][10]/P0001 , \wishbone_bd_ram_mem1_reg[201][11]/P0001 , \wishbone_bd_ram_mem1_reg[201][12]/P0001 , \wishbone_bd_ram_mem1_reg[201][13]/P0001 , \wishbone_bd_ram_mem1_reg[201][14]/P0001 , \wishbone_bd_ram_mem1_reg[201][15]/P0001 , \wishbone_bd_ram_mem1_reg[201][8]/P0001 , \wishbone_bd_ram_mem1_reg[201][9]/P0001 , \wishbone_bd_ram_mem1_reg[202][10]/P0001 , \wishbone_bd_ram_mem1_reg[202][11]/P0001 , \wishbone_bd_ram_mem1_reg[202][12]/P0001 , \wishbone_bd_ram_mem1_reg[202][13]/P0001 , \wishbone_bd_ram_mem1_reg[202][14]/P0001 , \wishbone_bd_ram_mem1_reg[202][15]/P0001 , \wishbone_bd_ram_mem1_reg[202][8]/P0001 , \wishbone_bd_ram_mem1_reg[202][9]/P0001 , \wishbone_bd_ram_mem1_reg[203][10]/P0001 , \wishbone_bd_ram_mem1_reg[203][11]/P0001 , \wishbone_bd_ram_mem1_reg[203][12]/P0001 , \wishbone_bd_ram_mem1_reg[203][13]/P0001 , \wishbone_bd_ram_mem1_reg[203][14]/P0001 , \wishbone_bd_ram_mem1_reg[203][15]/P0001 , \wishbone_bd_ram_mem1_reg[203][8]/P0001 , \wishbone_bd_ram_mem1_reg[203][9]/P0001 , \wishbone_bd_ram_mem1_reg[204][10]/P0001 , \wishbone_bd_ram_mem1_reg[204][11]/P0001 , \wishbone_bd_ram_mem1_reg[204][12]/P0001 , \wishbone_bd_ram_mem1_reg[204][13]/P0001 , \wishbone_bd_ram_mem1_reg[204][14]/P0001 , \wishbone_bd_ram_mem1_reg[204][15]/P0001 , \wishbone_bd_ram_mem1_reg[204][8]/P0001 , \wishbone_bd_ram_mem1_reg[204][9]/P0001 , \wishbone_bd_ram_mem1_reg[205][10]/P0001 , \wishbone_bd_ram_mem1_reg[205][11]/P0001 , \wishbone_bd_ram_mem1_reg[205][12]/P0001 , \wishbone_bd_ram_mem1_reg[205][13]/P0001 , \wishbone_bd_ram_mem1_reg[205][14]/P0001 , \wishbone_bd_ram_mem1_reg[205][15]/P0001 , \wishbone_bd_ram_mem1_reg[205][8]/P0001 , \wishbone_bd_ram_mem1_reg[205][9]/P0001 , \wishbone_bd_ram_mem1_reg[206][10]/P0001 , \wishbone_bd_ram_mem1_reg[206][11]/P0001 , \wishbone_bd_ram_mem1_reg[206][12]/P0001 , \wishbone_bd_ram_mem1_reg[206][13]/P0001 , \wishbone_bd_ram_mem1_reg[206][14]/P0001 , \wishbone_bd_ram_mem1_reg[206][15]/P0001 , \wishbone_bd_ram_mem1_reg[206][8]/P0001 , \wishbone_bd_ram_mem1_reg[206][9]/P0001 , \wishbone_bd_ram_mem1_reg[207][10]/P0001 , \wishbone_bd_ram_mem1_reg[207][11]/P0001 , \wishbone_bd_ram_mem1_reg[207][12]/P0001 , \wishbone_bd_ram_mem1_reg[207][13]/P0001 , \wishbone_bd_ram_mem1_reg[207][14]/P0001 , \wishbone_bd_ram_mem1_reg[207][15]/P0001 , \wishbone_bd_ram_mem1_reg[207][8]/P0001 , \wishbone_bd_ram_mem1_reg[207][9]/P0001 , \wishbone_bd_ram_mem1_reg[208][10]/P0001 , \wishbone_bd_ram_mem1_reg[208][11]/P0001 , \wishbone_bd_ram_mem1_reg[208][12]/P0001 , \wishbone_bd_ram_mem1_reg[208][13]/P0001 , \wishbone_bd_ram_mem1_reg[208][14]/P0001 , \wishbone_bd_ram_mem1_reg[208][15]/P0001 , \wishbone_bd_ram_mem1_reg[208][8]/P0001 , \wishbone_bd_ram_mem1_reg[208][9]/P0001 , \wishbone_bd_ram_mem1_reg[209][10]/P0001 , \wishbone_bd_ram_mem1_reg[209][11]/P0001 , \wishbone_bd_ram_mem1_reg[209][12]/P0001 , \wishbone_bd_ram_mem1_reg[209][13]/P0001 , \wishbone_bd_ram_mem1_reg[209][14]/P0001 , \wishbone_bd_ram_mem1_reg[209][15]/P0001 , \wishbone_bd_ram_mem1_reg[209][8]/P0001 , \wishbone_bd_ram_mem1_reg[209][9]/P0001 , \wishbone_bd_ram_mem1_reg[20][10]/P0001 , \wishbone_bd_ram_mem1_reg[20][11]/P0001 , \wishbone_bd_ram_mem1_reg[20][12]/P0001 , \wishbone_bd_ram_mem1_reg[20][13]/P0001 , \wishbone_bd_ram_mem1_reg[20][14]/P0001 , \wishbone_bd_ram_mem1_reg[20][15]/P0001 , \wishbone_bd_ram_mem1_reg[20][8]/P0001 , \wishbone_bd_ram_mem1_reg[20][9]/P0001 , \wishbone_bd_ram_mem1_reg[210][10]/P0001 , \wishbone_bd_ram_mem1_reg[210][11]/P0001 , \wishbone_bd_ram_mem1_reg[210][12]/P0001 , \wishbone_bd_ram_mem1_reg[210][13]/P0001 , \wishbone_bd_ram_mem1_reg[210][14]/P0001 , \wishbone_bd_ram_mem1_reg[210][15]/P0001 , \wishbone_bd_ram_mem1_reg[210][8]/P0001 , \wishbone_bd_ram_mem1_reg[210][9]/P0001 , \wishbone_bd_ram_mem1_reg[211][10]/P0001 , \wishbone_bd_ram_mem1_reg[211][11]/P0001 , \wishbone_bd_ram_mem1_reg[211][12]/P0001 , \wishbone_bd_ram_mem1_reg[211][13]/P0001 , \wishbone_bd_ram_mem1_reg[211][14]/P0001 , \wishbone_bd_ram_mem1_reg[211][15]/P0001 , \wishbone_bd_ram_mem1_reg[211][8]/P0001 , \wishbone_bd_ram_mem1_reg[211][9]/P0001 , \wishbone_bd_ram_mem1_reg[212][10]/P0001 , \wishbone_bd_ram_mem1_reg[212][11]/P0001 , \wishbone_bd_ram_mem1_reg[212][12]/P0001 , \wishbone_bd_ram_mem1_reg[212][13]/P0001 , \wishbone_bd_ram_mem1_reg[212][14]/P0001 , \wishbone_bd_ram_mem1_reg[212][15]/P0001 , \wishbone_bd_ram_mem1_reg[212][8]/P0001 , \wishbone_bd_ram_mem1_reg[212][9]/P0001 , \wishbone_bd_ram_mem1_reg[213][10]/P0001 , \wishbone_bd_ram_mem1_reg[213][11]/P0001 , \wishbone_bd_ram_mem1_reg[213][12]/P0001 , \wishbone_bd_ram_mem1_reg[213][13]/P0001 , \wishbone_bd_ram_mem1_reg[213][14]/P0001 , \wishbone_bd_ram_mem1_reg[213][15]/P0001 , \wishbone_bd_ram_mem1_reg[213][8]/P0001 , \wishbone_bd_ram_mem1_reg[213][9]/P0001 , \wishbone_bd_ram_mem1_reg[214][10]/P0001 , \wishbone_bd_ram_mem1_reg[214][11]/P0001 , \wishbone_bd_ram_mem1_reg[214][12]/P0001 , \wishbone_bd_ram_mem1_reg[214][13]/P0001 , \wishbone_bd_ram_mem1_reg[214][14]/P0001 , \wishbone_bd_ram_mem1_reg[214][15]/P0001 , \wishbone_bd_ram_mem1_reg[214][8]/P0001 , \wishbone_bd_ram_mem1_reg[214][9]/P0001 , \wishbone_bd_ram_mem1_reg[215][10]/P0001 , \wishbone_bd_ram_mem1_reg[215][11]/P0001 , \wishbone_bd_ram_mem1_reg[215][12]/P0001 , \wishbone_bd_ram_mem1_reg[215][13]/P0001 , \wishbone_bd_ram_mem1_reg[215][14]/P0001 , \wishbone_bd_ram_mem1_reg[215][15]/P0001 , \wishbone_bd_ram_mem1_reg[215][8]/P0001 , \wishbone_bd_ram_mem1_reg[215][9]/P0001 , \wishbone_bd_ram_mem1_reg[216][10]/P0001 , \wishbone_bd_ram_mem1_reg[216][11]/P0001 , \wishbone_bd_ram_mem1_reg[216][12]/P0001 , \wishbone_bd_ram_mem1_reg[216][13]/P0001 , \wishbone_bd_ram_mem1_reg[216][14]/P0001 , \wishbone_bd_ram_mem1_reg[216][15]/P0001 , \wishbone_bd_ram_mem1_reg[216][8]/P0001 , \wishbone_bd_ram_mem1_reg[216][9]/P0001 , \wishbone_bd_ram_mem1_reg[217][10]/P0001 , \wishbone_bd_ram_mem1_reg[217][11]/P0001 , \wishbone_bd_ram_mem1_reg[217][12]/P0001 , \wishbone_bd_ram_mem1_reg[217][13]/P0001 , \wishbone_bd_ram_mem1_reg[217][14]/P0001 , \wishbone_bd_ram_mem1_reg[217][15]/P0001 , \wishbone_bd_ram_mem1_reg[217][8]/P0001 , \wishbone_bd_ram_mem1_reg[217][9]/P0001 , \wishbone_bd_ram_mem1_reg[218][10]/P0001 , \wishbone_bd_ram_mem1_reg[218][11]/P0001 , \wishbone_bd_ram_mem1_reg[218][12]/P0001 , \wishbone_bd_ram_mem1_reg[218][13]/P0001 , \wishbone_bd_ram_mem1_reg[218][14]/P0001 , \wishbone_bd_ram_mem1_reg[218][15]/P0001 , \wishbone_bd_ram_mem1_reg[218][8]/P0001 , \wishbone_bd_ram_mem1_reg[218][9]/P0001 , \wishbone_bd_ram_mem1_reg[219][10]/P0001 , \wishbone_bd_ram_mem1_reg[219][11]/P0001 , \wishbone_bd_ram_mem1_reg[219][12]/P0001 , \wishbone_bd_ram_mem1_reg[219][13]/P0001 , \wishbone_bd_ram_mem1_reg[219][14]/P0001 , \wishbone_bd_ram_mem1_reg[219][15]/P0001 , \wishbone_bd_ram_mem1_reg[219][8]/P0001 , \wishbone_bd_ram_mem1_reg[219][9]/P0001 , \wishbone_bd_ram_mem1_reg[21][10]/P0001 , \wishbone_bd_ram_mem1_reg[21][11]/P0001 , \wishbone_bd_ram_mem1_reg[21][12]/P0001 , \wishbone_bd_ram_mem1_reg[21][13]/P0001 , \wishbone_bd_ram_mem1_reg[21][14]/P0001 , \wishbone_bd_ram_mem1_reg[21][15]/P0001 , \wishbone_bd_ram_mem1_reg[21][8]/P0001 , \wishbone_bd_ram_mem1_reg[21][9]/P0001 , \wishbone_bd_ram_mem1_reg[220][10]/P0001 , \wishbone_bd_ram_mem1_reg[220][11]/P0001 , \wishbone_bd_ram_mem1_reg[220][12]/P0001 , \wishbone_bd_ram_mem1_reg[220][13]/P0001 , \wishbone_bd_ram_mem1_reg[220][14]/P0001 , \wishbone_bd_ram_mem1_reg[220][15]/P0001 , \wishbone_bd_ram_mem1_reg[220][8]/P0001 , \wishbone_bd_ram_mem1_reg[220][9]/P0001 , \wishbone_bd_ram_mem1_reg[221][10]/P0001 , \wishbone_bd_ram_mem1_reg[221][11]/P0001 , \wishbone_bd_ram_mem1_reg[221][12]/P0001 , \wishbone_bd_ram_mem1_reg[221][13]/P0001 , \wishbone_bd_ram_mem1_reg[221][14]/P0001 , \wishbone_bd_ram_mem1_reg[221][15]/P0001 , \wishbone_bd_ram_mem1_reg[221][8]/P0001 , \wishbone_bd_ram_mem1_reg[221][9]/P0001 , \wishbone_bd_ram_mem1_reg[222][10]/P0001 , \wishbone_bd_ram_mem1_reg[222][11]/P0001 , \wishbone_bd_ram_mem1_reg[222][12]/P0001 , \wishbone_bd_ram_mem1_reg[222][13]/P0001 , \wishbone_bd_ram_mem1_reg[222][14]/P0001 , \wishbone_bd_ram_mem1_reg[222][15]/P0001 , \wishbone_bd_ram_mem1_reg[222][8]/P0001 , \wishbone_bd_ram_mem1_reg[222][9]/P0001 , \wishbone_bd_ram_mem1_reg[223][10]/P0001 , \wishbone_bd_ram_mem1_reg[223][11]/P0001 , \wishbone_bd_ram_mem1_reg[223][12]/P0001 , \wishbone_bd_ram_mem1_reg[223][13]/P0001 , \wishbone_bd_ram_mem1_reg[223][14]/P0001 , \wishbone_bd_ram_mem1_reg[223][15]/P0001 , \wishbone_bd_ram_mem1_reg[223][8]/P0001 , \wishbone_bd_ram_mem1_reg[223][9]/P0001 , \wishbone_bd_ram_mem1_reg[224][10]/P0001 , \wishbone_bd_ram_mem1_reg[224][11]/P0001 , \wishbone_bd_ram_mem1_reg[224][12]/P0001 , \wishbone_bd_ram_mem1_reg[224][13]/P0001 , \wishbone_bd_ram_mem1_reg[224][14]/P0001 , \wishbone_bd_ram_mem1_reg[224][15]/P0001 , \wishbone_bd_ram_mem1_reg[224][8]/P0001 , \wishbone_bd_ram_mem1_reg[224][9]/P0001 , \wishbone_bd_ram_mem1_reg[225][10]/P0001 , \wishbone_bd_ram_mem1_reg[225][11]/P0001 , \wishbone_bd_ram_mem1_reg[225][12]/P0001 , \wishbone_bd_ram_mem1_reg[225][13]/P0001 , \wishbone_bd_ram_mem1_reg[225][14]/P0001 , \wishbone_bd_ram_mem1_reg[225][15]/P0001 , \wishbone_bd_ram_mem1_reg[225][8]/P0001 , \wishbone_bd_ram_mem1_reg[225][9]/P0001 , \wishbone_bd_ram_mem1_reg[226][10]/P0001 , \wishbone_bd_ram_mem1_reg[226][11]/P0001 , \wishbone_bd_ram_mem1_reg[226][12]/P0001 , \wishbone_bd_ram_mem1_reg[226][13]/P0001 , \wishbone_bd_ram_mem1_reg[226][14]/P0001 , \wishbone_bd_ram_mem1_reg[226][15]/P0001 , \wishbone_bd_ram_mem1_reg[226][8]/P0001 , \wishbone_bd_ram_mem1_reg[226][9]/P0001 , \wishbone_bd_ram_mem1_reg[227][10]/P0001 , \wishbone_bd_ram_mem1_reg[227][11]/P0001 , \wishbone_bd_ram_mem1_reg[227][12]/P0001 , \wishbone_bd_ram_mem1_reg[227][13]/P0001 , \wishbone_bd_ram_mem1_reg[227][14]/P0001 , \wishbone_bd_ram_mem1_reg[227][15]/P0001 , \wishbone_bd_ram_mem1_reg[227][8]/P0001 , \wishbone_bd_ram_mem1_reg[227][9]/P0001 , \wishbone_bd_ram_mem1_reg[228][10]/P0001 , \wishbone_bd_ram_mem1_reg[228][11]/P0001 , \wishbone_bd_ram_mem1_reg[228][12]/P0001 , \wishbone_bd_ram_mem1_reg[228][13]/P0001 , \wishbone_bd_ram_mem1_reg[228][14]/P0001 , \wishbone_bd_ram_mem1_reg[228][15]/P0001 , \wishbone_bd_ram_mem1_reg[228][8]/P0001 , \wishbone_bd_ram_mem1_reg[228][9]/P0001 , \wishbone_bd_ram_mem1_reg[229][10]/P0001 , \wishbone_bd_ram_mem1_reg[229][11]/P0001 , \wishbone_bd_ram_mem1_reg[229][12]/P0001 , \wishbone_bd_ram_mem1_reg[229][13]/P0001 , \wishbone_bd_ram_mem1_reg[229][14]/P0001 , \wishbone_bd_ram_mem1_reg[229][15]/P0001 , \wishbone_bd_ram_mem1_reg[229][8]/P0001 , \wishbone_bd_ram_mem1_reg[229][9]/P0001 , \wishbone_bd_ram_mem1_reg[22][10]/P0001 , \wishbone_bd_ram_mem1_reg[22][11]/P0001 , \wishbone_bd_ram_mem1_reg[22][12]/P0001 , \wishbone_bd_ram_mem1_reg[22][13]/P0001 , \wishbone_bd_ram_mem1_reg[22][14]/P0001 , \wishbone_bd_ram_mem1_reg[22][15]/P0001 , \wishbone_bd_ram_mem1_reg[22][8]/P0001 , \wishbone_bd_ram_mem1_reg[22][9]/P0001 , \wishbone_bd_ram_mem1_reg[230][10]/P0001 , \wishbone_bd_ram_mem1_reg[230][11]/P0001 , \wishbone_bd_ram_mem1_reg[230][12]/P0001 , \wishbone_bd_ram_mem1_reg[230][13]/P0001 , \wishbone_bd_ram_mem1_reg[230][14]/P0001 , \wishbone_bd_ram_mem1_reg[230][15]/P0001 , \wishbone_bd_ram_mem1_reg[230][8]/P0001 , \wishbone_bd_ram_mem1_reg[230][9]/P0001 , \wishbone_bd_ram_mem1_reg[231][10]/P0001 , \wishbone_bd_ram_mem1_reg[231][11]/P0001 , \wishbone_bd_ram_mem1_reg[231][12]/P0001 , \wishbone_bd_ram_mem1_reg[231][13]/P0001 , \wishbone_bd_ram_mem1_reg[231][14]/P0001 , \wishbone_bd_ram_mem1_reg[231][15]/P0001 , \wishbone_bd_ram_mem1_reg[231][8]/P0001 , \wishbone_bd_ram_mem1_reg[231][9]/P0001 , \wishbone_bd_ram_mem1_reg[232][10]/P0001 , \wishbone_bd_ram_mem1_reg[232][11]/P0001 , \wishbone_bd_ram_mem1_reg[232][12]/P0001 , \wishbone_bd_ram_mem1_reg[232][13]/P0001 , \wishbone_bd_ram_mem1_reg[232][14]/P0001 , \wishbone_bd_ram_mem1_reg[232][15]/P0001 , \wishbone_bd_ram_mem1_reg[232][8]/P0001 , \wishbone_bd_ram_mem1_reg[232][9]/P0001 , \wishbone_bd_ram_mem1_reg[233][10]/P0001 , \wishbone_bd_ram_mem1_reg[233][11]/P0001 , \wishbone_bd_ram_mem1_reg[233][12]/P0001 , \wishbone_bd_ram_mem1_reg[233][13]/P0001 , \wishbone_bd_ram_mem1_reg[233][14]/P0001 , \wishbone_bd_ram_mem1_reg[233][15]/P0001 , \wishbone_bd_ram_mem1_reg[233][8]/P0001 , \wishbone_bd_ram_mem1_reg[233][9]/P0001 , \wishbone_bd_ram_mem1_reg[234][10]/P0001 , \wishbone_bd_ram_mem1_reg[234][11]/P0001 , \wishbone_bd_ram_mem1_reg[234][12]/P0001 , \wishbone_bd_ram_mem1_reg[234][13]/P0001 , \wishbone_bd_ram_mem1_reg[234][14]/P0001 , \wishbone_bd_ram_mem1_reg[234][15]/P0001 , \wishbone_bd_ram_mem1_reg[234][8]/P0001 , \wishbone_bd_ram_mem1_reg[234][9]/P0001 , \wishbone_bd_ram_mem1_reg[235][10]/P0001 , \wishbone_bd_ram_mem1_reg[235][11]/P0001 , \wishbone_bd_ram_mem1_reg[235][12]/P0001 , \wishbone_bd_ram_mem1_reg[235][13]/P0001 , \wishbone_bd_ram_mem1_reg[235][14]/P0001 , \wishbone_bd_ram_mem1_reg[235][15]/P0001 , \wishbone_bd_ram_mem1_reg[235][8]/P0001 , \wishbone_bd_ram_mem1_reg[235][9]/P0001 , \wishbone_bd_ram_mem1_reg[236][10]/P0001 , \wishbone_bd_ram_mem1_reg[236][11]/P0001 , \wishbone_bd_ram_mem1_reg[236][12]/P0001 , \wishbone_bd_ram_mem1_reg[236][13]/P0001 , \wishbone_bd_ram_mem1_reg[236][14]/P0001 , \wishbone_bd_ram_mem1_reg[236][15]/P0001 , \wishbone_bd_ram_mem1_reg[236][8]/P0001 , \wishbone_bd_ram_mem1_reg[236][9]/P0001 , \wishbone_bd_ram_mem1_reg[237][10]/P0001 , \wishbone_bd_ram_mem1_reg[237][11]/P0001 , \wishbone_bd_ram_mem1_reg[237][12]/P0001 , \wishbone_bd_ram_mem1_reg[237][13]/P0001 , \wishbone_bd_ram_mem1_reg[237][14]/P0001 , \wishbone_bd_ram_mem1_reg[237][15]/P0001 , \wishbone_bd_ram_mem1_reg[237][8]/P0001 , \wishbone_bd_ram_mem1_reg[237][9]/P0001 , \wishbone_bd_ram_mem1_reg[238][10]/P0001 , \wishbone_bd_ram_mem1_reg[238][11]/P0001 , \wishbone_bd_ram_mem1_reg[238][12]/P0001 , \wishbone_bd_ram_mem1_reg[238][13]/P0001 , \wishbone_bd_ram_mem1_reg[238][14]/P0001 , \wishbone_bd_ram_mem1_reg[238][15]/P0001 , \wishbone_bd_ram_mem1_reg[238][8]/P0001 , \wishbone_bd_ram_mem1_reg[238][9]/P0001 , \wishbone_bd_ram_mem1_reg[239][10]/P0001 , \wishbone_bd_ram_mem1_reg[239][11]/P0001 , \wishbone_bd_ram_mem1_reg[239][12]/P0001 , \wishbone_bd_ram_mem1_reg[239][13]/P0001 , \wishbone_bd_ram_mem1_reg[239][14]/P0001 , \wishbone_bd_ram_mem1_reg[239][15]/P0001 , \wishbone_bd_ram_mem1_reg[239][8]/P0001 , \wishbone_bd_ram_mem1_reg[239][9]/P0001 , \wishbone_bd_ram_mem1_reg[23][10]/P0001 , \wishbone_bd_ram_mem1_reg[23][11]/P0001 , \wishbone_bd_ram_mem1_reg[23][12]/P0001 , \wishbone_bd_ram_mem1_reg[23][13]/P0001 , \wishbone_bd_ram_mem1_reg[23][14]/P0001 , \wishbone_bd_ram_mem1_reg[23][15]/P0001 , \wishbone_bd_ram_mem1_reg[23][8]/P0001 , \wishbone_bd_ram_mem1_reg[23][9]/P0001 , \wishbone_bd_ram_mem1_reg[240][10]/P0001 , \wishbone_bd_ram_mem1_reg[240][11]/P0001 , \wishbone_bd_ram_mem1_reg[240][12]/P0001 , \wishbone_bd_ram_mem1_reg[240][13]/P0001 , \wishbone_bd_ram_mem1_reg[240][14]/P0001 , \wishbone_bd_ram_mem1_reg[240][15]/P0001 , \wishbone_bd_ram_mem1_reg[240][8]/P0001 , \wishbone_bd_ram_mem1_reg[240][9]/P0001 , \wishbone_bd_ram_mem1_reg[241][10]/P0001 , \wishbone_bd_ram_mem1_reg[241][11]/P0001 , \wishbone_bd_ram_mem1_reg[241][12]/P0001 , \wishbone_bd_ram_mem1_reg[241][13]/P0001 , \wishbone_bd_ram_mem1_reg[241][14]/P0001 , \wishbone_bd_ram_mem1_reg[241][15]/P0001 , \wishbone_bd_ram_mem1_reg[241][8]/P0001 , \wishbone_bd_ram_mem1_reg[241][9]/P0001 , \wishbone_bd_ram_mem1_reg[242][10]/P0001 , \wishbone_bd_ram_mem1_reg[242][11]/P0001 , \wishbone_bd_ram_mem1_reg[242][12]/P0001 , \wishbone_bd_ram_mem1_reg[242][13]/P0001 , \wishbone_bd_ram_mem1_reg[242][14]/P0001 , \wishbone_bd_ram_mem1_reg[242][15]/P0001 , \wishbone_bd_ram_mem1_reg[242][8]/P0001 , \wishbone_bd_ram_mem1_reg[242][9]/P0001 , \wishbone_bd_ram_mem1_reg[243][10]/P0001 , \wishbone_bd_ram_mem1_reg[243][11]/P0001 , \wishbone_bd_ram_mem1_reg[243][12]/P0001 , \wishbone_bd_ram_mem1_reg[243][13]/P0001 , \wishbone_bd_ram_mem1_reg[243][14]/P0001 , \wishbone_bd_ram_mem1_reg[243][15]/P0001 , \wishbone_bd_ram_mem1_reg[243][8]/P0001 , \wishbone_bd_ram_mem1_reg[243][9]/P0001 , \wishbone_bd_ram_mem1_reg[244][10]/P0001 , \wishbone_bd_ram_mem1_reg[244][11]/P0001 , \wishbone_bd_ram_mem1_reg[244][12]/P0001 , \wishbone_bd_ram_mem1_reg[244][13]/P0001 , \wishbone_bd_ram_mem1_reg[244][14]/P0001 , \wishbone_bd_ram_mem1_reg[244][15]/P0001 , \wishbone_bd_ram_mem1_reg[244][8]/P0001 , \wishbone_bd_ram_mem1_reg[244][9]/P0001 , \wishbone_bd_ram_mem1_reg[245][10]/P0001 , \wishbone_bd_ram_mem1_reg[245][11]/P0001 , \wishbone_bd_ram_mem1_reg[245][12]/P0001 , \wishbone_bd_ram_mem1_reg[245][13]/P0001 , \wishbone_bd_ram_mem1_reg[245][14]/P0001 , \wishbone_bd_ram_mem1_reg[245][15]/P0001 , \wishbone_bd_ram_mem1_reg[245][8]/P0001 , \wishbone_bd_ram_mem1_reg[245][9]/P0001 , \wishbone_bd_ram_mem1_reg[246][10]/P0001 , \wishbone_bd_ram_mem1_reg[246][11]/P0001 , \wishbone_bd_ram_mem1_reg[246][12]/P0001 , \wishbone_bd_ram_mem1_reg[246][13]/P0001 , \wishbone_bd_ram_mem1_reg[246][14]/P0001 , \wishbone_bd_ram_mem1_reg[246][15]/P0001 , \wishbone_bd_ram_mem1_reg[246][8]/P0001 , \wishbone_bd_ram_mem1_reg[246][9]/P0001 , \wishbone_bd_ram_mem1_reg[247][10]/P0001 , \wishbone_bd_ram_mem1_reg[247][11]/P0001 , \wishbone_bd_ram_mem1_reg[247][12]/P0001 , \wishbone_bd_ram_mem1_reg[247][13]/P0001 , \wishbone_bd_ram_mem1_reg[247][14]/P0001 , \wishbone_bd_ram_mem1_reg[247][15]/P0001 , \wishbone_bd_ram_mem1_reg[247][8]/P0001 , \wishbone_bd_ram_mem1_reg[247][9]/P0001 , \wishbone_bd_ram_mem1_reg[248][10]/P0001 , \wishbone_bd_ram_mem1_reg[248][11]/P0001 , \wishbone_bd_ram_mem1_reg[248][12]/P0001 , \wishbone_bd_ram_mem1_reg[248][13]/P0001 , \wishbone_bd_ram_mem1_reg[248][14]/P0001 , \wishbone_bd_ram_mem1_reg[248][15]/P0001 , \wishbone_bd_ram_mem1_reg[248][8]/P0001 , \wishbone_bd_ram_mem1_reg[248][9]/P0001 , \wishbone_bd_ram_mem1_reg[249][10]/P0001 , \wishbone_bd_ram_mem1_reg[249][11]/P0001 , \wishbone_bd_ram_mem1_reg[249][12]/P0001 , \wishbone_bd_ram_mem1_reg[249][13]/P0001 , \wishbone_bd_ram_mem1_reg[249][14]/P0001 , \wishbone_bd_ram_mem1_reg[249][15]/P0001 , \wishbone_bd_ram_mem1_reg[249][8]/P0001 , \wishbone_bd_ram_mem1_reg[249][9]/P0001 , \wishbone_bd_ram_mem1_reg[24][10]/P0001 , \wishbone_bd_ram_mem1_reg[24][11]/P0001 , \wishbone_bd_ram_mem1_reg[24][12]/P0001 , \wishbone_bd_ram_mem1_reg[24][13]/P0001 , \wishbone_bd_ram_mem1_reg[24][14]/P0001 , \wishbone_bd_ram_mem1_reg[24][15]/P0001 , \wishbone_bd_ram_mem1_reg[24][8]/P0001 , \wishbone_bd_ram_mem1_reg[24][9]/P0001 , \wishbone_bd_ram_mem1_reg[250][10]/P0001 , \wishbone_bd_ram_mem1_reg[250][11]/P0001 , \wishbone_bd_ram_mem1_reg[250][12]/P0001 , \wishbone_bd_ram_mem1_reg[250][13]/P0001 , \wishbone_bd_ram_mem1_reg[250][14]/P0001 , \wishbone_bd_ram_mem1_reg[250][15]/P0001 , \wishbone_bd_ram_mem1_reg[250][8]/P0001 , \wishbone_bd_ram_mem1_reg[250][9]/P0001 , \wishbone_bd_ram_mem1_reg[251][10]/P0001 , \wishbone_bd_ram_mem1_reg[251][11]/P0001 , \wishbone_bd_ram_mem1_reg[251][12]/P0001 , \wishbone_bd_ram_mem1_reg[251][13]/P0001 , \wishbone_bd_ram_mem1_reg[251][14]/P0001 , \wishbone_bd_ram_mem1_reg[251][15]/P0001 , \wishbone_bd_ram_mem1_reg[251][8]/P0001 , \wishbone_bd_ram_mem1_reg[251][9]/P0001 , \wishbone_bd_ram_mem1_reg[252][10]/P0001 , \wishbone_bd_ram_mem1_reg[252][11]/P0001 , \wishbone_bd_ram_mem1_reg[252][12]/P0001 , \wishbone_bd_ram_mem1_reg[252][13]/P0001 , \wishbone_bd_ram_mem1_reg[252][14]/P0001 , \wishbone_bd_ram_mem1_reg[252][15]/P0001 , \wishbone_bd_ram_mem1_reg[252][8]/P0001 , \wishbone_bd_ram_mem1_reg[252][9]/P0001 , \wishbone_bd_ram_mem1_reg[253][10]/P0001 , \wishbone_bd_ram_mem1_reg[253][11]/P0001 , \wishbone_bd_ram_mem1_reg[253][12]/P0001 , \wishbone_bd_ram_mem1_reg[253][13]/P0001 , \wishbone_bd_ram_mem1_reg[253][14]/P0001 , \wishbone_bd_ram_mem1_reg[253][15]/P0001 , \wishbone_bd_ram_mem1_reg[253][8]/P0001 , \wishbone_bd_ram_mem1_reg[253][9]/P0001 , \wishbone_bd_ram_mem1_reg[254][10]/P0001 , \wishbone_bd_ram_mem1_reg[254][11]/P0001 , \wishbone_bd_ram_mem1_reg[254][12]/P0001 , \wishbone_bd_ram_mem1_reg[254][13]/P0001 , \wishbone_bd_ram_mem1_reg[254][14]/P0001 , \wishbone_bd_ram_mem1_reg[254][15]/P0001 , \wishbone_bd_ram_mem1_reg[254][8]/P0001 , \wishbone_bd_ram_mem1_reg[254][9]/P0001 , \wishbone_bd_ram_mem1_reg[255][10]/P0001 , \wishbone_bd_ram_mem1_reg[255][11]/P0001 , \wishbone_bd_ram_mem1_reg[255][12]/P0001 , \wishbone_bd_ram_mem1_reg[255][13]/P0001 , \wishbone_bd_ram_mem1_reg[255][14]/P0001 , \wishbone_bd_ram_mem1_reg[255][15]/P0001 , \wishbone_bd_ram_mem1_reg[255][8]/P0001 , \wishbone_bd_ram_mem1_reg[255][9]/P0001 , \wishbone_bd_ram_mem1_reg[25][10]/P0001 , \wishbone_bd_ram_mem1_reg[25][11]/P0001 , \wishbone_bd_ram_mem1_reg[25][12]/P0001 , \wishbone_bd_ram_mem1_reg[25][13]/P0001 , \wishbone_bd_ram_mem1_reg[25][14]/P0001 , \wishbone_bd_ram_mem1_reg[25][15]/P0001 , \wishbone_bd_ram_mem1_reg[25][8]/P0001 , \wishbone_bd_ram_mem1_reg[25][9]/P0001 , \wishbone_bd_ram_mem1_reg[26][10]/P0001 , \wishbone_bd_ram_mem1_reg[26][11]/P0001 , \wishbone_bd_ram_mem1_reg[26][12]/P0001 , \wishbone_bd_ram_mem1_reg[26][13]/P0001 , \wishbone_bd_ram_mem1_reg[26][14]/P0001 , \wishbone_bd_ram_mem1_reg[26][15]/P0001 , \wishbone_bd_ram_mem1_reg[26][8]/P0001 , \wishbone_bd_ram_mem1_reg[26][9]/P0001 , \wishbone_bd_ram_mem1_reg[27][10]/P0001 , \wishbone_bd_ram_mem1_reg[27][11]/P0001 , \wishbone_bd_ram_mem1_reg[27][12]/P0001 , \wishbone_bd_ram_mem1_reg[27][13]/P0001 , \wishbone_bd_ram_mem1_reg[27][14]/P0001 , \wishbone_bd_ram_mem1_reg[27][15]/P0001 , \wishbone_bd_ram_mem1_reg[27][8]/P0001 , \wishbone_bd_ram_mem1_reg[27][9]/P0001 , \wishbone_bd_ram_mem1_reg[28][10]/P0001 , \wishbone_bd_ram_mem1_reg[28][11]/P0001 , \wishbone_bd_ram_mem1_reg[28][12]/P0001 , \wishbone_bd_ram_mem1_reg[28][13]/P0001 , \wishbone_bd_ram_mem1_reg[28][14]/P0001 , \wishbone_bd_ram_mem1_reg[28][15]/P0001 , \wishbone_bd_ram_mem1_reg[28][8]/P0001 , \wishbone_bd_ram_mem1_reg[28][9]/P0001 , \wishbone_bd_ram_mem1_reg[29][10]/P0001 , \wishbone_bd_ram_mem1_reg[29][11]/P0001 , \wishbone_bd_ram_mem1_reg[29][12]/P0001 , \wishbone_bd_ram_mem1_reg[29][13]/P0001 , \wishbone_bd_ram_mem1_reg[29][14]/P0001 , \wishbone_bd_ram_mem1_reg[29][15]/P0001 , \wishbone_bd_ram_mem1_reg[29][8]/P0001 , \wishbone_bd_ram_mem1_reg[29][9]/P0001 , \wishbone_bd_ram_mem1_reg[2][10]/P0001 , \wishbone_bd_ram_mem1_reg[2][11]/P0001 , \wishbone_bd_ram_mem1_reg[2][12]/P0001 , \wishbone_bd_ram_mem1_reg[2][13]/P0001 , \wishbone_bd_ram_mem1_reg[2][14]/P0001 , \wishbone_bd_ram_mem1_reg[2][15]/P0001 , \wishbone_bd_ram_mem1_reg[2][8]/P0001 , \wishbone_bd_ram_mem1_reg[2][9]/P0001 , \wishbone_bd_ram_mem1_reg[30][10]/P0001 , \wishbone_bd_ram_mem1_reg[30][11]/P0001 , \wishbone_bd_ram_mem1_reg[30][12]/P0001 , \wishbone_bd_ram_mem1_reg[30][13]/P0001 , \wishbone_bd_ram_mem1_reg[30][14]/P0001 , \wishbone_bd_ram_mem1_reg[30][15]/P0001 , \wishbone_bd_ram_mem1_reg[30][8]/P0001 , \wishbone_bd_ram_mem1_reg[30][9]/P0001 , \wishbone_bd_ram_mem1_reg[31][10]/P0001 , \wishbone_bd_ram_mem1_reg[31][11]/P0001 , \wishbone_bd_ram_mem1_reg[31][12]/P0001 , \wishbone_bd_ram_mem1_reg[31][13]/P0001 , \wishbone_bd_ram_mem1_reg[31][14]/P0001 , \wishbone_bd_ram_mem1_reg[31][15]/P0001 , \wishbone_bd_ram_mem1_reg[31][8]/P0001 , \wishbone_bd_ram_mem1_reg[31][9]/P0001 , \wishbone_bd_ram_mem1_reg[32][10]/P0001 , \wishbone_bd_ram_mem1_reg[32][11]/P0001 , \wishbone_bd_ram_mem1_reg[32][12]/P0001 , \wishbone_bd_ram_mem1_reg[32][13]/P0001 , \wishbone_bd_ram_mem1_reg[32][14]/P0001 , \wishbone_bd_ram_mem1_reg[32][15]/P0001 , \wishbone_bd_ram_mem1_reg[32][8]/P0001 , \wishbone_bd_ram_mem1_reg[32][9]/P0001 , \wishbone_bd_ram_mem1_reg[33][10]/P0001 , \wishbone_bd_ram_mem1_reg[33][11]/P0001 , \wishbone_bd_ram_mem1_reg[33][12]/P0001 , \wishbone_bd_ram_mem1_reg[33][13]/P0001 , \wishbone_bd_ram_mem1_reg[33][14]/P0001 , \wishbone_bd_ram_mem1_reg[33][15]/P0001 , \wishbone_bd_ram_mem1_reg[33][8]/P0001 , \wishbone_bd_ram_mem1_reg[33][9]/P0001 , \wishbone_bd_ram_mem1_reg[34][10]/P0001 , \wishbone_bd_ram_mem1_reg[34][11]/P0001 , \wishbone_bd_ram_mem1_reg[34][12]/P0001 , \wishbone_bd_ram_mem1_reg[34][13]/P0001 , \wishbone_bd_ram_mem1_reg[34][14]/P0001 , \wishbone_bd_ram_mem1_reg[34][15]/P0001 , \wishbone_bd_ram_mem1_reg[34][8]/P0001 , \wishbone_bd_ram_mem1_reg[34][9]/P0001 , \wishbone_bd_ram_mem1_reg[35][10]/P0001 , \wishbone_bd_ram_mem1_reg[35][11]/P0001 , \wishbone_bd_ram_mem1_reg[35][12]/P0001 , \wishbone_bd_ram_mem1_reg[35][13]/P0001 , \wishbone_bd_ram_mem1_reg[35][14]/P0001 , \wishbone_bd_ram_mem1_reg[35][15]/P0001 , \wishbone_bd_ram_mem1_reg[35][8]/P0001 , \wishbone_bd_ram_mem1_reg[35][9]/P0001 , \wishbone_bd_ram_mem1_reg[36][10]/P0001 , \wishbone_bd_ram_mem1_reg[36][11]/P0001 , \wishbone_bd_ram_mem1_reg[36][12]/P0001 , \wishbone_bd_ram_mem1_reg[36][13]/P0001 , \wishbone_bd_ram_mem1_reg[36][14]/P0001 , \wishbone_bd_ram_mem1_reg[36][15]/P0001 , \wishbone_bd_ram_mem1_reg[36][8]/P0001 , \wishbone_bd_ram_mem1_reg[36][9]/P0001 , \wishbone_bd_ram_mem1_reg[37][10]/P0001 , \wishbone_bd_ram_mem1_reg[37][11]/P0001 , \wishbone_bd_ram_mem1_reg[37][12]/P0001 , \wishbone_bd_ram_mem1_reg[37][13]/P0001 , \wishbone_bd_ram_mem1_reg[37][14]/P0001 , \wishbone_bd_ram_mem1_reg[37][15]/P0001 , \wishbone_bd_ram_mem1_reg[37][8]/P0001 , \wishbone_bd_ram_mem1_reg[37][9]/P0001 , \wishbone_bd_ram_mem1_reg[38][10]/P0001 , \wishbone_bd_ram_mem1_reg[38][11]/P0001 , \wishbone_bd_ram_mem1_reg[38][12]/P0001 , \wishbone_bd_ram_mem1_reg[38][13]/P0001 , \wishbone_bd_ram_mem1_reg[38][14]/P0001 , \wishbone_bd_ram_mem1_reg[38][15]/P0001 , \wishbone_bd_ram_mem1_reg[38][8]/P0001 , \wishbone_bd_ram_mem1_reg[38][9]/P0001 , \wishbone_bd_ram_mem1_reg[39][10]/P0001 , \wishbone_bd_ram_mem1_reg[39][11]/P0001 , \wishbone_bd_ram_mem1_reg[39][12]/P0001 , \wishbone_bd_ram_mem1_reg[39][13]/P0001 , \wishbone_bd_ram_mem1_reg[39][14]/P0001 , \wishbone_bd_ram_mem1_reg[39][15]/P0001 , \wishbone_bd_ram_mem1_reg[39][8]/P0001 , \wishbone_bd_ram_mem1_reg[39][9]/P0001 , \wishbone_bd_ram_mem1_reg[3][10]/P0001 , \wishbone_bd_ram_mem1_reg[3][11]/P0001 , \wishbone_bd_ram_mem1_reg[3][12]/P0001 , \wishbone_bd_ram_mem1_reg[3][13]/P0001 , \wishbone_bd_ram_mem1_reg[3][14]/P0001 , \wishbone_bd_ram_mem1_reg[3][15]/P0001 , \wishbone_bd_ram_mem1_reg[3][8]/P0001 , \wishbone_bd_ram_mem1_reg[3][9]/P0001 , \wishbone_bd_ram_mem1_reg[40][10]/P0001 , \wishbone_bd_ram_mem1_reg[40][11]/P0001 , \wishbone_bd_ram_mem1_reg[40][12]/P0001 , \wishbone_bd_ram_mem1_reg[40][13]/P0001 , \wishbone_bd_ram_mem1_reg[40][14]/P0001 , \wishbone_bd_ram_mem1_reg[40][15]/P0001 , \wishbone_bd_ram_mem1_reg[40][8]/P0001 , \wishbone_bd_ram_mem1_reg[40][9]/P0001 , \wishbone_bd_ram_mem1_reg[41][10]/P0001 , \wishbone_bd_ram_mem1_reg[41][11]/P0001 , \wishbone_bd_ram_mem1_reg[41][12]/P0001 , \wishbone_bd_ram_mem1_reg[41][13]/P0001 , \wishbone_bd_ram_mem1_reg[41][14]/P0001 , \wishbone_bd_ram_mem1_reg[41][15]/P0001 , \wishbone_bd_ram_mem1_reg[41][8]/P0001 , \wishbone_bd_ram_mem1_reg[41][9]/P0001 , \wishbone_bd_ram_mem1_reg[42][10]/P0001 , \wishbone_bd_ram_mem1_reg[42][11]/P0001 , \wishbone_bd_ram_mem1_reg[42][12]/P0001 , \wishbone_bd_ram_mem1_reg[42][13]/P0001 , \wishbone_bd_ram_mem1_reg[42][14]/P0001 , \wishbone_bd_ram_mem1_reg[42][15]/P0001 , \wishbone_bd_ram_mem1_reg[42][8]/P0001 , \wishbone_bd_ram_mem1_reg[42][9]/P0001 , \wishbone_bd_ram_mem1_reg[43][10]/P0001 , \wishbone_bd_ram_mem1_reg[43][11]/P0001 , \wishbone_bd_ram_mem1_reg[43][12]/P0001 , \wishbone_bd_ram_mem1_reg[43][13]/P0001 , \wishbone_bd_ram_mem1_reg[43][14]/P0001 , \wishbone_bd_ram_mem1_reg[43][15]/P0001 , \wishbone_bd_ram_mem1_reg[43][8]/P0001 , \wishbone_bd_ram_mem1_reg[43][9]/P0001 , \wishbone_bd_ram_mem1_reg[44][10]/P0001 , \wishbone_bd_ram_mem1_reg[44][11]/P0001 , \wishbone_bd_ram_mem1_reg[44][12]/P0001 , \wishbone_bd_ram_mem1_reg[44][13]/P0001 , \wishbone_bd_ram_mem1_reg[44][14]/P0001 , \wishbone_bd_ram_mem1_reg[44][15]/P0001 , \wishbone_bd_ram_mem1_reg[44][8]/P0001 , \wishbone_bd_ram_mem1_reg[44][9]/P0001 , \wishbone_bd_ram_mem1_reg[45][10]/P0001 , \wishbone_bd_ram_mem1_reg[45][11]/P0001 , \wishbone_bd_ram_mem1_reg[45][12]/P0001 , \wishbone_bd_ram_mem1_reg[45][13]/P0001 , \wishbone_bd_ram_mem1_reg[45][14]/P0001 , \wishbone_bd_ram_mem1_reg[45][15]/P0001 , \wishbone_bd_ram_mem1_reg[45][8]/P0001 , \wishbone_bd_ram_mem1_reg[45][9]/P0001 , \wishbone_bd_ram_mem1_reg[46][10]/P0001 , \wishbone_bd_ram_mem1_reg[46][11]/P0001 , \wishbone_bd_ram_mem1_reg[46][12]/P0001 , \wishbone_bd_ram_mem1_reg[46][13]/P0001 , \wishbone_bd_ram_mem1_reg[46][14]/P0001 , \wishbone_bd_ram_mem1_reg[46][15]/P0001 , \wishbone_bd_ram_mem1_reg[46][8]/P0001 , \wishbone_bd_ram_mem1_reg[46][9]/P0001 , \wishbone_bd_ram_mem1_reg[47][10]/P0001 , \wishbone_bd_ram_mem1_reg[47][11]/P0001 , \wishbone_bd_ram_mem1_reg[47][12]/P0001 , \wishbone_bd_ram_mem1_reg[47][13]/P0001 , \wishbone_bd_ram_mem1_reg[47][14]/P0001 , \wishbone_bd_ram_mem1_reg[47][15]/P0001 , \wishbone_bd_ram_mem1_reg[47][8]/P0001 , \wishbone_bd_ram_mem1_reg[47][9]/P0001 , \wishbone_bd_ram_mem1_reg[48][10]/P0001 , \wishbone_bd_ram_mem1_reg[48][11]/P0001 , \wishbone_bd_ram_mem1_reg[48][12]/P0001 , \wishbone_bd_ram_mem1_reg[48][13]/P0001 , \wishbone_bd_ram_mem1_reg[48][14]/P0001 , \wishbone_bd_ram_mem1_reg[48][15]/P0001 , \wishbone_bd_ram_mem1_reg[48][8]/P0001 , \wishbone_bd_ram_mem1_reg[48][9]/P0001 , \wishbone_bd_ram_mem1_reg[49][10]/P0001 , \wishbone_bd_ram_mem1_reg[49][11]/P0001 , \wishbone_bd_ram_mem1_reg[49][12]/P0001 , \wishbone_bd_ram_mem1_reg[49][13]/P0001 , \wishbone_bd_ram_mem1_reg[49][14]/P0001 , \wishbone_bd_ram_mem1_reg[49][15]/P0001 , \wishbone_bd_ram_mem1_reg[49][8]/P0001 , \wishbone_bd_ram_mem1_reg[49][9]/P0001 , \wishbone_bd_ram_mem1_reg[4][10]/P0001 , \wishbone_bd_ram_mem1_reg[4][11]/P0001 , \wishbone_bd_ram_mem1_reg[4][12]/P0001 , \wishbone_bd_ram_mem1_reg[4][13]/P0001 , \wishbone_bd_ram_mem1_reg[4][14]/P0001 , \wishbone_bd_ram_mem1_reg[4][15]/P0001 , \wishbone_bd_ram_mem1_reg[4][8]/P0001 , \wishbone_bd_ram_mem1_reg[4][9]/P0001 , \wishbone_bd_ram_mem1_reg[50][10]/P0001 , \wishbone_bd_ram_mem1_reg[50][11]/P0001 , \wishbone_bd_ram_mem1_reg[50][12]/P0001 , \wishbone_bd_ram_mem1_reg[50][13]/P0001 , \wishbone_bd_ram_mem1_reg[50][14]/P0001 , \wishbone_bd_ram_mem1_reg[50][15]/P0001 , \wishbone_bd_ram_mem1_reg[50][8]/P0001 , \wishbone_bd_ram_mem1_reg[50][9]/P0001 , \wishbone_bd_ram_mem1_reg[51][10]/P0001 , \wishbone_bd_ram_mem1_reg[51][11]/P0001 , \wishbone_bd_ram_mem1_reg[51][12]/P0001 , \wishbone_bd_ram_mem1_reg[51][13]/P0001 , \wishbone_bd_ram_mem1_reg[51][14]/P0001 , \wishbone_bd_ram_mem1_reg[51][15]/P0001 , \wishbone_bd_ram_mem1_reg[51][8]/P0001 , \wishbone_bd_ram_mem1_reg[51][9]/P0001 , \wishbone_bd_ram_mem1_reg[52][10]/P0001 , \wishbone_bd_ram_mem1_reg[52][11]/P0001 , \wishbone_bd_ram_mem1_reg[52][12]/P0001 , \wishbone_bd_ram_mem1_reg[52][13]/P0001 , \wishbone_bd_ram_mem1_reg[52][14]/P0001 , \wishbone_bd_ram_mem1_reg[52][15]/P0001 , \wishbone_bd_ram_mem1_reg[52][8]/P0001 , \wishbone_bd_ram_mem1_reg[52][9]/P0001 , \wishbone_bd_ram_mem1_reg[53][10]/P0001 , \wishbone_bd_ram_mem1_reg[53][11]/P0001 , \wishbone_bd_ram_mem1_reg[53][12]/P0001 , \wishbone_bd_ram_mem1_reg[53][13]/P0001 , \wishbone_bd_ram_mem1_reg[53][14]/P0001 , \wishbone_bd_ram_mem1_reg[53][15]/P0001 , \wishbone_bd_ram_mem1_reg[53][8]/P0001 , \wishbone_bd_ram_mem1_reg[53][9]/P0001 , \wishbone_bd_ram_mem1_reg[54][10]/P0001 , \wishbone_bd_ram_mem1_reg[54][11]/P0001 , \wishbone_bd_ram_mem1_reg[54][12]/P0001 , \wishbone_bd_ram_mem1_reg[54][13]/P0001 , \wishbone_bd_ram_mem1_reg[54][14]/P0001 , \wishbone_bd_ram_mem1_reg[54][15]/P0001 , \wishbone_bd_ram_mem1_reg[54][8]/P0001 , \wishbone_bd_ram_mem1_reg[54][9]/P0001 , \wishbone_bd_ram_mem1_reg[55][10]/P0001 , \wishbone_bd_ram_mem1_reg[55][11]/P0001 , \wishbone_bd_ram_mem1_reg[55][12]/P0001 , \wishbone_bd_ram_mem1_reg[55][13]/P0001 , \wishbone_bd_ram_mem1_reg[55][14]/P0001 , \wishbone_bd_ram_mem1_reg[55][15]/P0001 , \wishbone_bd_ram_mem1_reg[55][8]/P0001 , \wishbone_bd_ram_mem1_reg[55][9]/P0001 , \wishbone_bd_ram_mem1_reg[56][10]/P0001 , \wishbone_bd_ram_mem1_reg[56][11]/P0001 , \wishbone_bd_ram_mem1_reg[56][12]/P0001 , \wishbone_bd_ram_mem1_reg[56][13]/P0001 , \wishbone_bd_ram_mem1_reg[56][14]/P0001 , \wishbone_bd_ram_mem1_reg[56][15]/P0001 , \wishbone_bd_ram_mem1_reg[56][8]/P0001 , \wishbone_bd_ram_mem1_reg[56][9]/P0001 , \wishbone_bd_ram_mem1_reg[57][10]/P0001 , \wishbone_bd_ram_mem1_reg[57][11]/P0001 , \wishbone_bd_ram_mem1_reg[57][12]/P0001 , \wishbone_bd_ram_mem1_reg[57][13]/P0001 , \wishbone_bd_ram_mem1_reg[57][14]/P0001 , \wishbone_bd_ram_mem1_reg[57][15]/P0001 , \wishbone_bd_ram_mem1_reg[57][8]/P0001 , \wishbone_bd_ram_mem1_reg[57][9]/P0001 , \wishbone_bd_ram_mem1_reg[58][10]/P0001 , \wishbone_bd_ram_mem1_reg[58][11]/P0001 , \wishbone_bd_ram_mem1_reg[58][12]/P0001 , \wishbone_bd_ram_mem1_reg[58][13]/P0001 , \wishbone_bd_ram_mem1_reg[58][14]/P0001 , \wishbone_bd_ram_mem1_reg[58][15]/P0001 , \wishbone_bd_ram_mem1_reg[58][8]/P0001 , \wishbone_bd_ram_mem1_reg[58][9]/P0001 , \wishbone_bd_ram_mem1_reg[59][10]/P0001 , \wishbone_bd_ram_mem1_reg[59][11]/P0001 , \wishbone_bd_ram_mem1_reg[59][12]/P0001 , \wishbone_bd_ram_mem1_reg[59][13]/P0001 , \wishbone_bd_ram_mem1_reg[59][14]/P0001 , \wishbone_bd_ram_mem1_reg[59][15]/P0001 , \wishbone_bd_ram_mem1_reg[59][8]/P0001 , \wishbone_bd_ram_mem1_reg[59][9]/P0001 , \wishbone_bd_ram_mem1_reg[5][10]/P0001 , \wishbone_bd_ram_mem1_reg[5][11]/P0001 , \wishbone_bd_ram_mem1_reg[5][12]/P0001 , \wishbone_bd_ram_mem1_reg[5][13]/P0001 , \wishbone_bd_ram_mem1_reg[5][14]/P0001 , \wishbone_bd_ram_mem1_reg[5][15]/P0001 , \wishbone_bd_ram_mem1_reg[5][8]/P0001 , \wishbone_bd_ram_mem1_reg[5][9]/P0001 , \wishbone_bd_ram_mem1_reg[60][10]/P0001 , \wishbone_bd_ram_mem1_reg[60][11]/P0001 , \wishbone_bd_ram_mem1_reg[60][12]/P0001 , \wishbone_bd_ram_mem1_reg[60][13]/P0001 , \wishbone_bd_ram_mem1_reg[60][14]/P0001 , \wishbone_bd_ram_mem1_reg[60][15]/P0001 , \wishbone_bd_ram_mem1_reg[60][8]/P0001 , \wishbone_bd_ram_mem1_reg[60][9]/P0001 , \wishbone_bd_ram_mem1_reg[61][10]/P0001 , \wishbone_bd_ram_mem1_reg[61][11]/P0001 , \wishbone_bd_ram_mem1_reg[61][12]/P0001 , \wishbone_bd_ram_mem1_reg[61][13]/P0001 , \wishbone_bd_ram_mem1_reg[61][14]/P0001 , \wishbone_bd_ram_mem1_reg[61][15]/P0001 , \wishbone_bd_ram_mem1_reg[61][8]/P0001 , \wishbone_bd_ram_mem1_reg[61][9]/P0001 , \wishbone_bd_ram_mem1_reg[62][10]/P0001 , \wishbone_bd_ram_mem1_reg[62][11]/P0001 , \wishbone_bd_ram_mem1_reg[62][12]/P0001 , \wishbone_bd_ram_mem1_reg[62][13]/P0001 , \wishbone_bd_ram_mem1_reg[62][14]/P0001 , \wishbone_bd_ram_mem1_reg[62][15]/P0001 , \wishbone_bd_ram_mem1_reg[62][8]/P0001 , \wishbone_bd_ram_mem1_reg[62][9]/P0001 , \wishbone_bd_ram_mem1_reg[63][10]/P0001 , \wishbone_bd_ram_mem1_reg[63][11]/P0001 , \wishbone_bd_ram_mem1_reg[63][12]/P0001 , \wishbone_bd_ram_mem1_reg[63][13]/P0001 , \wishbone_bd_ram_mem1_reg[63][14]/P0001 , \wishbone_bd_ram_mem1_reg[63][15]/P0001 , \wishbone_bd_ram_mem1_reg[63][8]/P0001 , \wishbone_bd_ram_mem1_reg[63][9]/P0001 , \wishbone_bd_ram_mem1_reg[64][10]/P0001 , \wishbone_bd_ram_mem1_reg[64][11]/P0001 , \wishbone_bd_ram_mem1_reg[64][12]/P0001 , \wishbone_bd_ram_mem1_reg[64][13]/P0001 , \wishbone_bd_ram_mem1_reg[64][14]/P0001 , \wishbone_bd_ram_mem1_reg[64][15]/P0001 , \wishbone_bd_ram_mem1_reg[64][8]/P0001 , \wishbone_bd_ram_mem1_reg[64][9]/P0001 , \wishbone_bd_ram_mem1_reg[65][10]/P0001 , \wishbone_bd_ram_mem1_reg[65][11]/P0001 , \wishbone_bd_ram_mem1_reg[65][12]/P0001 , \wishbone_bd_ram_mem1_reg[65][13]/P0001 , \wishbone_bd_ram_mem1_reg[65][14]/P0001 , \wishbone_bd_ram_mem1_reg[65][15]/P0001 , \wishbone_bd_ram_mem1_reg[65][8]/P0001 , \wishbone_bd_ram_mem1_reg[65][9]/P0001 , \wishbone_bd_ram_mem1_reg[66][10]/P0001 , \wishbone_bd_ram_mem1_reg[66][11]/P0001 , \wishbone_bd_ram_mem1_reg[66][12]/P0001 , \wishbone_bd_ram_mem1_reg[66][13]/P0001 , \wishbone_bd_ram_mem1_reg[66][14]/P0001 , \wishbone_bd_ram_mem1_reg[66][15]/P0001 , \wishbone_bd_ram_mem1_reg[66][8]/P0001 , \wishbone_bd_ram_mem1_reg[66][9]/P0001 , \wishbone_bd_ram_mem1_reg[67][10]/P0001 , \wishbone_bd_ram_mem1_reg[67][11]/P0001 , \wishbone_bd_ram_mem1_reg[67][12]/P0001 , \wishbone_bd_ram_mem1_reg[67][13]/P0001 , \wishbone_bd_ram_mem1_reg[67][14]/P0001 , \wishbone_bd_ram_mem1_reg[67][15]/P0001 , \wishbone_bd_ram_mem1_reg[67][8]/P0001 , \wishbone_bd_ram_mem1_reg[67][9]/P0001 , \wishbone_bd_ram_mem1_reg[68][10]/P0001 , \wishbone_bd_ram_mem1_reg[68][11]/P0001 , \wishbone_bd_ram_mem1_reg[68][12]/P0001 , \wishbone_bd_ram_mem1_reg[68][13]/P0001 , \wishbone_bd_ram_mem1_reg[68][14]/P0001 , \wishbone_bd_ram_mem1_reg[68][15]/P0001 , \wishbone_bd_ram_mem1_reg[68][8]/P0001 , \wishbone_bd_ram_mem1_reg[68][9]/P0001 , \wishbone_bd_ram_mem1_reg[69][10]/P0001 , \wishbone_bd_ram_mem1_reg[69][11]/P0001 , \wishbone_bd_ram_mem1_reg[69][12]/P0001 , \wishbone_bd_ram_mem1_reg[69][13]/P0001 , \wishbone_bd_ram_mem1_reg[69][14]/P0001 , \wishbone_bd_ram_mem1_reg[69][15]/P0001 , \wishbone_bd_ram_mem1_reg[69][8]/P0001 , \wishbone_bd_ram_mem1_reg[69][9]/P0001 , \wishbone_bd_ram_mem1_reg[6][10]/P0001 , \wishbone_bd_ram_mem1_reg[6][11]/P0001 , \wishbone_bd_ram_mem1_reg[6][12]/P0001 , \wishbone_bd_ram_mem1_reg[6][13]/P0001 , \wishbone_bd_ram_mem1_reg[6][14]/P0001 , \wishbone_bd_ram_mem1_reg[6][15]/P0001 , \wishbone_bd_ram_mem1_reg[6][8]/P0001 , \wishbone_bd_ram_mem1_reg[6][9]/P0001 , \wishbone_bd_ram_mem1_reg[70][10]/P0001 , \wishbone_bd_ram_mem1_reg[70][11]/P0001 , \wishbone_bd_ram_mem1_reg[70][12]/P0001 , \wishbone_bd_ram_mem1_reg[70][13]/P0001 , \wishbone_bd_ram_mem1_reg[70][14]/P0001 , \wishbone_bd_ram_mem1_reg[70][15]/P0001 , \wishbone_bd_ram_mem1_reg[70][8]/P0001 , \wishbone_bd_ram_mem1_reg[70][9]/P0001 , \wishbone_bd_ram_mem1_reg[71][10]/P0001 , \wishbone_bd_ram_mem1_reg[71][11]/P0001 , \wishbone_bd_ram_mem1_reg[71][12]/P0001 , \wishbone_bd_ram_mem1_reg[71][13]/P0001 , \wishbone_bd_ram_mem1_reg[71][14]/P0001 , \wishbone_bd_ram_mem1_reg[71][15]/P0001 , \wishbone_bd_ram_mem1_reg[71][8]/P0001 , \wishbone_bd_ram_mem1_reg[71][9]/P0001 , \wishbone_bd_ram_mem1_reg[72][10]/P0001 , \wishbone_bd_ram_mem1_reg[72][11]/P0001 , \wishbone_bd_ram_mem1_reg[72][12]/P0001 , \wishbone_bd_ram_mem1_reg[72][13]/P0001 , \wishbone_bd_ram_mem1_reg[72][14]/P0001 , \wishbone_bd_ram_mem1_reg[72][15]/P0001 , \wishbone_bd_ram_mem1_reg[72][8]/P0001 , \wishbone_bd_ram_mem1_reg[72][9]/P0001 , \wishbone_bd_ram_mem1_reg[73][10]/P0001 , \wishbone_bd_ram_mem1_reg[73][11]/P0001 , \wishbone_bd_ram_mem1_reg[73][12]/P0001 , \wishbone_bd_ram_mem1_reg[73][13]/P0001 , \wishbone_bd_ram_mem1_reg[73][14]/P0001 , \wishbone_bd_ram_mem1_reg[73][15]/P0001 , \wishbone_bd_ram_mem1_reg[73][8]/P0001 , \wishbone_bd_ram_mem1_reg[73][9]/P0001 , \wishbone_bd_ram_mem1_reg[74][10]/P0001 , \wishbone_bd_ram_mem1_reg[74][11]/P0001 , \wishbone_bd_ram_mem1_reg[74][12]/P0001 , \wishbone_bd_ram_mem1_reg[74][13]/P0001 , \wishbone_bd_ram_mem1_reg[74][14]/P0001 , \wishbone_bd_ram_mem1_reg[74][15]/P0001 , \wishbone_bd_ram_mem1_reg[74][8]/P0001 , \wishbone_bd_ram_mem1_reg[74][9]/P0001 , \wishbone_bd_ram_mem1_reg[75][10]/P0001 , \wishbone_bd_ram_mem1_reg[75][11]/P0001 , \wishbone_bd_ram_mem1_reg[75][12]/P0001 , \wishbone_bd_ram_mem1_reg[75][13]/P0001 , \wishbone_bd_ram_mem1_reg[75][14]/P0001 , \wishbone_bd_ram_mem1_reg[75][15]/P0001 , \wishbone_bd_ram_mem1_reg[75][8]/P0001 , \wishbone_bd_ram_mem1_reg[75][9]/P0001 , \wishbone_bd_ram_mem1_reg[76][10]/P0001 , \wishbone_bd_ram_mem1_reg[76][11]/P0001 , \wishbone_bd_ram_mem1_reg[76][12]/P0001 , \wishbone_bd_ram_mem1_reg[76][13]/P0001 , \wishbone_bd_ram_mem1_reg[76][14]/P0001 , \wishbone_bd_ram_mem1_reg[76][15]/P0001 , \wishbone_bd_ram_mem1_reg[76][8]/P0001 , \wishbone_bd_ram_mem1_reg[76][9]/P0001 , \wishbone_bd_ram_mem1_reg[77][10]/P0001 , \wishbone_bd_ram_mem1_reg[77][11]/P0001 , \wishbone_bd_ram_mem1_reg[77][12]/P0001 , \wishbone_bd_ram_mem1_reg[77][13]/P0001 , \wishbone_bd_ram_mem1_reg[77][14]/P0001 , \wishbone_bd_ram_mem1_reg[77][15]/P0001 , \wishbone_bd_ram_mem1_reg[77][8]/P0001 , \wishbone_bd_ram_mem1_reg[77][9]/P0001 , \wishbone_bd_ram_mem1_reg[78][10]/P0001 , \wishbone_bd_ram_mem1_reg[78][11]/P0001 , \wishbone_bd_ram_mem1_reg[78][12]/P0001 , \wishbone_bd_ram_mem1_reg[78][13]/P0001 , \wishbone_bd_ram_mem1_reg[78][14]/P0001 , \wishbone_bd_ram_mem1_reg[78][15]/P0001 , \wishbone_bd_ram_mem1_reg[78][8]/P0001 , \wishbone_bd_ram_mem1_reg[78][9]/P0001 , \wishbone_bd_ram_mem1_reg[79][10]/P0001 , \wishbone_bd_ram_mem1_reg[79][11]/P0001 , \wishbone_bd_ram_mem1_reg[79][12]/P0001 , \wishbone_bd_ram_mem1_reg[79][13]/P0001 , \wishbone_bd_ram_mem1_reg[79][14]/P0001 , \wishbone_bd_ram_mem1_reg[79][15]/P0001 , \wishbone_bd_ram_mem1_reg[79][8]/P0001 , \wishbone_bd_ram_mem1_reg[79][9]/P0001 , \wishbone_bd_ram_mem1_reg[7][10]/P0001 , \wishbone_bd_ram_mem1_reg[7][11]/P0001 , \wishbone_bd_ram_mem1_reg[7][12]/P0001 , \wishbone_bd_ram_mem1_reg[7][13]/P0001 , \wishbone_bd_ram_mem1_reg[7][14]/P0001 , \wishbone_bd_ram_mem1_reg[7][15]/P0001 , \wishbone_bd_ram_mem1_reg[7][8]/P0001 , \wishbone_bd_ram_mem1_reg[7][9]/P0001 , \wishbone_bd_ram_mem1_reg[80][10]/P0001 , \wishbone_bd_ram_mem1_reg[80][11]/P0001 , \wishbone_bd_ram_mem1_reg[80][12]/P0001 , \wishbone_bd_ram_mem1_reg[80][13]/P0001 , \wishbone_bd_ram_mem1_reg[80][14]/P0001 , \wishbone_bd_ram_mem1_reg[80][15]/P0001 , \wishbone_bd_ram_mem1_reg[80][8]/P0001 , \wishbone_bd_ram_mem1_reg[80][9]/P0001 , \wishbone_bd_ram_mem1_reg[81][10]/P0001 , \wishbone_bd_ram_mem1_reg[81][11]/P0001 , \wishbone_bd_ram_mem1_reg[81][12]/P0001 , \wishbone_bd_ram_mem1_reg[81][13]/P0001 , \wishbone_bd_ram_mem1_reg[81][14]/P0001 , \wishbone_bd_ram_mem1_reg[81][15]/P0001 , \wishbone_bd_ram_mem1_reg[81][8]/P0001 , \wishbone_bd_ram_mem1_reg[81][9]/P0001 , \wishbone_bd_ram_mem1_reg[82][10]/P0001 , \wishbone_bd_ram_mem1_reg[82][11]/P0001 , \wishbone_bd_ram_mem1_reg[82][12]/P0001 , \wishbone_bd_ram_mem1_reg[82][13]/P0001 , \wishbone_bd_ram_mem1_reg[82][14]/P0001 , \wishbone_bd_ram_mem1_reg[82][15]/P0001 , \wishbone_bd_ram_mem1_reg[82][8]/P0001 , \wishbone_bd_ram_mem1_reg[82][9]/P0001 , \wishbone_bd_ram_mem1_reg[83][10]/P0001 , \wishbone_bd_ram_mem1_reg[83][11]/P0001 , \wishbone_bd_ram_mem1_reg[83][12]/P0001 , \wishbone_bd_ram_mem1_reg[83][13]/P0001 , \wishbone_bd_ram_mem1_reg[83][14]/P0001 , \wishbone_bd_ram_mem1_reg[83][15]/P0001 , \wishbone_bd_ram_mem1_reg[83][8]/P0001 , \wishbone_bd_ram_mem1_reg[83][9]/P0001 , \wishbone_bd_ram_mem1_reg[84][10]/P0001 , \wishbone_bd_ram_mem1_reg[84][11]/P0001 , \wishbone_bd_ram_mem1_reg[84][12]/P0001 , \wishbone_bd_ram_mem1_reg[84][13]/P0001 , \wishbone_bd_ram_mem1_reg[84][14]/P0001 , \wishbone_bd_ram_mem1_reg[84][15]/P0001 , \wishbone_bd_ram_mem1_reg[84][8]/P0001 , \wishbone_bd_ram_mem1_reg[84][9]/P0001 , \wishbone_bd_ram_mem1_reg[85][10]/P0001 , \wishbone_bd_ram_mem1_reg[85][11]/P0001 , \wishbone_bd_ram_mem1_reg[85][12]/P0001 , \wishbone_bd_ram_mem1_reg[85][13]/P0001 , \wishbone_bd_ram_mem1_reg[85][14]/P0001 , \wishbone_bd_ram_mem1_reg[85][15]/P0001 , \wishbone_bd_ram_mem1_reg[85][8]/P0001 , \wishbone_bd_ram_mem1_reg[85][9]/P0001 , \wishbone_bd_ram_mem1_reg[86][10]/P0001 , \wishbone_bd_ram_mem1_reg[86][11]/P0001 , \wishbone_bd_ram_mem1_reg[86][12]/P0001 , \wishbone_bd_ram_mem1_reg[86][13]/P0001 , \wishbone_bd_ram_mem1_reg[86][14]/P0001 , \wishbone_bd_ram_mem1_reg[86][15]/P0001 , \wishbone_bd_ram_mem1_reg[86][8]/P0001 , \wishbone_bd_ram_mem1_reg[86][9]/P0001 , \wishbone_bd_ram_mem1_reg[87][10]/P0001 , \wishbone_bd_ram_mem1_reg[87][11]/P0001 , \wishbone_bd_ram_mem1_reg[87][12]/P0001 , \wishbone_bd_ram_mem1_reg[87][13]/P0001 , \wishbone_bd_ram_mem1_reg[87][14]/P0001 , \wishbone_bd_ram_mem1_reg[87][15]/P0001 , \wishbone_bd_ram_mem1_reg[87][8]/P0001 , \wishbone_bd_ram_mem1_reg[87][9]/P0001 , \wishbone_bd_ram_mem1_reg[88][10]/P0001 , \wishbone_bd_ram_mem1_reg[88][11]/P0001 , \wishbone_bd_ram_mem1_reg[88][12]/P0001 , \wishbone_bd_ram_mem1_reg[88][13]/P0001 , \wishbone_bd_ram_mem1_reg[88][14]/P0001 , \wishbone_bd_ram_mem1_reg[88][15]/P0001 , \wishbone_bd_ram_mem1_reg[88][8]/P0001 , \wishbone_bd_ram_mem1_reg[88][9]/P0001 , \wishbone_bd_ram_mem1_reg[89][10]/P0001 , \wishbone_bd_ram_mem1_reg[89][11]/P0001 , \wishbone_bd_ram_mem1_reg[89][12]/P0001 , \wishbone_bd_ram_mem1_reg[89][13]/P0001 , \wishbone_bd_ram_mem1_reg[89][14]/P0001 , \wishbone_bd_ram_mem1_reg[89][15]/P0001 , \wishbone_bd_ram_mem1_reg[89][8]/P0001 , \wishbone_bd_ram_mem1_reg[89][9]/P0001 , \wishbone_bd_ram_mem1_reg[8][10]/P0001 , \wishbone_bd_ram_mem1_reg[8][11]/P0001 , \wishbone_bd_ram_mem1_reg[8][12]/P0001 , \wishbone_bd_ram_mem1_reg[8][13]/P0001 , \wishbone_bd_ram_mem1_reg[8][14]/P0001 , \wishbone_bd_ram_mem1_reg[8][15]/P0001 , \wishbone_bd_ram_mem1_reg[8][8]/P0001 , \wishbone_bd_ram_mem1_reg[8][9]/P0001 , \wishbone_bd_ram_mem1_reg[90][10]/P0001 , \wishbone_bd_ram_mem1_reg[90][11]/P0001 , \wishbone_bd_ram_mem1_reg[90][12]/P0001 , \wishbone_bd_ram_mem1_reg[90][13]/P0001 , \wishbone_bd_ram_mem1_reg[90][14]/P0001 , \wishbone_bd_ram_mem1_reg[90][15]/P0001 , \wishbone_bd_ram_mem1_reg[90][8]/P0001 , \wishbone_bd_ram_mem1_reg[90][9]/P0001 , \wishbone_bd_ram_mem1_reg[91][10]/P0001 , \wishbone_bd_ram_mem1_reg[91][11]/P0001 , \wishbone_bd_ram_mem1_reg[91][12]/P0001 , \wishbone_bd_ram_mem1_reg[91][13]/P0001 , \wishbone_bd_ram_mem1_reg[91][14]/P0001 , \wishbone_bd_ram_mem1_reg[91][15]/P0001 , \wishbone_bd_ram_mem1_reg[91][8]/P0001 , \wishbone_bd_ram_mem1_reg[91][9]/P0001 , \wishbone_bd_ram_mem1_reg[92][10]/P0001 , \wishbone_bd_ram_mem1_reg[92][11]/P0001 , \wishbone_bd_ram_mem1_reg[92][12]/P0001 , \wishbone_bd_ram_mem1_reg[92][13]/P0001 , \wishbone_bd_ram_mem1_reg[92][14]/P0001 , \wishbone_bd_ram_mem1_reg[92][15]/P0001 , \wishbone_bd_ram_mem1_reg[92][8]/P0001 , \wishbone_bd_ram_mem1_reg[92][9]/P0001 , \wishbone_bd_ram_mem1_reg[93][10]/P0001 , \wishbone_bd_ram_mem1_reg[93][11]/P0001 , \wishbone_bd_ram_mem1_reg[93][12]/P0001 , \wishbone_bd_ram_mem1_reg[93][13]/P0001 , \wishbone_bd_ram_mem1_reg[93][14]/P0001 , \wishbone_bd_ram_mem1_reg[93][15]/P0001 , \wishbone_bd_ram_mem1_reg[93][8]/P0001 , \wishbone_bd_ram_mem1_reg[93][9]/P0001 , \wishbone_bd_ram_mem1_reg[94][10]/P0001 , \wishbone_bd_ram_mem1_reg[94][11]/P0001 , \wishbone_bd_ram_mem1_reg[94][12]/P0001 , \wishbone_bd_ram_mem1_reg[94][13]/P0001 , \wishbone_bd_ram_mem1_reg[94][14]/P0001 , \wishbone_bd_ram_mem1_reg[94][15]/P0001 , \wishbone_bd_ram_mem1_reg[94][8]/P0001 , \wishbone_bd_ram_mem1_reg[94][9]/P0001 , \wishbone_bd_ram_mem1_reg[95][10]/P0001 , \wishbone_bd_ram_mem1_reg[95][11]/P0001 , \wishbone_bd_ram_mem1_reg[95][12]/P0001 , \wishbone_bd_ram_mem1_reg[95][13]/P0001 , \wishbone_bd_ram_mem1_reg[95][14]/P0001 , \wishbone_bd_ram_mem1_reg[95][15]/P0001 , \wishbone_bd_ram_mem1_reg[95][8]/P0001 , \wishbone_bd_ram_mem1_reg[95][9]/P0001 , \wishbone_bd_ram_mem1_reg[96][10]/P0001 , \wishbone_bd_ram_mem1_reg[96][11]/P0001 , \wishbone_bd_ram_mem1_reg[96][12]/P0001 , \wishbone_bd_ram_mem1_reg[96][13]/P0001 , \wishbone_bd_ram_mem1_reg[96][14]/P0001 , \wishbone_bd_ram_mem1_reg[96][15]/P0001 , \wishbone_bd_ram_mem1_reg[96][8]/P0001 , \wishbone_bd_ram_mem1_reg[96][9]/P0001 , \wishbone_bd_ram_mem1_reg[97][10]/P0001 , \wishbone_bd_ram_mem1_reg[97][11]/P0001 , \wishbone_bd_ram_mem1_reg[97][12]/P0001 , \wishbone_bd_ram_mem1_reg[97][13]/P0001 , \wishbone_bd_ram_mem1_reg[97][14]/P0001 , \wishbone_bd_ram_mem1_reg[97][15]/P0001 , \wishbone_bd_ram_mem1_reg[97][8]/P0001 , \wishbone_bd_ram_mem1_reg[97][9]/P0001 , \wishbone_bd_ram_mem1_reg[98][10]/P0001 , \wishbone_bd_ram_mem1_reg[98][11]/P0001 , \wishbone_bd_ram_mem1_reg[98][12]/P0001 , \wishbone_bd_ram_mem1_reg[98][13]/P0001 , \wishbone_bd_ram_mem1_reg[98][14]/P0001 , \wishbone_bd_ram_mem1_reg[98][15]/P0001 , \wishbone_bd_ram_mem1_reg[98][8]/P0001 , \wishbone_bd_ram_mem1_reg[98][9]/P0001 , \wishbone_bd_ram_mem1_reg[99][10]/P0001 , \wishbone_bd_ram_mem1_reg[99][11]/P0001 , \wishbone_bd_ram_mem1_reg[99][12]/P0001 , \wishbone_bd_ram_mem1_reg[99][13]/P0001 , \wishbone_bd_ram_mem1_reg[99][14]/P0001 , \wishbone_bd_ram_mem1_reg[99][15]/P0001 , \wishbone_bd_ram_mem1_reg[99][8]/P0001 , \wishbone_bd_ram_mem1_reg[99][9]/P0001 , \wishbone_bd_ram_mem1_reg[9][10]/P0001 , \wishbone_bd_ram_mem1_reg[9][11]/P0001 , \wishbone_bd_ram_mem1_reg[9][12]/P0001 , \wishbone_bd_ram_mem1_reg[9][13]/P0001 , \wishbone_bd_ram_mem1_reg[9][14]/P0001 , \wishbone_bd_ram_mem1_reg[9][15]/P0001 , \wishbone_bd_ram_mem1_reg[9][8]/P0001 , \wishbone_bd_ram_mem1_reg[9][9]/P0001 , \wishbone_bd_ram_mem2_reg[0][16]/P0001 , \wishbone_bd_ram_mem2_reg[0][17]/P0001 , \wishbone_bd_ram_mem2_reg[0][18]/P0001 , \wishbone_bd_ram_mem2_reg[0][19]/P0001 , \wishbone_bd_ram_mem2_reg[0][20]/P0001 , \wishbone_bd_ram_mem2_reg[0][21]/P0001 , \wishbone_bd_ram_mem2_reg[0][22]/P0001 , \wishbone_bd_ram_mem2_reg[0][23]/P0001 , \wishbone_bd_ram_mem2_reg[100][16]/P0001 , \wishbone_bd_ram_mem2_reg[100][17]/P0001 , \wishbone_bd_ram_mem2_reg[100][18]/P0001 , \wishbone_bd_ram_mem2_reg[100][19]/P0001 , \wishbone_bd_ram_mem2_reg[100][20]/P0001 , \wishbone_bd_ram_mem2_reg[100][21]/P0001 , \wishbone_bd_ram_mem2_reg[100][22]/P0001 , \wishbone_bd_ram_mem2_reg[100][23]/P0001 , \wishbone_bd_ram_mem2_reg[101][16]/P0001 , \wishbone_bd_ram_mem2_reg[101][17]/P0001 , \wishbone_bd_ram_mem2_reg[101][18]/P0001 , \wishbone_bd_ram_mem2_reg[101][19]/P0001 , \wishbone_bd_ram_mem2_reg[101][20]/P0001 , \wishbone_bd_ram_mem2_reg[101][21]/P0001 , \wishbone_bd_ram_mem2_reg[101][22]/P0001 , \wishbone_bd_ram_mem2_reg[101][23]/P0001 , \wishbone_bd_ram_mem2_reg[102][16]/P0001 , \wishbone_bd_ram_mem2_reg[102][17]/P0001 , \wishbone_bd_ram_mem2_reg[102][18]/P0001 , \wishbone_bd_ram_mem2_reg[102][19]/P0001 , \wishbone_bd_ram_mem2_reg[102][20]/P0001 , \wishbone_bd_ram_mem2_reg[102][21]/P0001 , \wishbone_bd_ram_mem2_reg[102][22]/P0001 , \wishbone_bd_ram_mem2_reg[102][23]/P0001 , \wishbone_bd_ram_mem2_reg[103][16]/P0001 , \wishbone_bd_ram_mem2_reg[103][17]/P0001 , \wishbone_bd_ram_mem2_reg[103][18]/P0001 , \wishbone_bd_ram_mem2_reg[103][19]/P0001 , \wishbone_bd_ram_mem2_reg[103][20]/P0001 , \wishbone_bd_ram_mem2_reg[103][21]/P0001 , \wishbone_bd_ram_mem2_reg[103][22]/P0001 , \wishbone_bd_ram_mem2_reg[103][23]/P0001 , \wishbone_bd_ram_mem2_reg[104][16]/P0001 , \wishbone_bd_ram_mem2_reg[104][17]/P0001 , \wishbone_bd_ram_mem2_reg[104][18]/P0001 , \wishbone_bd_ram_mem2_reg[104][19]/P0001 , \wishbone_bd_ram_mem2_reg[104][20]/P0001 , \wishbone_bd_ram_mem2_reg[104][21]/P0001 , \wishbone_bd_ram_mem2_reg[104][22]/P0001 , \wishbone_bd_ram_mem2_reg[104][23]/P0001 , \wishbone_bd_ram_mem2_reg[105][16]/P0001 , \wishbone_bd_ram_mem2_reg[105][17]/P0001 , \wishbone_bd_ram_mem2_reg[105][18]/P0001 , \wishbone_bd_ram_mem2_reg[105][19]/P0001 , \wishbone_bd_ram_mem2_reg[105][20]/P0001 , \wishbone_bd_ram_mem2_reg[105][21]/P0001 , \wishbone_bd_ram_mem2_reg[105][22]/P0001 , \wishbone_bd_ram_mem2_reg[105][23]/P0001 , \wishbone_bd_ram_mem2_reg[106][16]/P0001 , \wishbone_bd_ram_mem2_reg[106][17]/P0001 , \wishbone_bd_ram_mem2_reg[106][18]/P0001 , \wishbone_bd_ram_mem2_reg[106][19]/P0001 , \wishbone_bd_ram_mem2_reg[106][20]/P0001 , \wishbone_bd_ram_mem2_reg[106][21]/P0001 , \wishbone_bd_ram_mem2_reg[106][22]/P0001 , \wishbone_bd_ram_mem2_reg[106][23]/P0001 , \wishbone_bd_ram_mem2_reg[107][16]/P0001 , \wishbone_bd_ram_mem2_reg[107][17]/P0001 , \wishbone_bd_ram_mem2_reg[107][18]/P0001 , \wishbone_bd_ram_mem2_reg[107][19]/P0001 , \wishbone_bd_ram_mem2_reg[107][20]/P0001 , \wishbone_bd_ram_mem2_reg[107][21]/P0001 , \wishbone_bd_ram_mem2_reg[107][22]/P0001 , \wishbone_bd_ram_mem2_reg[107][23]/P0001 , \wishbone_bd_ram_mem2_reg[108][16]/P0001 , \wishbone_bd_ram_mem2_reg[108][17]/P0001 , \wishbone_bd_ram_mem2_reg[108][18]/P0001 , \wishbone_bd_ram_mem2_reg[108][19]/P0001 , \wishbone_bd_ram_mem2_reg[108][20]/P0001 , \wishbone_bd_ram_mem2_reg[108][21]/P0001 , \wishbone_bd_ram_mem2_reg[108][22]/P0001 , \wishbone_bd_ram_mem2_reg[108][23]/P0001 , \wishbone_bd_ram_mem2_reg[109][16]/P0001 , \wishbone_bd_ram_mem2_reg[109][17]/P0001 , \wishbone_bd_ram_mem2_reg[109][18]/P0001 , \wishbone_bd_ram_mem2_reg[109][19]/P0001 , \wishbone_bd_ram_mem2_reg[109][20]/P0001 , \wishbone_bd_ram_mem2_reg[109][21]/P0001 , \wishbone_bd_ram_mem2_reg[109][22]/P0001 , \wishbone_bd_ram_mem2_reg[109][23]/P0001 , \wishbone_bd_ram_mem2_reg[10][16]/P0001 , \wishbone_bd_ram_mem2_reg[10][17]/P0001 , \wishbone_bd_ram_mem2_reg[10][18]/P0001 , \wishbone_bd_ram_mem2_reg[10][19]/P0001 , \wishbone_bd_ram_mem2_reg[10][20]/P0001 , \wishbone_bd_ram_mem2_reg[10][21]/P0001 , \wishbone_bd_ram_mem2_reg[10][22]/P0001 , \wishbone_bd_ram_mem2_reg[10][23]/P0001 , \wishbone_bd_ram_mem2_reg[110][16]/P0001 , \wishbone_bd_ram_mem2_reg[110][17]/P0001 , \wishbone_bd_ram_mem2_reg[110][18]/P0001 , \wishbone_bd_ram_mem2_reg[110][19]/P0001 , \wishbone_bd_ram_mem2_reg[110][20]/P0001 , \wishbone_bd_ram_mem2_reg[110][21]/P0001 , \wishbone_bd_ram_mem2_reg[110][22]/P0001 , \wishbone_bd_ram_mem2_reg[110][23]/P0001 , \wishbone_bd_ram_mem2_reg[111][16]/P0001 , \wishbone_bd_ram_mem2_reg[111][17]/P0001 , \wishbone_bd_ram_mem2_reg[111][18]/P0001 , \wishbone_bd_ram_mem2_reg[111][19]/P0001 , \wishbone_bd_ram_mem2_reg[111][20]/P0001 , \wishbone_bd_ram_mem2_reg[111][21]/P0001 , \wishbone_bd_ram_mem2_reg[111][22]/P0001 , \wishbone_bd_ram_mem2_reg[111][23]/P0001 , \wishbone_bd_ram_mem2_reg[112][16]/P0001 , \wishbone_bd_ram_mem2_reg[112][17]/P0001 , \wishbone_bd_ram_mem2_reg[112][18]/P0001 , \wishbone_bd_ram_mem2_reg[112][19]/P0001 , \wishbone_bd_ram_mem2_reg[112][20]/P0001 , \wishbone_bd_ram_mem2_reg[112][21]/P0001 , \wishbone_bd_ram_mem2_reg[112][22]/P0001 , \wishbone_bd_ram_mem2_reg[112][23]/P0001 , \wishbone_bd_ram_mem2_reg[113][16]/P0001 , \wishbone_bd_ram_mem2_reg[113][17]/P0001 , \wishbone_bd_ram_mem2_reg[113][18]/P0001 , \wishbone_bd_ram_mem2_reg[113][19]/P0001 , \wishbone_bd_ram_mem2_reg[113][20]/P0001 , \wishbone_bd_ram_mem2_reg[113][21]/P0001 , \wishbone_bd_ram_mem2_reg[113][22]/P0001 , \wishbone_bd_ram_mem2_reg[113][23]/P0001 , \wishbone_bd_ram_mem2_reg[114][16]/P0001 , \wishbone_bd_ram_mem2_reg[114][17]/P0001 , \wishbone_bd_ram_mem2_reg[114][18]/P0001 , \wishbone_bd_ram_mem2_reg[114][19]/P0001 , \wishbone_bd_ram_mem2_reg[114][20]/P0001 , \wishbone_bd_ram_mem2_reg[114][21]/P0001 , \wishbone_bd_ram_mem2_reg[114][22]/P0001 , \wishbone_bd_ram_mem2_reg[114][23]/P0001 , \wishbone_bd_ram_mem2_reg[115][16]/P0001 , \wishbone_bd_ram_mem2_reg[115][17]/P0001 , \wishbone_bd_ram_mem2_reg[115][18]/P0001 , \wishbone_bd_ram_mem2_reg[115][19]/P0001 , \wishbone_bd_ram_mem2_reg[115][20]/P0001 , \wishbone_bd_ram_mem2_reg[115][21]/P0001 , \wishbone_bd_ram_mem2_reg[115][22]/P0001 , \wishbone_bd_ram_mem2_reg[115][23]/P0001 , \wishbone_bd_ram_mem2_reg[116][16]/P0001 , \wishbone_bd_ram_mem2_reg[116][17]/P0001 , \wishbone_bd_ram_mem2_reg[116][18]/P0001 , \wishbone_bd_ram_mem2_reg[116][19]/P0001 , \wishbone_bd_ram_mem2_reg[116][20]/P0001 , \wishbone_bd_ram_mem2_reg[116][21]/P0001 , \wishbone_bd_ram_mem2_reg[116][22]/P0001 , \wishbone_bd_ram_mem2_reg[116][23]/P0001 , \wishbone_bd_ram_mem2_reg[117][16]/P0001 , \wishbone_bd_ram_mem2_reg[117][17]/P0001 , \wishbone_bd_ram_mem2_reg[117][18]/P0001 , \wishbone_bd_ram_mem2_reg[117][19]/P0001 , \wishbone_bd_ram_mem2_reg[117][20]/P0001 , \wishbone_bd_ram_mem2_reg[117][21]/P0001 , \wishbone_bd_ram_mem2_reg[117][22]/P0001 , \wishbone_bd_ram_mem2_reg[117][23]/P0001 , \wishbone_bd_ram_mem2_reg[118][16]/P0001 , \wishbone_bd_ram_mem2_reg[118][17]/P0001 , \wishbone_bd_ram_mem2_reg[118][18]/P0001 , \wishbone_bd_ram_mem2_reg[118][19]/P0001 , \wishbone_bd_ram_mem2_reg[118][20]/P0001 , \wishbone_bd_ram_mem2_reg[118][21]/P0001 , \wishbone_bd_ram_mem2_reg[118][22]/P0001 , \wishbone_bd_ram_mem2_reg[118][23]/P0001 , \wishbone_bd_ram_mem2_reg[119][16]/P0001 , \wishbone_bd_ram_mem2_reg[119][17]/P0001 , \wishbone_bd_ram_mem2_reg[119][18]/P0001 , \wishbone_bd_ram_mem2_reg[119][19]/P0001 , \wishbone_bd_ram_mem2_reg[119][20]/P0001 , \wishbone_bd_ram_mem2_reg[119][21]/P0001 , \wishbone_bd_ram_mem2_reg[119][22]/P0001 , \wishbone_bd_ram_mem2_reg[119][23]/P0001 , \wishbone_bd_ram_mem2_reg[11][16]/P0001 , \wishbone_bd_ram_mem2_reg[11][17]/P0001 , \wishbone_bd_ram_mem2_reg[11][18]/P0001 , \wishbone_bd_ram_mem2_reg[11][19]/P0001 , \wishbone_bd_ram_mem2_reg[11][20]/P0001 , \wishbone_bd_ram_mem2_reg[11][21]/P0001 , \wishbone_bd_ram_mem2_reg[11][22]/P0001 , \wishbone_bd_ram_mem2_reg[11][23]/P0001 , \wishbone_bd_ram_mem2_reg[120][16]/P0001 , \wishbone_bd_ram_mem2_reg[120][17]/P0001 , \wishbone_bd_ram_mem2_reg[120][18]/P0001 , \wishbone_bd_ram_mem2_reg[120][19]/P0001 , \wishbone_bd_ram_mem2_reg[120][20]/P0001 , \wishbone_bd_ram_mem2_reg[120][21]/P0001 , \wishbone_bd_ram_mem2_reg[120][22]/P0001 , \wishbone_bd_ram_mem2_reg[120][23]/P0001 , \wishbone_bd_ram_mem2_reg[121][16]/P0001 , \wishbone_bd_ram_mem2_reg[121][17]/P0001 , \wishbone_bd_ram_mem2_reg[121][18]/P0001 , \wishbone_bd_ram_mem2_reg[121][19]/P0001 , \wishbone_bd_ram_mem2_reg[121][20]/P0001 , \wishbone_bd_ram_mem2_reg[121][21]/P0001 , \wishbone_bd_ram_mem2_reg[121][22]/P0001 , \wishbone_bd_ram_mem2_reg[121][23]/P0001 , \wishbone_bd_ram_mem2_reg[122][16]/P0001 , \wishbone_bd_ram_mem2_reg[122][17]/P0001 , \wishbone_bd_ram_mem2_reg[122][18]/P0001 , \wishbone_bd_ram_mem2_reg[122][19]/P0001 , \wishbone_bd_ram_mem2_reg[122][20]/P0001 , \wishbone_bd_ram_mem2_reg[122][21]/P0001 , \wishbone_bd_ram_mem2_reg[122][22]/P0001 , \wishbone_bd_ram_mem2_reg[122][23]/P0001 , \wishbone_bd_ram_mem2_reg[123][16]/P0001 , \wishbone_bd_ram_mem2_reg[123][17]/P0001 , \wishbone_bd_ram_mem2_reg[123][18]/P0001 , \wishbone_bd_ram_mem2_reg[123][19]/P0001 , \wishbone_bd_ram_mem2_reg[123][20]/P0001 , \wishbone_bd_ram_mem2_reg[123][21]/P0001 , \wishbone_bd_ram_mem2_reg[123][22]/P0001 , \wishbone_bd_ram_mem2_reg[123][23]/P0001 , \wishbone_bd_ram_mem2_reg[124][16]/P0001 , \wishbone_bd_ram_mem2_reg[124][17]/P0001 , \wishbone_bd_ram_mem2_reg[124][18]/P0001 , \wishbone_bd_ram_mem2_reg[124][19]/P0001 , \wishbone_bd_ram_mem2_reg[124][20]/P0001 , \wishbone_bd_ram_mem2_reg[124][21]/P0001 , \wishbone_bd_ram_mem2_reg[124][22]/P0001 , \wishbone_bd_ram_mem2_reg[124][23]/P0001 , \wishbone_bd_ram_mem2_reg[125][16]/P0001 , \wishbone_bd_ram_mem2_reg[125][17]/P0001 , \wishbone_bd_ram_mem2_reg[125][18]/P0001 , \wishbone_bd_ram_mem2_reg[125][19]/P0001 , \wishbone_bd_ram_mem2_reg[125][20]/P0001 , \wishbone_bd_ram_mem2_reg[125][21]/P0001 , \wishbone_bd_ram_mem2_reg[125][22]/P0001 , \wishbone_bd_ram_mem2_reg[125][23]/P0001 , \wishbone_bd_ram_mem2_reg[126][16]/P0001 , \wishbone_bd_ram_mem2_reg[126][17]/P0001 , \wishbone_bd_ram_mem2_reg[126][18]/P0001 , \wishbone_bd_ram_mem2_reg[126][19]/P0001 , \wishbone_bd_ram_mem2_reg[126][20]/P0001 , \wishbone_bd_ram_mem2_reg[126][21]/P0001 , \wishbone_bd_ram_mem2_reg[126][22]/P0001 , \wishbone_bd_ram_mem2_reg[126][23]/P0001 , \wishbone_bd_ram_mem2_reg[127][16]/P0001 , \wishbone_bd_ram_mem2_reg[127][17]/P0001 , \wishbone_bd_ram_mem2_reg[127][18]/P0001 , \wishbone_bd_ram_mem2_reg[127][19]/P0001 , \wishbone_bd_ram_mem2_reg[127][20]/P0001 , \wishbone_bd_ram_mem2_reg[127][21]/P0001 , \wishbone_bd_ram_mem2_reg[127][22]/P0001 , \wishbone_bd_ram_mem2_reg[127][23]/P0001 , \wishbone_bd_ram_mem2_reg[128][16]/P0001 , \wishbone_bd_ram_mem2_reg[128][17]/P0001 , \wishbone_bd_ram_mem2_reg[128][18]/P0001 , \wishbone_bd_ram_mem2_reg[128][19]/P0001 , \wishbone_bd_ram_mem2_reg[128][20]/P0001 , \wishbone_bd_ram_mem2_reg[128][21]/P0001 , \wishbone_bd_ram_mem2_reg[128][22]/P0001 , \wishbone_bd_ram_mem2_reg[128][23]/P0001 , \wishbone_bd_ram_mem2_reg[129][16]/P0001 , \wishbone_bd_ram_mem2_reg[129][17]/P0001 , \wishbone_bd_ram_mem2_reg[129][18]/P0001 , \wishbone_bd_ram_mem2_reg[129][19]/P0001 , \wishbone_bd_ram_mem2_reg[129][20]/P0001 , \wishbone_bd_ram_mem2_reg[129][21]/P0001 , \wishbone_bd_ram_mem2_reg[129][22]/P0001 , \wishbone_bd_ram_mem2_reg[129][23]/P0001 , \wishbone_bd_ram_mem2_reg[12][16]/P0001 , \wishbone_bd_ram_mem2_reg[12][17]/P0001 , \wishbone_bd_ram_mem2_reg[12][18]/P0001 , \wishbone_bd_ram_mem2_reg[12][19]/P0001 , \wishbone_bd_ram_mem2_reg[12][20]/P0001 , \wishbone_bd_ram_mem2_reg[12][21]/P0001 , \wishbone_bd_ram_mem2_reg[12][22]/P0001 , \wishbone_bd_ram_mem2_reg[12][23]/P0001 , \wishbone_bd_ram_mem2_reg[130][16]/P0001 , \wishbone_bd_ram_mem2_reg[130][17]/P0001 , \wishbone_bd_ram_mem2_reg[130][18]/P0001 , \wishbone_bd_ram_mem2_reg[130][19]/P0001 , \wishbone_bd_ram_mem2_reg[130][20]/P0001 , \wishbone_bd_ram_mem2_reg[130][21]/P0001 , \wishbone_bd_ram_mem2_reg[130][22]/P0001 , \wishbone_bd_ram_mem2_reg[130][23]/P0001 , \wishbone_bd_ram_mem2_reg[131][16]/P0001 , \wishbone_bd_ram_mem2_reg[131][17]/P0001 , \wishbone_bd_ram_mem2_reg[131][18]/P0001 , \wishbone_bd_ram_mem2_reg[131][19]/P0001 , \wishbone_bd_ram_mem2_reg[131][20]/P0001 , \wishbone_bd_ram_mem2_reg[131][21]/P0001 , \wishbone_bd_ram_mem2_reg[131][22]/P0001 , \wishbone_bd_ram_mem2_reg[131][23]/P0001 , \wishbone_bd_ram_mem2_reg[132][16]/P0001 , \wishbone_bd_ram_mem2_reg[132][17]/P0001 , \wishbone_bd_ram_mem2_reg[132][18]/P0001 , \wishbone_bd_ram_mem2_reg[132][19]/P0001 , \wishbone_bd_ram_mem2_reg[132][20]/P0001 , \wishbone_bd_ram_mem2_reg[132][21]/P0001 , \wishbone_bd_ram_mem2_reg[132][22]/P0001 , \wishbone_bd_ram_mem2_reg[132][23]/P0001 , \wishbone_bd_ram_mem2_reg[133][16]/P0001 , \wishbone_bd_ram_mem2_reg[133][17]/P0001 , \wishbone_bd_ram_mem2_reg[133][18]/P0001 , \wishbone_bd_ram_mem2_reg[133][19]/P0001 , \wishbone_bd_ram_mem2_reg[133][20]/P0001 , \wishbone_bd_ram_mem2_reg[133][21]/P0001 , \wishbone_bd_ram_mem2_reg[133][22]/P0001 , \wishbone_bd_ram_mem2_reg[133][23]/P0001 , \wishbone_bd_ram_mem2_reg[134][16]/P0001 , \wishbone_bd_ram_mem2_reg[134][17]/P0001 , \wishbone_bd_ram_mem2_reg[134][18]/P0001 , \wishbone_bd_ram_mem2_reg[134][19]/P0001 , \wishbone_bd_ram_mem2_reg[134][20]/P0001 , \wishbone_bd_ram_mem2_reg[134][21]/P0001 , \wishbone_bd_ram_mem2_reg[134][22]/P0001 , \wishbone_bd_ram_mem2_reg[134][23]/P0001 , \wishbone_bd_ram_mem2_reg[135][16]/P0001 , \wishbone_bd_ram_mem2_reg[135][17]/P0001 , \wishbone_bd_ram_mem2_reg[135][18]/P0001 , \wishbone_bd_ram_mem2_reg[135][19]/P0001 , \wishbone_bd_ram_mem2_reg[135][20]/P0001 , \wishbone_bd_ram_mem2_reg[135][21]/P0001 , \wishbone_bd_ram_mem2_reg[135][22]/P0001 , \wishbone_bd_ram_mem2_reg[135][23]/P0001 , \wishbone_bd_ram_mem2_reg[136][16]/P0001 , \wishbone_bd_ram_mem2_reg[136][17]/P0001 , \wishbone_bd_ram_mem2_reg[136][18]/P0001 , \wishbone_bd_ram_mem2_reg[136][19]/P0001 , \wishbone_bd_ram_mem2_reg[136][20]/P0001 , \wishbone_bd_ram_mem2_reg[136][21]/P0001 , \wishbone_bd_ram_mem2_reg[136][22]/P0001 , \wishbone_bd_ram_mem2_reg[136][23]/P0001 , \wishbone_bd_ram_mem2_reg[137][16]/P0001 , \wishbone_bd_ram_mem2_reg[137][17]/P0001 , \wishbone_bd_ram_mem2_reg[137][18]/P0001 , \wishbone_bd_ram_mem2_reg[137][19]/P0001 , \wishbone_bd_ram_mem2_reg[137][20]/P0001 , \wishbone_bd_ram_mem2_reg[137][21]/P0001 , \wishbone_bd_ram_mem2_reg[137][22]/P0001 , \wishbone_bd_ram_mem2_reg[137][23]/P0001 , \wishbone_bd_ram_mem2_reg[138][16]/P0001 , \wishbone_bd_ram_mem2_reg[138][17]/P0001 , \wishbone_bd_ram_mem2_reg[138][18]/P0001 , \wishbone_bd_ram_mem2_reg[138][19]/P0001 , \wishbone_bd_ram_mem2_reg[138][20]/P0001 , \wishbone_bd_ram_mem2_reg[138][21]/P0001 , \wishbone_bd_ram_mem2_reg[138][22]/P0001 , \wishbone_bd_ram_mem2_reg[138][23]/P0001 , \wishbone_bd_ram_mem2_reg[139][16]/P0001 , \wishbone_bd_ram_mem2_reg[139][17]/P0001 , \wishbone_bd_ram_mem2_reg[139][18]/P0001 , \wishbone_bd_ram_mem2_reg[139][19]/P0001 , \wishbone_bd_ram_mem2_reg[139][20]/P0001 , \wishbone_bd_ram_mem2_reg[139][21]/P0001 , \wishbone_bd_ram_mem2_reg[139][22]/P0001 , \wishbone_bd_ram_mem2_reg[139][23]/P0001 , \wishbone_bd_ram_mem2_reg[13][16]/P0001 , \wishbone_bd_ram_mem2_reg[13][17]/P0001 , \wishbone_bd_ram_mem2_reg[13][18]/P0001 , \wishbone_bd_ram_mem2_reg[13][19]/P0001 , \wishbone_bd_ram_mem2_reg[13][20]/P0001 , \wishbone_bd_ram_mem2_reg[13][21]/P0001 , \wishbone_bd_ram_mem2_reg[13][22]/P0001 , \wishbone_bd_ram_mem2_reg[13][23]/P0001 , \wishbone_bd_ram_mem2_reg[140][16]/P0001 , \wishbone_bd_ram_mem2_reg[140][17]/P0001 , \wishbone_bd_ram_mem2_reg[140][18]/P0001 , \wishbone_bd_ram_mem2_reg[140][19]/P0001 , \wishbone_bd_ram_mem2_reg[140][20]/P0001 , \wishbone_bd_ram_mem2_reg[140][21]/P0001 , \wishbone_bd_ram_mem2_reg[140][22]/P0001 , \wishbone_bd_ram_mem2_reg[140][23]/P0001 , \wishbone_bd_ram_mem2_reg[141][16]/P0001 , \wishbone_bd_ram_mem2_reg[141][17]/P0001 , \wishbone_bd_ram_mem2_reg[141][18]/P0001 , \wishbone_bd_ram_mem2_reg[141][19]/P0001 , \wishbone_bd_ram_mem2_reg[141][20]/P0001 , \wishbone_bd_ram_mem2_reg[141][21]/P0001 , \wishbone_bd_ram_mem2_reg[141][22]/P0001 , \wishbone_bd_ram_mem2_reg[141][23]/P0001 , \wishbone_bd_ram_mem2_reg[142][16]/P0001 , \wishbone_bd_ram_mem2_reg[142][17]/P0001 , \wishbone_bd_ram_mem2_reg[142][18]/P0001 , \wishbone_bd_ram_mem2_reg[142][19]/P0001 , \wishbone_bd_ram_mem2_reg[142][20]/P0001 , \wishbone_bd_ram_mem2_reg[142][21]/P0001 , \wishbone_bd_ram_mem2_reg[142][22]/P0001 , \wishbone_bd_ram_mem2_reg[142][23]/P0001 , \wishbone_bd_ram_mem2_reg[143][16]/P0001 , \wishbone_bd_ram_mem2_reg[143][17]/P0001 , \wishbone_bd_ram_mem2_reg[143][18]/P0001 , \wishbone_bd_ram_mem2_reg[143][19]/P0001 , \wishbone_bd_ram_mem2_reg[143][20]/P0001 , \wishbone_bd_ram_mem2_reg[143][21]/P0001 , \wishbone_bd_ram_mem2_reg[143][22]/P0001 , \wishbone_bd_ram_mem2_reg[143][23]/P0001 , \wishbone_bd_ram_mem2_reg[144][16]/P0001 , \wishbone_bd_ram_mem2_reg[144][17]/P0001 , \wishbone_bd_ram_mem2_reg[144][18]/P0001 , \wishbone_bd_ram_mem2_reg[144][19]/P0001 , \wishbone_bd_ram_mem2_reg[144][20]/P0001 , \wishbone_bd_ram_mem2_reg[144][21]/P0001 , \wishbone_bd_ram_mem2_reg[144][22]/P0001 , \wishbone_bd_ram_mem2_reg[144][23]/P0001 , \wishbone_bd_ram_mem2_reg[145][16]/P0001 , \wishbone_bd_ram_mem2_reg[145][17]/P0001 , \wishbone_bd_ram_mem2_reg[145][18]/P0001 , \wishbone_bd_ram_mem2_reg[145][19]/P0001 , \wishbone_bd_ram_mem2_reg[145][20]/P0001 , \wishbone_bd_ram_mem2_reg[145][21]/P0001 , \wishbone_bd_ram_mem2_reg[145][22]/P0001 , \wishbone_bd_ram_mem2_reg[145][23]/P0001 , \wishbone_bd_ram_mem2_reg[146][16]/P0001 , \wishbone_bd_ram_mem2_reg[146][17]/P0001 , \wishbone_bd_ram_mem2_reg[146][18]/P0001 , \wishbone_bd_ram_mem2_reg[146][19]/P0001 , \wishbone_bd_ram_mem2_reg[146][20]/P0001 , \wishbone_bd_ram_mem2_reg[146][21]/P0001 , \wishbone_bd_ram_mem2_reg[146][22]/P0001 , \wishbone_bd_ram_mem2_reg[146][23]/P0001 , \wishbone_bd_ram_mem2_reg[147][16]/P0001 , \wishbone_bd_ram_mem2_reg[147][17]/P0001 , \wishbone_bd_ram_mem2_reg[147][18]/P0001 , \wishbone_bd_ram_mem2_reg[147][19]/P0001 , \wishbone_bd_ram_mem2_reg[147][20]/P0001 , \wishbone_bd_ram_mem2_reg[147][21]/P0001 , \wishbone_bd_ram_mem2_reg[147][22]/P0001 , \wishbone_bd_ram_mem2_reg[147][23]/P0001 , \wishbone_bd_ram_mem2_reg[148][16]/P0001 , \wishbone_bd_ram_mem2_reg[148][17]/P0001 , \wishbone_bd_ram_mem2_reg[148][18]/P0001 , \wishbone_bd_ram_mem2_reg[148][19]/P0001 , \wishbone_bd_ram_mem2_reg[148][20]/P0001 , \wishbone_bd_ram_mem2_reg[148][21]/P0001 , \wishbone_bd_ram_mem2_reg[148][22]/P0001 , \wishbone_bd_ram_mem2_reg[148][23]/P0001 , \wishbone_bd_ram_mem2_reg[149][16]/P0001 , \wishbone_bd_ram_mem2_reg[149][17]/P0001 , \wishbone_bd_ram_mem2_reg[149][18]/P0001 , \wishbone_bd_ram_mem2_reg[149][19]/P0001 , \wishbone_bd_ram_mem2_reg[149][20]/P0001 , \wishbone_bd_ram_mem2_reg[149][21]/P0001 , \wishbone_bd_ram_mem2_reg[149][22]/P0001 , \wishbone_bd_ram_mem2_reg[149][23]/P0001 , \wishbone_bd_ram_mem2_reg[14][16]/P0001 , \wishbone_bd_ram_mem2_reg[14][17]/P0001 , \wishbone_bd_ram_mem2_reg[14][18]/P0001 , \wishbone_bd_ram_mem2_reg[14][19]/P0001 , \wishbone_bd_ram_mem2_reg[14][20]/P0001 , \wishbone_bd_ram_mem2_reg[14][21]/P0001 , \wishbone_bd_ram_mem2_reg[14][22]/P0001 , \wishbone_bd_ram_mem2_reg[14][23]/P0001 , \wishbone_bd_ram_mem2_reg[150][16]/P0001 , \wishbone_bd_ram_mem2_reg[150][17]/P0001 , \wishbone_bd_ram_mem2_reg[150][18]/P0001 , \wishbone_bd_ram_mem2_reg[150][19]/P0001 , \wishbone_bd_ram_mem2_reg[150][20]/P0001 , \wishbone_bd_ram_mem2_reg[150][21]/P0001 , \wishbone_bd_ram_mem2_reg[150][22]/P0001 , \wishbone_bd_ram_mem2_reg[150][23]/P0001 , \wishbone_bd_ram_mem2_reg[151][16]/P0001 , \wishbone_bd_ram_mem2_reg[151][17]/P0001 , \wishbone_bd_ram_mem2_reg[151][18]/P0001 , \wishbone_bd_ram_mem2_reg[151][19]/P0001 , \wishbone_bd_ram_mem2_reg[151][20]/P0001 , \wishbone_bd_ram_mem2_reg[151][21]/P0001 , \wishbone_bd_ram_mem2_reg[151][22]/P0001 , \wishbone_bd_ram_mem2_reg[151][23]/P0001 , \wishbone_bd_ram_mem2_reg[152][16]/P0001 , \wishbone_bd_ram_mem2_reg[152][17]/P0001 , \wishbone_bd_ram_mem2_reg[152][18]/P0001 , \wishbone_bd_ram_mem2_reg[152][19]/P0001 , \wishbone_bd_ram_mem2_reg[152][20]/P0001 , \wishbone_bd_ram_mem2_reg[152][21]/P0001 , \wishbone_bd_ram_mem2_reg[152][22]/P0001 , \wishbone_bd_ram_mem2_reg[152][23]/P0001 , \wishbone_bd_ram_mem2_reg[153][16]/P0001 , \wishbone_bd_ram_mem2_reg[153][17]/P0001 , \wishbone_bd_ram_mem2_reg[153][18]/P0001 , \wishbone_bd_ram_mem2_reg[153][19]/P0001 , \wishbone_bd_ram_mem2_reg[153][20]/P0001 , \wishbone_bd_ram_mem2_reg[153][21]/P0001 , \wishbone_bd_ram_mem2_reg[153][22]/P0001 , \wishbone_bd_ram_mem2_reg[153][23]/P0001 , \wishbone_bd_ram_mem2_reg[154][16]/P0001 , \wishbone_bd_ram_mem2_reg[154][17]/P0001 , \wishbone_bd_ram_mem2_reg[154][18]/P0001 , \wishbone_bd_ram_mem2_reg[154][19]/P0001 , \wishbone_bd_ram_mem2_reg[154][20]/P0001 , \wishbone_bd_ram_mem2_reg[154][21]/P0001 , \wishbone_bd_ram_mem2_reg[154][22]/P0001 , \wishbone_bd_ram_mem2_reg[154][23]/P0001 , \wishbone_bd_ram_mem2_reg[155][16]/P0001 , \wishbone_bd_ram_mem2_reg[155][17]/P0001 , \wishbone_bd_ram_mem2_reg[155][18]/P0001 , \wishbone_bd_ram_mem2_reg[155][19]/P0001 , \wishbone_bd_ram_mem2_reg[155][20]/P0001 , \wishbone_bd_ram_mem2_reg[155][21]/P0001 , \wishbone_bd_ram_mem2_reg[155][22]/P0001 , \wishbone_bd_ram_mem2_reg[155][23]/P0001 , \wishbone_bd_ram_mem2_reg[156][16]/P0001 , \wishbone_bd_ram_mem2_reg[156][17]/P0001 , \wishbone_bd_ram_mem2_reg[156][18]/P0001 , \wishbone_bd_ram_mem2_reg[156][19]/P0001 , \wishbone_bd_ram_mem2_reg[156][20]/P0001 , \wishbone_bd_ram_mem2_reg[156][21]/P0001 , \wishbone_bd_ram_mem2_reg[156][22]/P0001 , \wishbone_bd_ram_mem2_reg[156][23]/P0001 , \wishbone_bd_ram_mem2_reg[157][16]/P0001 , \wishbone_bd_ram_mem2_reg[157][17]/P0001 , \wishbone_bd_ram_mem2_reg[157][18]/P0001 , \wishbone_bd_ram_mem2_reg[157][19]/P0001 , \wishbone_bd_ram_mem2_reg[157][20]/P0001 , \wishbone_bd_ram_mem2_reg[157][21]/P0001 , \wishbone_bd_ram_mem2_reg[157][22]/P0001 , \wishbone_bd_ram_mem2_reg[157][23]/P0001 , \wishbone_bd_ram_mem2_reg[158][16]/P0001 , \wishbone_bd_ram_mem2_reg[158][17]/P0001 , \wishbone_bd_ram_mem2_reg[158][18]/P0001 , \wishbone_bd_ram_mem2_reg[158][19]/P0001 , \wishbone_bd_ram_mem2_reg[158][20]/P0001 , \wishbone_bd_ram_mem2_reg[158][21]/P0001 , \wishbone_bd_ram_mem2_reg[158][22]/P0001 , \wishbone_bd_ram_mem2_reg[158][23]/P0001 , \wishbone_bd_ram_mem2_reg[159][16]/P0001 , \wishbone_bd_ram_mem2_reg[159][17]/P0001 , \wishbone_bd_ram_mem2_reg[159][18]/P0001 , \wishbone_bd_ram_mem2_reg[159][19]/P0001 , \wishbone_bd_ram_mem2_reg[159][20]/P0001 , \wishbone_bd_ram_mem2_reg[159][21]/P0001 , \wishbone_bd_ram_mem2_reg[159][22]/P0001 , \wishbone_bd_ram_mem2_reg[159][23]/P0001 , \wishbone_bd_ram_mem2_reg[15][16]/P0001 , \wishbone_bd_ram_mem2_reg[15][17]/P0001 , \wishbone_bd_ram_mem2_reg[15][18]/P0001 , \wishbone_bd_ram_mem2_reg[15][19]/P0001 , \wishbone_bd_ram_mem2_reg[15][20]/P0001 , \wishbone_bd_ram_mem2_reg[15][21]/P0001 , \wishbone_bd_ram_mem2_reg[15][22]/P0001 , \wishbone_bd_ram_mem2_reg[15][23]/P0001 , \wishbone_bd_ram_mem2_reg[160][16]/P0001 , \wishbone_bd_ram_mem2_reg[160][17]/P0001 , \wishbone_bd_ram_mem2_reg[160][18]/P0001 , \wishbone_bd_ram_mem2_reg[160][19]/P0001 , \wishbone_bd_ram_mem2_reg[160][20]/P0001 , \wishbone_bd_ram_mem2_reg[160][21]/P0001 , \wishbone_bd_ram_mem2_reg[160][22]/P0001 , \wishbone_bd_ram_mem2_reg[160][23]/P0001 , \wishbone_bd_ram_mem2_reg[161][16]/P0001 , \wishbone_bd_ram_mem2_reg[161][17]/P0001 , \wishbone_bd_ram_mem2_reg[161][18]/P0001 , \wishbone_bd_ram_mem2_reg[161][19]/P0001 , \wishbone_bd_ram_mem2_reg[161][20]/P0001 , \wishbone_bd_ram_mem2_reg[161][21]/P0001 , \wishbone_bd_ram_mem2_reg[161][22]/P0001 , \wishbone_bd_ram_mem2_reg[161][23]/P0001 , \wishbone_bd_ram_mem2_reg[162][16]/P0001 , \wishbone_bd_ram_mem2_reg[162][17]/P0001 , \wishbone_bd_ram_mem2_reg[162][18]/P0001 , \wishbone_bd_ram_mem2_reg[162][19]/P0001 , \wishbone_bd_ram_mem2_reg[162][20]/P0001 , \wishbone_bd_ram_mem2_reg[162][21]/P0001 , \wishbone_bd_ram_mem2_reg[162][22]/P0001 , \wishbone_bd_ram_mem2_reg[162][23]/P0001 , \wishbone_bd_ram_mem2_reg[163][16]/P0001 , \wishbone_bd_ram_mem2_reg[163][17]/P0001 , \wishbone_bd_ram_mem2_reg[163][18]/P0001 , \wishbone_bd_ram_mem2_reg[163][19]/P0001 , \wishbone_bd_ram_mem2_reg[163][20]/P0001 , \wishbone_bd_ram_mem2_reg[163][21]/P0001 , \wishbone_bd_ram_mem2_reg[163][22]/P0001 , \wishbone_bd_ram_mem2_reg[163][23]/P0001 , \wishbone_bd_ram_mem2_reg[164][16]/P0001 , \wishbone_bd_ram_mem2_reg[164][17]/P0001 , \wishbone_bd_ram_mem2_reg[164][18]/P0001 , \wishbone_bd_ram_mem2_reg[164][19]/P0001 , \wishbone_bd_ram_mem2_reg[164][20]/P0001 , \wishbone_bd_ram_mem2_reg[164][21]/P0001 , \wishbone_bd_ram_mem2_reg[164][22]/P0001 , \wishbone_bd_ram_mem2_reg[164][23]/P0001 , \wishbone_bd_ram_mem2_reg[165][16]/P0001 , \wishbone_bd_ram_mem2_reg[165][17]/P0001 , \wishbone_bd_ram_mem2_reg[165][18]/P0001 , \wishbone_bd_ram_mem2_reg[165][19]/P0001 , \wishbone_bd_ram_mem2_reg[165][20]/P0001 , \wishbone_bd_ram_mem2_reg[165][21]/P0001 , \wishbone_bd_ram_mem2_reg[165][22]/P0001 , \wishbone_bd_ram_mem2_reg[165][23]/P0001 , \wishbone_bd_ram_mem2_reg[166][16]/P0001 , \wishbone_bd_ram_mem2_reg[166][17]/P0001 , \wishbone_bd_ram_mem2_reg[166][18]/P0001 , \wishbone_bd_ram_mem2_reg[166][19]/P0001 , \wishbone_bd_ram_mem2_reg[166][20]/P0001 , \wishbone_bd_ram_mem2_reg[166][21]/P0001 , \wishbone_bd_ram_mem2_reg[166][22]/P0001 , \wishbone_bd_ram_mem2_reg[166][23]/P0001 , \wishbone_bd_ram_mem2_reg[167][16]/P0001 , \wishbone_bd_ram_mem2_reg[167][17]/P0001 , \wishbone_bd_ram_mem2_reg[167][18]/P0001 , \wishbone_bd_ram_mem2_reg[167][19]/P0001 , \wishbone_bd_ram_mem2_reg[167][20]/P0001 , \wishbone_bd_ram_mem2_reg[167][21]/P0001 , \wishbone_bd_ram_mem2_reg[167][22]/P0001 , \wishbone_bd_ram_mem2_reg[167][23]/P0001 , \wishbone_bd_ram_mem2_reg[168][16]/P0001 , \wishbone_bd_ram_mem2_reg[168][17]/P0001 , \wishbone_bd_ram_mem2_reg[168][18]/P0001 , \wishbone_bd_ram_mem2_reg[168][19]/P0001 , \wishbone_bd_ram_mem2_reg[168][20]/P0001 , \wishbone_bd_ram_mem2_reg[168][21]/P0001 , \wishbone_bd_ram_mem2_reg[168][22]/P0001 , \wishbone_bd_ram_mem2_reg[168][23]/P0001 , \wishbone_bd_ram_mem2_reg[169][16]/P0001 , \wishbone_bd_ram_mem2_reg[169][17]/P0001 , \wishbone_bd_ram_mem2_reg[169][18]/P0001 , \wishbone_bd_ram_mem2_reg[169][19]/P0001 , \wishbone_bd_ram_mem2_reg[169][20]/P0001 , \wishbone_bd_ram_mem2_reg[169][21]/P0001 , \wishbone_bd_ram_mem2_reg[169][22]/P0001 , \wishbone_bd_ram_mem2_reg[169][23]/P0001 , \wishbone_bd_ram_mem2_reg[16][16]/P0001 , \wishbone_bd_ram_mem2_reg[16][17]/P0001 , \wishbone_bd_ram_mem2_reg[16][18]/P0001 , \wishbone_bd_ram_mem2_reg[16][19]/P0001 , \wishbone_bd_ram_mem2_reg[16][20]/P0001 , \wishbone_bd_ram_mem2_reg[16][21]/P0001 , \wishbone_bd_ram_mem2_reg[16][22]/P0001 , \wishbone_bd_ram_mem2_reg[16][23]/P0001 , \wishbone_bd_ram_mem2_reg[170][16]/P0001 , \wishbone_bd_ram_mem2_reg[170][17]/P0001 , \wishbone_bd_ram_mem2_reg[170][18]/P0001 , \wishbone_bd_ram_mem2_reg[170][19]/P0001 , \wishbone_bd_ram_mem2_reg[170][20]/P0001 , \wishbone_bd_ram_mem2_reg[170][21]/P0001 , \wishbone_bd_ram_mem2_reg[170][22]/P0001 , \wishbone_bd_ram_mem2_reg[170][23]/P0001 , \wishbone_bd_ram_mem2_reg[171][16]/P0001 , \wishbone_bd_ram_mem2_reg[171][17]/P0001 , \wishbone_bd_ram_mem2_reg[171][18]/P0001 , \wishbone_bd_ram_mem2_reg[171][19]/P0001 , \wishbone_bd_ram_mem2_reg[171][20]/P0001 , \wishbone_bd_ram_mem2_reg[171][21]/P0001 , \wishbone_bd_ram_mem2_reg[171][22]/P0001 , \wishbone_bd_ram_mem2_reg[171][23]/P0001 , \wishbone_bd_ram_mem2_reg[172][16]/P0001 , \wishbone_bd_ram_mem2_reg[172][17]/P0001 , \wishbone_bd_ram_mem2_reg[172][18]/P0001 , \wishbone_bd_ram_mem2_reg[172][19]/P0001 , \wishbone_bd_ram_mem2_reg[172][20]/P0001 , \wishbone_bd_ram_mem2_reg[172][21]/P0001 , \wishbone_bd_ram_mem2_reg[172][22]/P0001 , \wishbone_bd_ram_mem2_reg[172][23]/P0001 , \wishbone_bd_ram_mem2_reg[173][16]/P0001 , \wishbone_bd_ram_mem2_reg[173][17]/P0001 , \wishbone_bd_ram_mem2_reg[173][18]/P0001 , \wishbone_bd_ram_mem2_reg[173][19]/P0001 , \wishbone_bd_ram_mem2_reg[173][20]/P0001 , \wishbone_bd_ram_mem2_reg[173][21]/P0001 , \wishbone_bd_ram_mem2_reg[173][22]/P0001 , \wishbone_bd_ram_mem2_reg[173][23]/P0001 , \wishbone_bd_ram_mem2_reg[174][16]/P0001 , \wishbone_bd_ram_mem2_reg[174][17]/P0001 , \wishbone_bd_ram_mem2_reg[174][18]/P0001 , \wishbone_bd_ram_mem2_reg[174][19]/P0001 , \wishbone_bd_ram_mem2_reg[174][20]/P0001 , \wishbone_bd_ram_mem2_reg[174][21]/P0001 , \wishbone_bd_ram_mem2_reg[174][22]/P0001 , \wishbone_bd_ram_mem2_reg[174][23]/P0001 , \wishbone_bd_ram_mem2_reg[175][16]/P0001 , \wishbone_bd_ram_mem2_reg[175][17]/P0001 , \wishbone_bd_ram_mem2_reg[175][18]/P0001 , \wishbone_bd_ram_mem2_reg[175][19]/P0001 , \wishbone_bd_ram_mem2_reg[175][20]/P0001 , \wishbone_bd_ram_mem2_reg[175][21]/P0001 , \wishbone_bd_ram_mem2_reg[175][22]/P0001 , \wishbone_bd_ram_mem2_reg[175][23]/P0001 , \wishbone_bd_ram_mem2_reg[176][16]/P0001 , \wishbone_bd_ram_mem2_reg[176][17]/P0001 , \wishbone_bd_ram_mem2_reg[176][18]/P0001 , \wishbone_bd_ram_mem2_reg[176][19]/P0001 , \wishbone_bd_ram_mem2_reg[176][20]/P0001 , \wishbone_bd_ram_mem2_reg[176][21]/P0001 , \wishbone_bd_ram_mem2_reg[176][22]/P0001 , \wishbone_bd_ram_mem2_reg[176][23]/P0001 , \wishbone_bd_ram_mem2_reg[177][16]/P0001 , \wishbone_bd_ram_mem2_reg[177][17]/P0001 , \wishbone_bd_ram_mem2_reg[177][18]/P0001 , \wishbone_bd_ram_mem2_reg[177][19]/P0001 , \wishbone_bd_ram_mem2_reg[177][20]/P0001 , \wishbone_bd_ram_mem2_reg[177][21]/P0001 , \wishbone_bd_ram_mem2_reg[177][22]/P0001 , \wishbone_bd_ram_mem2_reg[177][23]/P0001 , \wishbone_bd_ram_mem2_reg[178][16]/P0001 , \wishbone_bd_ram_mem2_reg[178][17]/P0001 , \wishbone_bd_ram_mem2_reg[178][18]/P0001 , \wishbone_bd_ram_mem2_reg[178][19]/P0001 , \wishbone_bd_ram_mem2_reg[178][20]/P0001 , \wishbone_bd_ram_mem2_reg[178][21]/P0001 , \wishbone_bd_ram_mem2_reg[178][22]/P0001 , \wishbone_bd_ram_mem2_reg[178][23]/P0001 , \wishbone_bd_ram_mem2_reg[179][16]/P0001 , \wishbone_bd_ram_mem2_reg[179][17]/P0001 , \wishbone_bd_ram_mem2_reg[179][18]/P0001 , \wishbone_bd_ram_mem2_reg[179][19]/P0001 , \wishbone_bd_ram_mem2_reg[179][20]/P0001 , \wishbone_bd_ram_mem2_reg[179][21]/P0001 , \wishbone_bd_ram_mem2_reg[179][22]/P0001 , \wishbone_bd_ram_mem2_reg[179][23]/P0001 , \wishbone_bd_ram_mem2_reg[17][16]/P0001 , \wishbone_bd_ram_mem2_reg[17][17]/P0001 , \wishbone_bd_ram_mem2_reg[17][18]/P0001 , \wishbone_bd_ram_mem2_reg[17][19]/P0001 , \wishbone_bd_ram_mem2_reg[17][20]/P0001 , \wishbone_bd_ram_mem2_reg[17][21]/P0001 , \wishbone_bd_ram_mem2_reg[17][22]/P0001 , \wishbone_bd_ram_mem2_reg[17][23]/P0001 , \wishbone_bd_ram_mem2_reg[180][16]/P0001 , \wishbone_bd_ram_mem2_reg[180][17]/P0001 , \wishbone_bd_ram_mem2_reg[180][18]/P0001 , \wishbone_bd_ram_mem2_reg[180][19]/P0001 , \wishbone_bd_ram_mem2_reg[180][20]/P0001 , \wishbone_bd_ram_mem2_reg[180][21]/P0001 , \wishbone_bd_ram_mem2_reg[180][22]/P0001 , \wishbone_bd_ram_mem2_reg[180][23]/P0001 , \wishbone_bd_ram_mem2_reg[181][16]/P0001 , \wishbone_bd_ram_mem2_reg[181][17]/P0001 , \wishbone_bd_ram_mem2_reg[181][18]/P0001 , \wishbone_bd_ram_mem2_reg[181][19]/P0001 , \wishbone_bd_ram_mem2_reg[181][20]/P0001 , \wishbone_bd_ram_mem2_reg[181][21]/P0001 , \wishbone_bd_ram_mem2_reg[181][22]/P0001 , \wishbone_bd_ram_mem2_reg[181][23]/P0001 , \wishbone_bd_ram_mem2_reg[182][16]/P0001 , \wishbone_bd_ram_mem2_reg[182][17]/P0001 , \wishbone_bd_ram_mem2_reg[182][18]/P0001 , \wishbone_bd_ram_mem2_reg[182][19]/P0001 , \wishbone_bd_ram_mem2_reg[182][20]/P0001 , \wishbone_bd_ram_mem2_reg[182][21]/P0001 , \wishbone_bd_ram_mem2_reg[182][22]/P0001 , \wishbone_bd_ram_mem2_reg[182][23]/P0001 , \wishbone_bd_ram_mem2_reg[183][16]/P0001 , \wishbone_bd_ram_mem2_reg[183][17]/P0001 , \wishbone_bd_ram_mem2_reg[183][18]/P0001 , \wishbone_bd_ram_mem2_reg[183][19]/P0001 , \wishbone_bd_ram_mem2_reg[183][20]/P0001 , \wishbone_bd_ram_mem2_reg[183][21]/P0001 , \wishbone_bd_ram_mem2_reg[183][22]/P0001 , \wishbone_bd_ram_mem2_reg[183][23]/P0001 , \wishbone_bd_ram_mem2_reg[184][16]/P0001 , \wishbone_bd_ram_mem2_reg[184][17]/P0001 , \wishbone_bd_ram_mem2_reg[184][18]/P0001 , \wishbone_bd_ram_mem2_reg[184][19]/P0001 , \wishbone_bd_ram_mem2_reg[184][20]/P0001 , \wishbone_bd_ram_mem2_reg[184][21]/P0001 , \wishbone_bd_ram_mem2_reg[184][22]/P0001 , \wishbone_bd_ram_mem2_reg[184][23]/P0001 , \wishbone_bd_ram_mem2_reg[185][16]/P0001 , \wishbone_bd_ram_mem2_reg[185][17]/P0001 , \wishbone_bd_ram_mem2_reg[185][18]/P0001 , \wishbone_bd_ram_mem2_reg[185][19]/P0001 , \wishbone_bd_ram_mem2_reg[185][20]/P0001 , \wishbone_bd_ram_mem2_reg[185][21]/P0001 , \wishbone_bd_ram_mem2_reg[185][22]/P0001 , \wishbone_bd_ram_mem2_reg[185][23]/P0001 , \wishbone_bd_ram_mem2_reg[186][16]/P0001 , \wishbone_bd_ram_mem2_reg[186][17]/P0001 , \wishbone_bd_ram_mem2_reg[186][18]/P0001 , \wishbone_bd_ram_mem2_reg[186][19]/P0001 , \wishbone_bd_ram_mem2_reg[186][20]/P0001 , \wishbone_bd_ram_mem2_reg[186][21]/P0001 , \wishbone_bd_ram_mem2_reg[186][22]/P0001 , \wishbone_bd_ram_mem2_reg[186][23]/P0001 , \wishbone_bd_ram_mem2_reg[187][16]/P0001 , \wishbone_bd_ram_mem2_reg[187][17]/P0001 , \wishbone_bd_ram_mem2_reg[187][18]/P0001 , \wishbone_bd_ram_mem2_reg[187][19]/P0001 , \wishbone_bd_ram_mem2_reg[187][20]/P0001 , \wishbone_bd_ram_mem2_reg[187][21]/P0001 , \wishbone_bd_ram_mem2_reg[187][22]/P0001 , \wishbone_bd_ram_mem2_reg[187][23]/P0001 , \wishbone_bd_ram_mem2_reg[188][16]/P0001 , \wishbone_bd_ram_mem2_reg[188][17]/P0001 , \wishbone_bd_ram_mem2_reg[188][18]/P0001 , \wishbone_bd_ram_mem2_reg[188][19]/P0001 , \wishbone_bd_ram_mem2_reg[188][20]/P0001 , \wishbone_bd_ram_mem2_reg[188][21]/P0001 , \wishbone_bd_ram_mem2_reg[188][22]/P0001 , \wishbone_bd_ram_mem2_reg[188][23]/P0001 , \wishbone_bd_ram_mem2_reg[189][16]/P0001 , \wishbone_bd_ram_mem2_reg[189][17]/P0001 , \wishbone_bd_ram_mem2_reg[189][18]/P0001 , \wishbone_bd_ram_mem2_reg[189][19]/P0001 , \wishbone_bd_ram_mem2_reg[189][20]/P0001 , \wishbone_bd_ram_mem2_reg[189][21]/P0001 , \wishbone_bd_ram_mem2_reg[189][22]/P0001 , \wishbone_bd_ram_mem2_reg[189][23]/P0001 , \wishbone_bd_ram_mem2_reg[18][16]/P0001 , \wishbone_bd_ram_mem2_reg[18][17]/P0001 , \wishbone_bd_ram_mem2_reg[18][18]/P0001 , \wishbone_bd_ram_mem2_reg[18][19]/P0001 , \wishbone_bd_ram_mem2_reg[18][20]/P0001 , \wishbone_bd_ram_mem2_reg[18][21]/P0001 , \wishbone_bd_ram_mem2_reg[18][22]/P0001 , \wishbone_bd_ram_mem2_reg[18][23]/P0001 , \wishbone_bd_ram_mem2_reg[190][16]/P0001 , \wishbone_bd_ram_mem2_reg[190][17]/P0001 , \wishbone_bd_ram_mem2_reg[190][18]/P0001 , \wishbone_bd_ram_mem2_reg[190][19]/P0001 , \wishbone_bd_ram_mem2_reg[190][20]/P0001 , \wishbone_bd_ram_mem2_reg[190][21]/P0001 , \wishbone_bd_ram_mem2_reg[190][22]/P0001 , \wishbone_bd_ram_mem2_reg[190][23]/P0001 , \wishbone_bd_ram_mem2_reg[191][16]/P0001 , \wishbone_bd_ram_mem2_reg[191][17]/P0001 , \wishbone_bd_ram_mem2_reg[191][18]/P0001 , \wishbone_bd_ram_mem2_reg[191][19]/P0001 , \wishbone_bd_ram_mem2_reg[191][20]/P0001 , \wishbone_bd_ram_mem2_reg[191][21]/P0001 , \wishbone_bd_ram_mem2_reg[191][22]/P0001 , \wishbone_bd_ram_mem2_reg[191][23]/P0001 , \wishbone_bd_ram_mem2_reg[192][16]/P0001 , \wishbone_bd_ram_mem2_reg[192][17]/P0001 , \wishbone_bd_ram_mem2_reg[192][18]/P0001 , \wishbone_bd_ram_mem2_reg[192][19]/P0001 , \wishbone_bd_ram_mem2_reg[192][20]/P0001 , \wishbone_bd_ram_mem2_reg[192][21]/P0001 , \wishbone_bd_ram_mem2_reg[192][22]/P0001 , \wishbone_bd_ram_mem2_reg[192][23]/P0001 , \wishbone_bd_ram_mem2_reg[193][16]/P0001 , \wishbone_bd_ram_mem2_reg[193][17]/P0001 , \wishbone_bd_ram_mem2_reg[193][18]/P0001 , \wishbone_bd_ram_mem2_reg[193][19]/P0001 , \wishbone_bd_ram_mem2_reg[193][20]/P0001 , \wishbone_bd_ram_mem2_reg[193][21]/P0001 , \wishbone_bd_ram_mem2_reg[193][22]/P0001 , \wishbone_bd_ram_mem2_reg[193][23]/P0001 , \wishbone_bd_ram_mem2_reg[194][16]/P0001 , \wishbone_bd_ram_mem2_reg[194][17]/P0001 , \wishbone_bd_ram_mem2_reg[194][18]/P0001 , \wishbone_bd_ram_mem2_reg[194][19]/P0001 , \wishbone_bd_ram_mem2_reg[194][20]/P0001 , \wishbone_bd_ram_mem2_reg[194][21]/P0001 , \wishbone_bd_ram_mem2_reg[194][22]/P0001 , \wishbone_bd_ram_mem2_reg[194][23]/P0001 , \wishbone_bd_ram_mem2_reg[195][16]/P0001 , \wishbone_bd_ram_mem2_reg[195][17]/P0001 , \wishbone_bd_ram_mem2_reg[195][18]/P0001 , \wishbone_bd_ram_mem2_reg[195][19]/P0001 , \wishbone_bd_ram_mem2_reg[195][20]/P0001 , \wishbone_bd_ram_mem2_reg[195][21]/P0001 , \wishbone_bd_ram_mem2_reg[195][22]/P0001 , \wishbone_bd_ram_mem2_reg[195][23]/P0001 , \wishbone_bd_ram_mem2_reg[196][16]/P0001 , \wishbone_bd_ram_mem2_reg[196][17]/P0001 , \wishbone_bd_ram_mem2_reg[196][18]/P0001 , \wishbone_bd_ram_mem2_reg[196][19]/P0001 , \wishbone_bd_ram_mem2_reg[196][20]/P0001 , \wishbone_bd_ram_mem2_reg[196][21]/P0001 , \wishbone_bd_ram_mem2_reg[196][22]/P0001 , \wishbone_bd_ram_mem2_reg[196][23]/P0001 , \wishbone_bd_ram_mem2_reg[197][16]/P0001 , \wishbone_bd_ram_mem2_reg[197][17]/P0001 , \wishbone_bd_ram_mem2_reg[197][18]/P0001 , \wishbone_bd_ram_mem2_reg[197][19]/P0001 , \wishbone_bd_ram_mem2_reg[197][20]/P0001 , \wishbone_bd_ram_mem2_reg[197][21]/P0001 , \wishbone_bd_ram_mem2_reg[197][22]/P0001 , \wishbone_bd_ram_mem2_reg[197][23]/P0001 , \wishbone_bd_ram_mem2_reg[198][16]/P0001 , \wishbone_bd_ram_mem2_reg[198][17]/P0001 , \wishbone_bd_ram_mem2_reg[198][18]/P0001 , \wishbone_bd_ram_mem2_reg[198][19]/P0001 , \wishbone_bd_ram_mem2_reg[198][20]/P0001 , \wishbone_bd_ram_mem2_reg[198][21]/P0001 , \wishbone_bd_ram_mem2_reg[198][22]/P0001 , \wishbone_bd_ram_mem2_reg[198][23]/P0001 , \wishbone_bd_ram_mem2_reg[199][16]/P0001 , \wishbone_bd_ram_mem2_reg[199][17]/P0001 , \wishbone_bd_ram_mem2_reg[199][18]/P0001 , \wishbone_bd_ram_mem2_reg[199][19]/P0001 , \wishbone_bd_ram_mem2_reg[199][20]/P0001 , \wishbone_bd_ram_mem2_reg[199][21]/P0001 , \wishbone_bd_ram_mem2_reg[199][22]/P0001 , \wishbone_bd_ram_mem2_reg[199][23]/P0001 , \wishbone_bd_ram_mem2_reg[19][16]/P0001 , \wishbone_bd_ram_mem2_reg[19][17]/P0001 , \wishbone_bd_ram_mem2_reg[19][18]/P0001 , \wishbone_bd_ram_mem2_reg[19][19]/P0001 , \wishbone_bd_ram_mem2_reg[19][20]/P0001 , \wishbone_bd_ram_mem2_reg[19][21]/P0001 , \wishbone_bd_ram_mem2_reg[19][22]/P0001 , \wishbone_bd_ram_mem2_reg[19][23]/P0001 , \wishbone_bd_ram_mem2_reg[1][16]/P0001 , \wishbone_bd_ram_mem2_reg[1][17]/P0001 , \wishbone_bd_ram_mem2_reg[1][18]/P0001 , \wishbone_bd_ram_mem2_reg[1][19]/P0001 , \wishbone_bd_ram_mem2_reg[1][20]/P0001 , \wishbone_bd_ram_mem2_reg[1][21]/P0001 , \wishbone_bd_ram_mem2_reg[1][22]/P0001 , \wishbone_bd_ram_mem2_reg[1][23]/P0001 , \wishbone_bd_ram_mem2_reg[200][16]/P0001 , \wishbone_bd_ram_mem2_reg[200][17]/P0001 , \wishbone_bd_ram_mem2_reg[200][18]/P0001 , \wishbone_bd_ram_mem2_reg[200][19]/P0001 , \wishbone_bd_ram_mem2_reg[200][20]/P0001 , \wishbone_bd_ram_mem2_reg[200][21]/P0001 , \wishbone_bd_ram_mem2_reg[200][22]/P0001 , \wishbone_bd_ram_mem2_reg[200][23]/P0001 , \wishbone_bd_ram_mem2_reg[201][16]/P0001 , \wishbone_bd_ram_mem2_reg[201][17]/P0001 , \wishbone_bd_ram_mem2_reg[201][18]/P0001 , \wishbone_bd_ram_mem2_reg[201][19]/P0001 , \wishbone_bd_ram_mem2_reg[201][20]/P0001 , \wishbone_bd_ram_mem2_reg[201][21]/P0001 , \wishbone_bd_ram_mem2_reg[201][22]/P0001 , \wishbone_bd_ram_mem2_reg[201][23]/P0001 , \wishbone_bd_ram_mem2_reg[202][16]/P0001 , \wishbone_bd_ram_mem2_reg[202][17]/P0001 , \wishbone_bd_ram_mem2_reg[202][18]/P0001 , \wishbone_bd_ram_mem2_reg[202][19]/P0001 , \wishbone_bd_ram_mem2_reg[202][20]/P0001 , \wishbone_bd_ram_mem2_reg[202][21]/P0001 , \wishbone_bd_ram_mem2_reg[202][22]/P0001 , \wishbone_bd_ram_mem2_reg[202][23]/P0001 , \wishbone_bd_ram_mem2_reg[203][16]/P0001 , \wishbone_bd_ram_mem2_reg[203][17]/P0001 , \wishbone_bd_ram_mem2_reg[203][18]/P0001 , \wishbone_bd_ram_mem2_reg[203][19]/P0001 , \wishbone_bd_ram_mem2_reg[203][20]/P0001 , \wishbone_bd_ram_mem2_reg[203][21]/P0001 , \wishbone_bd_ram_mem2_reg[203][22]/P0001 , \wishbone_bd_ram_mem2_reg[203][23]/P0001 , \wishbone_bd_ram_mem2_reg[204][16]/P0001 , \wishbone_bd_ram_mem2_reg[204][17]/P0001 , \wishbone_bd_ram_mem2_reg[204][18]/P0001 , \wishbone_bd_ram_mem2_reg[204][19]/P0001 , \wishbone_bd_ram_mem2_reg[204][20]/P0001 , \wishbone_bd_ram_mem2_reg[204][21]/P0001 , \wishbone_bd_ram_mem2_reg[204][22]/P0001 , \wishbone_bd_ram_mem2_reg[204][23]/P0001 , \wishbone_bd_ram_mem2_reg[205][16]/P0001 , \wishbone_bd_ram_mem2_reg[205][17]/P0001 , \wishbone_bd_ram_mem2_reg[205][18]/P0001 , \wishbone_bd_ram_mem2_reg[205][19]/P0001 , \wishbone_bd_ram_mem2_reg[205][20]/P0001 , \wishbone_bd_ram_mem2_reg[205][21]/P0001 , \wishbone_bd_ram_mem2_reg[205][22]/P0001 , \wishbone_bd_ram_mem2_reg[205][23]/P0001 , \wishbone_bd_ram_mem2_reg[206][16]/P0001 , \wishbone_bd_ram_mem2_reg[206][17]/P0001 , \wishbone_bd_ram_mem2_reg[206][18]/P0001 , \wishbone_bd_ram_mem2_reg[206][19]/P0001 , \wishbone_bd_ram_mem2_reg[206][20]/P0001 , \wishbone_bd_ram_mem2_reg[206][21]/P0001 , \wishbone_bd_ram_mem2_reg[206][22]/P0001 , \wishbone_bd_ram_mem2_reg[206][23]/P0001 , \wishbone_bd_ram_mem2_reg[207][16]/P0001 , \wishbone_bd_ram_mem2_reg[207][17]/P0001 , \wishbone_bd_ram_mem2_reg[207][18]/P0001 , \wishbone_bd_ram_mem2_reg[207][19]/P0001 , \wishbone_bd_ram_mem2_reg[207][20]/P0001 , \wishbone_bd_ram_mem2_reg[207][21]/P0001 , \wishbone_bd_ram_mem2_reg[207][22]/P0001 , \wishbone_bd_ram_mem2_reg[207][23]/P0001 , \wishbone_bd_ram_mem2_reg[208][16]/P0001 , \wishbone_bd_ram_mem2_reg[208][17]/P0001 , \wishbone_bd_ram_mem2_reg[208][18]/P0001 , \wishbone_bd_ram_mem2_reg[208][19]/P0001 , \wishbone_bd_ram_mem2_reg[208][20]/P0001 , \wishbone_bd_ram_mem2_reg[208][21]/P0001 , \wishbone_bd_ram_mem2_reg[208][22]/P0001 , \wishbone_bd_ram_mem2_reg[208][23]/P0001 , \wishbone_bd_ram_mem2_reg[209][16]/P0001 , \wishbone_bd_ram_mem2_reg[209][17]/P0001 , \wishbone_bd_ram_mem2_reg[209][18]/P0001 , \wishbone_bd_ram_mem2_reg[209][19]/P0001 , \wishbone_bd_ram_mem2_reg[209][20]/P0001 , \wishbone_bd_ram_mem2_reg[209][21]/P0001 , \wishbone_bd_ram_mem2_reg[209][22]/P0001 , \wishbone_bd_ram_mem2_reg[209][23]/P0001 , \wishbone_bd_ram_mem2_reg[20][16]/P0001 , \wishbone_bd_ram_mem2_reg[20][17]/P0001 , \wishbone_bd_ram_mem2_reg[20][18]/P0001 , \wishbone_bd_ram_mem2_reg[20][19]/P0001 , \wishbone_bd_ram_mem2_reg[20][20]/P0001 , \wishbone_bd_ram_mem2_reg[20][21]/P0001 , \wishbone_bd_ram_mem2_reg[20][22]/P0001 , \wishbone_bd_ram_mem2_reg[20][23]/P0001 , \wishbone_bd_ram_mem2_reg[210][16]/P0001 , \wishbone_bd_ram_mem2_reg[210][17]/P0001 , \wishbone_bd_ram_mem2_reg[210][18]/P0001 , \wishbone_bd_ram_mem2_reg[210][19]/P0001 , \wishbone_bd_ram_mem2_reg[210][20]/P0001 , \wishbone_bd_ram_mem2_reg[210][21]/P0001 , \wishbone_bd_ram_mem2_reg[210][22]/P0001 , \wishbone_bd_ram_mem2_reg[210][23]/P0001 , \wishbone_bd_ram_mem2_reg[211][16]/P0001 , \wishbone_bd_ram_mem2_reg[211][17]/P0001 , \wishbone_bd_ram_mem2_reg[211][18]/P0001 , \wishbone_bd_ram_mem2_reg[211][19]/P0001 , \wishbone_bd_ram_mem2_reg[211][20]/P0001 , \wishbone_bd_ram_mem2_reg[211][21]/P0001 , \wishbone_bd_ram_mem2_reg[211][22]/P0001 , \wishbone_bd_ram_mem2_reg[211][23]/P0001 , \wishbone_bd_ram_mem2_reg[212][16]/P0001 , \wishbone_bd_ram_mem2_reg[212][17]/P0001 , \wishbone_bd_ram_mem2_reg[212][18]/P0001 , \wishbone_bd_ram_mem2_reg[212][19]/P0001 , \wishbone_bd_ram_mem2_reg[212][20]/P0001 , \wishbone_bd_ram_mem2_reg[212][21]/P0001 , \wishbone_bd_ram_mem2_reg[212][22]/P0001 , \wishbone_bd_ram_mem2_reg[212][23]/P0001 , \wishbone_bd_ram_mem2_reg[213][16]/P0001 , \wishbone_bd_ram_mem2_reg[213][17]/P0001 , \wishbone_bd_ram_mem2_reg[213][18]/P0001 , \wishbone_bd_ram_mem2_reg[213][19]/P0001 , \wishbone_bd_ram_mem2_reg[213][20]/P0001 , \wishbone_bd_ram_mem2_reg[213][21]/P0001 , \wishbone_bd_ram_mem2_reg[213][22]/P0001 , \wishbone_bd_ram_mem2_reg[213][23]/P0001 , \wishbone_bd_ram_mem2_reg[214][16]/P0001 , \wishbone_bd_ram_mem2_reg[214][17]/P0001 , \wishbone_bd_ram_mem2_reg[214][18]/P0001 , \wishbone_bd_ram_mem2_reg[214][19]/P0001 , \wishbone_bd_ram_mem2_reg[214][20]/P0001 , \wishbone_bd_ram_mem2_reg[214][21]/P0001 , \wishbone_bd_ram_mem2_reg[214][22]/P0001 , \wishbone_bd_ram_mem2_reg[214][23]/P0001 , \wishbone_bd_ram_mem2_reg[215][16]/P0001 , \wishbone_bd_ram_mem2_reg[215][17]/P0001 , \wishbone_bd_ram_mem2_reg[215][18]/P0001 , \wishbone_bd_ram_mem2_reg[215][19]/P0001 , \wishbone_bd_ram_mem2_reg[215][20]/P0001 , \wishbone_bd_ram_mem2_reg[215][21]/P0001 , \wishbone_bd_ram_mem2_reg[215][22]/P0001 , \wishbone_bd_ram_mem2_reg[215][23]/P0001 , \wishbone_bd_ram_mem2_reg[216][16]/P0001 , \wishbone_bd_ram_mem2_reg[216][17]/P0001 , \wishbone_bd_ram_mem2_reg[216][18]/P0001 , \wishbone_bd_ram_mem2_reg[216][19]/P0001 , \wishbone_bd_ram_mem2_reg[216][20]/P0001 , \wishbone_bd_ram_mem2_reg[216][21]/P0001 , \wishbone_bd_ram_mem2_reg[216][22]/P0001 , \wishbone_bd_ram_mem2_reg[216][23]/P0001 , \wishbone_bd_ram_mem2_reg[217][16]/P0001 , \wishbone_bd_ram_mem2_reg[217][17]/P0001 , \wishbone_bd_ram_mem2_reg[217][18]/P0001 , \wishbone_bd_ram_mem2_reg[217][19]/P0001 , \wishbone_bd_ram_mem2_reg[217][20]/P0001 , \wishbone_bd_ram_mem2_reg[217][21]/P0001 , \wishbone_bd_ram_mem2_reg[217][22]/P0001 , \wishbone_bd_ram_mem2_reg[217][23]/P0001 , \wishbone_bd_ram_mem2_reg[218][16]/P0001 , \wishbone_bd_ram_mem2_reg[218][17]/P0001 , \wishbone_bd_ram_mem2_reg[218][18]/P0001 , \wishbone_bd_ram_mem2_reg[218][19]/P0001 , \wishbone_bd_ram_mem2_reg[218][20]/P0001 , \wishbone_bd_ram_mem2_reg[218][21]/P0001 , \wishbone_bd_ram_mem2_reg[218][22]/P0001 , \wishbone_bd_ram_mem2_reg[218][23]/P0001 , \wishbone_bd_ram_mem2_reg[219][16]/P0001 , \wishbone_bd_ram_mem2_reg[219][17]/P0001 , \wishbone_bd_ram_mem2_reg[219][18]/P0001 , \wishbone_bd_ram_mem2_reg[219][19]/P0001 , \wishbone_bd_ram_mem2_reg[219][20]/P0001 , \wishbone_bd_ram_mem2_reg[219][21]/P0001 , \wishbone_bd_ram_mem2_reg[219][22]/P0001 , \wishbone_bd_ram_mem2_reg[219][23]/P0001 , \wishbone_bd_ram_mem2_reg[21][16]/P0001 , \wishbone_bd_ram_mem2_reg[21][17]/P0001 , \wishbone_bd_ram_mem2_reg[21][18]/P0001 , \wishbone_bd_ram_mem2_reg[21][19]/P0001 , \wishbone_bd_ram_mem2_reg[21][20]/P0001 , \wishbone_bd_ram_mem2_reg[21][21]/P0001 , \wishbone_bd_ram_mem2_reg[21][22]/P0001 , \wishbone_bd_ram_mem2_reg[21][23]/P0001 , \wishbone_bd_ram_mem2_reg[220][16]/P0001 , \wishbone_bd_ram_mem2_reg[220][17]/P0001 , \wishbone_bd_ram_mem2_reg[220][18]/P0001 , \wishbone_bd_ram_mem2_reg[220][19]/P0001 , \wishbone_bd_ram_mem2_reg[220][20]/P0001 , \wishbone_bd_ram_mem2_reg[220][21]/P0001 , \wishbone_bd_ram_mem2_reg[220][22]/P0001 , \wishbone_bd_ram_mem2_reg[220][23]/P0001 , \wishbone_bd_ram_mem2_reg[221][16]/P0001 , \wishbone_bd_ram_mem2_reg[221][17]/P0001 , \wishbone_bd_ram_mem2_reg[221][18]/P0001 , \wishbone_bd_ram_mem2_reg[221][19]/P0001 , \wishbone_bd_ram_mem2_reg[221][20]/P0001 , \wishbone_bd_ram_mem2_reg[221][21]/P0001 , \wishbone_bd_ram_mem2_reg[221][22]/P0001 , \wishbone_bd_ram_mem2_reg[221][23]/P0001 , \wishbone_bd_ram_mem2_reg[222][16]/P0001 , \wishbone_bd_ram_mem2_reg[222][17]/P0001 , \wishbone_bd_ram_mem2_reg[222][18]/P0001 , \wishbone_bd_ram_mem2_reg[222][19]/P0001 , \wishbone_bd_ram_mem2_reg[222][20]/P0001 , \wishbone_bd_ram_mem2_reg[222][21]/P0001 , \wishbone_bd_ram_mem2_reg[222][22]/P0001 , \wishbone_bd_ram_mem2_reg[222][23]/P0001 , \wishbone_bd_ram_mem2_reg[223][16]/P0001 , \wishbone_bd_ram_mem2_reg[223][17]/P0001 , \wishbone_bd_ram_mem2_reg[223][18]/P0001 , \wishbone_bd_ram_mem2_reg[223][19]/P0001 , \wishbone_bd_ram_mem2_reg[223][20]/P0001 , \wishbone_bd_ram_mem2_reg[223][21]/P0001 , \wishbone_bd_ram_mem2_reg[223][22]/P0001 , \wishbone_bd_ram_mem2_reg[223][23]/P0001 , \wishbone_bd_ram_mem2_reg[224][16]/P0001 , \wishbone_bd_ram_mem2_reg[224][17]/P0001 , \wishbone_bd_ram_mem2_reg[224][18]/P0001 , \wishbone_bd_ram_mem2_reg[224][19]/P0001 , \wishbone_bd_ram_mem2_reg[224][20]/P0001 , \wishbone_bd_ram_mem2_reg[224][21]/P0001 , \wishbone_bd_ram_mem2_reg[224][22]/P0001 , \wishbone_bd_ram_mem2_reg[224][23]/P0001 , \wishbone_bd_ram_mem2_reg[225][16]/P0001 , \wishbone_bd_ram_mem2_reg[225][17]/P0001 , \wishbone_bd_ram_mem2_reg[225][18]/P0001 , \wishbone_bd_ram_mem2_reg[225][19]/P0001 , \wishbone_bd_ram_mem2_reg[225][20]/P0001 , \wishbone_bd_ram_mem2_reg[225][21]/P0001 , \wishbone_bd_ram_mem2_reg[225][22]/P0001 , \wishbone_bd_ram_mem2_reg[225][23]/P0001 , \wishbone_bd_ram_mem2_reg[226][16]/P0001 , \wishbone_bd_ram_mem2_reg[226][17]/P0001 , \wishbone_bd_ram_mem2_reg[226][18]/P0001 , \wishbone_bd_ram_mem2_reg[226][19]/P0001 , \wishbone_bd_ram_mem2_reg[226][20]/P0001 , \wishbone_bd_ram_mem2_reg[226][21]/P0001 , \wishbone_bd_ram_mem2_reg[226][22]/P0001 , \wishbone_bd_ram_mem2_reg[226][23]/P0001 , \wishbone_bd_ram_mem2_reg[227][16]/P0001 , \wishbone_bd_ram_mem2_reg[227][17]/P0001 , \wishbone_bd_ram_mem2_reg[227][18]/P0001 , \wishbone_bd_ram_mem2_reg[227][19]/P0001 , \wishbone_bd_ram_mem2_reg[227][20]/P0001 , \wishbone_bd_ram_mem2_reg[227][21]/P0001 , \wishbone_bd_ram_mem2_reg[227][22]/P0001 , \wishbone_bd_ram_mem2_reg[227][23]/P0001 , \wishbone_bd_ram_mem2_reg[228][16]/P0001 , \wishbone_bd_ram_mem2_reg[228][17]/P0001 , \wishbone_bd_ram_mem2_reg[228][18]/P0001 , \wishbone_bd_ram_mem2_reg[228][19]/P0001 , \wishbone_bd_ram_mem2_reg[228][20]/P0001 , \wishbone_bd_ram_mem2_reg[228][21]/P0001 , \wishbone_bd_ram_mem2_reg[228][22]/P0001 , \wishbone_bd_ram_mem2_reg[228][23]/P0001 , \wishbone_bd_ram_mem2_reg[229][16]/P0001 , \wishbone_bd_ram_mem2_reg[229][17]/P0001 , \wishbone_bd_ram_mem2_reg[229][18]/P0001 , \wishbone_bd_ram_mem2_reg[229][19]/P0001 , \wishbone_bd_ram_mem2_reg[229][20]/P0001 , \wishbone_bd_ram_mem2_reg[229][21]/P0001 , \wishbone_bd_ram_mem2_reg[229][22]/P0001 , \wishbone_bd_ram_mem2_reg[229][23]/P0001 , \wishbone_bd_ram_mem2_reg[22][16]/P0001 , \wishbone_bd_ram_mem2_reg[22][17]/P0001 , \wishbone_bd_ram_mem2_reg[22][18]/P0001 , \wishbone_bd_ram_mem2_reg[22][19]/P0001 , \wishbone_bd_ram_mem2_reg[22][20]/P0001 , \wishbone_bd_ram_mem2_reg[22][21]/P0001 , \wishbone_bd_ram_mem2_reg[22][22]/P0001 , \wishbone_bd_ram_mem2_reg[22][23]/P0001 , \wishbone_bd_ram_mem2_reg[230][16]/P0001 , \wishbone_bd_ram_mem2_reg[230][17]/P0001 , \wishbone_bd_ram_mem2_reg[230][18]/P0001 , \wishbone_bd_ram_mem2_reg[230][19]/P0001 , \wishbone_bd_ram_mem2_reg[230][20]/P0001 , \wishbone_bd_ram_mem2_reg[230][21]/P0001 , \wishbone_bd_ram_mem2_reg[230][22]/P0001 , \wishbone_bd_ram_mem2_reg[230][23]/P0001 , \wishbone_bd_ram_mem2_reg[231][16]/P0001 , \wishbone_bd_ram_mem2_reg[231][17]/P0001 , \wishbone_bd_ram_mem2_reg[231][18]/P0001 , \wishbone_bd_ram_mem2_reg[231][19]/P0001 , \wishbone_bd_ram_mem2_reg[231][20]/P0001 , \wishbone_bd_ram_mem2_reg[231][21]/P0001 , \wishbone_bd_ram_mem2_reg[231][22]/P0001 , \wishbone_bd_ram_mem2_reg[231][23]/P0001 , \wishbone_bd_ram_mem2_reg[232][16]/P0001 , \wishbone_bd_ram_mem2_reg[232][17]/P0001 , \wishbone_bd_ram_mem2_reg[232][18]/P0001 , \wishbone_bd_ram_mem2_reg[232][19]/P0001 , \wishbone_bd_ram_mem2_reg[232][20]/P0001 , \wishbone_bd_ram_mem2_reg[232][21]/P0001 , \wishbone_bd_ram_mem2_reg[232][22]/P0001 , \wishbone_bd_ram_mem2_reg[232][23]/P0001 , \wishbone_bd_ram_mem2_reg[233][16]/P0001 , \wishbone_bd_ram_mem2_reg[233][17]/P0001 , \wishbone_bd_ram_mem2_reg[233][18]/P0001 , \wishbone_bd_ram_mem2_reg[233][19]/P0001 , \wishbone_bd_ram_mem2_reg[233][20]/P0001 , \wishbone_bd_ram_mem2_reg[233][21]/P0001 , \wishbone_bd_ram_mem2_reg[233][22]/P0001 , \wishbone_bd_ram_mem2_reg[233][23]/P0001 , \wishbone_bd_ram_mem2_reg[234][16]/P0001 , \wishbone_bd_ram_mem2_reg[234][17]/P0001 , \wishbone_bd_ram_mem2_reg[234][18]/P0001 , \wishbone_bd_ram_mem2_reg[234][19]/P0001 , \wishbone_bd_ram_mem2_reg[234][20]/P0001 , \wishbone_bd_ram_mem2_reg[234][21]/P0001 , \wishbone_bd_ram_mem2_reg[234][22]/P0001 , \wishbone_bd_ram_mem2_reg[234][23]/P0001 , \wishbone_bd_ram_mem2_reg[235][16]/P0001 , \wishbone_bd_ram_mem2_reg[235][17]/P0001 , \wishbone_bd_ram_mem2_reg[235][18]/P0001 , \wishbone_bd_ram_mem2_reg[235][19]/P0001 , \wishbone_bd_ram_mem2_reg[235][20]/P0001 , \wishbone_bd_ram_mem2_reg[235][21]/P0001 , \wishbone_bd_ram_mem2_reg[235][22]/P0001 , \wishbone_bd_ram_mem2_reg[235][23]/P0001 , \wishbone_bd_ram_mem2_reg[236][16]/P0001 , \wishbone_bd_ram_mem2_reg[236][17]/P0001 , \wishbone_bd_ram_mem2_reg[236][18]/P0001 , \wishbone_bd_ram_mem2_reg[236][19]/P0001 , \wishbone_bd_ram_mem2_reg[236][20]/P0001 , \wishbone_bd_ram_mem2_reg[236][21]/P0001 , \wishbone_bd_ram_mem2_reg[236][22]/P0001 , \wishbone_bd_ram_mem2_reg[236][23]/P0001 , \wishbone_bd_ram_mem2_reg[237][16]/P0001 , \wishbone_bd_ram_mem2_reg[237][17]/P0001 , \wishbone_bd_ram_mem2_reg[237][18]/P0001 , \wishbone_bd_ram_mem2_reg[237][19]/P0001 , \wishbone_bd_ram_mem2_reg[237][20]/P0001 , \wishbone_bd_ram_mem2_reg[237][21]/P0001 , \wishbone_bd_ram_mem2_reg[237][22]/P0001 , \wishbone_bd_ram_mem2_reg[237][23]/P0001 , \wishbone_bd_ram_mem2_reg[238][16]/P0001 , \wishbone_bd_ram_mem2_reg[238][17]/P0001 , \wishbone_bd_ram_mem2_reg[238][18]/P0001 , \wishbone_bd_ram_mem2_reg[238][19]/P0001 , \wishbone_bd_ram_mem2_reg[238][20]/P0001 , \wishbone_bd_ram_mem2_reg[238][21]/P0001 , \wishbone_bd_ram_mem2_reg[238][22]/P0001 , \wishbone_bd_ram_mem2_reg[238][23]/P0001 , \wishbone_bd_ram_mem2_reg[239][16]/P0001 , \wishbone_bd_ram_mem2_reg[239][17]/P0001 , \wishbone_bd_ram_mem2_reg[239][18]/P0001 , \wishbone_bd_ram_mem2_reg[239][19]/P0001 , \wishbone_bd_ram_mem2_reg[239][20]/P0001 , \wishbone_bd_ram_mem2_reg[239][21]/P0001 , \wishbone_bd_ram_mem2_reg[239][22]/P0001 , \wishbone_bd_ram_mem2_reg[239][23]/P0001 , \wishbone_bd_ram_mem2_reg[23][16]/P0001 , \wishbone_bd_ram_mem2_reg[23][17]/P0001 , \wishbone_bd_ram_mem2_reg[23][18]/P0001 , \wishbone_bd_ram_mem2_reg[23][19]/P0001 , \wishbone_bd_ram_mem2_reg[23][20]/P0001 , \wishbone_bd_ram_mem2_reg[23][21]/P0001 , \wishbone_bd_ram_mem2_reg[23][22]/P0001 , \wishbone_bd_ram_mem2_reg[23][23]/P0001 , \wishbone_bd_ram_mem2_reg[240][16]/P0001 , \wishbone_bd_ram_mem2_reg[240][17]/P0001 , \wishbone_bd_ram_mem2_reg[240][18]/P0001 , \wishbone_bd_ram_mem2_reg[240][19]/P0001 , \wishbone_bd_ram_mem2_reg[240][20]/P0001 , \wishbone_bd_ram_mem2_reg[240][21]/P0001 , \wishbone_bd_ram_mem2_reg[240][22]/P0001 , \wishbone_bd_ram_mem2_reg[240][23]/P0001 , \wishbone_bd_ram_mem2_reg[241][16]/P0001 , \wishbone_bd_ram_mem2_reg[241][17]/P0001 , \wishbone_bd_ram_mem2_reg[241][18]/P0001 , \wishbone_bd_ram_mem2_reg[241][19]/P0001 , \wishbone_bd_ram_mem2_reg[241][20]/P0001 , \wishbone_bd_ram_mem2_reg[241][21]/P0001 , \wishbone_bd_ram_mem2_reg[241][22]/P0001 , \wishbone_bd_ram_mem2_reg[241][23]/P0001 , \wishbone_bd_ram_mem2_reg[242][16]/P0001 , \wishbone_bd_ram_mem2_reg[242][17]/P0001 , \wishbone_bd_ram_mem2_reg[242][18]/P0001 , \wishbone_bd_ram_mem2_reg[242][19]/P0001 , \wishbone_bd_ram_mem2_reg[242][20]/P0001 , \wishbone_bd_ram_mem2_reg[242][21]/P0001 , \wishbone_bd_ram_mem2_reg[242][22]/P0001 , \wishbone_bd_ram_mem2_reg[242][23]/P0001 , \wishbone_bd_ram_mem2_reg[243][16]/P0001 , \wishbone_bd_ram_mem2_reg[243][17]/P0001 , \wishbone_bd_ram_mem2_reg[243][18]/P0001 , \wishbone_bd_ram_mem2_reg[243][19]/P0001 , \wishbone_bd_ram_mem2_reg[243][20]/P0001 , \wishbone_bd_ram_mem2_reg[243][21]/P0001 , \wishbone_bd_ram_mem2_reg[243][22]/P0001 , \wishbone_bd_ram_mem2_reg[243][23]/P0001 , \wishbone_bd_ram_mem2_reg[244][16]/P0001 , \wishbone_bd_ram_mem2_reg[244][17]/P0001 , \wishbone_bd_ram_mem2_reg[244][18]/P0001 , \wishbone_bd_ram_mem2_reg[244][19]/P0001 , \wishbone_bd_ram_mem2_reg[244][20]/P0001 , \wishbone_bd_ram_mem2_reg[244][21]/P0001 , \wishbone_bd_ram_mem2_reg[244][22]/P0001 , \wishbone_bd_ram_mem2_reg[244][23]/P0001 , \wishbone_bd_ram_mem2_reg[245][16]/P0001 , \wishbone_bd_ram_mem2_reg[245][17]/P0001 , \wishbone_bd_ram_mem2_reg[245][18]/P0001 , \wishbone_bd_ram_mem2_reg[245][19]/P0001 , \wishbone_bd_ram_mem2_reg[245][20]/P0001 , \wishbone_bd_ram_mem2_reg[245][21]/P0001 , \wishbone_bd_ram_mem2_reg[245][22]/P0001 , \wishbone_bd_ram_mem2_reg[245][23]/P0001 , \wishbone_bd_ram_mem2_reg[246][16]/P0001 , \wishbone_bd_ram_mem2_reg[246][17]/P0001 , \wishbone_bd_ram_mem2_reg[246][18]/P0001 , \wishbone_bd_ram_mem2_reg[246][19]/P0001 , \wishbone_bd_ram_mem2_reg[246][20]/P0001 , \wishbone_bd_ram_mem2_reg[246][21]/P0001 , \wishbone_bd_ram_mem2_reg[246][22]/P0001 , \wishbone_bd_ram_mem2_reg[246][23]/P0001 , \wishbone_bd_ram_mem2_reg[247][16]/P0001 , \wishbone_bd_ram_mem2_reg[247][17]/P0001 , \wishbone_bd_ram_mem2_reg[247][18]/P0001 , \wishbone_bd_ram_mem2_reg[247][19]/P0001 , \wishbone_bd_ram_mem2_reg[247][20]/P0001 , \wishbone_bd_ram_mem2_reg[247][21]/P0001 , \wishbone_bd_ram_mem2_reg[247][22]/P0001 , \wishbone_bd_ram_mem2_reg[247][23]/P0001 , \wishbone_bd_ram_mem2_reg[248][16]/P0001 , \wishbone_bd_ram_mem2_reg[248][17]/P0001 , \wishbone_bd_ram_mem2_reg[248][18]/P0001 , \wishbone_bd_ram_mem2_reg[248][19]/P0001 , \wishbone_bd_ram_mem2_reg[248][20]/P0001 , \wishbone_bd_ram_mem2_reg[248][21]/P0001 , \wishbone_bd_ram_mem2_reg[248][22]/P0001 , \wishbone_bd_ram_mem2_reg[248][23]/P0001 , \wishbone_bd_ram_mem2_reg[249][16]/P0001 , \wishbone_bd_ram_mem2_reg[249][17]/P0001 , \wishbone_bd_ram_mem2_reg[249][18]/P0001 , \wishbone_bd_ram_mem2_reg[249][19]/P0001 , \wishbone_bd_ram_mem2_reg[249][20]/P0001 , \wishbone_bd_ram_mem2_reg[249][21]/P0001 , \wishbone_bd_ram_mem2_reg[249][22]/P0001 , \wishbone_bd_ram_mem2_reg[249][23]/P0001 , \wishbone_bd_ram_mem2_reg[24][16]/P0001 , \wishbone_bd_ram_mem2_reg[24][17]/P0001 , \wishbone_bd_ram_mem2_reg[24][18]/P0001 , \wishbone_bd_ram_mem2_reg[24][19]/P0001 , \wishbone_bd_ram_mem2_reg[24][20]/P0001 , \wishbone_bd_ram_mem2_reg[24][21]/P0001 , \wishbone_bd_ram_mem2_reg[24][22]/P0001 , \wishbone_bd_ram_mem2_reg[24][23]/P0001 , \wishbone_bd_ram_mem2_reg[250][16]/P0001 , \wishbone_bd_ram_mem2_reg[250][17]/P0001 , \wishbone_bd_ram_mem2_reg[250][18]/P0001 , \wishbone_bd_ram_mem2_reg[250][19]/P0001 , \wishbone_bd_ram_mem2_reg[250][20]/P0001 , \wishbone_bd_ram_mem2_reg[250][21]/P0001 , \wishbone_bd_ram_mem2_reg[250][22]/P0001 , \wishbone_bd_ram_mem2_reg[250][23]/P0001 , \wishbone_bd_ram_mem2_reg[251][16]/P0001 , \wishbone_bd_ram_mem2_reg[251][17]/P0001 , \wishbone_bd_ram_mem2_reg[251][18]/P0001 , \wishbone_bd_ram_mem2_reg[251][19]/P0001 , \wishbone_bd_ram_mem2_reg[251][20]/P0001 , \wishbone_bd_ram_mem2_reg[251][21]/P0001 , \wishbone_bd_ram_mem2_reg[251][22]/P0001 , \wishbone_bd_ram_mem2_reg[251][23]/P0001 , \wishbone_bd_ram_mem2_reg[252][16]/P0001 , \wishbone_bd_ram_mem2_reg[252][17]/P0001 , \wishbone_bd_ram_mem2_reg[252][18]/P0001 , \wishbone_bd_ram_mem2_reg[252][19]/P0001 , \wishbone_bd_ram_mem2_reg[252][20]/P0001 , \wishbone_bd_ram_mem2_reg[252][21]/P0001 , \wishbone_bd_ram_mem2_reg[252][22]/P0001 , \wishbone_bd_ram_mem2_reg[252][23]/P0001 , \wishbone_bd_ram_mem2_reg[253][16]/P0001 , \wishbone_bd_ram_mem2_reg[253][17]/P0001 , \wishbone_bd_ram_mem2_reg[253][18]/P0001 , \wishbone_bd_ram_mem2_reg[253][19]/P0001 , \wishbone_bd_ram_mem2_reg[253][20]/P0001 , \wishbone_bd_ram_mem2_reg[253][21]/P0001 , \wishbone_bd_ram_mem2_reg[253][22]/P0001 , \wishbone_bd_ram_mem2_reg[253][23]/P0001 , \wishbone_bd_ram_mem2_reg[254][16]/P0001 , \wishbone_bd_ram_mem2_reg[254][17]/P0001 , \wishbone_bd_ram_mem2_reg[254][18]/P0001 , \wishbone_bd_ram_mem2_reg[254][19]/P0001 , \wishbone_bd_ram_mem2_reg[254][20]/P0001 , \wishbone_bd_ram_mem2_reg[254][21]/P0001 , \wishbone_bd_ram_mem2_reg[254][22]/P0001 , \wishbone_bd_ram_mem2_reg[254][23]/P0001 , \wishbone_bd_ram_mem2_reg[255][16]/P0001 , \wishbone_bd_ram_mem2_reg[255][17]/P0001 , \wishbone_bd_ram_mem2_reg[255][18]/P0001 , \wishbone_bd_ram_mem2_reg[255][19]/P0001 , \wishbone_bd_ram_mem2_reg[255][20]/P0001 , \wishbone_bd_ram_mem2_reg[255][21]/P0001 , \wishbone_bd_ram_mem2_reg[255][22]/P0001 , \wishbone_bd_ram_mem2_reg[255][23]/P0001 , \wishbone_bd_ram_mem2_reg[25][16]/P0001 , \wishbone_bd_ram_mem2_reg[25][17]/P0001 , \wishbone_bd_ram_mem2_reg[25][18]/P0001 , \wishbone_bd_ram_mem2_reg[25][19]/P0001 , \wishbone_bd_ram_mem2_reg[25][20]/P0001 , \wishbone_bd_ram_mem2_reg[25][21]/P0001 , \wishbone_bd_ram_mem2_reg[25][22]/P0001 , \wishbone_bd_ram_mem2_reg[25][23]/P0001 , \wishbone_bd_ram_mem2_reg[26][16]/P0001 , \wishbone_bd_ram_mem2_reg[26][17]/P0001 , \wishbone_bd_ram_mem2_reg[26][18]/P0001 , \wishbone_bd_ram_mem2_reg[26][19]/P0001 , \wishbone_bd_ram_mem2_reg[26][20]/P0001 , \wishbone_bd_ram_mem2_reg[26][21]/P0001 , \wishbone_bd_ram_mem2_reg[26][22]/P0001 , \wishbone_bd_ram_mem2_reg[26][23]/P0001 , \wishbone_bd_ram_mem2_reg[27][16]/P0001 , \wishbone_bd_ram_mem2_reg[27][17]/P0001 , \wishbone_bd_ram_mem2_reg[27][18]/P0001 , \wishbone_bd_ram_mem2_reg[27][19]/P0001 , \wishbone_bd_ram_mem2_reg[27][20]/P0001 , \wishbone_bd_ram_mem2_reg[27][21]/P0001 , \wishbone_bd_ram_mem2_reg[27][22]/P0001 , \wishbone_bd_ram_mem2_reg[27][23]/P0001 , \wishbone_bd_ram_mem2_reg[28][16]/P0001 , \wishbone_bd_ram_mem2_reg[28][17]/P0001 , \wishbone_bd_ram_mem2_reg[28][18]/P0001 , \wishbone_bd_ram_mem2_reg[28][19]/P0001 , \wishbone_bd_ram_mem2_reg[28][20]/P0001 , \wishbone_bd_ram_mem2_reg[28][21]/P0001 , \wishbone_bd_ram_mem2_reg[28][22]/P0001 , \wishbone_bd_ram_mem2_reg[28][23]/P0001 , \wishbone_bd_ram_mem2_reg[29][16]/P0001 , \wishbone_bd_ram_mem2_reg[29][17]/P0001 , \wishbone_bd_ram_mem2_reg[29][18]/P0001 , \wishbone_bd_ram_mem2_reg[29][19]/P0001 , \wishbone_bd_ram_mem2_reg[29][20]/P0001 , \wishbone_bd_ram_mem2_reg[29][21]/P0001 , \wishbone_bd_ram_mem2_reg[29][22]/P0001 , \wishbone_bd_ram_mem2_reg[29][23]/P0001 , \wishbone_bd_ram_mem2_reg[2][16]/P0001 , \wishbone_bd_ram_mem2_reg[2][17]/P0001 , \wishbone_bd_ram_mem2_reg[2][18]/P0001 , \wishbone_bd_ram_mem2_reg[2][19]/P0001 , \wishbone_bd_ram_mem2_reg[2][20]/P0001 , \wishbone_bd_ram_mem2_reg[2][21]/P0001 , \wishbone_bd_ram_mem2_reg[2][22]/P0001 , \wishbone_bd_ram_mem2_reg[2][23]/P0001 , \wishbone_bd_ram_mem2_reg[30][16]/P0001 , \wishbone_bd_ram_mem2_reg[30][17]/P0001 , \wishbone_bd_ram_mem2_reg[30][18]/P0001 , \wishbone_bd_ram_mem2_reg[30][19]/P0001 , \wishbone_bd_ram_mem2_reg[30][20]/P0001 , \wishbone_bd_ram_mem2_reg[30][21]/P0001 , \wishbone_bd_ram_mem2_reg[30][22]/P0001 , \wishbone_bd_ram_mem2_reg[30][23]/P0001 , \wishbone_bd_ram_mem2_reg[31][16]/P0001 , \wishbone_bd_ram_mem2_reg[31][17]/P0001 , \wishbone_bd_ram_mem2_reg[31][18]/P0001 , \wishbone_bd_ram_mem2_reg[31][19]/P0001 , \wishbone_bd_ram_mem2_reg[31][20]/P0001 , \wishbone_bd_ram_mem2_reg[31][21]/P0001 , \wishbone_bd_ram_mem2_reg[31][22]/P0001 , \wishbone_bd_ram_mem2_reg[31][23]/P0001 , \wishbone_bd_ram_mem2_reg[32][16]/P0001 , \wishbone_bd_ram_mem2_reg[32][17]/P0001 , \wishbone_bd_ram_mem2_reg[32][18]/P0001 , \wishbone_bd_ram_mem2_reg[32][19]/P0001 , \wishbone_bd_ram_mem2_reg[32][20]/P0001 , \wishbone_bd_ram_mem2_reg[32][21]/P0001 , \wishbone_bd_ram_mem2_reg[32][22]/P0001 , \wishbone_bd_ram_mem2_reg[32][23]/P0001 , \wishbone_bd_ram_mem2_reg[33][16]/P0001 , \wishbone_bd_ram_mem2_reg[33][17]/P0001 , \wishbone_bd_ram_mem2_reg[33][18]/P0001 , \wishbone_bd_ram_mem2_reg[33][19]/P0001 , \wishbone_bd_ram_mem2_reg[33][20]/P0001 , \wishbone_bd_ram_mem2_reg[33][21]/P0001 , \wishbone_bd_ram_mem2_reg[33][22]/P0001 , \wishbone_bd_ram_mem2_reg[33][23]/P0001 , \wishbone_bd_ram_mem2_reg[34][16]/P0001 , \wishbone_bd_ram_mem2_reg[34][17]/P0001 , \wishbone_bd_ram_mem2_reg[34][18]/P0001 , \wishbone_bd_ram_mem2_reg[34][19]/P0001 , \wishbone_bd_ram_mem2_reg[34][20]/P0001 , \wishbone_bd_ram_mem2_reg[34][21]/P0001 , \wishbone_bd_ram_mem2_reg[34][22]/P0001 , \wishbone_bd_ram_mem2_reg[34][23]/P0001 , \wishbone_bd_ram_mem2_reg[35][16]/P0001 , \wishbone_bd_ram_mem2_reg[35][17]/P0001 , \wishbone_bd_ram_mem2_reg[35][18]/P0001 , \wishbone_bd_ram_mem2_reg[35][19]/P0001 , \wishbone_bd_ram_mem2_reg[35][20]/P0001 , \wishbone_bd_ram_mem2_reg[35][21]/P0001 , \wishbone_bd_ram_mem2_reg[35][22]/P0001 , \wishbone_bd_ram_mem2_reg[35][23]/P0001 , \wishbone_bd_ram_mem2_reg[36][16]/P0001 , \wishbone_bd_ram_mem2_reg[36][17]/P0001 , \wishbone_bd_ram_mem2_reg[36][18]/P0001 , \wishbone_bd_ram_mem2_reg[36][19]/P0001 , \wishbone_bd_ram_mem2_reg[36][20]/P0001 , \wishbone_bd_ram_mem2_reg[36][21]/P0001 , \wishbone_bd_ram_mem2_reg[36][22]/P0001 , \wishbone_bd_ram_mem2_reg[36][23]/P0001 , \wishbone_bd_ram_mem2_reg[37][16]/P0001 , \wishbone_bd_ram_mem2_reg[37][17]/P0001 , \wishbone_bd_ram_mem2_reg[37][18]/P0001 , \wishbone_bd_ram_mem2_reg[37][19]/P0001 , \wishbone_bd_ram_mem2_reg[37][20]/P0001 , \wishbone_bd_ram_mem2_reg[37][21]/P0001 , \wishbone_bd_ram_mem2_reg[37][22]/P0001 , \wishbone_bd_ram_mem2_reg[37][23]/P0001 , \wishbone_bd_ram_mem2_reg[38][16]/P0001 , \wishbone_bd_ram_mem2_reg[38][17]/P0001 , \wishbone_bd_ram_mem2_reg[38][18]/P0001 , \wishbone_bd_ram_mem2_reg[38][19]/P0001 , \wishbone_bd_ram_mem2_reg[38][20]/P0001 , \wishbone_bd_ram_mem2_reg[38][21]/P0001 , \wishbone_bd_ram_mem2_reg[38][22]/P0001 , \wishbone_bd_ram_mem2_reg[38][23]/P0001 , \wishbone_bd_ram_mem2_reg[39][16]/P0001 , \wishbone_bd_ram_mem2_reg[39][17]/P0001 , \wishbone_bd_ram_mem2_reg[39][18]/P0001 , \wishbone_bd_ram_mem2_reg[39][19]/P0001 , \wishbone_bd_ram_mem2_reg[39][20]/P0001 , \wishbone_bd_ram_mem2_reg[39][21]/P0001 , \wishbone_bd_ram_mem2_reg[39][22]/P0001 , \wishbone_bd_ram_mem2_reg[39][23]/P0001 , \wishbone_bd_ram_mem2_reg[3][16]/P0001 , \wishbone_bd_ram_mem2_reg[3][17]/P0001 , \wishbone_bd_ram_mem2_reg[3][18]/P0001 , \wishbone_bd_ram_mem2_reg[3][19]/P0001 , \wishbone_bd_ram_mem2_reg[3][20]/P0001 , \wishbone_bd_ram_mem2_reg[3][21]/P0001 , \wishbone_bd_ram_mem2_reg[3][22]/P0001 , \wishbone_bd_ram_mem2_reg[3][23]/P0001 , \wishbone_bd_ram_mem2_reg[40][16]/P0001 , \wishbone_bd_ram_mem2_reg[40][17]/P0001 , \wishbone_bd_ram_mem2_reg[40][18]/P0001 , \wishbone_bd_ram_mem2_reg[40][19]/P0001 , \wishbone_bd_ram_mem2_reg[40][20]/P0001 , \wishbone_bd_ram_mem2_reg[40][21]/P0001 , \wishbone_bd_ram_mem2_reg[40][22]/P0001 , \wishbone_bd_ram_mem2_reg[40][23]/P0001 , \wishbone_bd_ram_mem2_reg[41][16]/P0001 , \wishbone_bd_ram_mem2_reg[41][17]/P0001 , \wishbone_bd_ram_mem2_reg[41][18]/P0001 , \wishbone_bd_ram_mem2_reg[41][19]/P0001 , \wishbone_bd_ram_mem2_reg[41][20]/P0001 , \wishbone_bd_ram_mem2_reg[41][21]/P0001 , \wishbone_bd_ram_mem2_reg[41][22]/P0001 , \wishbone_bd_ram_mem2_reg[41][23]/P0001 , \wishbone_bd_ram_mem2_reg[42][16]/P0001 , \wishbone_bd_ram_mem2_reg[42][17]/P0001 , \wishbone_bd_ram_mem2_reg[42][18]/P0001 , \wishbone_bd_ram_mem2_reg[42][19]/P0001 , \wishbone_bd_ram_mem2_reg[42][20]/P0001 , \wishbone_bd_ram_mem2_reg[42][21]/P0001 , \wishbone_bd_ram_mem2_reg[42][22]/P0001 , \wishbone_bd_ram_mem2_reg[42][23]/P0001 , \wishbone_bd_ram_mem2_reg[43][16]/P0001 , \wishbone_bd_ram_mem2_reg[43][17]/P0001 , \wishbone_bd_ram_mem2_reg[43][18]/P0001 , \wishbone_bd_ram_mem2_reg[43][19]/P0001 , \wishbone_bd_ram_mem2_reg[43][20]/P0001 , \wishbone_bd_ram_mem2_reg[43][21]/P0001 , \wishbone_bd_ram_mem2_reg[43][22]/P0001 , \wishbone_bd_ram_mem2_reg[43][23]/P0001 , \wishbone_bd_ram_mem2_reg[44][16]/P0001 , \wishbone_bd_ram_mem2_reg[44][17]/P0001 , \wishbone_bd_ram_mem2_reg[44][18]/P0001 , \wishbone_bd_ram_mem2_reg[44][19]/P0001 , \wishbone_bd_ram_mem2_reg[44][20]/P0001 , \wishbone_bd_ram_mem2_reg[44][21]/P0001 , \wishbone_bd_ram_mem2_reg[44][22]/P0001 , \wishbone_bd_ram_mem2_reg[44][23]/P0001 , \wishbone_bd_ram_mem2_reg[45][16]/P0001 , \wishbone_bd_ram_mem2_reg[45][17]/P0001 , \wishbone_bd_ram_mem2_reg[45][18]/P0001 , \wishbone_bd_ram_mem2_reg[45][19]/P0001 , \wishbone_bd_ram_mem2_reg[45][20]/P0001 , \wishbone_bd_ram_mem2_reg[45][21]/P0001 , \wishbone_bd_ram_mem2_reg[45][22]/P0001 , \wishbone_bd_ram_mem2_reg[45][23]/P0001 , \wishbone_bd_ram_mem2_reg[46][16]/P0001 , \wishbone_bd_ram_mem2_reg[46][17]/P0001 , \wishbone_bd_ram_mem2_reg[46][18]/P0001 , \wishbone_bd_ram_mem2_reg[46][19]/P0001 , \wishbone_bd_ram_mem2_reg[46][20]/P0001 , \wishbone_bd_ram_mem2_reg[46][21]/P0001 , \wishbone_bd_ram_mem2_reg[46][22]/P0001 , \wishbone_bd_ram_mem2_reg[46][23]/P0001 , \wishbone_bd_ram_mem2_reg[47][16]/P0001 , \wishbone_bd_ram_mem2_reg[47][17]/P0001 , \wishbone_bd_ram_mem2_reg[47][18]/P0001 , \wishbone_bd_ram_mem2_reg[47][19]/P0001 , \wishbone_bd_ram_mem2_reg[47][20]/P0001 , \wishbone_bd_ram_mem2_reg[47][21]/P0001 , \wishbone_bd_ram_mem2_reg[47][22]/P0001 , \wishbone_bd_ram_mem2_reg[47][23]/P0001 , \wishbone_bd_ram_mem2_reg[48][16]/P0001 , \wishbone_bd_ram_mem2_reg[48][17]/P0001 , \wishbone_bd_ram_mem2_reg[48][18]/P0001 , \wishbone_bd_ram_mem2_reg[48][19]/P0001 , \wishbone_bd_ram_mem2_reg[48][20]/P0001 , \wishbone_bd_ram_mem2_reg[48][21]/P0001 , \wishbone_bd_ram_mem2_reg[48][22]/P0001 , \wishbone_bd_ram_mem2_reg[48][23]/P0001 , \wishbone_bd_ram_mem2_reg[49][16]/P0001 , \wishbone_bd_ram_mem2_reg[49][17]/P0001 , \wishbone_bd_ram_mem2_reg[49][18]/P0001 , \wishbone_bd_ram_mem2_reg[49][19]/P0001 , \wishbone_bd_ram_mem2_reg[49][20]/P0001 , \wishbone_bd_ram_mem2_reg[49][21]/P0001 , \wishbone_bd_ram_mem2_reg[49][22]/P0001 , \wishbone_bd_ram_mem2_reg[49][23]/P0001 , \wishbone_bd_ram_mem2_reg[4][16]/P0001 , \wishbone_bd_ram_mem2_reg[4][17]/P0001 , \wishbone_bd_ram_mem2_reg[4][18]/P0001 , \wishbone_bd_ram_mem2_reg[4][19]/P0001 , \wishbone_bd_ram_mem2_reg[4][20]/P0001 , \wishbone_bd_ram_mem2_reg[4][21]/P0001 , \wishbone_bd_ram_mem2_reg[4][22]/P0001 , \wishbone_bd_ram_mem2_reg[4][23]/P0001 , \wishbone_bd_ram_mem2_reg[50][16]/P0001 , \wishbone_bd_ram_mem2_reg[50][17]/P0001 , \wishbone_bd_ram_mem2_reg[50][18]/P0001 , \wishbone_bd_ram_mem2_reg[50][19]/P0001 , \wishbone_bd_ram_mem2_reg[50][20]/P0001 , \wishbone_bd_ram_mem2_reg[50][21]/P0001 , \wishbone_bd_ram_mem2_reg[50][22]/P0001 , \wishbone_bd_ram_mem2_reg[50][23]/P0001 , \wishbone_bd_ram_mem2_reg[51][16]/P0001 , \wishbone_bd_ram_mem2_reg[51][17]/P0001 , \wishbone_bd_ram_mem2_reg[51][18]/P0001 , \wishbone_bd_ram_mem2_reg[51][19]/P0001 , \wishbone_bd_ram_mem2_reg[51][20]/P0001 , \wishbone_bd_ram_mem2_reg[51][21]/P0001 , \wishbone_bd_ram_mem2_reg[51][22]/P0001 , \wishbone_bd_ram_mem2_reg[51][23]/P0001 , \wishbone_bd_ram_mem2_reg[52][16]/P0001 , \wishbone_bd_ram_mem2_reg[52][17]/P0001 , \wishbone_bd_ram_mem2_reg[52][18]/P0001 , \wishbone_bd_ram_mem2_reg[52][19]/P0001 , \wishbone_bd_ram_mem2_reg[52][20]/P0001 , \wishbone_bd_ram_mem2_reg[52][21]/P0001 , \wishbone_bd_ram_mem2_reg[52][22]/P0001 , \wishbone_bd_ram_mem2_reg[52][23]/P0001 , \wishbone_bd_ram_mem2_reg[53][16]/P0001 , \wishbone_bd_ram_mem2_reg[53][17]/P0001 , \wishbone_bd_ram_mem2_reg[53][18]/P0001 , \wishbone_bd_ram_mem2_reg[53][19]/P0001 , \wishbone_bd_ram_mem2_reg[53][20]/P0001 , \wishbone_bd_ram_mem2_reg[53][21]/P0001 , \wishbone_bd_ram_mem2_reg[53][22]/P0001 , \wishbone_bd_ram_mem2_reg[53][23]/P0001 , \wishbone_bd_ram_mem2_reg[54][16]/P0001 , \wishbone_bd_ram_mem2_reg[54][17]/P0001 , \wishbone_bd_ram_mem2_reg[54][18]/P0001 , \wishbone_bd_ram_mem2_reg[54][19]/P0001 , \wishbone_bd_ram_mem2_reg[54][20]/P0001 , \wishbone_bd_ram_mem2_reg[54][21]/P0001 , \wishbone_bd_ram_mem2_reg[54][22]/P0001 , \wishbone_bd_ram_mem2_reg[54][23]/P0001 , \wishbone_bd_ram_mem2_reg[55][16]/P0001 , \wishbone_bd_ram_mem2_reg[55][17]/P0001 , \wishbone_bd_ram_mem2_reg[55][18]/P0001 , \wishbone_bd_ram_mem2_reg[55][19]/P0001 , \wishbone_bd_ram_mem2_reg[55][20]/P0001 , \wishbone_bd_ram_mem2_reg[55][21]/P0001 , \wishbone_bd_ram_mem2_reg[55][22]/P0001 , \wishbone_bd_ram_mem2_reg[55][23]/P0001 , \wishbone_bd_ram_mem2_reg[56][16]/P0001 , \wishbone_bd_ram_mem2_reg[56][17]/P0001 , \wishbone_bd_ram_mem2_reg[56][18]/P0001 , \wishbone_bd_ram_mem2_reg[56][19]/P0001 , \wishbone_bd_ram_mem2_reg[56][20]/P0001 , \wishbone_bd_ram_mem2_reg[56][21]/P0001 , \wishbone_bd_ram_mem2_reg[56][22]/P0001 , \wishbone_bd_ram_mem2_reg[56][23]/P0001 , \wishbone_bd_ram_mem2_reg[57][16]/P0001 , \wishbone_bd_ram_mem2_reg[57][17]/P0001 , \wishbone_bd_ram_mem2_reg[57][18]/P0001 , \wishbone_bd_ram_mem2_reg[57][19]/P0001 , \wishbone_bd_ram_mem2_reg[57][20]/P0001 , \wishbone_bd_ram_mem2_reg[57][21]/P0001 , \wishbone_bd_ram_mem2_reg[57][22]/P0001 , \wishbone_bd_ram_mem2_reg[57][23]/P0001 , \wishbone_bd_ram_mem2_reg[58][16]/P0001 , \wishbone_bd_ram_mem2_reg[58][17]/P0001 , \wishbone_bd_ram_mem2_reg[58][18]/P0001 , \wishbone_bd_ram_mem2_reg[58][19]/P0001 , \wishbone_bd_ram_mem2_reg[58][20]/P0001 , \wishbone_bd_ram_mem2_reg[58][21]/P0001 , \wishbone_bd_ram_mem2_reg[58][22]/P0001 , \wishbone_bd_ram_mem2_reg[58][23]/P0001 , \wishbone_bd_ram_mem2_reg[59][16]/P0001 , \wishbone_bd_ram_mem2_reg[59][17]/P0001 , \wishbone_bd_ram_mem2_reg[59][18]/P0001 , \wishbone_bd_ram_mem2_reg[59][19]/P0001 , \wishbone_bd_ram_mem2_reg[59][20]/P0001 , \wishbone_bd_ram_mem2_reg[59][21]/P0001 , \wishbone_bd_ram_mem2_reg[59][22]/P0001 , \wishbone_bd_ram_mem2_reg[59][23]/P0001 , \wishbone_bd_ram_mem2_reg[5][16]/P0001 , \wishbone_bd_ram_mem2_reg[5][17]/P0001 , \wishbone_bd_ram_mem2_reg[5][18]/P0001 , \wishbone_bd_ram_mem2_reg[5][19]/P0001 , \wishbone_bd_ram_mem2_reg[5][20]/P0001 , \wishbone_bd_ram_mem2_reg[5][21]/P0001 , \wishbone_bd_ram_mem2_reg[5][22]/P0001 , \wishbone_bd_ram_mem2_reg[5][23]/P0001 , \wishbone_bd_ram_mem2_reg[60][16]/P0001 , \wishbone_bd_ram_mem2_reg[60][17]/P0001 , \wishbone_bd_ram_mem2_reg[60][18]/P0001 , \wishbone_bd_ram_mem2_reg[60][19]/P0001 , \wishbone_bd_ram_mem2_reg[60][20]/P0001 , \wishbone_bd_ram_mem2_reg[60][21]/P0001 , \wishbone_bd_ram_mem2_reg[60][22]/P0001 , \wishbone_bd_ram_mem2_reg[60][23]/P0001 , \wishbone_bd_ram_mem2_reg[61][16]/P0001 , \wishbone_bd_ram_mem2_reg[61][17]/P0001 , \wishbone_bd_ram_mem2_reg[61][18]/P0001 , \wishbone_bd_ram_mem2_reg[61][19]/P0001 , \wishbone_bd_ram_mem2_reg[61][20]/P0001 , \wishbone_bd_ram_mem2_reg[61][21]/P0001 , \wishbone_bd_ram_mem2_reg[61][22]/P0001 , \wishbone_bd_ram_mem2_reg[61][23]/P0001 , \wishbone_bd_ram_mem2_reg[62][16]/P0001 , \wishbone_bd_ram_mem2_reg[62][17]/P0001 , \wishbone_bd_ram_mem2_reg[62][18]/P0001 , \wishbone_bd_ram_mem2_reg[62][19]/P0001 , \wishbone_bd_ram_mem2_reg[62][20]/P0001 , \wishbone_bd_ram_mem2_reg[62][21]/P0001 , \wishbone_bd_ram_mem2_reg[62][22]/P0001 , \wishbone_bd_ram_mem2_reg[62][23]/P0001 , \wishbone_bd_ram_mem2_reg[63][16]/P0001 , \wishbone_bd_ram_mem2_reg[63][17]/P0001 , \wishbone_bd_ram_mem2_reg[63][18]/P0001 , \wishbone_bd_ram_mem2_reg[63][19]/P0001 , \wishbone_bd_ram_mem2_reg[63][20]/P0001 , \wishbone_bd_ram_mem2_reg[63][21]/P0001 , \wishbone_bd_ram_mem2_reg[63][22]/P0001 , \wishbone_bd_ram_mem2_reg[63][23]/P0001 , \wishbone_bd_ram_mem2_reg[64][16]/P0001 , \wishbone_bd_ram_mem2_reg[64][17]/P0001 , \wishbone_bd_ram_mem2_reg[64][18]/P0001 , \wishbone_bd_ram_mem2_reg[64][19]/P0001 , \wishbone_bd_ram_mem2_reg[64][20]/P0001 , \wishbone_bd_ram_mem2_reg[64][21]/P0001 , \wishbone_bd_ram_mem2_reg[64][22]/P0001 , \wishbone_bd_ram_mem2_reg[64][23]/P0001 , \wishbone_bd_ram_mem2_reg[65][16]/P0001 , \wishbone_bd_ram_mem2_reg[65][17]/P0001 , \wishbone_bd_ram_mem2_reg[65][18]/P0001 , \wishbone_bd_ram_mem2_reg[65][19]/P0001 , \wishbone_bd_ram_mem2_reg[65][20]/P0001 , \wishbone_bd_ram_mem2_reg[65][21]/P0001 , \wishbone_bd_ram_mem2_reg[65][22]/P0001 , \wishbone_bd_ram_mem2_reg[65][23]/P0001 , \wishbone_bd_ram_mem2_reg[66][16]/P0001 , \wishbone_bd_ram_mem2_reg[66][17]/P0001 , \wishbone_bd_ram_mem2_reg[66][18]/P0001 , \wishbone_bd_ram_mem2_reg[66][19]/P0001 , \wishbone_bd_ram_mem2_reg[66][20]/P0001 , \wishbone_bd_ram_mem2_reg[66][21]/P0001 , \wishbone_bd_ram_mem2_reg[66][22]/P0001 , \wishbone_bd_ram_mem2_reg[66][23]/P0001 , \wishbone_bd_ram_mem2_reg[67][16]/P0001 , \wishbone_bd_ram_mem2_reg[67][17]/P0001 , \wishbone_bd_ram_mem2_reg[67][18]/P0001 , \wishbone_bd_ram_mem2_reg[67][19]/P0001 , \wishbone_bd_ram_mem2_reg[67][20]/P0001 , \wishbone_bd_ram_mem2_reg[67][21]/P0001 , \wishbone_bd_ram_mem2_reg[67][22]/P0001 , \wishbone_bd_ram_mem2_reg[67][23]/P0001 , \wishbone_bd_ram_mem2_reg[68][16]/P0001 , \wishbone_bd_ram_mem2_reg[68][17]/P0001 , \wishbone_bd_ram_mem2_reg[68][18]/P0001 , \wishbone_bd_ram_mem2_reg[68][19]/P0001 , \wishbone_bd_ram_mem2_reg[68][20]/P0001 , \wishbone_bd_ram_mem2_reg[68][21]/P0001 , \wishbone_bd_ram_mem2_reg[68][22]/P0001 , \wishbone_bd_ram_mem2_reg[68][23]/P0001 , \wishbone_bd_ram_mem2_reg[69][16]/P0001 , \wishbone_bd_ram_mem2_reg[69][17]/P0001 , \wishbone_bd_ram_mem2_reg[69][18]/P0001 , \wishbone_bd_ram_mem2_reg[69][19]/P0001 , \wishbone_bd_ram_mem2_reg[69][20]/P0001 , \wishbone_bd_ram_mem2_reg[69][21]/P0001 , \wishbone_bd_ram_mem2_reg[69][22]/P0001 , \wishbone_bd_ram_mem2_reg[69][23]/P0001 , \wishbone_bd_ram_mem2_reg[6][16]/P0001 , \wishbone_bd_ram_mem2_reg[6][17]/P0001 , \wishbone_bd_ram_mem2_reg[6][18]/P0001 , \wishbone_bd_ram_mem2_reg[6][19]/P0001 , \wishbone_bd_ram_mem2_reg[6][20]/P0001 , \wishbone_bd_ram_mem2_reg[6][21]/P0001 , \wishbone_bd_ram_mem2_reg[6][22]/P0001 , \wishbone_bd_ram_mem2_reg[6][23]/P0001 , \wishbone_bd_ram_mem2_reg[70][16]/P0001 , \wishbone_bd_ram_mem2_reg[70][17]/P0001 , \wishbone_bd_ram_mem2_reg[70][18]/P0001 , \wishbone_bd_ram_mem2_reg[70][19]/P0001 , \wishbone_bd_ram_mem2_reg[70][20]/P0001 , \wishbone_bd_ram_mem2_reg[70][21]/P0001 , \wishbone_bd_ram_mem2_reg[70][22]/P0001 , \wishbone_bd_ram_mem2_reg[70][23]/P0001 , \wishbone_bd_ram_mem2_reg[71][16]/P0001 , \wishbone_bd_ram_mem2_reg[71][17]/P0001 , \wishbone_bd_ram_mem2_reg[71][18]/P0001 , \wishbone_bd_ram_mem2_reg[71][19]/P0001 , \wishbone_bd_ram_mem2_reg[71][20]/P0001 , \wishbone_bd_ram_mem2_reg[71][21]/P0001 , \wishbone_bd_ram_mem2_reg[71][22]/P0001 , \wishbone_bd_ram_mem2_reg[71][23]/P0001 , \wishbone_bd_ram_mem2_reg[72][16]/P0001 , \wishbone_bd_ram_mem2_reg[72][17]/P0001 , \wishbone_bd_ram_mem2_reg[72][18]/P0001 , \wishbone_bd_ram_mem2_reg[72][19]/P0001 , \wishbone_bd_ram_mem2_reg[72][20]/P0001 , \wishbone_bd_ram_mem2_reg[72][21]/P0001 , \wishbone_bd_ram_mem2_reg[72][22]/P0001 , \wishbone_bd_ram_mem2_reg[72][23]/P0001 , \wishbone_bd_ram_mem2_reg[73][16]/P0001 , \wishbone_bd_ram_mem2_reg[73][17]/P0001 , \wishbone_bd_ram_mem2_reg[73][18]/P0001 , \wishbone_bd_ram_mem2_reg[73][19]/P0001 , \wishbone_bd_ram_mem2_reg[73][20]/P0001 , \wishbone_bd_ram_mem2_reg[73][21]/P0001 , \wishbone_bd_ram_mem2_reg[73][22]/P0001 , \wishbone_bd_ram_mem2_reg[73][23]/P0001 , \wishbone_bd_ram_mem2_reg[74][16]/P0001 , \wishbone_bd_ram_mem2_reg[74][17]/P0001 , \wishbone_bd_ram_mem2_reg[74][18]/P0001 , \wishbone_bd_ram_mem2_reg[74][19]/P0001 , \wishbone_bd_ram_mem2_reg[74][20]/P0001 , \wishbone_bd_ram_mem2_reg[74][21]/P0001 , \wishbone_bd_ram_mem2_reg[74][22]/P0001 , \wishbone_bd_ram_mem2_reg[74][23]/P0001 , \wishbone_bd_ram_mem2_reg[75][16]/P0001 , \wishbone_bd_ram_mem2_reg[75][17]/P0001 , \wishbone_bd_ram_mem2_reg[75][18]/P0001 , \wishbone_bd_ram_mem2_reg[75][19]/P0001 , \wishbone_bd_ram_mem2_reg[75][20]/P0001 , \wishbone_bd_ram_mem2_reg[75][21]/P0001 , \wishbone_bd_ram_mem2_reg[75][22]/P0001 , \wishbone_bd_ram_mem2_reg[75][23]/P0001 , \wishbone_bd_ram_mem2_reg[76][16]/P0001 , \wishbone_bd_ram_mem2_reg[76][17]/P0001 , \wishbone_bd_ram_mem2_reg[76][18]/P0001 , \wishbone_bd_ram_mem2_reg[76][19]/P0001 , \wishbone_bd_ram_mem2_reg[76][20]/P0001 , \wishbone_bd_ram_mem2_reg[76][21]/P0001 , \wishbone_bd_ram_mem2_reg[76][22]/P0001 , \wishbone_bd_ram_mem2_reg[76][23]/P0001 , \wishbone_bd_ram_mem2_reg[77][16]/P0001 , \wishbone_bd_ram_mem2_reg[77][17]/P0001 , \wishbone_bd_ram_mem2_reg[77][18]/P0001 , \wishbone_bd_ram_mem2_reg[77][19]/P0001 , \wishbone_bd_ram_mem2_reg[77][20]/P0001 , \wishbone_bd_ram_mem2_reg[77][21]/P0001 , \wishbone_bd_ram_mem2_reg[77][22]/P0001 , \wishbone_bd_ram_mem2_reg[77][23]/P0001 , \wishbone_bd_ram_mem2_reg[78][16]/P0001 , \wishbone_bd_ram_mem2_reg[78][17]/P0001 , \wishbone_bd_ram_mem2_reg[78][18]/P0001 , \wishbone_bd_ram_mem2_reg[78][19]/P0001 , \wishbone_bd_ram_mem2_reg[78][20]/P0001 , \wishbone_bd_ram_mem2_reg[78][21]/P0001 , \wishbone_bd_ram_mem2_reg[78][22]/P0001 , \wishbone_bd_ram_mem2_reg[78][23]/P0001 , \wishbone_bd_ram_mem2_reg[79][16]/P0001 , \wishbone_bd_ram_mem2_reg[79][17]/P0001 , \wishbone_bd_ram_mem2_reg[79][18]/P0001 , \wishbone_bd_ram_mem2_reg[79][19]/P0001 , \wishbone_bd_ram_mem2_reg[79][20]/P0001 , \wishbone_bd_ram_mem2_reg[79][21]/P0001 , \wishbone_bd_ram_mem2_reg[79][22]/P0001 , \wishbone_bd_ram_mem2_reg[79][23]/P0001 , \wishbone_bd_ram_mem2_reg[7][16]/P0001 , \wishbone_bd_ram_mem2_reg[7][17]/P0001 , \wishbone_bd_ram_mem2_reg[7][18]/P0001 , \wishbone_bd_ram_mem2_reg[7][19]/P0001 , \wishbone_bd_ram_mem2_reg[7][20]/P0001 , \wishbone_bd_ram_mem2_reg[7][21]/P0001 , \wishbone_bd_ram_mem2_reg[7][22]/P0001 , \wishbone_bd_ram_mem2_reg[7][23]/P0001 , \wishbone_bd_ram_mem2_reg[80][16]/P0001 , \wishbone_bd_ram_mem2_reg[80][17]/P0001 , \wishbone_bd_ram_mem2_reg[80][18]/P0001 , \wishbone_bd_ram_mem2_reg[80][19]/P0001 , \wishbone_bd_ram_mem2_reg[80][20]/P0001 , \wishbone_bd_ram_mem2_reg[80][21]/P0001 , \wishbone_bd_ram_mem2_reg[80][22]/P0001 , \wishbone_bd_ram_mem2_reg[80][23]/P0001 , \wishbone_bd_ram_mem2_reg[81][16]/P0001 , \wishbone_bd_ram_mem2_reg[81][17]/P0001 , \wishbone_bd_ram_mem2_reg[81][18]/P0001 , \wishbone_bd_ram_mem2_reg[81][19]/P0001 , \wishbone_bd_ram_mem2_reg[81][20]/P0001 , \wishbone_bd_ram_mem2_reg[81][21]/P0001 , \wishbone_bd_ram_mem2_reg[81][22]/P0001 , \wishbone_bd_ram_mem2_reg[81][23]/P0001 , \wishbone_bd_ram_mem2_reg[82][16]/P0001 , \wishbone_bd_ram_mem2_reg[82][17]/P0001 , \wishbone_bd_ram_mem2_reg[82][18]/P0001 , \wishbone_bd_ram_mem2_reg[82][19]/P0001 , \wishbone_bd_ram_mem2_reg[82][20]/P0001 , \wishbone_bd_ram_mem2_reg[82][21]/P0001 , \wishbone_bd_ram_mem2_reg[82][22]/P0001 , \wishbone_bd_ram_mem2_reg[82][23]/P0001 , \wishbone_bd_ram_mem2_reg[83][16]/P0001 , \wishbone_bd_ram_mem2_reg[83][17]/P0001 , \wishbone_bd_ram_mem2_reg[83][18]/P0001 , \wishbone_bd_ram_mem2_reg[83][19]/P0001 , \wishbone_bd_ram_mem2_reg[83][20]/P0001 , \wishbone_bd_ram_mem2_reg[83][21]/P0001 , \wishbone_bd_ram_mem2_reg[83][22]/P0001 , \wishbone_bd_ram_mem2_reg[83][23]/P0001 , \wishbone_bd_ram_mem2_reg[84][16]/P0001 , \wishbone_bd_ram_mem2_reg[84][17]/P0001 , \wishbone_bd_ram_mem2_reg[84][18]/P0001 , \wishbone_bd_ram_mem2_reg[84][19]/P0001 , \wishbone_bd_ram_mem2_reg[84][20]/P0001 , \wishbone_bd_ram_mem2_reg[84][21]/P0001 , \wishbone_bd_ram_mem2_reg[84][22]/P0001 , \wishbone_bd_ram_mem2_reg[84][23]/P0001 , \wishbone_bd_ram_mem2_reg[85][16]/P0001 , \wishbone_bd_ram_mem2_reg[85][17]/P0001 , \wishbone_bd_ram_mem2_reg[85][18]/P0001 , \wishbone_bd_ram_mem2_reg[85][19]/P0001 , \wishbone_bd_ram_mem2_reg[85][20]/P0001 , \wishbone_bd_ram_mem2_reg[85][21]/P0001 , \wishbone_bd_ram_mem2_reg[85][22]/P0001 , \wishbone_bd_ram_mem2_reg[85][23]/P0001 , \wishbone_bd_ram_mem2_reg[86][16]/P0001 , \wishbone_bd_ram_mem2_reg[86][17]/P0001 , \wishbone_bd_ram_mem2_reg[86][18]/P0001 , \wishbone_bd_ram_mem2_reg[86][19]/P0001 , \wishbone_bd_ram_mem2_reg[86][20]/P0001 , \wishbone_bd_ram_mem2_reg[86][21]/P0001 , \wishbone_bd_ram_mem2_reg[86][22]/P0001 , \wishbone_bd_ram_mem2_reg[86][23]/P0001 , \wishbone_bd_ram_mem2_reg[87][16]/P0001 , \wishbone_bd_ram_mem2_reg[87][17]/P0001 , \wishbone_bd_ram_mem2_reg[87][18]/P0001 , \wishbone_bd_ram_mem2_reg[87][19]/P0001 , \wishbone_bd_ram_mem2_reg[87][20]/P0001 , \wishbone_bd_ram_mem2_reg[87][21]/P0001 , \wishbone_bd_ram_mem2_reg[87][22]/P0001 , \wishbone_bd_ram_mem2_reg[87][23]/P0001 , \wishbone_bd_ram_mem2_reg[88][16]/P0001 , \wishbone_bd_ram_mem2_reg[88][17]/P0001 , \wishbone_bd_ram_mem2_reg[88][18]/P0001 , \wishbone_bd_ram_mem2_reg[88][19]/P0001 , \wishbone_bd_ram_mem2_reg[88][20]/P0001 , \wishbone_bd_ram_mem2_reg[88][21]/P0001 , \wishbone_bd_ram_mem2_reg[88][22]/P0001 , \wishbone_bd_ram_mem2_reg[88][23]/P0001 , \wishbone_bd_ram_mem2_reg[89][16]/P0001 , \wishbone_bd_ram_mem2_reg[89][17]/P0001 , \wishbone_bd_ram_mem2_reg[89][18]/P0001 , \wishbone_bd_ram_mem2_reg[89][19]/P0001 , \wishbone_bd_ram_mem2_reg[89][20]/P0001 , \wishbone_bd_ram_mem2_reg[89][21]/P0001 , \wishbone_bd_ram_mem2_reg[89][22]/P0001 , \wishbone_bd_ram_mem2_reg[89][23]/P0001 , \wishbone_bd_ram_mem2_reg[8][16]/P0001 , \wishbone_bd_ram_mem2_reg[8][17]/P0001 , \wishbone_bd_ram_mem2_reg[8][18]/P0001 , \wishbone_bd_ram_mem2_reg[8][19]/P0001 , \wishbone_bd_ram_mem2_reg[8][20]/P0001 , \wishbone_bd_ram_mem2_reg[8][21]/P0001 , \wishbone_bd_ram_mem2_reg[8][22]/P0001 , \wishbone_bd_ram_mem2_reg[8][23]/P0001 , \wishbone_bd_ram_mem2_reg[90][16]/P0001 , \wishbone_bd_ram_mem2_reg[90][17]/P0001 , \wishbone_bd_ram_mem2_reg[90][18]/P0001 , \wishbone_bd_ram_mem2_reg[90][19]/P0001 , \wishbone_bd_ram_mem2_reg[90][20]/P0001 , \wishbone_bd_ram_mem2_reg[90][21]/P0001 , \wishbone_bd_ram_mem2_reg[90][22]/P0001 , \wishbone_bd_ram_mem2_reg[90][23]/P0001 , \wishbone_bd_ram_mem2_reg[91][16]/P0001 , \wishbone_bd_ram_mem2_reg[91][17]/P0001 , \wishbone_bd_ram_mem2_reg[91][18]/P0001 , \wishbone_bd_ram_mem2_reg[91][19]/P0001 , \wishbone_bd_ram_mem2_reg[91][20]/P0001 , \wishbone_bd_ram_mem2_reg[91][21]/P0001 , \wishbone_bd_ram_mem2_reg[91][22]/P0001 , \wishbone_bd_ram_mem2_reg[91][23]/P0001 , \wishbone_bd_ram_mem2_reg[92][16]/P0001 , \wishbone_bd_ram_mem2_reg[92][17]/P0001 , \wishbone_bd_ram_mem2_reg[92][18]/P0001 , \wishbone_bd_ram_mem2_reg[92][19]/P0001 , \wishbone_bd_ram_mem2_reg[92][20]/P0001 , \wishbone_bd_ram_mem2_reg[92][21]/P0001 , \wishbone_bd_ram_mem2_reg[92][22]/P0001 , \wishbone_bd_ram_mem2_reg[92][23]/P0001 , \wishbone_bd_ram_mem2_reg[93][16]/P0001 , \wishbone_bd_ram_mem2_reg[93][17]/P0001 , \wishbone_bd_ram_mem2_reg[93][18]/P0001 , \wishbone_bd_ram_mem2_reg[93][19]/P0001 , \wishbone_bd_ram_mem2_reg[93][20]/P0001 , \wishbone_bd_ram_mem2_reg[93][21]/P0001 , \wishbone_bd_ram_mem2_reg[93][22]/P0001 , \wishbone_bd_ram_mem2_reg[93][23]/P0001 , \wishbone_bd_ram_mem2_reg[94][16]/P0001 , \wishbone_bd_ram_mem2_reg[94][17]/P0001 , \wishbone_bd_ram_mem2_reg[94][18]/P0001 , \wishbone_bd_ram_mem2_reg[94][19]/P0001 , \wishbone_bd_ram_mem2_reg[94][20]/P0001 , \wishbone_bd_ram_mem2_reg[94][21]/P0001 , \wishbone_bd_ram_mem2_reg[94][22]/P0001 , \wishbone_bd_ram_mem2_reg[94][23]/P0001 , \wishbone_bd_ram_mem2_reg[95][16]/P0001 , \wishbone_bd_ram_mem2_reg[95][17]/P0001 , \wishbone_bd_ram_mem2_reg[95][18]/P0001 , \wishbone_bd_ram_mem2_reg[95][19]/P0001 , \wishbone_bd_ram_mem2_reg[95][20]/P0001 , \wishbone_bd_ram_mem2_reg[95][21]/P0001 , \wishbone_bd_ram_mem2_reg[95][22]/P0001 , \wishbone_bd_ram_mem2_reg[95][23]/P0001 , \wishbone_bd_ram_mem2_reg[96][16]/P0001 , \wishbone_bd_ram_mem2_reg[96][17]/P0001 , \wishbone_bd_ram_mem2_reg[96][18]/P0001 , \wishbone_bd_ram_mem2_reg[96][19]/P0001 , \wishbone_bd_ram_mem2_reg[96][20]/P0001 , \wishbone_bd_ram_mem2_reg[96][21]/P0001 , \wishbone_bd_ram_mem2_reg[96][22]/P0001 , \wishbone_bd_ram_mem2_reg[96][23]/P0001 , \wishbone_bd_ram_mem2_reg[97][16]/P0001 , \wishbone_bd_ram_mem2_reg[97][17]/P0001 , \wishbone_bd_ram_mem2_reg[97][18]/P0001 , \wishbone_bd_ram_mem2_reg[97][19]/P0001 , \wishbone_bd_ram_mem2_reg[97][20]/P0001 , \wishbone_bd_ram_mem2_reg[97][21]/P0001 , \wishbone_bd_ram_mem2_reg[97][22]/P0001 , \wishbone_bd_ram_mem2_reg[97][23]/P0001 , \wishbone_bd_ram_mem2_reg[98][16]/P0001 , \wishbone_bd_ram_mem2_reg[98][17]/P0001 , \wishbone_bd_ram_mem2_reg[98][18]/P0001 , \wishbone_bd_ram_mem2_reg[98][19]/P0001 , \wishbone_bd_ram_mem2_reg[98][20]/P0001 , \wishbone_bd_ram_mem2_reg[98][21]/P0001 , \wishbone_bd_ram_mem2_reg[98][22]/P0001 , \wishbone_bd_ram_mem2_reg[98][23]/P0001 , \wishbone_bd_ram_mem2_reg[99][16]/P0001 , \wishbone_bd_ram_mem2_reg[99][17]/P0001 , \wishbone_bd_ram_mem2_reg[99][18]/P0001 , \wishbone_bd_ram_mem2_reg[99][19]/P0001 , \wishbone_bd_ram_mem2_reg[99][20]/P0001 , \wishbone_bd_ram_mem2_reg[99][21]/P0001 , \wishbone_bd_ram_mem2_reg[99][22]/P0001 , \wishbone_bd_ram_mem2_reg[99][23]/P0001 , \wishbone_bd_ram_mem2_reg[9][16]/P0001 , \wishbone_bd_ram_mem2_reg[9][17]/P0001 , \wishbone_bd_ram_mem2_reg[9][18]/P0001 , \wishbone_bd_ram_mem2_reg[9][19]/P0001 , \wishbone_bd_ram_mem2_reg[9][20]/P0001 , \wishbone_bd_ram_mem2_reg[9][21]/P0001 , \wishbone_bd_ram_mem2_reg[9][22]/P0001 , \wishbone_bd_ram_mem2_reg[9][23]/P0001 , \wishbone_bd_ram_mem3_reg[0][24]/P0001 , \wishbone_bd_ram_mem3_reg[0][25]/P0001 , \wishbone_bd_ram_mem3_reg[0][26]/P0001 , \wishbone_bd_ram_mem3_reg[0][27]/P0001 , \wishbone_bd_ram_mem3_reg[0][28]/P0001 , \wishbone_bd_ram_mem3_reg[0][29]/P0001 , \wishbone_bd_ram_mem3_reg[0][30]/P0001 , \wishbone_bd_ram_mem3_reg[0][31]/P0001 , \wishbone_bd_ram_mem3_reg[100][24]/P0001 , \wishbone_bd_ram_mem3_reg[100][25]/P0001 , \wishbone_bd_ram_mem3_reg[100][26]/P0001 , \wishbone_bd_ram_mem3_reg[100][27]/P0001 , \wishbone_bd_ram_mem3_reg[100][28]/P0001 , \wishbone_bd_ram_mem3_reg[100][29]/P0001 , \wishbone_bd_ram_mem3_reg[100][30]/P0001 , \wishbone_bd_ram_mem3_reg[100][31]/P0001 , \wishbone_bd_ram_mem3_reg[101][24]/P0001 , \wishbone_bd_ram_mem3_reg[101][25]/P0001 , \wishbone_bd_ram_mem3_reg[101][26]/P0001 , \wishbone_bd_ram_mem3_reg[101][27]/P0001 , \wishbone_bd_ram_mem3_reg[101][28]/P0001 , \wishbone_bd_ram_mem3_reg[101][29]/P0001 , \wishbone_bd_ram_mem3_reg[101][30]/P0001 , \wishbone_bd_ram_mem3_reg[101][31]/P0001 , \wishbone_bd_ram_mem3_reg[102][24]/P0001 , \wishbone_bd_ram_mem3_reg[102][25]/P0001 , \wishbone_bd_ram_mem3_reg[102][26]/P0001 , \wishbone_bd_ram_mem3_reg[102][27]/P0001 , \wishbone_bd_ram_mem3_reg[102][28]/P0001 , \wishbone_bd_ram_mem3_reg[102][29]/P0001 , \wishbone_bd_ram_mem3_reg[102][30]/P0001 , \wishbone_bd_ram_mem3_reg[102][31]/P0001 , \wishbone_bd_ram_mem3_reg[103][24]/P0001 , \wishbone_bd_ram_mem3_reg[103][25]/P0001 , \wishbone_bd_ram_mem3_reg[103][26]/P0001 , \wishbone_bd_ram_mem3_reg[103][27]/P0001 , \wishbone_bd_ram_mem3_reg[103][28]/P0001 , \wishbone_bd_ram_mem3_reg[103][29]/P0001 , \wishbone_bd_ram_mem3_reg[103][30]/P0001 , \wishbone_bd_ram_mem3_reg[103][31]/P0001 , \wishbone_bd_ram_mem3_reg[104][24]/P0001 , \wishbone_bd_ram_mem3_reg[104][25]/P0001 , \wishbone_bd_ram_mem3_reg[104][26]/P0001 , \wishbone_bd_ram_mem3_reg[104][27]/P0001 , \wishbone_bd_ram_mem3_reg[104][28]/P0001 , \wishbone_bd_ram_mem3_reg[104][29]/P0001 , \wishbone_bd_ram_mem3_reg[104][30]/P0001 , \wishbone_bd_ram_mem3_reg[104][31]/P0001 , \wishbone_bd_ram_mem3_reg[105][24]/P0001 , \wishbone_bd_ram_mem3_reg[105][25]/P0001 , \wishbone_bd_ram_mem3_reg[105][26]/P0001 , \wishbone_bd_ram_mem3_reg[105][27]/P0001 , \wishbone_bd_ram_mem3_reg[105][28]/P0001 , \wishbone_bd_ram_mem3_reg[105][29]/P0001 , \wishbone_bd_ram_mem3_reg[105][30]/P0001 , \wishbone_bd_ram_mem3_reg[105][31]/P0001 , \wishbone_bd_ram_mem3_reg[106][24]/P0001 , \wishbone_bd_ram_mem3_reg[106][25]/P0001 , \wishbone_bd_ram_mem3_reg[106][26]/P0001 , \wishbone_bd_ram_mem3_reg[106][27]/P0001 , \wishbone_bd_ram_mem3_reg[106][28]/P0001 , \wishbone_bd_ram_mem3_reg[106][29]/P0001 , \wishbone_bd_ram_mem3_reg[106][30]/P0001 , \wishbone_bd_ram_mem3_reg[106][31]/P0001 , \wishbone_bd_ram_mem3_reg[107][24]/P0001 , \wishbone_bd_ram_mem3_reg[107][25]/P0001 , \wishbone_bd_ram_mem3_reg[107][26]/P0001 , \wishbone_bd_ram_mem3_reg[107][27]/P0001 , \wishbone_bd_ram_mem3_reg[107][28]/P0001 , \wishbone_bd_ram_mem3_reg[107][29]/P0001 , \wishbone_bd_ram_mem3_reg[107][30]/P0001 , \wishbone_bd_ram_mem3_reg[107][31]/P0001 , \wishbone_bd_ram_mem3_reg[108][24]/P0001 , \wishbone_bd_ram_mem3_reg[108][25]/P0001 , \wishbone_bd_ram_mem3_reg[108][26]/P0001 , \wishbone_bd_ram_mem3_reg[108][27]/P0001 , \wishbone_bd_ram_mem3_reg[108][28]/P0001 , \wishbone_bd_ram_mem3_reg[108][29]/P0001 , \wishbone_bd_ram_mem3_reg[108][30]/P0001 , \wishbone_bd_ram_mem3_reg[108][31]/P0001 , \wishbone_bd_ram_mem3_reg[109][24]/P0001 , \wishbone_bd_ram_mem3_reg[109][25]/P0001 , \wishbone_bd_ram_mem3_reg[109][26]/P0001 , \wishbone_bd_ram_mem3_reg[109][27]/P0001 , \wishbone_bd_ram_mem3_reg[109][28]/P0001 , \wishbone_bd_ram_mem3_reg[109][29]/P0001 , \wishbone_bd_ram_mem3_reg[109][30]/P0001 , \wishbone_bd_ram_mem3_reg[109][31]/P0001 , \wishbone_bd_ram_mem3_reg[10][24]/P0001 , \wishbone_bd_ram_mem3_reg[10][25]/P0001 , \wishbone_bd_ram_mem3_reg[10][26]/P0001 , \wishbone_bd_ram_mem3_reg[10][27]/P0001 , \wishbone_bd_ram_mem3_reg[10][28]/P0001 , \wishbone_bd_ram_mem3_reg[10][29]/P0001 , \wishbone_bd_ram_mem3_reg[10][30]/P0001 , \wishbone_bd_ram_mem3_reg[10][31]/P0001 , \wishbone_bd_ram_mem3_reg[110][24]/P0001 , \wishbone_bd_ram_mem3_reg[110][25]/P0001 , \wishbone_bd_ram_mem3_reg[110][26]/P0001 , \wishbone_bd_ram_mem3_reg[110][27]/P0001 , \wishbone_bd_ram_mem3_reg[110][28]/P0001 , \wishbone_bd_ram_mem3_reg[110][29]/P0001 , \wishbone_bd_ram_mem3_reg[110][30]/P0001 , \wishbone_bd_ram_mem3_reg[110][31]/P0001 , \wishbone_bd_ram_mem3_reg[111][24]/P0001 , \wishbone_bd_ram_mem3_reg[111][25]/P0001 , \wishbone_bd_ram_mem3_reg[111][26]/P0001 , \wishbone_bd_ram_mem3_reg[111][27]/P0001 , \wishbone_bd_ram_mem3_reg[111][28]/P0001 , \wishbone_bd_ram_mem3_reg[111][29]/P0001 , \wishbone_bd_ram_mem3_reg[111][30]/P0001 , \wishbone_bd_ram_mem3_reg[111][31]/P0001 , \wishbone_bd_ram_mem3_reg[112][24]/P0001 , \wishbone_bd_ram_mem3_reg[112][25]/P0001 , \wishbone_bd_ram_mem3_reg[112][26]/P0001 , \wishbone_bd_ram_mem3_reg[112][27]/P0001 , \wishbone_bd_ram_mem3_reg[112][28]/P0001 , \wishbone_bd_ram_mem3_reg[112][29]/P0001 , \wishbone_bd_ram_mem3_reg[112][30]/P0001 , \wishbone_bd_ram_mem3_reg[112][31]/P0001 , \wishbone_bd_ram_mem3_reg[113][24]/P0001 , \wishbone_bd_ram_mem3_reg[113][25]/P0001 , \wishbone_bd_ram_mem3_reg[113][26]/P0001 , \wishbone_bd_ram_mem3_reg[113][27]/P0001 , \wishbone_bd_ram_mem3_reg[113][28]/P0001 , \wishbone_bd_ram_mem3_reg[113][29]/P0001 , \wishbone_bd_ram_mem3_reg[113][30]/P0001 , \wishbone_bd_ram_mem3_reg[113][31]/P0001 , \wishbone_bd_ram_mem3_reg[114][24]/P0001 , \wishbone_bd_ram_mem3_reg[114][25]/P0001 , \wishbone_bd_ram_mem3_reg[114][26]/P0001 , \wishbone_bd_ram_mem3_reg[114][27]/P0001 , \wishbone_bd_ram_mem3_reg[114][28]/P0001 , \wishbone_bd_ram_mem3_reg[114][29]/P0001 , \wishbone_bd_ram_mem3_reg[114][30]/P0001 , \wishbone_bd_ram_mem3_reg[114][31]/P0001 , \wishbone_bd_ram_mem3_reg[115][24]/P0001 , \wishbone_bd_ram_mem3_reg[115][25]/P0001 , \wishbone_bd_ram_mem3_reg[115][26]/P0001 , \wishbone_bd_ram_mem3_reg[115][27]/P0001 , \wishbone_bd_ram_mem3_reg[115][28]/P0001 , \wishbone_bd_ram_mem3_reg[115][29]/P0001 , \wishbone_bd_ram_mem3_reg[115][30]/P0001 , \wishbone_bd_ram_mem3_reg[115][31]/P0001 , \wishbone_bd_ram_mem3_reg[116][24]/P0001 , \wishbone_bd_ram_mem3_reg[116][25]/P0001 , \wishbone_bd_ram_mem3_reg[116][26]/P0001 , \wishbone_bd_ram_mem3_reg[116][27]/P0001 , \wishbone_bd_ram_mem3_reg[116][28]/P0001 , \wishbone_bd_ram_mem3_reg[116][29]/P0001 , \wishbone_bd_ram_mem3_reg[116][30]/P0001 , \wishbone_bd_ram_mem3_reg[116][31]/P0001 , \wishbone_bd_ram_mem3_reg[117][24]/P0001 , \wishbone_bd_ram_mem3_reg[117][25]/P0001 , \wishbone_bd_ram_mem3_reg[117][26]/P0001 , \wishbone_bd_ram_mem3_reg[117][27]/P0001 , \wishbone_bd_ram_mem3_reg[117][28]/P0001 , \wishbone_bd_ram_mem3_reg[117][29]/P0001 , \wishbone_bd_ram_mem3_reg[117][30]/P0001 , \wishbone_bd_ram_mem3_reg[117][31]/P0001 , \wishbone_bd_ram_mem3_reg[118][24]/P0001 , \wishbone_bd_ram_mem3_reg[118][25]/P0001 , \wishbone_bd_ram_mem3_reg[118][26]/P0001 , \wishbone_bd_ram_mem3_reg[118][27]/P0001 , \wishbone_bd_ram_mem3_reg[118][28]/P0001 , \wishbone_bd_ram_mem3_reg[118][29]/P0001 , \wishbone_bd_ram_mem3_reg[118][30]/P0001 , \wishbone_bd_ram_mem3_reg[118][31]/P0001 , \wishbone_bd_ram_mem3_reg[119][24]/P0001 , \wishbone_bd_ram_mem3_reg[119][25]/P0001 , \wishbone_bd_ram_mem3_reg[119][26]/P0001 , \wishbone_bd_ram_mem3_reg[119][27]/P0001 , \wishbone_bd_ram_mem3_reg[119][28]/P0001 , \wishbone_bd_ram_mem3_reg[119][29]/P0001 , \wishbone_bd_ram_mem3_reg[119][30]/P0001 , \wishbone_bd_ram_mem3_reg[119][31]/P0001 , \wishbone_bd_ram_mem3_reg[11][24]/P0001 , \wishbone_bd_ram_mem3_reg[11][25]/P0001 , \wishbone_bd_ram_mem3_reg[11][26]/P0001 , \wishbone_bd_ram_mem3_reg[11][27]/P0001 , \wishbone_bd_ram_mem3_reg[11][28]/P0001 , \wishbone_bd_ram_mem3_reg[11][29]/P0001 , \wishbone_bd_ram_mem3_reg[11][30]/P0001 , \wishbone_bd_ram_mem3_reg[11][31]/P0001 , \wishbone_bd_ram_mem3_reg[120][24]/P0001 , \wishbone_bd_ram_mem3_reg[120][25]/P0001 , \wishbone_bd_ram_mem3_reg[120][26]/P0001 , \wishbone_bd_ram_mem3_reg[120][27]/P0001 , \wishbone_bd_ram_mem3_reg[120][28]/P0001 , \wishbone_bd_ram_mem3_reg[120][29]/P0001 , \wishbone_bd_ram_mem3_reg[120][30]/P0001 , \wishbone_bd_ram_mem3_reg[120][31]/P0001 , \wishbone_bd_ram_mem3_reg[121][24]/P0001 , \wishbone_bd_ram_mem3_reg[121][25]/P0001 , \wishbone_bd_ram_mem3_reg[121][26]/P0001 , \wishbone_bd_ram_mem3_reg[121][27]/P0001 , \wishbone_bd_ram_mem3_reg[121][28]/P0001 , \wishbone_bd_ram_mem3_reg[121][29]/P0001 , \wishbone_bd_ram_mem3_reg[121][30]/P0001 , \wishbone_bd_ram_mem3_reg[121][31]/P0001 , \wishbone_bd_ram_mem3_reg[122][24]/P0001 , \wishbone_bd_ram_mem3_reg[122][25]/P0001 , \wishbone_bd_ram_mem3_reg[122][26]/P0001 , \wishbone_bd_ram_mem3_reg[122][27]/P0001 , \wishbone_bd_ram_mem3_reg[122][28]/P0001 , \wishbone_bd_ram_mem3_reg[122][29]/P0001 , \wishbone_bd_ram_mem3_reg[122][30]/P0001 , \wishbone_bd_ram_mem3_reg[122][31]/P0001 , \wishbone_bd_ram_mem3_reg[123][24]/P0001 , \wishbone_bd_ram_mem3_reg[123][25]/P0001 , \wishbone_bd_ram_mem3_reg[123][26]/P0001 , \wishbone_bd_ram_mem3_reg[123][27]/P0001 , \wishbone_bd_ram_mem3_reg[123][28]/P0001 , \wishbone_bd_ram_mem3_reg[123][29]/P0001 , \wishbone_bd_ram_mem3_reg[123][30]/P0001 , \wishbone_bd_ram_mem3_reg[123][31]/P0001 , \wishbone_bd_ram_mem3_reg[124][24]/P0001 , \wishbone_bd_ram_mem3_reg[124][25]/P0001 , \wishbone_bd_ram_mem3_reg[124][26]/P0001 , \wishbone_bd_ram_mem3_reg[124][27]/P0001 , \wishbone_bd_ram_mem3_reg[124][28]/P0001 , \wishbone_bd_ram_mem3_reg[124][29]/P0001 , \wishbone_bd_ram_mem3_reg[124][30]/P0001 , \wishbone_bd_ram_mem3_reg[124][31]/P0001 , \wishbone_bd_ram_mem3_reg[125][24]/P0001 , \wishbone_bd_ram_mem3_reg[125][25]/P0001 , \wishbone_bd_ram_mem3_reg[125][26]/P0001 , \wishbone_bd_ram_mem3_reg[125][27]/P0001 , \wishbone_bd_ram_mem3_reg[125][28]/P0001 , \wishbone_bd_ram_mem3_reg[125][29]/P0001 , \wishbone_bd_ram_mem3_reg[125][30]/P0001 , \wishbone_bd_ram_mem3_reg[125][31]/P0001 , \wishbone_bd_ram_mem3_reg[126][24]/P0001 , \wishbone_bd_ram_mem3_reg[126][25]/P0001 , \wishbone_bd_ram_mem3_reg[126][26]/P0001 , \wishbone_bd_ram_mem3_reg[126][27]/P0001 , \wishbone_bd_ram_mem3_reg[126][28]/P0001 , \wishbone_bd_ram_mem3_reg[126][29]/P0001 , \wishbone_bd_ram_mem3_reg[126][30]/P0001 , \wishbone_bd_ram_mem3_reg[126][31]/P0001 , \wishbone_bd_ram_mem3_reg[127][24]/P0001 , \wishbone_bd_ram_mem3_reg[127][25]/P0001 , \wishbone_bd_ram_mem3_reg[127][26]/P0001 , \wishbone_bd_ram_mem3_reg[127][27]/P0001 , \wishbone_bd_ram_mem3_reg[127][28]/P0001 , \wishbone_bd_ram_mem3_reg[127][29]/P0001 , \wishbone_bd_ram_mem3_reg[127][30]/P0001 , \wishbone_bd_ram_mem3_reg[127][31]/P0001 , \wishbone_bd_ram_mem3_reg[128][24]/P0001 , \wishbone_bd_ram_mem3_reg[128][25]/P0001 , \wishbone_bd_ram_mem3_reg[128][26]/P0001 , \wishbone_bd_ram_mem3_reg[128][27]/P0001 , \wishbone_bd_ram_mem3_reg[128][28]/P0001 , \wishbone_bd_ram_mem3_reg[128][29]/P0001 , \wishbone_bd_ram_mem3_reg[128][30]/P0001 , \wishbone_bd_ram_mem3_reg[128][31]/P0001 , \wishbone_bd_ram_mem3_reg[129][24]/P0001 , \wishbone_bd_ram_mem3_reg[129][25]/P0001 , \wishbone_bd_ram_mem3_reg[129][26]/P0001 , \wishbone_bd_ram_mem3_reg[129][27]/P0001 , \wishbone_bd_ram_mem3_reg[129][28]/P0001 , \wishbone_bd_ram_mem3_reg[129][29]/P0001 , \wishbone_bd_ram_mem3_reg[129][30]/P0001 , \wishbone_bd_ram_mem3_reg[129][31]/P0001 , \wishbone_bd_ram_mem3_reg[12][24]/P0001 , \wishbone_bd_ram_mem3_reg[12][25]/P0001 , \wishbone_bd_ram_mem3_reg[12][26]/P0001 , \wishbone_bd_ram_mem3_reg[12][27]/P0001 , \wishbone_bd_ram_mem3_reg[12][28]/P0001 , \wishbone_bd_ram_mem3_reg[12][29]/P0001 , \wishbone_bd_ram_mem3_reg[12][30]/P0001 , \wishbone_bd_ram_mem3_reg[12][31]/P0001 , \wishbone_bd_ram_mem3_reg[130][24]/P0001 , \wishbone_bd_ram_mem3_reg[130][25]/P0001 , \wishbone_bd_ram_mem3_reg[130][26]/P0001 , \wishbone_bd_ram_mem3_reg[130][27]/P0001 , \wishbone_bd_ram_mem3_reg[130][28]/P0001 , \wishbone_bd_ram_mem3_reg[130][29]/P0001 , \wishbone_bd_ram_mem3_reg[130][30]/P0001 , \wishbone_bd_ram_mem3_reg[130][31]/P0001 , \wishbone_bd_ram_mem3_reg[131][24]/P0001 , \wishbone_bd_ram_mem3_reg[131][25]/P0001 , \wishbone_bd_ram_mem3_reg[131][26]/P0001 , \wishbone_bd_ram_mem3_reg[131][27]/P0001 , \wishbone_bd_ram_mem3_reg[131][28]/P0001 , \wishbone_bd_ram_mem3_reg[131][29]/P0001 , \wishbone_bd_ram_mem3_reg[131][30]/P0001 , \wishbone_bd_ram_mem3_reg[131][31]/P0001 , \wishbone_bd_ram_mem3_reg[132][24]/P0001 , \wishbone_bd_ram_mem3_reg[132][25]/P0001 , \wishbone_bd_ram_mem3_reg[132][26]/P0001 , \wishbone_bd_ram_mem3_reg[132][27]/P0001 , \wishbone_bd_ram_mem3_reg[132][28]/P0001 , \wishbone_bd_ram_mem3_reg[132][29]/P0001 , \wishbone_bd_ram_mem3_reg[132][30]/P0001 , \wishbone_bd_ram_mem3_reg[132][31]/P0001 , \wishbone_bd_ram_mem3_reg[133][24]/P0001 , \wishbone_bd_ram_mem3_reg[133][25]/P0001 , \wishbone_bd_ram_mem3_reg[133][26]/P0001 , \wishbone_bd_ram_mem3_reg[133][27]/P0001 , \wishbone_bd_ram_mem3_reg[133][28]/P0001 , \wishbone_bd_ram_mem3_reg[133][29]/P0001 , \wishbone_bd_ram_mem3_reg[133][30]/P0001 , \wishbone_bd_ram_mem3_reg[133][31]/P0001 , \wishbone_bd_ram_mem3_reg[134][24]/P0001 , \wishbone_bd_ram_mem3_reg[134][25]/P0001 , \wishbone_bd_ram_mem3_reg[134][26]/P0001 , \wishbone_bd_ram_mem3_reg[134][27]/P0001 , \wishbone_bd_ram_mem3_reg[134][28]/P0001 , \wishbone_bd_ram_mem3_reg[134][29]/P0001 , \wishbone_bd_ram_mem3_reg[134][30]/P0001 , \wishbone_bd_ram_mem3_reg[134][31]/P0001 , \wishbone_bd_ram_mem3_reg[135][24]/P0001 , \wishbone_bd_ram_mem3_reg[135][25]/P0001 , \wishbone_bd_ram_mem3_reg[135][26]/P0001 , \wishbone_bd_ram_mem3_reg[135][27]/P0001 , \wishbone_bd_ram_mem3_reg[135][28]/P0001 , \wishbone_bd_ram_mem3_reg[135][29]/P0001 , \wishbone_bd_ram_mem3_reg[135][30]/P0001 , \wishbone_bd_ram_mem3_reg[135][31]/P0001 , \wishbone_bd_ram_mem3_reg[136][24]/P0001 , \wishbone_bd_ram_mem3_reg[136][25]/P0001 , \wishbone_bd_ram_mem3_reg[136][26]/P0001 , \wishbone_bd_ram_mem3_reg[136][27]/P0001 , \wishbone_bd_ram_mem3_reg[136][28]/P0001 , \wishbone_bd_ram_mem3_reg[136][29]/P0001 , \wishbone_bd_ram_mem3_reg[136][30]/P0001 , \wishbone_bd_ram_mem3_reg[136][31]/P0001 , \wishbone_bd_ram_mem3_reg[137][24]/P0001 , \wishbone_bd_ram_mem3_reg[137][25]/P0001 , \wishbone_bd_ram_mem3_reg[137][26]/P0001 , \wishbone_bd_ram_mem3_reg[137][27]/P0001 , \wishbone_bd_ram_mem3_reg[137][28]/P0001 , \wishbone_bd_ram_mem3_reg[137][29]/P0001 , \wishbone_bd_ram_mem3_reg[137][30]/P0001 , \wishbone_bd_ram_mem3_reg[137][31]/P0001 , \wishbone_bd_ram_mem3_reg[138][24]/P0001 , \wishbone_bd_ram_mem3_reg[138][25]/P0001 , \wishbone_bd_ram_mem3_reg[138][26]/P0001 , \wishbone_bd_ram_mem3_reg[138][27]/P0001 , \wishbone_bd_ram_mem3_reg[138][28]/P0001 , \wishbone_bd_ram_mem3_reg[138][29]/P0001 , \wishbone_bd_ram_mem3_reg[138][30]/P0001 , \wishbone_bd_ram_mem3_reg[138][31]/P0001 , \wishbone_bd_ram_mem3_reg[139][24]/P0001 , \wishbone_bd_ram_mem3_reg[139][25]/P0001 , \wishbone_bd_ram_mem3_reg[139][26]/P0001 , \wishbone_bd_ram_mem3_reg[139][27]/P0001 , \wishbone_bd_ram_mem3_reg[139][28]/P0001 , \wishbone_bd_ram_mem3_reg[139][29]/P0001 , \wishbone_bd_ram_mem3_reg[139][30]/P0001 , \wishbone_bd_ram_mem3_reg[139][31]/P0001 , \wishbone_bd_ram_mem3_reg[13][24]/P0001 , \wishbone_bd_ram_mem3_reg[13][25]/P0001 , \wishbone_bd_ram_mem3_reg[13][26]/P0001 , \wishbone_bd_ram_mem3_reg[13][27]/P0001 , \wishbone_bd_ram_mem3_reg[13][28]/P0001 , \wishbone_bd_ram_mem3_reg[13][29]/P0001 , \wishbone_bd_ram_mem3_reg[13][30]/P0001 , \wishbone_bd_ram_mem3_reg[13][31]/P0001 , \wishbone_bd_ram_mem3_reg[140][24]/P0001 , \wishbone_bd_ram_mem3_reg[140][25]/P0001 , \wishbone_bd_ram_mem3_reg[140][26]/P0001 , \wishbone_bd_ram_mem3_reg[140][27]/P0001 , \wishbone_bd_ram_mem3_reg[140][28]/P0001 , \wishbone_bd_ram_mem3_reg[140][29]/P0001 , \wishbone_bd_ram_mem3_reg[140][30]/P0001 , \wishbone_bd_ram_mem3_reg[140][31]/P0001 , \wishbone_bd_ram_mem3_reg[141][24]/P0001 , \wishbone_bd_ram_mem3_reg[141][25]/P0001 , \wishbone_bd_ram_mem3_reg[141][26]/P0001 , \wishbone_bd_ram_mem3_reg[141][27]/P0001 , \wishbone_bd_ram_mem3_reg[141][28]/P0001 , \wishbone_bd_ram_mem3_reg[141][29]/P0001 , \wishbone_bd_ram_mem3_reg[141][30]/P0001 , \wishbone_bd_ram_mem3_reg[141][31]/P0001 , \wishbone_bd_ram_mem3_reg[142][24]/P0001 , \wishbone_bd_ram_mem3_reg[142][25]/P0001 , \wishbone_bd_ram_mem3_reg[142][26]/P0001 , \wishbone_bd_ram_mem3_reg[142][27]/P0001 , \wishbone_bd_ram_mem3_reg[142][28]/P0001 , \wishbone_bd_ram_mem3_reg[142][29]/P0001 , \wishbone_bd_ram_mem3_reg[142][30]/P0001 , \wishbone_bd_ram_mem3_reg[142][31]/P0001 , \wishbone_bd_ram_mem3_reg[143][24]/P0001 , \wishbone_bd_ram_mem3_reg[143][25]/P0001 , \wishbone_bd_ram_mem3_reg[143][26]/P0001 , \wishbone_bd_ram_mem3_reg[143][27]/P0001 , \wishbone_bd_ram_mem3_reg[143][28]/P0001 , \wishbone_bd_ram_mem3_reg[143][29]/P0001 , \wishbone_bd_ram_mem3_reg[143][30]/P0001 , \wishbone_bd_ram_mem3_reg[143][31]/P0001 , \wishbone_bd_ram_mem3_reg[144][24]/P0001 , \wishbone_bd_ram_mem3_reg[144][25]/P0001 , \wishbone_bd_ram_mem3_reg[144][26]/P0001 , \wishbone_bd_ram_mem3_reg[144][27]/P0001 , \wishbone_bd_ram_mem3_reg[144][28]/P0001 , \wishbone_bd_ram_mem3_reg[144][29]/P0001 , \wishbone_bd_ram_mem3_reg[144][30]/P0001 , \wishbone_bd_ram_mem3_reg[144][31]/P0001 , \wishbone_bd_ram_mem3_reg[145][24]/P0001 , \wishbone_bd_ram_mem3_reg[145][25]/P0001 , \wishbone_bd_ram_mem3_reg[145][26]/P0001 , \wishbone_bd_ram_mem3_reg[145][27]/P0001 , \wishbone_bd_ram_mem3_reg[145][28]/P0001 , \wishbone_bd_ram_mem3_reg[145][29]/P0001 , \wishbone_bd_ram_mem3_reg[145][30]/P0001 , \wishbone_bd_ram_mem3_reg[145][31]/P0001 , \wishbone_bd_ram_mem3_reg[146][24]/P0001 , \wishbone_bd_ram_mem3_reg[146][25]/P0001 , \wishbone_bd_ram_mem3_reg[146][26]/P0001 , \wishbone_bd_ram_mem3_reg[146][27]/P0001 , \wishbone_bd_ram_mem3_reg[146][28]/P0001 , \wishbone_bd_ram_mem3_reg[146][29]/P0001 , \wishbone_bd_ram_mem3_reg[146][30]/P0001 , \wishbone_bd_ram_mem3_reg[146][31]/P0001 , \wishbone_bd_ram_mem3_reg[147][24]/P0001 , \wishbone_bd_ram_mem3_reg[147][25]/P0001 , \wishbone_bd_ram_mem3_reg[147][26]/P0001 , \wishbone_bd_ram_mem3_reg[147][27]/P0001 , \wishbone_bd_ram_mem3_reg[147][28]/P0001 , \wishbone_bd_ram_mem3_reg[147][29]/P0001 , \wishbone_bd_ram_mem3_reg[147][30]/P0001 , \wishbone_bd_ram_mem3_reg[147][31]/P0001 , \wishbone_bd_ram_mem3_reg[148][24]/P0001 , \wishbone_bd_ram_mem3_reg[148][25]/P0001 , \wishbone_bd_ram_mem3_reg[148][26]/P0001 , \wishbone_bd_ram_mem3_reg[148][27]/P0001 , \wishbone_bd_ram_mem3_reg[148][28]/P0001 , \wishbone_bd_ram_mem3_reg[148][29]/P0001 , \wishbone_bd_ram_mem3_reg[148][30]/P0001 , \wishbone_bd_ram_mem3_reg[148][31]/P0001 , \wishbone_bd_ram_mem3_reg[149][24]/P0001 , \wishbone_bd_ram_mem3_reg[149][25]/P0001 , \wishbone_bd_ram_mem3_reg[149][26]/P0001 , \wishbone_bd_ram_mem3_reg[149][27]/P0001 , \wishbone_bd_ram_mem3_reg[149][28]/P0001 , \wishbone_bd_ram_mem3_reg[149][29]/P0001 , \wishbone_bd_ram_mem3_reg[149][30]/P0001 , \wishbone_bd_ram_mem3_reg[149][31]/P0001 , \wishbone_bd_ram_mem3_reg[14][24]/P0001 , \wishbone_bd_ram_mem3_reg[14][25]/P0001 , \wishbone_bd_ram_mem3_reg[14][26]/P0001 , \wishbone_bd_ram_mem3_reg[14][27]/P0001 , \wishbone_bd_ram_mem3_reg[14][28]/P0001 , \wishbone_bd_ram_mem3_reg[14][29]/P0001 , \wishbone_bd_ram_mem3_reg[14][30]/P0001 , \wishbone_bd_ram_mem3_reg[14][31]/P0001 , \wishbone_bd_ram_mem3_reg[150][24]/P0001 , \wishbone_bd_ram_mem3_reg[150][25]/P0001 , \wishbone_bd_ram_mem3_reg[150][26]/P0001 , \wishbone_bd_ram_mem3_reg[150][27]/P0001 , \wishbone_bd_ram_mem3_reg[150][28]/P0001 , \wishbone_bd_ram_mem3_reg[150][29]/P0001 , \wishbone_bd_ram_mem3_reg[150][30]/P0001 , \wishbone_bd_ram_mem3_reg[150][31]/P0001 , \wishbone_bd_ram_mem3_reg[151][24]/P0001 , \wishbone_bd_ram_mem3_reg[151][25]/P0001 , \wishbone_bd_ram_mem3_reg[151][26]/P0001 , \wishbone_bd_ram_mem3_reg[151][27]/P0001 , \wishbone_bd_ram_mem3_reg[151][28]/P0001 , \wishbone_bd_ram_mem3_reg[151][29]/P0001 , \wishbone_bd_ram_mem3_reg[151][30]/P0001 , \wishbone_bd_ram_mem3_reg[151][31]/P0001 , \wishbone_bd_ram_mem3_reg[152][24]/P0001 , \wishbone_bd_ram_mem3_reg[152][25]/P0001 , \wishbone_bd_ram_mem3_reg[152][26]/P0001 , \wishbone_bd_ram_mem3_reg[152][27]/P0001 , \wishbone_bd_ram_mem3_reg[152][28]/P0001 , \wishbone_bd_ram_mem3_reg[152][29]/P0001 , \wishbone_bd_ram_mem3_reg[152][30]/P0001 , \wishbone_bd_ram_mem3_reg[152][31]/P0001 , \wishbone_bd_ram_mem3_reg[153][24]/P0001 , \wishbone_bd_ram_mem3_reg[153][25]/P0001 , \wishbone_bd_ram_mem3_reg[153][26]/P0001 , \wishbone_bd_ram_mem3_reg[153][27]/P0001 , \wishbone_bd_ram_mem3_reg[153][28]/P0001 , \wishbone_bd_ram_mem3_reg[153][29]/P0001 , \wishbone_bd_ram_mem3_reg[153][30]/P0001 , \wishbone_bd_ram_mem3_reg[153][31]/P0001 , \wishbone_bd_ram_mem3_reg[154][24]/P0001 , \wishbone_bd_ram_mem3_reg[154][25]/P0001 , \wishbone_bd_ram_mem3_reg[154][26]/P0001 , \wishbone_bd_ram_mem3_reg[154][27]/P0001 , \wishbone_bd_ram_mem3_reg[154][28]/P0001 , \wishbone_bd_ram_mem3_reg[154][29]/P0001 , \wishbone_bd_ram_mem3_reg[154][30]/P0001 , \wishbone_bd_ram_mem3_reg[154][31]/P0001 , \wishbone_bd_ram_mem3_reg[155][24]/P0001 , \wishbone_bd_ram_mem3_reg[155][25]/P0001 , \wishbone_bd_ram_mem3_reg[155][26]/P0001 , \wishbone_bd_ram_mem3_reg[155][27]/P0001 , \wishbone_bd_ram_mem3_reg[155][28]/P0001 , \wishbone_bd_ram_mem3_reg[155][29]/P0001 , \wishbone_bd_ram_mem3_reg[155][30]/P0001 , \wishbone_bd_ram_mem3_reg[155][31]/P0001 , \wishbone_bd_ram_mem3_reg[156][24]/P0001 , \wishbone_bd_ram_mem3_reg[156][25]/P0001 , \wishbone_bd_ram_mem3_reg[156][26]/P0001 , \wishbone_bd_ram_mem3_reg[156][27]/P0001 , \wishbone_bd_ram_mem3_reg[156][28]/P0001 , \wishbone_bd_ram_mem3_reg[156][29]/P0001 , \wishbone_bd_ram_mem3_reg[156][30]/P0001 , \wishbone_bd_ram_mem3_reg[156][31]/P0001 , \wishbone_bd_ram_mem3_reg[157][24]/P0001 , \wishbone_bd_ram_mem3_reg[157][25]/P0001 , \wishbone_bd_ram_mem3_reg[157][26]/P0001 , \wishbone_bd_ram_mem3_reg[157][27]/P0001 , \wishbone_bd_ram_mem3_reg[157][28]/P0001 , \wishbone_bd_ram_mem3_reg[157][29]/P0001 , \wishbone_bd_ram_mem3_reg[157][30]/P0001 , \wishbone_bd_ram_mem3_reg[157][31]/P0001 , \wishbone_bd_ram_mem3_reg[158][24]/P0001 , \wishbone_bd_ram_mem3_reg[158][25]/P0001 , \wishbone_bd_ram_mem3_reg[158][26]/P0001 , \wishbone_bd_ram_mem3_reg[158][27]/P0001 , \wishbone_bd_ram_mem3_reg[158][28]/P0001 , \wishbone_bd_ram_mem3_reg[158][29]/P0001 , \wishbone_bd_ram_mem3_reg[158][30]/P0001 , \wishbone_bd_ram_mem3_reg[158][31]/P0001 , \wishbone_bd_ram_mem3_reg[159][24]/P0001 , \wishbone_bd_ram_mem3_reg[159][25]/P0001 , \wishbone_bd_ram_mem3_reg[159][26]/P0001 , \wishbone_bd_ram_mem3_reg[159][27]/P0001 , \wishbone_bd_ram_mem3_reg[159][28]/P0001 , \wishbone_bd_ram_mem3_reg[159][29]/P0001 , \wishbone_bd_ram_mem3_reg[159][30]/P0001 , \wishbone_bd_ram_mem3_reg[159][31]/P0001 , \wishbone_bd_ram_mem3_reg[15][24]/P0001 , \wishbone_bd_ram_mem3_reg[15][25]/P0001 , \wishbone_bd_ram_mem3_reg[15][26]/P0001 , \wishbone_bd_ram_mem3_reg[15][27]/P0001 , \wishbone_bd_ram_mem3_reg[15][28]/P0001 , \wishbone_bd_ram_mem3_reg[15][29]/P0001 , \wishbone_bd_ram_mem3_reg[15][30]/P0001 , \wishbone_bd_ram_mem3_reg[15][31]/P0001 , \wishbone_bd_ram_mem3_reg[160][24]/P0001 , \wishbone_bd_ram_mem3_reg[160][25]/P0001 , \wishbone_bd_ram_mem3_reg[160][26]/P0001 , \wishbone_bd_ram_mem3_reg[160][27]/P0001 , \wishbone_bd_ram_mem3_reg[160][28]/P0001 , \wishbone_bd_ram_mem3_reg[160][29]/P0001 , \wishbone_bd_ram_mem3_reg[160][30]/P0001 , \wishbone_bd_ram_mem3_reg[160][31]/P0001 , \wishbone_bd_ram_mem3_reg[161][24]/P0001 , \wishbone_bd_ram_mem3_reg[161][25]/P0001 , \wishbone_bd_ram_mem3_reg[161][26]/P0001 , \wishbone_bd_ram_mem3_reg[161][27]/P0001 , \wishbone_bd_ram_mem3_reg[161][28]/P0001 , \wishbone_bd_ram_mem3_reg[161][29]/P0001 , \wishbone_bd_ram_mem3_reg[161][30]/P0001 , \wishbone_bd_ram_mem3_reg[161][31]/P0001 , \wishbone_bd_ram_mem3_reg[162][24]/P0001 , \wishbone_bd_ram_mem3_reg[162][25]/P0001 , \wishbone_bd_ram_mem3_reg[162][26]/P0001 , \wishbone_bd_ram_mem3_reg[162][27]/P0001 , \wishbone_bd_ram_mem3_reg[162][28]/P0001 , \wishbone_bd_ram_mem3_reg[162][29]/P0001 , \wishbone_bd_ram_mem3_reg[162][30]/P0001 , \wishbone_bd_ram_mem3_reg[162][31]/P0001 , \wishbone_bd_ram_mem3_reg[163][24]/P0001 , \wishbone_bd_ram_mem3_reg[163][25]/P0001 , \wishbone_bd_ram_mem3_reg[163][26]/P0001 , \wishbone_bd_ram_mem3_reg[163][27]/P0001 , \wishbone_bd_ram_mem3_reg[163][28]/P0001 , \wishbone_bd_ram_mem3_reg[163][29]/P0001 , \wishbone_bd_ram_mem3_reg[163][30]/P0001 , \wishbone_bd_ram_mem3_reg[163][31]/P0001 , \wishbone_bd_ram_mem3_reg[164][24]/P0001 , \wishbone_bd_ram_mem3_reg[164][25]/P0001 , \wishbone_bd_ram_mem3_reg[164][26]/P0001 , \wishbone_bd_ram_mem3_reg[164][27]/P0001 , \wishbone_bd_ram_mem3_reg[164][28]/P0001 , \wishbone_bd_ram_mem3_reg[164][29]/P0001 , \wishbone_bd_ram_mem3_reg[164][30]/P0001 , \wishbone_bd_ram_mem3_reg[164][31]/P0001 , \wishbone_bd_ram_mem3_reg[165][24]/P0001 , \wishbone_bd_ram_mem3_reg[165][25]/P0001 , \wishbone_bd_ram_mem3_reg[165][26]/P0001 , \wishbone_bd_ram_mem3_reg[165][27]/P0001 , \wishbone_bd_ram_mem3_reg[165][28]/P0001 , \wishbone_bd_ram_mem3_reg[165][29]/P0001 , \wishbone_bd_ram_mem3_reg[165][30]/P0001 , \wishbone_bd_ram_mem3_reg[165][31]/P0001 , \wishbone_bd_ram_mem3_reg[166][24]/P0001 , \wishbone_bd_ram_mem3_reg[166][25]/P0001 , \wishbone_bd_ram_mem3_reg[166][26]/P0001 , \wishbone_bd_ram_mem3_reg[166][27]/P0001 , \wishbone_bd_ram_mem3_reg[166][28]/P0001 , \wishbone_bd_ram_mem3_reg[166][29]/P0001 , \wishbone_bd_ram_mem3_reg[166][30]/P0001 , \wishbone_bd_ram_mem3_reg[166][31]/P0001 , \wishbone_bd_ram_mem3_reg[167][24]/P0001 , \wishbone_bd_ram_mem3_reg[167][25]/P0001 , \wishbone_bd_ram_mem3_reg[167][26]/P0001 , \wishbone_bd_ram_mem3_reg[167][27]/P0001 , \wishbone_bd_ram_mem3_reg[167][28]/P0001 , \wishbone_bd_ram_mem3_reg[167][29]/P0001 , \wishbone_bd_ram_mem3_reg[167][30]/P0001 , \wishbone_bd_ram_mem3_reg[167][31]/P0001 , \wishbone_bd_ram_mem3_reg[168][24]/P0001 , \wishbone_bd_ram_mem3_reg[168][25]/P0001 , \wishbone_bd_ram_mem3_reg[168][26]/P0001 , \wishbone_bd_ram_mem3_reg[168][27]/P0001 , \wishbone_bd_ram_mem3_reg[168][28]/P0001 , \wishbone_bd_ram_mem3_reg[168][29]/P0001 , \wishbone_bd_ram_mem3_reg[168][30]/P0001 , \wishbone_bd_ram_mem3_reg[168][31]/P0001 , \wishbone_bd_ram_mem3_reg[169][24]/P0001 , \wishbone_bd_ram_mem3_reg[169][25]/P0001 , \wishbone_bd_ram_mem3_reg[169][26]/P0001 , \wishbone_bd_ram_mem3_reg[169][27]/P0001 , \wishbone_bd_ram_mem3_reg[169][28]/P0001 , \wishbone_bd_ram_mem3_reg[169][29]/P0001 , \wishbone_bd_ram_mem3_reg[169][30]/P0001 , \wishbone_bd_ram_mem3_reg[169][31]/P0001 , \wishbone_bd_ram_mem3_reg[16][24]/P0001 , \wishbone_bd_ram_mem3_reg[16][25]/P0001 , \wishbone_bd_ram_mem3_reg[16][26]/P0001 , \wishbone_bd_ram_mem3_reg[16][27]/P0001 , \wishbone_bd_ram_mem3_reg[16][28]/P0001 , \wishbone_bd_ram_mem3_reg[16][29]/P0001 , \wishbone_bd_ram_mem3_reg[16][30]/P0001 , \wishbone_bd_ram_mem3_reg[16][31]/P0001 , \wishbone_bd_ram_mem3_reg[170][24]/P0001 , \wishbone_bd_ram_mem3_reg[170][25]/P0001 , \wishbone_bd_ram_mem3_reg[170][26]/P0001 , \wishbone_bd_ram_mem3_reg[170][27]/P0001 , \wishbone_bd_ram_mem3_reg[170][28]/P0001 , \wishbone_bd_ram_mem3_reg[170][29]/P0001 , \wishbone_bd_ram_mem3_reg[170][30]/P0001 , \wishbone_bd_ram_mem3_reg[170][31]/P0001 , \wishbone_bd_ram_mem3_reg[171][24]/P0001 , \wishbone_bd_ram_mem3_reg[171][25]/P0001 , \wishbone_bd_ram_mem3_reg[171][26]/P0001 , \wishbone_bd_ram_mem3_reg[171][27]/P0001 , \wishbone_bd_ram_mem3_reg[171][28]/P0001 , \wishbone_bd_ram_mem3_reg[171][29]/P0001 , \wishbone_bd_ram_mem3_reg[171][30]/P0001 , \wishbone_bd_ram_mem3_reg[171][31]/P0001 , \wishbone_bd_ram_mem3_reg[172][24]/P0001 , \wishbone_bd_ram_mem3_reg[172][25]/P0001 , \wishbone_bd_ram_mem3_reg[172][26]/P0001 , \wishbone_bd_ram_mem3_reg[172][27]/P0001 , \wishbone_bd_ram_mem3_reg[172][28]/P0001 , \wishbone_bd_ram_mem3_reg[172][29]/P0001 , \wishbone_bd_ram_mem3_reg[172][30]/P0001 , \wishbone_bd_ram_mem3_reg[172][31]/P0001 , \wishbone_bd_ram_mem3_reg[173][24]/P0001 , \wishbone_bd_ram_mem3_reg[173][25]/P0001 , \wishbone_bd_ram_mem3_reg[173][26]/P0001 , \wishbone_bd_ram_mem3_reg[173][27]/P0001 , \wishbone_bd_ram_mem3_reg[173][28]/P0001 , \wishbone_bd_ram_mem3_reg[173][29]/P0001 , \wishbone_bd_ram_mem3_reg[173][30]/P0001 , \wishbone_bd_ram_mem3_reg[173][31]/P0001 , \wishbone_bd_ram_mem3_reg[174][24]/P0001 , \wishbone_bd_ram_mem3_reg[174][25]/P0001 , \wishbone_bd_ram_mem3_reg[174][26]/P0001 , \wishbone_bd_ram_mem3_reg[174][27]/P0001 , \wishbone_bd_ram_mem3_reg[174][28]/P0001 , \wishbone_bd_ram_mem3_reg[174][29]/P0001 , \wishbone_bd_ram_mem3_reg[174][30]/P0001 , \wishbone_bd_ram_mem3_reg[174][31]/P0001 , \wishbone_bd_ram_mem3_reg[175][24]/P0001 , \wishbone_bd_ram_mem3_reg[175][25]/P0001 , \wishbone_bd_ram_mem3_reg[175][26]/P0001 , \wishbone_bd_ram_mem3_reg[175][27]/P0001 , \wishbone_bd_ram_mem3_reg[175][28]/P0001 , \wishbone_bd_ram_mem3_reg[175][29]/P0001 , \wishbone_bd_ram_mem3_reg[175][30]/P0001 , \wishbone_bd_ram_mem3_reg[175][31]/P0001 , \wishbone_bd_ram_mem3_reg[176][24]/P0001 , \wishbone_bd_ram_mem3_reg[176][25]/P0001 , \wishbone_bd_ram_mem3_reg[176][26]/P0001 , \wishbone_bd_ram_mem3_reg[176][27]/P0001 , \wishbone_bd_ram_mem3_reg[176][28]/P0001 , \wishbone_bd_ram_mem3_reg[176][29]/P0001 , \wishbone_bd_ram_mem3_reg[176][30]/P0001 , \wishbone_bd_ram_mem3_reg[176][31]/P0001 , \wishbone_bd_ram_mem3_reg[177][24]/P0001 , \wishbone_bd_ram_mem3_reg[177][25]/P0001 , \wishbone_bd_ram_mem3_reg[177][26]/P0001 , \wishbone_bd_ram_mem3_reg[177][27]/P0001 , \wishbone_bd_ram_mem3_reg[177][28]/P0001 , \wishbone_bd_ram_mem3_reg[177][29]/P0001 , \wishbone_bd_ram_mem3_reg[177][30]/P0001 , \wishbone_bd_ram_mem3_reg[177][31]/P0001 , \wishbone_bd_ram_mem3_reg[178][24]/P0001 , \wishbone_bd_ram_mem3_reg[178][25]/P0001 , \wishbone_bd_ram_mem3_reg[178][26]/P0001 , \wishbone_bd_ram_mem3_reg[178][27]/P0001 , \wishbone_bd_ram_mem3_reg[178][28]/P0001 , \wishbone_bd_ram_mem3_reg[178][29]/P0001 , \wishbone_bd_ram_mem3_reg[178][30]/P0001 , \wishbone_bd_ram_mem3_reg[178][31]/P0001 , \wishbone_bd_ram_mem3_reg[179][24]/P0001 , \wishbone_bd_ram_mem3_reg[179][25]/P0001 , \wishbone_bd_ram_mem3_reg[179][26]/P0001 , \wishbone_bd_ram_mem3_reg[179][27]/P0001 , \wishbone_bd_ram_mem3_reg[179][28]/P0001 , \wishbone_bd_ram_mem3_reg[179][29]/P0001 , \wishbone_bd_ram_mem3_reg[179][30]/P0001 , \wishbone_bd_ram_mem3_reg[179][31]/P0001 , \wishbone_bd_ram_mem3_reg[17][24]/P0001 , \wishbone_bd_ram_mem3_reg[17][25]/P0001 , \wishbone_bd_ram_mem3_reg[17][26]/P0001 , \wishbone_bd_ram_mem3_reg[17][27]/P0001 , \wishbone_bd_ram_mem3_reg[17][28]/P0001 , \wishbone_bd_ram_mem3_reg[17][29]/P0001 , \wishbone_bd_ram_mem3_reg[17][30]/P0001 , \wishbone_bd_ram_mem3_reg[17][31]/P0001 , \wishbone_bd_ram_mem3_reg[180][24]/P0001 , \wishbone_bd_ram_mem3_reg[180][25]/P0001 , \wishbone_bd_ram_mem3_reg[180][26]/P0001 , \wishbone_bd_ram_mem3_reg[180][27]/P0001 , \wishbone_bd_ram_mem3_reg[180][28]/P0001 , \wishbone_bd_ram_mem3_reg[180][29]/P0001 , \wishbone_bd_ram_mem3_reg[180][30]/P0001 , \wishbone_bd_ram_mem3_reg[180][31]/P0001 , \wishbone_bd_ram_mem3_reg[181][24]/P0001 , \wishbone_bd_ram_mem3_reg[181][25]/P0001 , \wishbone_bd_ram_mem3_reg[181][26]/P0001 , \wishbone_bd_ram_mem3_reg[181][27]/P0001 , \wishbone_bd_ram_mem3_reg[181][28]/P0001 , \wishbone_bd_ram_mem3_reg[181][29]/P0001 , \wishbone_bd_ram_mem3_reg[181][30]/P0001 , \wishbone_bd_ram_mem3_reg[181][31]/P0001 , \wishbone_bd_ram_mem3_reg[182][24]/P0001 , \wishbone_bd_ram_mem3_reg[182][25]/P0001 , \wishbone_bd_ram_mem3_reg[182][26]/P0001 , \wishbone_bd_ram_mem3_reg[182][27]/P0001 , \wishbone_bd_ram_mem3_reg[182][28]/P0001 , \wishbone_bd_ram_mem3_reg[182][29]/P0001 , \wishbone_bd_ram_mem3_reg[182][30]/P0001 , \wishbone_bd_ram_mem3_reg[182][31]/P0001 , \wishbone_bd_ram_mem3_reg[183][24]/P0001 , \wishbone_bd_ram_mem3_reg[183][25]/P0001 , \wishbone_bd_ram_mem3_reg[183][26]/P0001 , \wishbone_bd_ram_mem3_reg[183][27]/P0001 , \wishbone_bd_ram_mem3_reg[183][28]/P0001 , \wishbone_bd_ram_mem3_reg[183][29]/P0001 , \wishbone_bd_ram_mem3_reg[183][30]/P0001 , \wishbone_bd_ram_mem3_reg[183][31]/P0001 , \wishbone_bd_ram_mem3_reg[184][24]/P0001 , \wishbone_bd_ram_mem3_reg[184][25]/P0001 , \wishbone_bd_ram_mem3_reg[184][26]/P0001 , \wishbone_bd_ram_mem3_reg[184][27]/P0001 , \wishbone_bd_ram_mem3_reg[184][28]/P0001 , \wishbone_bd_ram_mem3_reg[184][29]/P0001 , \wishbone_bd_ram_mem3_reg[184][30]/P0001 , \wishbone_bd_ram_mem3_reg[184][31]/P0001 , \wishbone_bd_ram_mem3_reg[185][24]/P0001 , \wishbone_bd_ram_mem3_reg[185][25]/P0001 , \wishbone_bd_ram_mem3_reg[185][26]/P0001 , \wishbone_bd_ram_mem3_reg[185][27]/P0001 , \wishbone_bd_ram_mem3_reg[185][28]/P0001 , \wishbone_bd_ram_mem3_reg[185][29]/P0001 , \wishbone_bd_ram_mem3_reg[185][30]/P0001 , \wishbone_bd_ram_mem3_reg[185][31]/P0001 , \wishbone_bd_ram_mem3_reg[186][24]/P0001 , \wishbone_bd_ram_mem3_reg[186][25]/P0001 , \wishbone_bd_ram_mem3_reg[186][26]/P0001 , \wishbone_bd_ram_mem3_reg[186][27]/P0001 , \wishbone_bd_ram_mem3_reg[186][28]/P0001 , \wishbone_bd_ram_mem3_reg[186][29]/P0001 , \wishbone_bd_ram_mem3_reg[186][30]/P0001 , \wishbone_bd_ram_mem3_reg[186][31]/P0001 , \wishbone_bd_ram_mem3_reg[187][24]/P0001 , \wishbone_bd_ram_mem3_reg[187][25]/P0001 , \wishbone_bd_ram_mem3_reg[187][26]/P0001 , \wishbone_bd_ram_mem3_reg[187][27]/P0001 , \wishbone_bd_ram_mem3_reg[187][28]/P0001 , \wishbone_bd_ram_mem3_reg[187][29]/P0001 , \wishbone_bd_ram_mem3_reg[187][30]/P0001 , \wishbone_bd_ram_mem3_reg[187][31]/P0001 , \wishbone_bd_ram_mem3_reg[188][24]/P0001 , \wishbone_bd_ram_mem3_reg[188][25]/P0001 , \wishbone_bd_ram_mem3_reg[188][26]/P0001 , \wishbone_bd_ram_mem3_reg[188][27]/P0001 , \wishbone_bd_ram_mem3_reg[188][28]/P0001 , \wishbone_bd_ram_mem3_reg[188][29]/P0001 , \wishbone_bd_ram_mem3_reg[188][30]/P0001 , \wishbone_bd_ram_mem3_reg[188][31]/P0001 , \wishbone_bd_ram_mem3_reg[189][24]/P0001 , \wishbone_bd_ram_mem3_reg[189][25]/P0001 , \wishbone_bd_ram_mem3_reg[189][26]/P0001 , \wishbone_bd_ram_mem3_reg[189][27]/P0001 , \wishbone_bd_ram_mem3_reg[189][28]/P0001 , \wishbone_bd_ram_mem3_reg[189][29]/P0001 , \wishbone_bd_ram_mem3_reg[189][30]/P0001 , \wishbone_bd_ram_mem3_reg[189][31]/P0001 , \wishbone_bd_ram_mem3_reg[18][24]/P0001 , \wishbone_bd_ram_mem3_reg[18][25]/P0001 , \wishbone_bd_ram_mem3_reg[18][26]/P0001 , \wishbone_bd_ram_mem3_reg[18][27]/P0001 , \wishbone_bd_ram_mem3_reg[18][28]/P0001 , \wishbone_bd_ram_mem3_reg[18][29]/P0001 , \wishbone_bd_ram_mem3_reg[18][30]/P0001 , \wishbone_bd_ram_mem3_reg[18][31]/P0001 , \wishbone_bd_ram_mem3_reg[190][24]/P0001 , \wishbone_bd_ram_mem3_reg[190][25]/P0001 , \wishbone_bd_ram_mem3_reg[190][26]/P0001 , \wishbone_bd_ram_mem3_reg[190][27]/P0001 , \wishbone_bd_ram_mem3_reg[190][28]/P0001 , \wishbone_bd_ram_mem3_reg[190][29]/P0001 , \wishbone_bd_ram_mem3_reg[190][30]/P0001 , \wishbone_bd_ram_mem3_reg[190][31]/P0001 , \wishbone_bd_ram_mem3_reg[191][24]/P0001 , \wishbone_bd_ram_mem3_reg[191][25]/P0001 , \wishbone_bd_ram_mem3_reg[191][26]/P0001 , \wishbone_bd_ram_mem3_reg[191][27]/P0001 , \wishbone_bd_ram_mem3_reg[191][28]/P0001 , \wishbone_bd_ram_mem3_reg[191][29]/P0001 , \wishbone_bd_ram_mem3_reg[191][30]/P0001 , \wishbone_bd_ram_mem3_reg[191][31]/P0001 , \wishbone_bd_ram_mem3_reg[192][24]/P0001 , \wishbone_bd_ram_mem3_reg[192][25]/P0001 , \wishbone_bd_ram_mem3_reg[192][26]/P0001 , \wishbone_bd_ram_mem3_reg[192][27]/P0001 , \wishbone_bd_ram_mem3_reg[192][28]/P0001 , \wishbone_bd_ram_mem3_reg[192][29]/P0001 , \wishbone_bd_ram_mem3_reg[192][30]/P0001 , \wishbone_bd_ram_mem3_reg[192][31]/P0001 , \wishbone_bd_ram_mem3_reg[193][24]/P0001 , \wishbone_bd_ram_mem3_reg[193][25]/P0001 , \wishbone_bd_ram_mem3_reg[193][26]/P0001 , \wishbone_bd_ram_mem3_reg[193][27]/P0001 , \wishbone_bd_ram_mem3_reg[193][28]/P0001 , \wishbone_bd_ram_mem3_reg[193][29]/P0001 , \wishbone_bd_ram_mem3_reg[193][30]/P0001 , \wishbone_bd_ram_mem3_reg[193][31]/P0001 , \wishbone_bd_ram_mem3_reg[194][24]/P0001 , \wishbone_bd_ram_mem3_reg[194][25]/P0001 , \wishbone_bd_ram_mem3_reg[194][26]/P0001 , \wishbone_bd_ram_mem3_reg[194][27]/P0001 , \wishbone_bd_ram_mem3_reg[194][28]/P0001 , \wishbone_bd_ram_mem3_reg[194][29]/P0001 , \wishbone_bd_ram_mem3_reg[194][30]/P0001 , \wishbone_bd_ram_mem3_reg[194][31]/P0001 , \wishbone_bd_ram_mem3_reg[195][24]/P0001 , \wishbone_bd_ram_mem3_reg[195][25]/P0001 , \wishbone_bd_ram_mem3_reg[195][26]/P0001 , \wishbone_bd_ram_mem3_reg[195][27]/P0001 , \wishbone_bd_ram_mem3_reg[195][28]/P0001 , \wishbone_bd_ram_mem3_reg[195][29]/P0001 , \wishbone_bd_ram_mem3_reg[195][30]/P0001 , \wishbone_bd_ram_mem3_reg[195][31]/P0001 , \wishbone_bd_ram_mem3_reg[196][24]/P0001 , \wishbone_bd_ram_mem3_reg[196][25]/P0001 , \wishbone_bd_ram_mem3_reg[196][26]/P0001 , \wishbone_bd_ram_mem3_reg[196][27]/P0001 , \wishbone_bd_ram_mem3_reg[196][28]/P0001 , \wishbone_bd_ram_mem3_reg[196][29]/P0001 , \wishbone_bd_ram_mem3_reg[196][30]/P0001 , \wishbone_bd_ram_mem3_reg[196][31]/P0001 , \wishbone_bd_ram_mem3_reg[197][24]/P0001 , \wishbone_bd_ram_mem3_reg[197][25]/P0001 , \wishbone_bd_ram_mem3_reg[197][26]/P0001 , \wishbone_bd_ram_mem3_reg[197][27]/P0001 , \wishbone_bd_ram_mem3_reg[197][28]/P0001 , \wishbone_bd_ram_mem3_reg[197][29]/P0001 , \wishbone_bd_ram_mem3_reg[197][30]/P0001 , \wishbone_bd_ram_mem3_reg[197][31]/P0001 , \wishbone_bd_ram_mem3_reg[198][24]/P0001 , \wishbone_bd_ram_mem3_reg[198][25]/P0001 , \wishbone_bd_ram_mem3_reg[198][26]/P0001 , \wishbone_bd_ram_mem3_reg[198][27]/P0001 , \wishbone_bd_ram_mem3_reg[198][28]/P0001 , \wishbone_bd_ram_mem3_reg[198][29]/P0001 , \wishbone_bd_ram_mem3_reg[198][30]/P0001 , \wishbone_bd_ram_mem3_reg[198][31]/P0001 , \wishbone_bd_ram_mem3_reg[199][24]/P0001 , \wishbone_bd_ram_mem3_reg[199][25]/P0001 , \wishbone_bd_ram_mem3_reg[199][26]/P0001 , \wishbone_bd_ram_mem3_reg[199][27]/P0001 , \wishbone_bd_ram_mem3_reg[199][28]/P0001 , \wishbone_bd_ram_mem3_reg[199][29]/P0001 , \wishbone_bd_ram_mem3_reg[199][30]/P0001 , \wishbone_bd_ram_mem3_reg[199][31]/P0001 , \wishbone_bd_ram_mem3_reg[19][24]/P0001 , \wishbone_bd_ram_mem3_reg[19][25]/P0001 , \wishbone_bd_ram_mem3_reg[19][26]/P0001 , \wishbone_bd_ram_mem3_reg[19][27]/P0001 , \wishbone_bd_ram_mem3_reg[19][28]/P0001 , \wishbone_bd_ram_mem3_reg[19][29]/P0001 , \wishbone_bd_ram_mem3_reg[19][30]/P0001 , \wishbone_bd_ram_mem3_reg[19][31]/P0001 , \wishbone_bd_ram_mem3_reg[1][24]/P0001 , \wishbone_bd_ram_mem3_reg[1][25]/P0001 , \wishbone_bd_ram_mem3_reg[1][26]/P0001 , \wishbone_bd_ram_mem3_reg[1][27]/P0001 , \wishbone_bd_ram_mem3_reg[1][28]/P0001 , \wishbone_bd_ram_mem3_reg[1][29]/P0001 , \wishbone_bd_ram_mem3_reg[1][30]/P0001 , \wishbone_bd_ram_mem3_reg[1][31]/P0001 , \wishbone_bd_ram_mem3_reg[200][24]/P0001 , \wishbone_bd_ram_mem3_reg[200][25]/P0001 , \wishbone_bd_ram_mem3_reg[200][26]/P0001 , \wishbone_bd_ram_mem3_reg[200][27]/P0001 , \wishbone_bd_ram_mem3_reg[200][28]/P0001 , \wishbone_bd_ram_mem3_reg[200][29]/P0001 , \wishbone_bd_ram_mem3_reg[200][30]/P0001 , \wishbone_bd_ram_mem3_reg[200][31]/P0001 , \wishbone_bd_ram_mem3_reg[201][24]/P0001 , \wishbone_bd_ram_mem3_reg[201][25]/P0001 , \wishbone_bd_ram_mem3_reg[201][26]/P0001 , \wishbone_bd_ram_mem3_reg[201][27]/P0001 , \wishbone_bd_ram_mem3_reg[201][28]/P0001 , \wishbone_bd_ram_mem3_reg[201][29]/P0001 , \wishbone_bd_ram_mem3_reg[201][30]/P0001 , \wishbone_bd_ram_mem3_reg[201][31]/P0001 , \wishbone_bd_ram_mem3_reg[202][24]/P0001 , \wishbone_bd_ram_mem3_reg[202][25]/P0001 , \wishbone_bd_ram_mem3_reg[202][26]/P0001 , \wishbone_bd_ram_mem3_reg[202][27]/P0001 , \wishbone_bd_ram_mem3_reg[202][28]/P0001 , \wishbone_bd_ram_mem3_reg[202][29]/P0001 , \wishbone_bd_ram_mem3_reg[202][30]/P0001 , \wishbone_bd_ram_mem3_reg[202][31]/P0001 , \wishbone_bd_ram_mem3_reg[203][24]/P0001 , \wishbone_bd_ram_mem3_reg[203][25]/P0001 , \wishbone_bd_ram_mem3_reg[203][26]/P0001 , \wishbone_bd_ram_mem3_reg[203][27]/P0001 , \wishbone_bd_ram_mem3_reg[203][28]/P0001 , \wishbone_bd_ram_mem3_reg[203][29]/P0001 , \wishbone_bd_ram_mem3_reg[203][30]/P0001 , \wishbone_bd_ram_mem3_reg[203][31]/P0001 , \wishbone_bd_ram_mem3_reg[204][24]/P0001 , \wishbone_bd_ram_mem3_reg[204][25]/P0001 , \wishbone_bd_ram_mem3_reg[204][26]/P0001 , \wishbone_bd_ram_mem3_reg[204][27]/P0001 , \wishbone_bd_ram_mem3_reg[204][28]/P0001 , \wishbone_bd_ram_mem3_reg[204][29]/P0001 , \wishbone_bd_ram_mem3_reg[204][30]/P0001 , \wishbone_bd_ram_mem3_reg[204][31]/P0001 , \wishbone_bd_ram_mem3_reg[205][24]/P0001 , \wishbone_bd_ram_mem3_reg[205][25]/P0001 , \wishbone_bd_ram_mem3_reg[205][26]/P0001 , \wishbone_bd_ram_mem3_reg[205][27]/P0001 , \wishbone_bd_ram_mem3_reg[205][28]/P0001 , \wishbone_bd_ram_mem3_reg[205][29]/P0001 , \wishbone_bd_ram_mem3_reg[205][30]/P0001 , \wishbone_bd_ram_mem3_reg[205][31]/P0001 , \wishbone_bd_ram_mem3_reg[206][24]/P0001 , \wishbone_bd_ram_mem3_reg[206][25]/P0001 , \wishbone_bd_ram_mem3_reg[206][26]/P0001 , \wishbone_bd_ram_mem3_reg[206][27]/P0001 , \wishbone_bd_ram_mem3_reg[206][28]/P0001 , \wishbone_bd_ram_mem3_reg[206][29]/P0001 , \wishbone_bd_ram_mem3_reg[206][30]/P0001 , \wishbone_bd_ram_mem3_reg[206][31]/P0001 , \wishbone_bd_ram_mem3_reg[207][24]/P0001 , \wishbone_bd_ram_mem3_reg[207][25]/P0001 , \wishbone_bd_ram_mem3_reg[207][26]/P0001 , \wishbone_bd_ram_mem3_reg[207][27]/P0001 , \wishbone_bd_ram_mem3_reg[207][28]/P0001 , \wishbone_bd_ram_mem3_reg[207][29]/P0001 , \wishbone_bd_ram_mem3_reg[207][30]/P0001 , \wishbone_bd_ram_mem3_reg[207][31]/P0001 , \wishbone_bd_ram_mem3_reg[208][24]/P0001 , \wishbone_bd_ram_mem3_reg[208][25]/P0001 , \wishbone_bd_ram_mem3_reg[208][26]/P0001 , \wishbone_bd_ram_mem3_reg[208][27]/P0001 , \wishbone_bd_ram_mem3_reg[208][28]/P0001 , \wishbone_bd_ram_mem3_reg[208][29]/P0001 , \wishbone_bd_ram_mem3_reg[208][30]/P0001 , \wishbone_bd_ram_mem3_reg[208][31]/P0001 , \wishbone_bd_ram_mem3_reg[209][24]/P0001 , \wishbone_bd_ram_mem3_reg[209][25]/P0001 , \wishbone_bd_ram_mem3_reg[209][26]/P0001 , \wishbone_bd_ram_mem3_reg[209][27]/P0001 , \wishbone_bd_ram_mem3_reg[209][28]/P0001 , \wishbone_bd_ram_mem3_reg[209][29]/P0001 , \wishbone_bd_ram_mem3_reg[209][30]/P0001 , \wishbone_bd_ram_mem3_reg[209][31]/P0001 , \wishbone_bd_ram_mem3_reg[20][24]/P0001 , \wishbone_bd_ram_mem3_reg[20][25]/P0001 , \wishbone_bd_ram_mem3_reg[20][26]/P0001 , \wishbone_bd_ram_mem3_reg[20][27]/P0001 , \wishbone_bd_ram_mem3_reg[20][28]/P0001 , \wishbone_bd_ram_mem3_reg[20][29]/P0001 , \wishbone_bd_ram_mem3_reg[20][30]/P0001 , \wishbone_bd_ram_mem3_reg[20][31]/P0001 , \wishbone_bd_ram_mem3_reg[210][24]/P0001 , \wishbone_bd_ram_mem3_reg[210][25]/P0001 , \wishbone_bd_ram_mem3_reg[210][26]/P0001 , \wishbone_bd_ram_mem3_reg[210][27]/P0001 , \wishbone_bd_ram_mem3_reg[210][28]/P0001 , \wishbone_bd_ram_mem3_reg[210][29]/P0001 , \wishbone_bd_ram_mem3_reg[210][30]/P0001 , \wishbone_bd_ram_mem3_reg[210][31]/P0001 , \wishbone_bd_ram_mem3_reg[211][24]/P0001 , \wishbone_bd_ram_mem3_reg[211][25]/P0001 , \wishbone_bd_ram_mem3_reg[211][26]/P0001 , \wishbone_bd_ram_mem3_reg[211][27]/P0001 , \wishbone_bd_ram_mem3_reg[211][28]/P0001 , \wishbone_bd_ram_mem3_reg[211][29]/P0001 , \wishbone_bd_ram_mem3_reg[211][30]/P0001 , \wishbone_bd_ram_mem3_reg[211][31]/P0001 , \wishbone_bd_ram_mem3_reg[212][24]/P0001 , \wishbone_bd_ram_mem3_reg[212][25]/P0001 , \wishbone_bd_ram_mem3_reg[212][26]/P0001 , \wishbone_bd_ram_mem3_reg[212][27]/P0001 , \wishbone_bd_ram_mem3_reg[212][28]/P0001 , \wishbone_bd_ram_mem3_reg[212][29]/P0001 , \wishbone_bd_ram_mem3_reg[212][30]/P0001 , \wishbone_bd_ram_mem3_reg[212][31]/P0001 , \wishbone_bd_ram_mem3_reg[213][24]/P0001 , \wishbone_bd_ram_mem3_reg[213][25]/P0001 , \wishbone_bd_ram_mem3_reg[213][26]/P0001 , \wishbone_bd_ram_mem3_reg[213][27]/P0001 , \wishbone_bd_ram_mem3_reg[213][28]/P0001 , \wishbone_bd_ram_mem3_reg[213][29]/P0001 , \wishbone_bd_ram_mem3_reg[213][30]/P0001 , \wishbone_bd_ram_mem3_reg[213][31]/P0001 , \wishbone_bd_ram_mem3_reg[214][24]/P0001 , \wishbone_bd_ram_mem3_reg[214][25]/P0001 , \wishbone_bd_ram_mem3_reg[214][26]/P0001 , \wishbone_bd_ram_mem3_reg[214][27]/P0001 , \wishbone_bd_ram_mem3_reg[214][28]/P0001 , \wishbone_bd_ram_mem3_reg[214][29]/P0001 , \wishbone_bd_ram_mem3_reg[214][30]/P0001 , \wishbone_bd_ram_mem3_reg[214][31]/P0001 , \wishbone_bd_ram_mem3_reg[215][24]/P0001 , \wishbone_bd_ram_mem3_reg[215][25]/P0001 , \wishbone_bd_ram_mem3_reg[215][26]/P0001 , \wishbone_bd_ram_mem3_reg[215][27]/P0001 , \wishbone_bd_ram_mem3_reg[215][28]/P0001 , \wishbone_bd_ram_mem3_reg[215][29]/P0001 , \wishbone_bd_ram_mem3_reg[215][30]/P0001 , \wishbone_bd_ram_mem3_reg[215][31]/P0001 , \wishbone_bd_ram_mem3_reg[216][24]/P0001 , \wishbone_bd_ram_mem3_reg[216][25]/P0001 , \wishbone_bd_ram_mem3_reg[216][26]/P0001 , \wishbone_bd_ram_mem3_reg[216][27]/P0001 , \wishbone_bd_ram_mem3_reg[216][28]/P0001 , \wishbone_bd_ram_mem3_reg[216][29]/P0001 , \wishbone_bd_ram_mem3_reg[216][30]/P0001 , \wishbone_bd_ram_mem3_reg[216][31]/P0001 , \wishbone_bd_ram_mem3_reg[217][24]/P0001 , \wishbone_bd_ram_mem3_reg[217][25]/P0001 , \wishbone_bd_ram_mem3_reg[217][26]/P0001 , \wishbone_bd_ram_mem3_reg[217][27]/P0001 , \wishbone_bd_ram_mem3_reg[217][28]/P0001 , \wishbone_bd_ram_mem3_reg[217][29]/P0001 , \wishbone_bd_ram_mem3_reg[217][30]/P0001 , \wishbone_bd_ram_mem3_reg[217][31]/P0001 , \wishbone_bd_ram_mem3_reg[218][24]/P0001 , \wishbone_bd_ram_mem3_reg[218][25]/P0001 , \wishbone_bd_ram_mem3_reg[218][26]/P0001 , \wishbone_bd_ram_mem3_reg[218][27]/P0001 , \wishbone_bd_ram_mem3_reg[218][28]/P0001 , \wishbone_bd_ram_mem3_reg[218][29]/P0001 , \wishbone_bd_ram_mem3_reg[218][30]/P0001 , \wishbone_bd_ram_mem3_reg[218][31]/P0001 , \wishbone_bd_ram_mem3_reg[219][24]/P0001 , \wishbone_bd_ram_mem3_reg[219][25]/P0001 , \wishbone_bd_ram_mem3_reg[219][26]/P0001 , \wishbone_bd_ram_mem3_reg[219][27]/P0001 , \wishbone_bd_ram_mem3_reg[219][28]/P0001 , \wishbone_bd_ram_mem3_reg[219][29]/P0001 , \wishbone_bd_ram_mem3_reg[219][30]/P0001 , \wishbone_bd_ram_mem3_reg[219][31]/P0001 , \wishbone_bd_ram_mem3_reg[21][24]/P0001 , \wishbone_bd_ram_mem3_reg[21][25]/P0001 , \wishbone_bd_ram_mem3_reg[21][26]/P0001 , \wishbone_bd_ram_mem3_reg[21][27]/P0001 , \wishbone_bd_ram_mem3_reg[21][28]/P0001 , \wishbone_bd_ram_mem3_reg[21][29]/P0001 , \wishbone_bd_ram_mem3_reg[21][30]/P0001 , \wishbone_bd_ram_mem3_reg[21][31]/P0001 , \wishbone_bd_ram_mem3_reg[220][24]/P0001 , \wishbone_bd_ram_mem3_reg[220][25]/P0001 , \wishbone_bd_ram_mem3_reg[220][26]/P0001 , \wishbone_bd_ram_mem3_reg[220][27]/P0001 , \wishbone_bd_ram_mem3_reg[220][28]/P0001 , \wishbone_bd_ram_mem3_reg[220][29]/P0001 , \wishbone_bd_ram_mem3_reg[220][30]/P0001 , \wishbone_bd_ram_mem3_reg[220][31]/P0001 , \wishbone_bd_ram_mem3_reg[221][24]/P0001 , \wishbone_bd_ram_mem3_reg[221][25]/P0001 , \wishbone_bd_ram_mem3_reg[221][26]/P0001 , \wishbone_bd_ram_mem3_reg[221][27]/P0001 , \wishbone_bd_ram_mem3_reg[221][28]/P0001 , \wishbone_bd_ram_mem3_reg[221][29]/P0001 , \wishbone_bd_ram_mem3_reg[221][30]/P0001 , \wishbone_bd_ram_mem3_reg[221][31]/P0001 , \wishbone_bd_ram_mem3_reg[222][24]/P0001 , \wishbone_bd_ram_mem3_reg[222][25]/P0001 , \wishbone_bd_ram_mem3_reg[222][26]/P0001 , \wishbone_bd_ram_mem3_reg[222][27]/P0001 , \wishbone_bd_ram_mem3_reg[222][28]/P0001 , \wishbone_bd_ram_mem3_reg[222][29]/P0001 , \wishbone_bd_ram_mem3_reg[222][30]/P0001 , \wishbone_bd_ram_mem3_reg[222][31]/P0001 , \wishbone_bd_ram_mem3_reg[223][24]/P0001 , \wishbone_bd_ram_mem3_reg[223][25]/P0001 , \wishbone_bd_ram_mem3_reg[223][26]/P0001 , \wishbone_bd_ram_mem3_reg[223][27]/P0001 , \wishbone_bd_ram_mem3_reg[223][28]/P0001 , \wishbone_bd_ram_mem3_reg[223][29]/P0001 , \wishbone_bd_ram_mem3_reg[223][30]/P0001 , \wishbone_bd_ram_mem3_reg[223][31]/P0001 , \wishbone_bd_ram_mem3_reg[224][24]/P0001 , \wishbone_bd_ram_mem3_reg[224][25]/P0001 , \wishbone_bd_ram_mem3_reg[224][26]/P0001 , \wishbone_bd_ram_mem3_reg[224][27]/P0001 , \wishbone_bd_ram_mem3_reg[224][28]/P0001 , \wishbone_bd_ram_mem3_reg[224][29]/P0001 , \wishbone_bd_ram_mem3_reg[224][30]/P0001 , \wishbone_bd_ram_mem3_reg[224][31]/P0001 , \wishbone_bd_ram_mem3_reg[225][24]/P0001 , \wishbone_bd_ram_mem3_reg[225][25]/P0001 , \wishbone_bd_ram_mem3_reg[225][26]/P0001 , \wishbone_bd_ram_mem3_reg[225][27]/P0001 , \wishbone_bd_ram_mem3_reg[225][28]/P0001 , \wishbone_bd_ram_mem3_reg[225][29]/P0001 , \wishbone_bd_ram_mem3_reg[225][30]/P0001 , \wishbone_bd_ram_mem3_reg[225][31]/P0001 , \wishbone_bd_ram_mem3_reg[226][24]/P0001 , \wishbone_bd_ram_mem3_reg[226][25]/P0001 , \wishbone_bd_ram_mem3_reg[226][26]/P0001 , \wishbone_bd_ram_mem3_reg[226][27]/P0001 , \wishbone_bd_ram_mem3_reg[226][28]/P0001 , \wishbone_bd_ram_mem3_reg[226][29]/P0001 , \wishbone_bd_ram_mem3_reg[226][30]/P0001 , \wishbone_bd_ram_mem3_reg[226][31]/P0001 , \wishbone_bd_ram_mem3_reg[227][24]/P0001 , \wishbone_bd_ram_mem3_reg[227][25]/P0001 , \wishbone_bd_ram_mem3_reg[227][26]/P0001 , \wishbone_bd_ram_mem3_reg[227][27]/P0001 , \wishbone_bd_ram_mem3_reg[227][28]/P0001 , \wishbone_bd_ram_mem3_reg[227][29]/P0001 , \wishbone_bd_ram_mem3_reg[227][30]/P0001 , \wishbone_bd_ram_mem3_reg[227][31]/P0001 , \wishbone_bd_ram_mem3_reg[228][24]/P0001 , \wishbone_bd_ram_mem3_reg[228][25]/P0001 , \wishbone_bd_ram_mem3_reg[228][26]/P0001 , \wishbone_bd_ram_mem3_reg[228][27]/P0001 , \wishbone_bd_ram_mem3_reg[228][28]/P0001 , \wishbone_bd_ram_mem3_reg[228][29]/P0001 , \wishbone_bd_ram_mem3_reg[228][30]/P0001 , \wishbone_bd_ram_mem3_reg[228][31]/P0001 , \wishbone_bd_ram_mem3_reg[229][24]/P0001 , \wishbone_bd_ram_mem3_reg[229][25]/P0001 , \wishbone_bd_ram_mem3_reg[229][26]/P0001 , \wishbone_bd_ram_mem3_reg[229][27]/P0001 , \wishbone_bd_ram_mem3_reg[229][28]/P0001 , \wishbone_bd_ram_mem3_reg[229][29]/P0001 , \wishbone_bd_ram_mem3_reg[229][30]/P0001 , \wishbone_bd_ram_mem3_reg[229][31]/P0001 , \wishbone_bd_ram_mem3_reg[22][24]/P0001 , \wishbone_bd_ram_mem3_reg[22][25]/P0001 , \wishbone_bd_ram_mem3_reg[22][26]/P0001 , \wishbone_bd_ram_mem3_reg[22][27]/P0001 , \wishbone_bd_ram_mem3_reg[22][28]/P0001 , \wishbone_bd_ram_mem3_reg[22][29]/P0001 , \wishbone_bd_ram_mem3_reg[22][30]/P0001 , \wishbone_bd_ram_mem3_reg[22][31]/P0001 , \wishbone_bd_ram_mem3_reg[230][24]/P0001 , \wishbone_bd_ram_mem3_reg[230][25]/P0001 , \wishbone_bd_ram_mem3_reg[230][26]/P0001 , \wishbone_bd_ram_mem3_reg[230][27]/P0001 , \wishbone_bd_ram_mem3_reg[230][28]/P0001 , \wishbone_bd_ram_mem3_reg[230][29]/P0001 , \wishbone_bd_ram_mem3_reg[230][30]/P0001 , \wishbone_bd_ram_mem3_reg[230][31]/P0001 , \wishbone_bd_ram_mem3_reg[231][24]/P0001 , \wishbone_bd_ram_mem3_reg[231][25]/P0001 , \wishbone_bd_ram_mem3_reg[231][26]/P0001 , \wishbone_bd_ram_mem3_reg[231][27]/P0001 , \wishbone_bd_ram_mem3_reg[231][28]/P0001 , \wishbone_bd_ram_mem3_reg[231][29]/P0001 , \wishbone_bd_ram_mem3_reg[231][30]/P0001 , \wishbone_bd_ram_mem3_reg[231][31]/P0001 , \wishbone_bd_ram_mem3_reg[232][24]/P0001 , \wishbone_bd_ram_mem3_reg[232][25]/P0001 , \wishbone_bd_ram_mem3_reg[232][26]/P0001 , \wishbone_bd_ram_mem3_reg[232][27]/P0001 , \wishbone_bd_ram_mem3_reg[232][28]/P0001 , \wishbone_bd_ram_mem3_reg[232][29]/P0001 , \wishbone_bd_ram_mem3_reg[232][30]/P0001 , \wishbone_bd_ram_mem3_reg[232][31]/P0001 , \wishbone_bd_ram_mem3_reg[233][24]/P0001 , \wishbone_bd_ram_mem3_reg[233][25]/P0001 , \wishbone_bd_ram_mem3_reg[233][26]/P0001 , \wishbone_bd_ram_mem3_reg[233][27]/P0001 , \wishbone_bd_ram_mem3_reg[233][28]/P0001 , \wishbone_bd_ram_mem3_reg[233][29]/P0001 , \wishbone_bd_ram_mem3_reg[233][30]/P0001 , \wishbone_bd_ram_mem3_reg[233][31]/P0001 , \wishbone_bd_ram_mem3_reg[234][24]/P0001 , \wishbone_bd_ram_mem3_reg[234][25]/P0001 , \wishbone_bd_ram_mem3_reg[234][26]/P0001 , \wishbone_bd_ram_mem3_reg[234][27]/P0001 , \wishbone_bd_ram_mem3_reg[234][28]/P0001 , \wishbone_bd_ram_mem3_reg[234][29]/P0001 , \wishbone_bd_ram_mem3_reg[234][30]/P0001 , \wishbone_bd_ram_mem3_reg[234][31]/P0001 , \wishbone_bd_ram_mem3_reg[235][24]/P0001 , \wishbone_bd_ram_mem3_reg[235][25]/P0001 , \wishbone_bd_ram_mem3_reg[235][26]/P0001 , \wishbone_bd_ram_mem3_reg[235][27]/P0001 , \wishbone_bd_ram_mem3_reg[235][28]/P0001 , \wishbone_bd_ram_mem3_reg[235][29]/P0001 , \wishbone_bd_ram_mem3_reg[235][30]/P0001 , \wishbone_bd_ram_mem3_reg[235][31]/P0001 , \wishbone_bd_ram_mem3_reg[236][24]/P0001 , \wishbone_bd_ram_mem3_reg[236][25]/P0001 , \wishbone_bd_ram_mem3_reg[236][26]/P0001 , \wishbone_bd_ram_mem3_reg[236][27]/P0001 , \wishbone_bd_ram_mem3_reg[236][28]/P0001 , \wishbone_bd_ram_mem3_reg[236][29]/P0001 , \wishbone_bd_ram_mem3_reg[236][30]/P0001 , \wishbone_bd_ram_mem3_reg[236][31]/P0001 , \wishbone_bd_ram_mem3_reg[237][24]/P0001 , \wishbone_bd_ram_mem3_reg[237][25]/P0001 , \wishbone_bd_ram_mem3_reg[237][26]/P0001 , \wishbone_bd_ram_mem3_reg[237][27]/P0001 , \wishbone_bd_ram_mem3_reg[237][28]/P0001 , \wishbone_bd_ram_mem3_reg[237][29]/P0001 , \wishbone_bd_ram_mem3_reg[237][30]/P0001 , \wishbone_bd_ram_mem3_reg[237][31]/P0001 , \wishbone_bd_ram_mem3_reg[238][24]/P0001 , \wishbone_bd_ram_mem3_reg[238][25]/P0001 , \wishbone_bd_ram_mem3_reg[238][26]/P0001 , \wishbone_bd_ram_mem3_reg[238][27]/P0001 , \wishbone_bd_ram_mem3_reg[238][28]/P0001 , \wishbone_bd_ram_mem3_reg[238][29]/P0001 , \wishbone_bd_ram_mem3_reg[238][30]/P0001 , \wishbone_bd_ram_mem3_reg[238][31]/P0001 , \wishbone_bd_ram_mem3_reg[239][24]/P0001 , \wishbone_bd_ram_mem3_reg[239][25]/P0001 , \wishbone_bd_ram_mem3_reg[239][26]/P0001 , \wishbone_bd_ram_mem3_reg[239][27]/P0001 , \wishbone_bd_ram_mem3_reg[239][28]/P0001 , \wishbone_bd_ram_mem3_reg[239][29]/P0001 , \wishbone_bd_ram_mem3_reg[239][30]/P0001 , \wishbone_bd_ram_mem3_reg[239][31]/P0001 , \wishbone_bd_ram_mem3_reg[23][24]/P0001 , \wishbone_bd_ram_mem3_reg[23][25]/P0001 , \wishbone_bd_ram_mem3_reg[23][26]/P0001 , \wishbone_bd_ram_mem3_reg[23][27]/P0001 , \wishbone_bd_ram_mem3_reg[23][28]/P0001 , \wishbone_bd_ram_mem3_reg[23][29]/P0001 , \wishbone_bd_ram_mem3_reg[23][30]/P0001 , \wishbone_bd_ram_mem3_reg[23][31]/P0001 , \wishbone_bd_ram_mem3_reg[240][24]/P0001 , \wishbone_bd_ram_mem3_reg[240][25]/P0001 , \wishbone_bd_ram_mem3_reg[240][26]/P0001 , \wishbone_bd_ram_mem3_reg[240][27]/P0001 , \wishbone_bd_ram_mem3_reg[240][28]/P0001 , \wishbone_bd_ram_mem3_reg[240][29]/P0001 , \wishbone_bd_ram_mem3_reg[240][30]/P0001 , \wishbone_bd_ram_mem3_reg[240][31]/P0001 , \wishbone_bd_ram_mem3_reg[241][24]/P0001 , \wishbone_bd_ram_mem3_reg[241][25]/P0001 , \wishbone_bd_ram_mem3_reg[241][26]/P0001 , \wishbone_bd_ram_mem3_reg[241][27]/P0001 , \wishbone_bd_ram_mem3_reg[241][28]/P0001 , \wishbone_bd_ram_mem3_reg[241][29]/P0001 , \wishbone_bd_ram_mem3_reg[241][30]/P0001 , \wishbone_bd_ram_mem3_reg[241][31]/P0001 , \wishbone_bd_ram_mem3_reg[242][24]/P0001 , \wishbone_bd_ram_mem3_reg[242][25]/P0001 , \wishbone_bd_ram_mem3_reg[242][26]/P0001 , \wishbone_bd_ram_mem3_reg[242][27]/P0001 , \wishbone_bd_ram_mem3_reg[242][28]/P0001 , \wishbone_bd_ram_mem3_reg[242][29]/P0001 , \wishbone_bd_ram_mem3_reg[242][30]/P0001 , \wishbone_bd_ram_mem3_reg[242][31]/P0001 , \wishbone_bd_ram_mem3_reg[243][24]/P0001 , \wishbone_bd_ram_mem3_reg[243][25]/P0001 , \wishbone_bd_ram_mem3_reg[243][26]/P0001 , \wishbone_bd_ram_mem3_reg[243][27]/P0001 , \wishbone_bd_ram_mem3_reg[243][28]/P0001 , \wishbone_bd_ram_mem3_reg[243][29]/P0001 , \wishbone_bd_ram_mem3_reg[243][30]/P0001 , \wishbone_bd_ram_mem3_reg[243][31]/P0001 , \wishbone_bd_ram_mem3_reg[244][24]/P0001 , \wishbone_bd_ram_mem3_reg[244][25]/P0001 , \wishbone_bd_ram_mem3_reg[244][26]/P0001 , \wishbone_bd_ram_mem3_reg[244][27]/P0001 , \wishbone_bd_ram_mem3_reg[244][28]/P0001 , \wishbone_bd_ram_mem3_reg[244][29]/P0001 , \wishbone_bd_ram_mem3_reg[244][30]/P0001 , \wishbone_bd_ram_mem3_reg[244][31]/P0001 , \wishbone_bd_ram_mem3_reg[245][24]/P0001 , \wishbone_bd_ram_mem3_reg[245][25]/P0001 , \wishbone_bd_ram_mem3_reg[245][26]/P0001 , \wishbone_bd_ram_mem3_reg[245][27]/P0001 , \wishbone_bd_ram_mem3_reg[245][28]/P0001 , \wishbone_bd_ram_mem3_reg[245][29]/P0001 , \wishbone_bd_ram_mem3_reg[245][30]/P0001 , \wishbone_bd_ram_mem3_reg[245][31]/P0001 , \wishbone_bd_ram_mem3_reg[246][24]/P0001 , \wishbone_bd_ram_mem3_reg[246][25]/P0001 , \wishbone_bd_ram_mem3_reg[246][26]/P0001 , \wishbone_bd_ram_mem3_reg[246][27]/P0001 , \wishbone_bd_ram_mem3_reg[246][28]/P0001 , \wishbone_bd_ram_mem3_reg[246][29]/P0001 , \wishbone_bd_ram_mem3_reg[246][30]/P0001 , \wishbone_bd_ram_mem3_reg[246][31]/P0001 , \wishbone_bd_ram_mem3_reg[247][24]/P0001 , \wishbone_bd_ram_mem3_reg[247][25]/P0001 , \wishbone_bd_ram_mem3_reg[247][26]/P0001 , \wishbone_bd_ram_mem3_reg[247][27]/P0001 , \wishbone_bd_ram_mem3_reg[247][28]/P0001 , \wishbone_bd_ram_mem3_reg[247][29]/P0001 , \wishbone_bd_ram_mem3_reg[247][30]/P0001 , \wishbone_bd_ram_mem3_reg[247][31]/P0001 , \wishbone_bd_ram_mem3_reg[248][24]/P0001 , \wishbone_bd_ram_mem3_reg[248][25]/P0001 , \wishbone_bd_ram_mem3_reg[248][26]/P0001 , \wishbone_bd_ram_mem3_reg[248][27]/P0001 , \wishbone_bd_ram_mem3_reg[248][28]/P0001 , \wishbone_bd_ram_mem3_reg[248][29]/P0001 , \wishbone_bd_ram_mem3_reg[248][30]/P0001 , \wishbone_bd_ram_mem3_reg[248][31]/P0001 , \wishbone_bd_ram_mem3_reg[249][24]/P0001 , \wishbone_bd_ram_mem3_reg[249][25]/P0001 , \wishbone_bd_ram_mem3_reg[249][26]/P0001 , \wishbone_bd_ram_mem3_reg[249][27]/P0001 , \wishbone_bd_ram_mem3_reg[249][28]/P0001 , \wishbone_bd_ram_mem3_reg[249][29]/P0001 , \wishbone_bd_ram_mem3_reg[249][30]/P0001 , \wishbone_bd_ram_mem3_reg[249][31]/P0001 , \wishbone_bd_ram_mem3_reg[24][24]/P0001 , \wishbone_bd_ram_mem3_reg[24][25]/P0001 , \wishbone_bd_ram_mem3_reg[24][26]/P0001 , \wishbone_bd_ram_mem3_reg[24][27]/P0001 , \wishbone_bd_ram_mem3_reg[24][28]/P0001 , \wishbone_bd_ram_mem3_reg[24][29]/P0001 , \wishbone_bd_ram_mem3_reg[24][30]/P0001 , \wishbone_bd_ram_mem3_reg[24][31]/P0001 , \wishbone_bd_ram_mem3_reg[250][24]/P0001 , \wishbone_bd_ram_mem3_reg[250][25]/P0001 , \wishbone_bd_ram_mem3_reg[250][26]/P0001 , \wishbone_bd_ram_mem3_reg[250][27]/P0001 , \wishbone_bd_ram_mem3_reg[250][28]/P0001 , \wishbone_bd_ram_mem3_reg[250][29]/P0001 , \wishbone_bd_ram_mem3_reg[250][30]/P0001 , \wishbone_bd_ram_mem3_reg[250][31]/P0001 , \wishbone_bd_ram_mem3_reg[251][24]/P0001 , \wishbone_bd_ram_mem3_reg[251][25]/P0001 , \wishbone_bd_ram_mem3_reg[251][26]/P0001 , \wishbone_bd_ram_mem3_reg[251][27]/P0001 , \wishbone_bd_ram_mem3_reg[251][28]/P0001 , \wishbone_bd_ram_mem3_reg[251][29]/P0001 , \wishbone_bd_ram_mem3_reg[251][30]/P0001 , \wishbone_bd_ram_mem3_reg[251][31]/P0001 , \wishbone_bd_ram_mem3_reg[252][24]/P0001 , \wishbone_bd_ram_mem3_reg[252][25]/P0001 , \wishbone_bd_ram_mem3_reg[252][26]/P0001 , \wishbone_bd_ram_mem3_reg[252][27]/P0001 , \wishbone_bd_ram_mem3_reg[252][28]/P0001 , \wishbone_bd_ram_mem3_reg[252][29]/P0001 , \wishbone_bd_ram_mem3_reg[252][30]/P0001 , \wishbone_bd_ram_mem3_reg[252][31]/P0001 , \wishbone_bd_ram_mem3_reg[253][24]/P0001 , \wishbone_bd_ram_mem3_reg[253][25]/P0001 , \wishbone_bd_ram_mem3_reg[253][26]/P0001 , \wishbone_bd_ram_mem3_reg[253][27]/P0001 , \wishbone_bd_ram_mem3_reg[253][28]/P0001 , \wishbone_bd_ram_mem3_reg[253][29]/P0001 , \wishbone_bd_ram_mem3_reg[253][30]/P0001 , \wishbone_bd_ram_mem3_reg[253][31]/P0001 , \wishbone_bd_ram_mem3_reg[254][24]/P0001 , \wishbone_bd_ram_mem3_reg[254][25]/P0001 , \wishbone_bd_ram_mem3_reg[254][26]/P0001 , \wishbone_bd_ram_mem3_reg[254][27]/P0001 , \wishbone_bd_ram_mem3_reg[254][28]/P0001 , \wishbone_bd_ram_mem3_reg[254][29]/P0001 , \wishbone_bd_ram_mem3_reg[254][30]/P0001 , \wishbone_bd_ram_mem3_reg[254][31]/P0001 , \wishbone_bd_ram_mem3_reg[255][24]/P0001 , \wishbone_bd_ram_mem3_reg[255][25]/P0001 , \wishbone_bd_ram_mem3_reg[255][26]/P0001 , \wishbone_bd_ram_mem3_reg[255][27]/P0001 , \wishbone_bd_ram_mem3_reg[255][28]/P0001 , \wishbone_bd_ram_mem3_reg[255][29]/P0001 , \wishbone_bd_ram_mem3_reg[255][30]/P0001 , \wishbone_bd_ram_mem3_reg[255][31]/P0001 , \wishbone_bd_ram_mem3_reg[25][24]/P0001 , \wishbone_bd_ram_mem3_reg[25][25]/P0001 , \wishbone_bd_ram_mem3_reg[25][26]/P0001 , \wishbone_bd_ram_mem3_reg[25][27]/P0001 , \wishbone_bd_ram_mem3_reg[25][28]/P0001 , \wishbone_bd_ram_mem3_reg[25][29]/P0001 , \wishbone_bd_ram_mem3_reg[25][30]/P0001 , \wishbone_bd_ram_mem3_reg[25][31]/P0001 , \wishbone_bd_ram_mem3_reg[26][24]/P0001 , \wishbone_bd_ram_mem3_reg[26][25]/P0001 , \wishbone_bd_ram_mem3_reg[26][26]/P0001 , \wishbone_bd_ram_mem3_reg[26][27]/P0001 , \wishbone_bd_ram_mem3_reg[26][28]/P0001 , \wishbone_bd_ram_mem3_reg[26][29]/P0001 , \wishbone_bd_ram_mem3_reg[26][30]/P0001 , \wishbone_bd_ram_mem3_reg[26][31]/P0001 , \wishbone_bd_ram_mem3_reg[27][24]/P0001 , \wishbone_bd_ram_mem3_reg[27][25]/P0001 , \wishbone_bd_ram_mem3_reg[27][26]/P0001 , \wishbone_bd_ram_mem3_reg[27][27]/P0001 , \wishbone_bd_ram_mem3_reg[27][28]/P0001 , \wishbone_bd_ram_mem3_reg[27][29]/P0001 , \wishbone_bd_ram_mem3_reg[27][30]/P0001 , \wishbone_bd_ram_mem3_reg[27][31]/P0001 , \wishbone_bd_ram_mem3_reg[28][24]/P0001 , \wishbone_bd_ram_mem3_reg[28][25]/P0001 , \wishbone_bd_ram_mem3_reg[28][26]/P0001 , \wishbone_bd_ram_mem3_reg[28][27]/P0001 , \wishbone_bd_ram_mem3_reg[28][28]/P0001 , \wishbone_bd_ram_mem3_reg[28][29]/P0001 , \wishbone_bd_ram_mem3_reg[28][30]/P0001 , \wishbone_bd_ram_mem3_reg[28][31]/P0001 , \wishbone_bd_ram_mem3_reg[29][24]/P0001 , \wishbone_bd_ram_mem3_reg[29][25]/P0001 , \wishbone_bd_ram_mem3_reg[29][26]/P0001 , \wishbone_bd_ram_mem3_reg[29][27]/P0001 , \wishbone_bd_ram_mem3_reg[29][28]/P0001 , \wishbone_bd_ram_mem3_reg[29][29]/P0001 , \wishbone_bd_ram_mem3_reg[29][30]/P0001 , \wishbone_bd_ram_mem3_reg[29][31]/P0001 , \wishbone_bd_ram_mem3_reg[2][24]/P0001 , \wishbone_bd_ram_mem3_reg[2][25]/P0001 , \wishbone_bd_ram_mem3_reg[2][26]/P0001 , \wishbone_bd_ram_mem3_reg[2][27]/P0001 , \wishbone_bd_ram_mem3_reg[2][28]/P0001 , \wishbone_bd_ram_mem3_reg[2][29]/P0001 , \wishbone_bd_ram_mem3_reg[2][30]/P0001 , \wishbone_bd_ram_mem3_reg[2][31]/P0001 , \wishbone_bd_ram_mem3_reg[30][24]/P0001 , \wishbone_bd_ram_mem3_reg[30][25]/P0001 , \wishbone_bd_ram_mem3_reg[30][26]/P0001 , \wishbone_bd_ram_mem3_reg[30][27]/P0001 , \wishbone_bd_ram_mem3_reg[30][28]/P0001 , \wishbone_bd_ram_mem3_reg[30][29]/P0001 , \wishbone_bd_ram_mem3_reg[30][30]/P0001 , \wishbone_bd_ram_mem3_reg[30][31]/P0001 , \wishbone_bd_ram_mem3_reg[31][24]/P0001 , \wishbone_bd_ram_mem3_reg[31][25]/P0001 , \wishbone_bd_ram_mem3_reg[31][26]/P0001 , \wishbone_bd_ram_mem3_reg[31][27]/P0001 , \wishbone_bd_ram_mem3_reg[31][28]/P0001 , \wishbone_bd_ram_mem3_reg[31][29]/P0001 , \wishbone_bd_ram_mem3_reg[31][30]/P0001 , \wishbone_bd_ram_mem3_reg[31][31]/P0001 , \wishbone_bd_ram_mem3_reg[32][24]/P0001 , \wishbone_bd_ram_mem3_reg[32][25]/P0001 , \wishbone_bd_ram_mem3_reg[32][26]/P0001 , \wishbone_bd_ram_mem3_reg[32][27]/P0001 , \wishbone_bd_ram_mem3_reg[32][28]/P0001 , \wishbone_bd_ram_mem3_reg[32][29]/P0001 , \wishbone_bd_ram_mem3_reg[32][30]/P0001 , \wishbone_bd_ram_mem3_reg[32][31]/P0001 , \wishbone_bd_ram_mem3_reg[33][24]/P0001 , \wishbone_bd_ram_mem3_reg[33][25]/P0001 , \wishbone_bd_ram_mem3_reg[33][26]/P0001 , \wishbone_bd_ram_mem3_reg[33][27]/P0001 , \wishbone_bd_ram_mem3_reg[33][28]/P0001 , \wishbone_bd_ram_mem3_reg[33][29]/P0001 , \wishbone_bd_ram_mem3_reg[33][30]/P0001 , \wishbone_bd_ram_mem3_reg[33][31]/P0001 , \wishbone_bd_ram_mem3_reg[34][24]/P0001 , \wishbone_bd_ram_mem3_reg[34][25]/P0001 , \wishbone_bd_ram_mem3_reg[34][26]/P0001 , \wishbone_bd_ram_mem3_reg[34][27]/P0001 , \wishbone_bd_ram_mem3_reg[34][28]/P0001 , \wishbone_bd_ram_mem3_reg[34][29]/P0001 , \wishbone_bd_ram_mem3_reg[34][30]/P0001 , \wishbone_bd_ram_mem3_reg[34][31]/P0001 , \wishbone_bd_ram_mem3_reg[35][24]/P0001 , \wishbone_bd_ram_mem3_reg[35][25]/P0001 , \wishbone_bd_ram_mem3_reg[35][26]/P0001 , \wishbone_bd_ram_mem3_reg[35][27]/P0001 , \wishbone_bd_ram_mem3_reg[35][28]/P0001 , \wishbone_bd_ram_mem3_reg[35][29]/P0001 , \wishbone_bd_ram_mem3_reg[35][30]/P0001 , \wishbone_bd_ram_mem3_reg[35][31]/P0001 , \wishbone_bd_ram_mem3_reg[36][24]/P0001 , \wishbone_bd_ram_mem3_reg[36][25]/P0001 , \wishbone_bd_ram_mem3_reg[36][26]/P0001 , \wishbone_bd_ram_mem3_reg[36][27]/P0001 , \wishbone_bd_ram_mem3_reg[36][28]/P0001 , \wishbone_bd_ram_mem3_reg[36][29]/P0001 , \wishbone_bd_ram_mem3_reg[36][30]/P0001 , \wishbone_bd_ram_mem3_reg[36][31]/P0001 , \wishbone_bd_ram_mem3_reg[37][24]/P0001 , \wishbone_bd_ram_mem3_reg[37][25]/P0001 , \wishbone_bd_ram_mem3_reg[37][26]/P0001 , \wishbone_bd_ram_mem3_reg[37][27]/P0001 , \wishbone_bd_ram_mem3_reg[37][28]/P0001 , \wishbone_bd_ram_mem3_reg[37][29]/P0001 , \wishbone_bd_ram_mem3_reg[37][30]/P0001 , \wishbone_bd_ram_mem3_reg[37][31]/P0001 , \wishbone_bd_ram_mem3_reg[38][24]/P0001 , \wishbone_bd_ram_mem3_reg[38][25]/P0001 , \wishbone_bd_ram_mem3_reg[38][26]/P0001 , \wishbone_bd_ram_mem3_reg[38][27]/P0001 , \wishbone_bd_ram_mem3_reg[38][28]/P0001 , \wishbone_bd_ram_mem3_reg[38][29]/P0001 , \wishbone_bd_ram_mem3_reg[38][30]/P0001 , \wishbone_bd_ram_mem3_reg[38][31]/P0001 , \wishbone_bd_ram_mem3_reg[39][24]/P0001 , \wishbone_bd_ram_mem3_reg[39][25]/P0001 , \wishbone_bd_ram_mem3_reg[39][26]/P0001 , \wishbone_bd_ram_mem3_reg[39][27]/P0001 , \wishbone_bd_ram_mem3_reg[39][28]/P0001 , \wishbone_bd_ram_mem3_reg[39][29]/P0001 , \wishbone_bd_ram_mem3_reg[39][30]/P0001 , \wishbone_bd_ram_mem3_reg[39][31]/P0001 , \wishbone_bd_ram_mem3_reg[3][24]/P0001 , \wishbone_bd_ram_mem3_reg[3][25]/P0001 , \wishbone_bd_ram_mem3_reg[3][26]/P0001 , \wishbone_bd_ram_mem3_reg[3][27]/P0001 , \wishbone_bd_ram_mem3_reg[3][28]/P0001 , \wishbone_bd_ram_mem3_reg[3][29]/P0001 , \wishbone_bd_ram_mem3_reg[3][30]/P0001 , \wishbone_bd_ram_mem3_reg[3][31]/P0001 , \wishbone_bd_ram_mem3_reg[40][24]/P0001 , \wishbone_bd_ram_mem3_reg[40][25]/P0001 , \wishbone_bd_ram_mem3_reg[40][26]/P0001 , \wishbone_bd_ram_mem3_reg[40][27]/P0001 , \wishbone_bd_ram_mem3_reg[40][28]/P0001 , \wishbone_bd_ram_mem3_reg[40][29]/P0001 , \wishbone_bd_ram_mem3_reg[40][30]/P0001 , \wishbone_bd_ram_mem3_reg[40][31]/P0001 , \wishbone_bd_ram_mem3_reg[41][24]/P0001 , \wishbone_bd_ram_mem3_reg[41][25]/P0001 , \wishbone_bd_ram_mem3_reg[41][26]/P0001 , \wishbone_bd_ram_mem3_reg[41][27]/P0001 , \wishbone_bd_ram_mem3_reg[41][28]/P0001 , \wishbone_bd_ram_mem3_reg[41][29]/P0001 , \wishbone_bd_ram_mem3_reg[41][30]/P0001 , \wishbone_bd_ram_mem3_reg[41][31]/P0001 , \wishbone_bd_ram_mem3_reg[42][24]/P0001 , \wishbone_bd_ram_mem3_reg[42][25]/P0001 , \wishbone_bd_ram_mem3_reg[42][26]/P0001 , \wishbone_bd_ram_mem3_reg[42][27]/P0001 , \wishbone_bd_ram_mem3_reg[42][28]/P0001 , \wishbone_bd_ram_mem3_reg[42][29]/P0001 , \wishbone_bd_ram_mem3_reg[42][30]/P0001 , \wishbone_bd_ram_mem3_reg[42][31]/P0001 , \wishbone_bd_ram_mem3_reg[43][24]/P0001 , \wishbone_bd_ram_mem3_reg[43][25]/P0001 , \wishbone_bd_ram_mem3_reg[43][26]/P0001 , \wishbone_bd_ram_mem3_reg[43][27]/P0001 , \wishbone_bd_ram_mem3_reg[43][28]/P0001 , \wishbone_bd_ram_mem3_reg[43][29]/P0001 , \wishbone_bd_ram_mem3_reg[43][30]/P0001 , \wishbone_bd_ram_mem3_reg[43][31]/P0001 , \wishbone_bd_ram_mem3_reg[44][24]/P0001 , \wishbone_bd_ram_mem3_reg[44][25]/P0001 , \wishbone_bd_ram_mem3_reg[44][26]/P0001 , \wishbone_bd_ram_mem3_reg[44][27]/P0001 , \wishbone_bd_ram_mem3_reg[44][28]/P0001 , \wishbone_bd_ram_mem3_reg[44][29]/P0001 , \wishbone_bd_ram_mem3_reg[44][30]/P0001 , \wishbone_bd_ram_mem3_reg[44][31]/P0001 , \wishbone_bd_ram_mem3_reg[45][24]/P0001 , \wishbone_bd_ram_mem3_reg[45][25]/P0001 , \wishbone_bd_ram_mem3_reg[45][26]/P0001 , \wishbone_bd_ram_mem3_reg[45][27]/P0001 , \wishbone_bd_ram_mem3_reg[45][28]/P0001 , \wishbone_bd_ram_mem3_reg[45][29]/P0001 , \wishbone_bd_ram_mem3_reg[45][30]/P0001 , \wishbone_bd_ram_mem3_reg[45][31]/P0001 , \wishbone_bd_ram_mem3_reg[46][24]/P0001 , \wishbone_bd_ram_mem3_reg[46][25]/P0001 , \wishbone_bd_ram_mem3_reg[46][26]/P0001 , \wishbone_bd_ram_mem3_reg[46][27]/P0001 , \wishbone_bd_ram_mem3_reg[46][28]/P0001 , \wishbone_bd_ram_mem3_reg[46][29]/P0001 , \wishbone_bd_ram_mem3_reg[46][30]/P0001 , \wishbone_bd_ram_mem3_reg[46][31]/P0001 , \wishbone_bd_ram_mem3_reg[47][24]/P0001 , \wishbone_bd_ram_mem3_reg[47][25]/P0001 , \wishbone_bd_ram_mem3_reg[47][26]/P0001 , \wishbone_bd_ram_mem3_reg[47][27]/P0001 , \wishbone_bd_ram_mem3_reg[47][28]/P0001 , \wishbone_bd_ram_mem3_reg[47][29]/P0001 , \wishbone_bd_ram_mem3_reg[47][30]/P0001 , \wishbone_bd_ram_mem3_reg[47][31]/P0001 , \wishbone_bd_ram_mem3_reg[48][24]/P0001 , \wishbone_bd_ram_mem3_reg[48][25]/P0001 , \wishbone_bd_ram_mem3_reg[48][26]/P0001 , \wishbone_bd_ram_mem3_reg[48][27]/P0001 , \wishbone_bd_ram_mem3_reg[48][28]/P0001 , \wishbone_bd_ram_mem3_reg[48][29]/P0001 , \wishbone_bd_ram_mem3_reg[48][30]/P0001 , \wishbone_bd_ram_mem3_reg[48][31]/P0001 , \wishbone_bd_ram_mem3_reg[49][24]/P0001 , \wishbone_bd_ram_mem3_reg[49][25]/P0001 , \wishbone_bd_ram_mem3_reg[49][26]/P0001 , \wishbone_bd_ram_mem3_reg[49][27]/P0001 , \wishbone_bd_ram_mem3_reg[49][28]/P0001 , \wishbone_bd_ram_mem3_reg[49][29]/P0001 , \wishbone_bd_ram_mem3_reg[49][30]/P0001 , \wishbone_bd_ram_mem3_reg[49][31]/P0001 , \wishbone_bd_ram_mem3_reg[4][24]/P0001 , \wishbone_bd_ram_mem3_reg[4][25]/P0001 , \wishbone_bd_ram_mem3_reg[4][26]/P0001 , \wishbone_bd_ram_mem3_reg[4][27]/P0001 , \wishbone_bd_ram_mem3_reg[4][28]/P0001 , \wishbone_bd_ram_mem3_reg[4][29]/P0001 , \wishbone_bd_ram_mem3_reg[4][30]/P0001 , \wishbone_bd_ram_mem3_reg[4][31]/P0001 , \wishbone_bd_ram_mem3_reg[50][24]/P0001 , \wishbone_bd_ram_mem3_reg[50][25]/P0001 , \wishbone_bd_ram_mem3_reg[50][26]/P0001 , \wishbone_bd_ram_mem3_reg[50][27]/P0001 , \wishbone_bd_ram_mem3_reg[50][28]/P0001 , \wishbone_bd_ram_mem3_reg[50][29]/P0001 , \wishbone_bd_ram_mem3_reg[50][30]/P0001 , \wishbone_bd_ram_mem3_reg[50][31]/P0001 , \wishbone_bd_ram_mem3_reg[51][24]/P0001 , \wishbone_bd_ram_mem3_reg[51][25]/P0001 , \wishbone_bd_ram_mem3_reg[51][26]/P0001 , \wishbone_bd_ram_mem3_reg[51][27]/P0001 , \wishbone_bd_ram_mem3_reg[51][28]/P0001 , \wishbone_bd_ram_mem3_reg[51][29]/P0001 , \wishbone_bd_ram_mem3_reg[51][30]/P0001 , \wishbone_bd_ram_mem3_reg[51][31]/P0001 , \wishbone_bd_ram_mem3_reg[52][24]/P0001 , \wishbone_bd_ram_mem3_reg[52][25]/P0001 , \wishbone_bd_ram_mem3_reg[52][26]/P0001 , \wishbone_bd_ram_mem3_reg[52][27]/P0001 , \wishbone_bd_ram_mem3_reg[52][28]/P0001 , \wishbone_bd_ram_mem3_reg[52][29]/P0001 , \wishbone_bd_ram_mem3_reg[52][30]/P0001 , \wishbone_bd_ram_mem3_reg[52][31]/P0001 , \wishbone_bd_ram_mem3_reg[53][24]/P0001 , \wishbone_bd_ram_mem3_reg[53][25]/P0001 , \wishbone_bd_ram_mem3_reg[53][26]/P0001 , \wishbone_bd_ram_mem3_reg[53][27]/P0001 , \wishbone_bd_ram_mem3_reg[53][28]/P0001 , \wishbone_bd_ram_mem3_reg[53][29]/P0001 , \wishbone_bd_ram_mem3_reg[53][30]/P0001 , \wishbone_bd_ram_mem3_reg[53][31]/P0001 , \wishbone_bd_ram_mem3_reg[54][24]/P0001 , \wishbone_bd_ram_mem3_reg[54][25]/P0001 , \wishbone_bd_ram_mem3_reg[54][26]/P0001 , \wishbone_bd_ram_mem3_reg[54][27]/P0001 , \wishbone_bd_ram_mem3_reg[54][28]/P0001 , \wishbone_bd_ram_mem3_reg[54][29]/P0001 , \wishbone_bd_ram_mem3_reg[54][30]/P0001 , \wishbone_bd_ram_mem3_reg[54][31]/P0001 , \wishbone_bd_ram_mem3_reg[55][24]/P0001 , \wishbone_bd_ram_mem3_reg[55][25]/P0001 , \wishbone_bd_ram_mem3_reg[55][26]/P0001 , \wishbone_bd_ram_mem3_reg[55][27]/P0001 , \wishbone_bd_ram_mem3_reg[55][28]/P0001 , \wishbone_bd_ram_mem3_reg[55][29]/P0001 , \wishbone_bd_ram_mem3_reg[55][30]/P0001 , \wishbone_bd_ram_mem3_reg[55][31]/P0001 , \wishbone_bd_ram_mem3_reg[56][24]/P0001 , \wishbone_bd_ram_mem3_reg[56][25]/P0001 , \wishbone_bd_ram_mem3_reg[56][26]/P0001 , \wishbone_bd_ram_mem3_reg[56][27]/P0001 , \wishbone_bd_ram_mem3_reg[56][28]/P0001 , \wishbone_bd_ram_mem3_reg[56][29]/P0001 , \wishbone_bd_ram_mem3_reg[56][30]/P0001 , \wishbone_bd_ram_mem3_reg[56][31]/P0001 , \wishbone_bd_ram_mem3_reg[57][24]/P0001 , \wishbone_bd_ram_mem3_reg[57][25]/P0001 , \wishbone_bd_ram_mem3_reg[57][26]/P0001 , \wishbone_bd_ram_mem3_reg[57][27]/P0001 , \wishbone_bd_ram_mem3_reg[57][28]/P0001 , \wishbone_bd_ram_mem3_reg[57][29]/P0001 , \wishbone_bd_ram_mem3_reg[57][30]/P0001 , \wishbone_bd_ram_mem3_reg[57][31]/P0001 , \wishbone_bd_ram_mem3_reg[58][24]/P0001 , \wishbone_bd_ram_mem3_reg[58][25]/P0001 , \wishbone_bd_ram_mem3_reg[58][26]/P0001 , \wishbone_bd_ram_mem3_reg[58][27]/P0001 , \wishbone_bd_ram_mem3_reg[58][28]/P0001 , \wishbone_bd_ram_mem3_reg[58][29]/P0001 , \wishbone_bd_ram_mem3_reg[58][30]/P0001 , \wishbone_bd_ram_mem3_reg[58][31]/P0001 , \wishbone_bd_ram_mem3_reg[59][24]/P0001 , \wishbone_bd_ram_mem3_reg[59][25]/P0001 , \wishbone_bd_ram_mem3_reg[59][26]/P0001 , \wishbone_bd_ram_mem3_reg[59][27]/P0001 , \wishbone_bd_ram_mem3_reg[59][28]/P0001 , \wishbone_bd_ram_mem3_reg[59][29]/P0001 , \wishbone_bd_ram_mem3_reg[59][30]/P0001 , \wishbone_bd_ram_mem3_reg[59][31]/P0001 , \wishbone_bd_ram_mem3_reg[5][24]/P0001 , \wishbone_bd_ram_mem3_reg[5][25]/P0001 , \wishbone_bd_ram_mem3_reg[5][26]/P0001 , \wishbone_bd_ram_mem3_reg[5][27]/P0001 , \wishbone_bd_ram_mem3_reg[5][28]/P0001 , \wishbone_bd_ram_mem3_reg[5][29]/P0001 , \wishbone_bd_ram_mem3_reg[5][30]/P0001 , \wishbone_bd_ram_mem3_reg[5][31]/P0001 , \wishbone_bd_ram_mem3_reg[60][24]/P0001 , \wishbone_bd_ram_mem3_reg[60][25]/P0001 , \wishbone_bd_ram_mem3_reg[60][26]/P0001 , \wishbone_bd_ram_mem3_reg[60][27]/P0001 , \wishbone_bd_ram_mem3_reg[60][28]/P0001 , \wishbone_bd_ram_mem3_reg[60][29]/P0001 , \wishbone_bd_ram_mem3_reg[60][30]/P0001 , \wishbone_bd_ram_mem3_reg[60][31]/P0001 , \wishbone_bd_ram_mem3_reg[61][24]/P0001 , \wishbone_bd_ram_mem3_reg[61][25]/P0001 , \wishbone_bd_ram_mem3_reg[61][26]/P0001 , \wishbone_bd_ram_mem3_reg[61][27]/P0001 , \wishbone_bd_ram_mem3_reg[61][28]/P0001 , \wishbone_bd_ram_mem3_reg[61][29]/P0001 , \wishbone_bd_ram_mem3_reg[61][30]/P0001 , \wishbone_bd_ram_mem3_reg[61][31]/P0001 , \wishbone_bd_ram_mem3_reg[62][24]/P0001 , \wishbone_bd_ram_mem3_reg[62][25]/P0001 , \wishbone_bd_ram_mem3_reg[62][26]/P0001 , \wishbone_bd_ram_mem3_reg[62][27]/P0001 , \wishbone_bd_ram_mem3_reg[62][28]/P0001 , \wishbone_bd_ram_mem3_reg[62][29]/P0001 , \wishbone_bd_ram_mem3_reg[62][30]/P0001 , \wishbone_bd_ram_mem3_reg[62][31]/P0001 , \wishbone_bd_ram_mem3_reg[63][24]/P0001 , \wishbone_bd_ram_mem3_reg[63][25]/P0001 , \wishbone_bd_ram_mem3_reg[63][26]/P0001 , \wishbone_bd_ram_mem3_reg[63][27]/P0001 , \wishbone_bd_ram_mem3_reg[63][28]/P0001 , \wishbone_bd_ram_mem3_reg[63][29]/P0001 , \wishbone_bd_ram_mem3_reg[63][30]/P0001 , \wishbone_bd_ram_mem3_reg[63][31]/P0001 , \wishbone_bd_ram_mem3_reg[64][24]/P0001 , \wishbone_bd_ram_mem3_reg[64][25]/P0001 , \wishbone_bd_ram_mem3_reg[64][26]/P0001 , \wishbone_bd_ram_mem3_reg[64][27]/P0001 , \wishbone_bd_ram_mem3_reg[64][28]/P0001 , \wishbone_bd_ram_mem3_reg[64][29]/P0001 , \wishbone_bd_ram_mem3_reg[64][30]/P0001 , \wishbone_bd_ram_mem3_reg[64][31]/P0001 , \wishbone_bd_ram_mem3_reg[65][24]/P0001 , \wishbone_bd_ram_mem3_reg[65][25]/P0001 , \wishbone_bd_ram_mem3_reg[65][26]/P0001 , \wishbone_bd_ram_mem3_reg[65][27]/P0001 , \wishbone_bd_ram_mem3_reg[65][28]/P0001 , \wishbone_bd_ram_mem3_reg[65][29]/P0001 , \wishbone_bd_ram_mem3_reg[65][30]/P0001 , \wishbone_bd_ram_mem3_reg[65][31]/P0001 , \wishbone_bd_ram_mem3_reg[66][24]/P0001 , \wishbone_bd_ram_mem3_reg[66][25]/P0001 , \wishbone_bd_ram_mem3_reg[66][26]/P0001 , \wishbone_bd_ram_mem3_reg[66][27]/P0001 , \wishbone_bd_ram_mem3_reg[66][28]/P0001 , \wishbone_bd_ram_mem3_reg[66][29]/P0001 , \wishbone_bd_ram_mem3_reg[66][30]/P0001 , \wishbone_bd_ram_mem3_reg[66][31]/P0001 , \wishbone_bd_ram_mem3_reg[67][24]/P0001 , \wishbone_bd_ram_mem3_reg[67][25]/P0001 , \wishbone_bd_ram_mem3_reg[67][26]/P0001 , \wishbone_bd_ram_mem3_reg[67][27]/P0001 , \wishbone_bd_ram_mem3_reg[67][28]/P0001 , \wishbone_bd_ram_mem3_reg[67][29]/P0001 , \wishbone_bd_ram_mem3_reg[67][30]/P0001 , \wishbone_bd_ram_mem3_reg[67][31]/P0001 , \wishbone_bd_ram_mem3_reg[68][24]/P0001 , \wishbone_bd_ram_mem3_reg[68][25]/P0001 , \wishbone_bd_ram_mem3_reg[68][26]/P0001 , \wishbone_bd_ram_mem3_reg[68][27]/P0001 , \wishbone_bd_ram_mem3_reg[68][28]/P0001 , \wishbone_bd_ram_mem3_reg[68][29]/P0001 , \wishbone_bd_ram_mem3_reg[68][30]/P0001 , \wishbone_bd_ram_mem3_reg[68][31]/P0001 , \wishbone_bd_ram_mem3_reg[69][24]/P0001 , \wishbone_bd_ram_mem3_reg[69][25]/P0001 , \wishbone_bd_ram_mem3_reg[69][26]/P0001 , \wishbone_bd_ram_mem3_reg[69][27]/P0001 , \wishbone_bd_ram_mem3_reg[69][28]/P0001 , \wishbone_bd_ram_mem3_reg[69][29]/P0001 , \wishbone_bd_ram_mem3_reg[69][30]/P0001 , \wishbone_bd_ram_mem3_reg[69][31]/P0001 , \wishbone_bd_ram_mem3_reg[6][24]/P0001 , \wishbone_bd_ram_mem3_reg[6][25]/P0001 , \wishbone_bd_ram_mem3_reg[6][26]/P0001 , \wishbone_bd_ram_mem3_reg[6][27]/P0001 , \wishbone_bd_ram_mem3_reg[6][28]/P0001 , \wishbone_bd_ram_mem3_reg[6][29]/P0001 , \wishbone_bd_ram_mem3_reg[6][30]/P0001 , \wishbone_bd_ram_mem3_reg[6][31]/P0001 , \wishbone_bd_ram_mem3_reg[70][24]/P0001 , \wishbone_bd_ram_mem3_reg[70][25]/P0001 , \wishbone_bd_ram_mem3_reg[70][26]/P0001 , \wishbone_bd_ram_mem3_reg[70][27]/P0001 , \wishbone_bd_ram_mem3_reg[70][28]/P0001 , \wishbone_bd_ram_mem3_reg[70][29]/P0001 , \wishbone_bd_ram_mem3_reg[70][30]/P0001 , \wishbone_bd_ram_mem3_reg[70][31]/P0001 , \wishbone_bd_ram_mem3_reg[71][24]/P0001 , \wishbone_bd_ram_mem3_reg[71][25]/P0001 , \wishbone_bd_ram_mem3_reg[71][26]/P0001 , \wishbone_bd_ram_mem3_reg[71][27]/P0001 , \wishbone_bd_ram_mem3_reg[71][28]/P0001 , \wishbone_bd_ram_mem3_reg[71][29]/P0001 , \wishbone_bd_ram_mem3_reg[71][30]/P0001 , \wishbone_bd_ram_mem3_reg[71][31]/P0001 , \wishbone_bd_ram_mem3_reg[72][24]/P0001 , \wishbone_bd_ram_mem3_reg[72][25]/P0001 , \wishbone_bd_ram_mem3_reg[72][26]/P0001 , \wishbone_bd_ram_mem3_reg[72][27]/P0001 , \wishbone_bd_ram_mem3_reg[72][28]/P0001 , \wishbone_bd_ram_mem3_reg[72][29]/P0001 , \wishbone_bd_ram_mem3_reg[72][30]/P0001 , \wishbone_bd_ram_mem3_reg[72][31]/P0001 , \wishbone_bd_ram_mem3_reg[73][24]/P0001 , \wishbone_bd_ram_mem3_reg[73][25]/P0001 , \wishbone_bd_ram_mem3_reg[73][26]/P0001 , \wishbone_bd_ram_mem3_reg[73][27]/P0001 , \wishbone_bd_ram_mem3_reg[73][28]/P0001 , \wishbone_bd_ram_mem3_reg[73][29]/P0001 , \wishbone_bd_ram_mem3_reg[73][30]/P0001 , \wishbone_bd_ram_mem3_reg[73][31]/P0001 , \wishbone_bd_ram_mem3_reg[74][24]/P0001 , \wishbone_bd_ram_mem3_reg[74][25]/P0001 , \wishbone_bd_ram_mem3_reg[74][26]/P0001 , \wishbone_bd_ram_mem3_reg[74][27]/P0001 , \wishbone_bd_ram_mem3_reg[74][28]/P0001 , \wishbone_bd_ram_mem3_reg[74][29]/P0001 , \wishbone_bd_ram_mem3_reg[74][30]/P0001 , \wishbone_bd_ram_mem3_reg[74][31]/P0001 , \wishbone_bd_ram_mem3_reg[75][24]/P0001 , \wishbone_bd_ram_mem3_reg[75][25]/P0001 , \wishbone_bd_ram_mem3_reg[75][26]/P0001 , \wishbone_bd_ram_mem3_reg[75][27]/P0001 , \wishbone_bd_ram_mem3_reg[75][28]/P0001 , \wishbone_bd_ram_mem3_reg[75][29]/P0001 , \wishbone_bd_ram_mem3_reg[75][30]/P0001 , \wishbone_bd_ram_mem3_reg[75][31]/P0001 , \wishbone_bd_ram_mem3_reg[76][24]/P0001 , \wishbone_bd_ram_mem3_reg[76][25]/P0001 , \wishbone_bd_ram_mem3_reg[76][26]/P0001 , \wishbone_bd_ram_mem3_reg[76][27]/P0001 , \wishbone_bd_ram_mem3_reg[76][28]/P0001 , \wishbone_bd_ram_mem3_reg[76][29]/P0001 , \wishbone_bd_ram_mem3_reg[76][30]/P0001 , \wishbone_bd_ram_mem3_reg[76][31]/P0001 , \wishbone_bd_ram_mem3_reg[77][24]/P0001 , \wishbone_bd_ram_mem3_reg[77][25]/P0001 , \wishbone_bd_ram_mem3_reg[77][26]/P0001 , \wishbone_bd_ram_mem3_reg[77][27]/P0001 , \wishbone_bd_ram_mem3_reg[77][28]/P0001 , \wishbone_bd_ram_mem3_reg[77][29]/P0001 , \wishbone_bd_ram_mem3_reg[77][30]/P0001 , \wishbone_bd_ram_mem3_reg[77][31]/P0001 , \wishbone_bd_ram_mem3_reg[78][24]/P0001 , \wishbone_bd_ram_mem3_reg[78][25]/P0001 , \wishbone_bd_ram_mem3_reg[78][26]/P0001 , \wishbone_bd_ram_mem3_reg[78][27]/P0001 , \wishbone_bd_ram_mem3_reg[78][28]/P0001 , \wishbone_bd_ram_mem3_reg[78][29]/P0001 , \wishbone_bd_ram_mem3_reg[78][30]/P0001 , \wishbone_bd_ram_mem3_reg[78][31]/P0001 , \wishbone_bd_ram_mem3_reg[79][24]/P0001 , \wishbone_bd_ram_mem3_reg[79][25]/P0001 , \wishbone_bd_ram_mem3_reg[79][26]/P0001 , \wishbone_bd_ram_mem3_reg[79][27]/P0001 , \wishbone_bd_ram_mem3_reg[79][28]/P0001 , \wishbone_bd_ram_mem3_reg[79][29]/P0001 , \wishbone_bd_ram_mem3_reg[79][30]/P0001 , \wishbone_bd_ram_mem3_reg[79][31]/P0001 , \wishbone_bd_ram_mem3_reg[7][24]/P0001 , \wishbone_bd_ram_mem3_reg[7][25]/P0001 , \wishbone_bd_ram_mem3_reg[7][26]/P0001 , \wishbone_bd_ram_mem3_reg[7][27]/P0001 , \wishbone_bd_ram_mem3_reg[7][28]/P0001 , \wishbone_bd_ram_mem3_reg[7][29]/P0001 , \wishbone_bd_ram_mem3_reg[7][30]/P0001 , \wishbone_bd_ram_mem3_reg[7][31]/P0001 , \wishbone_bd_ram_mem3_reg[80][24]/P0001 , \wishbone_bd_ram_mem3_reg[80][25]/P0001 , \wishbone_bd_ram_mem3_reg[80][26]/P0001 , \wishbone_bd_ram_mem3_reg[80][27]/P0001 , \wishbone_bd_ram_mem3_reg[80][28]/P0001 , \wishbone_bd_ram_mem3_reg[80][29]/P0001 , \wishbone_bd_ram_mem3_reg[80][30]/P0001 , \wishbone_bd_ram_mem3_reg[80][31]/P0001 , \wishbone_bd_ram_mem3_reg[81][24]/P0001 , \wishbone_bd_ram_mem3_reg[81][25]/P0001 , \wishbone_bd_ram_mem3_reg[81][26]/P0001 , \wishbone_bd_ram_mem3_reg[81][27]/P0001 , \wishbone_bd_ram_mem3_reg[81][28]/P0001 , \wishbone_bd_ram_mem3_reg[81][29]/P0001 , \wishbone_bd_ram_mem3_reg[81][30]/P0001 , \wishbone_bd_ram_mem3_reg[81][31]/P0001 , \wishbone_bd_ram_mem3_reg[82][24]/P0001 , \wishbone_bd_ram_mem3_reg[82][25]/P0001 , \wishbone_bd_ram_mem3_reg[82][26]/P0001 , \wishbone_bd_ram_mem3_reg[82][27]/P0001 , \wishbone_bd_ram_mem3_reg[82][28]/P0001 , \wishbone_bd_ram_mem3_reg[82][29]/P0001 , \wishbone_bd_ram_mem3_reg[82][30]/P0001 , \wishbone_bd_ram_mem3_reg[82][31]/P0001 , \wishbone_bd_ram_mem3_reg[83][24]/P0001 , \wishbone_bd_ram_mem3_reg[83][25]/P0001 , \wishbone_bd_ram_mem3_reg[83][26]/P0001 , \wishbone_bd_ram_mem3_reg[83][27]/P0001 , \wishbone_bd_ram_mem3_reg[83][28]/P0001 , \wishbone_bd_ram_mem3_reg[83][29]/P0001 , \wishbone_bd_ram_mem3_reg[83][30]/P0001 , \wishbone_bd_ram_mem3_reg[83][31]/P0001 , \wishbone_bd_ram_mem3_reg[84][24]/P0001 , \wishbone_bd_ram_mem3_reg[84][25]/P0001 , \wishbone_bd_ram_mem3_reg[84][26]/P0001 , \wishbone_bd_ram_mem3_reg[84][27]/P0001 , \wishbone_bd_ram_mem3_reg[84][28]/P0001 , \wishbone_bd_ram_mem3_reg[84][29]/P0001 , \wishbone_bd_ram_mem3_reg[84][30]/P0001 , \wishbone_bd_ram_mem3_reg[84][31]/P0001 , \wishbone_bd_ram_mem3_reg[85][24]/P0001 , \wishbone_bd_ram_mem3_reg[85][25]/P0001 , \wishbone_bd_ram_mem3_reg[85][26]/P0001 , \wishbone_bd_ram_mem3_reg[85][27]/P0001 , \wishbone_bd_ram_mem3_reg[85][28]/P0001 , \wishbone_bd_ram_mem3_reg[85][29]/P0001 , \wishbone_bd_ram_mem3_reg[85][30]/P0001 , \wishbone_bd_ram_mem3_reg[85][31]/P0001 , \wishbone_bd_ram_mem3_reg[86][24]/P0001 , \wishbone_bd_ram_mem3_reg[86][25]/P0001 , \wishbone_bd_ram_mem3_reg[86][26]/P0001 , \wishbone_bd_ram_mem3_reg[86][27]/P0001 , \wishbone_bd_ram_mem3_reg[86][28]/P0001 , \wishbone_bd_ram_mem3_reg[86][29]/P0001 , \wishbone_bd_ram_mem3_reg[86][30]/P0001 , \wishbone_bd_ram_mem3_reg[86][31]/P0001 , \wishbone_bd_ram_mem3_reg[87][24]/P0001 , \wishbone_bd_ram_mem3_reg[87][25]/P0001 , \wishbone_bd_ram_mem3_reg[87][26]/P0001 , \wishbone_bd_ram_mem3_reg[87][27]/P0001 , \wishbone_bd_ram_mem3_reg[87][28]/P0001 , \wishbone_bd_ram_mem3_reg[87][29]/P0001 , \wishbone_bd_ram_mem3_reg[87][30]/P0001 , \wishbone_bd_ram_mem3_reg[87][31]/P0001 , \wishbone_bd_ram_mem3_reg[88][24]/P0001 , \wishbone_bd_ram_mem3_reg[88][25]/P0001 , \wishbone_bd_ram_mem3_reg[88][26]/P0001 , \wishbone_bd_ram_mem3_reg[88][27]/P0001 , \wishbone_bd_ram_mem3_reg[88][28]/P0001 , \wishbone_bd_ram_mem3_reg[88][29]/P0001 , \wishbone_bd_ram_mem3_reg[88][30]/P0001 , \wishbone_bd_ram_mem3_reg[88][31]/P0001 , \wishbone_bd_ram_mem3_reg[89][24]/P0001 , \wishbone_bd_ram_mem3_reg[89][25]/P0001 , \wishbone_bd_ram_mem3_reg[89][26]/P0001 , \wishbone_bd_ram_mem3_reg[89][27]/P0001 , \wishbone_bd_ram_mem3_reg[89][28]/P0001 , \wishbone_bd_ram_mem3_reg[89][29]/P0001 , \wishbone_bd_ram_mem3_reg[89][30]/P0001 , \wishbone_bd_ram_mem3_reg[89][31]/P0001 , \wishbone_bd_ram_mem3_reg[8][24]/P0001 , \wishbone_bd_ram_mem3_reg[8][25]/P0001 , \wishbone_bd_ram_mem3_reg[8][26]/P0001 , \wishbone_bd_ram_mem3_reg[8][27]/P0001 , \wishbone_bd_ram_mem3_reg[8][28]/P0001 , \wishbone_bd_ram_mem3_reg[8][29]/P0001 , \wishbone_bd_ram_mem3_reg[8][30]/P0001 , \wishbone_bd_ram_mem3_reg[8][31]/P0001 , \wishbone_bd_ram_mem3_reg[90][24]/P0001 , \wishbone_bd_ram_mem3_reg[90][25]/P0001 , \wishbone_bd_ram_mem3_reg[90][26]/P0001 , \wishbone_bd_ram_mem3_reg[90][27]/P0001 , \wishbone_bd_ram_mem3_reg[90][28]/P0001 , \wishbone_bd_ram_mem3_reg[90][29]/P0001 , \wishbone_bd_ram_mem3_reg[90][30]/P0001 , \wishbone_bd_ram_mem3_reg[90][31]/P0001 , \wishbone_bd_ram_mem3_reg[91][24]/P0001 , \wishbone_bd_ram_mem3_reg[91][25]/P0001 , \wishbone_bd_ram_mem3_reg[91][26]/P0001 , \wishbone_bd_ram_mem3_reg[91][27]/P0001 , \wishbone_bd_ram_mem3_reg[91][28]/P0001 , \wishbone_bd_ram_mem3_reg[91][29]/P0001 , \wishbone_bd_ram_mem3_reg[91][30]/P0001 , \wishbone_bd_ram_mem3_reg[91][31]/P0001 , \wishbone_bd_ram_mem3_reg[92][24]/P0001 , \wishbone_bd_ram_mem3_reg[92][25]/P0001 , \wishbone_bd_ram_mem3_reg[92][26]/P0001 , \wishbone_bd_ram_mem3_reg[92][27]/P0001 , \wishbone_bd_ram_mem3_reg[92][28]/P0001 , \wishbone_bd_ram_mem3_reg[92][29]/P0001 , \wishbone_bd_ram_mem3_reg[92][30]/P0001 , \wishbone_bd_ram_mem3_reg[92][31]/P0001 , \wishbone_bd_ram_mem3_reg[93][24]/P0001 , \wishbone_bd_ram_mem3_reg[93][25]/P0001 , \wishbone_bd_ram_mem3_reg[93][26]/P0001 , \wishbone_bd_ram_mem3_reg[93][27]/P0001 , \wishbone_bd_ram_mem3_reg[93][28]/P0001 , \wishbone_bd_ram_mem3_reg[93][29]/P0001 , \wishbone_bd_ram_mem3_reg[93][30]/P0001 , \wishbone_bd_ram_mem3_reg[93][31]/P0001 , \wishbone_bd_ram_mem3_reg[94][24]/P0001 , \wishbone_bd_ram_mem3_reg[94][25]/P0001 , \wishbone_bd_ram_mem3_reg[94][26]/P0001 , \wishbone_bd_ram_mem3_reg[94][27]/P0001 , \wishbone_bd_ram_mem3_reg[94][28]/P0001 , \wishbone_bd_ram_mem3_reg[94][29]/P0001 , \wishbone_bd_ram_mem3_reg[94][30]/P0001 , \wishbone_bd_ram_mem3_reg[94][31]/P0001 , \wishbone_bd_ram_mem3_reg[95][24]/P0001 , \wishbone_bd_ram_mem3_reg[95][25]/P0001 , \wishbone_bd_ram_mem3_reg[95][26]/P0001 , \wishbone_bd_ram_mem3_reg[95][27]/P0001 , \wishbone_bd_ram_mem3_reg[95][28]/P0001 , \wishbone_bd_ram_mem3_reg[95][29]/P0001 , \wishbone_bd_ram_mem3_reg[95][30]/P0001 , \wishbone_bd_ram_mem3_reg[95][31]/P0001 , \wishbone_bd_ram_mem3_reg[96][24]/P0001 , \wishbone_bd_ram_mem3_reg[96][25]/P0001 , \wishbone_bd_ram_mem3_reg[96][26]/P0001 , \wishbone_bd_ram_mem3_reg[96][27]/P0001 , \wishbone_bd_ram_mem3_reg[96][28]/P0001 , \wishbone_bd_ram_mem3_reg[96][29]/P0001 , \wishbone_bd_ram_mem3_reg[96][30]/P0001 , \wishbone_bd_ram_mem3_reg[96][31]/P0001 , \wishbone_bd_ram_mem3_reg[97][24]/P0001 , \wishbone_bd_ram_mem3_reg[97][25]/P0001 , \wishbone_bd_ram_mem3_reg[97][26]/P0001 , \wishbone_bd_ram_mem3_reg[97][27]/P0001 , \wishbone_bd_ram_mem3_reg[97][28]/P0001 , \wishbone_bd_ram_mem3_reg[97][29]/P0001 , \wishbone_bd_ram_mem3_reg[97][30]/P0001 , \wishbone_bd_ram_mem3_reg[97][31]/P0001 , \wishbone_bd_ram_mem3_reg[98][24]/P0001 , \wishbone_bd_ram_mem3_reg[98][25]/P0001 , \wishbone_bd_ram_mem3_reg[98][26]/P0001 , \wishbone_bd_ram_mem3_reg[98][27]/P0001 , \wishbone_bd_ram_mem3_reg[98][28]/P0001 , \wishbone_bd_ram_mem3_reg[98][29]/P0001 , \wishbone_bd_ram_mem3_reg[98][30]/P0001 , \wishbone_bd_ram_mem3_reg[98][31]/P0001 , \wishbone_bd_ram_mem3_reg[99][24]/P0001 , \wishbone_bd_ram_mem3_reg[99][25]/P0001 , \wishbone_bd_ram_mem3_reg[99][26]/P0001 , \wishbone_bd_ram_mem3_reg[99][27]/P0001 , \wishbone_bd_ram_mem3_reg[99][28]/P0001 , \wishbone_bd_ram_mem3_reg[99][29]/P0001 , \wishbone_bd_ram_mem3_reg[99][30]/P0001 , \wishbone_bd_ram_mem3_reg[99][31]/P0001 , \wishbone_bd_ram_mem3_reg[9][24]/P0001 , \wishbone_bd_ram_mem3_reg[9][25]/P0001 , \wishbone_bd_ram_mem3_reg[9][26]/P0001 , \wishbone_bd_ram_mem3_reg[9][27]/P0001 , \wishbone_bd_ram_mem3_reg[9][28]/P0001 , \wishbone_bd_ram_mem3_reg[9][29]/P0001 , \wishbone_bd_ram_mem3_reg[9][30]/P0001 , \wishbone_bd_ram_mem3_reg[9][31]/P0001 , \wishbone_bd_ram_raddr_reg[0]/P0001 , \wishbone_bd_ram_raddr_reg[1]/NET0131 , \wishbone_bd_ram_raddr_reg[2]/NET0131 , \wishbone_bd_ram_raddr_reg[3]/P0001 , \wishbone_bd_ram_raddr_reg[4]/NET0131 , \wishbone_bd_ram_raddr_reg[5]/NET0131 , \wishbone_bd_ram_raddr_reg[6]/NET0131 , \wishbone_bd_ram_raddr_reg[7]/NET0131 , \wishbone_cyc_cleared_reg/NET0131 , \wishbone_r_RxEn_q_reg/NET0131 , \wishbone_r_TxEn_q_reg/NET0131 , \wishbone_ram_addr_reg[0]/NET0131 , \wishbone_ram_addr_reg[1]/NET0131 , \wishbone_ram_addr_reg[2]/NET0131 , \wishbone_ram_addr_reg[3]/NET0131 , \wishbone_ram_addr_reg[4]/NET0131 , \wishbone_ram_addr_reg[5]/NET0131 , \wishbone_ram_addr_reg[6]/NET0131 , \wishbone_ram_addr_reg[7]/NET0131 , \wishbone_ram_di_reg[0]/NET0131 , \wishbone_ram_di_reg[10]/NET0131 , \wishbone_ram_di_reg[11]/NET0131 , \wishbone_ram_di_reg[12]/NET0131 , \wishbone_ram_di_reg[13]/NET0131 , \wishbone_ram_di_reg[14]/NET0131 , \wishbone_ram_di_reg[15]/NET0131 , \wishbone_ram_di_reg[16]/NET0131 , \wishbone_ram_di_reg[17]/NET0131 , \wishbone_ram_di_reg[18]/NET0131 , \wishbone_ram_di_reg[19]/NET0131 , \wishbone_ram_di_reg[1]/NET0131 , \wishbone_ram_di_reg[20]/NET0131 , \wishbone_ram_di_reg[21]/NET0131 , \wishbone_ram_di_reg[22]/NET0131 , \wishbone_ram_di_reg[23]/NET0131 , \wishbone_ram_di_reg[24]/NET0131 , \wishbone_ram_di_reg[25]/NET0131 , \wishbone_ram_di_reg[26]/NET0131 , \wishbone_ram_di_reg[27]/NET0131 , \wishbone_ram_di_reg[28]/NET0131 , \wishbone_ram_di_reg[29]/NET0131 , \wishbone_ram_di_reg[2]/NET0131 , \wishbone_ram_di_reg[30]/NET0131 , \wishbone_ram_di_reg[31]/NET0131 , \wishbone_ram_di_reg[3]/NET0131 , \wishbone_ram_di_reg[4]/NET0131 , \wishbone_ram_di_reg[5]/NET0131 , \wishbone_ram_di_reg[6]/NET0131 , \wishbone_ram_di_reg[7]/NET0131 , \wishbone_ram_di_reg[8]/NET0131 , \wishbone_ram_di_reg[9]/NET0131 , \wishbone_rx_burst_cnt_reg[0]/NET0131 , \wishbone_rx_burst_cnt_reg[1]/NET0131 , \wishbone_rx_burst_cnt_reg[2]/NET0131 , \wishbone_rx_burst_en_reg/NET0131 , \wishbone_rx_fifo_cnt_reg[0]/NET0131 , \wishbone_rx_fifo_cnt_reg[1]/NET0131 , \wishbone_rx_fifo_cnt_reg[2]/NET0131 , \wishbone_rx_fifo_cnt_reg[3]/NET0131 , \wishbone_rx_fifo_cnt_reg[4]/NET0131 , \wishbone_rx_fifo_fifo_reg[0][0]/P0001 , \wishbone_rx_fifo_fifo_reg[0][10]/P0001 , \wishbone_rx_fifo_fifo_reg[0][11]/P0001 , \wishbone_rx_fifo_fifo_reg[0][12]/P0001 , \wishbone_rx_fifo_fifo_reg[0][13]/P0001 , \wishbone_rx_fifo_fifo_reg[0][14]/P0001 , \wishbone_rx_fifo_fifo_reg[0][15]/P0001 , \wishbone_rx_fifo_fifo_reg[0][16]/P0001 , \wishbone_rx_fifo_fifo_reg[0][17]/P0001 , \wishbone_rx_fifo_fifo_reg[0][18]/P0001 , \wishbone_rx_fifo_fifo_reg[0][19]/P0001 , \wishbone_rx_fifo_fifo_reg[0][1]/P0001 , \wishbone_rx_fifo_fifo_reg[0][20]/P0001 , \wishbone_rx_fifo_fifo_reg[0][21]/P0001 , \wishbone_rx_fifo_fifo_reg[0][22]/P0001 , \wishbone_rx_fifo_fifo_reg[0][23]/P0001 , \wishbone_rx_fifo_fifo_reg[0][24]/P0001 , \wishbone_rx_fifo_fifo_reg[0][25]/P0001 , \wishbone_rx_fifo_fifo_reg[0][26]/P0001 , \wishbone_rx_fifo_fifo_reg[0][27]/P0001 , \wishbone_rx_fifo_fifo_reg[0][28]/P0001 , \wishbone_rx_fifo_fifo_reg[0][29]/P0001 , \wishbone_rx_fifo_fifo_reg[0][2]/P0001 , \wishbone_rx_fifo_fifo_reg[0][30]/P0001 , \wishbone_rx_fifo_fifo_reg[0][31]/P0001 , \wishbone_rx_fifo_fifo_reg[0][3]/P0001 , \wishbone_rx_fifo_fifo_reg[0][4]/P0001 , \wishbone_rx_fifo_fifo_reg[0][5]/P0001 , \wishbone_rx_fifo_fifo_reg[0][6]/P0001 , \wishbone_rx_fifo_fifo_reg[0][7]/P0001 , \wishbone_rx_fifo_fifo_reg[0][8]/P0001 , \wishbone_rx_fifo_fifo_reg[0][9]/P0001 , \wishbone_rx_fifo_fifo_reg[10][0]/P0001 , \wishbone_rx_fifo_fifo_reg[10][10]/P0001 , \wishbone_rx_fifo_fifo_reg[10][11]/P0001 , \wishbone_rx_fifo_fifo_reg[10][12]/P0001 , \wishbone_rx_fifo_fifo_reg[10][13]/P0001 , \wishbone_rx_fifo_fifo_reg[10][14]/P0001 , \wishbone_rx_fifo_fifo_reg[10][15]/P0001 , \wishbone_rx_fifo_fifo_reg[10][16]/P0001 , \wishbone_rx_fifo_fifo_reg[10][17]/P0001 , \wishbone_rx_fifo_fifo_reg[10][18]/P0001 , \wishbone_rx_fifo_fifo_reg[10][19]/P0001 , \wishbone_rx_fifo_fifo_reg[10][1]/P0001 , \wishbone_rx_fifo_fifo_reg[10][20]/P0001 , \wishbone_rx_fifo_fifo_reg[10][21]/P0001 , \wishbone_rx_fifo_fifo_reg[10][22]/P0001 , \wishbone_rx_fifo_fifo_reg[10][23]/P0001 , \wishbone_rx_fifo_fifo_reg[10][24]/P0001 , \wishbone_rx_fifo_fifo_reg[10][25]/P0001 , \wishbone_rx_fifo_fifo_reg[10][26]/P0001 , \wishbone_rx_fifo_fifo_reg[10][27]/P0001 , \wishbone_rx_fifo_fifo_reg[10][28]/P0001 , \wishbone_rx_fifo_fifo_reg[10][29]/P0001 , \wishbone_rx_fifo_fifo_reg[10][2]/P0001 , \wishbone_rx_fifo_fifo_reg[10][30]/P0001 , \wishbone_rx_fifo_fifo_reg[10][31]/P0001 , \wishbone_rx_fifo_fifo_reg[10][3]/P0001 , \wishbone_rx_fifo_fifo_reg[10][4]/P0001 , \wishbone_rx_fifo_fifo_reg[10][5]/P0001 , \wishbone_rx_fifo_fifo_reg[10][6]/P0001 , \wishbone_rx_fifo_fifo_reg[10][7]/P0001 , \wishbone_rx_fifo_fifo_reg[10][8]/P0001 , \wishbone_rx_fifo_fifo_reg[10][9]/P0001 , \wishbone_rx_fifo_fifo_reg[11][0]/P0001 , \wishbone_rx_fifo_fifo_reg[11][10]/P0001 , \wishbone_rx_fifo_fifo_reg[11][11]/P0001 , \wishbone_rx_fifo_fifo_reg[11][12]/P0001 , \wishbone_rx_fifo_fifo_reg[11][13]/P0001 , \wishbone_rx_fifo_fifo_reg[11][14]/P0001 , \wishbone_rx_fifo_fifo_reg[11][15]/P0001 , \wishbone_rx_fifo_fifo_reg[11][16]/P0001 , \wishbone_rx_fifo_fifo_reg[11][17]/P0001 , \wishbone_rx_fifo_fifo_reg[11][18]/P0001 , \wishbone_rx_fifo_fifo_reg[11][19]/P0001 , \wishbone_rx_fifo_fifo_reg[11][1]/P0001 , \wishbone_rx_fifo_fifo_reg[11][20]/P0001 , \wishbone_rx_fifo_fifo_reg[11][21]/P0001 , \wishbone_rx_fifo_fifo_reg[11][22]/P0001 , \wishbone_rx_fifo_fifo_reg[11][23]/P0001 , \wishbone_rx_fifo_fifo_reg[11][24]/P0001 , \wishbone_rx_fifo_fifo_reg[11][25]/P0001 , \wishbone_rx_fifo_fifo_reg[11][26]/P0001 , \wishbone_rx_fifo_fifo_reg[11][27]/P0001 , \wishbone_rx_fifo_fifo_reg[11][28]/P0001 , \wishbone_rx_fifo_fifo_reg[11][29]/P0001 , \wishbone_rx_fifo_fifo_reg[11][2]/P0001 , \wishbone_rx_fifo_fifo_reg[11][30]/P0001 , \wishbone_rx_fifo_fifo_reg[11][31]/P0001 , \wishbone_rx_fifo_fifo_reg[11][3]/P0001 , \wishbone_rx_fifo_fifo_reg[11][4]/P0001 , \wishbone_rx_fifo_fifo_reg[11][5]/P0001 , \wishbone_rx_fifo_fifo_reg[11][6]/P0001 , \wishbone_rx_fifo_fifo_reg[11][7]/P0001 , \wishbone_rx_fifo_fifo_reg[11][8]/P0001 , \wishbone_rx_fifo_fifo_reg[11][9]/P0001 , \wishbone_rx_fifo_fifo_reg[12][0]/P0001 , \wishbone_rx_fifo_fifo_reg[12][10]/P0001 , \wishbone_rx_fifo_fifo_reg[12][11]/P0001 , \wishbone_rx_fifo_fifo_reg[12][12]/P0001 , \wishbone_rx_fifo_fifo_reg[12][13]/P0001 , \wishbone_rx_fifo_fifo_reg[12][14]/P0001 , \wishbone_rx_fifo_fifo_reg[12][15]/P0001 , \wishbone_rx_fifo_fifo_reg[12][16]/P0001 , \wishbone_rx_fifo_fifo_reg[12][17]/P0001 , \wishbone_rx_fifo_fifo_reg[12][18]/P0001 , \wishbone_rx_fifo_fifo_reg[12][19]/P0001 , \wishbone_rx_fifo_fifo_reg[12][1]/P0001 , \wishbone_rx_fifo_fifo_reg[12][20]/P0001 , \wishbone_rx_fifo_fifo_reg[12][21]/P0001 , \wishbone_rx_fifo_fifo_reg[12][22]/P0001 , \wishbone_rx_fifo_fifo_reg[12][23]/P0001 , \wishbone_rx_fifo_fifo_reg[12][24]/P0001 , \wishbone_rx_fifo_fifo_reg[12][25]/P0001 , \wishbone_rx_fifo_fifo_reg[12][26]/P0001 , \wishbone_rx_fifo_fifo_reg[12][27]/P0001 , \wishbone_rx_fifo_fifo_reg[12][28]/P0001 , \wishbone_rx_fifo_fifo_reg[12][29]/P0001 , \wishbone_rx_fifo_fifo_reg[12][2]/P0001 , \wishbone_rx_fifo_fifo_reg[12][30]/P0001 , \wishbone_rx_fifo_fifo_reg[12][31]/P0001 , \wishbone_rx_fifo_fifo_reg[12][3]/P0001 , \wishbone_rx_fifo_fifo_reg[12][4]/P0001 , \wishbone_rx_fifo_fifo_reg[12][5]/P0001 , \wishbone_rx_fifo_fifo_reg[12][6]/P0001 , \wishbone_rx_fifo_fifo_reg[12][7]/P0001 , \wishbone_rx_fifo_fifo_reg[12][8]/P0001 , \wishbone_rx_fifo_fifo_reg[12][9]/P0001 , \wishbone_rx_fifo_fifo_reg[13][0]/P0001 , \wishbone_rx_fifo_fifo_reg[13][10]/P0001 , \wishbone_rx_fifo_fifo_reg[13][11]/P0001 , \wishbone_rx_fifo_fifo_reg[13][12]/P0001 , \wishbone_rx_fifo_fifo_reg[13][13]/P0001 , \wishbone_rx_fifo_fifo_reg[13][14]/P0001 , \wishbone_rx_fifo_fifo_reg[13][15]/P0001 , \wishbone_rx_fifo_fifo_reg[13][16]/P0001 , \wishbone_rx_fifo_fifo_reg[13][17]/P0001 , \wishbone_rx_fifo_fifo_reg[13][18]/P0001 , \wishbone_rx_fifo_fifo_reg[13][19]/P0001 , \wishbone_rx_fifo_fifo_reg[13][1]/P0001 , \wishbone_rx_fifo_fifo_reg[13][20]/P0001 , \wishbone_rx_fifo_fifo_reg[13][21]/P0001 , \wishbone_rx_fifo_fifo_reg[13][22]/P0001 , \wishbone_rx_fifo_fifo_reg[13][23]/P0001 , \wishbone_rx_fifo_fifo_reg[13][24]/P0001 , \wishbone_rx_fifo_fifo_reg[13][25]/P0001 , \wishbone_rx_fifo_fifo_reg[13][26]/P0001 , \wishbone_rx_fifo_fifo_reg[13][27]/P0001 , \wishbone_rx_fifo_fifo_reg[13][28]/P0001 , \wishbone_rx_fifo_fifo_reg[13][29]/P0001 , \wishbone_rx_fifo_fifo_reg[13][2]/P0001 , \wishbone_rx_fifo_fifo_reg[13][30]/P0001 , \wishbone_rx_fifo_fifo_reg[13][31]/P0001 , \wishbone_rx_fifo_fifo_reg[13][3]/P0001 , \wishbone_rx_fifo_fifo_reg[13][4]/P0001 , \wishbone_rx_fifo_fifo_reg[13][5]/P0001 , \wishbone_rx_fifo_fifo_reg[13][6]/P0001 , \wishbone_rx_fifo_fifo_reg[13][7]/P0001 , \wishbone_rx_fifo_fifo_reg[13][8]/P0001 , \wishbone_rx_fifo_fifo_reg[13][9]/P0001 , \wishbone_rx_fifo_fifo_reg[14][0]/P0001 , \wishbone_rx_fifo_fifo_reg[14][10]/P0001 , \wishbone_rx_fifo_fifo_reg[14][11]/P0001 , \wishbone_rx_fifo_fifo_reg[14][12]/P0001 , \wishbone_rx_fifo_fifo_reg[14][13]/P0001 , \wishbone_rx_fifo_fifo_reg[14][14]/P0001 , \wishbone_rx_fifo_fifo_reg[14][15]/P0001 , \wishbone_rx_fifo_fifo_reg[14][16]/P0001 , \wishbone_rx_fifo_fifo_reg[14][17]/P0001 , \wishbone_rx_fifo_fifo_reg[14][18]/P0001 , \wishbone_rx_fifo_fifo_reg[14][19]/P0001 , \wishbone_rx_fifo_fifo_reg[14][1]/P0001 , \wishbone_rx_fifo_fifo_reg[14][20]/P0001 , \wishbone_rx_fifo_fifo_reg[14][21]/P0001 , \wishbone_rx_fifo_fifo_reg[14][22]/P0001 , \wishbone_rx_fifo_fifo_reg[14][23]/P0001 , \wishbone_rx_fifo_fifo_reg[14][24]/P0001 , \wishbone_rx_fifo_fifo_reg[14][25]/P0001 , \wishbone_rx_fifo_fifo_reg[14][26]/P0001 , \wishbone_rx_fifo_fifo_reg[14][27]/P0001 , \wishbone_rx_fifo_fifo_reg[14][28]/P0001 , \wishbone_rx_fifo_fifo_reg[14][29]/P0001 , \wishbone_rx_fifo_fifo_reg[14][2]/P0001 , \wishbone_rx_fifo_fifo_reg[14][30]/P0001 , \wishbone_rx_fifo_fifo_reg[14][31]/P0001 , \wishbone_rx_fifo_fifo_reg[14][3]/P0001 , \wishbone_rx_fifo_fifo_reg[14][4]/P0001 , \wishbone_rx_fifo_fifo_reg[14][5]/P0001 , \wishbone_rx_fifo_fifo_reg[14][6]/P0001 , \wishbone_rx_fifo_fifo_reg[14][7]/P0001 , \wishbone_rx_fifo_fifo_reg[14][8]/P0001 , \wishbone_rx_fifo_fifo_reg[14][9]/P0001 , \wishbone_rx_fifo_fifo_reg[15][0]/P0001 , \wishbone_rx_fifo_fifo_reg[15][10]/P0001 , \wishbone_rx_fifo_fifo_reg[15][11]/P0001 , \wishbone_rx_fifo_fifo_reg[15][12]/P0001 , \wishbone_rx_fifo_fifo_reg[15][13]/P0001 , \wishbone_rx_fifo_fifo_reg[15][14]/P0001 , \wishbone_rx_fifo_fifo_reg[15][15]/P0001 , \wishbone_rx_fifo_fifo_reg[15][16]/P0001 , \wishbone_rx_fifo_fifo_reg[15][17]/P0001 , \wishbone_rx_fifo_fifo_reg[15][18]/P0001 , \wishbone_rx_fifo_fifo_reg[15][19]/P0001 , \wishbone_rx_fifo_fifo_reg[15][1]/P0001 , \wishbone_rx_fifo_fifo_reg[15][20]/P0001 , \wishbone_rx_fifo_fifo_reg[15][21]/P0001 , \wishbone_rx_fifo_fifo_reg[15][22]/P0001 , \wishbone_rx_fifo_fifo_reg[15][23]/P0001 , \wishbone_rx_fifo_fifo_reg[15][24]/P0001 , \wishbone_rx_fifo_fifo_reg[15][25]/P0001 , \wishbone_rx_fifo_fifo_reg[15][26]/P0001 , \wishbone_rx_fifo_fifo_reg[15][27]/P0001 , \wishbone_rx_fifo_fifo_reg[15][28]/P0001 , \wishbone_rx_fifo_fifo_reg[15][29]/P0001 , \wishbone_rx_fifo_fifo_reg[15][2]/P0001 , \wishbone_rx_fifo_fifo_reg[15][30]/P0001 , \wishbone_rx_fifo_fifo_reg[15][31]/P0001 , \wishbone_rx_fifo_fifo_reg[15][3]/P0001 , \wishbone_rx_fifo_fifo_reg[15][4]/P0001 , \wishbone_rx_fifo_fifo_reg[15][5]/P0001 , \wishbone_rx_fifo_fifo_reg[15][6]/P0001 , \wishbone_rx_fifo_fifo_reg[15][7]/P0001 , \wishbone_rx_fifo_fifo_reg[15][8]/P0001 , \wishbone_rx_fifo_fifo_reg[15][9]/P0001 , \wishbone_rx_fifo_fifo_reg[1][0]/P0001 , \wishbone_rx_fifo_fifo_reg[1][10]/P0001 , \wishbone_rx_fifo_fifo_reg[1][11]/P0001 , \wishbone_rx_fifo_fifo_reg[1][12]/P0001 , \wishbone_rx_fifo_fifo_reg[1][13]/P0001 , \wishbone_rx_fifo_fifo_reg[1][14]/P0001 , \wishbone_rx_fifo_fifo_reg[1][15]/P0001 , \wishbone_rx_fifo_fifo_reg[1][16]/P0001 , \wishbone_rx_fifo_fifo_reg[1][17]/P0001 , \wishbone_rx_fifo_fifo_reg[1][18]/P0001 , \wishbone_rx_fifo_fifo_reg[1][19]/P0001 , \wishbone_rx_fifo_fifo_reg[1][1]/P0001 , \wishbone_rx_fifo_fifo_reg[1][20]/P0001 , \wishbone_rx_fifo_fifo_reg[1][21]/P0001 , \wishbone_rx_fifo_fifo_reg[1][22]/P0001 , \wishbone_rx_fifo_fifo_reg[1][23]/P0001 , \wishbone_rx_fifo_fifo_reg[1][24]/P0001 , \wishbone_rx_fifo_fifo_reg[1][25]/P0001 , \wishbone_rx_fifo_fifo_reg[1][26]/P0001 , \wishbone_rx_fifo_fifo_reg[1][27]/P0001 , \wishbone_rx_fifo_fifo_reg[1][28]/P0001 , \wishbone_rx_fifo_fifo_reg[1][29]/P0001 , \wishbone_rx_fifo_fifo_reg[1][2]/P0001 , \wishbone_rx_fifo_fifo_reg[1][30]/P0001 , \wishbone_rx_fifo_fifo_reg[1][31]/P0001 , \wishbone_rx_fifo_fifo_reg[1][3]/P0001 , \wishbone_rx_fifo_fifo_reg[1][4]/P0001 , \wishbone_rx_fifo_fifo_reg[1][5]/P0001 , \wishbone_rx_fifo_fifo_reg[1][6]/P0001 , \wishbone_rx_fifo_fifo_reg[1][7]/P0001 , \wishbone_rx_fifo_fifo_reg[1][8]/P0001 , \wishbone_rx_fifo_fifo_reg[1][9]/P0001 , \wishbone_rx_fifo_fifo_reg[2][0]/P0001 , \wishbone_rx_fifo_fifo_reg[2][10]/P0001 , \wishbone_rx_fifo_fifo_reg[2][11]/P0001 , \wishbone_rx_fifo_fifo_reg[2][12]/P0001 , \wishbone_rx_fifo_fifo_reg[2][13]/P0001 , \wishbone_rx_fifo_fifo_reg[2][14]/P0001 , \wishbone_rx_fifo_fifo_reg[2][15]/P0001 , \wishbone_rx_fifo_fifo_reg[2][16]/P0001 , \wishbone_rx_fifo_fifo_reg[2][17]/P0001 , \wishbone_rx_fifo_fifo_reg[2][18]/P0001 , \wishbone_rx_fifo_fifo_reg[2][19]/P0001 , \wishbone_rx_fifo_fifo_reg[2][1]/P0001 , \wishbone_rx_fifo_fifo_reg[2][20]/P0001 , \wishbone_rx_fifo_fifo_reg[2][21]/P0001 , \wishbone_rx_fifo_fifo_reg[2][22]/P0001 , \wishbone_rx_fifo_fifo_reg[2][23]/P0001 , \wishbone_rx_fifo_fifo_reg[2][24]/P0001 , \wishbone_rx_fifo_fifo_reg[2][25]/P0001 , \wishbone_rx_fifo_fifo_reg[2][26]/P0001 , \wishbone_rx_fifo_fifo_reg[2][27]/P0001 , \wishbone_rx_fifo_fifo_reg[2][28]/P0001 , \wishbone_rx_fifo_fifo_reg[2][29]/P0001 , \wishbone_rx_fifo_fifo_reg[2][2]/P0001 , \wishbone_rx_fifo_fifo_reg[2][30]/P0001 , \wishbone_rx_fifo_fifo_reg[2][31]/P0001 , \wishbone_rx_fifo_fifo_reg[2][3]/P0001 , \wishbone_rx_fifo_fifo_reg[2][4]/P0001 , \wishbone_rx_fifo_fifo_reg[2][5]/P0001 , \wishbone_rx_fifo_fifo_reg[2][6]/P0001 , \wishbone_rx_fifo_fifo_reg[2][7]/P0001 , \wishbone_rx_fifo_fifo_reg[2][8]/P0001 , \wishbone_rx_fifo_fifo_reg[2][9]/P0001 , \wishbone_rx_fifo_fifo_reg[3][0]/P0001 , \wishbone_rx_fifo_fifo_reg[3][10]/P0001 , \wishbone_rx_fifo_fifo_reg[3][11]/P0001 , \wishbone_rx_fifo_fifo_reg[3][12]/P0001 , \wishbone_rx_fifo_fifo_reg[3][13]/P0001 , \wishbone_rx_fifo_fifo_reg[3][14]/P0001 , \wishbone_rx_fifo_fifo_reg[3][15]/P0001 , \wishbone_rx_fifo_fifo_reg[3][16]/P0001 , \wishbone_rx_fifo_fifo_reg[3][17]/P0001 , \wishbone_rx_fifo_fifo_reg[3][18]/P0001 , \wishbone_rx_fifo_fifo_reg[3][19]/P0001 , \wishbone_rx_fifo_fifo_reg[3][1]/P0001 , \wishbone_rx_fifo_fifo_reg[3][20]/P0001 , \wishbone_rx_fifo_fifo_reg[3][21]/P0001 , \wishbone_rx_fifo_fifo_reg[3][22]/P0001 , \wishbone_rx_fifo_fifo_reg[3][23]/P0001 , \wishbone_rx_fifo_fifo_reg[3][24]/P0001 , \wishbone_rx_fifo_fifo_reg[3][25]/P0001 , \wishbone_rx_fifo_fifo_reg[3][26]/P0001 , \wishbone_rx_fifo_fifo_reg[3][27]/P0001 , \wishbone_rx_fifo_fifo_reg[3][28]/P0001 , \wishbone_rx_fifo_fifo_reg[3][29]/P0001 , \wishbone_rx_fifo_fifo_reg[3][2]/P0001 , \wishbone_rx_fifo_fifo_reg[3][30]/P0001 , \wishbone_rx_fifo_fifo_reg[3][31]/P0001 , \wishbone_rx_fifo_fifo_reg[3][3]/P0001 , \wishbone_rx_fifo_fifo_reg[3][4]/P0001 , \wishbone_rx_fifo_fifo_reg[3][5]/P0001 , \wishbone_rx_fifo_fifo_reg[3][6]/P0001 , \wishbone_rx_fifo_fifo_reg[3][7]/P0001 , \wishbone_rx_fifo_fifo_reg[3][8]/P0001 , \wishbone_rx_fifo_fifo_reg[3][9]/P0001 , \wishbone_rx_fifo_fifo_reg[4][0]/P0001 , \wishbone_rx_fifo_fifo_reg[4][10]/P0001 , \wishbone_rx_fifo_fifo_reg[4][11]/P0001 , \wishbone_rx_fifo_fifo_reg[4][12]/P0001 , \wishbone_rx_fifo_fifo_reg[4][13]/P0001 , \wishbone_rx_fifo_fifo_reg[4][14]/P0001 , \wishbone_rx_fifo_fifo_reg[4][15]/P0001 , \wishbone_rx_fifo_fifo_reg[4][16]/P0001 , \wishbone_rx_fifo_fifo_reg[4][17]/P0001 , \wishbone_rx_fifo_fifo_reg[4][18]/P0001 , \wishbone_rx_fifo_fifo_reg[4][19]/P0001 , \wishbone_rx_fifo_fifo_reg[4][1]/P0001 , \wishbone_rx_fifo_fifo_reg[4][20]/P0001 , \wishbone_rx_fifo_fifo_reg[4][21]/P0001 , \wishbone_rx_fifo_fifo_reg[4][22]/P0001 , \wishbone_rx_fifo_fifo_reg[4][23]/P0001 , \wishbone_rx_fifo_fifo_reg[4][24]/P0001 , \wishbone_rx_fifo_fifo_reg[4][25]/P0001 , \wishbone_rx_fifo_fifo_reg[4][26]/P0001 , \wishbone_rx_fifo_fifo_reg[4][27]/P0001 , \wishbone_rx_fifo_fifo_reg[4][28]/P0001 , \wishbone_rx_fifo_fifo_reg[4][29]/P0001 , \wishbone_rx_fifo_fifo_reg[4][2]/P0001 , \wishbone_rx_fifo_fifo_reg[4][30]/P0001 , \wishbone_rx_fifo_fifo_reg[4][31]/P0001 , \wishbone_rx_fifo_fifo_reg[4][3]/P0001 , \wishbone_rx_fifo_fifo_reg[4][4]/P0001 , \wishbone_rx_fifo_fifo_reg[4][5]/P0001 , \wishbone_rx_fifo_fifo_reg[4][6]/P0001 , \wishbone_rx_fifo_fifo_reg[4][7]/P0001 , \wishbone_rx_fifo_fifo_reg[4][8]/P0001 , \wishbone_rx_fifo_fifo_reg[4][9]/P0001 , \wishbone_rx_fifo_fifo_reg[5][0]/P0001 , \wishbone_rx_fifo_fifo_reg[5][10]/P0001 , \wishbone_rx_fifo_fifo_reg[5][11]/P0001 , \wishbone_rx_fifo_fifo_reg[5][12]/P0001 , \wishbone_rx_fifo_fifo_reg[5][13]/P0001 , \wishbone_rx_fifo_fifo_reg[5][14]/P0001 , \wishbone_rx_fifo_fifo_reg[5][15]/P0001 , \wishbone_rx_fifo_fifo_reg[5][16]/P0001 , \wishbone_rx_fifo_fifo_reg[5][17]/P0001 , \wishbone_rx_fifo_fifo_reg[5][18]/P0001 , \wishbone_rx_fifo_fifo_reg[5][19]/P0001 , \wishbone_rx_fifo_fifo_reg[5][1]/P0001 , \wishbone_rx_fifo_fifo_reg[5][20]/P0001 , \wishbone_rx_fifo_fifo_reg[5][21]/P0001 , \wishbone_rx_fifo_fifo_reg[5][22]/P0001 , \wishbone_rx_fifo_fifo_reg[5][23]/P0001 , \wishbone_rx_fifo_fifo_reg[5][24]/P0001 , \wishbone_rx_fifo_fifo_reg[5][25]/P0001 , \wishbone_rx_fifo_fifo_reg[5][26]/P0001 , \wishbone_rx_fifo_fifo_reg[5][27]/P0001 , \wishbone_rx_fifo_fifo_reg[5][28]/P0001 , \wishbone_rx_fifo_fifo_reg[5][29]/P0001 , \wishbone_rx_fifo_fifo_reg[5][2]/P0001 , \wishbone_rx_fifo_fifo_reg[5][30]/P0001 , \wishbone_rx_fifo_fifo_reg[5][31]/P0001 , \wishbone_rx_fifo_fifo_reg[5][3]/P0001 , \wishbone_rx_fifo_fifo_reg[5][4]/P0001 , \wishbone_rx_fifo_fifo_reg[5][5]/P0001 , \wishbone_rx_fifo_fifo_reg[5][6]/P0001 , \wishbone_rx_fifo_fifo_reg[5][7]/P0001 , \wishbone_rx_fifo_fifo_reg[5][8]/P0001 , \wishbone_rx_fifo_fifo_reg[5][9]/P0001 , \wishbone_rx_fifo_fifo_reg[6][0]/P0001 , \wishbone_rx_fifo_fifo_reg[6][10]/P0001 , \wishbone_rx_fifo_fifo_reg[6][11]/P0001 , \wishbone_rx_fifo_fifo_reg[6][12]/P0001 , \wishbone_rx_fifo_fifo_reg[6][13]/P0001 , \wishbone_rx_fifo_fifo_reg[6][14]/P0001 , \wishbone_rx_fifo_fifo_reg[6][15]/P0001 , \wishbone_rx_fifo_fifo_reg[6][16]/P0001 , \wishbone_rx_fifo_fifo_reg[6][17]/P0001 , \wishbone_rx_fifo_fifo_reg[6][18]/P0001 , \wishbone_rx_fifo_fifo_reg[6][19]/P0001 , \wishbone_rx_fifo_fifo_reg[6][1]/P0001 , \wishbone_rx_fifo_fifo_reg[6][20]/P0001 , \wishbone_rx_fifo_fifo_reg[6][21]/P0001 , \wishbone_rx_fifo_fifo_reg[6][22]/P0001 , \wishbone_rx_fifo_fifo_reg[6][23]/P0001 , \wishbone_rx_fifo_fifo_reg[6][24]/P0001 , \wishbone_rx_fifo_fifo_reg[6][25]/P0001 , \wishbone_rx_fifo_fifo_reg[6][26]/P0001 , \wishbone_rx_fifo_fifo_reg[6][27]/P0001 , \wishbone_rx_fifo_fifo_reg[6][28]/P0001 , \wishbone_rx_fifo_fifo_reg[6][29]/P0001 , \wishbone_rx_fifo_fifo_reg[6][2]/P0001 , \wishbone_rx_fifo_fifo_reg[6][30]/P0001 , \wishbone_rx_fifo_fifo_reg[6][31]/P0001 , \wishbone_rx_fifo_fifo_reg[6][3]/P0001 , \wishbone_rx_fifo_fifo_reg[6][4]/P0001 , \wishbone_rx_fifo_fifo_reg[6][5]/P0001 , \wishbone_rx_fifo_fifo_reg[6][6]/P0001 , \wishbone_rx_fifo_fifo_reg[6][7]/P0001 , \wishbone_rx_fifo_fifo_reg[6][8]/P0001 , \wishbone_rx_fifo_fifo_reg[6][9]/P0001 , \wishbone_rx_fifo_fifo_reg[7][0]/P0001 , \wishbone_rx_fifo_fifo_reg[7][10]/P0001 , \wishbone_rx_fifo_fifo_reg[7][11]/P0001 , \wishbone_rx_fifo_fifo_reg[7][12]/P0001 , \wishbone_rx_fifo_fifo_reg[7][13]/P0001 , \wishbone_rx_fifo_fifo_reg[7][14]/P0001 , \wishbone_rx_fifo_fifo_reg[7][15]/P0001 , \wishbone_rx_fifo_fifo_reg[7][16]/P0001 , \wishbone_rx_fifo_fifo_reg[7][17]/P0001 , \wishbone_rx_fifo_fifo_reg[7][18]/P0001 , \wishbone_rx_fifo_fifo_reg[7][19]/P0001 , \wishbone_rx_fifo_fifo_reg[7][1]/P0001 , \wishbone_rx_fifo_fifo_reg[7][20]/P0001 , \wishbone_rx_fifo_fifo_reg[7][21]/P0001 , \wishbone_rx_fifo_fifo_reg[7][22]/P0001 , \wishbone_rx_fifo_fifo_reg[7][23]/P0001 , \wishbone_rx_fifo_fifo_reg[7][24]/P0001 , \wishbone_rx_fifo_fifo_reg[7][25]/P0001 , \wishbone_rx_fifo_fifo_reg[7][26]/P0001 , \wishbone_rx_fifo_fifo_reg[7][27]/P0001 , \wishbone_rx_fifo_fifo_reg[7][28]/P0001 , \wishbone_rx_fifo_fifo_reg[7][29]/P0001 , \wishbone_rx_fifo_fifo_reg[7][2]/P0001 , \wishbone_rx_fifo_fifo_reg[7][30]/P0001 , \wishbone_rx_fifo_fifo_reg[7][31]/P0001 , \wishbone_rx_fifo_fifo_reg[7][3]/P0001 , \wishbone_rx_fifo_fifo_reg[7][4]/P0001 , \wishbone_rx_fifo_fifo_reg[7][5]/P0001 , \wishbone_rx_fifo_fifo_reg[7][6]/P0001 , \wishbone_rx_fifo_fifo_reg[7][7]/P0001 , \wishbone_rx_fifo_fifo_reg[7][8]/P0001 , \wishbone_rx_fifo_fifo_reg[7][9]/P0001 , \wishbone_rx_fifo_fifo_reg[8][0]/P0001 , \wishbone_rx_fifo_fifo_reg[8][10]/P0001 , \wishbone_rx_fifo_fifo_reg[8][11]/P0001 , \wishbone_rx_fifo_fifo_reg[8][12]/P0001 , \wishbone_rx_fifo_fifo_reg[8][13]/P0001 , \wishbone_rx_fifo_fifo_reg[8][14]/P0001 , \wishbone_rx_fifo_fifo_reg[8][15]/P0001 , \wishbone_rx_fifo_fifo_reg[8][16]/P0001 , \wishbone_rx_fifo_fifo_reg[8][17]/P0001 , \wishbone_rx_fifo_fifo_reg[8][18]/P0001 , \wishbone_rx_fifo_fifo_reg[8][19]/P0001 , \wishbone_rx_fifo_fifo_reg[8][1]/P0001 , \wishbone_rx_fifo_fifo_reg[8][20]/P0001 , \wishbone_rx_fifo_fifo_reg[8][21]/P0001 , \wishbone_rx_fifo_fifo_reg[8][22]/P0001 , \wishbone_rx_fifo_fifo_reg[8][23]/P0001 , \wishbone_rx_fifo_fifo_reg[8][24]/P0001 , \wishbone_rx_fifo_fifo_reg[8][25]/P0001 , \wishbone_rx_fifo_fifo_reg[8][26]/P0001 , \wishbone_rx_fifo_fifo_reg[8][27]/P0001 , \wishbone_rx_fifo_fifo_reg[8][28]/P0001 , \wishbone_rx_fifo_fifo_reg[8][29]/P0001 , \wishbone_rx_fifo_fifo_reg[8][2]/P0001 , \wishbone_rx_fifo_fifo_reg[8][30]/P0001 , \wishbone_rx_fifo_fifo_reg[8][31]/P0001 , \wishbone_rx_fifo_fifo_reg[8][3]/P0001 , \wishbone_rx_fifo_fifo_reg[8][4]/P0001 , \wishbone_rx_fifo_fifo_reg[8][5]/P0001 , \wishbone_rx_fifo_fifo_reg[8][6]/P0001 , \wishbone_rx_fifo_fifo_reg[8][7]/P0001 , \wishbone_rx_fifo_fifo_reg[8][8]/P0001 , \wishbone_rx_fifo_fifo_reg[8][9]/P0001 , \wishbone_rx_fifo_fifo_reg[9][0]/P0001 , \wishbone_rx_fifo_fifo_reg[9][10]/P0001 , \wishbone_rx_fifo_fifo_reg[9][11]/P0001 , \wishbone_rx_fifo_fifo_reg[9][12]/P0001 , \wishbone_rx_fifo_fifo_reg[9][13]/P0001 , \wishbone_rx_fifo_fifo_reg[9][14]/P0001 , \wishbone_rx_fifo_fifo_reg[9][15]/P0001 , \wishbone_rx_fifo_fifo_reg[9][16]/P0001 , \wishbone_rx_fifo_fifo_reg[9][17]/P0001 , \wishbone_rx_fifo_fifo_reg[9][18]/P0001 , \wishbone_rx_fifo_fifo_reg[9][19]/P0001 , \wishbone_rx_fifo_fifo_reg[9][1]/P0001 , \wishbone_rx_fifo_fifo_reg[9][20]/P0001 , \wishbone_rx_fifo_fifo_reg[9][21]/P0001 , \wishbone_rx_fifo_fifo_reg[9][22]/P0001 , \wishbone_rx_fifo_fifo_reg[9][23]/P0001 , \wishbone_rx_fifo_fifo_reg[9][24]/P0001 , \wishbone_rx_fifo_fifo_reg[9][25]/P0001 , \wishbone_rx_fifo_fifo_reg[9][26]/P0001 , \wishbone_rx_fifo_fifo_reg[9][27]/P0001 , \wishbone_rx_fifo_fifo_reg[9][28]/P0001 , \wishbone_rx_fifo_fifo_reg[9][29]/P0001 , \wishbone_rx_fifo_fifo_reg[9][2]/P0001 , \wishbone_rx_fifo_fifo_reg[9][30]/P0001 , \wishbone_rx_fifo_fifo_reg[9][31]/P0001 , \wishbone_rx_fifo_fifo_reg[9][3]/P0001 , \wishbone_rx_fifo_fifo_reg[9][4]/P0001 , \wishbone_rx_fifo_fifo_reg[9][5]/P0001 , \wishbone_rx_fifo_fifo_reg[9][6]/P0001 , \wishbone_rx_fifo_fifo_reg[9][7]/P0001 , \wishbone_rx_fifo_fifo_reg[9][8]/P0001 , \wishbone_rx_fifo_fifo_reg[9][9]/P0001 , \wishbone_rx_fifo_read_pointer_reg[0]/NET0131 , \wishbone_rx_fifo_read_pointer_reg[1]/NET0131 , \wishbone_rx_fifo_read_pointer_reg[2]/NET0131 , \wishbone_rx_fifo_read_pointer_reg[3]/NET0131 , \wishbone_rx_fifo_write_pointer_reg[0]/NET0131 , \wishbone_rx_fifo_write_pointer_reg[1]/NET0131 , \wishbone_rx_fifo_write_pointer_reg[2]/NET0131 , \wishbone_rx_fifo_write_pointer_reg[3]/NET0131 , \wishbone_tx_burst_cnt_reg[0]/NET0131 , \wishbone_tx_burst_cnt_reg[1]/NET0131 , \wishbone_tx_burst_cnt_reg[2]/NET0131 , \wishbone_tx_burst_en_reg/NET0131 , \wishbone_tx_fifo_cnt_reg[0]/NET0131 , \wishbone_tx_fifo_cnt_reg[1]/NET0131 , \wishbone_tx_fifo_cnt_reg[2]/NET0131 , \wishbone_tx_fifo_cnt_reg[3]/NET0131 , \wishbone_tx_fifo_cnt_reg[4]/NET0131 , \wishbone_tx_fifo_data_out_reg[0]/P0001 , \wishbone_tx_fifo_data_out_reg[10]/P0001 , \wishbone_tx_fifo_data_out_reg[11]/P0001 , \wishbone_tx_fifo_data_out_reg[12]/P0001 , \wishbone_tx_fifo_data_out_reg[13]/P0001 , \wishbone_tx_fifo_data_out_reg[14]/P0001 , \wishbone_tx_fifo_data_out_reg[15]/P0001 , \wishbone_tx_fifo_data_out_reg[16]/P0001 , \wishbone_tx_fifo_data_out_reg[17]/P0001 , \wishbone_tx_fifo_data_out_reg[18]/P0001 , \wishbone_tx_fifo_data_out_reg[19]/P0001 , \wishbone_tx_fifo_data_out_reg[1]/P0001 , \wishbone_tx_fifo_data_out_reg[20]/P0001 , \wishbone_tx_fifo_data_out_reg[21]/P0001 , \wishbone_tx_fifo_data_out_reg[22]/P0001 , \wishbone_tx_fifo_data_out_reg[23]/P0001 , \wishbone_tx_fifo_data_out_reg[24]/P0001 , \wishbone_tx_fifo_data_out_reg[25]/P0001 , \wishbone_tx_fifo_data_out_reg[26]/P0001 , \wishbone_tx_fifo_data_out_reg[27]/P0001 , \wishbone_tx_fifo_data_out_reg[28]/P0001 , \wishbone_tx_fifo_data_out_reg[29]/P0001 , \wishbone_tx_fifo_data_out_reg[2]/P0001 , \wishbone_tx_fifo_data_out_reg[30]/P0001 , \wishbone_tx_fifo_data_out_reg[31]/P0001 , \wishbone_tx_fifo_data_out_reg[3]/P0001 , \wishbone_tx_fifo_data_out_reg[4]/P0001 , \wishbone_tx_fifo_data_out_reg[5]/P0001 , \wishbone_tx_fifo_data_out_reg[6]/P0001 , \wishbone_tx_fifo_data_out_reg[7]/P0001 , \wishbone_tx_fifo_data_out_reg[8]/P0001 , \wishbone_tx_fifo_data_out_reg[9]/P0001 , \wishbone_tx_fifo_fifo_reg[0][0]/P0001 , \wishbone_tx_fifo_fifo_reg[0][10]/P0001 , \wishbone_tx_fifo_fifo_reg[0][11]/P0001 , \wishbone_tx_fifo_fifo_reg[0][12]/P0001 , \wishbone_tx_fifo_fifo_reg[0][13]/P0001 , \wishbone_tx_fifo_fifo_reg[0][14]/P0001 , \wishbone_tx_fifo_fifo_reg[0][15]/P0001 , \wishbone_tx_fifo_fifo_reg[0][16]/P0001 , \wishbone_tx_fifo_fifo_reg[0][17]/P0001 , \wishbone_tx_fifo_fifo_reg[0][18]/P0001 , \wishbone_tx_fifo_fifo_reg[0][19]/P0001 , \wishbone_tx_fifo_fifo_reg[0][1]/P0001 , \wishbone_tx_fifo_fifo_reg[0][20]/P0001 , \wishbone_tx_fifo_fifo_reg[0][21]/P0001 , \wishbone_tx_fifo_fifo_reg[0][22]/P0001 , \wishbone_tx_fifo_fifo_reg[0][23]/P0001 , \wishbone_tx_fifo_fifo_reg[0][24]/P0001 , \wishbone_tx_fifo_fifo_reg[0][25]/P0001 , \wishbone_tx_fifo_fifo_reg[0][26]/P0001 , \wishbone_tx_fifo_fifo_reg[0][27]/P0001 , \wishbone_tx_fifo_fifo_reg[0][28]/P0001 , \wishbone_tx_fifo_fifo_reg[0][29]/P0001 , \wishbone_tx_fifo_fifo_reg[0][2]/P0001 , \wishbone_tx_fifo_fifo_reg[0][30]/P0001 , \wishbone_tx_fifo_fifo_reg[0][31]/P0001 , \wishbone_tx_fifo_fifo_reg[0][3]/P0001 , \wishbone_tx_fifo_fifo_reg[0][4]/P0001 , \wishbone_tx_fifo_fifo_reg[0][5]/P0001 , \wishbone_tx_fifo_fifo_reg[0][6]/P0001 , \wishbone_tx_fifo_fifo_reg[0][7]/P0001 , \wishbone_tx_fifo_fifo_reg[0][8]/P0001 , \wishbone_tx_fifo_fifo_reg[0][9]/P0001 , \wishbone_tx_fifo_fifo_reg[10][0]/P0001 , \wishbone_tx_fifo_fifo_reg[10][10]/P0001 , \wishbone_tx_fifo_fifo_reg[10][11]/P0001 , \wishbone_tx_fifo_fifo_reg[10][12]/P0001 , \wishbone_tx_fifo_fifo_reg[10][13]/P0001 , \wishbone_tx_fifo_fifo_reg[10][14]/P0001 , \wishbone_tx_fifo_fifo_reg[10][15]/P0001 , \wishbone_tx_fifo_fifo_reg[10][16]/P0001 , \wishbone_tx_fifo_fifo_reg[10][17]/P0001 , \wishbone_tx_fifo_fifo_reg[10][18]/P0001 , \wishbone_tx_fifo_fifo_reg[10][19]/P0001 , \wishbone_tx_fifo_fifo_reg[10][1]/P0001 , \wishbone_tx_fifo_fifo_reg[10][20]/P0001 , \wishbone_tx_fifo_fifo_reg[10][21]/P0001 , \wishbone_tx_fifo_fifo_reg[10][22]/P0001 , \wishbone_tx_fifo_fifo_reg[10][23]/P0001 , \wishbone_tx_fifo_fifo_reg[10][24]/P0001 , \wishbone_tx_fifo_fifo_reg[10][25]/P0001 , \wishbone_tx_fifo_fifo_reg[10][26]/P0001 , \wishbone_tx_fifo_fifo_reg[10][27]/P0001 , \wishbone_tx_fifo_fifo_reg[10][28]/P0001 , \wishbone_tx_fifo_fifo_reg[10][29]/P0001 , \wishbone_tx_fifo_fifo_reg[10][2]/P0001 , \wishbone_tx_fifo_fifo_reg[10][30]/P0001 , \wishbone_tx_fifo_fifo_reg[10][31]/P0001 , \wishbone_tx_fifo_fifo_reg[10][3]/P0001 , \wishbone_tx_fifo_fifo_reg[10][4]/P0001 , \wishbone_tx_fifo_fifo_reg[10][5]/P0001 , \wishbone_tx_fifo_fifo_reg[10][6]/P0001 , \wishbone_tx_fifo_fifo_reg[10][7]/P0001 , \wishbone_tx_fifo_fifo_reg[10][8]/P0001 , \wishbone_tx_fifo_fifo_reg[10][9]/P0001 , \wishbone_tx_fifo_fifo_reg[11][0]/P0001 , \wishbone_tx_fifo_fifo_reg[11][10]/P0001 , \wishbone_tx_fifo_fifo_reg[11][11]/P0001 , \wishbone_tx_fifo_fifo_reg[11][12]/P0001 , \wishbone_tx_fifo_fifo_reg[11][13]/P0001 , \wishbone_tx_fifo_fifo_reg[11][14]/P0001 , \wishbone_tx_fifo_fifo_reg[11][15]/P0001 , \wishbone_tx_fifo_fifo_reg[11][16]/P0001 , \wishbone_tx_fifo_fifo_reg[11][17]/P0001 , \wishbone_tx_fifo_fifo_reg[11][18]/P0001 , \wishbone_tx_fifo_fifo_reg[11][19]/P0001 , \wishbone_tx_fifo_fifo_reg[11][1]/P0001 , \wishbone_tx_fifo_fifo_reg[11][20]/P0001 , \wishbone_tx_fifo_fifo_reg[11][21]/P0001 , \wishbone_tx_fifo_fifo_reg[11][22]/P0001 , \wishbone_tx_fifo_fifo_reg[11][23]/P0001 , \wishbone_tx_fifo_fifo_reg[11][24]/P0001 , \wishbone_tx_fifo_fifo_reg[11][25]/P0001 , \wishbone_tx_fifo_fifo_reg[11][26]/P0001 , \wishbone_tx_fifo_fifo_reg[11][27]/P0001 , \wishbone_tx_fifo_fifo_reg[11][28]/P0001 , \wishbone_tx_fifo_fifo_reg[11][29]/P0001 , \wishbone_tx_fifo_fifo_reg[11][2]/P0001 , \wishbone_tx_fifo_fifo_reg[11][30]/P0001 , \wishbone_tx_fifo_fifo_reg[11][31]/P0001 , \wishbone_tx_fifo_fifo_reg[11][3]/P0001 , \wishbone_tx_fifo_fifo_reg[11][4]/P0001 , \wishbone_tx_fifo_fifo_reg[11][5]/P0001 , \wishbone_tx_fifo_fifo_reg[11][6]/P0001 , \wishbone_tx_fifo_fifo_reg[11][7]/P0001 , \wishbone_tx_fifo_fifo_reg[11][8]/P0001 , \wishbone_tx_fifo_fifo_reg[11][9]/P0001 , \wishbone_tx_fifo_fifo_reg[12][0]/P0001 , \wishbone_tx_fifo_fifo_reg[12][10]/P0001 , \wishbone_tx_fifo_fifo_reg[12][11]/P0001 , \wishbone_tx_fifo_fifo_reg[12][12]/P0001 , \wishbone_tx_fifo_fifo_reg[12][13]/P0001 , \wishbone_tx_fifo_fifo_reg[12][14]/P0001 , \wishbone_tx_fifo_fifo_reg[12][15]/P0001 , \wishbone_tx_fifo_fifo_reg[12][16]/P0001 , \wishbone_tx_fifo_fifo_reg[12][17]/P0001 , \wishbone_tx_fifo_fifo_reg[12][18]/P0001 , \wishbone_tx_fifo_fifo_reg[12][19]/P0001 , \wishbone_tx_fifo_fifo_reg[12][1]/P0001 , \wishbone_tx_fifo_fifo_reg[12][20]/P0001 , \wishbone_tx_fifo_fifo_reg[12][21]/P0001 , \wishbone_tx_fifo_fifo_reg[12][22]/P0001 , \wishbone_tx_fifo_fifo_reg[12][23]/P0001 , \wishbone_tx_fifo_fifo_reg[12][24]/P0001 , \wishbone_tx_fifo_fifo_reg[12][25]/P0001 , \wishbone_tx_fifo_fifo_reg[12][26]/P0001 , \wishbone_tx_fifo_fifo_reg[12][27]/P0001 , \wishbone_tx_fifo_fifo_reg[12][28]/P0001 , \wishbone_tx_fifo_fifo_reg[12][29]/P0001 , \wishbone_tx_fifo_fifo_reg[12][2]/P0001 , \wishbone_tx_fifo_fifo_reg[12][30]/P0001 , \wishbone_tx_fifo_fifo_reg[12][31]/P0001 , \wishbone_tx_fifo_fifo_reg[12][3]/P0001 , \wishbone_tx_fifo_fifo_reg[12][4]/P0001 , \wishbone_tx_fifo_fifo_reg[12][5]/P0001 , \wishbone_tx_fifo_fifo_reg[12][6]/P0001 , \wishbone_tx_fifo_fifo_reg[12][7]/P0001 , \wishbone_tx_fifo_fifo_reg[12][8]/P0001 , \wishbone_tx_fifo_fifo_reg[12][9]/P0001 , \wishbone_tx_fifo_fifo_reg[13][0]/P0001 , \wishbone_tx_fifo_fifo_reg[13][10]/P0001 , \wishbone_tx_fifo_fifo_reg[13][11]/P0001 , \wishbone_tx_fifo_fifo_reg[13][12]/P0001 , \wishbone_tx_fifo_fifo_reg[13][13]/P0001 , \wishbone_tx_fifo_fifo_reg[13][14]/P0001 , \wishbone_tx_fifo_fifo_reg[13][15]/P0001 , \wishbone_tx_fifo_fifo_reg[13][16]/P0001 , \wishbone_tx_fifo_fifo_reg[13][17]/P0001 , \wishbone_tx_fifo_fifo_reg[13][18]/P0001 , \wishbone_tx_fifo_fifo_reg[13][19]/P0001 , \wishbone_tx_fifo_fifo_reg[13][1]/P0001 , \wishbone_tx_fifo_fifo_reg[13][20]/P0001 , \wishbone_tx_fifo_fifo_reg[13][21]/P0001 , \wishbone_tx_fifo_fifo_reg[13][22]/P0001 , \wishbone_tx_fifo_fifo_reg[13][23]/P0001 , \wishbone_tx_fifo_fifo_reg[13][24]/P0001 , \wishbone_tx_fifo_fifo_reg[13][25]/P0001 , \wishbone_tx_fifo_fifo_reg[13][26]/P0001 , \wishbone_tx_fifo_fifo_reg[13][27]/P0001 , \wishbone_tx_fifo_fifo_reg[13][28]/P0001 , \wishbone_tx_fifo_fifo_reg[13][29]/P0001 , \wishbone_tx_fifo_fifo_reg[13][2]/P0001 , \wishbone_tx_fifo_fifo_reg[13][30]/P0001 , \wishbone_tx_fifo_fifo_reg[13][31]/P0001 , \wishbone_tx_fifo_fifo_reg[13][3]/P0001 , \wishbone_tx_fifo_fifo_reg[13][4]/P0001 , \wishbone_tx_fifo_fifo_reg[13][5]/P0001 , \wishbone_tx_fifo_fifo_reg[13][6]/P0001 , \wishbone_tx_fifo_fifo_reg[13][7]/P0001 , \wishbone_tx_fifo_fifo_reg[13][8]/P0001 , \wishbone_tx_fifo_fifo_reg[13][9]/P0001 , \wishbone_tx_fifo_fifo_reg[14][0]/P0001 , \wishbone_tx_fifo_fifo_reg[14][10]/P0001 , \wishbone_tx_fifo_fifo_reg[14][11]/P0001 , \wishbone_tx_fifo_fifo_reg[14][12]/P0001 , \wishbone_tx_fifo_fifo_reg[14][13]/P0001 , \wishbone_tx_fifo_fifo_reg[14][14]/P0001 , \wishbone_tx_fifo_fifo_reg[14][15]/P0001 , \wishbone_tx_fifo_fifo_reg[14][16]/P0001 , \wishbone_tx_fifo_fifo_reg[14][17]/P0001 , \wishbone_tx_fifo_fifo_reg[14][18]/P0001 , \wishbone_tx_fifo_fifo_reg[14][19]/P0001 , \wishbone_tx_fifo_fifo_reg[14][1]/P0001 , \wishbone_tx_fifo_fifo_reg[14][20]/P0001 , \wishbone_tx_fifo_fifo_reg[14][21]/P0001 , \wishbone_tx_fifo_fifo_reg[14][22]/P0001 , \wishbone_tx_fifo_fifo_reg[14][23]/P0001 , \wishbone_tx_fifo_fifo_reg[14][24]/P0001 , \wishbone_tx_fifo_fifo_reg[14][25]/P0001 , \wishbone_tx_fifo_fifo_reg[14][26]/P0001 , \wishbone_tx_fifo_fifo_reg[14][27]/P0001 , \wishbone_tx_fifo_fifo_reg[14][28]/P0001 , \wishbone_tx_fifo_fifo_reg[14][29]/P0001 , \wishbone_tx_fifo_fifo_reg[14][2]/P0001 , \wishbone_tx_fifo_fifo_reg[14][30]/P0001 , \wishbone_tx_fifo_fifo_reg[14][31]/P0001 , \wishbone_tx_fifo_fifo_reg[14][3]/P0001 , \wishbone_tx_fifo_fifo_reg[14][4]/P0001 , \wishbone_tx_fifo_fifo_reg[14][5]/P0001 , \wishbone_tx_fifo_fifo_reg[14][6]/P0001 , \wishbone_tx_fifo_fifo_reg[14][7]/P0001 , \wishbone_tx_fifo_fifo_reg[14][8]/P0001 , \wishbone_tx_fifo_fifo_reg[14][9]/P0001 , \wishbone_tx_fifo_fifo_reg[15][0]/P0001 , \wishbone_tx_fifo_fifo_reg[15][10]/P0001 , \wishbone_tx_fifo_fifo_reg[15][11]/P0001 , \wishbone_tx_fifo_fifo_reg[15][12]/P0001 , \wishbone_tx_fifo_fifo_reg[15][13]/P0001 , \wishbone_tx_fifo_fifo_reg[15][14]/P0001 , \wishbone_tx_fifo_fifo_reg[15][15]/P0001 , \wishbone_tx_fifo_fifo_reg[15][16]/P0001 , \wishbone_tx_fifo_fifo_reg[15][17]/P0001 , \wishbone_tx_fifo_fifo_reg[15][18]/P0001 , \wishbone_tx_fifo_fifo_reg[15][19]/P0001 , \wishbone_tx_fifo_fifo_reg[15][1]/P0001 , \wishbone_tx_fifo_fifo_reg[15][20]/P0001 , \wishbone_tx_fifo_fifo_reg[15][21]/P0001 , \wishbone_tx_fifo_fifo_reg[15][22]/P0001 , \wishbone_tx_fifo_fifo_reg[15][23]/P0001 , \wishbone_tx_fifo_fifo_reg[15][24]/P0001 , \wishbone_tx_fifo_fifo_reg[15][25]/P0001 , \wishbone_tx_fifo_fifo_reg[15][26]/P0001 , \wishbone_tx_fifo_fifo_reg[15][27]/P0001 , \wishbone_tx_fifo_fifo_reg[15][28]/P0001 , \wishbone_tx_fifo_fifo_reg[15][29]/P0001 , \wishbone_tx_fifo_fifo_reg[15][2]/P0001 , \wishbone_tx_fifo_fifo_reg[15][30]/P0001 , \wishbone_tx_fifo_fifo_reg[15][31]/P0001 , \wishbone_tx_fifo_fifo_reg[15][3]/P0001 , \wishbone_tx_fifo_fifo_reg[15][4]/P0001 , \wishbone_tx_fifo_fifo_reg[15][5]/P0001 , \wishbone_tx_fifo_fifo_reg[15][6]/P0001 , \wishbone_tx_fifo_fifo_reg[15][7]/P0001 , \wishbone_tx_fifo_fifo_reg[15][8]/P0001 , \wishbone_tx_fifo_fifo_reg[15][9]/P0001 , \wishbone_tx_fifo_fifo_reg[1][0]/P0001 , \wishbone_tx_fifo_fifo_reg[1][10]/P0001 , \wishbone_tx_fifo_fifo_reg[1][11]/P0001 , \wishbone_tx_fifo_fifo_reg[1][12]/P0001 , \wishbone_tx_fifo_fifo_reg[1][13]/P0001 , \wishbone_tx_fifo_fifo_reg[1][14]/P0001 , \wishbone_tx_fifo_fifo_reg[1][15]/P0001 , \wishbone_tx_fifo_fifo_reg[1][16]/P0001 , \wishbone_tx_fifo_fifo_reg[1][17]/P0001 , \wishbone_tx_fifo_fifo_reg[1][18]/P0001 , \wishbone_tx_fifo_fifo_reg[1][19]/P0001 , \wishbone_tx_fifo_fifo_reg[1][1]/P0001 , \wishbone_tx_fifo_fifo_reg[1][20]/P0001 , \wishbone_tx_fifo_fifo_reg[1][21]/P0001 , \wishbone_tx_fifo_fifo_reg[1][22]/P0001 , \wishbone_tx_fifo_fifo_reg[1][23]/P0001 , \wishbone_tx_fifo_fifo_reg[1][24]/P0001 , \wishbone_tx_fifo_fifo_reg[1][25]/P0001 , \wishbone_tx_fifo_fifo_reg[1][26]/P0001 , \wishbone_tx_fifo_fifo_reg[1][27]/P0001 , \wishbone_tx_fifo_fifo_reg[1][28]/P0001 , \wishbone_tx_fifo_fifo_reg[1][29]/P0001 , \wishbone_tx_fifo_fifo_reg[1][2]/P0001 , \wishbone_tx_fifo_fifo_reg[1][30]/P0001 , \wishbone_tx_fifo_fifo_reg[1][31]/P0001 , \wishbone_tx_fifo_fifo_reg[1][3]/P0001 , \wishbone_tx_fifo_fifo_reg[1][4]/P0001 , \wishbone_tx_fifo_fifo_reg[1][5]/P0001 , \wishbone_tx_fifo_fifo_reg[1][6]/P0001 , \wishbone_tx_fifo_fifo_reg[1][7]/P0001 , \wishbone_tx_fifo_fifo_reg[1][8]/P0001 , \wishbone_tx_fifo_fifo_reg[1][9]/P0001 , \wishbone_tx_fifo_fifo_reg[2][0]/P0001 , \wishbone_tx_fifo_fifo_reg[2][10]/P0001 , \wishbone_tx_fifo_fifo_reg[2][11]/P0001 , \wishbone_tx_fifo_fifo_reg[2][12]/P0001 , \wishbone_tx_fifo_fifo_reg[2][13]/P0001 , \wishbone_tx_fifo_fifo_reg[2][14]/P0001 , \wishbone_tx_fifo_fifo_reg[2][15]/P0001 , \wishbone_tx_fifo_fifo_reg[2][16]/P0001 , \wishbone_tx_fifo_fifo_reg[2][17]/P0001 , \wishbone_tx_fifo_fifo_reg[2][18]/P0001 , \wishbone_tx_fifo_fifo_reg[2][19]/P0001 , \wishbone_tx_fifo_fifo_reg[2][1]/P0001 , \wishbone_tx_fifo_fifo_reg[2][20]/P0001 , \wishbone_tx_fifo_fifo_reg[2][21]/P0001 , \wishbone_tx_fifo_fifo_reg[2][22]/P0001 , \wishbone_tx_fifo_fifo_reg[2][23]/P0001 , \wishbone_tx_fifo_fifo_reg[2][24]/P0001 , \wishbone_tx_fifo_fifo_reg[2][25]/P0001 , \wishbone_tx_fifo_fifo_reg[2][26]/P0001 , \wishbone_tx_fifo_fifo_reg[2][27]/P0001 , \wishbone_tx_fifo_fifo_reg[2][28]/P0001 , \wishbone_tx_fifo_fifo_reg[2][29]/P0001 , \wishbone_tx_fifo_fifo_reg[2][2]/P0001 , \wishbone_tx_fifo_fifo_reg[2][30]/P0001 , \wishbone_tx_fifo_fifo_reg[2][31]/P0001 , \wishbone_tx_fifo_fifo_reg[2][3]/P0001 , \wishbone_tx_fifo_fifo_reg[2][4]/P0001 , \wishbone_tx_fifo_fifo_reg[2][5]/P0001 , \wishbone_tx_fifo_fifo_reg[2][6]/P0001 , \wishbone_tx_fifo_fifo_reg[2][7]/P0001 , \wishbone_tx_fifo_fifo_reg[2][8]/P0001 , \wishbone_tx_fifo_fifo_reg[2][9]/P0001 , \wishbone_tx_fifo_fifo_reg[3][0]/P0001 , \wishbone_tx_fifo_fifo_reg[3][10]/P0001 , \wishbone_tx_fifo_fifo_reg[3][11]/P0001 , \wishbone_tx_fifo_fifo_reg[3][12]/P0001 , \wishbone_tx_fifo_fifo_reg[3][13]/P0001 , \wishbone_tx_fifo_fifo_reg[3][14]/P0001 , \wishbone_tx_fifo_fifo_reg[3][15]/P0001 , \wishbone_tx_fifo_fifo_reg[3][16]/P0001 , \wishbone_tx_fifo_fifo_reg[3][17]/P0001 , \wishbone_tx_fifo_fifo_reg[3][18]/P0001 , \wishbone_tx_fifo_fifo_reg[3][19]/P0001 , \wishbone_tx_fifo_fifo_reg[3][1]/P0001 , \wishbone_tx_fifo_fifo_reg[3][20]/P0001 , \wishbone_tx_fifo_fifo_reg[3][21]/P0001 , \wishbone_tx_fifo_fifo_reg[3][22]/P0001 , \wishbone_tx_fifo_fifo_reg[3][23]/P0001 , \wishbone_tx_fifo_fifo_reg[3][24]/P0001 , \wishbone_tx_fifo_fifo_reg[3][25]/P0001 , \wishbone_tx_fifo_fifo_reg[3][26]/P0001 , \wishbone_tx_fifo_fifo_reg[3][27]/P0001 , \wishbone_tx_fifo_fifo_reg[3][28]/P0001 , \wishbone_tx_fifo_fifo_reg[3][29]/P0001 , \wishbone_tx_fifo_fifo_reg[3][2]/P0001 , \wishbone_tx_fifo_fifo_reg[3][30]/P0001 , \wishbone_tx_fifo_fifo_reg[3][31]/P0001 , \wishbone_tx_fifo_fifo_reg[3][3]/P0001 , \wishbone_tx_fifo_fifo_reg[3][4]/P0001 , \wishbone_tx_fifo_fifo_reg[3][5]/P0001 , \wishbone_tx_fifo_fifo_reg[3][6]/P0001 , \wishbone_tx_fifo_fifo_reg[3][7]/P0001 , \wishbone_tx_fifo_fifo_reg[3][8]/P0001 , \wishbone_tx_fifo_fifo_reg[3][9]/P0001 , \wishbone_tx_fifo_fifo_reg[4][0]/P0001 , \wishbone_tx_fifo_fifo_reg[4][10]/P0001 , \wishbone_tx_fifo_fifo_reg[4][11]/P0001 , \wishbone_tx_fifo_fifo_reg[4][12]/P0001 , \wishbone_tx_fifo_fifo_reg[4][13]/P0001 , \wishbone_tx_fifo_fifo_reg[4][14]/P0001 , \wishbone_tx_fifo_fifo_reg[4][15]/P0001 , \wishbone_tx_fifo_fifo_reg[4][16]/P0001 , \wishbone_tx_fifo_fifo_reg[4][17]/P0001 , \wishbone_tx_fifo_fifo_reg[4][18]/P0001 , \wishbone_tx_fifo_fifo_reg[4][19]/P0001 , \wishbone_tx_fifo_fifo_reg[4][1]/P0001 , \wishbone_tx_fifo_fifo_reg[4][20]/P0001 , \wishbone_tx_fifo_fifo_reg[4][21]/P0001 , \wishbone_tx_fifo_fifo_reg[4][22]/P0001 , \wishbone_tx_fifo_fifo_reg[4][23]/P0001 , \wishbone_tx_fifo_fifo_reg[4][24]/P0001 , \wishbone_tx_fifo_fifo_reg[4][25]/P0001 , \wishbone_tx_fifo_fifo_reg[4][26]/P0001 , \wishbone_tx_fifo_fifo_reg[4][27]/P0001 , \wishbone_tx_fifo_fifo_reg[4][28]/P0001 , \wishbone_tx_fifo_fifo_reg[4][29]/P0001 , \wishbone_tx_fifo_fifo_reg[4][2]/P0001 , \wishbone_tx_fifo_fifo_reg[4][30]/P0001 , \wishbone_tx_fifo_fifo_reg[4][31]/P0001 , \wishbone_tx_fifo_fifo_reg[4][3]/P0001 , \wishbone_tx_fifo_fifo_reg[4][4]/P0001 , \wishbone_tx_fifo_fifo_reg[4][5]/P0001 , \wishbone_tx_fifo_fifo_reg[4][6]/P0001 , \wishbone_tx_fifo_fifo_reg[4][7]/P0001 , \wishbone_tx_fifo_fifo_reg[4][8]/P0001 , \wishbone_tx_fifo_fifo_reg[4][9]/P0001 , \wishbone_tx_fifo_fifo_reg[5][0]/P0001 , \wishbone_tx_fifo_fifo_reg[5][10]/P0001 , \wishbone_tx_fifo_fifo_reg[5][11]/P0001 , \wishbone_tx_fifo_fifo_reg[5][12]/P0001 , \wishbone_tx_fifo_fifo_reg[5][13]/P0001 , \wishbone_tx_fifo_fifo_reg[5][14]/P0001 , \wishbone_tx_fifo_fifo_reg[5][15]/P0001 , \wishbone_tx_fifo_fifo_reg[5][16]/P0001 , \wishbone_tx_fifo_fifo_reg[5][17]/P0001 , \wishbone_tx_fifo_fifo_reg[5][18]/P0001 , \wishbone_tx_fifo_fifo_reg[5][19]/P0001 , \wishbone_tx_fifo_fifo_reg[5][1]/P0001 , \wishbone_tx_fifo_fifo_reg[5][20]/P0001 , \wishbone_tx_fifo_fifo_reg[5][21]/P0001 , \wishbone_tx_fifo_fifo_reg[5][22]/P0001 , \wishbone_tx_fifo_fifo_reg[5][23]/P0001 , \wishbone_tx_fifo_fifo_reg[5][24]/P0001 , \wishbone_tx_fifo_fifo_reg[5][25]/P0001 , \wishbone_tx_fifo_fifo_reg[5][26]/P0001 , \wishbone_tx_fifo_fifo_reg[5][27]/P0001 , \wishbone_tx_fifo_fifo_reg[5][28]/P0001 , \wishbone_tx_fifo_fifo_reg[5][29]/P0001 , \wishbone_tx_fifo_fifo_reg[5][2]/P0001 , \wishbone_tx_fifo_fifo_reg[5][30]/P0001 , \wishbone_tx_fifo_fifo_reg[5][31]/P0001 , \wishbone_tx_fifo_fifo_reg[5][3]/P0001 , \wishbone_tx_fifo_fifo_reg[5][4]/P0001 , \wishbone_tx_fifo_fifo_reg[5][5]/P0001 , \wishbone_tx_fifo_fifo_reg[5][6]/P0001 , \wishbone_tx_fifo_fifo_reg[5][7]/P0001 , \wishbone_tx_fifo_fifo_reg[5][8]/P0001 , \wishbone_tx_fifo_fifo_reg[5][9]/P0001 , \wishbone_tx_fifo_fifo_reg[6][0]/P0001 , \wishbone_tx_fifo_fifo_reg[6][10]/P0001 , \wishbone_tx_fifo_fifo_reg[6][11]/P0001 , \wishbone_tx_fifo_fifo_reg[6][12]/P0001 , \wishbone_tx_fifo_fifo_reg[6][13]/P0001 , \wishbone_tx_fifo_fifo_reg[6][14]/P0001 , \wishbone_tx_fifo_fifo_reg[6][15]/P0001 , \wishbone_tx_fifo_fifo_reg[6][16]/P0001 , \wishbone_tx_fifo_fifo_reg[6][17]/P0001 , \wishbone_tx_fifo_fifo_reg[6][18]/P0001 , \wishbone_tx_fifo_fifo_reg[6][19]/P0001 , \wishbone_tx_fifo_fifo_reg[6][1]/P0001 , \wishbone_tx_fifo_fifo_reg[6][20]/P0001 , \wishbone_tx_fifo_fifo_reg[6][21]/P0001 , \wishbone_tx_fifo_fifo_reg[6][22]/P0001 , \wishbone_tx_fifo_fifo_reg[6][23]/P0001 , \wishbone_tx_fifo_fifo_reg[6][24]/P0001 , \wishbone_tx_fifo_fifo_reg[6][25]/P0001 , \wishbone_tx_fifo_fifo_reg[6][26]/P0001 , \wishbone_tx_fifo_fifo_reg[6][27]/P0001 , \wishbone_tx_fifo_fifo_reg[6][28]/P0001 , \wishbone_tx_fifo_fifo_reg[6][29]/P0001 , \wishbone_tx_fifo_fifo_reg[6][2]/P0001 , \wishbone_tx_fifo_fifo_reg[6][30]/P0001 , \wishbone_tx_fifo_fifo_reg[6][31]/P0001 , \wishbone_tx_fifo_fifo_reg[6][3]/P0001 , \wishbone_tx_fifo_fifo_reg[6][4]/P0001 , \wishbone_tx_fifo_fifo_reg[6][5]/P0001 , \wishbone_tx_fifo_fifo_reg[6][6]/P0001 , \wishbone_tx_fifo_fifo_reg[6][7]/P0001 , \wishbone_tx_fifo_fifo_reg[6][8]/P0001 , \wishbone_tx_fifo_fifo_reg[6][9]/P0001 , \wishbone_tx_fifo_fifo_reg[7][0]/P0001 , \wishbone_tx_fifo_fifo_reg[7][10]/P0001 , \wishbone_tx_fifo_fifo_reg[7][11]/P0001 , \wishbone_tx_fifo_fifo_reg[7][12]/P0001 , \wishbone_tx_fifo_fifo_reg[7][13]/P0001 , \wishbone_tx_fifo_fifo_reg[7][14]/P0001 , \wishbone_tx_fifo_fifo_reg[7][15]/P0001 , \wishbone_tx_fifo_fifo_reg[7][16]/P0001 , \wishbone_tx_fifo_fifo_reg[7][17]/P0001 , \wishbone_tx_fifo_fifo_reg[7][18]/P0001 , \wishbone_tx_fifo_fifo_reg[7][19]/P0001 , \wishbone_tx_fifo_fifo_reg[7][1]/P0001 , \wishbone_tx_fifo_fifo_reg[7][20]/P0001 , \wishbone_tx_fifo_fifo_reg[7][21]/P0001 , \wishbone_tx_fifo_fifo_reg[7][22]/P0001 , \wishbone_tx_fifo_fifo_reg[7][23]/P0001 , \wishbone_tx_fifo_fifo_reg[7][24]/P0001 , \wishbone_tx_fifo_fifo_reg[7][25]/P0001 , \wishbone_tx_fifo_fifo_reg[7][26]/P0001 , \wishbone_tx_fifo_fifo_reg[7][27]/P0001 , \wishbone_tx_fifo_fifo_reg[7][28]/P0001 , \wishbone_tx_fifo_fifo_reg[7][29]/P0001 , \wishbone_tx_fifo_fifo_reg[7][2]/P0001 , \wishbone_tx_fifo_fifo_reg[7][30]/P0001 , \wishbone_tx_fifo_fifo_reg[7][31]/P0001 , \wishbone_tx_fifo_fifo_reg[7][3]/P0001 , \wishbone_tx_fifo_fifo_reg[7][4]/P0001 , \wishbone_tx_fifo_fifo_reg[7][5]/P0001 , \wishbone_tx_fifo_fifo_reg[7][6]/P0001 , \wishbone_tx_fifo_fifo_reg[7][7]/P0001 , \wishbone_tx_fifo_fifo_reg[7][8]/P0001 , \wishbone_tx_fifo_fifo_reg[7][9]/P0001 , \wishbone_tx_fifo_fifo_reg[8][0]/P0001 , \wishbone_tx_fifo_fifo_reg[8][10]/P0001 , \wishbone_tx_fifo_fifo_reg[8][11]/P0001 , \wishbone_tx_fifo_fifo_reg[8][12]/P0001 , \wishbone_tx_fifo_fifo_reg[8][13]/P0001 , \wishbone_tx_fifo_fifo_reg[8][14]/P0001 , \wishbone_tx_fifo_fifo_reg[8][15]/P0001 , \wishbone_tx_fifo_fifo_reg[8][16]/P0001 , \wishbone_tx_fifo_fifo_reg[8][17]/P0001 , \wishbone_tx_fifo_fifo_reg[8][18]/P0001 , \wishbone_tx_fifo_fifo_reg[8][19]/P0001 , \wishbone_tx_fifo_fifo_reg[8][1]/P0001 , \wishbone_tx_fifo_fifo_reg[8][20]/P0001 , \wishbone_tx_fifo_fifo_reg[8][21]/P0001 , \wishbone_tx_fifo_fifo_reg[8][22]/P0001 , \wishbone_tx_fifo_fifo_reg[8][23]/P0001 , \wishbone_tx_fifo_fifo_reg[8][24]/P0001 , \wishbone_tx_fifo_fifo_reg[8][25]/P0001 , \wishbone_tx_fifo_fifo_reg[8][26]/P0001 , \wishbone_tx_fifo_fifo_reg[8][27]/P0001 , \wishbone_tx_fifo_fifo_reg[8][28]/P0001 , \wishbone_tx_fifo_fifo_reg[8][29]/P0001 , \wishbone_tx_fifo_fifo_reg[8][2]/P0001 , \wishbone_tx_fifo_fifo_reg[8][30]/P0001 , \wishbone_tx_fifo_fifo_reg[8][31]/P0001 , \wishbone_tx_fifo_fifo_reg[8][3]/P0001 , \wishbone_tx_fifo_fifo_reg[8][4]/P0001 , \wishbone_tx_fifo_fifo_reg[8][5]/P0001 , \wishbone_tx_fifo_fifo_reg[8][6]/P0001 , \wishbone_tx_fifo_fifo_reg[8][7]/P0001 , \wishbone_tx_fifo_fifo_reg[8][8]/P0001 , \wishbone_tx_fifo_fifo_reg[8][9]/P0001 , \wishbone_tx_fifo_fifo_reg[9][0]/P0001 , \wishbone_tx_fifo_fifo_reg[9][10]/P0001 , \wishbone_tx_fifo_fifo_reg[9][11]/P0001 , \wishbone_tx_fifo_fifo_reg[9][12]/P0001 , \wishbone_tx_fifo_fifo_reg[9][13]/P0001 , \wishbone_tx_fifo_fifo_reg[9][14]/P0001 , \wishbone_tx_fifo_fifo_reg[9][15]/P0001 , \wishbone_tx_fifo_fifo_reg[9][16]/P0001 , \wishbone_tx_fifo_fifo_reg[9][17]/P0001 , \wishbone_tx_fifo_fifo_reg[9][18]/P0001 , \wishbone_tx_fifo_fifo_reg[9][19]/P0001 , \wishbone_tx_fifo_fifo_reg[9][1]/P0001 , \wishbone_tx_fifo_fifo_reg[9][20]/P0001 , \wishbone_tx_fifo_fifo_reg[9][21]/P0001 , \wishbone_tx_fifo_fifo_reg[9][22]/P0001 , \wishbone_tx_fifo_fifo_reg[9][23]/P0001 , \wishbone_tx_fifo_fifo_reg[9][24]/P0001 , \wishbone_tx_fifo_fifo_reg[9][25]/P0001 , \wishbone_tx_fifo_fifo_reg[9][26]/P0001 , \wishbone_tx_fifo_fifo_reg[9][27]/P0001 , \wishbone_tx_fifo_fifo_reg[9][28]/P0001 , \wishbone_tx_fifo_fifo_reg[9][29]/P0001 , \wishbone_tx_fifo_fifo_reg[9][2]/P0001 , \wishbone_tx_fifo_fifo_reg[9][30]/P0001 , \wishbone_tx_fifo_fifo_reg[9][31]/P0001 , \wishbone_tx_fifo_fifo_reg[9][3]/P0001 , \wishbone_tx_fifo_fifo_reg[9][4]/P0001 , \wishbone_tx_fifo_fifo_reg[9][5]/P0001 , \wishbone_tx_fifo_fifo_reg[9][6]/P0001 , \wishbone_tx_fifo_fifo_reg[9][7]/P0001 , \wishbone_tx_fifo_fifo_reg[9][8]/P0001 , \wishbone_tx_fifo_fifo_reg[9][9]/P0001 , \wishbone_tx_fifo_read_pointer_reg[0]/NET0131 , \wishbone_tx_fifo_read_pointer_reg[1]/NET0131 , \wishbone_tx_fifo_read_pointer_reg[2]/NET0131 , \wishbone_tx_fifo_read_pointer_reg[3]/NET0131 , \wishbone_tx_fifo_write_pointer_reg[0]/NET0131 , \wishbone_tx_fifo_write_pointer_reg[1]/NET0131 , \wishbone_tx_fifo_write_pointer_reg[2]/NET0131 , \wishbone_tx_fifo_write_pointer_reg[3]/NET0131 , \_al_n1 , \g215539/_0_ , \g215543/_0_ , \g215547/_0_ , \g215551/_0_ , \g215552/_0_ , \g215578/_0_ , \g215587/_1_ , \g215589/_1_ , \g215591/_1_ , \g215593/_1_ , \g215595/_1_ , \g215597/_1_ , \g215599/_1_ , \g215601/_1_ , \g215603/_1_ , \g215605/_1_ , \g215607/_1_ , \g215609/_1_ , \g215611/_1_ , \g215613/_1_ , \g215615/_1_ , \g215617/_1_ , \g215618/_0_ , \g215619/_0_ , \g215620/_0_ , \g215632/_1_ , \g215634/_0_ , \g215635/_0_ , \g215636/_0_ , \g215637/_0_ , \g215638/_0_ , \g215639/_0_ , \g215655/_1_ , \g215657/_1_ , \g215659/_1_ , \g215661/_1_ , \g215662/_0_ , \g215663/_0_ , \g215664/_0_ , \g215665/_0_ , \g215668/_0_ , \g215674/_0_ , \g215677/_0_ , \g215686/_0_ , \g215695/_0_ , \g215696/_0_ , \g215702/_1__syn_2 , \g215705/_0_ , \g215706/_0_ , \g215716/_0_ , \g215717/_0_ , \g215718/_0_ , \g215726/_0_ , \g215727/_0_ , \g215728/_0_ , \g215760/_0_ , \g215764/_0_ , \g215765/_0_ , \g215766/_0_ , \g215767/_3_ , \g215768/_3_ , \g215769/_3_ , \g215770/_3_ , \g215771/_3_ , \g215772/_3_ , \g215773/_3_ , \g215774/_3_ , \g215775/_3_ , \g215776/_3_ , \g215777/_3_ , \g215778/_3_ , \g215779/_3_ , \g215780/_3_ , \g215790/_0_ , \g215791/_0_ , \g215792/_0_ , \g215793/_0_ , \g215801/_0_ , \g215802/_0_ , \g215803/_0_ , \g215804/_0_ , \g215812/_0_ , \g215813/_0_ , \g215821/_0_ , \g215823/_0_ , \g215831/_0_ , \g215832/_0_ , \g215833/_0_ , \g215845/_0_ , \g215846/_0_ , \g215847/_0_ , \g215872/_0_ , \g215873/_0_ , \g215874/_0_ , \g215904/_0_ , \g215905/_0_ , \g215906/_0_ , \g215907/_0_ , \g215908/_0_ , \g215909/_0_ , \g215910/_0_ , \g215911/_0_ , \g215912/_0_ , \g215913/_0_ , \g215914/_0_ , \g215915/_0_ , \g215916/_0_ , \g215917/_0_ , \g215918/_0_ , \g215919/_0_ , \g215920/_0_ , \g215923/_0_ , \g215926/_0_ , \g215941/_0_ , \g215942/_0_ , \g215943/_0_ , \g215944/_0_ , \g215945/_0_ , \g215946/_0_ , \g215947/_0_ , \g215948/_0_ , \g215949/_0_ , \g215950/_0_ , \g215951/_0_ , \g215952/_0_ , \g215953/_0_ , \g215954/_0_ , \g215955/_0_ , \g215956/_0_ , \g215957/_0_ , \g215959/_00_ , \g215960/_0_ , \g215962/_0_ , \g215964/_0_ , \g215966/_0_ , \g215972/_0_ , \g216035/_0_ , \g216037/_0_ , \g216038/_0_ , \g216039/_0_ , \g216040/_0_ , \g216041/_0_ , \g216042/_0_ , \g216046/_0_ , \g216048/_0_ , \g216057/_0_ , \g216263/_0_ , \g216264/_0_ , \g216265/_0_ , \g216266/_0_ , \g216267/_0_ , \g216268/_0_ , \g216269/_0_ , \g216270/_0_ , \g216271/_0_ , \g216272/_0_ , \g216273/_0_ , \g216284/_0_ , \g216289/_0_ , \g216290/_0_ , \g216292/_0_ , \g216296/_0_ , \g216297/_0_ , \g216300/_0_ , \g216301/_0_ , \g216302/_0_ , \g216303/_0_ , \g216304/_0_ , \g216305/_0_ , \g216306/_0_ , \g216307/_0_ , \g216310/_3_ , \g216311/_3_ , \g216314/u3_syn_7 , \g216322/_3_ , \g216323/_3_ , \g216324/_3_ , \g216325/_3_ , \g216326/_3_ , \g216327/_3_ , \g216328/_3_ , \g216329/_3_ , \g216369/_0_ , \g216370/_0_ , \g216371/_0_ , \g216372/_0_ , \g216373/_0_ , \g216374/_0_ , \g216375/_0_ , \g216376/_0_ , \g216379/_0_ , \g216380/_0_ , \g216381/_0_ , \g216385/_0_ , \g216389/_0_ , \g216390/_0_ , \g216402/_0_ , \g216404/_0_ , \g216405/_0_ , \g216406/_0_ , \g216407/_0_ , \g216408/_0_ , \g216409/_0_ , \g216410/_0_ , \g216411/_0_ , \g216412/_0_ , \g216413/_0_ , \g216414/_0_ , \g216415/_0_ , \g216416/_0_ , \g216417/_0_ , \g216418/_0_ , \g216419/_0_ , \g216420/_0_ , \g216421/_0_ , \g216422/_0_ , \g216423/_0_ , \g216424/_0_ , \g216425/_0_ , \g216426/_0_ , \g216427/_0_ , \g216428/_0_ , \g216429/_0_ , \g216430/_0_ , \g216431/_0_ , \g216432/_0_ , \g216433/_0_ , \g216434/_0_ , \g216435/_0_ , \g216436/_0_ , \g216437/_0_ , \g216438/_0_ , \g216439/_3_ , \g216447/_3_ , \g216448/_3_ , \g216452/_0_ , \g216453/_0_ , \g216454/_0_ , \g216455/_0_ , \g216456/_0_ , \g216457/_0_ , \g216458/_3_ , \g216459/_3_ , \g216461/_3_ , \g216462/_3_ , \g216463/_3_ , \g216464/_3_ , \g216465/_3_ , \g216466/_0_ , \g216467/_3_ , \g216468/_3_ , \g216469/_3_ , \g216470/_3_ , \g216471/_3_ , \g216473/_3_ , \g216474/_3_ , \g216475/_3_ , \g216476/_3_ , \g216477/_3_ , \g216478/_0_ , \g216479/_3_ , \g216480/_3_ , \g216481/_3_ , \g216492/_0_ , \g216494/_0_ , \g216495/_3_ , \g216496/_3_ , \g216498/_3_ , \g216499/_3_ , \g216500/_3_ , \g216513/_3_ , \g216514/_3_ , \g216515/_3_ , \g216516/_3_ , \g216517/_3_ , \g216518/_3_ , \g216519/_3_ , \g216520/_3_ , \g216521/_3_ , \g216522/_3_ , \g216523/_3_ , \g216524/_3_ , \g216525/_3_ , \g216526/_3_ , \g216527/_3_ , \g216528/_3_ , \g216529/_3_ , \g216530/_3_ , \g216531/_3_ , \g216532/_3_ , \g216533/_3_ , \g216534/_3_ , \g216535/_3_ , \g216536/_3_ , \g216537/_3_ , \g216538/_3_ , \g216555/_3_ , \g216556/_3_ , \g216557/_3_ , \g216560/_3_ , \g216561/_3_ , \g216562/_3_ , \g216563/_3_ , \g216564/_3_ , \g216565/_3_ , \g216566/_3_ , \g216567/_3_ , \g216568/_3_ , \g216569/_3_ , \g216570/_3_ , \g216571/_3_ , \g216575/_3_ , \g216576/_3_ , \g216577/_3_ , \g216578/_3_ , \g216579/_3_ , \g216580/_3_ , \g216581/_3_ , \g216582/_3_ , \g216583/_3_ , \g216586/_3_ , \g216587/_3_ , \g216588/_3_ , \g216589/_3_ , \g216590/_3_ , \g216591/_3_ , \g216592/_3_ , \g216593/_3_ , \g216594/_3_ , \g216595/_3_ , \g216600/_3_ , \g216683/_0_ , \g216689/_0_ , \g216693/_0_ , \g216694/_0_ , \g216727/_0_ , \g216728/_0_ , \g216729/_0_ , \g216732/_0_ , \g216733/_0_ , \g216734/_0_ , \g216735/_0_ , \g216736/_0_ , \g216737/_0_ , \g216738/_0_ , \g216739/_0_ , \g216740/_0_ , \g216741/_0_ , \g216742/_0_ , \g216743/_0_ , \g216744/_0_ , \g216745/_0_ , \g216746/_0_ , \g216748/_0_ , \g216751/_0_ , \g216754/_0_ , \g216762/_0_ , \g216934/_2_ , \g216952/_0_ , \g216955/_0_ , \g216969/_0_ , \g216979/_0_ , \g216984/_0_ , \g216996/_0_ , \g217002/_0_ , \g217014/_0_ , \g217015/_0_ , \g217016/_0_ , \g217017/_0_ , \g217018/_0_ , \g217019/_0_ , \g217023/_0_ , \g217116/_0_ , \g217146/_3_ , \g217149/_0_ , \g217151/_0_ , \g217160/_0_ , \g217167/_0_ , \g217168/_0_ , \g217169/_0_ , \g217170/_0_ , \g217171/_0_ , \g217172/_0_ , \g217173/_0_ , \g217174/_0_ , \g217175/_0_ , \g217176/_0_ , \g217177/_0_ , \g217178/_0_ , \g217179/_0_ , \g217180/_0_ , \g217181/_0_ , \g217182/_0_ , \g217183/_0_ , \g217187/_0_ , \g217188/_0_ , \g217189/_0_ , \g217193/_0_ , \g217194/_0_ , \g217195/_0_ , \g217196/_0_ , \g217202/_0_ , \g217205/_0_ , \g217206/_0_ , \g217207/_0_ , \g217208/_0_ , \g217209/_0_ , \g217210/_0_ , \g217211/_0_ , \g217212/_0_ , \g217213/_0_ , \g217214/_0_ , \g217215/_0_ , \g217216/_0_ , \g217217/_0_ , \g217218/_0_ , \g217219/_0_ , \g217220/_0_ , \g217223/_0_ , \g217231/_0_ , \g217237/_0_ , \g217238/_0_ , \g217242/_0_ , \g217243/_0_ , \g217250/_3_ , \g217251/_3_ , \g217252/_3_ , \g217253/_3_ , \g217254/_3_ , \g217255/_3_ , \g217256/_3_ , \g217257/_3_ , \g217258/_3_ , \g217259/_3_ , \g217260/_3_ , \g217261/_3_ , \g217262/_3_ , \g217263/_3_ , \g217264/_3_ , \g217265/_3_ , \g217266/_3_ , \g217267/_3_ , \g217268/_3_ , \g217269/_3_ , \g217270/_3_ , \g217271/_3_ , \g217272/_3_ , \g217273/_3_ , \g217274/_3_ , \g217275/_3_ , \g217276/_3_ , \g217277/_3_ , \g217278/_3_ , \g217279/_3_ , \g217280/_3_ , \g217281/_3_ , \g217282/_3_ , \g217283/_3_ , \g217284/_3_ , \g217285/_3_ , \g217286/_3_ , \g217287/_3_ , \g217288/_3_ , \g217289/_3_ , \g217290/_3_ , \g217291/_3_ , \g217292/_3_ , \g217293/_3_ , \g217294/_3_ , \g217295/_3_ , \g217296/_3_ , \g217297/_3_ , \g217298/_3_ , \g217299/_3_ , \g217300/_3_ , \g217301/_3_ , \g217302/_3_ , \g217303/_3_ , \g217304/_3_ , \g217305/_3_ , \g217306/_3_ , \g217307/_3_ , \g217308/_3_ , \g217309/_3_ , \g217310/_3_ , \g217311/_3_ , \g217312/_3_ , \g217313/_3_ , \g217318/_0_ , \g217662/_0_ , \g217663/_0_ , \g217682/_0_ , \g217697/_0_ , \g217698/_0_ , \g217699/_0_ , \g217700/_0_ , \g217701/_0_ , \g217705/_0_ , \g217711/_0_ , \g217747/_0_ , \g217753/_00_ , \g217775/_0_ , \g217781/_0_ , \g217784/_0_ , \g217785/_0_ , \g217786/_0_ , \g217787/_0_ , \g217788/_0_ , \g217790/_0_ , \g217815/_0_ , \g217817/_0_ , \g218145/_0_ , \g218148/_0_ , \g218150/_0_ , \g218167/_0_ , \g218168/_0_ , \g218234/_0_ , \g218235/_0_ , \g218236/_0_ , \g218238/_0_ , \g218242/_0_ , \g218332/_0_ , \g218335/_0_ , \g218336/_0_ , \g218337/_0_ , \g218338/_0_ , \g218339/_0_ , \g218340/_0_ , \g218341/_0_ , \g218342/_0_ , \g218343/_0_ , \g218344/_0_ , \g218345/_0_ , \g218346/_0_ , \g218347/_0_ , \g218348/_0_ , \g218349/_0_ , \g218350/_0_ , \g218351/_0_ , \g218352/_0_ , \g218353/_0_ , \g218354/_0_ , \g218355/_0_ , \g218356/_0_ , \g218357/_0_ , \g218358/_0_ , \g218359/_0_ , \g218360/_0_ , \g218398/_3_ , \g218430/_0_ , \g218440/_0_ , \g218452/u3_syn_4 , \g218495/u3_syn_4 , \g218517/u3_syn_4 , \g218554/u3_syn_4 , \g218575/u3_syn_4 , \g218600/u3_syn_4 , \g218621/u3_syn_4 , \g218638/u3_syn_4 , \g218659/u3_syn_4 , \g218673/u3_syn_4 , \g218707/u3_syn_4 , \g218735/_3_ , \g219186/_0_ , \g219187/_0_ , \g219188/_0_ , \g219189/_0_ , \g219190/_0_ , \g219196/_0_ , \g219198/_0_ , \g219199/_0_ , \g219200/_0_ , \g219308/_0_ , \g219314/_0_ , \g219326/_0_ , \g219328/_0_ , \g219348/_0_ , \g219351/_0_ , \g219363/_0_ , \g219364/_0_ , \g219365/_0_ , \g219366/_0_ , \g219367/_0_ , \g219368/_0_ , \g219369/_0_ , \g219376/_0_ , \g219381/_0_ , \g219382/_0_ , \g219384/_0_ , \g219385/_0_ , \g219391/_0_ , \g219394/_0_ , \g219395/_0_ , \g219396/_0_ , \g219397/_0_ , \g219398/_0_ , \g219399/_0_ , \g219400/_0_ , \g219401/_0_ , \g219402/_0_ , \g219403/_0_ , \g219404/_0_ , \g219405/_0_ , \g219406/_0_ , \g219407/_0_ , \g219408/_0_ , \g219409/_0_ , \g219410/_0_ , \g219411/_0_ , \g219412/_0_ , \g219413/_0_ , \g219414/_0_ , \g219415/_0_ , \g219416/_0_ , \g219417/_0_ , \g219418/_0_ , \g219419/_0_ , \g219420/_0_ , \g219421/_0_ , \g219422/_0_ , \g219423/_0_ , \g219424/_0_ , \g219425/_0_ , \g219426/_0_ , \g219427/_0_ , \g219428/_0_ , \g219429/_0_ , \g219430/_0_ , \g219431/_0_ , \g219432/_0_ , \g219433/_0_ , \g219434/_0_ , \g219435/_0_ , \g219436/_0_ , \g219437/_0_ , \g219438/_0_ , \g219439/_0_ , \g219440/_0_ , \g219441/_0_ , \g219442/_0_ , \g219443/_0_ , \g219444/_0_ , \g219445/_0_ , \g219446/_0_ , \g219447/_0_ , \g219449/_0_ , \g219450/_0_ , \g219451/_0_ , \g219452/_0_ , \g219453/_0_ , \g219454/_0_ , \g219455/_0_ , \g219456/_0_ , \g219457/_0_ , \g219458/_0_ , \g219464/u3_syn_7 , \g219496/u3_syn_4 , \g219512/u3_syn_4 , \g219526/u3_syn_4 , \g219549/u3_syn_4 , \g219571/u3_syn_4 , \g219588/u3_syn_4 , \g219603/u3_syn_4 , \g219621/u3_syn_4 , \g219636/_3_ , \g219652/u3_syn_4 , \g219676/_3_ , \g219686/_0_ , \g219689/_0_ , \g219694/_3_ , \g220062/_0_ , \g220068/_0_ , \g220069/_0_ , \g220072/_0_ , \g220084/_0_ , \g220149/_0_ , \g220162/_0_ , \g220317/_0_ , \g220360/_2_ , \g220368/_2_ , \g220369/_0_ , \g220370/_0_ , \g220371/_0_ , \g220372/_0_ , \g220376/_0_ , \g220390/_0_ , \g220395/_0_ , \g220499/_0_ , \g220500/_0_ , \g220501/_0_ , \g220502/_0_ , \g220503/_0_ , \g220504/_0_ , \g220505/_0_ , \g220506/_0_ , \g220507/_0_ , \g220508/_0_ , \g220509/_0_ , \g220510/_0_ , \g220511/_0_ , \g220512/_0_ , \g220513/_0_ , \g220514/_0_ , \g220515/_0_ , \g220516/_0_ , \g220517/_0_ , \g220518/_0_ , \g220519/_0_ , \g220520/_0_ , \g220521/_0_ , \g220522/_0_ , \g220523/_0_ , \g220524/_0_ , \g220525/_0_ , \g220526/_0_ , \g220527/_0_ , \g220528/_0_ , \g220529/_0_ , \g220530/_0_ , \g220531/_0_ , \g220532/_0_ , \g220533/_0_ , \g220534/_0_ , \g220535/_0_ , \g220557/_0_ , \g220558/_0_ , \g220559/_0_ , \g220560/_0_ , \g220561/_0_ , \g220562/_0_ , \g220563/_0_ , \g220564/_0_ , \g220565/_0_ , \g220566/_0_ , \g220567/_0_ , \g220568/_0_ , \g220569/_0_ , \g220570/_0_ , \g220571/_0_ , \g220572/_0_ , \g220573/_0_ , \g220574/_0_ , \g220575/_0_ , \g220576/_0_ , \g220577/_0_ , \g220578/_0_ , \g220579/_0_ , \g220580/_0_ , \g220581/_0_ , \g220582/_0_ , \g220583/_0_ , \g220584/_0_ , \g220585/_0_ , \g220586/_0_ , \g220587/_0_ , \g220588/_0_ , \g220589/_0_ , \g220590/_0_ , \g220591/_0_ , \g220592/_0_ , \g220593/_0_ , \g220594/_0_ , \g220595/_0_ , \g220596/_0_ , \g220597/_0_ , \g220598/_0_ , \g220599/_0_ , \g220600/_0_ , \g220601/_0_ , \g220602/_0_ , \g220603/_0_ , \g220604/_0_ , \g220605/_0_ , \g220606/_0_ , \g220607/_0_ , \g220608/_0_ , \g220609/_0_ , \g220610/_0_ , \g220611/_0_ , \g220612/_0_ , \g220613/_0_ , \g220614/_0_ , \g220615/_0_ , \g220616/_0_ , \g220617/_0_ , \g220618/_0_ , \g220619/_0_ , \g220620/_0_ , \g220621/_0_ , \g220622/_0_ , \g220623/_0_ , \g220624/_0_ , \g220625/_0_ , \g220626/_0_ , \g220627/_0_ , \g220628/_0_ , \g220629/_0_ , \g220630/_0_ , \g220631/_0_ , \g220632/_0_ , \g220633/_0_ , \g220634/_0_ , \g220635/_0_ , \g220636/_0_ , \g220637/_0_ , \g220638/_0_ , \g220639/_0_ , \g220640/_0_ , \g220641/_0_ , \g220642/_0_ , \g220643/_0_ , \g220644/_0_ , \g220645/_0_ , \g220646/_0_ , \g220647/_0_ , \g220648/_0_ , \g220649/_0_ , \g220650/_0_ , \g220651/_0_ , \g220652/_0_ , \g220653/_0_ , \g220654/_0_ , \g220655/_0_ , \g220656/_0_ , \g220657/_0_ , \g220658/_0_ , \g220659/_0_ , \g220660/_0_ , \g220661/_0_ , \g220662/_0_ , \g220663/_0_ , \g220664/_0_ , \g220665/_0_ , \g220666/_0_ , \g220674/_0_ , \g220679/u3_syn_7 , \g220711/u3_syn_4 , \g220726/u3_syn_4 , \g220739/u3_syn_4 , \g220751/u3_syn_4 , \g220759/u3_syn_4 , \g220773/u3_syn_4 , \g220782/u3_syn_4 , \g220805/u3_syn_4 , \g220828/u3_syn_4 , \g220921/_0_ , \g220930/u3_syn_4 , \g220949/_3_ , \g220994/_3_ , \g221207/_0_ , \g221213/_0_ , \g221223/_0_ , \g221224/_0_ , \g221225/_0_ , \g221226/_0_ , \g221231/_0_ , \g221232/_0_ , \g221234/_0_ , \g221235/_0_ , \g221246/_2_ , \g221249/_2_ , \g221265/_0_ , \g221287/_0_ , \g221325/_0_ , \g221326/_0_ , \g221447/_0_ , \g221449/_0_ , \g221452/_0_ , \g221469/_0_ , \g221473/_0_ , \g221503/_0_ , \g221510/_0_ , \g221512/_0_ , \g221516/_0_ , \g221517/_0_ , \g221524/_0_ , \g221530/_0_ , \g221592/_0_ , \g221593/_0_ , \g221634/u3_syn_4 , \g221669/u3_syn_4 , \g221789/u3_syn_4 , \g221813/u3_syn_4 , \g221829/u3_syn_4 , \g221861/u3_syn_4 , \g221876/_0_ , \g221935/_0_ , \g221944/_3_ , \g230200/_0_ , \g230201/_0_ , \g230205/_0_ , \g230295/_0_ , \g230297/_0_ , \g230298/_0_ , \g230300/_0_ , \g230302/_0_ , \g230303/_0_ , \g230343/_0_ , \g230368/_0_ , \g230511/_0_ , \g230531/_0_ , \g230635/_2_ , \g230661/_0_ , \g230715/_1__syn_2 , \g230731/_0_ , \g230766/_0_ , \g230784/_0_ , \g230785/_0_ , \g230786/_0_ , \g230787/_0_ , \g230797/_0_ , \g230798/_0_ , \g230803/_0_ , \g230804/_00_ , \g230805/_00_ , \g230806/_00_ , \g230807/_00_ , \g230808/_00_ , \g230809/_00_ , \g230815/_0_ , \g230816/_2_ , \g230817/_2_ , \g230829/_0_ , \g230834/_0_ , \g230835/_0_ , \g230836/_0_ , \g230837/_0_ , \g230844/_0_ , \g230863/_3_ , \g230864/_3_ , \g230870/_0_ , \g230988/_3_ , \g231010/_3_ , \g231016/_3_ , \g231042/_3_ , \g231471/_0_ , \g231472/_0_ , \g231476/_3_ , \g231480/_3_ , \g231484/_3_ , \g231504/_0_ , \g231532/_0_ , \g231542/_0_ , \g231560/_1_ , \g231578/_1_ , \g231580/_0_ , \g231590/_1__syn_2 , \g231615/_0_ , \g231623/_1_ , \g231634/_2_ , \g231635/_0_ , \g231638/_2_ , \g231640/_0_ , \g231653/_2_ , \g231787/_0_ , \g231931/_0_ , \g231939/_3_ , \g231940/_0_ , \g231951/_0_ , \g231955/_0_ , \g231956/_0_ , \g231959/_2_ , \g231960/_0_ , \g231964/_0_ , \g231965/_0_ , \g231975/_0_ , \g231986/_1_ , \g231987/_1_ , \g231989/_1_ , \g231990/_1_ , \g231991/_0_ , \g231992/_0_ , \g231995/_0_ , \g231998/_0_ , \g231999/_0_ , \g232002/_3_ , \g232035/u3_syn_4 , \g232038/u3_syn_4 , \g232046/u3_syn_4 , \g232054/u3_syn_4 , \g232062/u3_syn_4 , \g232070/u3_syn_4 , \g232078/u3_syn_4 , \g232079/u3_syn_4 , \g232087/u3_syn_4 , \g232096/u3_syn_4 , \g232104/u3_syn_4 , \g232112/u3_syn_4 , \g232120/u3_syn_4 , \g232128/u3_syn_4 , \g232136/u3_syn_4 , \g232144/u3_syn_4 , \g232152/u3_syn_4 , \g232161/u3_syn_4 , \g232169/u3_syn_4 , \g232177/u3_syn_4 , \g232185/u3_syn_4 , \g232186/u3_syn_4 , \g232194/u3_syn_4 , \g232202/u3_syn_4 , \g232210/u3_syn_4 , \g232218/u3_syn_4 , \g232226/u3_syn_4 , \g232234/u3_syn_4 , \g232242/u3_syn_4 , \g232251/u3_syn_4 , \g232259/u3_syn_4 , \g232267/u3_syn_4 , \g232275/u3_syn_4 , \g232283/u3_syn_4 , \g232291/u3_syn_4 , \g232299/u3_syn_4 , \g232307/u3_syn_4 , \g232315/u3_syn_4 , \g232324/u3_syn_4 , \g232332/u3_syn_4 , \g232341/u3_syn_4 , \g232349/u3_syn_4 , \g232357/u3_syn_4 , \g232366/u3_syn_4 , \g232374/u3_syn_4 , \g232382/u3_syn_4 , \g232390/u3_syn_4 , \g232398/u3_syn_4 , \g232406/u3_syn_4 , \g232414/u3_syn_4 , \g232422/u3_syn_4 , \g232427/u3_syn_4 , \g232431/u3_syn_4 , \g232439/u3_syn_4 , \g232444/u3_syn_4 , \g232452/u3_syn_4 , \g232461/u3_syn_4 , \g232471/u3_syn_4 , \g232479/u3_syn_4 , \g232487/u3_syn_4 , \g232495/u3_syn_4 , \g232503/u3_syn_4 , \g232506/u3_syn_4 , \g232514/u3_syn_4 , \g232527/u3_syn_4 , \g232530/u3_syn_4 , \g232536/u3_syn_4 , \g232544/u3_syn_4 , \g232551/u3_syn_4 , \g232557/u3_syn_4 , \g232568/u3_syn_4 , \g232576/u3_syn_4 , \g232585/u3_syn_4 , \g232593/u3_syn_4 , \g232597/u3_syn_4 , \g232609/u3_syn_4 , \g232617/u3_syn_4 , \g232625/u3_syn_4 , \g232633/u3_syn_4 , \g232641/u3_syn_4 , \g232649/u3_syn_4 , \g232657/u3_syn_4 , \g232665/u3_syn_4 , \g232673/u3_syn_4 , \g232681/u3_syn_4 , \g232689/u3_syn_4 , \g232697/u3_syn_4 , \g232705/u3_syn_4 , \g232713/u3_syn_4 , \g232717/u3_syn_4 , \g232729/u3_syn_4 , \g232737/u3_syn_4 , \g232745/u3_syn_4 , \g232749/u3_syn_4 , \g232761/u3_syn_4 , \g232768/u3_syn_4 , \g232777/u3_syn_4 , \g232785/u3_syn_4 , \g232793/u3_syn_4 , \g232801/u3_syn_4 , \g232809/u3_syn_4 , \g232815/u3_syn_4 , \g232823/u3_syn_4 , \g232833/u3_syn_4 , \g232841/u3_syn_4 , \g232846/u3_syn_4 , \g232851/u3_syn_4 , \g232865/u3_syn_4 , \g232873/u3_syn_4 , \g232881/u3_syn_4 , \g232882/u3_syn_4 , \g232895/u3_syn_4 , \g232904/u3_syn_4 , \g232913/u3_syn_4 , \g232921/u3_syn_4 , \g232928/u3_syn_4 , \g232934/u3_syn_4 , \g232945/u3_syn_4 , \g232953/u3_syn_4 , \g232954/u3_syn_4 , \g232969/u3_syn_4 , \g232977/u3_syn_4 , \g232981/u3_syn_4 , \g232993/u3_syn_4 , \g232995/u3_syn_4 , \g233009/u3_syn_4 , \g233017/u3_syn_4 , \g233025/u3_syn_4 , \g233033/u3_syn_4 , \g233041/u3_syn_4 , \g233047/u3_syn_4 , \g233057/u3_syn_4 , \g233065/u3_syn_4 , \g233073/u3_syn_4 , \g233081/u3_syn_4 , \g233087/u3_syn_4 , \g233097/u3_syn_4 , \g233105/u3_syn_4 , \g233113/u3_syn_4 , \g233121/u3_syn_4 , \g233128/u3_syn_4 , \g233134/u3_syn_4 , \g233144/u3_syn_4 , \g233153/u3_syn_4 , \g233161/u3_syn_4 , \g233169/u3_syn_4 , \g233177/u3_syn_4 , \g233185/u3_syn_4 , \g233193/u3_syn_4 , \g233201/u3_syn_4 , \g233209/u3_syn_4 , \g233217/u3_syn_4 , \g233219/u3_syn_4 , \g233229/u3_syn_4 , \g233241/u3_syn_4 , \g233249/u3_syn_4 , \g233257/u3_syn_4 , \g233265/u3_syn_4 , \g233273/u3_syn_4 , \g233281/u3_syn_4 , \g233289/u3_syn_4 , \g233297/u3_syn_4 , \g233305/u3_syn_4 , \g233313/u3_syn_4 , \g233321/u3_syn_4 , \g233329/u3_syn_4 , \g233337/u3_syn_4 , \g233345/u3_syn_4 , \g233353/u3_syn_4 , \g233361/u3_syn_4 , \g233369/u3_syn_4 , \g233377/u3_syn_4 , \g233382/u3_syn_4 , \g233392/u3_syn_4 , \g233394/u3_syn_4 , \g233409/u3_syn_4 , \g233417/u3_syn_4 , \g233425/u3_syn_4 , \g233433/u3_syn_4 , \g233441/u3_syn_4 , \g233449/u3_syn_4 , \g233453/u3_syn_4 , \g233465/u3_syn_4 , \g233473/u3_syn_4 , \g233481/u3_syn_4 , \g233489/u3_syn_4 , \g233497/u3_syn_4 , \g233505/u3_syn_4 , \g233513/u3_syn_4 , \g233516/u3_syn_4 , \g233529/u3_syn_4 , \g233531/u3_syn_4 , \g233546/u3_syn_4 , \g233554/u3_syn_4 , \g233562/u3_syn_4 , \g233570/u3_syn_4 , \g233578/u3_syn_4 , \g233586/u3_syn_4 , \g233594/u3_syn_4 , \g233602/u3_syn_4 , \g233603/u3_syn_4 , \g233618/u3_syn_4 , \g233626/u3_syn_4 , \g233634/u3_syn_4 , \g233642/u3_syn_4 , \g233650/u3_syn_4 , \g233658/u3_syn_4 , \g233666/u3_syn_4 , \g233674/u3_syn_4 , \g233682/u3_syn_4 , \g233690/u3_syn_4 , \g233698/u3_syn_4 , \g233706/u3_syn_4 , \g233714/u3_syn_4 , \g233722/u3_syn_4 , \g233730/u3_syn_4 , \g233738/u3_syn_4 , \g233746/u3_syn_4 , \g233754/u3_syn_4 , \g233762/u3_syn_4 , \g233770/u3_syn_4 , \g233778/u3_syn_4 , \g233783/u3_syn_4 , \g233794/u3_syn_4 , \g233802/u3_syn_4 , \g233806/u3_syn_4 , \g233818/u3_syn_4 , \g233826/u3_syn_4 , \g233828/u3_syn_4 , \g233838/u3_syn_4 , \g233850/u3_syn_4 , \g233858/u3_syn_4 , \g233860/u3_syn_4 , \g233870/u3_syn_4 , \g233881/u3_syn_4 , \g233890/u3_syn_4 , \g233899/u3_syn_4 , \g233908/u3_syn_4 , \g233917/u3_syn_4 , \g233919/u3_syn_4 , \g233927/u3_syn_4 , \g233935/u3_syn_4 , \g233943/u3_syn_4 , \g233945/u3_syn_4 , \g233953/u3_syn_4 , \g233961/u3_syn_4 , \g233969/u3_syn_4 , \g233977/u3_syn_4 , \g233985/u3_syn_4 , \g233993/u3_syn_4 , \g234001/u3_syn_4 , \g234008/u3_syn_4 , \g234009/u3_syn_4 , \g234024/u3_syn_4 , \g234032/u3_syn_4 , \g234038/u3_syn_4 , \g234056/u3_syn_4 , \g234063/u3_syn_4 , \g234071/u3_syn_4 , \g234079/u3_syn_4 , \g234098/u3_syn_4 , \g234106/u3_syn_4 , \g234114/u3_syn_4 , \g234122/u3_syn_4 , \g234130/u3_syn_4 , \g234138/u3_syn_4 , \g234145/u3_syn_4 , \g234156/u3_syn_4 , \g234162/u3_syn_4 , \g234171/u3_syn_4 , \g234183/u3_syn_4 , \g234248/u3_syn_4 , \g234265/u3_syn_4 , \g234273/u3_syn_4 , \g234281/u3_syn_4 , \g234289/u3_syn_4 , \g234297/u3_syn_4 , \g234306/u3_syn_4 , \g234314/u3_syn_4 , \g234322/u3_syn_4 , \g234331/u3_syn_4 , \g234339/u3_syn_4 , \g234347/u3_syn_4 , \g234355/u3_syn_4 , \g234363/u3_syn_4 , \g234371/u3_syn_4 , \g234379/u3_syn_4 , \g234387/u3_syn_4 , \g234395/u3_syn_4 , \g234403/u3_syn_4 , \g234411/u3_syn_4 , \g234419/u3_syn_4 , \g234427/u3_syn_4 , \g234435/u3_syn_4 , \g234443/u3_syn_4 , \g234451/u3_syn_4 , \g234459/u3_syn_4 , \g234467/u3_syn_4 , \g234475/u3_syn_4 , \g234483/u3_syn_4 , \g234491/u3_syn_4 , \g234499/u3_syn_4 , \g234507/u3_syn_4 , \g234515/u3_syn_4 , \g234523/u3_syn_4 , \g234531/u3_syn_4 , \g234539/u3_syn_4 , \g234547/u3_syn_4 , \g234555/u3_syn_4 , \g234563/u3_syn_4 , \g234571/u3_syn_4 , \g234579/u3_syn_4 , \g234587/u3_syn_4 , \g234595/u3_syn_4 , \g234604/u3_syn_4 , \g234612/u3_syn_4 , \g234620/u3_syn_4 , \g234628/u3_syn_4 , \g234636/u3_syn_4 , \g234644/u3_syn_4 , \g234652/u3_syn_4 , \g234660/u3_syn_4 , \g234668/u3_syn_4 , \g234676/u3_syn_4 , \g234684/u3_syn_4 , \g234692/u3_syn_4 , \g234700/u3_syn_4 , \g234708/u3_syn_4 , \g234716/u3_syn_4 , \g234725/u3_syn_4 , \g234733/u3_syn_4 , \g234741/u3_syn_4 , \g234749/u3_syn_4 , \g234757/u3_syn_4 , \g234765/u3_syn_4 , \g234773/u3_syn_4 , \g234781/u3_syn_4 , \g234789/u3_syn_4 , \g234798/u3_syn_4 , \g234806/u3_syn_4 , \g234814/u3_syn_4 , \g234822/u3_syn_4 , \g234830/u3_syn_4 , \g234838/u3_syn_4 , \g235911/u3_syn_4 , \g235912/u3_syn_4 , \g235920/u3_syn_4 , \g235928/u3_syn_4 , \g235936/u3_syn_4 , \g235944/u3_syn_4 , \g235952/u3_syn_4 , \g235960/u3_syn_4 , \g235968/u3_syn_4 , \g235976/u3_syn_4 , \g235984/u3_syn_4 , \g235992/u3_syn_4 , \g236000/u3_syn_4 , \g236008/u3_syn_4 , \g236016/u3_syn_4 , \g236021/u3_syn_4 , \g236025/u3_syn_4 , \g236033/u3_syn_4 , \g236041/u3_syn_4 , \g236049/u3_syn_4 , \g236057/u3_syn_4 , \g236065/u3_syn_4 , \g236073/u3_syn_4 , \g236081/u3_syn_4 , \g236089/u3_syn_4 , \g236097/u3_syn_4 , \g236105/u3_syn_4 , \g236113/u3_syn_4 , \g236121/u3_syn_4 , \g236129/u3_syn_4 , \g236137/u3_syn_4 , \g236145/u3_syn_4 , \g236153/u3_syn_4 , \g236161/u3_syn_4 , \g236169/u3_syn_4 , \g236177/u3_syn_4 , \g236185/u3_syn_4 , \g236193/u3_syn_4 , \g236196/u3_syn_4 , \g236198/u3_syn_4 , \g236203/u3_syn_4 , \g236211/u3_syn_4 , \g236219/u3_syn_4 , \g236220/u3_syn_4 , \g236229/u3_syn_4 , \g236232/u3_syn_4 , \g236238/u3_syn_4 , \g236246/u3_syn_4 , \g236255/u3_syn_4 , \g236263/u3_syn_4 , \g236271/u3_syn_4 , \g236275/u3_syn_4 , \g236280/u3_syn_4 , \g236288/u3_syn_4 , \g236296/u3_syn_4 , \g236304/u3_syn_4 , \g236305/u3_syn_4 , \g236306/u3_syn_4 , \g236315/u3_syn_4 , \g236323/u3_syn_4 , \g236331/u3_syn_4 , \g236334/u3_syn_4 , \g236340/u3_syn_4 , \g236348/u3_syn_4 , \g236357/u3_syn_4 , \g236359/u3_syn_4 , \g236367/u3_syn_4 , \g236374/u3_syn_4 , \g236376/u3_syn_4 , \g236377/u3_syn_4 , \g236385/u3_syn_4 , \g236393/u3_syn_4 , \g236402/u3_syn_4 , \g236410/u3_syn_4 , \g236419/u3_syn_4 , \g236427/u3_syn_4 , \g236433/u3_syn_4 , \g236436/u3_syn_4 , \g236444/u3_syn_4 , \g236452/u3_syn_4 , \g236460/u3_syn_4 , \g236468/u3_syn_4 , \g236476/u3_syn_4 , \g236484/u3_syn_4 , \g236492/u3_syn_4 , \g236500/u3_syn_4 , \g236508/u3_syn_4 , \g236516/u3_syn_4 , \g236518/u3_syn_4 , \g236525/u3_syn_4 , \g236533/u3_syn_4 , \g236542/u3_syn_4 , \g236550/u3_syn_4 , \g236559/u3_syn_4 , \g236567/u3_syn_4 , \g236575/u3_syn_4 , \g236583/u3_syn_4 , \g236591/u3_syn_4 , \g236599/u3_syn_4 , \g236607/u3_syn_4 , \g236608/u3_syn_4 , \g236616/u3_syn_4 , \g236624/u3_syn_4 , \g236632/u3_syn_4 , \g236640/u3_syn_4 , \g236647/u3_syn_4 , \g236649/u3_syn_4 , \g236659/u3_syn_4 , \g236671/u3_syn_4 , \g236677/u3_syn_4 , \g236688/u3_syn_4 , \g236696/u3_syn_4 , \g236705/u3_syn_4 , \g236712/u3_syn_4 , \g236718/u3_syn_4 , \g236729/u3_syn_4 , \g236732/u3_syn_4 , \g236745/u3_syn_4 , \g236753/u3_syn_4 , \g236761/u3_syn_4 , \g236769/u3_syn_4 , \g236777/u3_syn_4 , \g236779/u3_syn_4 , \g236788/u3_syn_4 , \g236800/u3_syn_4 , \g236802/u3_syn_4 , \g236805/u3_syn_4 , \g236813/u3_syn_4 , \g236825/u3_syn_4 , \g236829/u3_syn_4 , \g236837/u3_syn_4 , \g236849/u3_syn_4 , \g236854/u3_syn_4 , \g236860/u3_syn_4 , \g236872/u3_syn_4 , \g236878/u3_syn_4 , \g236884/u3_syn_4 , \g236896/u3_syn_4 , \g236903/u3_syn_4 , \g236908/u3_syn_4 , \g236920/u3_syn_4 , \g236930/u3_syn_4 , \g236939/u3_syn_4 , \g236947/u3_syn_4 , \g236949/u3_syn_4 , \g236956/u3_syn_4 , \g236962/u3_syn_4 , \g236965/u3_syn_4 , \g236980/u3_syn_4 , \g236988/u3_syn_4 , \g236989/u3_syn_4 , \g237004/u3_syn_4 , \g237005/u3_syn_4 , \g237020/u3_syn_4 , \g237021/u3_syn_4 , \g237033/u3_syn_4 , \g237044/u3_syn_4 , \g237045/u3_syn_4 , \g237056/u3_syn_4 , \g237068/u3_syn_4 , \g237076/u3_syn_4 , \g237084/u3_syn_4 , \g237092/u3_syn_4 , \g237095/u3_syn_4 , \g237107/u3_syn_4 , \g237110/u3_syn_4 , \g237119/u3_syn_4 , \g237131/u3_syn_4 , \g237135/u3_syn_4 , \g237148/u3_syn_4 , \g237152/u3_syn_4 , \g237165/u3_syn_4 , \g237168/u3_syn_4 , \g237180/u3_syn_4 , \g237185/u3_syn_4 , \g237192/u3_syn_4 , \g237204/u3_syn_4 , \g237209/u3_syn_4 , \g237215/u3_syn_4 , \g237229/u3_syn_4 , \g237231/u3_syn_4 , \g237245/u3_syn_4 , \g237251/u3_syn_4 , \g237260/u3_syn_4 , \g237262/u3_syn_4 , \g237277/u3_syn_4 , \g237281/u3_syn_4 , \g237293/u3_syn_4 , \g237294/u3_syn_4 , \g237310/u3_syn_4 , \g237311/u3_syn_4 , \g237323/u3_syn_4 , \g237334/u3_syn_4 , \g237342/u3_syn_4 , \g237350/u3_syn_4 , \g237353/u3_syn_4 , \g237359/u3_syn_4 , \g237367/u3_syn_4 , \g237368/u3_syn_4 , \g237378/u3_syn_4 , \g237391/u3_syn_4 , \g237392/u3_syn_4 , \g237403/u3_syn_4 , \g237415/u3_syn_4 , \g237417/u3_syn_4 , \g237431/u3_syn_4 , \g237439/u3_syn_4 , \g237440/u3_syn_4 , \g237454/u3_syn_4 , \g237457/u3_syn_4 , \g237472/u3_syn_4 , \g237480/u3_syn_4 , \g237488/u3_syn_4 , \g237496/u3_syn_4 , \g237499/u3_syn_4 , \g237512/u3_syn_4 , \g237515/u3_syn_4 , \g237525/u3_syn_4 , \g237529/u3_syn_4 , \g237535/u3_syn_4 , \g237541/u3_syn_4 , \g237553/u3_syn_4 , \g237561/u3_syn_4 , \g237569/u3_syn_4 , \g237575/u3_syn_4 , \g237578/u3_syn_4 , \g237581/u3_syn_4 , \g237591/u3_syn_4 , \g237602/u3_syn_4 , \g237610/u3_syn_4 , \g237617/u3_syn_4 , \g237623/u3_syn_4 , \g237633/u3_syn_4 , \g237635/u3_syn_4 , \g237648/u3_syn_4 , \g237658/u3_syn_4 , \g237659/u3_syn_4 , \g237660/u3_syn_4 , \g237668/u3_syn_4 , \g237675/u3_syn_4 , \g237684/u3_syn_4 , \g237692/u3_syn_4 , \g237693/u3_syn_4 , \g237705/u3_syn_4 , \g237716/u3_syn_4 , \g237717/u3_syn_4 , \g237729/u3_syn_4 , \g237740/u3_syn_4 , \g237741/u3_syn_4 , \g237756/u3_syn_4 , \g237764/u3_syn_4 , \g237768/u3_syn_4 , \g237780/u3_syn_4 , \g237782/u3_syn_4 , \g237792/u3_syn_4 , \g237804/u3_syn_4 , \g237812/u3_syn_4 , \g237820/u3_syn_4 , \g237828/u3_syn_4 , \g237836/u3_syn_4 , \g237844/u3_syn_4 , \g237852/u3_syn_4 , \g237860/u3_syn_4 , \g237868/u3_syn_4 , \g237876/u3_syn_4 , \g237884/u3_syn_4 , \g237888/u3_syn_4 , \g237895/u3_syn_4 , \g237907/u3_syn_4 , \g237916/u3_syn_4 , \g237924/u3_syn_4 , \g237931/u3_syn_4 , \g237940/u3_syn_4 , \g237949/u3_syn_4 , \g237950/u3_syn_4 , \g237955/u3_syn_4 , \g237961/u3_syn_4 , \g237965/u3_syn_4 , \g237975/u3_syn_4 , \g237983/u3_syn_4 , \g237989/u3_syn_4 , \g237999/u3_syn_4 , \g238007/u3_syn_4 , \g238015/u3_syn_4 , \g238017/u3_syn_4 , \g238033/u3_syn_4 , \g238035/u3_syn_4 , \g238049/u3_syn_4 , \g238057/u3_syn_4 , \g238065/u3_syn_4 , \g238072/u3_syn_4 , \g238081/u3_syn_4 , \g238082/u3_syn_4 , \g238097/u3_syn_4 , \g238105/u3_syn_4 , \g238113/u3_syn_4 , \g238114/u3_syn_4 , \g238129/u3_syn_4 , \g238137/u3_syn_4 , \g238145/u3_syn_4 , \g238153/u3_syn_4 , \g238161/u3_syn_4 , \g238163/u3_syn_4 , \g238177/u3_syn_4 , \g238179/u3_syn_4 , \g238194/u3_syn_4 , \g238197/u3_syn_4 , \g238209/u3_syn_4 , \g238213/u3_syn_4 , \g238225/u3_syn_4 , \g238229/u3_syn_4 , \g238237/u3_syn_4 , \g238250/u3_syn_4 , \g238257/u3_syn_4 , \g238263/u3_syn_4 , \g238269/u3_syn_4 , \g238282/u3_syn_4 , \g238285/u3_syn_4 , \g238298/u3_syn_4 , \g238301/u3_syn_4 , \g238314/u3_syn_4 , \g238316/u3_syn_4 , \g238329/u3_syn_4 , \g238338/u3_syn_4 , \g238346/u3_syn_4 , \g238351/u3_syn_4 , \g238356/u3_syn_4 , \g238368/u3_syn_4 , \g238378/u3_syn_4 , \g238386/u3_syn_4 , \g238394/u3_syn_4 , \g238402/u3_syn_4 , \g238409/u3_syn_4 , \g238412/u3_syn_4 , \g238427/u3_syn_4 , \g238429/u3_syn_4 , \g238443/u3_syn_4 , \g238448/u3_syn_4 , \g238457/u3_syn_4 , \g238460/u3_syn_4 , \g238472/u3_syn_4 , \g238484/u3_syn_4 , \g238492/u3_syn_4 , \g238500/u3_syn_4 , \g238505/u3_syn_4 , \g238516/u3_syn_4 , \g238524/u3_syn_4 , \g238532/u3_syn_4 , \g238534/u3_syn_4 , \g238544/u3_syn_4 , \g238549/u3_syn_4 , \g238550/u3_syn_4 , \g238565/u3_syn_4 , \g238566/u3_syn_4 , \g238582/u3_syn_4 , \g238583/u3_syn_4 , \g238594/u3_syn_4 , \g238606/u3_syn_4 , \g238614/u3_syn_4 , \g238615/u3_syn_4 , \g238619/u3_syn_4 , \g238631/u3_syn_4 , \g238639/u3_syn_4 , \g238647/u3_syn_4 , \g238649/u3_syn_4 , \g238659/u3_syn_4 , \g238670/u3_syn_4 , \g238671/u3_syn_4 , \g238680/u3_syn_4 , \g238688/u3_syn_4 , \g238691/u3_syn_4 , \g238696/u3_syn_4 , \g238705/u3_syn_4 , \g238708/u3_syn_4 , \g238721/u3_syn_4 , \g238724/u3_syn_4 , \g238736/u3_syn_4 , \g238745/u3_syn_4 , \g238753/u3_syn_4 , \g238757/u3_syn_4 , \g238764/u3_syn_4 , \g238776/u3_syn_4 , \g238781/u3_syn_4 , \g238787/u3_syn_4 , \g238799/u3_syn_4 , \g238807/u3_syn_4 , \g238811/u3_syn_4 , \g238824/u3_syn_4 , \g238830/u3_syn_4 , \g238841/u3_syn_4 , \g238843/u3_syn_4 , \g238855/u3_syn_4 , \g238859/u3_syn_4 , \g238863/u3_syn_4 , \g238868/u3_syn_4 , \g238880/u3_syn_4 , \g238888/u3_syn_4 , \g238892/u3_syn_4 , \g238903/u3_syn_4 , \g238911/u3_syn_4 , \g238915/u3_syn_4 , \g238927/u3_syn_4 , \g238937/u3_syn_4 , \g238945/u3_syn_4 , \g238953/u3_syn_4 , \g238961/u3_syn_4 , \g238970/u3_syn_4 , \g238971/u3_syn_4 , \g238983/u3_syn_4 , \g238994/u3_syn_4 , \g239002/u3_syn_4 , \g239009/u3_syn_4 , \g239015/u3_syn_4 , \g239025/u3_syn_4 , \g239030/u3_syn_4 , \g239041/u3_syn_4 , \g239048/u3_syn_4 , \g239053/u3_syn_4 , \g239065/u3_syn_4 , \g239073/u3_syn_4 , \g239081/u3_syn_4 , \g239082/u3_syn_4 , \g239093/u3_syn_4 , \g239105/u3_syn_4 , \g239108/u3_syn_4 , \g239117/u3_syn_4 , \g239129/u3_syn_4 , \g239137/u3_syn_4 , \g239139/u3_syn_4 , \g239148/u3_syn_4 , \g239160/u3_syn_4 , \g239162/u3_syn_4 , \g239172/u3_syn_4 , \g239184/u3_syn_4 , \g239187/u3_syn_4 , \g239189/u3_syn_4 , \g239201/u3_syn_4 , \g239208/u3_syn_4 , \g239217/u3_syn_4 , \g239219/u3_syn_4 , \g239226/u3_syn_4 , \g239234/u3_syn_4 , \g239242/u3_syn_4 , \g239246/u3_syn_4 , \g239257/u3_syn_4 , \g239258/u3_syn_4 , \g239263/u3_syn_4 , \g239275/u3_syn_4 , \g239277/u3_syn_4 , \g239291/u3_syn_4 , \g239296/u3_syn_4 , \g239308/u3_syn_4 , \g239311/u3_syn_4 , \g239322/u3_syn_4 , \g239329/u3_syn_4 , \g239338/u3_syn_4 , \g239339/u3_syn_4 , \g239346/u3_syn_4 , \g239351/u3_syn_4 , \g239363/u3_syn_4 , \g239370/u3_syn_4 , \g239375/u3_syn_4 , \g239387/u3_syn_4 , \g239395/u3_syn_4 , \g239418/u3_syn_4 , \g239439/u3_syn_4 , \g239442/u3_syn_4 , \g239454/u3_syn_4 , \g239464/u3_syn_4 , \g239470/u3_syn_4 , \g239481/u3_syn_4 , \g239487/u3_syn_4 , \g239497/u3_syn_4 , \g239520/u3_syn_4 , \g239532/u3_syn_4 , \g239543/u3_syn_4 , \g239551/u3_syn_4 , \g239552/u3_syn_4 , \g239567/u3_syn_4 , \g239575/u3_syn_4 , \g239579/u3_syn_4 , \g239592/u3_syn_4 , \g239594/u3_syn_4 , \g239608/u3_syn_4 , \g239626/u3_syn_4 , \g239634/u3_syn_4 , \g239646/u3_syn_4 , \g239649/u3_syn_4 , \g239657/u3_syn_4 , \g239670/u3_syn_4 , \g239673/u3_syn_4 , \g239686/u3_syn_4 , \g239694/u3_syn_4 , \g239695/u3_syn_4 , \g239701/u3_syn_4 , \g239705/u3_syn_4 , \g239709/u3_syn_4 , \g239715/u3_syn_4 , \g239717/u3_syn_4 , \g239726/u3_syn_4 , \g239734/u3_syn_4 , \g239735/u3_syn_4 , \g239743/u3_syn_4 , \g239760/u3_syn_4 , \g239768/u3_syn_4 , \g239776/u3_syn_4 , \g239784/u3_syn_4 , \g239793/u3_syn_4 , \g239801/u3_syn_4 , \g239817/u3_syn_4 , \g239818/u3_syn_4 , \g239848/u3_syn_4 , \g239856/u3_syn_4 , \g239872/u3_syn_4 , \g239880/u3_syn_4 , \g239888/u3_syn_4 , \g239896/u3_syn_4 , \g239904/u3_syn_4 , \g239912/u3_syn_4 , \g239920/u3_syn_4 , \g239928/u3_syn_4 , \g239936/u3_syn_4 , \g239951/u3_syn_4 , \g239963/u3_syn_4 , \g239979/u3_syn_4 , \g239986/u3_syn_4 , \g239999/u3_syn_4 , \g240000/u3_syn_4 , \g240008/u3_syn_4 , \g240012/u3_syn_4 , \g240018/u3_syn_4 , \g240026/u3_syn_4 , \g240034/u3_syn_4 , \g240042/u3_syn_4 , \g240050/u3_syn_4 , \g240074/u3_syn_4 , \g240091/u3_syn_4 , \g240122/u3_syn_4 , \g240147/u3_syn_4 , \g240209/u3_syn_4 , \g240219/u3_syn_4 , \g240259/u3_syn_4 , \g240334/u3_syn_4 , \g240406/u3_syn_4 , \g240416/u3_syn_4 , \g240424/u3_syn_4 , \g240432/u3_syn_4 , \g240440/u3_syn_4 , \g240448/u3_syn_4 , \g240456/u3_syn_4 , \g240464/u3_syn_4 , \g240472/u3_syn_4 , \g240480/u3_syn_4 , \g240488/u3_syn_4 , \g240496/u3_syn_4 , \g240504/u3_syn_4 , \g240512/u3_syn_4 , \g240520/u3_syn_4 , \g240530/u3_syn_4 , \g240538/u3_syn_4 , \g240547/u3_syn_4 , \g240555/u3_syn_4 , \g240563/u3_syn_4 , \g240571/u3_syn_4 , \g240579/u3_syn_4 , \g240587/u3_syn_4 , \g240595/u3_syn_4 , \g240603/u3_syn_4 , \g240611/u3_syn_4 , \g240619/u3_syn_4 , \g240627/u3_syn_4 , \g240635/u3_syn_4 , \g240643/u3_syn_4 , \g240651/u3_syn_4 , \g240659/u3_syn_4 , \g240667/u3_syn_4 , \g240675/u3_syn_4 , \g240683/u3_syn_4 , \g240691/u3_syn_4 , \g240699/u3_syn_4 , \g240707/u3_syn_4 , \g240715/u3_syn_4 , \g240723/u3_syn_4 , \g240731/u3_syn_4 , \g240739/u3_syn_4 , \g240747/u3_syn_4 , \g240755/u3_syn_4 , \g240763/u3_syn_4 , \g240771/u3_syn_4 , \g240779/u3_syn_4 , \g240787/u3_syn_4 , \g240795/u3_syn_4 , \g240803/u3_syn_4 , \g240811/u3_syn_4 , \g240819/u3_syn_4 , \g240827/u3_syn_4 , \g240835/u3_syn_4 , \g240843/u3_syn_4 , \g240851/u3_syn_4 , \g240859/u3_syn_4 , \g240867/u3_syn_4 , \g240875/u3_syn_4 , \g240883/u3_syn_4 , \g240891/u3_syn_4 , \g240899/u3_syn_4 , \g240907/u3_syn_4 , \g240915/u3_syn_4 , \g240923/u3_syn_4 , \g240931/u3_syn_4 , \g240939/u3_syn_4 , \g240947/u3_syn_4 , \g240955/u3_syn_4 , \g240963/u3_syn_4 , \g240971/u3_syn_4 , \g240979/u3_syn_4 , \g240987/u3_syn_4 , \g240995/u3_syn_4 , \g241003/u3_syn_4 , \g241011/u3_syn_4 , \g241019/u3_syn_4 , \g241027/u3_syn_4 , \g241036/u3_syn_4 , \g241044/u3_syn_4 , \g241052/u3_syn_4 , \g241060/u3_syn_4 , \g241068/u3_syn_4 , \g241076/u3_syn_4 , \g241084/u3_syn_4 , \g241092/u3_syn_4 , \g241100/u3_syn_4 , \g241108/u3_syn_4 , \g241116/u3_syn_4 , \g241124/u3_syn_4 , \g241132/u3_syn_4 , \g241140/u3_syn_4 , \g241148/u3_syn_4 , \g241156/u3_syn_4 , \g241164/u3_syn_4 , \g241172/u3_syn_4 , \g241180/u3_syn_4 , \g241188/u3_syn_4 , \g241196/u3_syn_4 , \g241205/u3_syn_4 , \g241213/u3_syn_4 , \g241221/u3_syn_4 , \g241229/u3_syn_4 , \g241237/u3_syn_4 , \g241245/u3_syn_4 , \g241253/u3_syn_4 , \g241261/u3_syn_4 , \g241269/u3_syn_4 , \g241277/u3_syn_4 , \g241285/u3_syn_4 , \g241293/u3_syn_4 , \g241301/u3_syn_4 , \g241309/u3_syn_4 , \g241317/u3_syn_4 , \g241325/u3_syn_4 , \g241333/u3_syn_4 , \g241341/u3_syn_4 , \g241349/u3_syn_4 , \g241358/u3_syn_4 , \g241366/u3_syn_4 , \g241374/u3_syn_4 , \g241382/u3_syn_4 , \g241390/u3_syn_4 , \g241398/u3_syn_4 , \g241406/u3_syn_4 , \g241415/u3_syn_4 , \g241424/u3_syn_4 , \g241433/u3_syn_4 , \g241441/u3_syn_4 , \g241449/u3_syn_4 , \g241459/u3_syn_4 , \g241470/u3_syn_4 , \g241480/u3_syn_4 , \g241489/u3_syn_4 , \g241497/u3_syn_4 , \g241505/u3_syn_4 , \g241513/u3_syn_4 , \g241545/_3_ , \g241580/_00_ , \g241737/_0_ , \g241752/_0_ , \g241755/_0_ , \g241767/_2__syn_2 , \g241781/_1__syn_2 , \g241782/_0_ , \g241803/_1__syn_2 , \g241805/_0_ , \g241812/_1__syn_2 , \g241814/_1__syn_2 , \g241816/_1__syn_2 , \g241819/_1__syn_2 , \g241822/_1__syn_2 , \g241823/_0_ , \g241833/_1__syn_2 , \g241843/_1__syn_2 , \g241844/_1__syn_2 , \g241848/_1__syn_2 , \g241855/_1__syn_2 , \g241868/_1__syn_2 , \g242013/_1__syn_2 , \g242015/_1__syn_2 , \g242017/_1__syn_2 , \g242021/_1__syn_2 , \g242039/_1__syn_2 , \g242081/_0_ , \g242086/_0_ , \g242101/_3_ , \g242116/_0_ , \g242135/_2_ , \g242147/_0_ , \g242158/_0_ , \g242196/_0_ , \g242202/_0_ , \g242203/_0_ , \g242204/_0_ , \g242212/_0_ , \g242226/_01_ , \g242281/_0_ , \g242407/_0_ , \g242410/_0_ , \g242426/_0_ , \g242438/_2_ , \g242466/_0_ , \g242530/_0_ , \g242532/_0_ , \g243397/_0_ , \g245925/_0_ , \g245932/_0_ , \g245933/_0_ , \g245986/_3_ , \g250157/_3_ , \g250202/_0_ , \g250246/_1_ , \g250248/_0_ , \g250250/_0_ , \g250305/_0_ , \g250323/_0_ , \g250373/_0_ , \g250377/_0_ , \g250412/_0_ , \g250413/_0_ , \g250418/_0_ , \g250419/_0_ , \g250421/_0_ , \g250433/_0_ , \g250448/_3_ , \g250567/_3_ , \g258965/_0_ , \g259006/_0_ , \g259471/_0_ , \g259473/_2_ , \g260557/_0_ , \g261035/_0_ , \g261095/_3_ , \g261207/_2__syn_2 , \g261754/_0_ , \g262017/_0_ , \g262045/_0_ , \g262046/_0_ , \g262100/_3_ , \g263539/_1_ , \g263574/_0_ , \g263858/_0_ , \g264104/_1_ , \g264107/_1_ , \g264117/_0_ , \g264282/_0_ , \g264511/_0_ , \g264541/_0_ , \g264562/_0_ , \g264618/_0_ , \g264660/_0_ , \g264681/_3_ , \g264727/_0_ , \g265013/_0_ , \g265084/_0_ , \g265378/_0_ , \g265413/_0_ , \g265446/_0_ , \g265486/_0_ , \g265524/_3_ , \g265528/_3_ , \g265548/_3_ , \g265579/_0_ , \g265768/_0_ , \g265801/_0_ , \g265819/_1_ , \g265853/_0_ , \g265933/_0_ , \g266022/_0_ , \g266183/_1_ , \g281909/_0_ , \g281965/_1_ , \g282284/_1_ , \g282639/_1_ , \g283047/_0_ , \g283157/_1_ , \g283184/_0_ , \g283334/_3_ , int_o_pad, \m_wb_adr_o[0]_pad , \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131_syn_2 , \wishbone_tx_fifo_fifo_reg[2][15]/P0001_reg_syn_3 , \wishbone_tx_fifo_fifo_reg[2][16]/P0001_reg_syn_3 , \wishbone_tx_fifo_fifo_reg[2][17]/P0001_reg_syn_3 , \wishbone_tx_fifo_fifo_reg[2][22]/P0001_reg_syn_3 , \wishbone_tx_fifo_fifo_reg[2][23]/P0001_reg_syn_3 , \wishbone_tx_fifo_fifo_reg[2][25]/P0001_reg_syn_3 , \wishbone_tx_fifo_fifo_reg[2][2]/P0001_reg_syn_3 );
	input \CarrierSense_Tx2_reg/NET0131  ;
	input \Collision_Tx1_reg/NET0131  ;
	input \Collision_Tx2_reg/NET0131  ;
	input \RstTxPauseRq_reg/NET0131  ;
	input \RxAbortRst_reg/NET0131  ;
	input \RxAbort_latch_reg/NET0131  ;
	input \RxAbort_wb_reg/NET0131  ;
	input \RxEnSync_reg/NET0131  ;
	input \TPauseRq_reg/NET0131  ;
	input \TxPauseRq_sync2_reg/NET0131  ;
	input \TxPauseRq_sync3_reg/NET0131  ;
	input \WillSendControlFrame_sync2_reg/NET0131  ;
	input \WillSendControlFrame_sync3_reg/NET0131  ;
	input \WillTransmit_q2_reg/P0001  ;
	input \ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_COLLCONF_2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_COLLCONF_2_DataOut_reg[1]/NET0131  ;
	input \ethreg1_COLLCONF_2_DataOut_reg[2]/NET0131  ;
	input \ethreg1_COLLCONF_2_DataOut_reg[3]/NET0131  ;
	input \ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_INT_MASK_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_INT_MASK_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_INT_MASK_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_INT_MASK_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_INT_MASK_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_INT_MASK_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_INT_MASK_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_IPGR1_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_IPGR1_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_IPGR1_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_IPGR1_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_IPGR1_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_IPGR1_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_IPGR1_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_IPGR2_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_IPGR2_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_IPGR2_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_IPGR2_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_IPGR2_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_IPGR2_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_IPGR2_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_IPGT_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_IPGT_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_IPGT_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_IPGT_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_IPGT_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_IPGT_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_IPGT_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MIIADDRESS_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIIADDRESS_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MIIADDRESS_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MIIADDRESS_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MIIADDRESS_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MIIADDRESS_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIIADDRESS_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MIIADDRESS_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MIIADDRESS_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MIIADDRESS_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MIICOMMAND0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIICOMMAND1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIICOMMAND2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MIIMODER_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[10]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[11]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[12]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[13]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[14]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[15]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[8]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[9]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MODER_2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[7]/NET0131  ;
	input \ethreg1_ResetRxCIrq_sync2_reg/NET0131  ;
	input \ethreg1_ResetRxCIrq_sync3_reg/NET0131  ;
	input \ethreg1_ResetTxCIrq_sync2_reg/NET0131  ;
	input \ethreg1_SetRxCIrq_reg/NET0131  ;
	input \ethreg1_SetRxCIrq_rxclk_reg/NET0131  ;
	input \ethreg1_SetRxCIrq_sync2_reg/NET0131  ;
	input \ethreg1_SetRxCIrq_sync3_reg/NET0131  ;
	input \ethreg1_SetTxCIrq_reg/NET0131  ;
	input \ethreg1_SetTxCIrq_sync2_reg/NET0131  ;
	input \ethreg1_SetTxCIrq_sync3_reg/NET0131  ;
	input \ethreg1_SetTxCIrq_txclk_reg/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_TXCTRL_2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_irq_busy_reg/NET0131  ;
	input \ethreg1_irq_rxb_reg/NET0131  ;
	input \ethreg1_irq_rxc_reg/NET0131  ;
	input \ethreg1_irq_rxe_reg/NET0131  ;
	input \ethreg1_irq_txb_reg/NET0131  ;
	input \ethreg1_irq_txc_reg/NET0131  ;
	input \ethreg1_irq_txe_reg/NET0131  ;
	input m_wb_ack_i_pad ;
	input \m_wb_adr_o[10]_pad  ;
	input \m_wb_adr_o[11]_pad  ;
	input \m_wb_adr_o[12]_pad  ;
	input \m_wb_adr_o[13]_pad  ;
	input \m_wb_adr_o[14]_pad  ;
	input \m_wb_adr_o[15]_pad  ;
	input \m_wb_adr_o[16]_pad  ;
	input \m_wb_adr_o[17]_pad  ;
	input \m_wb_adr_o[18]_pad  ;
	input \m_wb_adr_o[19]_pad  ;
	input \m_wb_adr_o[20]_pad  ;
	input \m_wb_adr_o[21]_pad  ;
	input \m_wb_adr_o[22]_pad  ;
	input \m_wb_adr_o[23]_pad  ;
	input \m_wb_adr_o[24]_pad  ;
	input \m_wb_adr_o[25]_pad  ;
	input \m_wb_adr_o[26]_pad  ;
	input \m_wb_adr_o[27]_pad  ;
	input \m_wb_adr_o[28]_pad  ;
	input \m_wb_adr_o[29]_pad  ;
	input \m_wb_adr_o[2]_pad  ;
	input \m_wb_adr_o[30]_pad  ;
	input \m_wb_adr_o[31]_pad  ;
	input \m_wb_adr_o[3]_pad  ;
	input \m_wb_adr_o[4]_pad  ;
	input \m_wb_adr_o[5]_pad  ;
	input \m_wb_adr_o[6]_pad  ;
	input \m_wb_adr_o[7]_pad  ;
	input \m_wb_adr_o[8]_pad  ;
	input \m_wb_adr_o[9]_pad  ;
	input \m_wb_dat_i[10]_pad  ;
	input \m_wb_dat_i[11]_pad  ;
	input \m_wb_dat_i[12]_pad  ;
	input \m_wb_dat_i[13]_pad  ;
	input \m_wb_dat_i[14]_pad  ;
	input \m_wb_dat_i[15]_pad  ;
	input \m_wb_dat_i[16]_pad  ;
	input \m_wb_dat_i[17]_pad  ;
	input \m_wb_dat_i[18]_pad  ;
	input \m_wb_dat_i[19]_pad  ;
	input \m_wb_dat_i[1]_pad  ;
	input \m_wb_dat_i[20]_pad  ;
	input \m_wb_dat_i[22]_pad  ;
	input \m_wb_dat_i[23]_pad  ;
	input \m_wb_dat_i[24]_pad  ;
	input \m_wb_dat_i[25]_pad  ;
	input \m_wb_dat_i[26]_pad  ;
	input \m_wb_dat_i[27]_pad  ;
	input \m_wb_dat_i[28]_pad  ;
	input \m_wb_dat_i[29]_pad  ;
	input \m_wb_dat_i[2]_pad  ;
	input \m_wb_dat_i[30]_pad  ;
	input \m_wb_dat_i[31]_pad  ;
	input \m_wb_dat_i[3]_pad  ;
	input \m_wb_dat_i[4]_pad  ;
	input \m_wb_dat_i[5]_pad  ;
	input \m_wb_dat_i[6]_pad  ;
	input \m_wb_dat_i[7]_pad  ;
	input \m_wb_dat_i[8]_pad  ;
	input m_wb_err_i_pad ;
	input \m_wb_sel_o[0]_pad  ;
	input \m_wb_sel_o[1]_pad  ;
	input \m_wb_sel_o[2]_pad  ;
	input \m_wb_sel_o[3]_pad  ;
	input m_wb_stb_o_pad ;
	input m_wb_we_o_pad ;
	input \maccontrol1_MuxedAbort_reg/NET0131  ;
	input \maccontrol1_MuxedDone_reg/NET0131  ;
	input \maccontrol1_TxAbortInLatched_reg/NET0131  ;
	input \maccontrol1_TxDoneInLatched_reg/NET0131  ;
	input \maccontrol1_TxUsedDataOutDetected_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_AddressOK_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[0]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[10]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[11]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[12]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[13]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[14]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[15]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[1]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[2]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[3]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[4]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[5]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[6]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[7]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[8]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[9]/NET0131  ;
	input \maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131  ;
	input \maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131  ;
	input \maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131  ;
	input \maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131  ;
	input \maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131  ;
	input \maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_Divider2_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_DlyCrcCnt_reg[0]/NET0131  ;
	input \maccontrol1_receivecontrol1_DlyCrcCnt_reg[1]/NET0131  ;
	input \maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[0]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[10]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[11]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[12]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[13]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[14]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[15]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[1]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[2]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[3]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[4]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[5]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[6]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[7]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[8]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[9]/NET0131  ;
	input \maccontrol1_receivecontrol1_OpCodeOK_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimerEq0_sync2_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[11]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[12]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[14]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[15]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[1]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[5]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[8]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131  ;
	input \maccontrol1_receivecontrol1_Pause_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_SlotTimer_reg[0]/NET0131  ;
	input \maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131  ;
	input \maccontrol1_receivecontrol1_SlotTimer_reg[2]/NET0131  ;
	input \maccontrol1_receivecontrol1_SlotTimer_reg[3]/NET0131  ;
	input \maccontrol1_receivecontrol1_SlotTimer_reg[4]/NET0131  ;
	input \maccontrol1_receivecontrol1_SlotTimer_reg[5]/NET0131  ;
	input \maccontrol1_receivecontrol1_TypeLengthOK_reg/NET0131  ;
	input \maccontrol1_transmitcontrol1_BlockTxDone_reg/NET0131  ;
	input \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[0]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[1]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[2]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[3]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[4]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[5]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[6]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[7]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlEnd_q_reg/P0001  ;
	input \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  ;
	input \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131  ;
	input \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[1]/NET0131  ;
	input \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131  ;
	input \maccontrol1_transmitcontrol1_SendingCtrlFrm_reg/NET0131  ;
	input \maccontrol1_transmitcontrol1_TxCtrlEndFrm_reg/NET0131  ;
	input \maccontrol1_transmitcontrol1_TxCtrlStartFrm_q_reg/P0001  ;
	input \maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131  ;
	input \maccontrol1_transmitcontrol1_TxUsedDataIn_q_reg/NET0131  ;
	input \maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131  ;
	input \macstatus1_CarrierSenseLost_reg/NET0131  ;
	input \macstatus1_DeferLatched_reg/NET0131  ;
	input \macstatus1_DribbleNibble_reg/NET0131  ;
	input \macstatus1_InvalidSymbol_reg/NET0131  ;
	input \macstatus1_LatchedCrcError_reg/NET0131  ;
	input \macstatus1_LatchedMRxErr_reg/NET0131  ;
	input \macstatus1_LateCollLatched_reg/P0002  ;
	input \macstatus1_LoadRxStatus_reg/NET0131  ;
	input \macstatus1_ReceiveEnd_reg/NET0131  ;
	input \macstatus1_ReceivedPacketTooBig_reg/NET0131  ;
	input \macstatus1_RetryCntLatched_reg[0]/P0002  ;
	input \macstatus1_RetryCntLatched_reg[1]/P0002  ;
	input \macstatus1_RetryCntLatched_reg[2]/P0002  ;
	input \macstatus1_RetryCntLatched_reg[3]/P0002  ;
	input \macstatus1_RetryLimit_reg/P0002  ;
	input \macstatus1_RxColWindow_reg/NET0131  ;
	input \macstatus1_RxLateCollision_reg/NET0131  ;
	input \macstatus1_ShortFrame_reg/NET0131  ;
	input mcoll_pad_i_pad ;
	input md_pad_i_pad ;
	input mdc_pad_o_pad ;
	input \miim1_BitCounter_reg[0]/NET0131  ;
	input \miim1_BitCounter_reg[1]/NET0131  ;
	input \miim1_BitCounter_reg[2]/NET0131  ;
	input \miim1_BitCounter_reg[3]/NET0131  ;
	input \miim1_BitCounter_reg[4]/NET0131  ;
	input \miim1_BitCounter_reg[5]/NET0131  ;
	input \miim1_BitCounter_reg[6]/NET0131  ;
	input \miim1_EndBusy_reg/NET0131  ;
	input \miim1_InProgress_q1_reg/NET0131  ;
	input \miim1_InProgress_q2_reg/NET0131  ;
	input \miim1_InProgress_q3_reg/NET0131  ;
	input \miim1_InProgress_reg/NET0131  ;
	input \miim1_LatchByte0_d_reg/NET0131  ;
	input \miim1_LatchByte1_d_reg/NET0131  ;
	input \miim1_LatchByte_reg[0]/NET0131  ;
	input \miim1_LatchByte_reg[1]/NET0131  ;
	input \miim1_Nvalid_reg/NET0131  ;
	input \miim1_RStatStart_q1_reg/NET0131  ;
	input \miim1_RStatStart_q2_reg/NET0131  ;
	input \miim1_RStatStart_reg/NET0131  ;
	input \miim1_RStat_q2_reg/NET0131  ;
	input \miim1_RStat_q3_reg/NET0131  ;
	input \miim1_ScanStat_q2_reg/NET0131  ;
	input \miim1_SyncStatMdcEn_reg/NET0131  ;
	input \miim1_WCtrlDataStart_q1_reg/NET0131  ;
	input \miim1_WCtrlDataStart_q2_reg/NET0131  ;
	input \miim1_WCtrlDataStart_q_reg/NET0131  ;
	input \miim1_WCtrlDataStart_reg/NET0131  ;
	input \miim1_WCtrlData_q2_reg/NET0131  ;
	input \miim1_WCtrlData_q3_reg/NET0131  ;
	input \miim1_WriteOp_reg/NET0131  ;
	input \miim1_clkgen_Counter_reg[0]/NET0131  ;
	input \miim1_clkgen_Counter_reg[1]/NET0131  ;
	input \miim1_clkgen_Counter_reg[2]/NET0131  ;
	input \miim1_clkgen_Counter_reg[3]/NET0131  ;
	input \miim1_clkgen_Counter_reg[4]/NET0131  ;
	input \miim1_clkgen_Counter_reg[5]/NET0131  ;
	input \miim1_clkgen_Counter_reg[6]/NET0131  ;
	input \miim1_outctrl_Mdo_2d_reg/NET0131  ;
	input \miim1_shftrg_LinkFail_reg/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[0]/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[1]/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[2]/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[3]/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[4]/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[5]/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[6]/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[7]/NET0131  ;
	input \mrxd_pad_i[0]_pad  ;
	input \mrxd_pad_i[1]_pad  ;
	input \mrxd_pad_i[2]_pad  ;
	input \mrxd_pad_i[3]_pad  ;
	input mrxdv_pad_i_pad ;
	input mrxerr_pad_i_pad ;
	input \mtxd_pad_o[0]_pad  ;
	input \mtxd_pad_o[1]_pad  ;
	input \mtxd_pad_o[2]_pad  ;
	input \mtxd_pad_o[3]_pad  ;
	input mtxen_pad_o_pad ;
	input mtxerr_pad_o_pad ;
	input \rxethmac1_Broadcast_reg/NET0131  ;
	input \rxethmac1_CrcHashGood_reg/P0001  ;
	input \rxethmac1_CrcHash_reg[0]/P0001  ;
	input \rxethmac1_CrcHash_reg[1]/P0001  ;
	input \rxethmac1_CrcHash_reg[2]/P0001  ;
	input \rxethmac1_CrcHash_reg[3]/P0001  ;
	input \rxethmac1_CrcHash_reg[4]/P0001  ;
	input \rxethmac1_CrcHash_reg[5]/P0001  ;
	input \rxethmac1_DelayData_reg/NET0131  ;
	input \rxethmac1_LatchedByte_reg[0]/NET0131  ;
	input \rxethmac1_LatchedByte_reg[1]/NET0131  ;
	input \rxethmac1_LatchedByte_reg[2]/NET0131  ;
	input \rxethmac1_LatchedByte_reg[3]/NET0131  ;
	input \rxethmac1_LatchedByte_reg[4]/NET0131  ;
	input \rxethmac1_LatchedByte_reg[5]/NET0131  ;
	input \rxethmac1_LatchedByte_reg[6]/NET0131  ;
	input \rxethmac1_LatchedByte_reg[7]/NET0131  ;
	input \rxethmac1_Multicast_reg/NET0131  ;
	input \rxethmac1_RxData_d_reg[0]/NET0131  ;
	input \rxethmac1_RxData_d_reg[1]/NET0131  ;
	input \rxethmac1_RxData_d_reg[2]/NET0131  ;
	input \rxethmac1_RxData_d_reg[3]/NET0131  ;
	input \rxethmac1_RxData_d_reg[4]/NET0131  ;
	input \rxethmac1_RxData_d_reg[5]/NET0131  ;
	input \rxethmac1_RxData_d_reg[6]/NET0131  ;
	input \rxethmac1_RxData_d_reg[7]/NET0131  ;
	input \rxethmac1_RxData_reg[0]/NET0131  ;
	input \rxethmac1_RxData_reg[1]/NET0131  ;
	input \rxethmac1_RxData_reg[2]/NET0131  ;
	input \rxethmac1_RxData_reg[3]/NET0131  ;
	input \rxethmac1_RxData_reg[4]/NET0131  ;
	input \rxethmac1_RxData_reg[5]/NET0131  ;
	input \rxethmac1_RxData_reg[6]/NET0131  ;
	input \rxethmac1_RxData_reg[7]/NET0131  ;
	input \rxethmac1_RxEndFrm_d_reg/NET0131  ;
	input \rxethmac1_RxEndFrm_reg/NET0131  ;
	input \rxethmac1_RxStartFrm_reg/NET0131  ;
	input \rxethmac1_RxValid_reg/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[0]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[10]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[11]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[12]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[13]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[14]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[15]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[16]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[17]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[18]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[19]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[1]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[20]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[21]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[22]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[23]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[24]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[25]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[26]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[27]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[28]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[29]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[2]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[30]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[31]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[3]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[4]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[5]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[6]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[7]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[8]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[9]/NET0131  ;
	input \rxethmac1_rxaddrcheck1_AddressMiss_reg/NET0131  ;
	input \rxethmac1_rxaddrcheck1_MulticastOK_reg/NET0131  ;
	input \rxethmac1_rxaddrcheck1_RxAbort_reg/NET0131  ;
	input \rxethmac1_rxaddrcheck1_UnicastOK_reg/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  ;
	input \rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131  ;
	input \rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131  ;
	input \rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131  ;
	input \rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131  ;
	input \rxethmac1_rxcounters1_IFGCounter_reg[0]/NET0131  ;
	input \rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131  ;
	input \rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131  ;
	input \rxethmac1_rxcounters1_IFGCounter_reg[3]/NET0131  ;
	input \rxethmac1_rxcounters1_IFGCounter_reg[4]/NET0131  ;
	input \rxethmac1_rxstatem1_StateData0_reg/NET0131  ;
	input \rxethmac1_rxstatem1_StateData1_reg/NET0131  ;
	input \rxethmac1_rxstatem1_StateDrop_reg/NET0131  ;
	input \rxethmac1_rxstatem1_StateIdle_reg/NET0131  ;
	input \rxethmac1_rxstatem1_StatePreamble_reg/NET0131  ;
	input \rxethmac1_rxstatem1_StateSFD_reg/NET0131  ;
	input \txethmac1_ColWindow_reg/NET0131  ;
	input \txethmac1_PacketFinished_q_reg/NET0131  ;
	input \txethmac1_RetryCnt_reg[0]/NET0131  ;
	input \txethmac1_RetryCnt_reg[1]/NET0131  ;
	input \txethmac1_RetryCnt_reg[2]/NET0131  ;
	input \txethmac1_RetryCnt_reg[3]/NET0131  ;
	input \txethmac1_StatusLatch_reg/NET0131  ;
	input \txethmac1_StopExcessiveDeferOccured_reg/NET0131  ;
	input \txethmac1_TxAbort_reg/NET0131  ;
	input \txethmac1_TxDone_reg/NET0131  ;
	input \txethmac1_TxRetry_reg/NET0131  ;
	input \txethmac1_TxUsedData_reg/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[0]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[1]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[2]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[3]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[4]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[5]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[6]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[7]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[8]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[9]/NET0131  ;
	input \txethmac1_random1_x_reg[1]/NET0131  ;
	input \txethmac1_random1_x_reg[2]/NET0131  ;
	input \txethmac1_random1_x_reg[3]/NET0131  ;
	input \txethmac1_random1_x_reg[4]/NET0131  ;
	input \txethmac1_random1_x_reg[5]/NET0131  ;
	input \txethmac1_random1_x_reg[6]/NET0131  ;
	input \txethmac1_random1_x_reg[7]/NET0131  ;
	input \txethmac1_random1_x_reg[8]/NET0131  ;
	input \txethmac1_random1_x_reg[9]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[0]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[10]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[11]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[12]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[13]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[14]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[15]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[1]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[2]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[4]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[5]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[6]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[7]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[8]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[9]/NET0131  ;
	input \txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131  ;
	input \txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131  ;
	input \txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[0]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[10]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[11]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[12]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[13]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[14]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[15]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[1]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[2]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[3]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[4]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[5]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[6]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[7]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[8]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[9]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[0]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[10]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[11]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[12]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[13]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[14]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[15]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[16]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[17]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[18]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[19]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[1]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[20]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[21]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[22]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[23]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[24]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[25]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[26]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[27]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[28]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[29]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[2]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[30]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[31]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[3]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[4]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[5]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[6]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[7]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[8]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[9]/NET0131  ;
	input \txethmac1_txstatem1_Rule1_reg/NET0131  ;
	input \txethmac1_txstatem1_StateBackOff_reg/NET0131  ;
	input \txethmac1_txstatem1_StateData_reg[0]/NET0131  ;
	input \txethmac1_txstatem1_StateData_reg[1]/NET0131  ;
	input \txethmac1_txstatem1_StateDefer_reg/NET0131  ;
	input \txethmac1_txstatem1_StateFCS_reg/NET0131  ;
	input \txethmac1_txstatem1_StateIPG_reg/NET0131  ;
	input \txethmac1_txstatem1_StateIdle_reg/NET0131  ;
	input \txethmac1_txstatem1_StateJam_q_reg/NET0131  ;
	input \txethmac1_txstatem1_StateJam_reg/NET0131  ;
	input \txethmac1_txstatem1_StatePAD_reg/NET0131  ;
	input \txethmac1_txstatem1_StatePreamble_reg/NET0131  ;
	input wb_ack_o_pad ;
	input \wb_adr_i[10]_pad  ;
	input \wb_adr_i[11]_pad  ;
	input \wb_adr_i[2]_pad  ;
	input \wb_adr_i[3]_pad  ;
	input \wb_adr_i[4]_pad  ;
	input \wb_adr_i[5]_pad  ;
	input \wb_adr_i[6]_pad  ;
	input \wb_adr_i[7]_pad  ;
	input \wb_adr_i[8]_pad  ;
	input \wb_adr_i[9]_pad  ;
	input wb_cyc_i_pad ;
	input \wb_dat_i[0]_pad  ;
	input \wb_dat_i[10]_pad  ;
	input \wb_dat_i[11]_pad  ;
	input \wb_dat_i[12]_pad  ;
	input \wb_dat_i[13]_pad  ;
	input \wb_dat_i[14]_pad  ;
	input \wb_dat_i[15]_pad  ;
	input \wb_dat_i[16]_pad  ;
	input \wb_dat_i[17]_pad  ;
	input \wb_dat_i[18]_pad  ;
	input \wb_dat_i[19]_pad  ;
	input \wb_dat_i[1]_pad  ;
	input \wb_dat_i[20]_pad  ;
	input \wb_dat_i[21]_pad  ;
	input \wb_dat_i[22]_pad  ;
	input \wb_dat_i[23]_pad  ;
	input \wb_dat_i[24]_pad  ;
	input \wb_dat_i[25]_pad  ;
	input \wb_dat_i[26]_pad  ;
	input \wb_dat_i[27]_pad  ;
	input \wb_dat_i[28]_pad  ;
	input \wb_dat_i[29]_pad  ;
	input \wb_dat_i[2]_pad  ;
	input \wb_dat_i[30]_pad  ;
	input \wb_dat_i[31]_pad  ;
	input \wb_dat_i[3]_pad  ;
	input \wb_dat_i[4]_pad  ;
	input \wb_dat_i[5]_pad  ;
	input \wb_dat_i[6]_pad  ;
	input \wb_dat_i[7]_pad  ;
	input \wb_dat_i[8]_pad  ;
	input \wb_dat_i[9]_pad  ;
	input wb_err_o_pad ;
	input wb_rst_i_pad ;
	input \wb_sel_i[0]_pad  ;
	input \wb_sel_i[1]_pad  ;
	input \wb_sel_i[2]_pad  ;
	input \wb_sel_i[3]_pad  ;
	input wb_stb_i_pad ;
	input wb_we_i_pad ;
	input \wishbone_BDRead_reg/NET0131  ;
	input \wishbone_BDWrite_reg[0]/NET0131  ;
	input \wishbone_BDWrite_reg[1]/NET0131  ;
	input \wishbone_BDWrite_reg[2]/NET0131  ;
	input \wishbone_BDWrite_reg[3]/NET0131  ;
	input \wishbone_BlockReadTxDataFromMemory_reg/NET0131  ;
	input \wishbone_BlockingIncrementTxPointer_reg/NET0131  ;
	input \wishbone_BlockingTxBDRead_reg/NET0131  ;
	input \wishbone_BlockingTxStatusWrite_reg/NET0131  ;
	input \wishbone_BlockingTxStatusWrite_sync2_reg/NET0131  ;
	input \wishbone_BlockingTxStatusWrite_sync3_reg/NET0131  ;
	input \wishbone_Busy_IRQ_rck_reg/NET0131  ;
	input \wishbone_Busy_IRQ_sync2_reg/P0001  ;
	input \wishbone_Busy_IRQ_sync3_reg/P0001  ;
	input \wishbone_Busy_IRQ_syncb2_reg/P0001  ;
	input \wishbone_Flop_reg/NET0131  ;
	input \wishbone_IncrTxPointer_reg/NET0131  ;
	input \wishbone_LastByteIn_reg/NET0131  ;
	input \wishbone_LastWord_reg/NET0131  ;
	input \wishbone_LatchValidBytes_q_reg/NET0131  ;
	input \wishbone_LatchValidBytes_reg/NET0131  ;
	input \wishbone_LatchedRxLength_reg[0]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[10]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[11]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[12]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[13]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[14]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[15]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[1]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[2]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[3]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[4]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[5]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[6]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[7]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[8]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[9]/NET0131  ;
	input \wishbone_LatchedRxStartFrm_reg/NET0131  ;
	input \wishbone_LatchedTxLength_reg[0]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[10]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[11]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[12]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[13]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[14]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[15]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[1]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[2]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[3]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[4]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[5]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[6]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[7]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[8]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[9]/NET0131  ;
	input \wishbone_MasterWbRX_reg/NET0131  ;
	input \wishbone_MasterWbTX_reg/NET0131  ;
	input \wishbone_ReadTxDataFromFifo_sync2_reg/NET0131  ;
	input \wishbone_ReadTxDataFromFifo_sync3_reg/NET0131  ;
	input \wishbone_ReadTxDataFromFifo_syncb2_reg/NET0131  ;
	input \wishbone_ReadTxDataFromFifo_syncb3_reg/NET0131  ;
	input \wishbone_ReadTxDataFromFifo_tck_reg/NET0131  ;
	input \wishbone_ReadTxDataFromMemory_reg/NET0131  ;
	input \wishbone_RxAbortLatched_reg/NET0131  ;
	input \wishbone_RxAbortSync2_reg/NET0131  ;
	input \wishbone_RxAbortSync3_reg/NET0131  ;
	input \wishbone_RxAbortSync4_reg/NET0131  ;
	input \wishbone_RxAbortSyncb2_reg/NET0131  ;
	input \wishbone_RxBDAddress_reg[1]/NET0131  ;
	input \wishbone_RxBDAddress_reg[2]/NET0131  ;
	input \wishbone_RxBDAddress_reg[3]/NET0131  ;
	input \wishbone_RxBDAddress_reg[4]/NET0131  ;
	input \wishbone_RxBDAddress_reg[5]/NET0131  ;
	input \wishbone_RxBDAddress_reg[6]/NET0131  ;
	input \wishbone_RxBDAddress_reg[7]/NET0131  ;
	input \wishbone_RxBDRead_reg/NET0131  ;
	input \wishbone_RxBDReady_reg/NET0131  ;
	input \wishbone_RxB_IRQ_reg/NET0131  ;
	input \wishbone_RxByteCnt_reg[0]/NET0131  ;
	input \wishbone_RxByteCnt_reg[1]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[10]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[11]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[12]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[13]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[14]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[15]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[16]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[17]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[18]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[19]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[20]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[21]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[22]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[23]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[24]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[25]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[26]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[27]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[28]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[29]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[30]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[31]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[8]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[9]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[0]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[10]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[11]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[12]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[13]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[14]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[15]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[16]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[17]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[18]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[19]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[1]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[20]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[21]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[22]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[23]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[24]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[25]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[26]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[27]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[28]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[29]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[2]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[30]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[31]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[3]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[4]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[5]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[6]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[7]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[8]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[9]/NET0131  ;
	input \wishbone_RxE_IRQ_reg/NET0131  ;
	input \wishbone_RxEn_needed_reg/NET0131  ;
	input \wishbone_RxEn_q_reg/NET0131  ;
	input \wishbone_RxEn_reg/NET0131  ;
	input \wishbone_RxEnableWindow_reg/NET0131  ;
	input \wishbone_RxOverrun_reg/NET0131  ;
	input \wishbone_RxPointerLSB_rst_reg[0]/NET0131  ;
	input \wishbone_RxPointerLSB_rst_reg[1]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[10]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[11]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[12]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[13]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[14]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[15]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[16]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[17]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[18]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[19]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[20]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[21]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[22]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[23]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[24]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[25]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[26]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[27]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[28]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[29]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[2]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[30]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[31]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[3]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[4]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[5]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[6]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[7]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[8]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[9]/NET0131  ;
	input \wishbone_RxPointerRead_reg/NET0131  ;
	input \wishbone_RxReady_reg/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[0]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[1]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[2]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[3]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[4]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[5]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[6]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[7]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[8]/NET0131  ;
	input \wishbone_RxStatusWriteLatched_reg/NET0131  ;
	input \wishbone_RxStatusWriteLatched_sync2_reg/NET0131  ;
	input \wishbone_RxStatusWriteLatched_syncb2_reg/NET0131  ;
	input \wishbone_RxStatus_reg[13]/NET0131  ;
	input \wishbone_RxStatus_reg[14]/NET0131  ;
	input \wishbone_RxValidBytes_reg[0]/NET0131  ;
	input \wishbone_RxValidBytes_reg[1]/NET0131  ;
	input \wishbone_ShiftEndedSync1_reg/NET0131  ;
	input \wishbone_ShiftEndedSync2_reg/NET0131  ;
	input \wishbone_ShiftEndedSync3_reg/NET0131  ;
	input \wishbone_ShiftEndedSync_c1_reg/NET0131  ;
	input \wishbone_ShiftEndedSync_c2_reg/NET0131  ;
	input \wishbone_ShiftEnded_rck_reg/NET0131  ;
	input \wishbone_ShiftEnded_reg/NET0131  ;
	input \wishbone_ShiftWillEnd_reg/NET0131  ;
	input \wishbone_StartOccured_reg/NET0131  ;
	input \wishbone_SyncRxStartFrm_q2_reg/NET0131  ;
	input \wishbone_SyncRxStartFrm_q_reg/NET0131  ;
	input \wishbone_TxAbortPacketBlocked_reg/NET0131  ;
	input \wishbone_TxAbortPacket_NotCleared_reg/NET0131  ;
	input \wishbone_TxAbortPacket_reg/NET0131  ;
	input \wishbone_TxAbort_q_reg/NET0131  ;
	input \wishbone_TxAbort_wb_q_reg/NET0131  ;
	input \wishbone_TxAbort_wb_reg/NET0131  ;
	input \wishbone_TxBDAddress_reg[1]/NET0131  ;
	input \wishbone_TxBDAddress_reg[2]/NET0131  ;
	input \wishbone_TxBDAddress_reg[3]/NET0131  ;
	input \wishbone_TxBDAddress_reg[4]/NET0131  ;
	input \wishbone_TxBDAddress_reg[5]/NET0131  ;
	input \wishbone_TxBDAddress_reg[6]/NET0131  ;
	input \wishbone_TxBDAddress_reg[7]/NET0131  ;
	input \wishbone_TxBDRead_reg/NET0131  ;
	input \wishbone_TxBDReady_reg/NET0131  ;
	input \wishbone_TxB_IRQ_reg/NET0131  ;
	input \wishbone_TxByteCnt_reg[0]/NET0131  ;
	input \wishbone_TxByteCnt_reg[1]/NET0131  ;
	input \wishbone_TxDataLatched_reg[0]/NET0131  ;
	input \wishbone_TxDataLatched_reg[10]/NET0131  ;
	input \wishbone_TxDataLatched_reg[11]/NET0131  ;
	input \wishbone_TxDataLatched_reg[12]/NET0131  ;
	input \wishbone_TxDataLatched_reg[13]/NET0131  ;
	input \wishbone_TxDataLatched_reg[14]/NET0131  ;
	input \wishbone_TxDataLatched_reg[15]/NET0131  ;
	input \wishbone_TxDataLatched_reg[16]/NET0131  ;
	input \wishbone_TxDataLatched_reg[17]/NET0131  ;
	input \wishbone_TxDataLatched_reg[18]/NET0131  ;
	input \wishbone_TxDataLatched_reg[19]/NET0131  ;
	input \wishbone_TxDataLatched_reg[1]/NET0131  ;
	input \wishbone_TxDataLatched_reg[20]/NET0131  ;
	input \wishbone_TxDataLatched_reg[21]/NET0131  ;
	input \wishbone_TxDataLatched_reg[22]/NET0131  ;
	input \wishbone_TxDataLatched_reg[23]/NET0131  ;
	input \wishbone_TxDataLatched_reg[24]/NET0131  ;
	input \wishbone_TxDataLatched_reg[25]/NET0131  ;
	input \wishbone_TxDataLatched_reg[26]/NET0131  ;
	input \wishbone_TxDataLatched_reg[27]/NET0131  ;
	input \wishbone_TxDataLatched_reg[28]/NET0131  ;
	input \wishbone_TxDataLatched_reg[29]/NET0131  ;
	input \wishbone_TxDataLatched_reg[2]/NET0131  ;
	input \wishbone_TxDataLatched_reg[30]/NET0131  ;
	input \wishbone_TxDataLatched_reg[31]/NET0131  ;
	input \wishbone_TxDataLatched_reg[3]/NET0131  ;
	input \wishbone_TxDataLatched_reg[4]/NET0131  ;
	input \wishbone_TxDataLatched_reg[5]/NET0131  ;
	input \wishbone_TxDataLatched_reg[6]/NET0131  ;
	input \wishbone_TxDataLatched_reg[7]/NET0131  ;
	input \wishbone_TxDataLatched_reg[8]/NET0131  ;
	input \wishbone_TxDataLatched_reg[9]/NET0131  ;
	input \wishbone_TxData_reg[0]/NET0131  ;
	input \wishbone_TxData_reg[1]/NET0131  ;
	input \wishbone_TxData_reg[2]/NET0131  ;
	input \wishbone_TxData_reg[3]/NET0131  ;
	input \wishbone_TxData_reg[4]/NET0131  ;
	input \wishbone_TxData_reg[5]/NET0131  ;
	input \wishbone_TxData_reg[6]/NET0131  ;
	input \wishbone_TxData_reg[7]/NET0131  ;
	input \wishbone_TxDonePacketBlocked_reg/NET0131  ;
	input \wishbone_TxDonePacket_NotCleared_reg/NET0131  ;
	input \wishbone_TxDonePacket_reg/NET0131  ;
	input \wishbone_TxDone_wb_q_reg/NET0131  ;
	input \wishbone_TxDone_wb_reg/NET0131  ;
	input \wishbone_TxE_IRQ_reg/NET0131  ;
	input \wishbone_TxEn_needed_reg/NET0131  ;
	input \wishbone_TxEn_q_reg/NET0131  ;
	input \wishbone_TxEn_reg/NET0131  ;
	input \wishbone_TxEndFrm_reg/NET0131  ;
	input \wishbone_TxEndFrm_wb_reg/NET0131  ;
	input \wishbone_TxLength_reg[0]/NET0131  ;
	input \wishbone_TxLength_reg[10]/NET0131  ;
	input \wishbone_TxLength_reg[11]/NET0131  ;
	input \wishbone_TxLength_reg[12]/NET0131  ;
	input \wishbone_TxLength_reg[13]/NET0131  ;
	input \wishbone_TxLength_reg[14]/NET0131  ;
	input \wishbone_TxLength_reg[15]/NET0131  ;
	input \wishbone_TxLength_reg[1]/NET0131  ;
	input \wishbone_TxLength_reg[2]/NET0131  ;
	input \wishbone_TxLength_reg[3]/NET0131  ;
	input \wishbone_TxLength_reg[4]/NET0131  ;
	input \wishbone_TxLength_reg[5]/NET0131  ;
	input \wishbone_TxLength_reg[6]/NET0131  ;
	input \wishbone_TxLength_reg[7]/NET0131  ;
	input \wishbone_TxLength_reg[8]/NET0131  ;
	input \wishbone_TxLength_reg[9]/NET0131  ;
	input \wishbone_TxPointerLSB_reg[0]/NET0131  ;
	input \wishbone_TxPointerLSB_reg[1]/NET0131  ;
	input \wishbone_TxPointerLSB_rst_reg[0]/NET0131  ;
	input \wishbone_TxPointerLSB_rst_reg[1]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[10]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[11]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[12]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[13]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[14]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[15]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[16]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[17]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[18]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[19]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[20]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[21]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[22]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[23]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[24]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[25]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[26]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[27]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[28]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[29]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[2]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[30]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[31]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[3]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[4]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[5]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[6]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[7]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[8]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[9]/NET0131  ;
	input \wishbone_TxPointerRead_reg/NET0131  ;
	input \wishbone_TxRetryPacketBlocked_reg/NET0131  ;
	input \wishbone_TxRetryPacket_NotCleared_reg/NET0131  ;
	input \wishbone_TxRetryPacket_reg/NET0131  ;
	input \wishbone_TxRetry_q_reg/NET0131  ;
	input \wishbone_TxRetry_wb_q_reg/NET0131  ;
	input \wishbone_TxRetry_wb_reg/NET0131  ;
	input \wishbone_TxStartFrm_reg/NET0131  ;
	input \wishbone_TxStartFrm_sync2_reg/NET0131  ;
	input \wishbone_TxStartFrm_syncb2_reg/NET0131  ;
	input \wishbone_TxStartFrm_wb_reg/NET0131  ;
	input \wishbone_TxStatus_reg[11]/NET0131  ;
	input \wishbone_TxStatus_reg[12]/NET0131  ;
	input \wishbone_TxStatus_reg[13]/NET0131  ;
	input \wishbone_TxStatus_reg[14]/NET0131  ;
	input \wishbone_TxUnderRun_reg/NET0131  ;
	input \wishbone_TxUnderRun_sync1_reg/NET0131  ;
	input \wishbone_TxUnderRun_wb_reg/NET0131  ;
	input \wishbone_TxUsedData_q_reg/NET0131  ;
	input \wishbone_TxValidBytesLatched_reg[0]/NET0131  ;
	input \wishbone_TxValidBytesLatched_reg[1]/NET0131  ;
	input \wishbone_WB_ACK_O_reg/P0001  ;
	input \wishbone_WbEn_q_reg/NET0131  ;
	input \wishbone_WbEn_reg/NET0131  ;
	input \wishbone_WriteRxDataToFifoSync2_reg/NET0131  ;
	input \wishbone_WriteRxDataToFifoSync3_reg/NET0131  ;
	input \wishbone_WriteRxDataToFifo_reg/NET0131  ;
	input \wishbone_bd_ram_mem0_reg[0][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[0][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[0][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[0][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[0][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[0][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[0][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[0][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][7]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][9]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][23]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][31]/P0001  ;
	input \wishbone_bd_ram_raddr_reg[0]/P0001  ;
	input \wishbone_bd_ram_raddr_reg[1]/NET0131  ;
	input \wishbone_bd_ram_raddr_reg[2]/NET0131  ;
	input \wishbone_bd_ram_raddr_reg[3]/P0001  ;
	input \wishbone_bd_ram_raddr_reg[4]/NET0131  ;
	input \wishbone_bd_ram_raddr_reg[5]/NET0131  ;
	input \wishbone_bd_ram_raddr_reg[6]/NET0131  ;
	input \wishbone_bd_ram_raddr_reg[7]/NET0131  ;
	input \wishbone_cyc_cleared_reg/NET0131  ;
	input \wishbone_r_RxEn_q_reg/NET0131  ;
	input \wishbone_r_TxEn_q_reg/NET0131  ;
	input \wishbone_ram_addr_reg[0]/NET0131  ;
	input \wishbone_ram_addr_reg[1]/NET0131  ;
	input \wishbone_ram_addr_reg[2]/NET0131  ;
	input \wishbone_ram_addr_reg[3]/NET0131  ;
	input \wishbone_ram_addr_reg[4]/NET0131  ;
	input \wishbone_ram_addr_reg[5]/NET0131  ;
	input \wishbone_ram_addr_reg[6]/NET0131  ;
	input \wishbone_ram_addr_reg[7]/NET0131  ;
	input \wishbone_ram_di_reg[0]/NET0131  ;
	input \wishbone_ram_di_reg[10]/NET0131  ;
	input \wishbone_ram_di_reg[11]/NET0131  ;
	input \wishbone_ram_di_reg[12]/NET0131  ;
	input \wishbone_ram_di_reg[13]/NET0131  ;
	input \wishbone_ram_di_reg[14]/NET0131  ;
	input \wishbone_ram_di_reg[15]/NET0131  ;
	input \wishbone_ram_di_reg[16]/NET0131  ;
	input \wishbone_ram_di_reg[17]/NET0131  ;
	input \wishbone_ram_di_reg[18]/NET0131  ;
	input \wishbone_ram_di_reg[19]/NET0131  ;
	input \wishbone_ram_di_reg[1]/NET0131  ;
	input \wishbone_ram_di_reg[20]/NET0131  ;
	input \wishbone_ram_di_reg[21]/NET0131  ;
	input \wishbone_ram_di_reg[22]/NET0131  ;
	input \wishbone_ram_di_reg[23]/NET0131  ;
	input \wishbone_ram_di_reg[24]/NET0131  ;
	input \wishbone_ram_di_reg[25]/NET0131  ;
	input \wishbone_ram_di_reg[26]/NET0131  ;
	input \wishbone_ram_di_reg[27]/NET0131  ;
	input \wishbone_ram_di_reg[28]/NET0131  ;
	input \wishbone_ram_di_reg[29]/NET0131  ;
	input \wishbone_ram_di_reg[2]/NET0131  ;
	input \wishbone_ram_di_reg[30]/NET0131  ;
	input \wishbone_ram_di_reg[31]/NET0131  ;
	input \wishbone_ram_di_reg[3]/NET0131  ;
	input \wishbone_ram_di_reg[4]/NET0131  ;
	input \wishbone_ram_di_reg[5]/NET0131  ;
	input \wishbone_ram_di_reg[6]/NET0131  ;
	input \wishbone_ram_di_reg[7]/NET0131  ;
	input \wishbone_ram_di_reg[8]/NET0131  ;
	input \wishbone_ram_di_reg[9]/NET0131  ;
	input \wishbone_rx_burst_cnt_reg[0]/NET0131  ;
	input \wishbone_rx_burst_cnt_reg[1]/NET0131  ;
	input \wishbone_rx_burst_cnt_reg[2]/NET0131  ;
	input \wishbone_rx_burst_en_reg/NET0131  ;
	input \wishbone_rx_fifo_cnt_reg[0]/NET0131  ;
	input \wishbone_rx_fifo_cnt_reg[1]/NET0131  ;
	input \wishbone_rx_fifo_cnt_reg[2]/NET0131  ;
	input \wishbone_rx_fifo_cnt_reg[3]/NET0131  ;
	input \wishbone_rx_fifo_cnt_reg[4]/NET0131  ;
	input \wishbone_rx_fifo_fifo_reg[0][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][9]/P0001  ;
	input \wishbone_rx_fifo_read_pointer_reg[0]/NET0131  ;
	input \wishbone_rx_fifo_read_pointer_reg[1]/NET0131  ;
	input \wishbone_rx_fifo_read_pointer_reg[2]/NET0131  ;
	input \wishbone_rx_fifo_read_pointer_reg[3]/NET0131  ;
	input \wishbone_rx_fifo_write_pointer_reg[0]/NET0131  ;
	input \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
	input \wishbone_rx_fifo_write_pointer_reg[2]/NET0131  ;
	input \wishbone_rx_fifo_write_pointer_reg[3]/NET0131  ;
	input \wishbone_tx_burst_cnt_reg[0]/NET0131  ;
	input \wishbone_tx_burst_cnt_reg[1]/NET0131  ;
	input \wishbone_tx_burst_cnt_reg[2]/NET0131  ;
	input \wishbone_tx_burst_en_reg/NET0131  ;
	input \wishbone_tx_fifo_cnt_reg[0]/NET0131  ;
	input \wishbone_tx_fifo_cnt_reg[1]/NET0131  ;
	input \wishbone_tx_fifo_cnt_reg[2]/NET0131  ;
	input \wishbone_tx_fifo_cnt_reg[3]/NET0131  ;
	input \wishbone_tx_fifo_cnt_reg[4]/NET0131  ;
	input \wishbone_tx_fifo_data_out_reg[0]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[10]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[11]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[12]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[13]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[14]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[15]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[16]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[17]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[18]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[19]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[1]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[20]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[21]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[22]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[23]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[24]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[25]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[26]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[27]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[28]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[29]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[2]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[30]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[31]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[3]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[4]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[5]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[6]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[7]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[8]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][9]/P0001  ;
	input \wishbone_tx_fifo_read_pointer_reg[0]/NET0131  ;
	input \wishbone_tx_fifo_read_pointer_reg[1]/NET0131  ;
	input \wishbone_tx_fifo_read_pointer_reg[2]/NET0131  ;
	input \wishbone_tx_fifo_read_pointer_reg[3]/NET0131  ;
	input \wishbone_tx_fifo_write_pointer_reg[0]/NET0131  ;
	input \wishbone_tx_fifo_write_pointer_reg[1]/NET0131  ;
	input \wishbone_tx_fifo_write_pointer_reg[2]/NET0131  ;
	input \wishbone_tx_fifo_write_pointer_reg[3]/NET0131  ;
	output \_al_n1  ;
	output \g215539/_0_  ;
	output \g215543/_0_  ;
	output \g215547/_0_  ;
	output \g215551/_0_  ;
	output \g215552/_0_  ;
	output \g215578/_0_  ;
	output \g215587/_1_  ;
	output \g215589/_1_  ;
	output \g215591/_1_  ;
	output \g215593/_1_  ;
	output \g215595/_1_  ;
	output \g215597/_1_  ;
	output \g215599/_1_  ;
	output \g215601/_1_  ;
	output \g215603/_1_  ;
	output \g215605/_1_  ;
	output \g215607/_1_  ;
	output \g215609/_1_  ;
	output \g215611/_1_  ;
	output \g215613/_1_  ;
	output \g215615/_1_  ;
	output \g215617/_1_  ;
	output \g215618/_0_  ;
	output \g215619/_0_  ;
	output \g215620/_0_  ;
	output \g215632/_1_  ;
	output \g215634/_0_  ;
	output \g215635/_0_  ;
	output \g215636/_0_  ;
	output \g215637/_0_  ;
	output \g215638/_0_  ;
	output \g215639/_0_  ;
	output \g215655/_1_  ;
	output \g215657/_1_  ;
	output \g215659/_1_  ;
	output \g215661/_1_  ;
	output \g215662/_0_  ;
	output \g215663/_0_  ;
	output \g215664/_0_  ;
	output \g215665/_0_  ;
	output \g215668/_0_  ;
	output \g215674/_0_  ;
	output \g215677/_0_  ;
	output \g215686/_0_  ;
	output \g215695/_0_  ;
	output \g215696/_0_  ;
	output \g215702/_1__syn_2  ;
	output \g215705/_0_  ;
	output \g215706/_0_  ;
	output \g215716/_0_  ;
	output \g215717/_0_  ;
	output \g215718/_0_  ;
	output \g215726/_0_  ;
	output \g215727/_0_  ;
	output \g215728/_0_  ;
	output \g215760/_0_  ;
	output \g215764/_0_  ;
	output \g215765/_0_  ;
	output \g215766/_0_  ;
	output \g215767/_3_  ;
	output \g215768/_3_  ;
	output \g215769/_3_  ;
	output \g215770/_3_  ;
	output \g215771/_3_  ;
	output \g215772/_3_  ;
	output \g215773/_3_  ;
	output \g215774/_3_  ;
	output \g215775/_3_  ;
	output \g215776/_3_  ;
	output \g215777/_3_  ;
	output \g215778/_3_  ;
	output \g215779/_3_  ;
	output \g215780/_3_  ;
	output \g215790/_0_  ;
	output \g215791/_0_  ;
	output \g215792/_0_  ;
	output \g215793/_0_  ;
	output \g215801/_0_  ;
	output \g215802/_0_  ;
	output \g215803/_0_  ;
	output \g215804/_0_  ;
	output \g215812/_0_  ;
	output \g215813/_0_  ;
	output \g215821/_0_  ;
	output \g215823/_0_  ;
	output \g215831/_0_  ;
	output \g215832/_0_  ;
	output \g215833/_0_  ;
	output \g215845/_0_  ;
	output \g215846/_0_  ;
	output \g215847/_0_  ;
	output \g215872/_0_  ;
	output \g215873/_0_  ;
	output \g215874/_0_  ;
	output \g215904/_0_  ;
	output \g215905/_0_  ;
	output \g215906/_0_  ;
	output \g215907/_0_  ;
	output \g215908/_0_  ;
	output \g215909/_0_  ;
	output \g215910/_0_  ;
	output \g215911/_0_  ;
	output \g215912/_0_  ;
	output \g215913/_0_  ;
	output \g215914/_0_  ;
	output \g215915/_0_  ;
	output \g215916/_0_  ;
	output \g215917/_0_  ;
	output \g215918/_0_  ;
	output \g215919/_0_  ;
	output \g215920/_0_  ;
	output \g215923/_0_  ;
	output \g215926/_0_  ;
	output \g215941/_0_  ;
	output \g215942/_0_  ;
	output \g215943/_0_  ;
	output \g215944/_0_  ;
	output \g215945/_0_  ;
	output \g215946/_0_  ;
	output \g215947/_0_  ;
	output \g215948/_0_  ;
	output \g215949/_0_  ;
	output \g215950/_0_  ;
	output \g215951/_0_  ;
	output \g215952/_0_  ;
	output \g215953/_0_  ;
	output \g215954/_0_  ;
	output \g215955/_0_  ;
	output \g215956/_0_  ;
	output \g215957/_0_  ;
	output \g215959/_00_  ;
	output \g215960/_0_  ;
	output \g215962/_0_  ;
	output \g215964/_0_  ;
	output \g215966/_0_  ;
	output \g215972/_0_  ;
	output \g216035/_0_  ;
	output \g216037/_0_  ;
	output \g216038/_0_  ;
	output \g216039/_0_  ;
	output \g216040/_0_  ;
	output \g216041/_0_  ;
	output \g216042/_0_  ;
	output \g216046/_0_  ;
	output \g216048/_0_  ;
	output \g216057/_0_  ;
	output \g216263/_0_  ;
	output \g216264/_0_  ;
	output \g216265/_0_  ;
	output \g216266/_0_  ;
	output \g216267/_0_  ;
	output \g216268/_0_  ;
	output \g216269/_0_  ;
	output \g216270/_0_  ;
	output \g216271/_0_  ;
	output \g216272/_0_  ;
	output \g216273/_0_  ;
	output \g216284/_0_  ;
	output \g216289/_0_  ;
	output \g216290/_0_  ;
	output \g216292/_0_  ;
	output \g216296/_0_  ;
	output \g216297/_0_  ;
	output \g216300/_0_  ;
	output \g216301/_0_  ;
	output \g216302/_0_  ;
	output \g216303/_0_  ;
	output \g216304/_0_  ;
	output \g216305/_0_  ;
	output \g216306/_0_  ;
	output \g216307/_0_  ;
	output \g216310/_3_  ;
	output \g216311/_3_  ;
	output \g216314/u3_syn_7  ;
	output \g216322/_3_  ;
	output \g216323/_3_  ;
	output \g216324/_3_  ;
	output \g216325/_3_  ;
	output \g216326/_3_  ;
	output \g216327/_3_  ;
	output \g216328/_3_  ;
	output \g216329/_3_  ;
	output \g216369/_0_  ;
	output \g216370/_0_  ;
	output \g216371/_0_  ;
	output \g216372/_0_  ;
	output \g216373/_0_  ;
	output \g216374/_0_  ;
	output \g216375/_0_  ;
	output \g216376/_0_  ;
	output \g216379/_0_  ;
	output \g216380/_0_  ;
	output \g216381/_0_  ;
	output \g216385/_0_  ;
	output \g216389/_0_  ;
	output \g216390/_0_  ;
	output \g216402/_0_  ;
	output \g216404/_0_  ;
	output \g216405/_0_  ;
	output \g216406/_0_  ;
	output \g216407/_0_  ;
	output \g216408/_0_  ;
	output \g216409/_0_  ;
	output \g216410/_0_  ;
	output \g216411/_0_  ;
	output \g216412/_0_  ;
	output \g216413/_0_  ;
	output \g216414/_0_  ;
	output \g216415/_0_  ;
	output \g216416/_0_  ;
	output \g216417/_0_  ;
	output \g216418/_0_  ;
	output \g216419/_0_  ;
	output \g216420/_0_  ;
	output \g216421/_0_  ;
	output \g216422/_0_  ;
	output \g216423/_0_  ;
	output \g216424/_0_  ;
	output \g216425/_0_  ;
	output \g216426/_0_  ;
	output \g216427/_0_  ;
	output \g216428/_0_  ;
	output \g216429/_0_  ;
	output \g216430/_0_  ;
	output \g216431/_0_  ;
	output \g216432/_0_  ;
	output \g216433/_0_  ;
	output \g216434/_0_  ;
	output \g216435/_0_  ;
	output \g216436/_0_  ;
	output \g216437/_0_  ;
	output \g216438/_0_  ;
	output \g216439/_3_  ;
	output \g216447/_3_  ;
	output \g216448/_3_  ;
	output \g216452/_0_  ;
	output \g216453/_0_  ;
	output \g216454/_0_  ;
	output \g216455/_0_  ;
	output \g216456/_0_  ;
	output \g216457/_0_  ;
	output \g216458/_3_  ;
	output \g216459/_3_  ;
	output \g216461/_3_  ;
	output \g216462/_3_  ;
	output \g216463/_3_  ;
	output \g216464/_3_  ;
	output \g216465/_3_  ;
	output \g216466/_0_  ;
	output \g216467/_3_  ;
	output \g216468/_3_  ;
	output \g216469/_3_  ;
	output \g216470/_3_  ;
	output \g216471/_3_  ;
	output \g216473/_3_  ;
	output \g216474/_3_  ;
	output \g216475/_3_  ;
	output \g216476/_3_  ;
	output \g216477/_3_  ;
	output \g216478/_0_  ;
	output \g216479/_3_  ;
	output \g216480/_3_  ;
	output \g216481/_3_  ;
	output \g216492/_0_  ;
	output \g216494/_0_  ;
	output \g216495/_3_  ;
	output \g216496/_3_  ;
	output \g216498/_3_  ;
	output \g216499/_3_  ;
	output \g216500/_3_  ;
	output \g216513/_3_  ;
	output \g216514/_3_  ;
	output \g216515/_3_  ;
	output \g216516/_3_  ;
	output \g216517/_3_  ;
	output \g216518/_3_  ;
	output \g216519/_3_  ;
	output \g216520/_3_  ;
	output \g216521/_3_  ;
	output \g216522/_3_  ;
	output \g216523/_3_  ;
	output \g216524/_3_  ;
	output \g216525/_3_  ;
	output \g216526/_3_  ;
	output \g216527/_3_  ;
	output \g216528/_3_  ;
	output \g216529/_3_  ;
	output \g216530/_3_  ;
	output \g216531/_3_  ;
	output \g216532/_3_  ;
	output \g216533/_3_  ;
	output \g216534/_3_  ;
	output \g216535/_3_  ;
	output \g216536/_3_  ;
	output \g216537/_3_  ;
	output \g216538/_3_  ;
	output \g216555/_3_  ;
	output \g216556/_3_  ;
	output \g216557/_3_  ;
	output \g216560/_3_  ;
	output \g216561/_3_  ;
	output \g216562/_3_  ;
	output \g216563/_3_  ;
	output \g216564/_3_  ;
	output \g216565/_3_  ;
	output \g216566/_3_  ;
	output \g216567/_3_  ;
	output \g216568/_3_  ;
	output \g216569/_3_  ;
	output \g216570/_3_  ;
	output \g216571/_3_  ;
	output \g216575/_3_  ;
	output \g216576/_3_  ;
	output \g216577/_3_  ;
	output \g216578/_3_  ;
	output \g216579/_3_  ;
	output \g216580/_3_  ;
	output \g216581/_3_  ;
	output \g216582/_3_  ;
	output \g216583/_3_  ;
	output \g216586/_3_  ;
	output \g216587/_3_  ;
	output \g216588/_3_  ;
	output \g216589/_3_  ;
	output \g216590/_3_  ;
	output \g216591/_3_  ;
	output \g216592/_3_  ;
	output \g216593/_3_  ;
	output \g216594/_3_  ;
	output \g216595/_3_  ;
	output \g216600/_3_  ;
	output \g216683/_0_  ;
	output \g216689/_0_  ;
	output \g216693/_0_  ;
	output \g216694/_0_  ;
	output \g216727/_0_  ;
	output \g216728/_0_  ;
	output \g216729/_0_  ;
	output \g216732/_0_  ;
	output \g216733/_0_  ;
	output \g216734/_0_  ;
	output \g216735/_0_  ;
	output \g216736/_0_  ;
	output \g216737/_0_  ;
	output \g216738/_0_  ;
	output \g216739/_0_  ;
	output \g216740/_0_  ;
	output \g216741/_0_  ;
	output \g216742/_0_  ;
	output \g216743/_0_  ;
	output \g216744/_0_  ;
	output \g216745/_0_  ;
	output \g216746/_0_  ;
	output \g216748/_0_  ;
	output \g216751/_0_  ;
	output \g216754/_0_  ;
	output \g216762/_0_  ;
	output \g216934/_2_  ;
	output \g216952/_0_  ;
	output \g216955/_0_  ;
	output \g216969/_0_  ;
	output \g216979/_0_  ;
	output \g216984/_0_  ;
	output \g216996/_0_  ;
	output \g217002/_0_  ;
	output \g217014/_0_  ;
	output \g217015/_0_  ;
	output \g217016/_0_  ;
	output \g217017/_0_  ;
	output \g217018/_0_  ;
	output \g217019/_0_  ;
	output \g217023/_0_  ;
	output \g217116/_0_  ;
	output \g217146/_3_  ;
	output \g217149/_0_  ;
	output \g217151/_0_  ;
	output \g217160/_0_  ;
	output \g217167/_0_  ;
	output \g217168/_0_  ;
	output \g217169/_0_  ;
	output \g217170/_0_  ;
	output \g217171/_0_  ;
	output \g217172/_0_  ;
	output \g217173/_0_  ;
	output \g217174/_0_  ;
	output \g217175/_0_  ;
	output \g217176/_0_  ;
	output \g217177/_0_  ;
	output \g217178/_0_  ;
	output \g217179/_0_  ;
	output \g217180/_0_  ;
	output \g217181/_0_  ;
	output \g217182/_0_  ;
	output \g217183/_0_  ;
	output \g217187/_0_  ;
	output \g217188/_0_  ;
	output \g217189/_0_  ;
	output \g217193/_0_  ;
	output \g217194/_0_  ;
	output \g217195/_0_  ;
	output \g217196/_0_  ;
	output \g217202/_0_  ;
	output \g217205/_0_  ;
	output \g217206/_0_  ;
	output \g217207/_0_  ;
	output \g217208/_0_  ;
	output \g217209/_0_  ;
	output \g217210/_0_  ;
	output \g217211/_0_  ;
	output \g217212/_0_  ;
	output \g217213/_0_  ;
	output \g217214/_0_  ;
	output \g217215/_0_  ;
	output \g217216/_0_  ;
	output \g217217/_0_  ;
	output \g217218/_0_  ;
	output \g217219/_0_  ;
	output \g217220/_0_  ;
	output \g217223/_0_  ;
	output \g217231/_0_  ;
	output \g217237/_0_  ;
	output \g217238/_0_  ;
	output \g217242/_0_  ;
	output \g217243/_0_  ;
	output \g217250/_3_  ;
	output \g217251/_3_  ;
	output \g217252/_3_  ;
	output \g217253/_3_  ;
	output \g217254/_3_  ;
	output \g217255/_3_  ;
	output \g217256/_3_  ;
	output \g217257/_3_  ;
	output \g217258/_3_  ;
	output \g217259/_3_  ;
	output \g217260/_3_  ;
	output \g217261/_3_  ;
	output \g217262/_3_  ;
	output \g217263/_3_  ;
	output \g217264/_3_  ;
	output \g217265/_3_  ;
	output \g217266/_3_  ;
	output \g217267/_3_  ;
	output \g217268/_3_  ;
	output \g217269/_3_  ;
	output \g217270/_3_  ;
	output \g217271/_3_  ;
	output \g217272/_3_  ;
	output \g217273/_3_  ;
	output \g217274/_3_  ;
	output \g217275/_3_  ;
	output \g217276/_3_  ;
	output \g217277/_3_  ;
	output \g217278/_3_  ;
	output \g217279/_3_  ;
	output \g217280/_3_  ;
	output \g217281/_3_  ;
	output \g217282/_3_  ;
	output \g217283/_3_  ;
	output \g217284/_3_  ;
	output \g217285/_3_  ;
	output \g217286/_3_  ;
	output \g217287/_3_  ;
	output \g217288/_3_  ;
	output \g217289/_3_  ;
	output \g217290/_3_  ;
	output \g217291/_3_  ;
	output \g217292/_3_  ;
	output \g217293/_3_  ;
	output \g217294/_3_  ;
	output \g217295/_3_  ;
	output \g217296/_3_  ;
	output \g217297/_3_  ;
	output \g217298/_3_  ;
	output \g217299/_3_  ;
	output \g217300/_3_  ;
	output \g217301/_3_  ;
	output \g217302/_3_  ;
	output \g217303/_3_  ;
	output \g217304/_3_  ;
	output \g217305/_3_  ;
	output \g217306/_3_  ;
	output \g217307/_3_  ;
	output \g217308/_3_  ;
	output \g217309/_3_  ;
	output \g217310/_3_  ;
	output \g217311/_3_  ;
	output \g217312/_3_  ;
	output \g217313/_3_  ;
	output \g217318/_0_  ;
	output \g217662/_0_  ;
	output \g217663/_0_  ;
	output \g217682/_0_  ;
	output \g217697/_0_  ;
	output \g217698/_0_  ;
	output \g217699/_0_  ;
	output \g217700/_0_  ;
	output \g217701/_0_  ;
	output \g217705/_0_  ;
	output \g217711/_0_  ;
	output \g217747/_0_  ;
	output \g217753/_00_  ;
	output \g217775/_0_  ;
	output \g217781/_0_  ;
	output \g217784/_0_  ;
	output \g217785/_0_  ;
	output \g217786/_0_  ;
	output \g217787/_0_  ;
	output \g217788/_0_  ;
	output \g217790/_0_  ;
	output \g217815/_0_  ;
	output \g217817/_0_  ;
	output \g218145/_0_  ;
	output \g218148/_0_  ;
	output \g218150/_0_  ;
	output \g218167/_0_  ;
	output \g218168/_0_  ;
	output \g218234/_0_  ;
	output \g218235/_0_  ;
	output \g218236/_0_  ;
	output \g218238/_0_  ;
	output \g218242/_0_  ;
	output \g218332/_0_  ;
	output \g218335/_0_  ;
	output \g218336/_0_  ;
	output \g218337/_0_  ;
	output \g218338/_0_  ;
	output \g218339/_0_  ;
	output \g218340/_0_  ;
	output \g218341/_0_  ;
	output \g218342/_0_  ;
	output \g218343/_0_  ;
	output \g218344/_0_  ;
	output \g218345/_0_  ;
	output \g218346/_0_  ;
	output \g218347/_0_  ;
	output \g218348/_0_  ;
	output \g218349/_0_  ;
	output \g218350/_0_  ;
	output \g218351/_0_  ;
	output \g218352/_0_  ;
	output \g218353/_0_  ;
	output \g218354/_0_  ;
	output \g218355/_0_  ;
	output \g218356/_0_  ;
	output \g218357/_0_  ;
	output \g218358/_0_  ;
	output \g218359/_0_  ;
	output \g218360/_0_  ;
	output \g218398/_3_  ;
	output \g218430/_0_  ;
	output \g218440/_0_  ;
	output \g218452/u3_syn_4  ;
	output \g218495/u3_syn_4  ;
	output \g218517/u3_syn_4  ;
	output \g218554/u3_syn_4  ;
	output \g218575/u3_syn_4  ;
	output \g218600/u3_syn_4  ;
	output \g218621/u3_syn_4  ;
	output \g218638/u3_syn_4  ;
	output \g218659/u3_syn_4  ;
	output \g218673/u3_syn_4  ;
	output \g218707/u3_syn_4  ;
	output \g218735/_3_  ;
	output \g219186/_0_  ;
	output \g219187/_0_  ;
	output \g219188/_0_  ;
	output \g219189/_0_  ;
	output \g219190/_0_  ;
	output \g219196/_0_  ;
	output \g219198/_0_  ;
	output \g219199/_0_  ;
	output \g219200/_0_  ;
	output \g219308/_0_  ;
	output \g219314/_0_  ;
	output \g219326/_0_  ;
	output \g219328/_0_  ;
	output \g219348/_0_  ;
	output \g219351/_0_  ;
	output \g219363/_0_  ;
	output \g219364/_0_  ;
	output \g219365/_0_  ;
	output \g219366/_0_  ;
	output \g219367/_0_  ;
	output \g219368/_0_  ;
	output \g219369/_0_  ;
	output \g219376/_0_  ;
	output \g219381/_0_  ;
	output \g219382/_0_  ;
	output \g219384/_0_  ;
	output \g219385/_0_  ;
	output \g219391/_0_  ;
	output \g219394/_0_  ;
	output \g219395/_0_  ;
	output \g219396/_0_  ;
	output \g219397/_0_  ;
	output \g219398/_0_  ;
	output \g219399/_0_  ;
	output \g219400/_0_  ;
	output \g219401/_0_  ;
	output \g219402/_0_  ;
	output \g219403/_0_  ;
	output \g219404/_0_  ;
	output \g219405/_0_  ;
	output \g219406/_0_  ;
	output \g219407/_0_  ;
	output \g219408/_0_  ;
	output \g219409/_0_  ;
	output \g219410/_0_  ;
	output \g219411/_0_  ;
	output \g219412/_0_  ;
	output \g219413/_0_  ;
	output \g219414/_0_  ;
	output \g219415/_0_  ;
	output \g219416/_0_  ;
	output \g219417/_0_  ;
	output \g219418/_0_  ;
	output \g219419/_0_  ;
	output \g219420/_0_  ;
	output \g219421/_0_  ;
	output \g219422/_0_  ;
	output \g219423/_0_  ;
	output \g219424/_0_  ;
	output \g219425/_0_  ;
	output \g219426/_0_  ;
	output \g219427/_0_  ;
	output \g219428/_0_  ;
	output \g219429/_0_  ;
	output \g219430/_0_  ;
	output \g219431/_0_  ;
	output \g219432/_0_  ;
	output \g219433/_0_  ;
	output \g219434/_0_  ;
	output \g219435/_0_  ;
	output \g219436/_0_  ;
	output \g219437/_0_  ;
	output \g219438/_0_  ;
	output \g219439/_0_  ;
	output \g219440/_0_  ;
	output \g219441/_0_  ;
	output \g219442/_0_  ;
	output \g219443/_0_  ;
	output \g219444/_0_  ;
	output \g219445/_0_  ;
	output \g219446/_0_  ;
	output \g219447/_0_  ;
	output \g219449/_0_  ;
	output \g219450/_0_  ;
	output \g219451/_0_  ;
	output \g219452/_0_  ;
	output \g219453/_0_  ;
	output \g219454/_0_  ;
	output \g219455/_0_  ;
	output \g219456/_0_  ;
	output \g219457/_0_  ;
	output \g219458/_0_  ;
	output \g219464/u3_syn_7  ;
	output \g219496/u3_syn_4  ;
	output \g219512/u3_syn_4  ;
	output \g219526/u3_syn_4  ;
	output \g219549/u3_syn_4  ;
	output \g219571/u3_syn_4  ;
	output \g219588/u3_syn_4  ;
	output \g219603/u3_syn_4  ;
	output \g219621/u3_syn_4  ;
	output \g219636/_3_  ;
	output \g219652/u3_syn_4  ;
	output \g219676/_3_  ;
	output \g219686/_0_  ;
	output \g219689/_0_  ;
	output \g219694/_3_  ;
	output \g220062/_0_  ;
	output \g220068/_0_  ;
	output \g220069/_0_  ;
	output \g220072/_0_  ;
	output \g220084/_0_  ;
	output \g220149/_0_  ;
	output \g220162/_0_  ;
	output \g220317/_0_  ;
	output \g220360/_2_  ;
	output \g220368/_2_  ;
	output \g220369/_0_  ;
	output \g220370/_0_  ;
	output \g220371/_0_  ;
	output \g220372/_0_  ;
	output \g220376/_0_  ;
	output \g220390/_0_  ;
	output \g220395/_0_  ;
	output \g220499/_0_  ;
	output \g220500/_0_  ;
	output \g220501/_0_  ;
	output \g220502/_0_  ;
	output \g220503/_0_  ;
	output \g220504/_0_  ;
	output \g220505/_0_  ;
	output \g220506/_0_  ;
	output \g220507/_0_  ;
	output \g220508/_0_  ;
	output \g220509/_0_  ;
	output \g220510/_0_  ;
	output \g220511/_0_  ;
	output \g220512/_0_  ;
	output \g220513/_0_  ;
	output \g220514/_0_  ;
	output \g220515/_0_  ;
	output \g220516/_0_  ;
	output \g220517/_0_  ;
	output \g220518/_0_  ;
	output \g220519/_0_  ;
	output \g220520/_0_  ;
	output \g220521/_0_  ;
	output \g220522/_0_  ;
	output \g220523/_0_  ;
	output \g220524/_0_  ;
	output \g220525/_0_  ;
	output \g220526/_0_  ;
	output \g220527/_0_  ;
	output \g220528/_0_  ;
	output \g220529/_0_  ;
	output \g220530/_0_  ;
	output \g220531/_0_  ;
	output \g220532/_0_  ;
	output \g220533/_0_  ;
	output \g220534/_0_  ;
	output \g220535/_0_  ;
	output \g220557/_0_  ;
	output \g220558/_0_  ;
	output \g220559/_0_  ;
	output \g220560/_0_  ;
	output \g220561/_0_  ;
	output \g220562/_0_  ;
	output \g220563/_0_  ;
	output \g220564/_0_  ;
	output \g220565/_0_  ;
	output \g220566/_0_  ;
	output \g220567/_0_  ;
	output \g220568/_0_  ;
	output \g220569/_0_  ;
	output \g220570/_0_  ;
	output \g220571/_0_  ;
	output \g220572/_0_  ;
	output \g220573/_0_  ;
	output \g220574/_0_  ;
	output \g220575/_0_  ;
	output \g220576/_0_  ;
	output \g220577/_0_  ;
	output \g220578/_0_  ;
	output \g220579/_0_  ;
	output \g220580/_0_  ;
	output \g220581/_0_  ;
	output \g220582/_0_  ;
	output \g220583/_0_  ;
	output \g220584/_0_  ;
	output \g220585/_0_  ;
	output \g220586/_0_  ;
	output \g220587/_0_  ;
	output \g220588/_0_  ;
	output \g220589/_0_  ;
	output \g220590/_0_  ;
	output \g220591/_0_  ;
	output \g220592/_0_  ;
	output \g220593/_0_  ;
	output \g220594/_0_  ;
	output \g220595/_0_  ;
	output \g220596/_0_  ;
	output \g220597/_0_  ;
	output \g220598/_0_  ;
	output \g220599/_0_  ;
	output \g220600/_0_  ;
	output \g220601/_0_  ;
	output \g220602/_0_  ;
	output \g220603/_0_  ;
	output \g220604/_0_  ;
	output \g220605/_0_  ;
	output \g220606/_0_  ;
	output \g220607/_0_  ;
	output \g220608/_0_  ;
	output \g220609/_0_  ;
	output \g220610/_0_  ;
	output \g220611/_0_  ;
	output \g220612/_0_  ;
	output \g220613/_0_  ;
	output \g220614/_0_  ;
	output \g220615/_0_  ;
	output \g220616/_0_  ;
	output \g220617/_0_  ;
	output \g220618/_0_  ;
	output \g220619/_0_  ;
	output \g220620/_0_  ;
	output \g220621/_0_  ;
	output \g220622/_0_  ;
	output \g220623/_0_  ;
	output \g220624/_0_  ;
	output \g220625/_0_  ;
	output \g220626/_0_  ;
	output \g220627/_0_  ;
	output \g220628/_0_  ;
	output \g220629/_0_  ;
	output \g220630/_0_  ;
	output \g220631/_0_  ;
	output \g220632/_0_  ;
	output \g220633/_0_  ;
	output \g220634/_0_  ;
	output \g220635/_0_  ;
	output \g220636/_0_  ;
	output \g220637/_0_  ;
	output \g220638/_0_  ;
	output \g220639/_0_  ;
	output \g220640/_0_  ;
	output \g220641/_0_  ;
	output \g220642/_0_  ;
	output \g220643/_0_  ;
	output \g220644/_0_  ;
	output \g220645/_0_  ;
	output \g220646/_0_  ;
	output \g220647/_0_  ;
	output \g220648/_0_  ;
	output \g220649/_0_  ;
	output \g220650/_0_  ;
	output \g220651/_0_  ;
	output \g220652/_0_  ;
	output \g220653/_0_  ;
	output \g220654/_0_  ;
	output \g220655/_0_  ;
	output \g220656/_0_  ;
	output \g220657/_0_  ;
	output \g220658/_0_  ;
	output \g220659/_0_  ;
	output \g220660/_0_  ;
	output \g220661/_0_  ;
	output \g220662/_0_  ;
	output \g220663/_0_  ;
	output \g220664/_0_  ;
	output \g220665/_0_  ;
	output \g220666/_0_  ;
	output \g220674/_0_  ;
	output \g220679/u3_syn_7  ;
	output \g220711/u3_syn_4  ;
	output \g220726/u3_syn_4  ;
	output \g220739/u3_syn_4  ;
	output \g220751/u3_syn_4  ;
	output \g220759/u3_syn_4  ;
	output \g220773/u3_syn_4  ;
	output \g220782/u3_syn_4  ;
	output \g220805/u3_syn_4  ;
	output \g220828/u3_syn_4  ;
	output \g220921/_0_  ;
	output \g220930/u3_syn_4  ;
	output \g220949/_3_  ;
	output \g220994/_3_  ;
	output \g221207/_0_  ;
	output \g221213/_0_  ;
	output \g221223/_0_  ;
	output \g221224/_0_  ;
	output \g221225/_0_  ;
	output \g221226/_0_  ;
	output \g221231/_0_  ;
	output \g221232/_0_  ;
	output \g221234/_0_  ;
	output \g221235/_0_  ;
	output \g221246/_2_  ;
	output \g221249/_2_  ;
	output \g221265/_0_  ;
	output \g221287/_0_  ;
	output \g221325/_0_  ;
	output \g221326/_0_  ;
	output \g221447/_0_  ;
	output \g221449/_0_  ;
	output \g221452/_0_  ;
	output \g221469/_0_  ;
	output \g221473/_0_  ;
	output \g221503/_0_  ;
	output \g221510/_0_  ;
	output \g221512/_0_  ;
	output \g221516/_0_  ;
	output \g221517/_0_  ;
	output \g221524/_0_  ;
	output \g221530/_0_  ;
	output \g221592/_0_  ;
	output \g221593/_0_  ;
	output \g221634/u3_syn_4  ;
	output \g221669/u3_syn_4  ;
	output \g221789/u3_syn_4  ;
	output \g221813/u3_syn_4  ;
	output \g221829/u3_syn_4  ;
	output \g221861/u3_syn_4  ;
	output \g221876/_0_  ;
	output \g221935/_0_  ;
	output \g221944/_3_  ;
	output \g230200/_0_  ;
	output \g230201/_0_  ;
	output \g230205/_0_  ;
	output \g230295/_0_  ;
	output \g230297/_0_  ;
	output \g230298/_0_  ;
	output \g230300/_0_  ;
	output \g230302/_0_  ;
	output \g230303/_0_  ;
	output \g230343/_0_  ;
	output \g230368/_0_  ;
	output \g230511/_0_  ;
	output \g230531/_0_  ;
	output \g230635/_2_  ;
	output \g230661/_0_  ;
	output \g230715/_1__syn_2  ;
	output \g230731/_0_  ;
	output \g230766/_0_  ;
	output \g230784/_0_  ;
	output \g230785/_0_  ;
	output \g230786/_0_  ;
	output \g230787/_0_  ;
	output \g230797/_0_  ;
	output \g230798/_0_  ;
	output \g230803/_0_  ;
	output \g230804/_00_  ;
	output \g230805/_00_  ;
	output \g230806/_00_  ;
	output \g230807/_00_  ;
	output \g230808/_00_  ;
	output \g230809/_00_  ;
	output \g230815/_0_  ;
	output \g230816/_2_  ;
	output \g230817/_2_  ;
	output \g230829/_0_  ;
	output \g230834/_0_  ;
	output \g230835/_0_  ;
	output \g230836/_0_  ;
	output \g230837/_0_  ;
	output \g230844/_0_  ;
	output \g230863/_3_  ;
	output \g230864/_3_  ;
	output \g230870/_0_  ;
	output \g230988/_3_  ;
	output \g231010/_3_  ;
	output \g231016/_3_  ;
	output \g231042/_3_  ;
	output \g231471/_0_  ;
	output \g231472/_0_  ;
	output \g231476/_3_  ;
	output \g231480/_3_  ;
	output \g231484/_3_  ;
	output \g231504/_0_  ;
	output \g231532/_0_  ;
	output \g231542/_0_  ;
	output \g231560/_1_  ;
	output \g231578/_1_  ;
	output \g231580/_0_  ;
	output \g231590/_1__syn_2  ;
	output \g231615/_0_  ;
	output \g231623/_1_  ;
	output \g231634/_2_  ;
	output \g231635/_0_  ;
	output \g231638/_2_  ;
	output \g231640/_0_  ;
	output \g231653/_2_  ;
	output \g231787/_0_  ;
	output \g231931/_0_  ;
	output \g231939/_3_  ;
	output \g231940/_0_  ;
	output \g231951/_0_  ;
	output \g231955/_0_  ;
	output \g231956/_0_  ;
	output \g231959/_2_  ;
	output \g231960/_0_  ;
	output \g231964/_0_  ;
	output \g231965/_0_  ;
	output \g231975/_0_  ;
	output \g231986/_1_  ;
	output \g231987/_1_  ;
	output \g231989/_1_  ;
	output \g231990/_1_  ;
	output \g231991/_0_  ;
	output \g231992/_0_  ;
	output \g231995/_0_  ;
	output \g231998/_0_  ;
	output \g231999/_0_  ;
	output \g232002/_3_  ;
	output \g232035/u3_syn_4  ;
	output \g232038/u3_syn_4  ;
	output \g232046/u3_syn_4  ;
	output \g232054/u3_syn_4  ;
	output \g232062/u3_syn_4  ;
	output \g232070/u3_syn_4  ;
	output \g232078/u3_syn_4  ;
	output \g232079/u3_syn_4  ;
	output \g232087/u3_syn_4  ;
	output \g232096/u3_syn_4  ;
	output \g232104/u3_syn_4  ;
	output \g232112/u3_syn_4  ;
	output \g232120/u3_syn_4  ;
	output \g232128/u3_syn_4  ;
	output \g232136/u3_syn_4  ;
	output \g232144/u3_syn_4  ;
	output \g232152/u3_syn_4  ;
	output \g232161/u3_syn_4  ;
	output \g232169/u3_syn_4  ;
	output \g232177/u3_syn_4  ;
	output \g232185/u3_syn_4  ;
	output \g232186/u3_syn_4  ;
	output \g232194/u3_syn_4  ;
	output \g232202/u3_syn_4  ;
	output \g232210/u3_syn_4  ;
	output \g232218/u3_syn_4  ;
	output \g232226/u3_syn_4  ;
	output \g232234/u3_syn_4  ;
	output \g232242/u3_syn_4  ;
	output \g232251/u3_syn_4  ;
	output \g232259/u3_syn_4  ;
	output \g232267/u3_syn_4  ;
	output \g232275/u3_syn_4  ;
	output \g232283/u3_syn_4  ;
	output \g232291/u3_syn_4  ;
	output \g232299/u3_syn_4  ;
	output \g232307/u3_syn_4  ;
	output \g232315/u3_syn_4  ;
	output \g232324/u3_syn_4  ;
	output \g232332/u3_syn_4  ;
	output \g232341/u3_syn_4  ;
	output \g232349/u3_syn_4  ;
	output \g232357/u3_syn_4  ;
	output \g232366/u3_syn_4  ;
	output \g232374/u3_syn_4  ;
	output \g232382/u3_syn_4  ;
	output \g232390/u3_syn_4  ;
	output \g232398/u3_syn_4  ;
	output \g232406/u3_syn_4  ;
	output \g232414/u3_syn_4  ;
	output \g232422/u3_syn_4  ;
	output \g232427/u3_syn_4  ;
	output \g232431/u3_syn_4  ;
	output \g232439/u3_syn_4  ;
	output \g232444/u3_syn_4  ;
	output \g232452/u3_syn_4  ;
	output \g232461/u3_syn_4  ;
	output \g232471/u3_syn_4  ;
	output \g232479/u3_syn_4  ;
	output \g232487/u3_syn_4  ;
	output \g232495/u3_syn_4  ;
	output \g232503/u3_syn_4  ;
	output \g232506/u3_syn_4  ;
	output \g232514/u3_syn_4  ;
	output \g232527/u3_syn_4  ;
	output \g232530/u3_syn_4  ;
	output \g232536/u3_syn_4  ;
	output \g232544/u3_syn_4  ;
	output \g232551/u3_syn_4  ;
	output \g232557/u3_syn_4  ;
	output \g232568/u3_syn_4  ;
	output \g232576/u3_syn_4  ;
	output \g232585/u3_syn_4  ;
	output \g232593/u3_syn_4  ;
	output \g232597/u3_syn_4  ;
	output \g232609/u3_syn_4  ;
	output \g232617/u3_syn_4  ;
	output \g232625/u3_syn_4  ;
	output \g232633/u3_syn_4  ;
	output \g232641/u3_syn_4  ;
	output \g232649/u3_syn_4  ;
	output \g232657/u3_syn_4  ;
	output \g232665/u3_syn_4  ;
	output \g232673/u3_syn_4  ;
	output \g232681/u3_syn_4  ;
	output \g232689/u3_syn_4  ;
	output \g232697/u3_syn_4  ;
	output \g232705/u3_syn_4  ;
	output \g232713/u3_syn_4  ;
	output \g232717/u3_syn_4  ;
	output \g232729/u3_syn_4  ;
	output \g232737/u3_syn_4  ;
	output \g232745/u3_syn_4  ;
	output \g232749/u3_syn_4  ;
	output \g232761/u3_syn_4  ;
	output \g232768/u3_syn_4  ;
	output \g232777/u3_syn_4  ;
	output \g232785/u3_syn_4  ;
	output \g232793/u3_syn_4  ;
	output \g232801/u3_syn_4  ;
	output \g232809/u3_syn_4  ;
	output \g232815/u3_syn_4  ;
	output \g232823/u3_syn_4  ;
	output \g232833/u3_syn_4  ;
	output \g232841/u3_syn_4  ;
	output \g232846/u3_syn_4  ;
	output \g232851/u3_syn_4  ;
	output \g232865/u3_syn_4  ;
	output \g232873/u3_syn_4  ;
	output \g232881/u3_syn_4  ;
	output \g232882/u3_syn_4  ;
	output \g232895/u3_syn_4  ;
	output \g232904/u3_syn_4  ;
	output \g232913/u3_syn_4  ;
	output \g232921/u3_syn_4  ;
	output \g232928/u3_syn_4  ;
	output \g232934/u3_syn_4  ;
	output \g232945/u3_syn_4  ;
	output \g232953/u3_syn_4  ;
	output \g232954/u3_syn_4  ;
	output \g232969/u3_syn_4  ;
	output \g232977/u3_syn_4  ;
	output \g232981/u3_syn_4  ;
	output \g232993/u3_syn_4  ;
	output \g232995/u3_syn_4  ;
	output \g233009/u3_syn_4  ;
	output \g233017/u3_syn_4  ;
	output \g233025/u3_syn_4  ;
	output \g233033/u3_syn_4  ;
	output \g233041/u3_syn_4  ;
	output \g233047/u3_syn_4  ;
	output \g233057/u3_syn_4  ;
	output \g233065/u3_syn_4  ;
	output \g233073/u3_syn_4  ;
	output \g233081/u3_syn_4  ;
	output \g233087/u3_syn_4  ;
	output \g233097/u3_syn_4  ;
	output \g233105/u3_syn_4  ;
	output \g233113/u3_syn_4  ;
	output \g233121/u3_syn_4  ;
	output \g233128/u3_syn_4  ;
	output \g233134/u3_syn_4  ;
	output \g233144/u3_syn_4  ;
	output \g233153/u3_syn_4  ;
	output \g233161/u3_syn_4  ;
	output \g233169/u3_syn_4  ;
	output \g233177/u3_syn_4  ;
	output \g233185/u3_syn_4  ;
	output \g233193/u3_syn_4  ;
	output \g233201/u3_syn_4  ;
	output \g233209/u3_syn_4  ;
	output \g233217/u3_syn_4  ;
	output \g233219/u3_syn_4  ;
	output \g233229/u3_syn_4  ;
	output \g233241/u3_syn_4  ;
	output \g233249/u3_syn_4  ;
	output \g233257/u3_syn_4  ;
	output \g233265/u3_syn_4  ;
	output \g233273/u3_syn_4  ;
	output \g233281/u3_syn_4  ;
	output \g233289/u3_syn_4  ;
	output \g233297/u3_syn_4  ;
	output \g233305/u3_syn_4  ;
	output \g233313/u3_syn_4  ;
	output \g233321/u3_syn_4  ;
	output \g233329/u3_syn_4  ;
	output \g233337/u3_syn_4  ;
	output \g233345/u3_syn_4  ;
	output \g233353/u3_syn_4  ;
	output \g233361/u3_syn_4  ;
	output \g233369/u3_syn_4  ;
	output \g233377/u3_syn_4  ;
	output \g233382/u3_syn_4  ;
	output \g233392/u3_syn_4  ;
	output \g233394/u3_syn_4  ;
	output \g233409/u3_syn_4  ;
	output \g233417/u3_syn_4  ;
	output \g233425/u3_syn_4  ;
	output \g233433/u3_syn_4  ;
	output \g233441/u3_syn_4  ;
	output \g233449/u3_syn_4  ;
	output \g233453/u3_syn_4  ;
	output \g233465/u3_syn_4  ;
	output \g233473/u3_syn_4  ;
	output \g233481/u3_syn_4  ;
	output \g233489/u3_syn_4  ;
	output \g233497/u3_syn_4  ;
	output \g233505/u3_syn_4  ;
	output \g233513/u3_syn_4  ;
	output \g233516/u3_syn_4  ;
	output \g233529/u3_syn_4  ;
	output \g233531/u3_syn_4  ;
	output \g233546/u3_syn_4  ;
	output \g233554/u3_syn_4  ;
	output \g233562/u3_syn_4  ;
	output \g233570/u3_syn_4  ;
	output \g233578/u3_syn_4  ;
	output \g233586/u3_syn_4  ;
	output \g233594/u3_syn_4  ;
	output \g233602/u3_syn_4  ;
	output \g233603/u3_syn_4  ;
	output \g233618/u3_syn_4  ;
	output \g233626/u3_syn_4  ;
	output \g233634/u3_syn_4  ;
	output \g233642/u3_syn_4  ;
	output \g233650/u3_syn_4  ;
	output \g233658/u3_syn_4  ;
	output \g233666/u3_syn_4  ;
	output \g233674/u3_syn_4  ;
	output \g233682/u3_syn_4  ;
	output \g233690/u3_syn_4  ;
	output \g233698/u3_syn_4  ;
	output \g233706/u3_syn_4  ;
	output \g233714/u3_syn_4  ;
	output \g233722/u3_syn_4  ;
	output \g233730/u3_syn_4  ;
	output \g233738/u3_syn_4  ;
	output \g233746/u3_syn_4  ;
	output \g233754/u3_syn_4  ;
	output \g233762/u3_syn_4  ;
	output \g233770/u3_syn_4  ;
	output \g233778/u3_syn_4  ;
	output \g233783/u3_syn_4  ;
	output \g233794/u3_syn_4  ;
	output \g233802/u3_syn_4  ;
	output \g233806/u3_syn_4  ;
	output \g233818/u3_syn_4  ;
	output \g233826/u3_syn_4  ;
	output \g233828/u3_syn_4  ;
	output \g233838/u3_syn_4  ;
	output \g233850/u3_syn_4  ;
	output \g233858/u3_syn_4  ;
	output \g233860/u3_syn_4  ;
	output \g233870/u3_syn_4  ;
	output \g233881/u3_syn_4  ;
	output \g233890/u3_syn_4  ;
	output \g233899/u3_syn_4  ;
	output \g233908/u3_syn_4  ;
	output \g233917/u3_syn_4  ;
	output \g233919/u3_syn_4  ;
	output \g233927/u3_syn_4  ;
	output \g233935/u3_syn_4  ;
	output \g233943/u3_syn_4  ;
	output \g233945/u3_syn_4  ;
	output \g233953/u3_syn_4  ;
	output \g233961/u3_syn_4  ;
	output \g233969/u3_syn_4  ;
	output \g233977/u3_syn_4  ;
	output \g233985/u3_syn_4  ;
	output \g233993/u3_syn_4  ;
	output \g234001/u3_syn_4  ;
	output \g234008/u3_syn_4  ;
	output \g234009/u3_syn_4  ;
	output \g234024/u3_syn_4  ;
	output \g234032/u3_syn_4  ;
	output \g234038/u3_syn_4  ;
	output \g234056/u3_syn_4  ;
	output \g234063/u3_syn_4  ;
	output \g234071/u3_syn_4  ;
	output \g234079/u3_syn_4  ;
	output \g234098/u3_syn_4  ;
	output \g234106/u3_syn_4  ;
	output \g234114/u3_syn_4  ;
	output \g234122/u3_syn_4  ;
	output \g234130/u3_syn_4  ;
	output \g234138/u3_syn_4  ;
	output \g234145/u3_syn_4  ;
	output \g234156/u3_syn_4  ;
	output \g234162/u3_syn_4  ;
	output \g234171/u3_syn_4  ;
	output \g234183/u3_syn_4  ;
	output \g234248/u3_syn_4  ;
	output \g234265/u3_syn_4  ;
	output \g234273/u3_syn_4  ;
	output \g234281/u3_syn_4  ;
	output \g234289/u3_syn_4  ;
	output \g234297/u3_syn_4  ;
	output \g234306/u3_syn_4  ;
	output \g234314/u3_syn_4  ;
	output \g234322/u3_syn_4  ;
	output \g234331/u3_syn_4  ;
	output \g234339/u3_syn_4  ;
	output \g234347/u3_syn_4  ;
	output \g234355/u3_syn_4  ;
	output \g234363/u3_syn_4  ;
	output \g234371/u3_syn_4  ;
	output \g234379/u3_syn_4  ;
	output \g234387/u3_syn_4  ;
	output \g234395/u3_syn_4  ;
	output \g234403/u3_syn_4  ;
	output \g234411/u3_syn_4  ;
	output \g234419/u3_syn_4  ;
	output \g234427/u3_syn_4  ;
	output \g234435/u3_syn_4  ;
	output \g234443/u3_syn_4  ;
	output \g234451/u3_syn_4  ;
	output \g234459/u3_syn_4  ;
	output \g234467/u3_syn_4  ;
	output \g234475/u3_syn_4  ;
	output \g234483/u3_syn_4  ;
	output \g234491/u3_syn_4  ;
	output \g234499/u3_syn_4  ;
	output \g234507/u3_syn_4  ;
	output \g234515/u3_syn_4  ;
	output \g234523/u3_syn_4  ;
	output \g234531/u3_syn_4  ;
	output \g234539/u3_syn_4  ;
	output \g234547/u3_syn_4  ;
	output \g234555/u3_syn_4  ;
	output \g234563/u3_syn_4  ;
	output \g234571/u3_syn_4  ;
	output \g234579/u3_syn_4  ;
	output \g234587/u3_syn_4  ;
	output \g234595/u3_syn_4  ;
	output \g234604/u3_syn_4  ;
	output \g234612/u3_syn_4  ;
	output \g234620/u3_syn_4  ;
	output \g234628/u3_syn_4  ;
	output \g234636/u3_syn_4  ;
	output \g234644/u3_syn_4  ;
	output \g234652/u3_syn_4  ;
	output \g234660/u3_syn_4  ;
	output \g234668/u3_syn_4  ;
	output \g234676/u3_syn_4  ;
	output \g234684/u3_syn_4  ;
	output \g234692/u3_syn_4  ;
	output \g234700/u3_syn_4  ;
	output \g234708/u3_syn_4  ;
	output \g234716/u3_syn_4  ;
	output \g234725/u3_syn_4  ;
	output \g234733/u3_syn_4  ;
	output \g234741/u3_syn_4  ;
	output \g234749/u3_syn_4  ;
	output \g234757/u3_syn_4  ;
	output \g234765/u3_syn_4  ;
	output \g234773/u3_syn_4  ;
	output \g234781/u3_syn_4  ;
	output \g234789/u3_syn_4  ;
	output \g234798/u3_syn_4  ;
	output \g234806/u3_syn_4  ;
	output \g234814/u3_syn_4  ;
	output \g234822/u3_syn_4  ;
	output \g234830/u3_syn_4  ;
	output \g234838/u3_syn_4  ;
	output \g235911/u3_syn_4  ;
	output \g235912/u3_syn_4  ;
	output \g235920/u3_syn_4  ;
	output \g235928/u3_syn_4  ;
	output \g235936/u3_syn_4  ;
	output \g235944/u3_syn_4  ;
	output \g235952/u3_syn_4  ;
	output \g235960/u3_syn_4  ;
	output \g235968/u3_syn_4  ;
	output \g235976/u3_syn_4  ;
	output \g235984/u3_syn_4  ;
	output \g235992/u3_syn_4  ;
	output \g236000/u3_syn_4  ;
	output \g236008/u3_syn_4  ;
	output \g236016/u3_syn_4  ;
	output \g236021/u3_syn_4  ;
	output \g236025/u3_syn_4  ;
	output \g236033/u3_syn_4  ;
	output \g236041/u3_syn_4  ;
	output \g236049/u3_syn_4  ;
	output \g236057/u3_syn_4  ;
	output \g236065/u3_syn_4  ;
	output \g236073/u3_syn_4  ;
	output \g236081/u3_syn_4  ;
	output \g236089/u3_syn_4  ;
	output \g236097/u3_syn_4  ;
	output \g236105/u3_syn_4  ;
	output \g236113/u3_syn_4  ;
	output \g236121/u3_syn_4  ;
	output \g236129/u3_syn_4  ;
	output \g236137/u3_syn_4  ;
	output \g236145/u3_syn_4  ;
	output \g236153/u3_syn_4  ;
	output \g236161/u3_syn_4  ;
	output \g236169/u3_syn_4  ;
	output \g236177/u3_syn_4  ;
	output \g236185/u3_syn_4  ;
	output \g236193/u3_syn_4  ;
	output \g236196/u3_syn_4  ;
	output \g236198/u3_syn_4  ;
	output \g236203/u3_syn_4  ;
	output \g236211/u3_syn_4  ;
	output \g236219/u3_syn_4  ;
	output \g236220/u3_syn_4  ;
	output \g236229/u3_syn_4  ;
	output \g236232/u3_syn_4  ;
	output \g236238/u3_syn_4  ;
	output \g236246/u3_syn_4  ;
	output \g236255/u3_syn_4  ;
	output \g236263/u3_syn_4  ;
	output \g236271/u3_syn_4  ;
	output \g236275/u3_syn_4  ;
	output \g236280/u3_syn_4  ;
	output \g236288/u3_syn_4  ;
	output \g236296/u3_syn_4  ;
	output \g236304/u3_syn_4  ;
	output \g236305/u3_syn_4  ;
	output \g236306/u3_syn_4  ;
	output \g236315/u3_syn_4  ;
	output \g236323/u3_syn_4  ;
	output \g236331/u3_syn_4  ;
	output \g236334/u3_syn_4  ;
	output \g236340/u3_syn_4  ;
	output \g236348/u3_syn_4  ;
	output \g236357/u3_syn_4  ;
	output \g236359/u3_syn_4  ;
	output \g236367/u3_syn_4  ;
	output \g236374/u3_syn_4  ;
	output \g236376/u3_syn_4  ;
	output \g236377/u3_syn_4  ;
	output \g236385/u3_syn_4  ;
	output \g236393/u3_syn_4  ;
	output \g236402/u3_syn_4  ;
	output \g236410/u3_syn_4  ;
	output \g236419/u3_syn_4  ;
	output \g236427/u3_syn_4  ;
	output \g236433/u3_syn_4  ;
	output \g236436/u3_syn_4  ;
	output \g236444/u3_syn_4  ;
	output \g236452/u3_syn_4  ;
	output \g236460/u3_syn_4  ;
	output \g236468/u3_syn_4  ;
	output \g236476/u3_syn_4  ;
	output \g236484/u3_syn_4  ;
	output \g236492/u3_syn_4  ;
	output \g236500/u3_syn_4  ;
	output \g236508/u3_syn_4  ;
	output \g236516/u3_syn_4  ;
	output \g236518/u3_syn_4  ;
	output \g236525/u3_syn_4  ;
	output \g236533/u3_syn_4  ;
	output \g236542/u3_syn_4  ;
	output \g236550/u3_syn_4  ;
	output \g236559/u3_syn_4  ;
	output \g236567/u3_syn_4  ;
	output \g236575/u3_syn_4  ;
	output \g236583/u3_syn_4  ;
	output \g236591/u3_syn_4  ;
	output \g236599/u3_syn_4  ;
	output \g236607/u3_syn_4  ;
	output \g236608/u3_syn_4  ;
	output \g236616/u3_syn_4  ;
	output \g236624/u3_syn_4  ;
	output \g236632/u3_syn_4  ;
	output \g236640/u3_syn_4  ;
	output \g236647/u3_syn_4  ;
	output \g236649/u3_syn_4  ;
	output \g236659/u3_syn_4  ;
	output \g236671/u3_syn_4  ;
	output \g236677/u3_syn_4  ;
	output \g236688/u3_syn_4  ;
	output \g236696/u3_syn_4  ;
	output \g236705/u3_syn_4  ;
	output \g236712/u3_syn_4  ;
	output \g236718/u3_syn_4  ;
	output \g236729/u3_syn_4  ;
	output \g236732/u3_syn_4  ;
	output \g236745/u3_syn_4  ;
	output \g236753/u3_syn_4  ;
	output \g236761/u3_syn_4  ;
	output \g236769/u3_syn_4  ;
	output \g236777/u3_syn_4  ;
	output \g236779/u3_syn_4  ;
	output \g236788/u3_syn_4  ;
	output \g236800/u3_syn_4  ;
	output \g236802/u3_syn_4  ;
	output \g236805/u3_syn_4  ;
	output \g236813/u3_syn_4  ;
	output \g236825/u3_syn_4  ;
	output \g236829/u3_syn_4  ;
	output \g236837/u3_syn_4  ;
	output \g236849/u3_syn_4  ;
	output \g236854/u3_syn_4  ;
	output \g236860/u3_syn_4  ;
	output \g236872/u3_syn_4  ;
	output \g236878/u3_syn_4  ;
	output \g236884/u3_syn_4  ;
	output \g236896/u3_syn_4  ;
	output \g236903/u3_syn_4  ;
	output \g236908/u3_syn_4  ;
	output \g236920/u3_syn_4  ;
	output \g236930/u3_syn_4  ;
	output \g236939/u3_syn_4  ;
	output \g236947/u3_syn_4  ;
	output \g236949/u3_syn_4  ;
	output \g236956/u3_syn_4  ;
	output \g236962/u3_syn_4  ;
	output \g236965/u3_syn_4  ;
	output \g236980/u3_syn_4  ;
	output \g236988/u3_syn_4  ;
	output \g236989/u3_syn_4  ;
	output \g237004/u3_syn_4  ;
	output \g237005/u3_syn_4  ;
	output \g237020/u3_syn_4  ;
	output \g237021/u3_syn_4  ;
	output \g237033/u3_syn_4  ;
	output \g237044/u3_syn_4  ;
	output \g237045/u3_syn_4  ;
	output \g237056/u3_syn_4  ;
	output \g237068/u3_syn_4  ;
	output \g237076/u3_syn_4  ;
	output \g237084/u3_syn_4  ;
	output \g237092/u3_syn_4  ;
	output \g237095/u3_syn_4  ;
	output \g237107/u3_syn_4  ;
	output \g237110/u3_syn_4  ;
	output \g237119/u3_syn_4  ;
	output \g237131/u3_syn_4  ;
	output \g237135/u3_syn_4  ;
	output \g237148/u3_syn_4  ;
	output \g237152/u3_syn_4  ;
	output \g237165/u3_syn_4  ;
	output \g237168/u3_syn_4  ;
	output \g237180/u3_syn_4  ;
	output \g237185/u3_syn_4  ;
	output \g237192/u3_syn_4  ;
	output \g237204/u3_syn_4  ;
	output \g237209/u3_syn_4  ;
	output \g237215/u3_syn_4  ;
	output \g237229/u3_syn_4  ;
	output \g237231/u3_syn_4  ;
	output \g237245/u3_syn_4  ;
	output \g237251/u3_syn_4  ;
	output \g237260/u3_syn_4  ;
	output \g237262/u3_syn_4  ;
	output \g237277/u3_syn_4  ;
	output \g237281/u3_syn_4  ;
	output \g237293/u3_syn_4  ;
	output \g237294/u3_syn_4  ;
	output \g237310/u3_syn_4  ;
	output \g237311/u3_syn_4  ;
	output \g237323/u3_syn_4  ;
	output \g237334/u3_syn_4  ;
	output \g237342/u3_syn_4  ;
	output \g237350/u3_syn_4  ;
	output \g237353/u3_syn_4  ;
	output \g237359/u3_syn_4  ;
	output \g237367/u3_syn_4  ;
	output \g237368/u3_syn_4  ;
	output \g237378/u3_syn_4  ;
	output \g237391/u3_syn_4  ;
	output \g237392/u3_syn_4  ;
	output \g237403/u3_syn_4  ;
	output \g237415/u3_syn_4  ;
	output \g237417/u3_syn_4  ;
	output \g237431/u3_syn_4  ;
	output \g237439/u3_syn_4  ;
	output \g237440/u3_syn_4  ;
	output \g237454/u3_syn_4  ;
	output \g237457/u3_syn_4  ;
	output \g237472/u3_syn_4  ;
	output \g237480/u3_syn_4  ;
	output \g237488/u3_syn_4  ;
	output \g237496/u3_syn_4  ;
	output \g237499/u3_syn_4  ;
	output \g237512/u3_syn_4  ;
	output \g237515/u3_syn_4  ;
	output \g237525/u3_syn_4  ;
	output \g237529/u3_syn_4  ;
	output \g237535/u3_syn_4  ;
	output \g237541/u3_syn_4  ;
	output \g237553/u3_syn_4  ;
	output \g237561/u3_syn_4  ;
	output \g237569/u3_syn_4  ;
	output \g237575/u3_syn_4  ;
	output \g237578/u3_syn_4  ;
	output \g237581/u3_syn_4  ;
	output \g237591/u3_syn_4  ;
	output \g237602/u3_syn_4  ;
	output \g237610/u3_syn_4  ;
	output \g237617/u3_syn_4  ;
	output \g237623/u3_syn_4  ;
	output \g237633/u3_syn_4  ;
	output \g237635/u3_syn_4  ;
	output \g237648/u3_syn_4  ;
	output \g237658/u3_syn_4  ;
	output \g237659/u3_syn_4  ;
	output \g237660/u3_syn_4  ;
	output \g237668/u3_syn_4  ;
	output \g237675/u3_syn_4  ;
	output \g237684/u3_syn_4  ;
	output \g237692/u3_syn_4  ;
	output \g237693/u3_syn_4  ;
	output \g237705/u3_syn_4  ;
	output \g237716/u3_syn_4  ;
	output \g237717/u3_syn_4  ;
	output \g237729/u3_syn_4  ;
	output \g237740/u3_syn_4  ;
	output \g237741/u3_syn_4  ;
	output \g237756/u3_syn_4  ;
	output \g237764/u3_syn_4  ;
	output \g237768/u3_syn_4  ;
	output \g237780/u3_syn_4  ;
	output \g237782/u3_syn_4  ;
	output \g237792/u3_syn_4  ;
	output \g237804/u3_syn_4  ;
	output \g237812/u3_syn_4  ;
	output \g237820/u3_syn_4  ;
	output \g237828/u3_syn_4  ;
	output \g237836/u3_syn_4  ;
	output \g237844/u3_syn_4  ;
	output \g237852/u3_syn_4  ;
	output \g237860/u3_syn_4  ;
	output \g237868/u3_syn_4  ;
	output \g237876/u3_syn_4  ;
	output \g237884/u3_syn_4  ;
	output \g237888/u3_syn_4  ;
	output \g237895/u3_syn_4  ;
	output \g237907/u3_syn_4  ;
	output \g237916/u3_syn_4  ;
	output \g237924/u3_syn_4  ;
	output \g237931/u3_syn_4  ;
	output \g237940/u3_syn_4  ;
	output \g237949/u3_syn_4  ;
	output \g237950/u3_syn_4  ;
	output \g237955/u3_syn_4  ;
	output \g237961/u3_syn_4  ;
	output \g237965/u3_syn_4  ;
	output \g237975/u3_syn_4  ;
	output \g237983/u3_syn_4  ;
	output \g237989/u3_syn_4  ;
	output \g237999/u3_syn_4  ;
	output \g238007/u3_syn_4  ;
	output \g238015/u3_syn_4  ;
	output \g238017/u3_syn_4  ;
	output \g238033/u3_syn_4  ;
	output \g238035/u3_syn_4  ;
	output \g238049/u3_syn_4  ;
	output \g238057/u3_syn_4  ;
	output \g238065/u3_syn_4  ;
	output \g238072/u3_syn_4  ;
	output \g238081/u3_syn_4  ;
	output \g238082/u3_syn_4  ;
	output \g238097/u3_syn_4  ;
	output \g238105/u3_syn_4  ;
	output \g238113/u3_syn_4  ;
	output \g238114/u3_syn_4  ;
	output \g238129/u3_syn_4  ;
	output \g238137/u3_syn_4  ;
	output \g238145/u3_syn_4  ;
	output \g238153/u3_syn_4  ;
	output \g238161/u3_syn_4  ;
	output \g238163/u3_syn_4  ;
	output \g238177/u3_syn_4  ;
	output \g238179/u3_syn_4  ;
	output \g238194/u3_syn_4  ;
	output \g238197/u3_syn_4  ;
	output \g238209/u3_syn_4  ;
	output \g238213/u3_syn_4  ;
	output \g238225/u3_syn_4  ;
	output \g238229/u3_syn_4  ;
	output \g238237/u3_syn_4  ;
	output \g238250/u3_syn_4  ;
	output \g238257/u3_syn_4  ;
	output \g238263/u3_syn_4  ;
	output \g238269/u3_syn_4  ;
	output \g238282/u3_syn_4  ;
	output \g238285/u3_syn_4  ;
	output \g238298/u3_syn_4  ;
	output \g238301/u3_syn_4  ;
	output \g238314/u3_syn_4  ;
	output \g238316/u3_syn_4  ;
	output \g238329/u3_syn_4  ;
	output \g238338/u3_syn_4  ;
	output \g238346/u3_syn_4  ;
	output \g238351/u3_syn_4  ;
	output \g238356/u3_syn_4  ;
	output \g238368/u3_syn_4  ;
	output \g238378/u3_syn_4  ;
	output \g238386/u3_syn_4  ;
	output \g238394/u3_syn_4  ;
	output \g238402/u3_syn_4  ;
	output \g238409/u3_syn_4  ;
	output \g238412/u3_syn_4  ;
	output \g238427/u3_syn_4  ;
	output \g238429/u3_syn_4  ;
	output \g238443/u3_syn_4  ;
	output \g238448/u3_syn_4  ;
	output \g238457/u3_syn_4  ;
	output \g238460/u3_syn_4  ;
	output \g238472/u3_syn_4  ;
	output \g238484/u3_syn_4  ;
	output \g238492/u3_syn_4  ;
	output \g238500/u3_syn_4  ;
	output \g238505/u3_syn_4  ;
	output \g238516/u3_syn_4  ;
	output \g238524/u3_syn_4  ;
	output \g238532/u3_syn_4  ;
	output \g238534/u3_syn_4  ;
	output \g238544/u3_syn_4  ;
	output \g238549/u3_syn_4  ;
	output \g238550/u3_syn_4  ;
	output \g238565/u3_syn_4  ;
	output \g238566/u3_syn_4  ;
	output \g238582/u3_syn_4  ;
	output \g238583/u3_syn_4  ;
	output \g238594/u3_syn_4  ;
	output \g238606/u3_syn_4  ;
	output \g238614/u3_syn_4  ;
	output \g238615/u3_syn_4  ;
	output \g238619/u3_syn_4  ;
	output \g238631/u3_syn_4  ;
	output \g238639/u3_syn_4  ;
	output \g238647/u3_syn_4  ;
	output \g238649/u3_syn_4  ;
	output \g238659/u3_syn_4  ;
	output \g238670/u3_syn_4  ;
	output \g238671/u3_syn_4  ;
	output \g238680/u3_syn_4  ;
	output \g238688/u3_syn_4  ;
	output \g238691/u3_syn_4  ;
	output \g238696/u3_syn_4  ;
	output \g238705/u3_syn_4  ;
	output \g238708/u3_syn_4  ;
	output \g238721/u3_syn_4  ;
	output \g238724/u3_syn_4  ;
	output \g238736/u3_syn_4  ;
	output \g238745/u3_syn_4  ;
	output \g238753/u3_syn_4  ;
	output \g238757/u3_syn_4  ;
	output \g238764/u3_syn_4  ;
	output \g238776/u3_syn_4  ;
	output \g238781/u3_syn_4  ;
	output \g238787/u3_syn_4  ;
	output \g238799/u3_syn_4  ;
	output \g238807/u3_syn_4  ;
	output \g238811/u3_syn_4  ;
	output \g238824/u3_syn_4  ;
	output \g238830/u3_syn_4  ;
	output \g238841/u3_syn_4  ;
	output \g238843/u3_syn_4  ;
	output \g238855/u3_syn_4  ;
	output \g238859/u3_syn_4  ;
	output \g238863/u3_syn_4  ;
	output \g238868/u3_syn_4  ;
	output \g238880/u3_syn_4  ;
	output \g238888/u3_syn_4  ;
	output \g238892/u3_syn_4  ;
	output \g238903/u3_syn_4  ;
	output \g238911/u3_syn_4  ;
	output \g238915/u3_syn_4  ;
	output \g238927/u3_syn_4  ;
	output \g238937/u3_syn_4  ;
	output \g238945/u3_syn_4  ;
	output \g238953/u3_syn_4  ;
	output \g238961/u3_syn_4  ;
	output \g238970/u3_syn_4  ;
	output \g238971/u3_syn_4  ;
	output \g238983/u3_syn_4  ;
	output \g238994/u3_syn_4  ;
	output \g239002/u3_syn_4  ;
	output \g239009/u3_syn_4  ;
	output \g239015/u3_syn_4  ;
	output \g239025/u3_syn_4  ;
	output \g239030/u3_syn_4  ;
	output \g239041/u3_syn_4  ;
	output \g239048/u3_syn_4  ;
	output \g239053/u3_syn_4  ;
	output \g239065/u3_syn_4  ;
	output \g239073/u3_syn_4  ;
	output \g239081/u3_syn_4  ;
	output \g239082/u3_syn_4  ;
	output \g239093/u3_syn_4  ;
	output \g239105/u3_syn_4  ;
	output \g239108/u3_syn_4  ;
	output \g239117/u3_syn_4  ;
	output \g239129/u3_syn_4  ;
	output \g239137/u3_syn_4  ;
	output \g239139/u3_syn_4  ;
	output \g239148/u3_syn_4  ;
	output \g239160/u3_syn_4  ;
	output \g239162/u3_syn_4  ;
	output \g239172/u3_syn_4  ;
	output \g239184/u3_syn_4  ;
	output \g239187/u3_syn_4  ;
	output \g239189/u3_syn_4  ;
	output \g239201/u3_syn_4  ;
	output \g239208/u3_syn_4  ;
	output \g239217/u3_syn_4  ;
	output \g239219/u3_syn_4  ;
	output \g239226/u3_syn_4  ;
	output \g239234/u3_syn_4  ;
	output \g239242/u3_syn_4  ;
	output \g239246/u3_syn_4  ;
	output \g239257/u3_syn_4  ;
	output \g239258/u3_syn_4  ;
	output \g239263/u3_syn_4  ;
	output \g239275/u3_syn_4  ;
	output \g239277/u3_syn_4  ;
	output \g239291/u3_syn_4  ;
	output \g239296/u3_syn_4  ;
	output \g239308/u3_syn_4  ;
	output \g239311/u3_syn_4  ;
	output \g239322/u3_syn_4  ;
	output \g239329/u3_syn_4  ;
	output \g239338/u3_syn_4  ;
	output \g239339/u3_syn_4  ;
	output \g239346/u3_syn_4  ;
	output \g239351/u3_syn_4  ;
	output \g239363/u3_syn_4  ;
	output \g239370/u3_syn_4  ;
	output \g239375/u3_syn_4  ;
	output \g239387/u3_syn_4  ;
	output \g239395/u3_syn_4  ;
	output \g239418/u3_syn_4  ;
	output \g239439/u3_syn_4  ;
	output \g239442/u3_syn_4  ;
	output \g239454/u3_syn_4  ;
	output \g239464/u3_syn_4  ;
	output \g239470/u3_syn_4  ;
	output \g239481/u3_syn_4  ;
	output \g239487/u3_syn_4  ;
	output \g239497/u3_syn_4  ;
	output \g239520/u3_syn_4  ;
	output \g239532/u3_syn_4  ;
	output \g239543/u3_syn_4  ;
	output \g239551/u3_syn_4  ;
	output \g239552/u3_syn_4  ;
	output \g239567/u3_syn_4  ;
	output \g239575/u3_syn_4  ;
	output \g239579/u3_syn_4  ;
	output \g239592/u3_syn_4  ;
	output \g239594/u3_syn_4  ;
	output \g239608/u3_syn_4  ;
	output \g239626/u3_syn_4  ;
	output \g239634/u3_syn_4  ;
	output \g239646/u3_syn_4  ;
	output \g239649/u3_syn_4  ;
	output \g239657/u3_syn_4  ;
	output \g239670/u3_syn_4  ;
	output \g239673/u3_syn_4  ;
	output \g239686/u3_syn_4  ;
	output \g239694/u3_syn_4  ;
	output \g239695/u3_syn_4  ;
	output \g239701/u3_syn_4  ;
	output \g239705/u3_syn_4  ;
	output \g239709/u3_syn_4  ;
	output \g239715/u3_syn_4  ;
	output \g239717/u3_syn_4  ;
	output \g239726/u3_syn_4  ;
	output \g239734/u3_syn_4  ;
	output \g239735/u3_syn_4  ;
	output \g239743/u3_syn_4  ;
	output \g239760/u3_syn_4  ;
	output \g239768/u3_syn_4  ;
	output \g239776/u3_syn_4  ;
	output \g239784/u3_syn_4  ;
	output \g239793/u3_syn_4  ;
	output \g239801/u3_syn_4  ;
	output \g239817/u3_syn_4  ;
	output \g239818/u3_syn_4  ;
	output \g239848/u3_syn_4  ;
	output \g239856/u3_syn_4  ;
	output \g239872/u3_syn_4  ;
	output \g239880/u3_syn_4  ;
	output \g239888/u3_syn_4  ;
	output \g239896/u3_syn_4  ;
	output \g239904/u3_syn_4  ;
	output \g239912/u3_syn_4  ;
	output \g239920/u3_syn_4  ;
	output \g239928/u3_syn_4  ;
	output \g239936/u3_syn_4  ;
	output \g239951/u3_syn_4  ;
	output \g239963/u3_syn_4  ;
	output \g239979/u3_syn_4  ;
	output \g239986/u3_syn_4  ;
	output \g239999/u3_syn_4  ;
	output \g240000/u3_syn_4  ;
	output \g240008/u3_syn_4  ;
	output \g240012/u3_syn_4  ;
	output \g240018/u3_syn_4  ;
	output \g240026/u3_syn_4  ;
	output \g240034/u3_syn_4  ;
	output \g240042/u3_syn_4  ;
	output \g240050/u3_syn_4  ;
	output \g240074/u3_syn_4  ;
	output \g240091/u3_syn_4  ;
	output \g240122/u3_syn_4  ;
	output \g240147/u3_syn_4  ;
	output \g240209/u3_syn_4  ;
	output \g240219/u3_syn_4  ;
	output \g240259/u3_syn_4  ;
	output \g240334/u3_syn_4  ;
	output \g240406/u3_syn_4  ;
	output \g240416/u3_syn_4  ;
	output \g240424/u3_syn_4  ;
	output \g240432/u3_syn_4  ;
	output \g240440/u3_syn_4  ;
	output \g240448/u3_syn_4  ;
	output \g240456/u3_syn_4  ;
	output \g240464/u3_syn_4  ;
	output \g240472/u3_syn_4  ;
	output \g240480/u3_syn_4  ;
	output \g240488/u3_syn_4  ;
	output \g240496/u3_syn_4  ;
	output \g240504/u3_syn_4  ;
	output \g240512/u3_syn_4  ;
	output \g240520/u3_syn_4  ;
	output \g240530/u3_syn_4  ;
	output \g240538/u3_syn_4  ;
	output \g240547/u3_syn_4  ;
	output \g240555/u3_syn_4  ;
	output \g240563/u3_syn_4  ;
	output \g240571/u3_syn_4  ;
	output \g240579/u3_syn_4  ;
	output \g240587/u3_syn_4  ;
	output \g240595/u3_syn_4  ;
	output \g240603/u3_syn_4  ;
	output \g240611/u3_syn_4  ;
	output \g240619/u3_syn_4  ;
	output \g240627/u3_syn_4  ;
	output \g240635/u3_syn_4  ;
	output \g240643/u3_syn_4  ;
	output \g240651/u3_syn_4  ;
	output \g240659/u3_syn_4  ;
	output \g240667/u3_syn_4  ;
	output \g240675/u3_syn_4  ;
	output \g240683/u3_syn_4  ;
	output \g240691/u3_syn_4  ;
	output \g240699/u3_syn_4  ;
	output \g240707/u3_syn_4  ;
	output \g240715/u3_syn_4  ;
	output \g240723/u3_syn_4  ;
	output \g240731/u3_syn_4  ;
	output \g240739/u3_syn_4  ;
	output \g240747/u3_syn_4  ;
	output \g240755/u3_syn_4  ;
	output \g240763/u3_syn_4  ;
	output \g240771/u3_syn_4  ;
	output \g240779/u3_syn_4  ;
	output \g240787/u3_syn_4  ;
	output \g240795/u3_syn_4  ;
	output \g240803/u3_syn_4  ;
	output \g240811/u3_syn_4  ;
	output \g240819/u3_syn_4  ;
	output \g240827/u3_syn_4  ;
	output \g240835/u3_syn_4  ;
	output \g240843/u3_syn_4  ;
	output \g240851/u3_syn_4  ;
	output \g240859/u3_syn_4  ;
	output \g240867/u3_syn_4  ;
	output \g240875/u3_syn_4  ;
	output \g240883/u3_syn_4  ;
	output \g240891/u3_syn_4  ;
	output \g240899/u3_syn_4  ;
	output \g240907/u3_syn_4  ;
	output \g240915/u3_syn_4  ;
	output \g240923/u3_syn_4  ;
	output \g240931/u3_syn_4  ;
	output \g240939/u3_syn_4  ;
	output \g240947/u3_syn_4  ;
	output \g240955/u3_syn_4  ;
	output \g240963/u3_syn_4  ;
	output \g240971/u3_syn_4  ;
	output \g240979/u3_syn_4  ;
	output \g240987/u3_syn_4  ;
	output \g240995/u3_syn_4  ;
	output \g241003/u3_syn_4  ;
	output \g241011/u3_syn_4  ;
	output \g241019/u3_syn_4  ;
	output \g241027/u3_syn_4  ;
	output \g241036/u3_syn_4  ;
	output \g241044/u3_syn_4  ;
	output \g241052/u3_syn_4  ;
	output \g241060/u3_syn_4  ;
	output \g241068/u3_syn_4  ;
	output \g241076/u3_syn_4  ;
	output \g241084/u3_syn_4  ;
	output \g241092/u3_syn_4  ;
	output \g241100/u3_syn_4  ;
	output \g241108/u3_syn_4  ;
	output \g241116/u3_syn_4  ;
	output \g241124/u3_syn_4  ;
	output \g241132/u3_syn_4  ;
	output \g241140/u3_syn_4  ;
	output \g241148/u3_syn_4  ;
	output \g241156/u3_syn_4  ;
	output \g241164/u3_syn_4  ;
	output \g241172/u3_syn_4  ;
	output \g241180/u3_syn_4  ;
	output \g241188/u3_syn_4  ;
	output \g241196/u3_syn_4  ;
	output \g241205/u3_syn_4  ;
	output \g241213/u3_syn_4  ;
	output \g241221/u3_syn_4  ;
	output \g241229/u3_syn_4  ;
	output \g241237/u3_syn_4  ;
	output \g241245/u3_syn_4  ;
	output \g241253/u3_syn_4  ;
	output \g241261/u3_syn_4  ;
	output \g241269/u3_syn_4  ;
	output \g241277/u3_syn_4  ;
	output \g241285/u3_syn_4  ;
	output \g241293/u3_syn_4  ;
	output \g241301/u3_syn_4  ;
	output \g241309/u3_syn_4  ;
	output \g241317/u3_syn_4  ;
	output \g241325/u3_syn_4  ;
	output \g241333/u3_syn_4  ;
	output \g241341/u3_syn_4  ;
	output \g241349/u3_syn_4  ;
	output \g241358/u3_syn_4  ;
	output \g241366/u3_syn_4  ;
	output \g241374/u3_syn_4  ;
	output \g241382/u3_syn_4  ;
	output \g241390/u3_syn_4  ;
	output \g241398/u3_syn_4  ;
	output \g241406/u3_syn_4  ;
	output \g241415/u3_syn_4  ;
	output \g241424/u3_syn_4  ;
	output \g241433/u3_syn_4  ;
	output \g241441/u3_syn_4  ;
	output \g241449/u3_syn_4  ;
	output \g241459/u3_syn_4  ;
	output \g241470/u3_syn_4  ;
	output \g241480/u3_syn_4  ;
	output \g241489/u3_syn_4  ;
	output \g241497/u3_syn_4  ;
	output \g241505/u3_syn_4  ;
	output \g241513/u3_syn_4  ;
	output \g241545/_3_  ;
	output \g241580/_00_  ;
	output \g241737/_0_  ;
	output \g241752/_0_  ;
	output \g241755/_0_  ;
	output \g241767/_2__syn_2  ;
	output \g241781/_1__syn_2  ;
	output \g241782/_0_  ;
	output \g241803/_1__syn_2  ;
	output \g241805/_0_  ;
	output \g241812/_1__syn_2  ;
	output \g241814/_1__syn_2  ;
	output \g241816/_1__syn_2  ;
	output \g241819/_1__syn_2  ;
	output \g241822/_1__syn_2  ;
	output \g241823/_0_  ;
	output \g241833/_1__syn_2  ;
	output \g241843/_1__syn_2  ;
	output \g241844/_1__syn_2  ;
	output \g241848/_1__syn_2  ;
	output \g241855/_1__syn_2  ;
	output \g241868/_1__syn_2  ;
	output \g242013/_1__syn_2  ;
	output \g242015/_1__syn_2  ;
	output \g242017/_1__syn_2  ;
	output \g242021/_1__syn_2  ;
	output \g242039/_1__syn_2  ;
	output \g242081/_0_  ;
	output \g242086/_0_  ;
	output \g242101/_3_  ;
	output \g242116/_0_  ;
	output \g242135/_2_  ;
	output \g242147/_0_  ;
	output \g242158/_0_  ;
	output \g242196/_0_  ;
	output \g242202/_0_  ;
	output \g242203/_0_  ;
	output \g242204/_0_  ;
	output \g242212/_0_  ;
	output \g242226/_01_  ;
	output \g242281/_0_  ;
	output \g242407/_0_  ;
	output \g242410/_0_  ;
	output \g242426/_0_  ;
	output \g242438/_2_  ;
	output \g242466/_0_  ;
	output \g242530/_0_  ;
	output \g242532/_0_  ;
	output \g243397/_0_  ;
	output \g245925/_0_  ;
	output \g245932/_0_  ;
	output \g245933/_0_  ;
	output \g245986/_3_  ;
	output \g250157/_3_  ;
	output \g250202/_0_  ;
	output \g250246/_1_  ;
	output \g250248/_0_  ;
	output \g250250/_0_  ;
	output \g250305/_0_  ;
	output \g250323/_0_  ;
	output \g250373/_0_  ;
	output \g250377/_0_  ;
	output \g250412/_0_  ;
	output \g250413/_0_  ;
	output \g250418/_0_  ;
	output \g250419/_0_  ;
	output \g250421/_0_  ;
	output \g250433/_0_  ;
	output \g250448/_3_  ;
	output \g250567/_3_  ;
	output \g258965/_0_  ;
	output \g259006/_0_  ;
	output \g259471/_0_  ;
	output \g259473/_2_  ;
	output \g260557/_0_  ;
	output \g261035/_0_  ;
	output \g261095/_3_  ;
	output \g261207/_2__syn_2  ;
	output \g261754/_0_  ;
	output \g262017/_0_  ;
	output \g262045/_0_  ;
	output \g262046/_0_  ;
	output \g262100/_3_  ;
	output \g263539/_1_  ;
	output \g263574/_0_  ;
	output \g263858/_0_  ;
	output \g264104/_1_  ;
	output \g264107/_1_  ;
	output \g264117/_0_  ;
	output \g264282/_0_  ;
	output \g264511/_0_  ;
	output \g264541/_0_  ;
	output \g264562/_0_  ;
	output \g264618/_0_  ;
	output \g264660/_0_  ;
	output \g264681/_3_  ;
	output \g264727/_0_  ;
	output \g265013/_0_  ;
	output \g265084/_0_  ;
	output \g265378/_0_  ;
	output \g265413/_0_  ;
	output \g265446/_0_  ;
	output \g265486/_0_  ;
	output \g265524/_3_  ;
	output \g265528/_3_  ;
	output \g265548/_3_  ;
	output \g265579/_0_  ;
	output \g265768/_0_  ;
	output \g265801/_0_  ;
	output \g265819/_1_  ;
	output \g265853/_0_  ;
	output \g265933/_0_  ;
	output \g266022/_0_  ;
	output \g266183/_1_  ;
	output \g281909/_0_  ;
	output \g281965/_1_  ;
	output \g282284/_1_  ;
	output \g282639/_1_  ;
	output \g283047/_0_  ;
	output \g283157/_1_  ;
	output \g283184/_0_  ;
	output \g283334/_3_  ;
	output int_o_pad ;
	output \m_wb_adr_o[0]_pad  ;
	output \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131_syn_2  ;
	output \wishbone_tx_fifo_fifo_reg[2][15]/P0001_reg_syn_3  ;
	output \wishbone_tx_fifo_fifo_reg[2][16]/P0001_reg_syn_3  ;
	output \wishbone_tx_fifo_fifo_reg[2][17]/P0001_reg_syn_3  ;
	output \wishbone_tx_fifo_fifo_reg[2][22]/P0001_reg_syn_3  ;
	output \wishbone_tx_fifo_fifo_reg[2][23]/P0001_reg_syn_3  ;
	output \wishbone_tx_fifo_fifo_reg[2][25]/P0001_reg_syn_3  ;
	output \wishbone_tx_fifo_fifo_reg[2][2]/P0001_reg_syn_3  ;
	wire _w28866_ ;
	wire _w28865_ ;
	wire _w28864_ ;
	wire _w28863_ ;
	wire _w28862_ ;
	wire _w28861_ ;
	wire _w28860_ ;
	wire _w28859_ ;
	wire _w28858_ ;
	wire _w28857_ ;
	wire _w28856_ ;
	wire _w28855_ ;
	wire _w28854_ ;
	wire _w28853_ ;
	wire _w28852_ ;
	wire _w28851_ ;
	wire _w28850_ ;
	wire _w28849_ ;
	wire _w28848_ ;
	wire _w28847_ ;
	wire _w28846_ ;
	wire _w28845_ ;
	wire _w28844_ ;
	wire _w28843_ ;
	wire _w28842_ ;
	wire _w28841_ ;
	wire _w28840_ ;
	wire _w28839_ ;
	wire _w28838_ ;
	wire _w28837_ ;
	wire _w28836_ ;
	wire _w28835_ ;
	wire _w28834_ ;
	wire _w28833_ ;
	wire _w28832_ ;
	wire _w28831_ ;
	wire _w28830_ ;
	wire _w28829_ ;
	wire _w28828_ ;
	wire _w28827_ ;
	wire _w28826_ ;
	wire _w28825_ ;
	wire _w28824_ ;
	wire _w28823_ ;
	wire _w28822_ ;
	wire _w28821_ ;
	wire _w28820_ ;
	wire _w28819_ ;
	wire _w28818_ ;
	wire _w28817_ ;
	wire _w28816_ ;
	wire _w28815_ ;
	wire _w28814_ ;
	wire _w28813_ ;
	wire _w28812_ ;
	wire _w28811_ ;
	wire _w28810_ ;
	wire _w28809_ ;
	wire _w28808_ ;
	wire _w28807_ ;
	wire _w28806_ ;
	wire _w28805_ ;
	wire _w28804_ ;
	wire _w28803_ ;
	wire _w28802_ ;
	wire _w28801_ ;
	wire _w28800_ ;
	wire _w28799_ ;
	wire _w28798_ ;
	wire _w28797_ ;
	wire _w28796_ ;
	wire _w28795_ ;
	wire _w28794_ ;
	wire _w28793_ ;
	wire _w28792_ ;
	wire _w28791_ ;
	wire _w28790_ ;
	wire _w28789_ ;
	wire _w28788_ ;
	wire _w28787_ ;
	wire _w28786_ ;
	wire _w28785_ ;
	wire _w28784_ ;
	wire _w28783_ ;
	wire _w28782_ ;
	wire _w28781_ ;
	wire _w28780_ ;
	wire _w28779_ ;
	wire _w28778_ ;
	wire _w28777_ ;
	wire _w28776_ ;
	wire _w28775_ ;
	wire _w28774_ ;
	wire _w28773_ ;
	wire _w28772_ ;
	wire _w28771_ ;
	wire _w28770_ ;
	wire _w28769_ ;
	wire _w28768_ ;
	wire _w28767_ ;
	wire _w28766_ ;
	wire _w28765_ ;
	wire _w28764_ ;
	wire _w28763_ ;
	wire _w28762_ ;
	wire _w28761_ ;
	wire _w28760_ ;
	wire _w28759_ ;
	wire _w28758_ ;
	wire _w28757_ ;
	wire _w28756_ ;
	wire _w28755_ ;
	wire _w28754_ ;
	wire _w28753_ ;
	wire _w28752_ ;
	wire _w28751_ ;
	wire _w28750_ ;
	wire _w28749_ ;
	wire _w28748_ ;
	wire _w28747_ ;
	wire _w28746_ ;
	wire _w28745_ ;
	wire _w28744_ ;
	wire _w28743_ ;
	wire _w28742_ ;
	wire _w28741_ ;
	wire _w28740_ ;
	wire _w28739_ ;
	wire _w28738_ ;
	wire _w28737_ ;
	wire _w28736_ ;
	wire _w28735_ ;
	wire _w28734_ ;
	wire _w28733_ ;
	wire _w28732_ ;
	wire _w28731_ ;
	wire _w28730_ ;
	wire _w28729_ ;
	wire _w28728_ ;
	wire _w28727_ ;
	wire _w28726_ ;
	wire _w28725_ ;
	wire _w28724_ ;
	wire _w28723_ ;
	wire _w28722_ ;
	wire _w28721_ ;
	wire _w28720_ ;
	wire _w28719_ ;
	wire _w28718_ ;
	wire _w28717_ ;
	wire _w28716_ ;
	wire _w28715_ ;
	wire _w28714_ ;
	wire _w28713_ ;
	wire _w28712_ ;
	wire _w28711_ ;
	wire _w28710_ ;
	wire _w28709_ ;
	wire _w28708_ ;
	wire _w28707_ ;
	wire _w28706_ ;
	wire _w28705_ ;
	wire _w28704_ ;
	wire _w28703_ ;
	wire _w28702_ ;
	wire _w28701_ ;
	wire _w28700_ ;
	wire _w28699_ ;
	wire _w28698_ ;
	wire _w28697_ ;
	wire _w28696_ ;
	wire _w28695_ ;
	wire _w28694_ ;
	wire _w28693_ ;
	wire _w28692_ ;
	wire _w28691_ ;
	wire _w28690_ ;
	wire _w28689_ ;
	wire _w28688_ ;
	wire _w28687_ ;
	wire _w28686_ ;
	wire _w28685_ ;
	wire _w28684_ ;
	wire _w28683_ ;
	wire _w28682_ ;
	wire _w28681_ ;
	wire _w28680_ ;
	wire _w28679_ ;
	wire _w28678_ ;
	wire _w28677_ ;
	wire _w28676_ ;
	wire _w28675_ ;
	wire _w28674_ ;
	wire _w28673_ ;
	wire _w28672_ ;
	wire _w28671_ ;
	wire _w28670_ ;
	wire _w28669_ ;
	wire _w28668_ ;
	wire _w28667_ ;
	wire _w28666_ ;
	wire _w28665_ ;
	wire _w28664_ ;
	wire _w28663_ ;
	wire _w28662_ ;
	wire _w28661_ ;
	wire _w28660_ ;
	wire _w28659_ ;
	wire _w28658_ ;
	wire _w28657_ ;
	wire _w28656_ ;
	wire _w28655_ ;
	wire _w28654_ ;
	wire _w28653_ ;
	wire _w28652_ ;
	wire _w28651_ ;
	wire _w28650_ ;
	wire _w28649_ ;
	wire _w28648_ ;
	wire _w28647_ ;
	wire _w28646_ ;
	wire _w28645_ ;
	wire _w28644_ ;
	wire _w28643_ ;
	wire _w28642_ ;
	wire _w28641_ ;
	wire _w28640_ ;
	wire _w28639_ ;
	wire _w28638_ ;
	wire _w28637_ ;
	wire _w28636_ ;
	wire _w28635_ ;
	wire _w28634_ ;
	wire _w28633_ ;
	wire _w28632_ ;
	wire _w28631_ ;
	wire _w28630_ ;
	wire _w28629_ ;
	wire _w28628_ ;
	wire _w28627_ ;
	wire _w28626_ ;
	wire _w28625_ ;
	wire _w28624_ ;
	wire _w28623_ ;
	wire _w28622_ ;
	wire _w28621_ ;
	wire _w28620_ ;
	wire _w28619_ ;
	wire _w28618_ ;
	wire _w28617_ ;
	wire _w28616_ ;
	wire _w28615_ ;
	wire _w28614_ ;
	wire _w28613_ ;
	wire _w28612_ ;
	wire _w28611_ ;
	wire _w28610_ ;
	wire _w28609_ ;
	wire _w28608_ ;
	wire _w28607_ ;
	wire _w28606_ ;
	wire _w28605_ ;
	wire _w28604_ ;
	wire _w28603_ ;
	wire _w28602_ ;
	wire _w28601_ ;
	wire _w28600_ ;
	wire _w28599_ ;
	wire _w28598_ ;
	wire _w28597_ ;
	wire _w28596_ ;
	wire _w28595_ ;
	wire _w28594_ ;
	wire _w28593_ ;
	wire _w28592_ ;
	wire _w28591_ ;
	wire _w28590_ ;
	wire _w28589_ ;
	wire _w28588_ ;
	wire _w28587_ ;
	wire _w28586_ ;
	wire _w28585_ ;
	wire _w28584_ ;
	wire _w28583_ ;
	wire _w28582_ ;
	wire _w28581_ ;
	wire _w28580_ ;
	wire _w28579_ ;
	wire _w28578_ ;
	wire _w28577_ ;
	wire _w28576_ ;
	wire _w28575_ ;
	wire _w28574_ ;
	wire _w28573_ ;
	wire _w28572_ ;
	wire _w28571_ ;
	wire _w28570_ ;
	wire _w28569_ ;
	wire _w28568_ ;
	wire _w28567_ ;
	wire _w28566_ ;
	wire _w28565_ ;
	wire _w28564_ ;
	wire _w28563_ ;
	wire _w28562_ ;
	wire _w28561_ ;
	wire _w28560_ ;
	wire _w28559_ ;
	wire _w28558_ ;
	wire _w28557_ ;
	wire _w28556_ ;
	wire _w28555_ ;
	wire _w28554_ ;
	wire _w28553_ ;
	wire _w28552_ ;
	wire _w28551_ ;
	wire _w28550_ ;
	wire _w28549_ ;
	wire _w28548_ ;
	wire _w28547_ ;
	wire _w28546_ ;
	wire _w28545_ ;
	wire _w28544_ ;
	wire _w28543_ ;
	wire _w28542_ ;
	wire _w28541_ ;
	wire _w28540_ ;
	wire _w28539_ ;
	wire _w28538_ ;
	wire _w28537_ ;
	wire _w28536_ ;
	wire _w28535_ ;
	wire _w28534_ ;
	wire _w28533_ ;
	wire _w28532_ ;
	wire _w28531_ ;
	wire _w28530_ ;
	wire _w28529_ ;
	wire _w28528_ ;
	wire _w28527_ ;
	wire _w28526_ ;
	wire _w28525_ ;
	wire _w28524_ ;
	wire _w28523_ ;
	wire _w28522_ ;
	wire _w28521_ ;
	wire _w28520_ ;
	wire _w28519_ ;
	wire _w28518_ ;
	wire _w28517_ ;
	wire _w28516_ ;
	wire _w28515_ ;
	wire _w28514_ ;
	wire _w28513_ ;
	wire _w28512_ ;
	wire _w28511_ ;
	wire _w28510_ ;
	wire _w28509_ ;
	wire _w28508_ ;
	wire _w28507_ ;
	wire _w28506_ ;
	wire _w28505_ ;
	wire _w28504_ ;
	wire _w28503_ ;
	wire _w28502_ ;
	wire _w28501_ ;
	wire _w28500_ ;
	wire _w28499_ ;
	wire _w28498_ ;
	wire _w28497_ ;
	wire _w28496_ ;
	wire _w28495_ ;
	wire _w28494_ ;
	wire _w28493_ ;
	wire _w28492_ ;
	wire _w28491_ ;
	wire _w28490_ ;
	wire _w28489_ ;
	wire _w28488_ ;
	wire _w28487_ ;
	wire _w28486_ ;
	wire _w28485_ ;
	wire _w28484_ ;
	wire _w28483_ ;
	wire _w28482_ ;
	wire _w28481_ ;
	wire _w28480_ ;
	wire _w28479_ ;
	wire _w28478_ ;
	wire _w28477_ ;
	wire _w28476_ ;
	wire _w28475_ ;
	wire _w28474_ ;
	wire _w28473_ ;
	wire _w28472_ ;
	wire _w28471_ ;
	wire _w28470_ ;
	wire _w28469_ ;
	wire _w28468_ ;
	wire _w28467_ ;
	wire _w28466_ ;
	wire _w28465_ ;
	wire _w28464_ ;
	wire _w28463_ ;
	wire _w28462_ ;
	wire _w28461_ ;
	wire _w28460_ ;
	wire _w28459_ ;
	wire _w28458_ ;
	wire _w28457_ ;
	wire _w28456_ ;
	wire _w28455_ ;
	wire _w28454_ ;
	wire _w28453_ ;
	wire _w28452_ ;
	wire _w28451_ ;
	wire _w28450_ ;
	wire _w28449_ ;
	wire _w28448_ ;
	wire _w28447_ ;
	wire _w28446_ ;
	wire _w28445_ ;
	wire _w28444_ ;
	wire _w28443_ ;
	wire _w28442_ ;
	wire _w28441_ ;
	wire _w28440_ ;
	wire _w28439_ ;
	wire _w28438_ ;
	wire _w28437_ ;
	wire _w28436_ ;
	wire _w28435_ ;
	wire _w28434_ ;
	wire _w28433_ ;
	wire _w28432_ ;
	wire _w28431_ ;
	wire _w28430_ ;
	wire _w28429_ ;
	wire _w28428_ ;
	wire _w28427_ ;
	wire _w28426_ ;
	wire _w28425_ ;
	wire _w28424_ ;
	wire _w28423_ ;
	wire _w28422_ ;
	wire _w28421_ ;
	wire _w28420_ ;
	wire _w28419_ ;
	wire _w28418_ ;
	wire _w28417_ ;
	wire _w28416_ ;
	wire _w28415_ ;
	wire _w28414_ ;
	wire _w28413_ ;
	wire _w28412_ ;
	wire _w28411_ ;
	wire _w28410_ ;
	wire _w28409_ ;
	wire _w28408_ ;
	wire _w28407_ ;
	wire _w28406_ ;
	wire _w28405_ ;
	wire _w28404_ ;
	wire _w28403_ ;
	wire _w28402_ ;
	wire _w28401_ ;
	wire _w28400_ ;
	wire _w28399_ ;
	wire _w28398_ ;
	wire _w28397_ ;
	wire _w28396_ ;
	wire _w28395_ ;
	wire _w28394_ ;
	wire _w28393_ ;
	wire _w28392_ ;
	wire _w28391_ ;
	wire _w28390_ ;
	wire _w28389_ ;
	wire _w28388_ ;
	wire _w28387_ ;
	wire _w28386_ ;
	wire _w28385_ ;
	wire _w28384_ ;
	wire _w28383_ ;
	wire _w28382_ ;
	wire _w28381_ ;
	wire _w28380_ ;
	wire _w28379_ ;
	wire _w28378_ ;
	wire _w28377_ ;
	wire _w28376_ ;
	wire _w28375_ ;
	wire _w28374_ ;
	wire _w28373_ ;
	wire _w28372_ ;
	wire _w28371_ ;
	wire _w28370_ ;
	wire _w28369_ ;
	wire _w28368_ ;
	wire _w28367_ ;
	wire _w28366_ ;
	wire _w28365_ ;
	wire _w28364_ ;
	wire _w28363_ ;
	wire _w28362_ ;
	wire _w28361_ ;
	wire _w28360_ ;
	wire _w28359_ ;
	wire _w28358_ ;
	wire _w28357_ ;
	wire _w28356_ ;
	wire _w28355_ ;
	wire _w28354_ ;
	wire _w28353_ ;
	wire _w28352_ ;
	wire _w28351_ ;
	wire _w28350_ ;
	wire _w28349_ ;
	wire _w28348_ ;
	wire _w28347_ ;
	wire _w28346_ ;
	wire _w28345_ ;
	wire _w28344_ ;
	wire _w28343_ ;
	wire _w28342_ ;
	wire _w28341_ ;
	wire _w28340_ ;
	wire _w28339_ ;
	wire _w28338_ ;
	wire _w28337_ ;
	wire _w28336_ ;
	wire _w28335_ ;
	wire _w28334_ ;
	wire _w28333_ ;
	wire _w28332_ ;
	wire _w28331_ ;
	wire _w28330_ ;
	wire _w28329_ ;
	wire _w28328_ ;
	wire _w28327_ ;
	wire _w28326_ ;
	wire _w28325_ ;
	wire _w28324_ ;
	wire _w28323_ ;
	wire _w28322_ ;
	wire _w28321_ ;
	wire _w28320_ ;
	wire _w28319_ ;
	wire _w28318_ ;
	wire _w28317_ ;
	wire _w28316_ ;
	wire _w28315_ ;
	wire _w28314_ ;
	wire _w28313_ ;
	wire _w28312_ ;
	wire _w28311_ ;
	wire _w28310_ ;
	wire _w28309_ ;
	wire _w28308_ ;
	wire _w28307_ ;
	wire _w28306_ ;
	wire _w28305_ ;
	wire _w28304_ ;
	wire _w28303_ ;
	wire _w28302_ ;
	wire _w28301_ ;
	wire _w28300_ ;
	wire _w28299_ ;
	wire _w28298_ ;
	wire _w28297_ ;
	wire _w28296_ ;
	wire _w28295_ ;
	wire _w28294_ ;
	wire _w28293_ ;
	wire _w28292_ ;
	wire _w28291_ ;
	wire _w28290_ ;
	wire _w28289_ ;
	wire _w28288_ ;
	wire _w28287_ ;
	wire _w28286_ ;
	wire _w28285_ ;
	wire _w28284_ ;
	wire _w28283_ ;
	wire _w28282_ ;
	wire _w28281_ ;
	wire _w28280_ ;
	wire _w28279_ ;
	wire _w28278_ ;
	wire _w28277_ ;
	wire _w28276_ ;
	wire _w28275_ ;
	wire _w28274_ ;
	wire _w28273_ ;
	wire _w28272_ ;
	wire _w28271_ ;
	wire _w28270_ ;
	wire _w28269_ ;
	wire _w28268_ ;
	wire _w28267_ ;
	wire _w28266_ ;
	wire _w28265_ ;
	wire _w28264_ ;
	wire _w28263_ ;
	wire _w28262_ ;
	wire _w28261_ ;
	wire _w28260_ ;
	wire _w28259_ ;
	wire _w28258_ ;
	wire _w28257_ ;
	wire _w28256_ ;
	wire _w28255_ ;
	wire _w28254_ ;
	wire _w28253_ ;
	wire _w28252_ ;
	wire _w28251_ ;
	wire _w28250_ ;
	wire _w28249_ ;
	wire _w28248_ ;
	wire _w28247_ ;
	wire _w28246_ ;
	wire _w28245_ ;
	wire _w28244_ ;
	wire _w28243_ ;
	wire _w28242_ ;
	wire _w28241_ ;
	wire _w28240_ ;
	wire _w28239_ ;
	wire _w28238_ ;
	wire _w28237_ ;
	wire _w28236_ ;
	wire _w28235_ ;
	wire _w28234_ ;
	wire _w28233_ ;
	wire _w28232_ ;
	wire _w28231_ ;
	wire _w28230_ ;
	wire _w28229_ ;
	wire _w28228_ ;
	wire _w28227_ ;
	wire _w28226_ ;
	wire _w28225_ ;
	wire _w28224_ ;
	wire _w28223_ ;
	wire _w28222_ ;
	wire _w28221_ ;
	wire _w28220_ ;
	wire _w28219_ ;
	wire _w28218_ ;
	wire _w28217_ ;
	wire _w28216_ ;
	wire _w28215_ ;
	wire _w28214_ ;
	wire _w28213_ ;
	wire _w28212_ ;
	wire _w28211_ ;
	wire _w28210_ ;
	wire _w28209_ ;
	wire _w28208_ ;
	wire _w28207_ ;
	wire _w28206_ ;
	wire _w28205_ ;
	wire _w28204_ ;
	wire _w28203_ ;
	wire _w28202_ ;
	wire _w28201_ ;
	wire _w28200_ ;
	wire _w28199_ ;
	wire _w28198_ ;
	wire _w28197_ ;
	wire _w28196_ ;
	wire _w28195_ ;
	wire _w28194_ ;
	wire _w28193_ ;
	wire _w28192_ ;
	wire _w28191_ ;
	wire _w28190_ ;
	wire _w28189_ ;
	wire _w28188_ ;
	wire _w28187_ ;
	wire _w28186_ ;
	wire _w28185_ ;
	wire _w28184_ ;
	wire _w28183_ ;
	wire _w28182_ ;
	wire _w28181_ ;
	wire _w28180_ ;
	wire _w28179_ ;
	wire _w28178_ ;
	wire _w28177_ ;
	wire _w28176_ ;
	wire _w28175_ ;
	wire _w28174_ ;
	wire _w28173_ ;
	wire _w28172_ ;
	wire _w28171_ ;
	wire _w28170_ ;
	wire _w28169_ ;
	wire _w28168_ ;
	wire _w28167_ ;
	wire _w28166_ ;
	wire _w28165_ ;
	wire _w28164_ ;
	wire _w28163_ ;
	wire _w28162_ ;
	wire _w28161_ ;
	wire _w28160_ ;
	wire _w28159_ ;
	wire _w28158_ ;
	wire _w28157_ ;
	wire _w28156_ ;
	wire _w28155_ ;
	wire _w28154_ ;
	wire _w28153_ ;
	wire _w28152_ ;
	wire _w28151_ ;
	wire _w28150_ ;
	wire _w28149_ ;
	wire _w28148_ ;
	wire _w28147_ ;
	wire _w28146_ ;
	wire _w28145_ ;
	wire _w28144_ ;
	wire _w28143_ ;
	wire _w28142_ ;
	wire _w28141_ ;
	wire _w28140_ ;
	wire _w28139_ ;
	wire _w28138_ ;
	wire _w28137_ ;
	wire _w28136_ ;
	wire _w28135_ ;
	wire _w28134_ ;
	wire _w28133_ ;
	wire _w28132_ ;
	wire _w28131_ ;
	wire _w28130_ ;
	wire _w28129_ ;
	wire _w28128_ ;
	wire _w28127_ ;
	wire _w28126_ ;
	wire _w28125_ ;
	wire _w28124_ ;
	wire _w28123_ ;
	wire _w28122_ ;
	wire _w28121_ ;
	wire _w28120_ ;
	wire _w28119_ ;
	wire _w28118_ ;
	wire _w28117_ ;
	wire _w28116_ ;
	wire _w28115_ ;
	wire _w28114_ ;
	wire _w28113_ ;
	wire _w28112_ ;
	wire _w28111_ ;
	wire _w28110_ ;
	wire _w28109_ ;
	wire _w28108_ ;
	wire _w28107_ ;
	wire _w28106_ ;
	wire _w28105_ ;
	wire _w28104_ ;
	wire _w28103_ ;
	wire _w28102_ ;
	wire _w28101_ ;
	wire _w28100_ ;
	wire _w28099_ ;
	wire _w28098_ ;
	wire _w28097_ ;
	wire _w28096_ ;
	wire _w28095_ ;
	wire _w28094_ ;
	wire _w28093_ ;
	wire _w28092_ ;
	wire _w28091_ ;
	wire _w28090_ ;
	wire _w28089_ ;
	wire _w28088_ ;
	wire _w28087_ ;
	wire _w28086_ ;
	wire _w28085_ ;
	wire _w28084_ ;
	wire _w28083_ ;
	wire _w28082_ ;
	wire _w28081_ ;
	wire _w28080_ ;
	wire _w28079_ ;
	wire _w28078_ ;
	wire _w28077_ ;
	wire _w28076_ ;
	wire _w28075_ ;
	wire _w28074_ ;
	wire _w28073_ ;
	wire _w28072_ ;
	wire _w28071_ ;
	wire _w28070_ ;
	wire _w28069_ ;
	wire _w28068_ ;
	wire _w28067_ ;
	wire _w28066_ ;
	wire _w28065_ ;
	wire _w28064_ ;
	wire _w28063_ ;
	wire _w28062_ ;
	wire _w28061_ ;
	wire _w28060_ ;
	wire _w28059_ ;
	wire _w28058_ ;
	wire _w28057_ ;
	wire _w28056_ ;
	wire _w28055_ ;
	wire _w28054_ ;
	wire _w28053_ ;
	wire _w28052_ ;
	wire _w28051_ ;
	wire _w28050_ ;
	wire _w28049_ ;
	wire _w28048_ ;
	wire _w28047_ ;
	wire _w28046_ ;
	wire _w28045_ ;
	wire _w28044_ ;
	wire _w28043_ ;
	wire _w28042_ ;
	wire _w28041_ ;
	wire _w28040_ ;
	wire _w28039_ ;
	wire _w28038_ ;
	wire _w28037_ ;
	wire _w28036_ ;
	wire _w28035_ ;
	wire _w28034_ ;
	wire _w28033_ ;
	wire _w28032_ ;
	wire _w28031_ ;
	wire _w28030_ ;
	wire _w28029_ ;
	wire _w28028_ ;
	wire _w28027_ ;
	wire _w28026_ ;
	wire _w28025_ ;
	wire _w28024_ ;
	wire _w28023_ ;
	wire _w28022_ ;
	wire _w28021_ ;
	wire _w28020_ ;
	wire _w28019_ ;
	wire _w28018_ ;
	wire _w28017_ ;
	wire _w28016_ ;
	wire _w28015_ ;
	wire _w28014_ ;
	wire _w28013_ ;
	wire _w28012_ ;
	wire _w28011_ ;
	wire _w28010_ ;
	wire _w28009_ ;
	wire _w28008_ ;
	wire _w28007_ ;
	wire _w28006_ ;
	wire _w28005_ ;
	wire _w28004_ ;
	wire _w28003_ ;
	wire _w28002_ ;
	wire _w28001_ ;
	wire _w28000_ ;
	wire _w27999_ ;
	wire _w27998_ ;
	wire _w27997_ ;
	wire _w27996_ ;
	wire _w27995_ ;
	wire _w27994_ ;
	wire _w27993_ ;
	wire _w27992_ ;
	wire _w27991_ ;
	wire _w27990_ ;
	wire _w27989_ ;
	wire _w27988_ ;
	wire _w27987_ ;
	wire _w27986_ ;
	wire _w27985_ ;
	wire _w27984_ ;
	wire _w27983_ ;
	wire _w27982_ ;
	wire _w27981_ ;
	wire _w27980_ ;
	wire _w27979_ ;
	wire _w27978_ ;
	wire _w27977_ ;
	wire _w27976_ ;
	wire _w27975_ ;
	wire _w27974_ ;
	wire _w27973_ ;
	wire _w27972_ ;
	wire _w27971_ ;
	wire _w27970_ ;
	wire _w27969_ ;
	wire _w27968_ ;
	wire _w27967_ ;
	wire _w27966_ ;
	wire _w27965_ ;
	wire _w27964_ ;
	wire _w27963_ ;
	wire _w27962_ ;
	wire _w27961_ ;
	wire _w27960_ ;
	wire _w27959_ ;
	wire _w27958_ ;
	wire _w27957_ ;
	wire _w27956_ ;
	wire _w27955_ ;
	wire _w27954_ ;
	wire _w27953_ ;
	wire _w27952_ ;
	wire _w27951_ ;
	wire _w27950_ ;
	wire _w27949_ ;
	wire _w27948_ ;
	wire _w27947_ ;
	wire _w27946_ ;
	wire _w27945_ ;
	wire _w27944_ ;
	wire _w27943_ ;
	wire _w27942_ ;
	wire _w27941_ ;
	wire _w27940_ ;
	wire _w27939_ ;
	wire _w27938_ ;
	wire _w27937_ ;
	wire _w27936_ ;
	wire _w27935_ ;
	wire _w27934_ ;
	wire _w27933_ ;
	wire _w27932_ ;
	wire _w27931_ ;
	wire _w27930_ ;
	wire _w27929_ ;
	wire _w27928_ ;
	wire _w27927_ ;
	wire _w27926_ ;
	wire _w27925_ ;
	wire _w27924_ ;
	wire _w27923_ ;
	wire _w27922_ ;
	wire _w27921_ ;
	wire _w27920_ ;
	wire _w27919_ ;
	wire _w27918_ ;
	wire _w27917_ ;
	wire _w27916_ ;
	wire _w27915_ ;
	wire _w27914_ ;
	wire _w27913_ ;
	wire _w27912_ ;
	wire _w27911_ ;
	wire _w27910_ ;
	wire _w27909_ ;
	wire _w27908_ ;
	wire _w27907_ ;
	wire _w27906_ ;
	wire _w27905_ ;
	wire _w27904_ ;
	wire _w27903_ ;
	wire _w27902_ ;
	wire _w27901_ ;
	wire _w27900_ ;
	wire _w27899_ ;
	wire _w27898_ ;
	wire _w27897_ ;
	wire _w27896_ ;
	wire _w27895_ ;
	wire _w27894_ ;
	wire _w27893_ ;
	wire _w27892_ ;
	wire _w27891_ ;
	wire _w27890_ ;
	wire _w27889_ ;
	wire _w27888_ ;
	wire _w27887_ ;
	wire _w27886_ ;
	wire _w27885_ ;
	wire _w27884_ ;
	wire _w27883_ ;
	wire _w27882_ ;
	wire _w27881_ ;
	wire _w27880_ ;
	wire _w27879_ ;
	wire _w27878_ ;
	wire _w27877_ ;
	wire _w27876_ ;
	wire _w27875_ ;
	wire _w27874_ ;
	wire _w27873_ ;
	wire _w27872_ ;
	wire _w27871_ ;
	wire _w27870_ ;
	wire _w27869_ ;
	wire _w27868_ ;
	wire _w27867_ ;
	wire _w27866_ ;
	wire _w27865_ ;
	wire _w27864_ ;
	wire _w27863_ ;
	wire _w27862_ ;
	wire _w27861_ ;
	wire _w27860_ ;
	wire _w27859_ ;
	wire _w27858_ ;
	wire _w27857_ ;
	wire _w27856_ ;
	wire _w27855_ ;
	wire _w27854_ ;
	wire _w27853_ ;
	wire _w27852_ ;
	wire _w27851_ ;
	wire _w27850_ ;
	wire _w27849_ ;
	wire _w27848_ ;
	wire _w27847_ ;
	wire _w27846_ ;
	wire _w27845_ ;
	wire _w27844_ ;
	wire _w27843_ ;
	wire _w27842_ ;
	wire _w27841_ ;
	wire _w27840_ ;
	wire _w27839_ ;
	wire _w27838_ ;
	wire _w27837_ ;
	wire _w27836_ ;
	wire _w27835_ ;
	wire _w27834_ ;
	wire _w27833_ ;
	wire _w27832_ ;
	wire _w27831_ ;
	wire _w27830_ ;
	wire _w27829_ ;
	wire _w27828_ ;
	wire _w27827_ ;
	wire _w27826_ ;
	wire _w27825_ ;
	wire _w27824_ ;
	wire _w27823_ ;
	wire _w27822_ ;
	wire _w27821_ ;
	wire _w27820_ ;
	wire _w27819_ ;
	wire _w27818_ ;
	wire _w27817_ ;
	wire _w27816_ ;
	wire _w27815_ ;
	wire _w27814_ ;
	wire _w27813_ ;
	wire _w27812_ ;
	wire _w27811_ ;
	wire _w27810_ ;
	wire _w27809_ ;
	wire _w27808_ ;
	wire _w27807_ ;
	wire _w27806_ ;
	wire _w27805_ ;
	wire _w27804_ ;
	wire _w27803_ ;
	wire _w27802_ ;
	wire _w27801_ ;
	wire _w27800_ ;
	wire _w27799_ ;
	wire _w27798_ ;
	wire _w27797_ ;
	wire _w27796_ ;
	wire _w27795_ ;
	wire _w27794_ ;
	wire _w27793_ ;
	wire _w27792_ ;
	wire _w27791_ ;
	wire _w27790_ ;
	wire _w27789_ ;
	wire _w27788_ ;
	wire _w27787_ ;
	wire _w27786_ ;
	wire _w27785_ ;
	wire _w27784_ ;
	wire _w27783_ ;
	wire _w27782_ ;
	wire _w27781_ ;
	wire _w27780_ ;
	wire _w27779_ ;
	wire _w27778_ ;
	wire _w27777_ ;
	wire _w27776_ ;
	wire _w27775_ ;
	wire _w27774_ ;
	wire _w27773_ ;
	wire _w27772_ ;
	wire _w27771_ ;
	wire _w27770_ ;
	wire _w27769_ ;
	wire _w27768_ ;
	wire _w27767_ ;
	wire _w27766_ ;
	wire _w27765_ ;
	wire _w27764_ ;
	wire _w27763_ ;
	wire _w27762_ ;
	wire _w27761_ ;
	wire _w27760_ ;
	wire _w27759_ ;
	wire _w27758_ ;
	wire _w27757_ ;
	wire _w27756_ ;
	wire _w27755_ ;
	wire _w27754_ ;
	wire _w27753_ ;
	wire _w27752_ ;
	wire _w27751_ ;
	wire _w27750_ ;
	wire _w27749_ ;
	wire _w27748_ ;
	wire _w27747_ ;
	wire _w27746_ ;
	wire _w27745_ ;
	wire _w27744_ ;
	wire _w27743_ ;
	wire _w27742_ ;
	wire _w27741_ ;
	wire _w27740_ ;
	wire _w27739_ ;
	wire _w27738_ ;
	wire _w27737_ ;
	wire _w27736_ ;
	wire _w27735_ ;
	wire _w27734_ ;
	wire _w27733_ ;
	wire _w27732_ ;
	wire _w27731_ ;
	wire _w27730_ ;
	wire _w27729_ ;
	wire _w27728_ ;
	wire _w27727_ ;
	wire _w27726_ ;
	wire _w27725_ ;
	wire _w27724_ ;
	wire _w27723_ ;
	wire _w27722_ ;
	wire _w27721_ ;
	wire _w27720_ ;
	wire _w27719_ ;
	wire _w27718_ ;
	wire _w27717_ ;
	wire _w27716_ ;
	wire _w27715_ ;
	wire _w27714_ ;
	wire _w27713_ ;
	wire _w27712_ ;
	wire _w27711_ ;
	wire _w27710_ ;
	wire _w27709_ ;
	wire _w27708_ ;
	wire _w27707_ ;
	wire _w27706_ ;
	wire _w27705_ ;
	wire _w27704_ ;
	wire _w27703_ ;
	wire _w27702_ ;
	wire _w27701_ ;
	wire _w27700_ ;
	wire _w27699_ ;
	wire _w27698_ ;
	wire _w27697_ ;
	wire _w27696_ ;
	wire _w27695_ ;
	wire _w27694_ ;
	wire _w27693_ ;
	wire _w27692_ ;
	wire _w27691_ ;
	wire _w27690_ ;
	wire _w27689_ ;
	wire _w27688_ ;
	wire _w27687_ ;
	wire _w27686_ ;
	wire _w27685_ ;
	wire _w27684_ ;
	wire _w27683_ ;
	wire _w27682_ ;
	wire _w27681_ ;
	wire _w27680_ ;
	wire _w27679_ ;
	wire _w27678_ ;
	wire _w27677_ ;
	wire _w27676_ ;
	wire _w27675_ ;
	wire _w27674_ ;
	wire _w27673_ ;
	wire _w27672_ ;
	wire _w27671_ ;
	wire _w27670_ ;
	wire _w27669_ ;
	wire _w27668_ ;
	wire _w27667_ ;
	wire _w27666_ ;
	wire _w27665_ ;
	wire _w27664_ ;
	wire _w27663_ ;
	wire _w27662_ ;
	wire _w27661_ ;
	wire _w27660_ ;
	wire _w27659_ ;
	wire _w27658_ ;
	wire _w27657_ ;
	wire _w27656_ ;
	wire _w27655_ ;
	wire _w27654_ ;
	wire _w27653_ ;
	wire _w27652_ ;
	wire _w27651_ ;
	wire _w27650_ ;
	wire _w27649_ ;
	wire _w27648_ ;
	wire _w27647_ ;
	wire _w27646_ ;
	wire _w27645_ ;
	wire _w27644_ ;
	wire _w27643_ ;
	wire _w27642_ ;
	wire _w27641_ ;
	wire _w27640_ ;
	wire _w27639_ ;
	wire _w27638_ ;
	wire _w27637_ ;
	wire _w27636_ ;
	wire _w27635_ ;
	wire _w27634_ ;
	wire _w27633_ ;
	wire _w27632_ ;
	wire _w27631_ ;
	wire _w27630_ ;
	wire _w27629_ ;
	wire _w27628_ ;
	wire _w27627_ ;
	wire _w27626_ ;
	wire _w27625_ ;
	wire _w27624_ ;
	wire _w27623_ ;
	wire _w27622_ ;
	wire _w27621_ ;
	wire _w27620_ ;
	wire _w27619_ ;
	wire _w27618_ ;
	wire _w27617_ ;
	wire _w27616_ ;
	wire _w27615_ ;
	wire _w27614_ ;
	wire _w27613_ ;
	wire _w27612_ ;
	wire _w27611_ ;
	wire _w27610_ ;
	wire _w27609_ ;
	wire _w27608_ ;
	wire _w27607_ ;
	wire _w27606_ ;
	wire _w27605_ ;
	wire _w27604_ ;
	wire _w27603_ ;
	wire _w27602_ ;
	wire _w27601_ ;
	wire _w27600_ ;
	wire _w27599_ ;
	wire _w27598_ ;
	wire _w27597_ ;
	wire _w27596_ ;
	wire _w27595_ ;
	wire _w27594_ ;
	wire _w27593_ ;
	wire _w27592_ ;
	wire _w27591_ ;
	wire _w27590_ ;
	wire _w27589_ ;
	wire _w27588_ ;
	wire _w27587_ ;
	wire _w27586_ ;
	wire _w27585_ ;
	wire _w27584_ ;
	wire _w27583_ ;
	wire _w27582_ ;
	wire _w27581_ ;
	wire _w27580_ ;
	wire _w27579_ ;
	wire _w27578_ ;
	wire _w27577_ ;
	wire _w27576_ ;
	wire _w27575_ ;
	wire _w27574_ ;
	wire _w27573_ ;
	wire _w27572_ ;
	wire _w27571_ ;
	wire _w27570_ ;
	wire _w27569_ ;
	wire _w27568_ ;
	wire _w27567_ ;
	wire _w27566_ ;
	wire _w27565_ ;
	wire _w27564_ ;
	wire _w27563_ ;
	wire _w27562_ ;
	wire _w27561_ ;
	wire _w27560_ ;
	wire _w27559_ ;
	wire _w27558_ ;
	wire _w27557_ ;
	wire _w27556_ ;
	wire _w27555_ ;
	wire _w27554_ ;
	wire _w27553_ ;
	wire _w27552_ ;
	wire _w27551_ ;
	wire _w27550_ ;
	wire _w27549_ ;
	wire _w27548_ ;
	wire _w27547_ ;
	wire _w27546_ ;
	wire _w27545_ ;
	wire _w27544_ ;
	wire _w27543_ ;
	wire _w27542_ ;
	wire _w27541_ ;
	wire _w27540_ ;
	wire _w27539_ ;
	wire _w27538_ ;
	wire _w27537_ ;
	wire _w27536_ ;
	wire _w27535_ ;
	wire _w27534_ ;
	wire _w27533_ ;
	wire _w27532_ ;
	wire _w27531_ ;
	wire _w27530_ ;
	wire _w27529_ ;
	wire _w27528_ ;
	wire _w27527_ ;
	wire _w27526_ ;
	wire _w27525_ ;
	wire _w27524_ ;
	wire _w27523_ ;
	wire _w27522_ ;
	wire _w27521_ ;
	wire _w27520_ ;
	wire _w27519_ ;
	wire _w27518_ ;
	wire _w27517_ ;
	wire _w27516_ ;
	wire _w27515_ ;
	wire _w27514_ ;
	wire _w27513_ ;
	wire _w27512_ ;
	wire _w27511_ ;
	wire _w27510_ ;
	wire _w27509_ ;
	wire _w27508_ ;
	wire _w27507_ ;
	wire _w27506_ ;
	wire _w27505_ ;
	wire _w27504_ ;
	wire _w27503_ ;
	wire _w27502_ ;
	wire _w27501_ ;
	wire _w27500_ ;
	wire _w27499_ ;
	wire _w27498_ ;
	wire _w27497_ ;
	wire _w27496_ ;
	wire _w27495_ ;
	wire _w27494_ ;
	wire _w27493_ ;
	wire _w27492_ ;
	wire _w27491_ ;
	wire _w27490_ ;
	wire _w27489_ ;
	wire _w27488_ ;
	wire _w27487_ ;
	wire _w27486_ ;
	wire _w27485_ ;
	wire _w27484_ ;
	wire _w27483_ ;
	wire _w27482_ ;
	wire _w27481_ ;
	wire _w27480_ ;
	wire _w27479_ ;
	wire _w27478_ ;
	wire _w27477_ ;
	wire _w27476_ ;
	wire _w27475_ ;
	wire _w27474_ ;
	wire _w27473_ ;
	wire _w27472_ ;
	wire _w27471_ ;
	wire _w27470_ ;
	wire _w27469_ ;
	wire _w27468_ ;
	wire _w27467_ ;
	wire _w27466_ ;
	wire _w27465_ ;
	wire _w27464_ ;
	wire _w27463_ ;
	wire _w27462_ ;
	wire _w27461_ ;
	wire _w27460_ ;
	wire _w27459_ ;
	wire _w27458_ ;
	wire _w27457_ ;
	wire _w27456_ ;
	wire _w27455_ ;
	wire _w27454_ ;
	wire _w27453_ ;
	wire _w27452_ ;
	wire _w27451_ ;
	wire _w27450_ ;
	wire _w27449_ ;
	wire _w27448_ ;
	wire _w27447_ ;
	wire _w27446_ ;
	wire _w27445_ ;
	wire _w27444_ ;
	wire _w27443_ ;
	wire _w27442_ ;
	wire _w27441_ ;
	wire _w27440_ ;
	wire _w27439_ ;
	wire _w27438_ ;
	wire _w27437_ ;
	wire _w27436_ ;
	wire _w27435_ ;
	wire _w27434_ ;
	wire _w27433_ ;
	wire _w27432_ ;
	wire _w27431_ ;
	wire _w27430_ ;
	wire _w27429_ ;
	wire _w27428_ ;
	wire _w27427_ ;
	wire _w27426_ ;
	wire _w27425_ ;
	wire _w27424_ ;
	wire _w27423_ ;
	wire _w27422_ ;
	wire _w27421_ ;
	wire _w27420_ ;
	wire _w27419_ ;
	wire _w27418_ ;
	wire _w27417_ ;
	wire _w27416_ ;
	wire _w27415_ ;
	wire _w27414_ ;
	wire _w27413_ ;
	wire _w27412_ ;
	wire _w27411_ ;
	wire _w27410_ ;
	wire _w27409_ ;
	wire _w27408_ ;
	wire _w27407_ ;
	wire _w27406_ ;
	wire _w27405_ ;
	wire _w27404_ ;
	wire _w27403_ ;
	wire _w27402_ ;
	wire _w27401_ ;
	wire _w27400_ ;
	wire _w27399_ ;
	wire _w27398_ ;
	wire _w27397_ ;
	wire _w27396_ ;
	wire _w27395_ ;
	wire _w27394_ ;
	wire _w27393_ ;
	wire _w27392_ ;
	wire _w27391_ ;
	wire _w27390_ ;
	wire _w27389_ ;
	wire _w27388_ ;
	wire _w27387_ ;
	wire _w27386_ ;
	wire _w27385_ ;
	wire _w27384_ ;
	wire _w27383_ ;
	wire _w27382_ ;
	wire _w27381_ ;
	wire _w27380_ ;
	wire _w27379_ ;
	wire _w27378_ ;
	wire _w27377_ ;
	wire _w27376_ ;
	wire _w27375_ ;
	wire _w27374_ ;
	wire _w27373_ ;
	wire _w27372_ ;
	wire _w27371_ ;
	wire _w27370_ ;
	wire _w27369_ ;
	wire _w27368_ ;
	wire _w27367_ ;
	wire _w27366_ ;
	wire _w27365_ ;
	wire _w27364_ ;
	wire _w27363_ ;
	wire _w27362_ ;
	wire _w27361_ ;
	wire _w27360_ ;
	wire _w27359_ ;
	wire _w27358_ ;
	wire _w27357_ ;
	wire _w27356_ ;
	wire _w27355_ ;
	wire _w27354_ ;
	wire _w27353_ ;
	wire _w27352_ ;
	wire _w27351_ ;
	wire _w27350_ ;
	wire _w27349_ ;
	wire _w27348_ ;
	wire _w27347_ ;
	wire _w27346_ ;
	wire _w27345_ ;
	wire _w27344_ ;
	wire _w27343_ ;
	wire _w27342_ ;
	wire _w27341_ ;
	wire _w27340_ ;
	wire _w27339_ ;
	wire _w27338_ ;
	wire _w27337_ ;
	wire _w27336_ ;
	wire _w27335_ ;
	wire _w27334_ ;
	wire _w27333_ ;
	wire _w27332_ ;
	wire _w27331_ ;
	wire _w27330_ ;
	wire _w27329_ ;
	wire _w27328_ ;
	wire _w27327_ ;
	wire _w27326_ ;
	wire _w27325_ ;
	wire _w27324_ ;
	wire _w27323_ ;
	wire _w27322_ ;
	wire _w27321_ ;
	wire _w27320_ ;
	wire _w27319_ ;
	wire _w27318_ ;
	wire _w27317_ ;
	wire _w27316_ ;
	wire _w27315_ ;
	wire _w27314_ ;
	wire _w27313_ ;
	wire _w27312_ ;
	wire _w27311_ ;
	wire _w27310_ ;
	wire _w27309_ ;
	wire _w27308_ ;
	wire _w27307_ ;
	wire _w27306_ ;
	wire _w27305_ ;
	wire _w27304_ ;
	wire _w27303_ ;
	wire _w27302_ ;
	wire _w27301_ ;
	wire _w27300_ ;
	wire _w27299_ ;
	wire _w27298_ ;
	wire _w27297_ ;
	wire _w27296_ ;
	wire _w27295_ ;
	wire _w27294_ ;
	wire _w27293_ ;
	wire _w27292_ ;
	wire _w27291_ ;
	wire _w27290_ ;
	wire _w27289_ ;
	wire _w27288_ ;
	wire _w27287_ ;
	wire _w27286_ ;
	wire _w27285_ ;
	wire _w27284_ ;
	wire _w27283_ ;
	wire _w27282_ ;
	wire _w27281_ ;
	wire _w27280_ ;
	wire _w27279_ ;
	wire _w27278_ ;
	wire _w27277_ ;
	wire _w27276_ ;
	wire _w27275_ ;
	wire _w27274_ ;
	wire _w27273_ ;
	wire _w27272_ ;
	wire _w27271_ ;
	wire _w27270_ ;
	wire _w27269_ ;
	wire _w27268_ ;
	wire _w27267_ ;
	wire _w27266_ ;
	wire _w27265_ ;
	wire _w27264_ ;
	wire _w27263_ ;
	wire _w27262_ ;
	wire _w27261_ ;
	wire _w27260_ ;
	wire _w27259_ ;
	wire _w27258_ ;
	wire _w27257_ ;
	wire _w27256_ ;
	wire _w27255_ ;
	wire _w27254_ ;
	wire _w27253_ ;
	wire _w27252_ ;
	wire _w27251_ ;
	wire _w27250_ ;
	wire _w27249_ ;
	wire _w27248_ ;
	wire _w27247_ ;
	wire _w27246_ ;
	wire _w27245_ ;
	wire _w27244_ ;
	wire _w27243_ ;
	wire _w27242_ ;
	wire _w27241_ ;
	wire _w27240_ ;
	wire _w27239_ ;
	wire _w27238_ ;
	wire _w27237_ ;
	wire _w27236_ ;
	wire _w27235_ ;
	wire _w27234_ ;
	wire _w27233_ ;
	wire _w27232_ ;
	wire _w27231_ ;
	wire _w27230_ ;
	wire _w27229_ ;
	wire _w27228_ ;
	wire _w27227_ ;
	wire _w27226_ ;
	wire _w27225_ ;
	wire _w27224_ ;
	wire _w27223_ ;
	wire _w27222_ ;
	wire _w27221_ ;
	wire _w27220_ ;
	wire _w27219_ ;
	wire _w27218_ ;
	wire _w27217_ ;
	wire _w27216_ ;
	wire _w27215_ ;
	wire _w27214_ ;
	wire _w27213_ ;
	wire _w27212_ ;
	wire _w27211_ ;
	wire _w27210_ ;
	wire _w27209_ ;
	wire _w27208_ ;
	wire _w27207_ ;
	wire _w27206_ ;
	wire _w27205_ ;
	wire _w27204_ ;
	wire _w27203_ ;
	wire _w27202_ ;
	wire _w27201_ ;
	wire _w27200_ ;
	wire _w27199_ ;
	wire _w27198_ ;
	wire _w27197_ ;
	wire _w27196_ ;
	wire _w27195_ ;
	wire _w27194_ ;
	wire _w27193_ ;
	wire _w27192_ ;
	wire _w27191_ ;
	wire _w27190_ ;
	wire _w27189_ ;
	wire _w27188_ ;
	wire _w27187_ ;
	wire _w27186_ ;
	wire _w27185_ ;
	wire _w27184_ ;
	wire _w27183_ ;
	wire _w27182_ ;
	wire _w27181_ ;
	wire _w27180_ ;
	wire _w27179_ ;
	wire _w27178_ ;
	wire _w27177_ ;
	wire _w27176_ ;
	wire _w27175_ ;
	wire _w27174_ ;
	wire _w27173_ ;
	wire _w27172_ ;
	wire _w27171_ ;
	wire _w27170_ ;
	wire _w27169_ ;
	wire _w27168_ ;
	wire _w27167_ ;
	wire _w27166_ ;
	wire _w27165_ ;
	wire _w27164_ ;
	wire _w27163_ ;
	wire _w27162_ ;
	wire _w27161_ ;
	wire _w27160_ ;
	wire _w27159_ ;
	wire _w27158_ ;
	wire _w27157_ ;
	wire _w27156_ ;
	wire _w27155_ ;
	wire _w27154_ ;
	wire _w27153_ ;
	wire _w27152_ ;
	wire _w27151_ ;
	wire _w27150_ ;
	wire _w27149_ ;
	wire _w27148_ ;
	wire _w27147_ ;
	wire _w27146_ ;
	wire _w27145_ ;
	wire _w27144_ ;
	wire _w27143_ ;
	wire _w27142_ ;
	wire _w27141_ ;
	wire _w27140_ ;
	wire _w27139_ ;
	wire _w27138_ ;
	wire _w27137_ ;
	wire _w27136_ ;
	wire _w27135_ ;
	wire _w27134_ ;
	wire _w27133_ ;
	wire _w27132_ ;
	wire _w27131_ ;
	wire _w27130_ ;
	wire _w27129_ ;
	wire _w27128_ ;
	wire _w27127_ ;
	wire _w27126_ ;
	wire _w27125_ ;
	wire _w27124_ ;
	wire _w27123_ ;
	wire _w27122_ ;
	wire _w27121_ ;
	wire _w27120_ ;
	wire _w27119_ ;
	wire _w27118_ ;
	wire _w27117_ ;
	wire _w27116_ ;
	wire _w27115_ ;
	wire _w27114_ ;
	wire _w27113_ ;
	wire _w27112_ ;
	wire _w27111_ ;
	wire _w27110_ ;
	wire _w27109_ ;
	wire _w27108_ ;
	wire _w27107_ ;
	wire _w27106_ ;
	wire _w27105_ ;
	wire _w27104_ ;
	wire _w27103_ ;
	wire _w27102_ ;
	wire _w27101_ ;
	wire _w27100_ ;
	wire _w27099_ ;
	wire _w27098_ ;
	wire _w27097_ ;
	wire _w27096_ ;
	wire _w27095_ ;
	wire _w27094_ ;
	wire _w27093_ ;
	wire _w27092_ ;
	wire _w27091_ ;
	wire _w27090_ ;
	wire _w27089_ ;
	wire _w27088_ ;
	wire _w27087_ ;
	wire _w27086_ ;
	wire _w27085_ ;
	wire _w27084_ ;
	wire _w27083_ ;
	wire _w27082_ ;
	wire _w27081_ ;
	wire _w27080_ ;
	wire _w27079_ ;
	wire _w27078_ ;
	wire _w27077_ ;
	wire _w27076_ ;
	wire _w27075_ ;
	wire _w27074_ ;
	wire _w27073_ ;
	wire _w27072_ ;
	wire _w27071_ ;
	wire _w27070_ ;
	wire _w27069_ ;
	wire _w27068_ ;
	wire _w27067_ ;
	wire _w27066_ ;
	wire _w27065_ ;
	wire _w27064_ ;
	wire _w27063_ ;
	wire _w27062_ ;
	wire _w27061_ ;
	wire _w27060_ ;
	wire _w27059_ ;
	wire _w27058_ ;
	wire _w27057_ ;
	wire _w27056_ ;
	wire _w27055_ ;
	wire _w27054_ ;
	wire _w27053_ ;
	wire _w27052_ ;
	wire _w27051_ ;
	wire _w27050_ ;
	wire _w27049_ ;
	wire _w27048_ ;
	wire _w27047_ ;
	wire _w27046_ ;
	wire _w27045_ ;
	wire _w27044_ ;
	wire _w27043_ ;
	wire _w27042_ ;
	wire _w27041_ ;
	wire _w27040_ ;
	wire _w27039_ ;
	wire _w27038_ ;
	wire _w27037_ ;
	wire _w27036_ ;
	wire _w27035_ ;
	wire _w27034_ ;
	wire _w27033_ ;
	wire _w27032_ ;
	wire _w27031_ ;
	wire _w27030_ ;
	wire _w27029_ ;
	wire _w27028_ ;
	wire _w27027_ ;
	wire _w27026_ ;
	wire _w27025_ ;
	wire _w27024_ ;
	wire _w27023_ ;
	wire _w27022_ ;
	wire _w27021_ ;
	wire _w27020_ ;
	wire _w27019_ ;
	wire _w27018_ ;
	wire _w27017_ ;
	wire _w27016_ ;
	wire _w27015_ ;
	wire _w27014_ ;
	wire _w27013_ ;
	wire _w27012_ ;
	wire _w27011_ ;
	wire _w27010_ ;
	wire _w27009_ ;
	wire _w27008_ ;
	wire _w27007_ ;
	wire _w27006_ ;
	wire _w27005_ ;
	wire _w27004_ ;
	wire _w27003_ ;
	wire _w27002_ ;
	wire _w27001_ ;
	wire _w27000_ ;
	wire _w26999_ ;
	wire _w26998_ ;
	wire _w26997_ ;
	wire _w26996_ ;
	wire _w26995_ ;
	wire _w26994_ ;
	wire _w26993_ ;
	wire _w26992_ ;
	wire _w26991_ ;
	wire _w26990_ ;
	wire _w26989_ ;
	wire _w26988_ ;
	wire _w26987_ ;
	wire _w26986_ ;
	wire _w26985_ ;
	wire _w26984_ ;
	wire _w26983_ ;
	wire _w26982_ ;
	wire _w26981_ ;
	wire _w26980_ ;
	wire _w26979_ ;
	wire _w26978_ ;
	wire _w26977_ ;
	wire _w26976_ ;
	wire _w26975_ ;
	wire _w26974_ ;
	wire _w26973_ ;
	wire _w26972_ ;
	wire _w26971_ ;
	wire _w26970_ ;
	wire _w26969_ ;
	wire _w26968_ ;
	wire _w26967_ ;
	wire _w26966_ ;
	wire _w26965_ ;
	wire _w26964_ ;
	wire _w26963_ ;
	wire _w26962_ ;
	wire _w26961_ ;
	wire _w26960_ ;
	wire _w26959_ ;
	wire _w26958_ ;
	wire _w26957_ ;
	wire _w26956_ ;
	wire _w26955_ ;
	wire _w26954_ ;
	wire _w26953_ ;
	wire _w26952_ ;
	wire _w26951_ ;
	wire _w26950_ ;
	wire _w26949_ ;
	wire _w26948_ ;
	wire _w26947_ ;
	wire _w26946_ ;
	wire _w26945_ ;
	wire _w26944_ ;
	wire _w26943_ ;
	wire _w26942_ ;
	wire _w26941_ ;
	wire _w26940_ ;
	wire _w26939_ ;
	wire _w26938_ ;
	wire _w26937_ ;
	wire _w26936_ ;
	wire _w26935_ ;
	wire _w26934_ ;
	wire _w26933_ ;
	wire _w26932_ ;
	wire _w26931_ ;
	wire _w26930_ ;
	wire _w26929_ ;
	wire _w26928_ ;
	wire _w26927_ ;
	wire _w26926_ ;
	wire _w26925_ ;
	wire _w26924_ ;
	wire _w26923_ ;
	wire _w26922_ ;
	wire _w26921_ ;
	wire _w26920_ ;
	wire _w26919_ ;
	wire _w26918_ ;
	wire _w26917_ ;
	wire _w26916_ ;
	wire _w26915_ ;
	wire _w26914_ ;
	wire _w26913_ ;
	wire _w26912_ ;
	wire _w26911_ ;
	wire _w26910_ ;
	wire _w26909_ ;
	wire _w26908_ ;
	wire _w26907_ ;
	wire _w26906_ ;
	wire _w26905_ ;
	wire _w26904_ ;
	wire _w26903_ ;
	wire _w26902_ ;
	wire _w26901_ ;
	wire _w26900_ ;
	wire _w26899_ ;
	wire _w26898_ ;
	wire _w26897_ ;
	wire _w26896_ ;
	wire _w26895_ ;
	wire _w26894_ ;
	wire _w26893_ ;
	wire _w26892_ ;
	wire _w26891_ ;
	wire _w26890_ ;
	wire _w26889_ ;
	wire _w26888_ ;
	wire _w26887_ ;
	wire _w26886_ ;
	wire _w26885_ ;
	wire _w26884_ ;
	wire _w26883_ ;
	wire _w26882_ ;
	wire _w26881_ ;
	wire _w26880_ ;
	wire _w26879_ ;
	wire _w26878_ ;
	wire _w26877_ ;
	wire _w26876_ ;
	wire _w26875_ ;
	wire _w26874_ ;
	wire _w26873_ ;
	wire _w26872_ ;
	wire _w26871_ ;
	wire _w26870_ ;
	wire _w26869_ ;
	wire _w26868_ ;
	wire _w26867_ ;
	wire _w26866_ ;
	wire _w26865_ ;
	wire _w26864_ ;
	wire _w26863_ ;
	wire _w26862_ ;
	wire _w26861_ ;
	wire _w26860_ ;
	wire _w26859_ ;
	wire _w26858_ ;
	wire _w26857_ ;
	wire _w26856_ ;
	wire _w26855_ ;
	wire _w26854_ ;
	wire _w26853_ ;
	wire _w26852_ ;
	wire _w26851_ ;
	wire _w26850_ ;
	wire _w26849_ ;
	wire _w26848_ ;
	wire _w26847_ ;
	wire _w26846_ ;
	wire _w26845_ ;
	wire _w26844_ ;
	wire _w26843_ ;
	wire _w26842_ ;
	wire _w26841_ ;
	wire _w26840_ ;
	wire _w26839_ ;
	wire _w26838_ ;
	wire _w26837_ ;
	wire _w26836_ ;
	wire _w26835_ ;
	wire _w26834_ ;
	wire _w26833_ ;
	wire _w26832_ ;
	wire _w26831_ ;
	wire _w26830_ ;
	wire _w26829_ ;
	wire _w26828_ ;
	wire _w26827_ ;
	wire _w26826_ ;
	wire _w26825_ ;
	wire _w26824_ ;
	wire _w26823_ ;
	wire _w26822_ ;
	wire _w26821_ ;
	wire _w26820_ ;
	wire _w26819_ ;
	wire _w26818_ ;
	wire _w26817_ ;
	wire _w26816_ ;
	wire _w26815_ ;
	wire _w26814_ ;
	wire _w26813_ ;
	wire _w26812_ ;
	wire _w26811_ ;
	wire _w26810_ ;
	wire _w26809_ ;
	wire _w26808_ ;
	wire _w26807_ ;
	wire _w26806_ ;
	wire _w26805_ ;
	wire _w26804_ ;
	wire _w26803_ ;
	wire _w26802_ ;
	wire _w26801_ ;
	wire _w26800_ ;
	wire _w26799_ ;
	wire _w26798_ ;
	wire _w26797_ ;
	wire _w26796_ ;
	wire _w26795_ ;
	wire _w26794_ ;
	wire _w26793_ ;
	wire _w26792_ ;
	wire _w26791_ ;
	wire _w26790_ ;
	wire _w26789_ ;
	wire _w26788_ ;
	wire _w26787_ ;
	wire _w26786_ ;
	wire _w26785_ ;
	wire _w26784_ ;
	wire _w26783_ ;
	wire _w26782_ ;
	wire _w26781_ ;
	wire _w26780_ ;
	wire _w26779_ ;
	wire _w26778_ ;
	wire _w26777_ ;
	wire _w26776_ ;
	wire _w26775_ ;
	wire _w26774_ ;
	wire _w26773_ ;
	wire _w26772_ ;
	wire _w26771_ ;
	wire _w26770_ ;
	wire _w26769_ ;
	wire _w26768_ ;
	wire _w26767_ ;
	wire _w26766_ ;
	wire _w26765_ ;
	wire _w26764_ ;
	wire _w26763_ ;
	wire _w26762_ ;
	wire _w26761_ ;
	wire _w26760_ ;
	wire _w26759_ ;
	wire _w26758_ ;
	wire _w26757_ ;
	wire _w26756_ ;
	wire _w26755_ ;
	wire _w26754_ ;
	wire _w26753_ ;
	wire _w26752_ ;
	wire _w26751_ ;
	wire _w26750_ ;
	wire _w26749_ ;
	wire _w26748_ ;
	wire _w26747_ ;
	wire _w26746_ ;
	wire _w26745_ ;
	wire _w26744_ ;
	wire _w26743_ ;
	wire _w26742_ ;
	wire _w26741_ ;
	wire _w26740_ ;
	wire _w26739_ ;
	wire _w26738_ ;
	wire _w26737_ ;
	wire _w26736_ ;
	wire _w26735_ ;
	wire _w26734_ ;
	wire _w26733_ ;
	wire _w26732_ ;
	wire _w26731_ ;
	wire _w26730_ ;
	wire _w26729_ ;
	wire _w26728_ ;
	wire _w26727_ ;
	wire _w26726_ ;
	wire _w26725_ ;
	wire _w26724_ ;
	wire _w26723_ ;
	wire _w26722_ ;
	wire _w26721_ ;
	wire _w26720_ ;
	wire _w26719_ ;
	wire _w26718_ ;
	wire _w26717_ ;
	wire _w26716_ ;
	wire _w26715_ ;
	wire _w26714_ ;
	wire _w26713_ ;
	wire _w26712_ ;
	wire _w26711_ ;
	wire _w26710_ ;
	wire _w26709_ ;
	wire _w26708_ ;
	wire _w26707_ ;
	wire _w26706_ ;
	wire _w26705_ ;
	wire _w26704_ ;
	wire _w26703_ ;
	wire _w26702_ ;
	wire _w26701_ ;
	wire _w26700_ ;
	wire _w26699_ ;
	wire _w26698_ ;
	wire _w26697_ ;
	wire _w26696_ ;
	wire _w26695_ ;
	wire _w26694_ ;
	wire _w26693_ ;
	wire _w26692_ ;
	wire _w26691_ ;
	wire _w26690_ ;
	wire _w26689_ ;
	wire _w26688_ ;
	wire _w26687_ ;
	wire _w26686_ ;
	wire _w26685_ ;
	wire _w26684_ ;
	wire _w26683_ ;
	wire _w26682_ ;
	wire _w26681_ ;
	wire _w26680_ ;
	wire _w26679_ ;
	wire _w26678_ ;
	wire _w26677_ ;
	wire _w26676_ ;
	wire _w26675_ ;
	wire _w26674_ ;
	wire _w26673_ ;
	wire _w26672_ ;
	wire _w26671_ ;
	wire _w26670_ ;
	wire _w26669_ ;
	wire _w26668_ ;
	wire _w26667_ ;
	wire _w26666_ ;
	wire _w26665_ ;
	wire _w26664_ ;
	wire _w26663_ ;
	wire _w26662_ ;
	wire _w26661_ ;
	wire _w26660_ ;
	wire _w26659_ ;
	wire _w26658_ ;
	wire _w26657_ ;
	wire _w26656_ ;
	wire _w26655_ ;
	wire _w26654_ ;
	wire _w26653_ ;
	wire _w26652_ ;
	wire _w26651_ ;
	wire _w26650_ ;
	wire _w26649_ ;
	wire _w26648_ ;
	wire _w26647_ ;
	wire _w26646_ ;
	wire _w26645_ ;
	wire _w26644_ ;
	wire _w26643_ ;
	wire _w26642_ ;
	wire _w26641_ ;
	wire _w26640_ ;
	wire _w26639_ ;
	wire _w26638_ ;
	wire _w26637_ ;
	wire _w26636_ ;
	wire _w26635_ ;
	wire _w26634_ ;
	wire _w26633_ ;
	wire _w26632_ ;
	wire _w26631_ ;
	wire _w26630_ ;
	wire _w26629_ ;
	wire _w26628_ ;
	wire _w26627_ ;
	wire _w26626_ ;
	wire _w26625_ ;
	wire _w26624_ ;
	wire _w26623_ ;
	wire _w26622_ ;
	wire _w26621_ ;
	wire _w26620_ ;
	wire _w26619_ ;
	wire _w26618_ ;
	wire _w26617_ ;
	wire _w26616_ ;
	wire _w26615_ ;
	wire _w26614_ ;
	wire _w26613_ ;
	wire _w26612_ ;
	wire _w26611_ ;
	wire _w26610_ ;
	wire _w26609_ ;
	wire _w26608_ ;
	wire _w26607_ ;
	wire _w26606_ ;
	wire _w26605_ ;
	wire _w26604_ ;
	wire _w26603_ ;
	wire _w26602_ ;
	wire _w26601_ ;
	wire _w26600_ ;
	wire _w26599_ ;
	wire _w26598_ ;
	wire _w26597_ ;
	wire _w26596_ ;
	wire _w26595_ ;
	wire _w26594_ ;
	wire _w26593_ ;
	wire _w26592_ ;
	wire _w26591_ ;
	wire _w26590_ ;
	wire _w26589_ ;
	wire _w26588_ ;
	wire _w26587_ ;
	wire _w26586_ ;
	wire _w26585_ ;
	wire _w26584_ ;
	wire _w26583_ ;
	wire _w26582_ ;
	wire _w26581_ ;
	wire _w26580_ ;
	wire _w26579_ ;
	wire _w26578_ ;
	wire _w26577_ ;
	wire _w26576_ ;
	wire _w26575_ ;
	wire _w26574_ ;
	wire _w26573_ ;
	wire _w26572_ ;
	wire _w26571_ ;
	wire _w26570_ ;
	wire _w26569_ ;
	wire _w26568_ ;
	wire _w26567_ ;
	wire _w26566_ ;
	wire _w26565_ ;
	wire _w26564_ ;
	wire _w26563_ ;
	wire _w26562_ ;
	wire _w26561_ ;
	wire _w26560_ ;
	wire _w26559_ ;
	wire _w26558_ ;
	wire _w26557_ ;
	wire _w26556_ ;
	wire _w26555_ ;
	wire _w26554_ ;
	wire _w26553_ ;
	wire _w26552_ ;
	wire _w26551_ ;
	wire _w26550_ ;
	wire _w26549_ ;
	wire _w26548_ ;
	wire _w26547_ ;
	wire _w26546_ ;
	wire _w26545_ ;
	wire _w26544_ ;
	wire _w26543_ ;
	wire _w26542_ ;
	wire _w26541_ ;
	wire _w26540_ ;
	wire _w26539_ ;
	wire _w26538_ ;
	wire _w26537_ ;
	wire _w26536_ ;
	wire _w26535_ ;
	wire _w26534_ ;
	wire _w26533_ ;
	wire _w26532_ ;
	wire _w26531_ ;
	wire _w26530_ ;
	wire _w26529_ ;
	wire _w26528_ ;
	wire _w26527_ ;
	wire _w26526_ ;
	wire _w26525_ ;
	wire _w26524_ ;
	wire _w26523_ ;
	wire _w26522_ ;
	wire _w26521_ ;
	wire _w26520_ ;
	wire _w26519_ ;
	wire _w26518_ ;
	wire _w26517_ ;
	wire _w26516_ ;
	wire _w26515_ ;
	wire _w26514_ ;
	wire _w26513_ ;
	wire _w26512_ ;
	wire _w26511_ ;
	wire _w26510_ ;
	wire _w26509_ ;
	wire _w26508_ ;
	wire _w26507_ ;
	wire _w26506_ ;
	wire _w26505_ ;
	wire _w26504_ ;
	wire _w26503_ ;
	wire _w26502_ ;
	wire _w26501_ ;
	wire _w26500_ ;
	wire _w26499_ ;
	wire _w26498_ ;
	wire _w26497_ ;
	wire _w26496_ ;
	wire _w26495_ ;
	wire _w26494_ ;
	wire _w26493_ ;
	wire _w26492_ ;
	wire _w26491_ ;
	wire _w26490_ ;
	wire _w26489_ ;
	wire _w26488_ ;
	wire _w26487_ ;
	wire _w26486_ ;
	wire _w26485_ ;
	wire _w26484_ ;
	wire _w26483_ ;
	wire _w26482_ ;
	wire _w26481_ ;
	wire _w26480_ ;
	wire _w26479_ ;
	wire _w26478_ ;
	wire _w26477_ ;
	wire _w26476_ ;
	wire _w26475_ ;
	wire _w26474_ ;
	wire _w26473_ ;
	wire _w26472_ ;
	wire _w26471_ ;
	wire _w26470_ ;
	wire _w26469_ ;
	wire _w26468_ ;
	wire _w26467_ ;
	wire _w26466_ ;
	wire _w26465_ ;
	wire _w26464_ ;
	wire _w26463_ ;
	wire _w26462_ ;
	wire _w26461_ ;
	wire _w26460_ ;
	wire _w26459_ ;
	wire _w26458_ ;
	wire _w26457_ ;
	wire _w26456_ ;
	wire _w26455_ ;
	wire _w26454_ ;
	wire _w26453_ ;
	wire _w26452_ ;
	wire _w26451_ ;
	wire _w26450_ ;
	wire _w26449_ ;
	wire _w26448_ ;
	wire _w26447_ ;
	wire _w26446_ ;
	wire _w26445_ ;
	wire _w26444_ ;
	wire _w26443_ ;
	wire _w26442_ ;
	wire _w26441_ ;
	wire _w26440_ ;
	wire _w26439_ ;
	wire _w26438_ ;
	wire _w26437_ ;
	wire _w26436_ ;
	wire _w26435_ ;
	wire _w26434_ ;
	wire _w26433_ ;
	wire _w26432_ ;
	wire _w26431_ ;
	wire _w26430_ ;
	wire _w26429_ ;
	wire _w26428_ ;
	wire _w26427_ ;
	wire _w26426_ ;
	wire _w26425_ ;
	wire _w26424_ ;
	wire _w26423_ ;
	wire _w26422_ ;
	wire _w26421_ ;
	wire _w26420_ ;
	wire _w26419_ ;
	wire _w26418_ ;
	wire _w26417_ ;
	wire _w26416_ ;
	wire _w26415_ ;
	wire _w26414_ ;
	wire _w26413_ ;
	wire _w26412_ ;
	wire _w26411_ ;
	wire _w26410_ ;
	wire _w26409_ ;
	wire _w26408_ ;
	wire _w26407_ ;
	wire _w26406_ ;
	wire _w26405_ ;
	wire _w26404_ ;
	wire _w26403_ ;
	wire _w26402_ ;
	wire _w26401_ ;
	wire _w26400_ ;
	wire _w26399_ ;
	wire _w26398_ ;
	wire _w26397_ ;
	wire _w26396_ ;
	wire _w26395_ ;
	wire _w26394_ ;
	wire _w26393_ ;
	wire _w26392_ ;
	wire _w26391_ ;
	wire _w26390_ ;
	wire _w26389_ ;
	wire _w26388_ ;
	wire _w26387_ ;
	wire _w26386_ ;
	wire _w26385_ ;
	wire _w26384_ ;
	wire _w26383_ ;
	wire _w26382_ ;
	wire _w26381_ ;
	wire _w26380_ ;
	wire _w26379_ ;
	wire _w26378_ ;
	wire _w26377_ ;
	wire _w26376_ ;
	wire _w26375_ ;
	wire _w26374_ ;
	wire _w26373_ ;
	wire _w26372_ ;
	wire _w26371_ ;
	wire _w26370_ ;
	wire _w26369_ ;
	wire _w26368_ ;
	wire _w26367_ ;
	wire _w26366_ ;
	wire _w26365_ ;
	wire _w26364_ ;
	wire _w26363_ ;
	wire _w26362_ ;
	wire _w26361_ ;
	wire _w26360_ ;
	wire _w26359_ ;
	wire _w26358_ ;
	wire _w26357_ ;
	wire _w26356_ ;
	wire _w26355_ ;
	wire _w26354_ ;
	wire _w26353_ ;
	wire _w26352_ ;
	wire _w26351_ ;
	wire _w26350_ ;
	wire _w26349_ ;
	wire _w26348_ ;
	wire _w26347_ ;
	wire _w26346_ ;
	wire _w26345_ ;
	wire _w26344_ ;
	wire _w26343_ ;
	wire _w26342_ ;
	wire _w26341_ ;
	wire _w26340_ ;
	wire _w26339_ ;
	wire _w26338_ ;
	wire _w26337_ ;
	wire _w26336_ ;
	wire _w26335_ ;
	wire _w26334_ ;
	wire _w26333_ ;
	wire _w26332_ ;
	wire _w26331_ ;
	wire _w26330_ ;
	wire _w26329_ ;
	wire _w26328_ ;
	wire _w26327_ ;
	wire _w26326_ ;
	wire _w26325_ ;
	wire _w26324_ ;
	wire _w26323_ ;
	wire _w26322_ ;
	wire _w26321_ ;
	wire _w26320_ ;
	wire _w26319_ ;
	wire _w26318_ ;
	wire _w26317_ ;
	wire _w26316_ ;
	wire _w26315_ ;
	wire _w26314_ ;
	wire _w26313_ ;
	wire _w26312_ ;
	wire _w26311_ ;
	wire _w26310_ ;
	wire _w26309_ ;
	wire _w26308_ ;
	wire _w26307_ ;
	wire _w26306_ ;
	wire _w26305_ ;
	wire _w26304_ ;
	wire _w26303_ ;
	wire _w26302_ ;
	wire _w26301_ ;
	wire _w26300_ ;
	wire _w26299_ ;
	wire _w26298_ ;
	wire _w26297_ ;
	wire _w26296_ ;
	wire _w26295_ ;
	wire _w26294_ ;
	wire _w26293_ ;
	wire _w26292_ ;
	wire _w26291_ ;
	wire _w26290_ ;
	wire _w26289_ ;
	wire _w26288_ ;
	wire _w26287_ ;
	wire _w26286_ ;
	wire _w26285_ ;
	wire _w26284_ ;
	wire _w26283_ ;
	wire _w26282_ ;
	wire _w26281_ ;
	wire _w26280_ ;
	wire _w26279_ ;
	wire _w26278_ ;
	wire _w26277_ ;
	wire _w26276_ ;
	wire _w26275_ ;
	wire _w26274_ ;
	wire _w26273_ ;
	wire _w26272_ ;
	wire _w26271_ ;
	wire _w26270_ ;
	wire _w26269_ ;
	wire _w26268_ ;
	wire _w26267_ ;
	wire _w26266_ ;
	wire _w26265_ ;
	wire _w26264_ ;
	wire _w26263_ ;
	wire _w26262_ ;
	wire _w26261_ ;
	wire _w26260_ ;
	wire _w26259_ ;
	wire _w26258_ ;
	wire _w26257_ ;
	wire _w26256_ ;
	wire _w26255_ ;
	wire _w26254_ ;
	wire _w26253_ ;
	wire _w26252_ ;
	wire _w26251_ ;
	wire _w26250_ ;
	wire _w26249_ ;
	wire _w26248_ ;
	wire _w26247_ ;
	wire _w26246_ ;
	wire _w26245_ ;
	wire _w26244_ ;
	wire _w26243_ ;
	wire _w26242_ ;
	wire _w26241_ ;
	wire _w26240_ ;
	wire _w26239_ ;
	wire _w26238_ ;
	wire _w26237_ ;
	wire _w26236_ ;
	wire _w26235_ ;
	wire _w26234_ ;
	wire _w26233_ ;
	wire _w26232_ ;
	wire _w26231_ ;
	wire _w26230_ ;
	wire _w26229_ ;
	wire _w26228_ ;
	wire _w26227_ ;
	wire _w26226_ ;
	wire _w26225_ ;
	wire _w26224_ ;
	wire _w26223_ ;
	wire _w26222_ ;
	wire _w26221_ ;
	wire _w26220_ ;
	wire _w26219_ ;
	wire _w26218_ ;
	wire _w26217_ ;
	wire _w26216_ ;
	wire _w26215_ ;
	wire _w26214_ ;
	wire _w26213_ ;
	wire _w26212_ ;
	wire _w26211_ ;
	wire _w26210_ ;
	wire _w26209_ ;
	wire _w26208_ ;
	wire _w26207_ ;
	wire _w26206_ ;
	wire _w26205_ ;
	wire _w26204_ ;
	wire _w26203_ ;
	wire _w26202_ ;
	wire _w26201_ ;
	wire _w26200_ ;
	wire _w26199_ ;
	wire _w26198_ ;
	wire _w26197_ ;
	wire _w26196_ ;
	wire _w26195_ ;
	wire _w26194_ ;
	wire _w26193_ ;
	wire _w26192_ ;
	wire _w26191_ ;
	wire _w26190_ ;
	wire _w26189_ ;
	wire _w26188_ ;
	wire _w26187_ ;
	wire _w26186_ ;
	wire _w26185_ ;
	wire _w26184_ ;
	wire _w26183_ ;
	wire _w26182_ ;
	wire _w26181_ ;
	wire _w26180_ ;
	wire _w26179_ ;
	wire _w26178_ ;
	wire _w26177_ ;
	wire _w26176_ ;
	wire _w26175_ ;
	wire _w26174_ ;
	wire _w26173_ ;
	wire _w26172_ ;
	wire _w26171_ ;
	wire _w26170_ ;
	wire _w26169_ ;
	wire _w26168_ ;
	wire _w26167_ ;
	wire _w26166_ ;
	wire _w26165_ ;
	wire _w26164_ ;
	wire _w26163_ ;
	wire _w26162_ ;
	wire _w26161_ ;
	wire _w26160_ ;
	wire _w26159_ ;
	wire _w26158_ ;
	wire _w26157_ ;
	wire _w26156_ ;
	wire _w26155_ ;
	wire _w26154_ ;
	wire _w26153_ ;
	wire _w26152_ ;
	wire _w26151_ ;
	wire _w26150_ ;
	wire _w26149_ ;
	wire _w26148_ ;
	wire _w26147_ ;
	wire _w26146_ ;
	wire _w26145_ ;
	wire _w26144_ ;
	wire _w26143_ ;
	wire _w26142_ ;
	wire _w26141_ ;
	wire _w26140_ ;
	wire _w26139_ ;
	wire _w26138_ ;
	wire _w26137_ ;
	wire _w26136_ ;
	wire _w26135_ ;
	wire _w26134_ ;
	wire _w26133_ ;
	wire _w26132_ ;
	wire _w26131_ ;
	wire _w26130_ ;
	wire _w26129_ ;
	wire _w26128_ ;
	wire _w26127_ ;
	wire _w26126_ ;
	wire _w26125_ ;
	wire _w26124_ ;
	wire _w26123_ ;
	wire _w26122_ ;
	wire _w26121_ ;
	wire _w26120_ ;
	wire _w26119_ ;
	wire _w26118_ ;
	wire _w26117_ ;
	wire _w26116_ ;
	wire _w26115_ ;
	wire _w26114_ ;
	wire _w26113_ ;
	wire _w26112_ ;
	wire _w26111_ ;
	wire _w26110_ ;
	wire _w26109_ ;
	wire _w26108_ ;
	wire _w26107_ ;
	wire _w26106_ ;
	wire _w26105_ ;
	wire _w26104_ ;
	wire _w26103_ ;
	wire _w26102_ ;
	wire _w26101_ ;
	wire _w26100_ ;
	wire _w26099_ ;
	wire _w26098_ ;
	wire _w26097_ ;
	wire _w26096_ ;
	wire _w26095_ ;
	wire _w26094_ ;
	wire _w26093_ ;
	wire _w26092_ ;
	wire _w26091_ ;
	wire _w26090_ ;
	wire _w26089_ ;
	wire _w26088_ ;
	wire _w26087_ ;
	wire _w26086_ ;
	wire _w26085_ ;
	wire _w26084_ ;
	wire _w26083_ ;
	wire _w26082_ ;
	wire _w26081_ ;
	wire _w26080_ ;
	wire _w26079_ ;
	wire _w26078_ ;
	wire _w26077_ ;
	wire _w26076_ ;
	wire _w26075_ ;
	wire _w26074_ ;
	wire _w26073_ ;
	wire _w26072_ ;
	wire _w26071_ ;
	wire _w26070_ ;
	wire _w26069_ ;
	wire _w26068_ ;
	wire _w26067_ ;
	wire _w26066_ ;
	wire _w26065_ ;
	wire _w26064_ ;
	wire _w26063_ ;
	wire _w26062_ ;
	wire _w26061_ ;
	wire _w26060_ ;
	wire _w26059_ ;
	wire _w26058_ ;
	wire _w26057_ ;
	wire _w26056_ ;
	wire _w26055_ ;
	wire _w26054_ ;
	wire _w26053_ ;
	wire _w26052_ ;
	wire _w26051_ ;
	wire _w26050_ ;
	wire _w26049_ ;
	wire _w26048_ ;
	wire _w26047_ ;
	wire _w26046_ ;
	wire _w26045_ ;
	wire _w26044_ ;
	wire _w26043_ ;
	wire _w26042_ ;
	wire _w26041_ ;
	wire _w26040_ ;
	wire _w26039_ ;
	wire _w26038_ ;
	wire _w26037_ ;
	wire _w26036_ ;
	wire _w26035_ ;
	wire _w26034_ ;
	wire _w26033_ ;
	wire _w26032_ ;
	wire _w26031_ ;
	wire _w26030_ ;
	wire _w26029_ ;
	wire _w26028_ ;
	wire _w26027_ ;
	wire _w26026_ ;
	wire _w26025_ ;
	wire _w26024_ ;
	wire _w26023_ ;
	wire _w26022_ ;
	wire _w26021_ ;
	wire _w26020_ ;
	wire _w26019_ ;
	wire _w26018_ ;
	wire _w26017_ ;
	wire _w26016_ ;
	wire _w26015_ ;
	wire _w26014_ ;
	wire _w26013_ ;
	wire _w26012_ ;
	wire _w26011_ ;
	wire _w26010_ ;
	wire _w26009_ ;
	wire _w26008_ ;
	wire _w26007_ ;
	wire _w26006_ ;
	wire _w26005_ ;
	wire _w26004_ ;
	wire _w26003_ ;
	wire _w26002_ ;
	wire _w26001_ ;
	wire _w26000_ ;
	wire _w25999_ ;
	wire _w25998_ ;
	wire _w25997_ ;
	wire _w25996_ ;
	wire _w25995_ ;
	wire _w25994_ ;
	wire _w25993_ ;
	wire _w25992_ ;
	wire _w25991_ ;
	wire _w25990_ ;
	wire _w25989_ ;
	wire _w25988_ ;
	wire _w25987_ ;
	wire _w25986_ ;
	wire _w25985_ ;
	wire _w25984_ ;
	wire _w25983_ ;
	wire _w25982_ ;
	wire _w25981_ ;
	wire _w25980_ ;
	wire _w25979_ ;
	wire _w25978_ ;
	wire _w25977_ ;
	wire _w25976_ ;
	wire _w25975_ ;
	wire _w25974_ ;
	wire _w25973_ ;
	wire _w25972_ ;
	wire _w25971_ ;
	wire _w25970_ ;
	wire _w25969_ ;
	wire _w25968_ ;
	wire _w25967_ ;
	wire _w25966_ ;
	wire _w25965_ ;
	wire _w25964_ ;
	wire _w25963_ ;
	wire _w25962_ ;
	wire _w25961_ ;
	wire _w25960_ ;
	wire _w25959_ ;
	wire _w25958_ ;
	wire _w25957_ ;
	wire _w25956_ ;
	wire _w25955_ ;
	wire _w25954_ ;
	wire _w25953_ ;
	wire _w25952_ ;
	wire _w25951_ ;
	wire _w25950_ ;
	wire _w25949_ ;
	wire _w25948_ ;
	wire _w25947_ ;
	wire _w25946_ ;
	wire _w25945_ ;
	wire _w25944_ ;
	wire _w25943_ ;
	wire _w25942_ ;
	wire _w25941_ ;
	wire _w25940_ ;
	wire _w25939_ ;
	wire _w25938_ ;
	wire _w25937_ ;
	wire _w25936_ ;
	wire _w25935_ ;
	wire _w25934_ ;
	wire _w25933_ ;
	wire _w25932_ ;
	wire _w25931_ ;
	wire _w25930_ ;
	wire _w25929_ ;
	wire _w25928_ ;
	wire _w25927_ ;
	wire _w25926_ ;
	wire _w25925_ ;
	wire _w25924_ ;
	wire _w25923_ ;
	wire _w25922_ ;
	wire _w25921_ ;
	wire _w25920_ ;
	wire _w25919_ ;
	wire _w25918_ ;
	wire _w25917_ ;
	wire _w25916_ ;
	wire _w25915_ ;
	wire _w25914_ ;
	wire _w25913_ ;
	wire _w25912_ ;
	wire _w25911_ ;
	wire _w25910_ ;
	wire _w25909_ ;
	wire _w25908_ ;
	wire _w25907_ ;
	wire _w25906_ ;
	wire _w25905_ ;
	wire _w25904_ ;
	wire _w25903_ ;
	wire _w25902_ ;
	wire _w25901_ ;
	wire _w25900_ ;
	wire _w25899_ ;
	wire _w25898_ ;
	wire _w25897_ ;
	wire _w25896_ ;
	wire _w25895_ ;
	wire _w25894_ ;
	wire _w25893_ ;
	wire _w25892_ ;
	wire _w25891_ ;
	wire _w25890_ ;
	wire _w25889_ ;
	wire _w25888_ ;
	wire _w25887_ ;
	wire _w25886_ ;
	wire _w25885_ ;
	wire _w25884_ ;
	wire _w25883_ ;
	wire _w25882_ ;
	wire _w25881_ ;
	wire _w25880_ ;
	wire _w25879_ ;
	wire _w25878_ ;
	wire _w25877_ ;
	wire _w25876_ ;
	wire _w25875_ ;
	wire _w25874_ ;
	wire _w25873_ ;
	wire _w25872_ ;
	wire _w25871_ ;
	wire _w25870_ ;
	wire _w25869_ ;
	wire _w25868_ ;
	wire _w25867_ ;
	wire _w25866_ ;
	wire _w25865_ ;
	wire _w25864_ ;
	wire _w25863_ ;
	wire _w25862_ ;
	wire _w25861_ ;
	wire _w25860_ ;
	wire _w25859_ ;
	wire _w25858_ ;
	wire _w25857_ ;
	wire _w25856_ ;
	wire _w25855_ ;
	wire _w25854_ ;
	wire _w25853_ ;
	wire _w25852_ ;
	wire _w25851_ ;
	wire _w25850_ ;
	wire _w25849_ ;
	wire _w25848_ ;
	wire _w25847_ ;
	wire _w25846_ ;
	wire _w25845_ ;
	wire _w25844_ ;
	wire _w25843_ ;
	wire _w25842_ ;
	wire _w25841_ ;
	wire _w25840_ ;
	wire _w25839_ ;
	wire _w25838_ ;
	wire _w25837_ ;
	wire _w25836_ ;
	wire _w25835_ ;
	wire _w25834_ ;
	wire _w25833_ ;
	wire _w25832_ ;
	wire _w25831_ ;
	wire _w25830_ ;
	wire _w25829_ ;
	wire _w25828_ ;
	wire _w25827_ ;
	wire _w25826_ ;
	wire _w25825_ ;
	wire _w25824_ ;
	wire _w25823_ ;
	wire _w25822_ ;
	wire _w25821_ ;
	wire _w25820_ ;
	wire _w25819_ ;
	wire _w25818_ ;
	wire _w25817_ ;
	wire _w25816_ ;
	wire _w25815_ ;
	wire _w25814_ ;
	wire _w25813_ ;
	wire _w25812_ ;
	wire _w25811_ ;
	wire _w25810_ ;
	wire _w25809_ ;
	wire _w25808_ ;
	wire _w25807_ ;
	wire _w25806_ ;
	wire _w25805_ ;
	wire _w25804_ ;
	wire _w25803_ ;
	wire _w25802_ ;
	wire _w25801_ ;
	wire _w25800_ ;
	wire _w25799_ ;
	wire _w25798_ ;
	wire _w25797_ ;
	wire _w25796_ ;
	wire _w25795_ ;
	wire _w25794_ ;
	wire _w25793_ ;
	wire _w25792_ ;
	wire _w25791_ ;
	wire _w25790_ ;
	wire _w25789_ ;
	wire _w25788_ ;
	wire _w25787_ ;
	wire _w25786_ ;
	wire _w25785_ ;
	wire _w25784_ ;
	wire _w25783_ ;
	wire _w25782_ ;
	wire _w25781_ ;
	wire _w25780_ ;
	wire _w25779_ ;
	wire _w25778_ ;
	wire _w25777_ ;
	wire _w25776_ ;
	wire _w25775_ ;
	wire _w25774_ ;
	wire _w25773_ ;
	wire _w25772_ ;
	wire _w25771_ ;
	wire _w25770_ ;
	wire _w25769_ ;
	wire _w25768_ ;
	wire _w25767_ ;
	wire _w25766_ ;
	wire _w25765_ ;
	wire _w25764_ ;
	wire _w25763_ ;
	wire _w25762_ ;
	wire _w25761_ ;
	wire _w25760_ ;
	wire _w25759_ ;
	wire _w25758_ ;
	wire _w25757_ ;
	wire _w25756_ ;
	wire _w25755_ ;
	wire _w25754_ ;
	wire _w25753_ ;
	wire _w25752_ ;
	wire _w25751_ ;
	wire _w25750_ ;
	wire _w25749_ ;
	wire _w25748_ ;
	wire _w25747_ ;
	wire _w25746_ ;
	wire _w25745_ ;
	wire _w25744_ ;
	wire _w25743_ ;
	wire _w25742_ ;
	wire _w25741_ ;
	wire _w25740_ ;
	wire _w25739_ ;
	wire _w25738_ ;
	wire _w25737_ ;
	wire _w25736_ ;
	wire _w25735_ ;
	wire _w25734_ ;
	wire _w25733_ ;
	wire _w25732_ ;
	wire _w25731_ ;
	wire _w25730_ ;
	wire _w25729_ ;
	wire _w25728_ ;
	wire _w25727_ ;
	wire _w25726_ ;
	wire _w25725_ ;
	wire _w25724_ ;
	wire _w25723_ ;
	wire _w25722_ ;
	wire _w25721_ ;
	wire _w25720_ ;
	wire _w25719_ ;
	wire _w25718_ ;
	wire _w25717_ ;
	wire _w25716_ ;
	wire _w25715_ ;
	wire _w25714_ ;
	wire _w25713_ ;
	wire _w25712_ ;
	wire _w25711_ ;
	wire _w25710_ ;
	wire _w25709_ ;
	wire _w25708_ ;
	wire _w25707_ ;
	wire _w25706_ ;
	wire _w25705_ ;
	wire _w25704_ ;
	wire _w25703_ ;
	wire _w25702_ ;
	wire _w25701_ ;
	wire _w25700_ ;
	wire _w25699_ ;
	wire _w25698_ ;
	wire _w25697_ ;
	wire _w25696_ ;
	wire _w25695_ ;
	wire _w25694_ ;
	wire _w25693_ ;
	wire _w25692_ ;
	wire _w25691_ ;
	wire _w25690_ ;
	wire _w25689_ ;
	wire _w25688_ ;
	wire _w25687_ ;
	wire _w25686_ ;
	wire _w25685_ ;
	wire _w25684_ ;
	wire _w25683_ ;
	wire _w25682_ ;
	wire _w25681_ ;
	wire _w25680_ ;
	wire _w25679_ ;
	wire _w25678_ ;
	wire _w25677_ ;
	wire _w25676_ ;
	wire _w25675_ ;
	wire _w25674_ ;
	wire _w25673_ ;
	wire _w25672_ ;
	wire _w25671_ ;
	wire _w25670_ ;
	wire _w25669_ ;
	wire _w25668_ ;
	wire _w25667_ ;
	wire _w25666_ ;
	wire _w25665_ ;
	wire _w25664_ ;
	wire _w25663_ ;
	wire _w25662_ ;
	wire _w25661_ ;
	wire _w25660_ ;
	wire _w25659_ ;
	wire _w25658_ ;
	wire _w25657_ ;
	wire _w25656_ ;
	wire _w25655_ ;
	wire _w25654_ ;
	wire _w25653_ ;
	wire _w25652_ ;
	wire _w25651_ ;
	wire _w25650_ ;
	wire _w25649_ ;
	wire _w25648_ ;
	wire _w25647_ ;
	wire _w25646_ ;
	wire _w25645_ ;
	wire _w25644_ ;
	wire _w25643_ ;
	wire _w25642_ ;
	wire _w25641_ ;
	wire _w25640_ ;
	wire _w25639_ ;
	wire _w25638_ ;
	wire _w25637_ ;
	wire _w25636_ ;
	wire _w25635_ ;
	wire _w25634_ ;
	wire _w25633_ ;
	wire _w25632_ ;
	wire _w25631_ ;
	wire _w25630_ ;
	wire _w25629_ ;
	wire _w25628_ ;
	wire _w25627_ ;
	wire _w25626_ ;
	wire _w25625_ ;
	wire _w25624_ ;
	wire _w25623_ ;
	wire _w25622_ ;
	wire _w25621_ ;
	wire _w25620_ ;
	wire _w25619_ ;
	wire _w25618_ ;
	wire _w25617_ ;
	wire _w25616_ ;
	wire _w25615_ ;
	wire _w25614_ ;
	wire _w25613_ ;
	wire _w25612_ ;
	wire _w25611_ ;
	wire _w25610_ ;
	wire _w25609_ ;
	wire _w25608_ ;
	wire _w25607_ ;
	wire _w25606_ ;
	wire _w25605_ ;
	wire _w25604_ ;
	wire _w25603_ ;
	wire _w25602_ ;
	wire _w25601_ ;
	wire _w25600_ ;
	wire _w25599_ ;
	wire _w25598_ ;
	wire _w25597_ ;
	wire _w25596_ ;
	wire _w25595_ ;
	wire _w25594_ ;
	wire _w25593_ ;
	wire _w25592_ ;
	wire _w25591_ ;
	wire _w25590_ ;
	wire _w25589_ ;
	wire _w25588_ ;
	wire _w25587_ ;
	wire _w25586_ ;
	wire _w25585_ ;
	wire _w25584_ ;
	wire _w25583_ ;
	wire _w25582_ ;
	wire _w25581_ ;
	wire _w25580_ ;
	wire _w25579_ ;
	wire _w25578_ ;
	wire _w25577_ ;
	wire _w25576_ ;
	wire _w25575_ ;
	wire _w25574_ ;
	wire _w25573_ ;
	wire _w25572_ ;
	wire _w25571_ ;
	wire _w25570_ ;
	wire _w25569_ ;
	wire _w25568_ ;
	wire _w25567_ ;
	wire _w25566_ ;
	wire _w25565_ ;
	wire _w25564_ ;
	wire _w25563_ ;
	wire _w25562_ ;
	wire _w25561_ ;
	wire _w25560_ ;
	wire _w25559_ ;
	wire _w25558_ ;
	wire _w25557_ ;
	wire _w25556_ ;
	wire _w25555_ ;
	wire _w25554_ ;
	wire _w25553_ ;
	wire _w25552_ ;
	wire _w25551_ ;
	wire _w25550_ ;
	wire _w25549_ ;
	wire _w25548_ ;
	wire _w25547_ ;
	wire _w25546_ ;
	wire _w25545_ ;
	wire _w25544_ ;
	wire _w25543_ ;
	wire _w25542_ ;
	wire _w25541_ ;
	wire _w25540_ ;
	wire _w25539_ ;
	wire _w25538_ ;
	wire _w25537_ ;
	wire _w25536_ ;
	wire _w25535_ ;
	wire _w25534_ ;
	wire _w25533_ ;
	wire _w25532_ ;
	wire _w25531_ ;
	wire _w25530_ ;
	wire _w25529_ ;
	wire _w25528_ ;
	wire _w25527_ ;
	wire _w25526_ ;
	wire _w25525_ ;
	wire _w25524_ ;
	wire _w25523_ ;
	wire _w25522_ ;
	wire _w25521_ ;
	wire _w25520_ ;
	wire _w25519_ ;
	wire _w25518_ ;
	wire _w25517_ ;
	wire _w25516_ ;
	wire _w25515_ ;
	wire _w25514_ ;
	wire _w25513_ ;
	wire _w25512_ ;
	wire _w25511_ ;
	wire _w25510_ ;
	wire _w25509_ ;
	wire _w25508_ ;
	wire _w25507_ ;
	wire _w25506_ ;
	wire _w25505_ ;
	wire _w25504_ ;
	wire _w25503_ ;
	wire _w25502_ ;
	wire _w25501_ ;
	wire _w25500_ ;
	wire _w25499_ ;
	wire _w25498_ ;
	wire _w25497_ ;
	wire _w25496_ ;
	wire _w25495_ ;
	wire _w25494_ ;
	wire _w25493_ ;
	wire _w25492_ ;
	wire _w25491_ ;
	wire _w25490_ ;
	wire _w25489_ ;
	wire _w25488_ ;
	wire _w25487_ ;
	wire _w25486_ ;
	wire _w25485_ ;
	wire _w25484_ ;
	wire _w25483_ ;
	wire _w25482_ ;
	wire _w25481_ ;
	wire _w25480_ ;
	wire _w25479_ ;
	wire _w25478_ ;
	wire _w25477_ ;
	wire _w25476_ ;
	wire _w25475_ ;
	wire _w25474_ ;
	wire _w25473_ ;
	wire _w25472_ ;
	wire _w25471_ ;
	wire _w25470_ ;
	wire _w25469_ ;
	wire _w25468_ ;
	wire _w25467_ ;
	wire _w25466_ ;
	wire _w25465_ ;
	wire _w25464_ ;
	wire _w25463_ ;
	wire _w25462_ ;
	wire _w25461_ ;
	wire _w25460_ ;
	wire _w25459_ ;
	wire _w25458_ ;
	wire _w25457_ ;
	wire _w25456_ ;
	wire _w25455_ ;
	wire _w25454_ ;
	wire _w25453_ ;
	wire _w25452_ ;
	wire _w25451_ ;
	wire _w25450_ ;
	wire _w25449_ ;
	wire _w25448_ ;
	wire _w25447_ ;
	wire _w25446_ ;
	wire _w25445_ ;
	wire _w25444_ ;
	wire _w25443_ ;
	wire _w25442_ ;
	wire _w25441_ ;
	wire _w25440_ ;
	wire _w25439_ ;
	wire _w25438_ ;
	wire _w25437_ ;
	wire _w25436_ ;
	wire _w25435_ ;
	wire _w25434_ ;
	wire _w25433_ ;
	wire _w25432_ ;
	wire _w25431_ ;
	wire _w25430_ ;
	wire _w25429_ ;
	wire _w25428_ ;
	wire _w25427_ ;
	wire _w25426_ ;
	wire _w25425_ ;
	wire _w25424_ ;
	wire _w25423_ ;
	wire _w25422_ ;
	wire _w25421_ ;
	wire _w25420_ ;
	wire _w25419_ ;
	wire _w25418_ ;
	wire _w25417_ ;
	wire _w25416_ ;
	wire _w25415_ ;
	wire _w25414_ ;
	wire _w25413_ ;
	wire _w25412_ ;
	wire _w25411_ ;
	wire _w25410_ ;
	wire _w25409_ ;
	wire _w25408_ ;
	wire _w25407_ ;
	wire _w25406_ ;
	wire _w25405_ ;
	wire _w25404_ ;
	wire _w25403_ ;
	wire _w25402_ ;
	wire _w25401_ ;
	wire _w25400_ ;
	wire _w25399_ ;
	wire _w25398_ ;
	wire _w25397_ ;
	wire _w25396_ ;
	wire _w25395_ ;
	wire _w25394_ ;
	wire _w25393_ ;
	wire _w25392_ ;
	wire _w25391_ ;
	wire _w25390_ ;
	wire _w25389_ ;
	wire _w25388_ ;
	wire _w25387_ ;
	wire _w25386_ ;
	wire _w25385_ ;
	wire _w25384_ ;
	wire _w25383_ ;
	wire _w25382_ ;
	wire _w25381_ ;
	wire _w25380_ ;
	wire _w25379_ ;
	wire _w25378_ ;
	wire _w25377_ ;
	wire _w25376_ ;
	wire _w25375_ ;
	wire _w25374_ ;
	wire _w25373_ ;
	wire _w25372_ ;
	wire _w25371_ ;
	wire _w25370_ ;
	wire _w25369_ ;
	wire _w25368_ ;
	wire _w25367_ ;
	wire _w25366_ ;
	wire _w25365_ ;
	wire _w25364_ ;
	wire _w25363_ ;
	wire _w25362_ ;
	wire _w25361_ ;
	wire _w25360_ ;
	wire _w25359_ ;
	wire _w25358_ ;
	wire _w25357_ ;
	wire _w25356_ ;
	wire _w25355_ ;
	wire _w25354_ ;
	wire _w25353_ ;
	wire _w25352_ ;
	wire _w25351_ ;
	wire _w25350_ ;
	wire _w25349_ ;
	wire _w25348_ ;
	wire _w25347_ ;
	wire _w25346_ ;
	wire _w25345_ ;
	wire _w25344_ ;
	wire _w25343_ ;
	wire _w25342_ ;
	wire _w25341_ ;
	wire _w25340_ ;
	wire _w25339_ ;
	wire _w25338_ ;
	wire _w25337_ ;
	wire _w25336_ ;
	wire _w25335_ ;
	wire _w25334_ ;
	wire _w25333_ ;
	wire _w25332_ ;
	wire _w25331_ ;
	wire _w25330_ ;
	wire _w25329_ ;
	wire _w25328_ ;
	wire _w25327_ ;
	wire _w25326_ ;
	wire _w25325_ ;
	wire _w25324_ ;
	wire _w25323_ ;
	wire _w25322_ ;
	wire _w25321_ ;
	wire _w25320_ ;
	wire _w25319_ ;
	wire _w25318_ ;
	wire _w25317_ ;
	wire _w25316_ ;
	wire _w25315_ ;
	wire _w25314_ ;
	wire _w25313_ ;
	wire _w25312_ ;
	wire _w25311_ ;
	wire _w25310_ ;
	wire _w25309_ ;
	wire _w25308_ ;
	wire _w25307_ ;
	wire _w25306_ ;
	wire _w25305_ ;
	wire _w25304_ ;
	wire _w25303_ ;
	wire _w25302_ ;
	wire _w25301_ ;
	wire _w25300_ ;
	wire _w25299_ ;
	wire _w25298_ ;
	wire _w25297_ ;
	wire _w25296_ ;
	wire _w25295_ ;
	wire _w25294_ ;
	wire _w25293_ ;
	wire _w25292_ ;
	wire _w25291_ ;
	wire _w25290_ ;
	wire _w25289_ ;
	wire _w25288_ ;
	wire _w25287_ ;
	wire _w25286_ ;
	wire _w25285_ ;
	wire _w25284_ ;
	wire _w25283_ ;
	wire _w25282_ ;
	wire _w25281_ ;
	wire _w25280_ ;
	wire _w25279_ ;
	wire _w25278_ ;
	wire _w25277_ ;
	wire _w25276_ ;
	wire _w25275_ ;
	wire _w25274_ ;
	wire _w25273_ ;
	wire _w25272_ ;
	wire _w25271_ ;
	wire _w25270_ ;
	wire _w25269_ ;
	wire _w25268_ ;
	wire _w25267_ ;
	wire _w25266_ ;
	wire _w25265_ ;
	wire _w25264_ ;
	wire _w25263_ ;
	wire _w25262_ ;
	wire _w25261_ ;
	wire _w25260_ ;
	wire _w25259_ ;
	wire _w25258_ ;
	wire _w25257_ ;
	wire _w25256_ ;
	wire _w25255_ ;
	wire _w25254_ ;
	wire _w25253_ ;
	wire _w25252_ ;
	wire _w25251_ ;
	wire _w25250_ ;
	wire _w25249_ ;
	wire _w25248_ ;
	wire _w25247_ ;
	wire _w25246_ ;
	wire _w25245_ ;
	wire _w25244_ ;
	wire _w25243_ ;
	wire _w25242_ ;
	wire _w25241_ ;
	wire _w25240_ ;
	wire _w25239_ ;
	wire _w25238_ ;
	wire _w25237_ ;
	wire _w25236_ ;
	wire _w25235_ ;
	wire _w25234_ ;
	wire _w25233_ ;
	wire _w25232_ ;
	wire _w25231_ ;
	wire _w25230_ ;
	wire _w25229_ ;
	wire _w25228_ ;
	wire _w25227_ ;
	wire _w25226_ ;
	wire _w25225_ ;
	wire _w25224_ ;
	wire _w25223_ ;
	wire _w25222_ ;
	wire _w25221_ ;
	wire _w25220_ ;
	wire _w25219_ ;
	wire _w25218_ ;
	wire _w25217_ ;
	wire _w25216_ ;
	wire _w25215_ ;
	wire _w25214_ ;
	wire _w25213_ ;
	wire _w25212_ ;
	wire _w25211_ ;
	wire _w25210_ ;
	wire _w25209_ ;
	wire _w25208_ ;
	wire _w25207_ ;
	wire _w25206_ ;
	wire _w25205_ ;
	wire _w25204_ ;
	wire _w25203_ ;
	wire _w25202_ ;
	wire _w25201_ ;
	wire _w25200_ ;
	wire _w25199_ ;
	wire _w25198_ ;
	wire _w25197_ ;
	wire _w25196_ ;
	wire _w25195_ ;
	wire _w25194_ ;
	wire _w25193_ ;
	wire _w25192_ ;
	wire _w25191_ ;
	wire _w25190_ ;
	wire _w25189_ ;
	wire _w25188_ ;
	wire _w25187_ ;
	wire _w25186_ ;
	wire _w25185_ ;
	wire _w25184_ ;
	wire _w25183_ ;
	wire _w25182_ ;
	wire _w25181_ ;
	wire _w25180_ ;
	wire _w25179_ ;
	wire _w25178_ ;
	wire _w25177_ ;
	wire _w25176_ ;
	wire _w25175_ ;
	wire _w25174_ ;
	wire _w25173_ ;
	wire _w25172_ ;
	wire _w25171_ ;
	wire _w25170_ ;
	wire _w25169_ ;
	wire _w25168_ ;
	wire _w25167_ ;
	wire _w25166_ ;
	wire _w25165_ ;
	wire _w25164_ ;
	wire _w25163_ ;
	wire _w25162_ ;
	wire _w25161_ ;
	wire _w25160_ ;
	wire _w25159_ ;
	wire _w25158_ ;
	wire _w25157_ ;
	wire _w25156_ ;
	wire _w25155_ ;
	wire _w25154_ ;
	wire _w25153_ ;
	wire _w25152_ ;
	wire _w25151_ ;
	wire _w25150_ ;
	wire _w25149_ ;
	wire _w25148_ ;
	wire _w25147_ ;
	wire _w25146_ ;
	wire _w25145_ ;
	wire _w25144_ ;
	wire _w25143_ ;
	wire _w25142_ ;
	wire _w25141_ ;
	wire _w25140_ ;
	wire _w25139_ ;
	wire _w25138_ ;
	wire _w25137_ ;
	wire _w25136_ ;
	wire _w25135_ ;
	wire _w25134_ ;
	wire _w25133_ ;
	wire _w25132_ ;
	wire _w25131_ ;
	wire _w25130_ ;
	wire _w25129_ ;
	wire _w25128_ ;
	wire _w25127_ ;
	wire _w25126_ ;
	wire _w25125_ ;
	wire _w25124_ ;
	wire _w25123_ ;
	wire _w25122_ ;
	wire _w25121_ ;
	wire _w25120_ ;
	wire _w25119_ ;
	wire _w25118_ ;
	wire _w25117_ ;
	wire _w25116_ ;
	wire _w25115_ ;
	wire _w25114_ ;
	wire _w25113_ ;
	wire _w25112_ ;
	wire _w25111_ ;
	wire _w25110_ ;
	wire _w25109_ ;
	wire _w25108_ ;
	wire _w25107_ ;
	wire _w25106_ ;
	wire _w25105_ ;
	wire _w25104_ ;
	wire _w25103_ ;
	wire _w25102_ ;
	wire _w25101_ ;
	wire _w25100_ ;
	wire _w25099_ ;
	wire _w25098_ ;
	wire _w25097_ ;
	wire _w25096_ ;
	wire _w25095_ ;
	wire _w25094_ ;
	wire _w25093_ ;
	wire _w25092_ ;
	wire _w25091_ ;
	wire _w25090_ ;
	wire _w25089_ ;
	wire _w25088_ ;
	wire _w25087_ ;
	wire _w25086_ ;
	wire _w25085_ ;
	wire _w25084_ ;
	wire _w25083_ ;
	wire _w25082_ ;
	wire _w25081_ ;
	wire _w25080_ ;
	wire _w25079_ ;
	wire _w25078_ ;
	wire _w25077_ ;
	wire _w25076_ ;
	wire _w25075_ ;
	wire _w25074_ ;
	wire _w25073_ ;
	wire _w25072_ ;
	wire _w25071_ ;
	wire _w25070_ ;
	wire _w25069_ ;
	wire _w25068_ ;
	wire _w25067_ ;
	wire _w25066_ ;
	wire _w25065_ ;
	wire _w25064_ ;
	wire _w25063_ ;
	wire _w25062_ ;
	wire _w25061_ ;
	wire _w25060_ ;
	wire _w25059_ ;
	wire _w25058_ ;
	wire _w25057_ ;
	wire _w25056_ ;
	wire _w25055_ ;
	wire _w25054_ ;
	wire _w25053_ ;
	wire _w25052_ ;
	wire _w25051_ ;
	wire _w25050_ ;
	wire _w25049_ ;
	wire _w25048_ ;
	wire _w25047_ ;
	wire _w25046_ ;
	wire _w25045_ ;
	wire _w25044_ ;
	wire _w25043_ ;
	wire _w25042_ ;
	wire _w25041_ ;
	wire _w25040_ ;
	wire _w25039_ ;
	wire _w25038_ ;
	wire _w25037_ ;
	wire _w25036_ ;
	wire _w25035_ ;
	wire _w25034_ ;
	wire _w25033_ ;
	wire _w25032_ ;
	wire _w25031_ ;
	wire _w25030_ ;
	wire _w25029_ ;
	wire _w25028_ ;
	wire _w25027_ ;
	wire _w25026_ ;
	wire _w25025_ ;
	wire _w25024_ ;
	wire _w25023_ ;
	wire _w25022_ ;
	wire _w25021_ ;
	wire _w25020_ ;
	wire _w25019_ ;
	wire _w25018_ ;
	wire _w25017_ ;
	wire _w25016_ ;
	wire _w25015_ ;
	wire _w25014_ ;
	wire _w25013_ ;
	wire _w25012_ ;
	wire _w25011_ ;
	wire _w25010_ ;
	wire _w25009_ ;
	wire _w25008_ ;
	wire _w25007_ ;
	wire _w25006_ ;
	wire _w25005_ ;
	wire _w25004_ ;
	wire _w25003_ ;
	wire _w25002_ ;
	wire _w25001_ ;
	wire _w25000_ ;
	wire _w24999_ ;
	wire _w24998_ ;
	wire _w24997_ ;
	wire _w24996_ ;
	wire _w24995_ ;
	wire _w24994_ ;
	wire _w24993_ ;
	wire _w24992_ ;
	wire _w24991_ ;
	wire _w24990_ ;
	wire _w24989_ ;
	wire _w24988_ ;
	wire _w24987_ ;
	wire _w24986_ ;
	wire _w24985_ ;
	wire _w24984_ ;
	wire _w24983_ ;
	wire _w24982_ ;
	wire _w24981_ ;
	wire _w24980_ ;
	wire _w24979_ ;
	wire _w24978_ ;
	wire _w24977_ ;
	wire _w24976_ ;
	wire _w24975_ ;
	wire _w24974_ ;
	wire _w24973_ ;
	wire _w24972_ ;
	wire _w24971_ ;
	wire _w24970_ ;
	wire _w24969_ ;
	wire _w24968_ ;
	wire _w24967_ ;
	wire _w24966_ ;
	wire _w24965_ ;
	wire _w24964_ ;
	wire _w24963_ ;
	wire _w24962_ ;
	wire _w24961_ ;
	wire _w24960_ ;
	wire _w24959_ ;
	wire _w24958_ ;
	wire _w24957_ ;
	wire _w24956_ ;
	wire _w24955_ ;
	wire _w24954_ ;
	wire _w24953_ ;
	wire _w24952_ ;
	wire _w24951_ ;
	wire _w24950_ ;
	wire _w24949_ ;
	wire _w24948_ ;
	wire _w24947_ ;
	wire _w24946_ ;
	wire _w24945_ ;
	wire _w24944_ ;
	wire _w24943_ ;
	wire _w24942_ ;
	wire _w24941_ ;
	wire _w24940_ ;
	wire _w24939_ ;
	wire _w24938_ ;
	wire _w24937_ ;
	wire _w24936_ ;
	wire _w24935_ ;
	wire _w24934_ ;
	wire _w24933_ ;
	wire _w24932_ ;
	wire _w24931_ ;
	wire _w24930_ ;
	wire _w24929_ ;
	wire _w24928_ ;
	wire _w24927_ ;
	wire _w24926_ ;
	wire _w24925_ ;
	wire _w24924_ ;
	wire _w24923_ ;
	wire _w24922_ ;
	wire _w24921_ ;
	wire _w24920_ ;
	wire _w24919_ ;
	wire _w24918_ ;
	wire _w24917_ ;
	wire _w24916_ ;
	wire _w24915_ ;
	wire _w24914_ ;
	wire _w24913_ ;
	wire _w24912_ ;
	wire _w24911_ ;
	wire _w24910_ ;
	wire _w24909_ ;
	wire _w24908_ ;
	wire _w24907_ ;
	wire _w24906_ ;
	wire _w24905_ ;
	wire _w24904_ ;
	wire _w24903_ ;
	wire _w24902_ ;
	wire _w24901_ ;
	wire _w24900_ ;
	wire _w24899_ ;
	wire _w24898_ ;
	wire _w24897_ ;
	wire _w24896_ ;
	wire _w24895_ ;
	wire _w24894_ ;
	wire _w24893_ ;
	wire _w24892_ ;
	wire _w24891_ ;
	wire _w24890_ ;
	wire _w24889_ ;
	wire _w24888_ ;
	wire _w24887_ ;
	wire _w24886_ ;
	wire _w24885_ ;
	wire _w24884_ ;
	wire _w24883_ ;
	wire _w24882_ ;
	wire _w24881_ ;
	wire _w24880_ ;
	wire _w24879_ ;
	wire _w24878_ ;
	wire _w24877_ ;
	wire _w24876_ ;
	wire _w24875_ ;
	wire _w24874_ ;
	wire _w24873_ ;
	wire _w24872_ ;
	wire _w24871_ ;
	wire _w24870_ ;
	wire _w24869_ ;
	wire _w24868_ ;
	wire _w24867_ ;
	wire _w24866_ ;
	wire _w24865_ ;
	wire _w24864_ ;
	wire _w24863_ ;
	wire _w24862_ ;
	wire _w24861_ ;
	wire _w24860_ ;
	wire _w24859_ ;
	wire _w24858_ ;
	wire _w24857_ ;
	wire _w24856_ ;
	wire _w24855_ ;
	wire _w24854_ ;
	wire _w24853_ ;
	wire _w24852_ ;
	wire _w24851_ ;
	wire _w24850_ ;
	wire _w24849_ ;
	wire _w24848_ ;
	wire _w24847_ ;
	wire _w24846_ ;
	wire _w24845_ ;
	wire _w24844_ ;
	wire _w24843_ ;
	wire _w24842_ ;
	wire _w24841_ ;
	wire _w24840_ ;
	wire _w24839_ ;
	wire _w24838_ ;
	wire _w24837_ ;
	wire _w24836_ ;
	wire _w24835_ ;
	wire _w24834_ ;
	wire _w24833_ ;
	wire _w24832_ ;
	wire _w24831_ ;
	wire _w24830_ ;
	wire _w24829_ ;
	wire _w24828_ ;
	wire _w24827_ ;
	wire _w24826_ ;
	wire _w24825_ ;
	wire _w24824_ ;
	wire _w24823_ ;
	wire _w24822_ ;
	wire _w24821_ ;
	wire _w24820_ ;
	wire _w24819_ ;
	wire _w24818_ ;
	wire _w24817_ ;
	wire _w24816_ ;
	wire _w24815_ ;
	wire _w24814_ ;
	wire _w24813_ ;
	wire _w24812_ ;
	wire _w24811_ ;
	wire _w24810_ ;
	wire _w24809_ ;
	wire _w24808_ ;
	wire _w24807_ ;
	wire _w24806_ ;
	wire _w24805_ ;
	wire _w24804_ ;
	wire _w24803_ ;
	wire _w24802_ ;
	wire _w24801_ ;
	wire _w24800_ ;
	wire _w24799_ ;
	wire _w24798_ ;
	wire _w24797_ ;
	wire _w24796_ ;
	wire _w24795_ ;
	wire _w24794_ ;
	wire _w24793_ ;
	wire _w24792_ ;
	wire _w24791_ ;
	wire _w24790_ ;
	wire _w24789_ ;
	wire _w24788_ ;
	wire _w24787_ ;
	wire _w24786_ ;
	wire _w24785_ ;
	wire _w24784_ ;
	wire _w24783_ ;
	wire _w24782_ ;
	wire _w24781_ ;
	wire _w24780_ ;
	wire _w24779_ ;
	wire _w24778_ ;
	wire _w24777_ ;
	wire _w24776_ ;
	wire _w24775_ ;
	wire _w24774_ ;
	wire _w24773_ ;
	wire _w24772_ ;
	wire _w24771_ ;
	wire _w24770_ ;
	wire _w24769_ ;
	wire _w24768_ ;
	wire _w24767_ ;
	wire _w24766_ ;
	wire _w24765_ ;
	wire _w24764_ ;
	wire _w24763_ ;
	wire _w24762_ ;
	wire _w24761_ ;
	wire _w24760_ ;
	wire _w24759_ ;
	wire _w24758_ ;
	wire _w24757_ ;
	wire _w24756_ ;
	wire _w24755_ ;
	wire _w24754_ ;
	wire _w24753_ ;
	wire _w24752_ ;
	wire _w24751_ ;
	wire _w24750_ ;
	wire _w24749_ ;
	wire _w24748_ ;
	wire _w24747_ ;
	wire _w24746_ ;
	wire _w24745_ ;
	wire _w24744_ ;
	wire _w24743_ ;
	wire _w24742_ ;
	wire _w24741_ ;
	wire _w24740_ ;
	wire _w24739_ ;
	wire _w24738_ ;
	wire _w24737_ ;
	wire _w24736_ ;
	wire _w24735_ ;
	wire _w24734_ ;
	wire _w24733_ ;
	wire _w24732_ ;
	wire _w24731_ ;
	wire _w24730_ ;
	wire _w24729_ ;
	wire _w24728_ ;
	wire _w24727_ ;
	wire _w24726_ ;
	wire _w24725_ ;
	wire _w24724_ ;
	wire _w24723_ ;
	wire _w24722_ ;
	wire _w24721_ ;
	wire _w24720_ ;
	wire _w24719_ ;
	wire _w24718_ ;
	wire _w24717_ ;
	wire _w24716_ ;
	wire _w24715_ ;
	wire _w24714_ ;
	wire _w24713_ ;
	wire _w24712_ ;
	wire _w24711_ ;
	wire _w24710_ ;
	wire _w24709_ ;
	wire _w24708_ ;
	wire _w24707_ ;
	wire _w24706_ ;
	wire _w24705_ ;
	wire _w24704_ ;
	wire _w24703_ ;
	wire _w24702_ ;
	wire _w24701_ ;
	wire _w24700_ ;
	wire _w24699_ ;
	wire _w24698_ ;
	wire _w24697_ ;
	wire _w24696_ ;
	wire _w24695_ ;
	wire _w24694_ ;
	wire _w24693_ ;
	wire _w24692_ ;
	wire _w24691_ ;
	wire _w24690_ ;
	wire _w24689_ ;
	wire _w24688_ ;
	wire _w24687_ ;
	wire _w24686_ ;
	wire _w24685_ ;
	wire _w24684_ ;
	wire _w24683_ ;
	wire _w24682_ ;
	wire _w24681_ ;
	wire _w24680_ ;
	wire _w24679_ ;
	wire _w24678_ ;
	wire _w24677_ ;
	wire _w24676_ ;
	wire _w24675_ ;
	wire _w24674_ ;
	wire _w24673_ ;
	wire _w24672_ ;
	wire _w24671_ ;
	wire _w24670_ ;
	wire _w24669_ ;
	wire _w24668_ ;
	wire _w24667_ ;
	wire _w24666_ ;
	wire _w24665_ ;
	wire _w24664_ ;
	wire _w24663_ ;
	wire _w24662_ ;
	wire _w24661_ ;
	wire _w24660_ ;
	wire _w24659_ ;
	wire _w24658_ ;
	wire _w24657_ ;
	wire _w24656_ ;
	wire _w24655_ ;
	wire _w24654_ ;
	wire _w24653_ ;
	wire _w24652_ ;
	wire _w24651_ ;
	wire _w24650_ ;
	wire _w24649_ ;
	wire _w24648_ ;
	wire _w24647_ ;
	wire _w24646_ ;
	wire _w24645_ ;
	wire _w24644_ ;
	wire _w24643_ ;
	wire _w24642_ ;
	wire _w24641_ ;
	wire _w24640_ ;
	wire _w24639_ ;
	wire _w24638_ ;
	wire _w24637_ ;
	wire _w24636_ ;
	wire _w24635_ ;
	wire _w24634_ ;
	wire _w24633_ ;
	wire _w24632_ ;
	wire _w24631_ ;
	wire _w24630_ ;
	wire _w24629_ ;
	wire _w24628_ ;
	wire _w24627_ ;
	wire _w24626_ ;
	wire _w24625_ ;
	wire _w24624_ ;
	wire _w24623_ ;
	wire _w24622_ ;
	wire _w24621_ ;
	wire _w24620_ ;
	wire _w24619_ ;
	wire _w24618_ ;
	wire _w24617_ ;
	wire _w24616_ ;
	wire _w24615_ ;
	wire _w24614_ ;
	wire _w24613_ ;
	wire _w24612_ ;
	wire _w24611_ ;
	wire _w24610_ ;
	wire _w24609_ ;
	wire _w24608_ ;
	wire _w24607_ ;
	wire _w24606_ ;
	wire _w24605_ ;
	wire _w24604_ ;
	wire _w24603_ ;
	wire _w24602_ ;
	wire _w24601_ ;
	wire _w24600_ ;
	wire _w24599_ ;
	wire _w24598_ ;
	wire _w24597_ ;
	wire _w24596_ ;
	wire _w24595_ ;
	wire _w24594_ ;
	wire _w24593_ ;
	wire _w24592_ ;
	wire _w24591_ ;
	wire _w24590_ ;
	wire _w24589_ ;
	wire _w24588_ ;
	wire _w24587_ ;
	wire _w24586_ ;
	wire _w24585_ ;
	wire _w24584_ ;
	wire _w24583_ ;
	wire _w24582_ ;
	wire _w24581_ ;
	wire _w24580_ ;
	wire _w24579_ ;
	wire _w24578_ ;
	wire _w24577_ ;
	wire _w24576_ ;
	wire _w24575_ ;
	wire _w24574_ ;
	wire _w24573_ ;
	wire _w24572_ ;
	wire _w24571_ ;
	wire _w24570_ ;
	wire _w24569_ ;
	wire _w24568_ ;
	wire _w24567_ ;
	wire _w24566_ ;
	wire _w24565_ ;
	wire _w24564_ ;
	wire _w24563_ ;
	wire _w24562_ ;
	wire _w24561_ ;
	wire _w24560_ ;
	wire _w24559_ ;
	wire _w24558_ ;
	wire _w24557_ ;
	wire _w24556_ ;
	wire _w24555_ ;
	wire _w24554_ ;
	wire _w24553_ ;
	wire _w24552_ ;
	wire _w24551_ ;
	wire _w24550_ ;
	wire _w24549_ ;
	wire _w24548_ ;
	wire _w24547_ ;
	wire _w24546_ ;
	wire _w24545_ ;
	wire _w24544_ ;
	wire _w24543_ ;
	wire _w24542_ ;
	wire _w24541_ ;
	wire _w24540_ ;
	wire _w24539_ ;
	wire _w24538_ ;
	wire _w24537_ ;
	wire _w24536_ ;
	wire _w24535_ ;
	wire _w24534_ ;
	wire _w24533_ ;
	wire _w24532_ ;
	wire _w24531_ ;
	wire _w24530_ ;
	wire _w24529_ ;
	wire _w24528_ ;
	wire _w24527_ ;
	wire _w24526_ ;
	wire _w24525_ ;
	wire _w24524_ ;
	wire _w24523_ ;
	wire _w24522_ ;
	wire _w24521_ ;
	wire _w24520_ ;
	wire _w24519_ ;
	wire _w24518_ ;
	wire _w24517_ ;
	wire _w24516_ ;
	wire _w24515_ ;
	wire _w24514_ ;
	wire _w24513_ ;
	wire _w24512_ ;
	wire _w24511_ ;
	wire _w24510_ ;
	wire _w24509_ ;
	wire _w24508_ ;
	wire _w24507_ ;
	wire _w24506_ ;
	wire _w24505_ ;
	wire _w24504_ ;
	wire _w24503_ ;
	wire _w24502_ ;
	wire _w24501_ ;
	wire _w24500_ ;
	wire _w24499_ ;
	wire _w24498_ ;
	wire _w24497_ ;
	wire _w24496_ ;
	wire _w24495_ ;
	wire _w24494_ ;
	wire _w24493_ ;
	wire _w24492_ ;
	wire _w24491_ ;
	wire _w24490_ ;
	wire _w24489_ ;
	wire _w24488_ ;
	wire _w24487_ ;
	wire _w24486_ ;
	wire _w24485_ ;
	wire _w24484_ ;
	wire _w24483_ ;
	wire _w24482_ ;
	wire _w24481_ ;
	wire _w24480_ ;
	wire _w24479_ ;
	wire _w24478_ ;
	wire _w24477_ ;
	wire _w24476_ ;
	wire _w24475_ ;
	wire _w24474_ ;
	wire _w24473_ ;
	wire _w24472_ ;
	wire _w24471_ ;
	wire _w24470_ ;
	wire _w24469_ ;
	wire _w24468_ ;
	wire _w24467_ ;
	wire _w24466_ ;
	wire _w24465_ ;
	wire _w24464_ ;
	wire _w24463_ ;
	wire _w24462_ ;
	wire _w24461_ ;
	wire _w24460_ ;
	wire _w24459_ ;
	wire _w24458_ ;
	wire _w24457_ ;
	wire _w24456_ ;
	wire _w24455_ ;
	wire _w24454_ ;
	wire _w24453_ ;
	wire _w24452_ ;
	wire _w24451_ ;
	wire _w24450_ ;
	wire _w24449_ ;
	wire _w24448_ ;
	wire _w24447_ ;
	wire _w24446_ ;
	wire _w24445_ ;
	wire _w24444_ ;
	wire _w24443_ ;
	wire _w24442_ ;
	wire _w24441_ ;
	wire _w24440_ ;
	wire _w24439_ ;
	wire _w24438_ ;
	wire _w24437_ ;
	wire _w24436_ ;
	wire _w24435_ ;
	wire _w24434_ ;
	wire _w24433_ ;
	wire _w24432_ ;
	wire _w24431_ ;
	wire _w24430_ ;
	wire _w24429_ ;
	wire _w24428_ ;
	wire _w24427_ ;
	wire _w24426_ ;
	wire _w24425_ ;
	wire _w24424_ ;
	wire _w24423_ ;
	wire _w24422_ ;
	wire _w24421_ ;
	wire _w24420_ ;
	wire _w24419_ ;
	wire _w24418_ ;
	wire _w24417_ ;
	wire _w24416_ ;
	wire _w24415_ ;
	wire _w24414_ ;
	wire _w24413_ ;
	wire _w24412_ ;
	wire _w24411_ ;
	wire _w24410_ ;
	wire _w24409_ ;
	wire _w24408_ ;
	wire _w24407_ ;
	wire _w24406_ ;
	wire _w24405_ ;
	wire _w24404_ ;
	wire _w24403_ ;
	wire _w24402_ ;
	wire _w24401_ ;
	wire _w24400_ ;
	wire _w24399_ ;
	wire _w24398_ ;
	wire _w24397_ ;
	wire _w24396_ ;
	wire _w24395_ ;
	wire _w24394_ ;
	wire _w24393_ ;
	wire _w24392_ ;
	wire _w24391_ ;
	wire _w24390_ ;
	wire _w24389_ ;
	wire _w24388_ ;
	wire _w24387_ ;
	wire _w24386_ ;
	wire _w24385_ ;
	wire _w24384_ ;
	wire _w24383_ ;
	wire _w24382_ ;
	wire _w24381_ ;
	wire _w24380_ ;
	wire _w24379_ ;
	wire _w24378_ ;
	wire _w24377_ ;
	wire _w24376_ ;
	wire _w24375_ ;
	wire _w24374_ ;
	wire _w24373_ ;
	wire _w24372_ ;
	wire _w24371_ ;
	wire _w24370_ ;
	wire _w24369_ ;
	wire _w24368_ ;
	wire _w24367_ ;
	wire _w24366_ ;
	wire _w24365_ ;
	wire _w24364_ ;
	wire _w24363_ ;
	wire _w24362_ ;
	wire _w24361_ ;
	wire _w24360_ ;
	wire _w24359_ ;
	wire _w24358_ ;
	wire _w24357_ ;
	wire _w24356_ ;
	wire _w24355_ ;
	wire _w24354_ ;
	wire _w24353_ ;
	wire _w24352_ ;
	wire _w24351_ ;
	wire _w24350_ ;
	wire _w24349_ ;
	wire _w24348_ ;
	wire _w24347_ ;
	wire _w24346_ ;
	wire _w24345_ ;
	wire _w24344_ ;
	wire _w24343_ ;
	wire _w24342_ ;
	wire _w24341_ ;
	wire _w24340_ ;
	wire _w24339_ ;
	wire _w24338_ ;
	wire _w24337_ ;
	wire _w24336_ ;
	wire _w24335_ ;
	wire _w24334_ ;
	wire _w24333_ ;
	wire _w24332_ ;
	wire _w24331_ ;
	wire _w24330_ ;
	wire _w24329_ ;
	wire _w24328_ ;
	wire _w24327_ ;
	wire _w24326_ ;
	wire _w24325_ ;
	wire _w24324_ ;
	wire _w24323_ ;
	wire _w24322_ ;
	wire _w24321_ ;
	wire _w24320_ ;
	wire _w24319_ ;
	wire _w24318_ ;
	wire _w24317_ ;
	wire _w24316_ ;
	wire _w24315_ ;
	wire _w24314_ ;
	wire _w24313_ ;
	wire _w24312_ ;
	wire _w24311_ ;
	wire _w24310_ ;
	wire _w24309_ ;
	wire _w24308_ ;
	wire _w24307_ ;
	wire _w24306_ ;
	wire _w24305_ ;
	wire _w24304_ ;
	wire _w24303_ ;
	wire _w24302_ ;
	wire _w24301_ ;
	wire _w24300_ ;
	wire _w24299_ ;
	wire _w24298_ ;
	wire _w24297_ ;
	wire _w24296_ ;
	wire _w24295_ ;
	wire _w24294_ ;
	wire _w24293_ ;
	wire _w24292_ ;
	wire _w24291_ ;
	wire _w24290_ ;
	wire _w24289_ ;
	wire _w24288_ ;
	wire _w24287_ ;
	wire _w24286_ ;
	wire _w24285_ ;
	wire _w24284_ ;
	wire _w24283_ ;
	wire _w24282_ ;
	wire _w24281_ ;
	wire _w24280_ ;
	wire _w24279_ ;
	wire _w24278_ ;
	wire _w24277_ ;
	wire _w24276_ ;
	wire _w24275_ ;
	wire _w24274_ ;
	wire _w24273_ ;
	wire _w24272_ ;
	wire _w24271_ ;
	wire _w24270_ ;
	wire _w24269_ ;
	wire _w24268_ ;
	wire _w24267_ ;
	wire _w24266_ ;
	wire _w24265_ ;
	wire _w24264_ ;
	wire _w24263_ ;
	wire _w24262_ ;
	wire _w24261_ ;
	wire _w24260_ ;
	wire _w24259_ ;
	wire _w24258_ ;
	wire _w24257_ ;
	wire _w24256_ ;
	wire _w24255_ ;
	wire _w24254_ ;
	wire _w24253_ ;
	wire _w24252_ ;
	wire _w24251_ ;
	wire _w24250_ ;
	wire _w24249_ ;
	wire _w24248_ ;
	wire _w24247_ ;
	wire _w24246_ ;
	wire _w24245_ ;
	wire _w24244_ ;
	wire _w24243_ ;
	wire _w24242_ ;
	wire _w24241_ ;
	wire _w24240_ ;
	wire _w24239_ ;
	wire _w24238_ ;
	wire _w24237_ ;
	wire _w24236_ ;
	wire _w24235_ ;
	wire _w24234_ ;
	wire _w24233_ ;
	wire _w24232_ ;
	wire _w24231_ ;
	wire _w24230_ ;
	wire _w24229_ ;
	wire _w24228_ ;
	wire _w24227_ ;
	wire _w24226_ ;
	wire _w24225_ ;
	wire _w24224_ ;
	wire _w24223_ ;
	wire _w24222_ ;
	wire _w24221_ ;
	wire _w24220_ ;
	wire _w24219_ ;
	wire _w24218_ ;
	wire _w24217_ ;
	wire _w24216_ ;
	wire _w24215_ ;
	wire _w24214_ ;
	wire _w24213_ ;
	wire _w24212_ ;
	wire _w24211_ ;
	wire _w24210_ ;
	wire _w24209_ ;
	wire _w24208_ ;
	wire _w24207_ ;
	wire _w24206_ ;
	wire _w24205_ ;
	wire _w24204_ ;
	wire _w24203_ ;
	wire _w24202_ ;
	wire _w24201_ ;
	wire _w24200_ ;
	wire _w24199_ ;
	wire _w24198_ ;
	wire _w24197_ ;
	wire _w24196_ ;
	wire _w24195_ ;
	wire _w24194_ ;
	wire _w24193_ ;
	wire _w24192_ ;
	wire _w24191_ ;
	wire _w24190_ ;
	wire _w24189_ ;
	wire _w24188_ ;
	wire _w24187_ ;
	wire _w24186_ ;
	wire _w24185_ ;
	wire _w24184_ ;
	wire _w24183_ ;
	wire _w24182_ ;
	wire _w24181_ ;
	wire _w24180_ ;
	wire _w24179_ ;
	wire _w24178_ ;
	wire _w24177_ ;
	wire _w24176_ ;
	wire _w24175_ ;
	wire _w24174_ ;
	wire _w24173_ ;
	wire _w24172_ ;
	wire _w24171_ ;
	wire _w24170_ ;
	wire _w24169_ ;
	wire _w24168_ ;
	wire _w24167_ ;
	wire _w24166_ ;
	wire _w24165_ ;
	wire _w24164_ ;
	wire _w24163_ ;
	wire _w24162_ ;
	wire _w24161_ ;
	wire _w24160_ ;
	wire _w24159_ ;
	wire _w24158_ ;
	wire _w24157_ ;
	wire _w24156_ ;
	wire _w24155_ ;
	wire _w24154_ ;
	wire _w24153_ ;
	wire _w24152_ ;
	wire _w24151_ ;
	wire _w24150_ ;
	wire _w24149_ ;
	wire _w24148_ ;
	wire _w24147_ ;
	wire _w24146_ ;
	wire _w24145_ ;
	wire _w24144_ ;
	wire _w24143_ ;
	wire _w24142_ ;
	wire _w24141_ ;
	wire _w24140_ ;
	wire _w24139_ ;
	wire _w24138_ ;
	wire _w24137_ ;
	wire _w24136_ ;
	wire _w24135_ ;
	wire _w24134_ ;
	wire _w24133_ ;
	wire _w24132_ ;
	wire _w24131_ ;
	wire _w24130_ ;
	wire _w24129_ ;
	wire _w24128_ ;
	wire _w24127_ ;
	wire _w24126_ ;
	wire _w24125_ ;
	wire _w24124_ ;
	wire _w24123_ ;
	wire _w24122_ ;
	wire _w24121_ ;
	wire _w24120_ ;
	wire _w24119_ ;
	wire _w24118_ ;
	wire _w24117_ ;
	wire _w24116_ ;
	wire _w24115_ ;
	wire _w24114_ ;
	wire _w24113_ ;
	wire _w24112_ ;
	wire _w24111_ ;
	wire _w24110_ ;
	wire _w24109_ ;
	wire _w24108_ ;
	wire _w24107_ ;
	wire _w24106_ ;
	wire _w24105_ ;
	wire _w24104_ ;
	wire _w24103_ ;
	wire _w24102_ ;
	wire _w24101_ ;
	wire _w24100_ ;
	wire _w24099_ ;
	wire _w24098_ ;
	wire _w24097_ ;
	wire _w24096_ ;
	wire _w24095_ ;
	wire _w24094_ ;
	wire _w24093_ ;
	wire _w24092_ ;
	wire _w24091_ ;
	wire _w24090_ ;
	wire _w24089_ ;
	wire _w24088_ ;
	wire _w24087_ ;
	wire _w24086_ ;
	wire _w24085_ ;
	wire _w24084_ ;
	wire _w24083_ ;
	wire _w24082_ ;
	wire _w24081_ ;
	wire _w24080_ ;
	wire _w24079_ ;
	wire _w24078_ ;
	wire _w24077_ ;
	wire _w24076_ ;
	wire _w24075_ ;
	wire _w24074_ ;
	wire _w24073_ ;
	wire _w24072_ ;
	wire _w24071_ ;
	wire _w24070_ ;
	wire _w24069_ ;
	wire _w24068_ ;
	wire _w24067_ ;
	wire _w24066_ ;
	wire _w24065_ ;
	wire _w24064_ ;
	wire _w24063_ ;
	wire _w24062_ ;
	wire _w24061_ ;
	wire _w24060_ ;
	wire _w24059_ ;
	wire _w24058_ ;
	wire _w24057_ ;
	wire _w24056_ ;
	wire _w24055_ ;
	wire _w24054_ ;
	wire _w24053_ ;
	wire _w24052_ ;
	wire _w24051_ ;
	wire _w24050_ ;
	wire _w24049_ ;
	wire _w24048_ ;
	wire _w24047_ ;
	wire _w24046_ ;
	wire _w24045_ ;
	wire _w24044_ ;
	wire _w24043_ ;
	wire _w24042_ ;
	wire _w24041_ ;
	wire _w24040_ ;
	wire _w24039_ ;
	wire _w24038_ ;
	wire _w24037_ ;
	wire _w24036_ ;
	wire _w24035_ ;
	wire _w24034_ ;
	wire _w24033_ ;
	wire _w24032_ ;
	wire _w24031_ ;
	wire _w24030_ ;
	wire _w24029_ ;
	wire _w24028_ ;
	wire _w24027_ ;
	wire _w24026_ ;
	wire _w24025_ ;
	wire _w24024_ ;
	wire _w24023_ ;
	wire _w24022_ ;
	wire _w24021_ ;
	wire _w24020_ ;
	wire _w24019_ ;
	wire _w24018_ ;
	wire _w24017_ ;
	wire _w24016_ ;
	wire _w24015_ ;
	wire _w24014_ ;
	wire _w24013_ ;
	wire _w24012_ ;
	wire _w24011_ ;
	wire _w24010_ ;
	wire _w24009_ ;
	wire _w24008_ ;
	wire _w24007_ ;
	wire _w24006_ ;
	wire _w24005_ ;
	wire _w24004_ ;
	wire _w24003_ ;
	wire _w24002_ ;
	wire _w24001_ ;
	wire _w24000_ ;
	wire _w23999_ ;
	wire _w23998_ ;
	wire _w23997_ ;
	wire _w23996_ ;
	wire _w23995_ ;
	wire _w23994_ ;
	wire _w23993_ ;
	wire _w23992_ ;
	wire _w23991_ ;
	wire _w23990_ ;
	wire _w23989_ ;
	wire _w23988_ ;
	wire _w23987_ ;
	wire _w23986_ ;
	wire _w23985_ ;
	wire _w23984_ ;
	wire _w23983_ ;
	wire _w23982_ ;
	wire _w23981_ ;
	wire _w23980_ ;
	wire _w23979_ ;
	wire _w23978_ ;
	wire _w23977_ ;
	wire _w23976_ ;
	wire _w23975_ ;
	wire _w23974_ ;
	wire _w23973_ ;
	wire _w23972_ ;
	wire _w23971_ ;
	wire _w23970_ ;
	wire _w23969_ ;
	wire _w23968_ ;
	wire _w23967_ ;
	wire _w23966_ ;
	wire _w23965_ ;
	wire _w23964_ ;
	wire _w23963_ ;
	wire _w23962_ ;
	wire _w23961_ ;
	wire _w23960_ ;
	wire _w23959_ ;
	wire _w23958_ ;
	wire _w23957_ ;
	wire _w23956_ ;
	wire _w23955_ ;
	wire _w23954_ ;
	wire _w23953_ ;
	wire _w23952_ ;
	wire _w23951_ ;
	wire _w23950_ ;
	wire _w23949_ ;
	wire _w23948_ ;
	wire _w23947_ ;
	wire _w23946_ ;
	wire _w23945_ ;
	wire _w23944_ ;
	wire _w23943_ ;
	wire _w23942_ ;
	wire _w23941_ ;
	wire _w23940_ ;
	wire _w23939_ ;
	wire _w23938_ ;
	wire _w23937_ ;
	wire _w23936_ ;
	wire _w23935_ ;
	wire _w23934_ ;
	wire _w23933_ ;
	wire _w23932_ ;
	wire _w23931_ ;
	wire _w23930_ ;
	wire _w23929_ ;
	wire _w23928_ ;
	wire _w23927_ ;
	wire _w23926_ ;
	wire _w23925_ ;
	wire _w23924_ ;
	wire _w23923_ ;
	wire _w23922_ ;
	wire _w23921_ ;
	wire _w23920_ ;
	wire _w23919_ ;
	wire _w23918_ ;
	wire _w23917_ ;
	wire _w23916_ ;
	wire _w23915_ ;
	wire _w23914_ ;
	wire _w23913_ ;
	wire _w23912_ ;
	wire _w23911_ ;
	wire _w23910_ ;
	wire _w23909_ ;
	wire _w23908_ ;
	wire _w23907_ ;
	wire _w23906_ ;
	wire _w23905_ ;
	wire _w23904_ ;
	wire _w23903_ ;
	wire _w23902_ ;
	wire _w23901_ ;
	wire _w23900_ ;
	wire _w23899_ ;
	wire _w23898_ ;
	wire _w23897_ ;
	wire _w23896_ ;
	wire _w23895_ ;
	wire _w23894_ ;
	wire _w23893_ ;
	wire _w23892_ ;
	wire _w23891_ ;
	wire _w23890_ ;
	wire _w23889_ ;
	wire _w23888_ ;
	wire _w23887_ ;
	wire _w23886_ ;
	wire _w23885_ ;
	wire _w23884_ ;
	wire _w23883_ ;
	wire _w23882_ ;
	wire _w23881_ ;
	wire _w23880_ ;
	wire _w23879_ ;
	wire _w23878_ ;
	wire _w23877_ ;
	wire _w23876_ ;
	wire _w23875_ ;
	wire _w23874_ ;
	wire _w23873_ ;
	wire _w23872_ ;
	wire _w23871_ ;
	wire _w23870_ ;
	wire _w23869_ ;
	wire _w23868_ ;
	wire _w23867_ ;
	wire _w23866_ ;
	wire _w23865_ ;
	wire _w23864_ ;
	wire _w23863_ ;
	wire _w23862_ ;
	wire _w23861_ ;
	wire _w23860_ ;
	wire _w23859_ ;
	wire _w23858_ ;
	wire _w23857_ ;
	wire _w23856_ ;
	wire _w23855_ ;
	wire _w23854_ ;
	wire _w23853_ ;
	wire _w23852_ ;
	wire _w23851_ ;
	wire _w23850_ ;
	wire _w23849_ ;
	wire _w23848_ ;
	wire _w23847_ ;
	wire _w23846_ ;
	wire _w23845_ ;
	wire _w23844_ ;
	wire _w23843_ ;
	wire _w23842_ ;
	wire _w23841_ ;
	wire _w23840_ ;
	wire _w23839_ ;
	wire _w23838_ ;
	wire _w23837_ ;
	wire _w23836_ ;
	wire _w23835_ ;
	wire _w23834_ ;
	wire _w23833_ ;
	wire _w23832_ ;
	wire _w23831_ ;
	wire _w23830_ ;
	wire _w23829_ ;
	wire _w23828_ ;
	wire _w23827_ ;
	wire _w23826_ ;
	wire _w23825_ ;
	wire _w23824_ ;
	wire _w23823_ ;
	wire _w23822_ ;
	wire _w23821_ ;
	wire _w23820_ ;
	wire _w23819_ ;
	wire _w23818_ ;
	wire _w23817_ ;
	wire _w23816_ ;
	wire _w23815_ ;
	wire _w23814_ ;
	wire _w23813_ ;
	wire _w23812_ ;
	wire _w23811_ ;
	wire _w23810_ ;
	wire _w23809_ ;
	wire _w23808_ ;
	wire _w23807_ ;
	wire _w23806_ ;
	wire _w23805_ ;
	wire _w23804_ ;
	wire _w23803_ ;
	wire _w23802_ ;
	wire _w23801_ ;
	wire _w23800_ ;
	wire _w23799_ ;
	wire _w23798_ ;
	wire _w23797_ ;
	wire _w23796_ ;
	wire _w23795_ ;
	wire _w23794_ ;
	wire _w23793_ ;
	wire _w23792_ ;
	wire _w23791_ ;
	wire _w23790_ ;
	wire _w23789_ ;
	wire _w23788_ ;
	wire _w23787_ ;
	wire _w23786_ ;
	wire _w23785_ ;
	wire _w23784_ ;
	wire _w23783_ ;
	wire _w23782_ ;
	wire _w23781_ ;
	wire _w23780_ ;
	wire _w23779_ ;
	wire _w23778_ ;
	wire _w23777_ ;
	wire _w23776_ ;
	wire _w23775_ ;
	wire _w23774_ ;
	wire _w23773_ ;
	wire _w23772_ ;
	wire _w23771_ ;
	wire _w23770_ ;
	wire _w23769_ ;
	wire _w23768_ ;
	wire _w23767_ ;
	wire _w23766_ ;
	wire _w23765_ ;
	wire _w23764_ ;
	wire _w23763_ ;
	wire _w23762_ ;
	wire _w23761_ ;
	wire _w23760_ ;
	wire _w23759_ ;
	wire _w23758_ ;
	wire _w23757_ ;
	wire _w23756_ ;
	wire _w23755_ ;
	wire _w23754_ ;
	wire _w23753_ ;
	wire _w23752_ ;
	wire _w23751_ ;
	wire _w23750_ ;
	wire _w23749_ ;
	wire _w23748_ ;
	wire _w23747_ ;
	wire _w23746_ ;
	wire _w23745_ ;
	wire _w23744_ ;
	wire _w23743_ ;
	wire _w23742_ ;
	wire _w23741_ ;
	wire _w23740_ ;
	wire _w23739_ ;
	wire _w23738_ ;
	wire _w23737_ ;
	wire _w23736_ ;
	wire _w23735_ ;
	wire _w23734_ ;
	wire _w23733_ ;
	wire _w23732_ ;
	wire _w23731_ ;
	wire _w23730_ ;
	wire _w23729_ ;
	wire _w23728_ ;
	wire _w23727_ ;
	wire _w23726_ ;
	wire _w23725_ ;
	wire _w23724_ ;
	wire _w23723_ ;
	wire _w23722_ ;
	wire _w23721_ ;
	wire _w23720_ ;
	wire _w23719_ ;
	wire _w23718_ ;
	wire _w23717_ ;
	wire _w23716_ ;
	wire _w23715_ ;
	wire _w23714_ ;
	wire _w23713_ ;
	wire _w23712_ ;
	wire _w23711_ ;
	wire _w23710_ ;
	wire _w23709_ ;
	wire _w23708_ ;
	wire _w23707_ ;
	wire _w23706_ ;
	wire _w23705_ ;
	wire _w23704_ ;
	wire _w23703_ ;
	wire _w23702_ ;
	wire _w23701_ ;
	wire _w23700_ ;
	wire _w23699_ ;
	wire _w23698_ ;
	wire _w23697_ ;
	wire _w23696_ ;
	wire _w23695_ ;
	wire _w23694_ ;
	wire _w23693_ ;
	wire _w23692_ ;
	wire _w23691_ ;
	wire _w23690_ ;
	wire _w23689_ ;
	wire _w23688_ ;
	wire _w23687_ ;
	wire _w23686_ ;
	wire _w23685_ ;
	wire _w23684_ ;
	wire _w23683_ ;
	wire _w23682_ ;
	wire _w23681_ ;
	wire _w23680_ ;
	wire _w23679_ ;
	wire _w23678_ ;
	wire _w23677_ ;
	wire _w23676_ ;
	wire _w23675_ ;
	wire _w23674_ ;
	wire _w23673_ ;
	wire _w23672_ ;
	wire _w23671_ ;
	wire _w23670_ ;
	wire _w23669_ ;
	wire _w23668_ ;
	wire _w23667_ ;
	wire _w23666_ ;
	wire _w23665_ ;
	wire _w23664_ ;
	wire _w23663_ ;
	wire _w23662_ ;
	wire _w23661_ ;
	wire _w23660_ ;
	wire _w23659_ ;
	wire _w23658_ ;
	wire _w23657_ ;
	wire _w23656_ ;
	wire _w23655_ ;
	wire _w23654_ ;
	wire _w23653_ ;
	wire _w23652_ ;
	wire _w23651_ ;
	wire _w23650_ ;
	wire _w23649_ ;
	wire _w23648_ ;
	wire _w23647_ ;
	wire _w23646_ ;
	wire _w23645_ ;
	wire _w23644_ ;
	wire _w23643_ ;
	wire _w23642_ ;
	wire _w23641_ ;
	wire _w23640_ ;
	wire _w23639_ ;
	wire _w23638_ ;
	wire _w23637_ ;
	wire _w23636_ ;
	wire _w23635_ ;
	wire _w23634_ ;
	wire _w23633_ ;
	wire _w23632_ ;
	wire _w23631_ ;
	wire _w23630_ ;
	wire _w23629_ ;
	wire _w23628_ ;
	wire _w23627_ ;
	wire _w23626_ ;
	wire _w23625_ ;
	wire _w23624_ ;
	wire _w23623_ ;
	wire _w23622_ ;
	wire _w23621_ ;
	wire _w23620_ ;
	wire _w23619_ ;
	wire _w23618_ ;
	wire _w23617_ ;
	wire _w23616_ ;
	wire _w23615_ ;
	wire _w23614_ ;
	wire _w23613_ ;
	wire _w23612_ ;
	wire _w23611_ ;
	wire _w23610_ ;
	wire _w23609_ ;
	wire _w23608_ ;
	wire _w23607_ ;
	wire _w23606_ ;
	wire _w23605_ ;
	wire _w23604_ ;
	wire _w23603_ ;
	wire _w23602_ ;
	wire _w23601_ ;
	wire _w23600_ ;
	wire _w23599_ ;
	wire _w23598_ ;
	wire _w23597_ ;
	wire _w23596_ ;
	wire _w23595_ ;
	wire _w23594_ ;
	wire _w23593_ ;
	wire _w23592_ ;
	wire _w23591_ ;
	wire _w23590_ ;
	wire _w23589_ ;
	wire _w23588_ ;
	wire _w23587_ ;
	wire _w23586_ ;
	wire _w23585_ ;
	wire _w23584_ ;
	wire _w23583_ ;
	wire _w23582_ ;
	wire _w23581_ ;
	wire _w23580_ ;
	wire _w23579_ ;
	wire _w23578_ ;
	wire _w23577_ ;
	wire _w23576_ ;
	wire _w23575_ ;
	wire _w23574_ ;
	wire _w23573_ ;
	wire _w23572_ ;
	wire _w23571_ ;
	wire _w23570_ ;
	wire _w23569_ ;
	wire _w23568_ ;
	wire _w23567_ ;
	wire _w23566_ ;
	wire _w23565_ ;
	wire _w23564_ ;
	wire _w23563_ ;
	wire _w23562_ ;
	wire _w23561_ ;
	wire _w23560_ ;
	wire _w23559_ ;
	wire _w23558_ ;
	wire _w23557_ ;
	wire _w23556_ ;
	wire _w23555_ ;
	wire _w23554_ ;
	wire _w23553_ ;
	wire _w23552_ ;
	wire _w23551_ ;
	wire _w23550_ ;
	wire _w23549_ ;
	wire _w23548_ ;
	wire _w23547_ ;
	wire _w23546_ ;
	wire _w23545_ ;
	wire _w23544_ ;
	wire _w23543_ ;
	wire _w23542_ ;
	wire _w23541_ ;
	wire _w23540_ ;
	wire _w23539_ ;
	wire _w23538_ ;
	wire _w23537_ ;
	wire _w23536_ ;
	wire _w23535_ ;
	wire _w23534_ ;
	wire _w23533_ ;
	wire _w23532_ ;
	wire _w23531_ ;
	wire _w23530_ ;
	wire _w23529_ ;
	wire _w23528_ ;
	wire _w23527_ ;
	wire _w23526_ ;
	wire _w23525_ ;
	wire _w23524_ ;
	wire _w23523_ ;
	wire _w23522_ ;
	wire _w23521_ ;
	wire _w23520_ ;
	wire _w23519_ ;
	wire _w23518_ ;
	wire _w23517_ ;
	wire _w23516_ ;
	wire _w23515_ ;
	wire _w23514_ ;
	wire _w23513_ ;
	wire _w23512_ ;
	wire _w23511_ ;
	wire _w23510_ ;
	wire _w23509_ ;
	wire _w23508_ ;
	wire _w23507_ ;
	wire _w23506_ ;
	wire _w23505_ ;
	wire _w23504_ ;
	wire _w23503_ ;
	wire _w23502_ ;
	wire _w23501_ ;
	wire _w23500_ ;
	wire _w23499_ ;
	wire _w23498_ ;
	wire _w23497_ ;
	wire _w23496_ ;
	wire _w23495_ ;
	wire _w23494_ ;
	wire _w23493_ ;
	wire _w23492_ ;
	wire _w23491_ ;
	wire _w23490_ ;
	wire _w23489_ ;
	wire _w23488_ ;
	wire _w23487_ ;
	wire _w23486_ ;
	wire _w23485_ ;
	wire _w23484_ ;
	wire _w23483_ ;
	wire _w23482_ ;
	wire _w23481_ ;
	wire _w23480_ ;
	wire _w23479_ ;
	wire _w23478_ ;
	wire _w23477_ ;
	wire _w23476_ ;
	wire _w23475_ ;
	wire _w23474_ ;
	wire _w23473_ ;
	wire _w23472_ ;
	wire _w23471_ ;
	wire _w23470_ ;
	wire _w23469_ ;
	wire _w23468_ ;
	wire _w23467_ ;
	wire _w23466_ ;
	wire _w23465_ ;
	wire _w23464_ ;
	wire _w23463_ ;
	wire _w23462_ ;
	wire _w23461_ ;
	wire _w23460_ ;
	wire _w23459_ ;
	wire _w23458_ ;
	wire _w23457_ ;
	wire _w23456_ ;
	wire _w23455_ ;
	wire _w23454_ ;
	wire _w23453_ ;
	wire _w23452_ ;
	wire _w23451_ ;
	wire _w23450_ ;
	wire _w23449_ ;
	wire _w23448_ ;
	wire _w23447_ ;
	wire _w23446_ ;
	wire _w23445_ ;
	wire _w23444_ ;
	wire _w23443_ ;
	wire _w23442_ ;
	wire _w23441_ ;
	wire _w23440_ ;
	wire _w23439_ ;
	wire _w23438_ ;
	wire _w23437_ ;
	wire _w23436_ ;
	wire _w23435_ ;
	wire _w23434_ ;
	wire _w23433_ ;
	wire _w23432_ ;
	wire _w23431_ ;
	wire _w23430_ ;
	wire _w23429_ ;
	wire _w23428_ ;
	wire _w23427_ ;
	wire _w23426_ ;
	wire _w23425_ ;
	wire _w23424_ ;
	wire _w23423_ ;
	wire _w23422_ ;
	wire _w23421_ ;
	wire _w23420_ ;
	wire _w23419_ ;
	wire _w23418_ ;
	wire _w23417_ ;
	wire _w23416_ ;
	wire _w23415_ ;
	wire _w23414_ ;
	wire _w23413_ ;
	wire _w23412_ ;
	wire _w23411_ ;
	wire _w23410_ ;
	wire _w23409_ ;
	wire _w23408_ ;
	wire _w23407_ ;
	wire _w23406_ ;
	wire _w23405_ ;
	wire _w23404_ ;
	wire _w23403_ ;
	wire _w23402_ ;
	wire _w23401_ ;
	wire _w23400_ ;
	wire _w23399_ ;
	wire _w23398_ ;
	wire _w23397_ ;
	wire _w23396_ ;
	wire _w23395_ ;
	wire _w23394_ ;
	wire _w23393_ ;
	wire _w23392_ ;
	wire _w23391_ ;
	wire _w23390_ ;
	wire _w23389_ ;
	wire _w23388_ ;
	wire _w23387_ ;
	wire _w23386_ ;
	wire _w23385_ ;
	wire _w23384_ ;
	wire _w23383_ ;
	wire _w23382_ ;
	wire _w23381_ ;
	wire _w23380_ ;
	wire _w23379_ ;
	wire _w23378_ ;
	wire _w23377_ ;
	wire _w23376_ ;
	wire _w23375_ ;
	wire _w23374_ ;
	wire _w23373_ ;
	wire _w23372_ ;
	wire _w23371_ ;
	wire _w23370_ ;
	wire _w23369_ ;
	wire _w23368_ ;
	wire _w23367_ ;
	wire _w23366_ ;
	wire _w23365_ ;
	wire _w23364_ ;
	wire _w23363_ ;
	wire _w23362_ ;
	wire _w23361_ ;
	wire _w23360_ ;
	wire _w23359_ ;
	wire _w23358_ ;
	wire _w23357_ ;
	wire _w23356_ ;
	wire _w23355_ ;
	wire _w23354_ ;
	wire _w23353_ ;
	wire _w23352_ ;
	wire _w23351_ ;
	wire _w23350_ ;
	wire _w23349_ ;
	wire _w23348_ ;
	wire _w23347_ ;
	wire _w23346_ ;
	wire _w23345_ ;
	wire _w23344_ ;
	wire _w23343_ ;
	wire _w23342_ ;
	wire _w23341_ ;
	wire _w23340_ ;
	wire _w23339_ ;
	wire _w23338_ ;
	wire _w23337_ ;
	wire _w23336_ ;
	wire _w23335_ ;
	wire _w23334_ ;
	wire _w23333_ ;
	wire _w23332_ ;
	wire _w23331_ ;
	wire _w23330_ ;
	wire _w23329_ ;
	wire _w23328_ ;
	wire _w23327_ ;
	wire _w23326_ ;
	wire _w23325_ ;
	wire _w23324_ ;
	wire _w23323_ ;
	wire _w23322_ ;
	wire _w23321_ ;
	wire _w23320_ ;
	wire _w23319_ ;
	wire _w23318_ ;
	wire _w23317_ ;
	wire _w23316_ ;
	wire _w23315_ ;
	wire _w23314_ ;
	wire _w23313_ ;
	wire _w23312_ ;
	wire _w23311_ ;
	wire _w23310_ ;
	wire _w23309_ ;
	wire _w23308_ ;
	wire _w23307_ ;
	wire _w23306_ ;
	wire _w23305_ ;
	wire _w23304_ ;
	wire _w23303_ ;
	wire _w23302_ ;
	wire _w23301_ ;
	wire _w23300_ ;
	wire _w23299_ ;
	wire _w23298_ ;
	wire _w23297_ ;
	wire _w23296_ ;
	wire _w23295_ ;
	wire _w23294_ ;
	wire _w23293_ ;
	wire _w23292_ ;
	wire _w23291_ ;
	wire _w23290_ ;
	wire _w23289_ ;
	wire _w23288_ ;
	wire _w23287_ ;
	wire _w23286_ ;
	wire _w23285_ ;
	wire _w23284_ ;
	wire _w23283_ ;
	wire _w23282_ ;
	wire _w23281_ ;
	wire _w23280_ ;
	wire _w23279_ ;
	wire _w23278_ ;
	wire _w23277_ ;
	wire _w23276_ ;
	wire _w23275_ ;
	wire _w23274_ ;
	wire _w23273_ ;
	wire _w23272_ ;
	wire _w23271_ ;
	wire _w23270_ ;
	wire _w23269_ ;
	wire _w23268_ ;
	wire _w23267_ ;
	wire _w23266_ ;
	wire _w23265_ ;
	wire _w23264_ ;
	wire _w23263_ ;
	wire _w23262_ ;
	wire _w23261_ ;
	wire _w23260_ ;
	wire _w23259_ ;
	wire _w23258_ ;
	wire _w23257_ ;
	wire _w23256_ ;
	wire _w23255_ ;
	wire _w23254_ ;
	wire _w23253_ ;
	wire _w23252_ ;
	wire _w23251_ ;
	wire _w23250_ ;
	wire _w23249_ ;
	wire _w23248_ ;
	wire _w23247_ ;
	wire _w23246_ ;
	wire _w23245_ ;
	wire _w23244_ ;
	wire _w23243_ ;
	wire _w23242_ ;
	wire _w23241_ ;
	wire _w23240_ ;
	wire _w23239_ ;
	wire _w23238_ ;
	wire _w23237_ ;
	wire _w23236_ ;
	wire _w23235_ ;
	wire _w23234_ ;
	wire _w23233_ ;
	wire _w23232_ ;
	wire _w23231_ ;
	wire _w23230_ ;
	wire _w23229_ ;
	wire _w23228_ ;
	wire _w23227_ ;
	wire _w23226_ ;
	wire _w23225_ ;
	wire _w23224_ ;
	wire _w23223_ ;
	wire _w23222_ ;
	wire _w23221_ ;
	wire _w23220_ ;
	wire _w23219_ ;
	wire _w23218_ ;
	wire _w23217_ ;
	wire _w23216_ ;
	wire _w23215_ ;
	wire _w23214_ ;
	wire _w23213_ ;
	wire _w23212_ ;
	wire _w23211_ ;
	wire _w23210_ ;
	wire _w23209_ ;
	wire _w23208_ ;
	wire _w23207_ ;
	wire _w23206_ ;
	wire _w23205_ ;
	wire _w23204_ ;
	wire _w23203_ ;
	wire _w23202_ ;
	wire _w23201_ ;
	wire _w23200_ ;
	wire _w23199_ ;
	wire _w23198_ ;
	wire _w23197_ ;
	wire _w23196_ ;
	wire _w23195_ ;
	wire _w23194_ ;
	wire _w23193_ ;
	wire _w23192_ ;
	wire _w23191_ ;
	wire _w23190_ ;
	wire _w23189_ ;
	wire _w23188_ ;
	wire _w23187_ ;
	wire _w23186_ ;
	wire _w23185_ ;
	wire _w23184_ ;
	wire _w23183_ ;
	wire _w23182_ ;
	wire _w23181_ ;
	wire _w23180_ ;
	wire _w23179_ ;
	wire _w23178_ ;
	wire _w23177_ ;
	wire _w23176_ ;
	wire _w23175_ ;
	wire _w23174_ ;
	wire _w23173_ ;
	wire _w23172_ ;
	wire _w23171_ ;
	wire _w23170_ ;
	wire _w23169_ ;
	wire _w23168_ ;
	wire _w23167_ ;
	wire _w23166_ ;
	wire _w23165_ ;
	wire _w23164_ ;
	wire _w23163_ ;
	wire _w23162_ ;
	wire _w23161_ ;
	wire _w23160_ ;
	wire _w23159_ ;
	wire _w23158_ ;
	wire _w23157_ ;
	wire _w23156_ ;
	wire _w23155_ ;
	wire _w23154_ ;
	wire _w23153_ ;
	wire _w23152_ ;
	wire _w23151_ ;
	wire _w23150_ ;
	wire _w23149_ ;
	wire _w23148_ ;
	wire _w23147_ ;
	wire _w23146_ ;
	wire _w23145_ ;
	wire _w23144_ ;
	wire _w23143_ ;
	wire _w23142_ ;
	wire _w23141_ ;
	wire _w23140_ ;
	wire _w23139_ ;
	wire _w23138_ ;
	wire _w23137_ ;
	wire _w23136_ ;
	wire _w23135_ ;
	wire _w23134_ ;
	wire _w23133_ ;
	wire _w23132_ ;
	wire _w23131_ ;
	wire _w23130_ ;
	wire _w23129_ ;
	wire _w23128_ ;
	wire _w23127_ ;
	wire _w23126_ ;
	wire _w23125_ ;
	wire _w23124_ ;
	wire _w23123_ ;
	wire _w23122_ ;
	wire _w23121_ ;
	wire _w23120_ ;
	wire _w23119_ ;
	wire _w23118_ ;
	wire _w23117_ ;
	wire _w23116_ ;
	wire _w23115_ ;
	wire _w23114_ ;
	wire _w23113_ ;
	wire _w23112_ ;
	wire _w23111_ ;
	wire _w23110_ ;
	wire _w23109_ ;
	wire _w23108_ ;
	wire _w23107_ ;
	wire _w23106_ ;
	wire _w23105_ ;
	wire _w23104_ ;
	wire _w23103_ ;
	wire _w23102_ ;
	wire _w23101_ ;
	wire _w23100_ ;
	wire _w23099_ ;
	wire _w23098_ ;
	wire _w23097_ ;
	wire _w23096_ ;
	wire _w23095_ ;
	wire _w23094_ ;
	wire _w23093_ ;
	wire _w23092_ ;
	wire _w23091_ ;
	wire _w23090_ ;
	wire _w23089_ ;
	wire _w23088_ ;
	wire _w23087_ ;
	wire _w23086_ ;
	wire _w23085_ ;
	wire _w23084_ ;
	wire _w23083_ ;
	wire _w23082_ ;
	wire _w23081_ ;
	wire _w23080_ ;
	wire _w23079_ ;
	wire _w23078_ ;
	wire _w23077_ ;
	wire _w23076_ ;
	wire _w23075_ ;
	wire _w23074_ ;
	wire _w23073_ ;
	wire _w23072_ ;
	wire _w23071_ ;
	wire _w23070_ ;
	wire _w23069_ ;
	wire _w23068_ ;
	wire _w23067_ ;
	wire _w23066_ ;
	wire _w23065_ ;
	wire _w23064_ ;
	wire _w23063_ ;
	wire _w23062_ ;
	wire _w23061_ ;
	wire _w23060_ ;
	wire _w23059_ ;
	wire _w23058_ ;
	wire _w23057_ ;
	wire _w23056_ ;
	wire _w23055_ ;
	wire _w23054_ ;
	wire _w23053_ ;
	wire _w23052_ ;
	wire _w23051_ ;
	wire _w23050_ ;
	wire _w23049_ ;
	wire _w23048_ ;
	wire _w23047_ ;
	wire _w23046_ ;
	wire _w23045_ ;
	wire _w23044_ ;
	wire _w23043_ ;
	wire _w23042_ ;
	wire _w23041_ ;
	wire _w23040_ ;
	wire _w23039_ ;
	wire _w23038_ ;
	wire _w23037_ ;
	wire _w23036_ ;
	wire _w23035_ ;
	wire _w23034_ ;
	wire _w23033_ ;
	wire _w23032_ ;
	wire _w23031_ ;
	wire _w23030_ ;
	wire _w23029_ ;
	wire _w23028_ ;
	wire _w23027_ ;
	wire _w23026_ ;
	wire _w23025_ ;
	wire _w23024_ ;
	wire _w23023_ ;
	wire _w23022_ ;
	wire _w23021_ ;
	wire _w23020_ ;
	wire _w23019_ ;
	wire _w23018_ ;
	wire _w23017_ ;
	wire _w23016_ ;
	wire _w23015_ ;
	wire _w23014_ ;
	wire _w23013_ ;
	wire _w23012_ ;
	wire _w23011_ ;
	wire _w23010_ ;
	wire _w23009_ ;
	wire _w23008_ ;
	wire _w23007_ ;
	wire _w23006_ ;
	wire _w23005_ ;
	wire _w23004_ ;
	wire _w23003_ ;
	wire _w23002_ ;
	wire _w23001_ ;
	wire _w23000_ ;
	wire _w22999_ ;
	wire _w22998_ ;
	wire _w22997_ ;
	wire _w22996_ ;
	wire _w22995_ ;
	wire _w22994_ ;
	wire _w22993_ ;
	wire _w22992_ ;
	wire _w22991_ ;
	wire _w22990_ ;
	wire _w22989_ ;
	wire _w22988_ ;
	wire _w22987_ ;
	wire _w22986_ ;
	wire _w22985_ ;
	wire _w22984_ ;
	wire _w22983_ ;
	wire _w22982_ ;
	wire _w22981_ ;
	wire _w22980_ ;
	wire _w22979_ ;
	wire _w22978_ ;
	wire _w22977_ ;
	wire _w22976_ ;
	wire _w22975_ ;
	wire _w22974_ ;
	wire _w22973_ ;
	wire _w22972_ ;
	wire _w22971_ ;
	wire _w22970_ ;
	wire _w22969_ ;
	wire _w22968_ ;
	wire _w22967_ ;
	wire _w22966_ ;
	wire _w22965_ ;
	wire _w22964_ ;
	wire _w22963_ ;
	wire _w22962_ ;
	wire _w22961_ ;
	wire _w22960_ ;
	wire _w22959_ ;
	wire _w22958_ ;
	wire _w22957_ ;
	wire _w22956_ ;
	wire _w22955_ ;
	wire _w22954_ ;
	wire _w22953_ ;
	wire _w22952_ ;
	wire _w22951_ ;
	wire _w22950_ ;
	wire _w22949_ ;
	wire _w22948_ ;
	wire _w22947_ ;
	wire _w22946_ ;
	wire _w22945_ ;
	wire _w22944_ ;
	wire _w22943_ ;
	wire _w22942_ ;
	wire _w22941_ ;
	wire _w22940_ ;
	wire _w22939_ ;
	wire _w22938_ ;
	wire _w22937_ ;
	wire _w22936_ ;
	wire _w22935_ ;
	wire _w22934_ ;
	wire _w22933_ ;
	wire _w22932_ ;
	wire _w22931_ ;
	wire _w22930_ ;
	wire _w22929_ ;
	wire _w22928_ ;
	wire _w22927_ ;
	wire _w22926_ ;
	wire _w22925_ ;
	wire _w22924_ ;
	wire _w22923_ ;
	wire _w22922_ ;
	wire _w22921_ ;
	wire _w22920_ ;
	wire _w22919_ ;
	wire _w22918_ ;
	wire _w22917_ ;
	wire _w22916_ ;
	wire _w22915_ ;
	wire _w22914_ ;
	wire _w22913_ ;
	wire _w22912_ ;
	wire _w22911_ ;
	wire _w22910_ ;
	wire _w22909_ ;
	wire _w22908_ ;
	wire _w22907_ ;
	wire _w22906_ ;
	wire _w22905_ ;
	wire _w22904_ ;
	wire _w22903_ ;
	wire _w22902_ ;
	wire _w22901_ ;
	wire _w22900_ ;
	wire _w22899_ ;
	wire _w22898_ ;
	wire _w22897_ ;
	wire _w22896_ ;
	wire _w22895_ ;
	wire _w22894_ ;
	wire _w22893_ ;
	wire _w22892_ ;
	wire _w22891_ ;
	wire _w22890_ ;
	wire _w22889_ ;
	wire _w22888_ ;
	wire _w22887_ ;
	wire _w22886_ ;
	wire _w22885_ ;
	wire _w22884_ ;
	wire _w22883_ ;
	wire _w22882_ ;
	wire _w22881_ ;
	wire _w22880_ ;
	wire _w22879_ ;
	wire _w22878_ ;
	wire _w22877_ ;
	wire _w22876_ ;
	wire _w22875_ ;
	wire _w22874_ ;
	wire _w22873_ ;
	wire _w22872_ ;
	wire _w22871_ ;
	wire _w22870_ ;
	wire _w22869_ ;
	wire _w22868_ ;
	wire _w22867_ ;
	wire _w22866_ ;
	wire _w22865_ ;
	wire _w22864_ ;
	wire _w22863_ ;
	wire _w22862_ ;
	wire _w22861_ ;
	wire _w22860_ ;
	wire _w22859_ ;
	wire _w22858_ ;
	wire _w22857_ ;
	wire _w22856_ ;
	wire _w22855_ ;
	wire _w22854_ ;
	wire _w22853_ ;
	wire _w22852_ ;
	wire _w22851_ ;
	wire _w22850_ ;
	wire _w22849_ ;
	wire _w22848_ ;
	wire _w22847_ ;
	wire _w22846_ ;
	wire _w22845_ ;
	wire _w22844_ ;
	wire _w22843_ ;
	wire _w22842_ ;
	wire _w22841_ ;
	wire _w22840_ ;
	wire _w22839_ ;
	wire _w22838_ ;
	wire _w22837_ ;
	wire _w22836_ ;
	wire _w22835_ ;
	wire _w22834_ ;
	wire _w22833_ ;
	wire _w22832_ ;
	wire _w22831_ ;
	wire _w22830_ ;
	wire _w22829_ ;
	wire _w22828_ ;
	wire _w22827_ ;
	wire _w22826_ ;
	wire _w22825_ ;
	wire _w22824_ ;
	wire _w22823_ ;
	wire _w22822_ ;
	wire _w22821_ ;
	wire _w22820_ ;
	wire _w22819_ ;
	wire _w22818_ ;
	wire _w22817_ ;
	wire _w22816_ ;
	wire _w22815_ ;
	wire _w22814_ ;
	wire _w22813_ ;
	wire _w22812_ ;
	wire _w22811_ ;
	wire _w22810_ ;
	wire _w22809_ ;
	wire _w22808_ ;
	wire _w22807_ ;
	wire _w22806_ ;
	wire _w22805_ ;
	wire _w22804_ ;
	wire _w22803_ ;
	wire _w22802_ ;
	wire _w22801_ ;
	wire _w22800_ ;
	wire _w22799_ ;
	wire _w22798_ ;
	wire _w22797_ ;
	wire _w22796_ ;
	wire _w22795_ ;
	wire _w22794_ ;
	wire _w22793_ ;
	wire _w22792_ ;
	wire _w22791_ ;
	wire _w22790_ ;
	wire _w22789_ ;
	wire _w22788_ ;
	wire _w22787_ ;
	wire _w22786_ ;
	wire _w22785_ ;
	wire _w22784_ ;
	wire _w22783_ ;
	wire _w22782_ ;
	wire _w22781_ ;
	wire _w22780_ ;
	wire _w22779_ ;
	wire _w22778_ ;
	wire _w22777_ ;
	wire _w22776_ ;
	wire _w22775_ ;
	wire _w22774_ ;
	wire _w22773_ ;
	wire _w22772_ ;
	wire _w22771_ ;
	wire _w22770_ ;
	wire _w22769_ ;
	wire _w22768_ ;
	wire _w22767_ ;
	wire _w22766_ ;
	wire _w22765_ ;
	wire _w22764_ ;
	wire _w22763_ ;
	wire _w22762_ ;
	wire _w22761_ ;
	wire _w22760_ ;
	wire _w22759_ ;
	wire _w22758_ ;
	wire _w22757_ ;
	wire _w22756_ ;
	wire _w22755_ ;
	wire _w22754_ ;
	wire _w22753_ ;
	wire _w22752_ ;
	wire _w22751_ ;
	wire _w22750_ ;
	wire _w22749_ ;
	wire _w22748_ ;
	wire _w22747_ ;
	wire _w22746_ ;
	wire _w22745_ ;
	wire _w22744_ ;
	wire _w22743_ ;
	wire _w22742_ ;
	wire _w22741_ ;
	wire _w22740_ ;
	wire _w22739_ ;
	wire _w22738_ ;
	wire _w22737_ ;
	wire _w22736_ ;
	wire _w22735_ ;
	wire _w22734_ ;
	wire _w22733_ ;
	wire _w22732_ ;
	wire _w22731_ ;
	wire _w22730_ ;
	wire _w22729_ ;
	wire _w22728_ ;
	wire _w22727_ ;
	wire _w22726_ ;
	wire _w22725_ ;
	wire _w22724_ ;
	wire _w22723_ ;
	wire _w22722_ ;
	wire _w22721_ ;
	wire _w22720_ ;
	wire _w22719_ ;
	wire _w22718_ ;
	wire _w22717_ ;
	wire _w22716_ ;
	wire _w22715_ ;
	wire _w22714_ ;
	wire _w22713_ ;
	wire _w22712_ ;
	wire _w22711_ ;
	wire _w22710_ ;
	wire _w22709_ ;
	wire _w22708_ ;
	wire _w22707_ ;
	wire _w22706_ ;
	wire _w22705_ ;
	wire _w22704_ ;
	wire _w22703_ ;
	wire _w22702_ ;
	wire _w22701_ ;
	wire _w22700_ ;
	wire _w22699_ ;
	wire _w22698_ ;
	wire _w22697_ ;
	wire _w22696_ ;
	wire _w22695_ ;
	wire _w22694_ ;
	wire _w22693_ ;
	wire _w22692_ ;
	wire _w22691_ ;
	wire _w22690_ ;
	wire _w22689_ ;
	wire _w22688_ ;
	wire _w22687_ ;
	wire _w22686_ ;
	wire _w22685_ ;
	wire _w22684_ ;
	wire _w22683_ ;
	wire _w22682_ ;
	wire _w22681_ ;
	wire _w22680_ ;
	wire _w22679_ ;
	wire _w22678_ ;
	wire _w22677_ ;
	wire _w22676_ ;
	wire _w22675_ ;
	wire _w22674_ ;
	wire _w22673_ ;
	wire _w22672_ ;
	wire _w22671_ ;
	wire _w22670_ ;
	wire _w22669_ ;
	wire _w22668_ ;
	wire _w22667_ ;
	wire _w22666_ ;
	wire _w22665_ ;
	wire _w22664_ ;
	wire _w22663_ ;
	wire _w22662_ ;
	wire _w22661_ ;
	wire _w22660_ ;
	wire _w22659_ ;
	wire _w22658_ ;
	wire _w22657_ ;
	wire _w22656_ ;
	wire _w22655_ ;
	wire _w22654_ ;
	wire _w22653_ ;
	wire _w22652_ ;
	wire _w22651_ ;
	wire _w22650_ ;
	wire _w22649_ ;
	wire _w22648_ ;
	wire _w22647_ ;
	wire _w22646_ ;
	wire _w22645_ ;
	wire _w22644_ ;
	wire _w22643_ ;
	wire _w22642_ ;
	wire _w22641_ ;
	wire _w22640_ ;
	wire _w22639_ ;
	wire _w22638_ ;
	wire _w22637_ ;
	wire _w22636_ ;
	wire _w22635_ ;
	wire _w22634_ ;
	wire _w22633_ ;
	wire _w22632_ ;
	wire _w22631_ ;
	wire _w22630_ ;
	wire _w22629_ ;
	wire _w22628_ ;
	wire _w22627_ ;
	wire _w22626_ ;
	wire _w22625_ ;
	wire _w22624_ ;
	wire _w22623_ ;
	wire _w22622_ ;
	wire _w22621_ ;
	wire _w22620_ ;
	wire _w22619_ ;
	wire _w22618_ ;
	wire _w22617_ ;
	wire _w22616_ ;
	wire _w22615_ ;
	wire _w22614_ ;
	wire _w22613_ ;
	wire _w22612_ ;
	wire _w22611_ ;
	wire _w22610_ ;
	wire _w22609_ ;
	wire _w22608_ ;
	wire _w22607_ ;
	wire _w22606_ ;
	wire _w22605_ ;
	wire _w22604_ ;
	wire _w22603_ ;
	wire _w22602_ ;
	wire _w22601_ ;
	wire _w22600_ ;
	wire _w22599_ ;
	wire _w22598_ ;
	wire _w22597_ ;
	wire _w22596_ ;
	wire _w22595_ ;
	wire _w22594_ ;
	wire _w22593_ ;
	wire _w22592_ ;
	wire _w22591_ ;
	wire _w22590_ ;
	wire _w22589_ ;
	wire _w22588_ ;
	wire _w22587_ ;
	wire _w22586_ ;
	wire _w22585_ ;
	wire _w22584_ ;
	wire _w22583_ ;
	wire _w22582_ ;
	wire _w22581_ ;
	wire _w22580_ ;
	wire _w22579_ ;
	wire _w22578_ ;
	wire _w22577_ ;
	wire _w22576_ ;
	wire _w22575_ ;
	wire _w22574_ ;
	wire _w22573_ ;
	wire _w22572_ ;
	wire _w22571_ ;
	wire _w22570_ ;
	wire _w22569_ ;
	wire _w22568_ ;
	wire _w22567_ ;
	wire _w22566_ ;
	wire _w22565_ ;
	wire _w22564_ ;
	wire _w22563_ ;
	wire _w22562_ ;
	wire _w22561_ ;
	wire _w22560_ ;
	wire _w22559_ ;
	wire _w22558_ ;
	wire _w22557_ ;
	wire _w22556_ ;
	wire _w22555_ ;
	wire _w22554_ ;
	wire _w22553_ ;
	wire _w22552_ ;
	wire _w22551_ ;
	wire _w22550_ ;
	wire _w22549_ ;
	wire _w22548_ ;
	wire _w22547_ ;
	wire _w22546_ ;
	wire _w22545_ ;
	wire _w22544_ ;
	wire _w22543_ ;
	wire _w22542_ ;
	wire _w22541_ ;
	wire _w22540_ ;
	wire _w22539_ ;
	wire _w22538_ ;
	wire _w22537_ ;
	wire _w22536_ ;
	wire _w22535_ ;
	wire _w22534_ ;
	wire _w22533_ ;
	wire _w22532_ ;
	wire _w22531_ ;
	wire _w22530_ ;
	wire _w22529_ ;
	wire _w22528_ ;
	wire _w22527_ ;
	wire _w22526_ ;
	wire _w22525_ ;
	wire _w22524_ ;
	wire _w22523_ ;
	wire _w22522_ ;
	wire _w22521_ ;
	wire _w22520_ ;
	wire _w22519_ ;
	wire _w22518_ ;
	wire _w22517_ ;
	wire _w22516_ ;
	wire _w22515_ ;
	wire _w22514_ ;
	wire _w22513_ ;
	wire _w22512_ ;
	wire _w22511_ ;
	wire _w22510_ ;
	wire _w22509_ ;
	wire _w22508_ ;
	wire _w22507_ ;
	wire _w22506_ ;
	wire _w22505_ ;
	wire _w22504_ ;
	wire _w22503_ ;
	wire _w22502_ ;
	wire _w22501_ ;
	wire _w22500_ ;
	wire _w22499_ ;
	wire _w22498_ ;
	wire _w22497_ ;
	wire _w22496_ ;
	wire _w22495_ ;
	wire _w22494_ ;
	wire _w22493_ ;
	wire _w22492_ ;
	wire _w22491_ ;
	wire _w22490_ ;
	wire _w22489_ ;
	wire _w22488_ ;
	wire _w22487_ ;
	wire _w22486_ ;
	wire _w22485_ ;
	wire _w22484_ ;
	wire _w22483_ ;
	wire _w22482_ ;
	wire _w22481_ ;
	wire _w22480_ ;
	wire _w22479_ ;
	wire _w22478_ ;
	wire _w22477_ ;
	wire _w22476_ ;
	wire _w22475_ ;
	wire _w22474_ ;
	wire _w22473_ ;
	wire _w22472_ ;
	wire _w22471_ ;
	wire _w22470_ ;
	wire _w22469_ ;
	wire _w22468_ ;
	wire _w22467_ ;
	wire _w22466_ ;
	wire _w22465_ ;
	wire _w22464_ ;
	wire _w22463_ ;
	wire _w22462_ ;
	wire _w22461_ ;
	wire _w22460_ ;
	wire _w22459_ ;
	wire _w22458_ ;
	wire _w22457_ ;
	wire _w22456_ ;
	wire _w22455_ ;
	wire _w22454_ ;
	wire _w22453_ ;
	wire _w22452_ ;
	wire _w22451_ ;
	wire _w22450_ ;
	wire _w22449_ ;
	wire _w22448_ ;
	wire _w22447_ ;
	wire _w22446_ ;
	wire _w22445_ ;
	wire _w22444_ ;
	wire _w22443_ ;
	wire _w22442_ ;
	wire _w22441_ ;
	wire _w22440_ ;
	wire _w22439_ ;
	wire _w22438_ ;
	wire _w22437_ ;
	wire _w22436_ ;
	wire _w22435_ ;
	wire _w22434_ ;
	wire _w22433_ ;
	wire _w22432_ ;
	wire _w22431_ ;
	wire _w22430_ ;
	wire _w22429_ ;
	wire _w22428_ ;
	wire _w22427_ ;
	wire _w22426_ ;
	wire _w22425_ ;
	wire _w22424_ ;
	wire _w22423_ ;
	wire _w22422_ ;
	wire _w22421_ ;
	wire _w22420_ ;
	wire _w22419_ ;
	wire _w22418_ ;
	wire _w22417_ ;
	wire _w22416_ ;
	wire _w22415_ ;
	wire _w22414_ ;
	wire _w22413_ ;
	wire _w22412_ ;
	wire _w22411_ ;
	wire _w22410_ ;
	wire _w22409_ ;
	wire _w22408_ ;
	wire _w22407_ ;
	wire _w22406_ ;
	wire _w22405_ ;
	wire _w22404_ ;
	wire _w22403_ ;
	wire _w22402_ ;
	wire _w22401_ ;
	wire _w22400_ ;
	wire _w22399_ ;
	wire _w22398_ ;
	wire _w22397_ ;
	wire _w22396_ ;
	wire _w22395_ ;
	wire _w22394_ ;
	wire _w22393_ ;
	wire _w22392_ ;
	wire _w22391_ ;
	wire _w22390_ ;
	wire _w22389_ ;
	wire _w22388_ ;
	wire _w22387_ ;
	wire _w22386_ ;
	wire _w22385_ ;
	wire _w22384_ ;
	wire _w22383_ ;
	wire _w22382_ ;
	wire _w22381_ ;
	wire _w22380_ ;
	wire _w22379_ ;
	wire _w22378_ ;
	wire _w22377_ ;
	wire _w22376_ ;
	wire _w22375_ ;
	wire _w22374_ ;
	wire _w22373_ ;
	wire _w22372_ ;
	wire _w22371_ ;
	wire _w22370_ ;
	wire _w22369_ ;
	wire _w22368_ ;
	wire _w22367_ ;
	wire _w22366_ ;
	wire _w22365_ ;
	wire _w22364_ ;
	wire _w22363_ ;
	wire _w22362_ ;
	wire _w22361_ ;
	wire _w22360_ ;
	wire _w22359_ ;
	wire _w22358_ ;
	wire _w22357_ ;
	wire _w22356_ ;
	wire _w22355_ ;
	wire _w22354_ ;
	wire _w22353_ ;
	wire _w22352_ ;
	wire _w22351_ ;
	wire _w22350_ ;
	wire _w22349_ ;
	wire _w22348_ ;
	wire _w22347_ ;
	wire _w22346_ ;
	wire _w22345_ ;
	wire _w22344_ ;
	wire _w22343_ ;
	wire _w22342_ ;
	wire _w22341_ ;
	wire _w22340_ ;
	wire _w22339_ ;
	wire _w22338_ ;
	wire _w22337_ ;
	wire _w22336_ ;
	wire _w22335_ ;
	wire _w22334_ ;
	wire _w22333_ ;
	wire _w22332_ ;
	wire _w22331_ ;
	wire _w22330_ ;
	wire _w22329_ ;
	wire _w22328_ ;
	wire _w22327_ ;
	wire _w22326_ ;
	wire _w22325_ ;
	wire _w22324_ ;
	wire _w22323_ ;
	wire _w22322_ ;
	wire _w22321_ ;
	wire _w22320_ ;
	wire _w22319_ ;
	wire _w22318_ ;
	wire _w22317_ ;
	wire _w22316_ ;
	wire _w22315_ ;
	wire _w22314_ ;
	wire _w22313_ ;
	wire _w22312_ ;
	wire _w22311_ ;
	wire _w22310_ ;
	wire _w22309_ ;
	wire _w22308_ ;
	wire _w22307_ ;
	wire _w22306_ ;
	wire _w22305_ ;
	wire _w22304_ ;
	wire _w22303_ ;
	wire _w22302_ ;
	wire _w22301_ ;
	wire _w22300_ ;
	wire _w22299_ ;
	wire _w22298_ ;
	wire _w22297_ ;
	wire _w22296_ ;
	wire _w22295_ ;
	wire _w22294_ ;
	wire _w22293_ ;
	wire _w22292_ ;
	wire _w22291_ ;
	wire _w22290_ ;
	wire _w22289_ ;
	wire _w22288_ ;
	wire _w22287_ ;
	wire _w22286_ ;
	wire _w22285_ ;
	wire _w22284_ ;
	wire _w22283_ ;
	wire _w22282_ ;
	wire _w22281_ ;
	wire _w22280_ ;
	wire _w22279_ ;
	wire _w22278_ ;
	wire _w22277_ ;
	wire _w22276_ ;
	wire _w22275_ ;
	wire _w22274_ ;
	wire _w22273_ ;
	wire _w22272_ ;
	wire _w22271_ ;
	wire _w22270_ ;
	wire _w22269_ ;
	wire _w22268_ ;
	wire _w22267_ ;
	wire _w22266_ ;
	wire _w22265_ ;
	wire _w22264_ ;
	wire _w22263_ ;
	wire _w22262_ ;
	wire _w22261_ ;
	wire _w22260_ ;
	wire _w22259_ ;
	wire _w22258_ ;
	wire _w22257_ ;
	wire _w22256_ ;
	wire _w22255_ ;
	wire _w22254_ ;
	wire _w22253_ ;
	wire _w22252_ ;
	wire _w22251_ ;
	wire _w22250_ ;
	wire _w22249_ ;
	wire _w22248_ ;
	wire _w22247_ ;
	wire _w22246_ ;
	wire _w22245_ ;
	wire _w22244_ ;
	wire _w22243_ ;
	wire _w22242_ ;
	wire _w22241_ ;
	wire _w22240_ ;
	wire _w22239_ ;
	wire _w22238_ ;
	wire _w22237_ ;
	wire _w22236_ ;
	wire _w22235_ ;
	wire _w22234_ ;
	wire _w22233_ ;
	wire _w22232_ ;
	wire _w22231_ ;
	wire _w22230_ ;
	wire _w22229_ ;
	wire _w22228_ ;
	wire _w22227_ ;
	wire _w22226_ ;
	wire _w22225_ ;
	wire _w22224_ ;
	wire _w22223_ ;
	wire _w22222_ ;
	wire _w22221_ ;
	wire _w22220_ ;
	wire _w22219_ ;
	wire _w22218_ ;
	wire _w22217_ ;
	wire _w22216_ ;
	wire _w22215_ ;
	wire _w22214_ ;
	wire _w22213_ ;
	wire _w22212_ ;
	wire _w22211_ ;
	wire _w22210_ ;
	wire _w22209_ ;
	wire _w22208_ ;
	wire _w22207_ ;
	wire _w22206_ ;
	wire _w22205_ ;
	wire _w22204_ ;
	wire _w22203_ ;
	wire _w22202_ ;
	wire _w22201_ ;
	wire _w22200_ ;
	wire _w22199_ ;
	wire _w22198_ ;
	wire _w22197_ ;
	wire _w22196_ ;
	wire _w22195_ ;
	wire _w22194_ ;
	wire _w22193_ ;
	wire _w22192_ ;
	wire _w22191_ ;
	wire _w22190_ ;
	wire _w22189_ ;
	wire _w22188_ ;
	wire _w22187_ ;
	wire _w22186_ ;
	wire _w22185_ ;
	wire _w22184_ ;
	wire _w22183_ ;
	wire _w22182_ ;
	wire _w22181_ ;
	wire _w22180_ ;
	wire _w22179_ ;
	wire _w22178_ ;
	wire _w22177_ ;
	wire _w22176_ ;
	wire _w22175_ ;
	wire _w22174_ ;
	wire _w22173_ ;
	wire _w22172_ ;
	wire _w22171_ ;
	wire _w22170_ ;
	wire _w22169_ ;
	wire _w22168_ ;
	wire _w22167_ ;
	wire _w22166_ ;
	wire _w22165_ ;
	wire _w22164_ ;
	wire _w22163_ ;
	wire _w22162_ ;
	wire _w22161_ ;
	wire _w22160_ ;
	wire _w22159_ ;
	wire _w22158_ ;
	wire _w22157_ ;
	wire _w22156_ ;
	wire _w22155_ ;
	wire _w22154_ ;
	wire _w22153_ ;
	wire _w22152_ ;
	wire _w22151_ ;
	wire _w22150_ ;
	wire _w22149_ ;
	wire _w22148_ ;
	wire _w22147_ ;
	wire _w22146_ ;
	wire _w22145_ ;
	wire _w22144_ ;
	wire _w22143_ ;
	wire _w22142_ ;
	wire _w22141_ ;
	wire _w22140_ ;
	wire _w22139_ ;
	wire _w22138_ ;
	wire _w22137_ ;
	wire _w22136_ ;
	wire _w22135_ ;
	wire _w22134_ ;
	wire _w22133_ ;
	wire _w22132_ ;
	wire _w22131_ ;
	wire _w22130_ ;
	wire _w22129_ ;
	wire _w22128_ ;
	wire _w22127_ ;
	wire _w22126_ ;
	wire _w22125_ ;
	wire _w22124_ ;
	wire _w22123_ ;
	wire _w22122_ ;
	wire _w22121_ ;
	wire _w22120_ ;
	wire _w22119_ ;
	wire _w22118_ ;
	wire _w22117_ ;
	wire _w22116_ ;
	wire _w22115_ ;
	wire _w22114_ ;
	wire _w22113_ ;
	wire _w22112_ ;
	wire _w22111_ ;
	wire _w22110_ ;
	wire _w22109_ ;
	wire _w22108_ ;
	wire _w22107_ ;
	wire _w22106_ ;
	wire _w22105_ ;
	wire _w22104_ ;
	wire _w22103_ ;
	wire _w22102_ ;
	wire _w22101_ ;
	wire _w22100_ ;
	wire _w22099_ ;
	wire _w22098_ ;
	wire _w22097_ ;
	wire _w22096_ ;
	wire _w22095_ ;
	wire _w22094_ ;
	wire _w22093_ ;
	wire _w22092_ ;
	wire _w22091_ ;
	wire _w22090_ ;
	wire _w22089_ ;
	wire _w22088_ ;
	wire _w22087_ ;
	wire _w22086_ ;
	wire _w22085_ ;
	wire _w22084_ ;
	wire _w22083_ ;
	wire _w22082_ ;
	wire _w22081_ ;
	wire _w22080_ ;
	wire _w22079_ ;
	wire _w22078_ ;
	wire _w22077_ ;
	wire _w22076_ ;
	wire _w22075_ ;
	wire _w22074_ ;
	wire _w22073_ ;
	wire _w22072_ ;
	wire _w22071_ ;
	wire _w22070_ ;
	wire _w22069_ ;
	wire _w22068_ ;
	wire _w22067_ ;
	wire _w22066_ ;
	wire _w22065_ ;
	wire _w22064_ ;
	wire _w22063_ ;
	wire _w22062_ ;
	wire _w22061_ ;
	wire _w22060_ ;
	wire _w22059_ ;
	wire _w22058_ ;
	wire _w22057_ ;
	wire _w22056_ ;
	wire _w22055_ ;
	wire _w22054_ ;
	wire _w22053_ ;
	wire _w22052_ ;
	wire _w22051_ ;
	wire _w22050_ ;
	wire _w22049_ ;
	wire _w22048_ ;
	wire _w22047_ ;
	wire _w22046_ ;
	wire _w22045_ ;
	wire _w22044_ ;
	wire _w22043_ ;
	wire _w22042_ ;
	wire _w22041_ ;
	wire _w22040_ ;
	wire _w22039_ ;
	wire _w22038_ ;
	wire _w22037_ ;
	wire _w22036_ ;
	wire _w22035_ ;
	wire _w22034_ ;
	wire _w22033_ ;
	wire _w22032_ ;
	wire _w22031_ ;
	wire _w22030_ ;
	wire _w22029_ ;
	wire _w22028_ ;
	wire _w22027_ ;
	wire _w22026_ ;
	wire _w22025_ ;
	wire _w22024_ ;
	wire _w22023_ ;
	wire _w22022_ ;
	wire _w22021_ ;
	wire _w22020_ ;
	wire _w22019_ ;
	wire _w22018_ ;
	wire _w22017_ ;
	wire _w22016_ ;
	wire _w22015_ ;
	wire _w22014_ ;
	wire _w22013_ ;
	wire _w22012_ ;
	wire _w22011_ ;
	wire _w22010_ ;
	wire _w22009_ ;
	wire _w22008_ ;
	wire _w22007_ ;
	wire _w22006_ ;
	wire _w22005_ ;
	wire _w22004_ ;
	wire _w22003_ ;
	wire _w22002_ ;
	wire _w22001_ ;
	wire _w22000_ ;
	wire _w21999_ ;
	wire _w21998_ ;
	wire _w21997_ ;
	wire _w21996_ ;
	wire _w21995_ ;
	wire _w21994_ ;
	wire _w21993_ ;
	wire _w21992_ ;
	wire _w21991_ ;
	wire _w21990_ ;
	wire _w21989_ ;
	wire _w21988_ ;
	wire _w21987_ ;
	wire _w21986_ ;
	wire _w21985_ ;
	wire _w21984_ ;
	wire _w21983_ ;
	wire _w21982_ ;
	wire _w21981_ ;
	wire _w21980_ ;
	wire _w21979_ ;
	wire _w21978_ ;
	wire _w21977_ ;
	wire _w21976_ ;
	wire _w21975_ ;
	wire _w21974_ ;
	wire _w21973_ ;
	wire _w21972_ ;
	wire _w21971_ ;
	wire _w21970_ ;
	wire _w21969_ ;
	wire _w21968_ ;
	wire _w21967_ ;
	wire _w21966_ ;
	wire _w21965_ ;
	wire _w21964_ ;
	wire _w21963_ ;
	wire _w21962_ ;
	wire _w21961_ ;
	wire _w21960_ ;
	wire _w21959_ ;
	wire _w21958_ ;
	wire _w21957_ ;
	wire _w21956_ ;
	wire _w21955_ ;
	wire _w21954_ ;
	wire _w21953_ ;
	wire _w21952_ ;
	wire _w21951_ ;
	wire _w21950_ ;
	wire _w21949_ ;
	wire _w21948_ ;
	wire _w21947_ ;
	wire _w21946_ ;
	wire _w21945_ ;
	wire _w21944_ ;
	wire _w21943_ ;
	wire _w21942_ ;
	wire _w21941_ ;
	wire _w21940_ ;
	wire _w21939_ ;
	wire _w21938_ ;
	wire _w21937_ ;
	wire _w21936_ ;
	wire _w21935_ ;
	wire _w21934_ ;
	wire _w21933_ ;
	wire _w21932_ ;
	wire _w21931_ ;
	wire _w21930_ ;
	wire _w21929_ ;
	wire _w21928_ ;
	wire _w21927_ ;
	wire _w21926_ ;
	wire _w21925_ ;
	wire _w21924_ ;
	wire _w21923_ ;
	wire _w21922_ ;
	wire _w21921_ ;
	wire _w21920_ ;
	wire _w21919_ ;
	wire _w21918_ ;
	wire _w21917_ ;
	wire _w21916_ ;
	wire _w21915_ ;
	wire _w21914_ ;
	wire _w21913_ ;
	wire _w21912_ ;
	wire _w21911_ ;
	wire _w21910_ ;
	wire _w21909_ ;
	wire _w21908_ ;
	wire _w21907_ ;
	wire _w21906_ ;
	wire _w21905_ ;
	wire _w21904_ ;
	wire _w21903_ ;
	wire _w21902_ ;
	wire _w21901_ ;
	wire _w21900_ ;
	wire _w21899_ ;
	wire _w21898_ ;
	wire _w21897_ ;
	wire _w21896_ ;
	wire _w21895_ ;
	wire _w21894_ ;
	wire _w21893_ ;
	wire _w21892_ ;
	wire _w21891_ ;
	wire _w21890_ ;
	wire _w21889_ ;
	wire _w21888_ ;
	wire _w21887_ ;
	wire _w21886_ ;
	wire _w21885_ ;
	wire _w21884_ ;
	wire _w21883_ ;
	wire _w21882_ ;
	wire _w21881_ ;
	wire _w21880_ ;
	wire _w21879_ ;
	wire _w21878_ ;
	wire _w21877_ ;
	wire _w21876_ ;
	wire _w21875_ ;
	wire _w21874_ ;
	wire _w21873_ ;
	wire _w21872_ ;
	wire _w21871_ ;
	wire _w21870_ ;
	wire _w21869_ ;
	wire _w21868_ ;
	wire _w21867_ ;
	wire _w21866_ ;
	wire _w21865_ ;
	wire _w21864_ ;
	wire _w21863_ ;
	wire _w21862_ ;
	wire _w21861_ ;
	wire _w21860_ ;
	wire _w21859_ ;
	wire _w21858_ ;
	wire _w21857_ ;
	wire _w21856_ ;
	wire _w21855_ ;
	wire _w21854_ ;
	wire _w21853_ ;
	wire _w21852_ ;
	wire _w21851_ ;
	wire _w21850_ ;
	wire _w21849_ ;
	wire _w21848_ ;
	wire _w21847_ ;
	wire _w21846_ ;
	wire _w21845_ ;
	wire _w21844_ ;
	wire _w21843_ ;
	wire _w21842_ ;
	wire _w21841_ ;
	wire _w21840_ ;
	wire _w21839_ ;
	wire _w21838_ ;
	wire _w21837_ ;
	wire _w21836_ ;
	wire _w21835_ ;
	wire _w21834_ ;
	wire _w21833_ ;
	wire _w21832_ ;
	wire _w21831_ ;
	wire _w21830_ ;
	wire _w21829_ ;
	wire _w21828_ ;
	wire _w21827_ ;
	wire _w21826_ ;
	wire _w21825_ ;
	wire _w21824_ ;
	wire _w21823_ ;
	wire _w21822_ ;
	wire _w21821_ ;
	wire _w21820_ ;
	wire _w21819_ ;
	wire _w21818_ ;
	wire _w21817_ ;
	wire _w21816_ ;
	wire _w21815_ ;
	wire _w21814_ ;
	wire _w21813_ ;
	wire _w21812_ ;
	wire _w21811_ ;
	wire _w21810_ ;
	wire _w21809_ ;
	wire _w21808_ ;
	wire _w21807_ ;
	wire _w21806_ ;
	wire _w21805_ ;
	wire _w21804_ ;
	wire _w21803_ ;
	wire _w21802_ ;
	wire _w21801_ ;
	wire _w21800_ ;
	wire _w21799_ ;
	wire _w21798_ ;
	wire _w21797_ ;
	wire _w21796_ ;
	wire _w21795_ ;
	wire _w21794_ ;
	wire _w21793_ ;
	wire _w21792_ ;
	wire _w21791_ ;
	wire _w21790_ ;
	wire _w21789_ ;
	wire _w21788_ ;
	wire _w21787_ ;
	wire _w21786_ ;
	wire _w21785_ ;
	wire _w21784_ ;
	wire _w21783_ ;
	wire _w21782_ ;
	wire _w21781_ ;
	wire _w21780_ ;
	wire _w21779_ ;
	wire _w21778_ ;
	wire _w21777_ ;
	wire _w21776_ ;
	wire _w21775_ ;
	wire _w21774_ ;
	wire _w21773_ ;
	wire _w21772_ ;
	wire _w21771_ ;
	wire _w21770_ ;
	wire _w21769_ ;
	wire _w21768_ ;
	wire _w21767_ ;
	wire _w21766_ ;
	wire _w21765_ ;
	wire _w21764_ ;
	wire _w21763_ ;
	wire _w21762_ ;
	wire _w21761_ ;
	wire _w21760_ ;
	wire _w21759_ ;
	wire _w21758_ ;
	wire _w21757_ ;
	wire _w21756_ ;
	wire _w21755_ ;
	wire _w21754_ ;
	wire _w21753_ ;
	wire _w21752_ ;
	wire _w21751_ ;
	wire _w21750_ ;
	wire _w21749_ ;
	wire _w21748_ ;
	wire _w21747_ ;
	wire _w21746_ ;
	wire _w21745_ ;
	wire _w21744_ ;
	wire _w21743_ ;
	wire _w21742_ ;
	wire _w21741_ ;
	wire _w21740_ ;
	wire _w21739_ ;
	wire _w21738_ ;
	wire _w21737_ ;
	wire _w21736_ ;
	wire _w21735_ ;
	wire _w21734_ ;
	wire _w21733_ ;
	wire _w21732_ ;
	wire _w21731_ ;
	wire _w21730_ ;
	wire _w21729_ ;
	wire _w21728_ ;
	wire _w21727_ ;
	wire _w21726_ ;
	wire _w21725_ ;
	wire _w21724_ ;
	wire _w21723_ ;
	wire _w21722_ ;
	wire _w21721_ ;
	wire _w21720_ ;
	wire _w21719_ ;
	wire _w21718_ ;
	wire _w21717_ ;
	wire _w21716_ ;
	wire _w21715_ ;
	wire _w21714_ ;
	wire _w21713_ ;
	wire _w21712_ ;
	wire _w21711_ ;
	wire _w21710_ ;
	wire _w21709_ ;
	wire _w21708_ ;
	wire _w21707_ ;
	wire _w21706_ ;
	wire _w21705_ ;
	wire _w21704_ ;
	wire _w21703_ ;
	wire _w21702_ ;
	wire _w21701_ ;
	wire _w21700_ ;
	wire _w21699_ ;
	wire _w21698_ ;
	wire _w21697_ ;
	wire _w21696_ ;
	wire _w21695_ ;
	wire _w21694_ ;
	wire _w21693_ ;
	wire _w21692_ ;
	wire _w21691_ ;
	wire _w21690_ ;
	wire _w21689_ ;
	wire _w21688_ ;
	wire _w21687_ ;
	wire _w21686_ ;
	wire _w21685_ ;
	wire _w21684_ ;
	wire _w21683_ ;
	wire _w21682_ ;
	wire _w21681_ ;
	wire _w21680_ ;
	wire _w21679_ ;
	wire _w21678_ ;
	wire _w21677_ ;
	wire _w21676_ ;
	wire _w21675_ ;
	wire _w21674_ ;
	wire _w21673_ ;
	wire _w21672_ ;
	wire _w21671_ ;
	wire _w21670_ ;
	wire _w21669_ ;
	wire _w21668_ ;
	wire _w21667_ ;
	wire _w21666_ ;
	wire _w21665_ ;
	wire _w21664_ ;
	wire _w21663_ ;
	wire _w21662_ ;
	wire _w21661_ ;
	wire _w21660_ ;
	wire _w21659_ ;
	wire _w21658_ ;
	wire _w21657_ ;
	wire _w21656_ ;
	wire _w21655_ ;
	wire _w21654_ ;
	wire _w21653_ ;
	wire _w21652_ ;
	wire _w21651_ ;
	wire _w21650_ ;
	wire _w21649_ ;
	wire _w21648_ ;
	wire _w21647_ ;
	wire _w21646_ ;
	wire _w21645_ ;
	wire _w21644_ ;
	wire _w21643_ ;
	wire _w21642_ ;
	wire _w21641_ ;
	wire _w21640_ ;
	wire _w21639_ ;
	wire _w21638_ ;
	wire _w21637_ ;
	wire _w21636_ ;
	wire _w21635_ ;
	wire _w21634_ ;
	wire _w21633_ ;
	wire _w21632_ ;
	wire _w21631_ ;
	wire _w21630_ ;
	wire _w21629_ ;
	wire _w21628_ ;
	wire _w21627_ ;
	wire _w21626_ ;
	wire _w21625_ ;
	wire _w21624_ ;
	wire _w21623_ ;
	wire _w21622_ ;
	wire _w21621_ ;
	wire _w21620_ ;
	wire _w21619_ ;
	wire _w21618_ ;
	wire _w21617_ ;
	wire _w21616_ ;
	wire _w21615_ ;
	wire _w21614_ ;
	wire _w21613_ ;
	wire _w21612_ ;
	wire _w21611_ ;
	wire _w21610_ ;
	wire _w21609_ ;
	wire _w21608_ ;
	wire _w21607_ ;
	wire _w21606_ ;
	wire _w21605_ ;
	wire _w21604_ ;
	wire _w21603_ ;
	wire _w21602_ ;
	wire _w21601_ ;
	wire _w21600_ ;
	wire _w21599_ ;
	wire _w21598_ ;
	wire _w21597_ ;
	wire _w21596_ ;
	wire _w21595_ ;
	wire _w21594_ ;
	wire _w21593_ ;
	wire _w21592_ ;
	wire _w21591_ ;
	wire _w21590_ ;
	wire _w21589_ ;
	wire _w21588_ ;
	wire _w21587_ ;
	wire _w21586_ ;
	wire _w21585_ ;
	wire _w21584_ ;
	wire _w21583_ ;
	wire _w21582_ ;
	wire _w21581_ ;
	wire _w21580_ ;
	wire _w21579_ ;
	wire _w21578_ ;
	wire _w21577_ ;
	wire _w21576_ ;
	wire _w21575_ ;
	wire _w21574_ ;
	wire _w21573_ ;
	wire _w21572_ ;
	wire _w21571_ ;
	wire _w21570_ ;
	wire _w21569_ ;
	wire _w21568_ ;
	wire _w21567_ ;
	wire _w21566_ ;
	wire _w21565_ ;
	wire _w21564_ ;
	wire _w21563_ ;
	wire _w21562_ ;
	wire _w21561_ ;
	wire _w21560_ ;
	wire _w21559_ ;
	wire _w21558_ ;
	wire _w21557_ ;
	wire _w21556_ ;
	wire _w21555_ ;
	wire _w21554_ ;
	wire _w21553_ ;
	wire _w21552_ ;
	wire _w21551_ ;
	wire _w21550_ ;
	wire _w21549_ ;
	wire _w21548_ ;
	wire _w21547_ ;
	wire _w21546_ ;
	wire _w21545_ ;
	wire _w21544_ ;
	wire _w21543_ ;
	wire _w21542_ ;
	wire _w21541_ ;
	wire _w21540_ ;
	wire _w21539_ ;
	wire _w21538_ ;
	wire _w21537_ ;
	wire _w21536_ ;
	wire _w21535_ ;
	wire _w21534_ ;
	wire _w21533_ ;
	wire _w21532_ ;
	wire _w21531_ ;
	wire _w21530_ ;
	wire _w21529_ ;
	wire _w21528_ ;
	wire _w21527_ ;
	wire _w21526_ ;
	wire _w21525_ ;
	wire _w21524_ ;
	wire _w21523_ ;
	wire _w21522_ ;
	wire _w21521_ ;
	wire _w21520_ ;
	wire _w21519_ ;
	wire _w21518_ ;
	wire _w21517_ ;
	wire _w21516_ ;
	wire _w21515_ ;
	wire _w21514_ ;
	wire _w21513_ ;
	wire _w21512_ ;
	wire _w21511_ ;
	wire _w21510_ ;
	wire _w21509_ ;
	wire _w21508_ ;
	wire _w21507_ ;
	wire _w21506_ ;
	wire _w21505_ ;
	wire _w21504_ ;
	wire _w21503_ ;
	wire _w21502_ ;
	wire _w21501_ ;
	wire _w21500_ ;
	wire _w21499_ ;
	wire _w21498_ ;
	wire _w21497_ ;
	wire _w21496_ ;
	wire _w21495_ ;
	wire _w21494_ ;
	wire _w21493_ ;
	wire _w21492_ ;
	wire _w21491_ ;
	wire _w21490_ ;
	wire _w21489_ ;
	wire _w21488_ ;
	wire _w21487_ ;
	wire _w21486_ ;
	wire _w21485_ ;
	wire _w21484_ ;
	wire _w21483_ ;
	wire _w21482_ ;
	wire _w21481_ ;
	wire _w21480_ ;
	wire _w21479_ ;
	wire _w21478_ ;
	wire _w21477_ ;
	wire _w21476_ ;
	wire _w21475_ ;
	wire _w21474_ ;
	wire _w21473_ ;
	wire _w21472_ ;
	wire _w21471_ ;
	wire _w21470_ ;
	wire _w21469_ ;
	wire _w21468_ ;
	wire _w21467_ ;
	wire _w21466_ ;
	wire _w21465_ ;
	wire _w21464_ ;
	wire _w21463_ ;
	wire _w21462_ ;
	wire _w21461_ ;
	wire _w21460_ ;
	wire _w21459_ ;
	wire _w21458_ ;
	wire _w21457_ ;
	wire _w21456_ ;
	wire _w21455_ ;
	wire _w21454_ ;
	wire _w21453_ ;
	wire _w21452_ ;
	wire _w21451_ ;
	wire _w21450_ ;
	wire _w21449_ ;
	wire _w21448_ ;
	wire _w21447_ ;
	wire _w21446_ ;
	wire _w21445_ ;
	wire _w21444_ ;
	wire _w21443_ ;
	wire _w21442_ ;
	wire _w21441_ ;
	wire _w21440_ ;
	wire _w21439_ ;
	wire _w21438_ ;
	wire _w21437_ ;
	wire _w21436_ ;
	wire _w21435_ ;
	wire _w21434_ ;
	wire _w21433_ ;
	wire _w21432_ ;
	wire _w21431_ ;
	wire _w21430_ ;
	wire _w21429_ ;
	wire _w21428_ ;
	wire _w21427_ ;
	wire _w21426_ ;
	wire _w21425_ ;
	wire _w21424_ ;
	wire _w21423_ ;
	wire _w21422_ ;
	wire _w21421_ ;
	wire _w21420_ ;
	wire _w21419_ ;
	wire _w21418_ ;
	wire _w21417_ ;
	wire _w21416_ ;
	wire _w21415_ ;
	wire _w21414_ ;
	wire _w21413_ ;
	wire _w21412_ ;
	wire _w21411_ ;
	wire _w21410_ ;
	wire _w21409_ ;
	wire _w21408_ ;
	wire _w21407_ ;
	wire _w21406_ ;
	wire _w21405_ ;
	wire _w21404_ ;
	wire _w21403_ ;
	wire _w21402_ ;
	wire _w21401_ ;
	wire _w21400_ ;
	wire _w21399_ ;
	wire _w21398_ ;
	wire _w21397_ ;
	wire _w21396_ ;
	wire _w21395_ ;
	wire _w21394_ ;
	wire _w21393_ ;
	wire _w21392_ ;
	wire _w21391_ ;
	wire _w21390_ ;
	wire _w21389_ ;
	wire _w21388_ ;
	wire _w21387_ ;
	wire _w21386_ ;
	wire _w21385_ ;
	wire _w21384_ ;
	wire _w21383_ ;
	wire _w21382_ ;
	wire _w21381_ ;
	wire _w21380_ ;
	wire _w21379_ ;
	wire _w21378_ ;
	wire _w21377_ ;
	wire _w21376_ ;
	wire _w21375_ ;
	wire _w21374_ ;
	wire _w21373_ ;
	wire _w21372_ ;
	wire _w21371_ ;
	wire _w21370_ ;
	wire _w21369_ ;
	wire _w21368_ ;
	wire _w21367_ ;
	wire _w21366_ ;
	wire _w21365_ ;
	wire _w21364_ ;
	wire _w21363_ ;
	wire _w21362_ ;
	wire _w21361_ ;
	wire _w21360_ ;
	wire _w21359_ ;
	wire _w21358_ ;
	wire _w21357_ ;
	wire _w21356_ ;
	wire _w21355_ ;
	wire _w21354_ ;
	wire _w21353_ ;
	wire _w21352_ ;
	wire _w21351_ ;
	wire _w21350_ ;
	wire _w21349_ ;
	wire _w21348_ ;
	wire _w21347_ ;
	wire _w21346_ ;
	wire _w21345_ ;
	wire _w21344_ ;
	wire _w21343_ ;
	wire _w21342_ ;
	wire _w21341_ ;
	wire _w21340_ ;
	wire _w21339_ ;
	wire _w21338_ ;
	wire _w21337_ ;
	wire _w21336_ ;
	wire _w21335_ ;
	wire _w21334_ ;
	wire _w21333_ ;
	wire _w21332_ ;
	wire _w21331_ ;
	wire _w21330_ ;
	wire _w21329_ ;
	wire _w21328_ ;
	wire _w21327_ ;
	wire _w21326_ ;
	wire _w21325_ ;
	wire _w21324_ ;
	wire _w21323_ ;
	wire _w21322_ ;
	wire _w21321_ ;
	wire _w21320_ ;
	wire _w21319_ ;
	wire _w21318_ ;
	wire _w21317_ ;
	wire _w21316_ ;
	wire _w21315_ ;
	wire _w21314_ ;
	wire _w21313_ ;
	wire _w21312_ ;
	wire _w21311_ ;
	wire _w21310_ ;
	wire _w21309_ ;
	wire _w21308_ ;
	wire _w21307_ ;
	wire _w21306_ ;
	wire _w21305_ ;
	wire _w21304_ ;
	wire _w21303_ ;
	wire _w21302_ ;
	wire _w21301_ ;
	wire _w21300_ ;
	wire _w21299_ ;
	wire _w21298_ ;
	wire _w21297_ ;
	wire _w21296_ ;
	wire _w21295_ ;
	wire _w21294_ ;
	wire _w21293_ ;
	wire _w21292_ ;
	wire _w21291_ ;
	wire _w21290_ ;
	wire _w21289_ ;
	wire _w21288_ ;
	wire _w21287_ ;
	wire _w21286_ ;
	wire _w21285_ ;
	wire _w21284_ ;
	wire _w21283_ ;
	wire _w21282_ ;
	wire _w21281_ ;
	wire _w21280_ ;
	wire _w21279_ ;
	wire _w21278_ ;
	wire _w21277_ ;
	wire _w21276_ ;
	wire _w21275_ ;
	wire _w21274_ ;
	wire _w21273_ ;
	wire _w21272_ ;
	wire _w21271_ ;
	wire _w21270_ ;
	wire _w21269_ ;
	wire _w21268_ ;
	wire _w21267_ ;
	wire _w21266_ ;
	wire _w21265_ ;
	wire _w21264_ ;
	wire _w21263_ ;
	wire _w21262_ ;
	wire _w21261_ ;
	wire _w21260_ ;
	wire _w21259_ ;
	wire _w21258_ ;
	wire _w21257_ ;
	wire _w21256_ ;
	wire _w21255_ ;
	wire _w21254_ ;
	wire _w21253_ ;
	wire _w21252_ ;
	wire _w21251_ ;
	wire _w21250_ ;
	wire _w21249_ ;
	wire _w21248_ ;
	wire _w21247_ ;
	wire _w21246_ ;
	wire _w21245_ ;
	wire _w21244_ ;
	wire _w21243_ ;
	wire _w21242_ ;
	wire _w21241_ ;
	wire _w21240_ ;
	wire _w21239_ ;
	wire _w21238_ ;
	wire _w21237_ ;
	wire _w21236_ ;
	wire _w21235_ ;
	wire _w21234_ ;
	wire _w21233_ ;
	wire _w21232_ ;
	wire _w21231_ ;
	wire _w21230_ ;
	wire _w21229_ ;
	wire _w21228_ ;
	wire _w21227_ ;
	wire _w21226_ ;
	wire _w21225_ ;
	wire _w21224_ ;
	wire _w21223_ ;
	wire _w21222_ ;
	wire _w21221_ ;
	wire _w21220_ ;
	wire _w21219_ ;
	wire _w21218_ ;
	wire _w21217_ ;
	wire _w21216_ ;
	wire _w21215_ ;
	wire _w21214_ ;
	wire _w21212_ ;
	wire _w21211_ ;
	wire _w21210_ ;
	wire _w21209_ ;
	wire _w21208_ ;
	wire _w21207_ ;
	wire _w21206_ ;
	wire _w21205_ ;
	wire _w21204_ ;
	wire _w21203_ ;
	wire _w21202_ ;
	wire _w21201_ ;
	wire _w21200_ ;
	wire _w21199_ ;
	wire _w21198_ ;
	wire _w21197_ ;
	wire _w21196_ ;
	wire _w21195_ ;
	wire _w21194_ ;
	wire _w21193_ ;
	wire _w21192_ ;
	wire _w21191_ ;
	wire _w21190_ ;
	wire _w21189_ ;
	wire _w21188_ ;
	wire _w21187_ ;
	wire _w21186_ ;
	wire _w21185_ ;
	wire _w21184_ ;
	wire _w21183_ ;
	wire _w21182_ ;
	wire _w21181_ ;
	wire _w21180_ ;
	wire _w21179_ ;
	wire _w21178_ ;
	wire _w21177_ ;
	wire _w21176_ ;
	wire _w21175_ ;
	wire _w21174_ ;
	wire _w21173_ ;
	wire _w21172_ ;
	wire _w21171_ ;
	wire _w21170_ ;
	wire _w21169_ ;
	wire _w21168_ ;
	wire _w21167_ ;
	wire _w21166_ ;
	wire _w21165_ ;
	wire _w21164_ ;
	wire _w21163_ ;
	wire _w21162_ ;
	wire _w21161_ ;
	wire _w21160_ ;
	wire _w21159_ ;
	wire _w21158_ ;
	wire _w21157_ ;
	wire _w21156_ ;
	wire _w21155_ ;
	wire _w21154_ ;
	wire _w21153_ ;
	wire _w21152_ ;
	wire _w21151_ ;
	wire _w21150_ ;
	wire _w21149_ ;
	wire _w21148_ ;
	wire _w21147_ ;
	wire _w21146_ ;
	wire _w21145_ ;
	wire _w21144_ ;
	wire _w21143_ ;
	wire _w21142_ ;
	wire _w21141_ ;
	wire _w21140_ ;
	wire _w21139_ ;
	wire _w21138_ ;
	wire _w21137_ ;
	wire _w21136_ ;
	wire _w21135_ ;
	wire _w21134_ ;
	wire _w21133_ ;
	wire _w21132_ ;
	wire _w21131_ ;
	wire _w21130_ ;
	wire _w21129_ ;
	wire _w21128_ ;
	wire _w21127_ ;
	wire _w21126_ ;
	wire _w21125_ ;
	wire _w21124_ ;
	wire _w21123_ ;
	wire _w21122_ ;
	wire _w21121_ ;
	wire _w21120_ ;
	wire _w21119_ ;
	wire _w21118_ ;
	wire _w21117_ ;
	wire _w21116_ ;
	wire _w21115_ ;
	wire _w21114_ ;
	wire _w21113_ ;
	wire _w21112_ ;
	wire _w21111_ ;
	wire _w21110_ ;
	wire _w21109_ ;
	wire _w21108_ ;
	wire _w21107_ ;
	wire _w21106_ ;
	wire _w21105_ ;
	wire _w21104_ ;
	wire _w21103_ ;
	wire _w21102_ ;
	wire _w21101_ ;
	wire _w21100_ ;
	wire _w21099_ ;
	wire _w21098_ ;
	wire _w21097_ ;
	wire _w21096_ ;
	wire _w21095_ ;
	wire _w21094_ ;
	wire _w21093_ ;
	wire _w21092_ ;
	wire _w21091_ ;
	wire _w21090_ ;
	wire _w21089_ ;
	wire _w21088_ ;
	wire _w21087_ ;
	wire _w21086_ ;
	wire _w21085_ ;
	wire _w21084_ ;
	wire _w21083_ ;
	wire _w21082_ ;
	wire _w21081_ ;
	wire _w21080_ ;
	wire _w21079_ ;
	wire _w21078_ ;
	wire _w21077_ ;
	wire _w21076_ ;
	wire _w21075_ ;
	wire _w21074_ ;
	wire _w21073_ ;
	wire _w21072_ ;
	wire _w21071_ ;
	wire _w21070_ ;
	wire _w21069_ ;
	wire _w21068_ ;
	wire _w21067_ ;
	wire _w21066_ ;
	wire _w21065_ ;
	wire _w21064_ ;
	wire _w21063_ ;
	wire _w21062_ ;
	wire _w21061_ ;
	wire _w21060_ ;
	wire _w21059_ ;
	wire _w21058_ ;
	wire _w21057_ ;
	wire _w21056_ ;
	wire _w21055_ ;
	wire _w21054_ ;
	wire _w21053_ ;
	wire _w21052_ ;
	wire _w21051_ ;
	wire _w21050_ ;
	wire _w21049_ ;
	wire _w21048_ ;
	wire _w21047_ ;
	wire _w21046_ ;
	wire _w21045_ ;
	wire _w21044_ ;
	wire _w21043_ ;
	wire _w21042_ ;
	wire _w21041_ ;
	wire _w21040_ ;
	wire _w21039_ ;
	wire _w21038_ ;
	wire _w21037_ ;
	wire _w21036_ ;
	wire _w21035_ ;
	wire _w21034_ ;
	wire _w21033_ ;
	wire _w21032_ ;
	wire _w21031_ ;
	wire _w21030_ ;
	wire _w21029_ ;
	wire _w21028_ ;
	wire _w21027_ ;
	wire _w21026_ ;
	wire _w21025_ ;
	wire _w21024_ ;
	wire _w21023_ ;
	wire _w21022_ ;
	wire _w21021_ ;
	wire _w21020_ ;
	wire _w21019_ ;
	wire _w21018_ ;
	wire _w21017_ ;
	wire _w21016_ ;
	wire _w21015_ ;
	wire _w21014_ ;
	wire _w21013_ ;
	wire _w21012_ ;
	wire _w21011_ ;
	wire _w21010_ ;
	wire _w21009_ ;
	wire _w21008_ ;
	wire _w21007_ ;
	wire _w21006_ ;
	wire _w21005_ ;
	wire _w21004_ ;
	wire _w21003_ ;
	wire _w21002_ ;
	wire _w21001_ ;
	wire _w21000_ ;
	wire _w20999_ ;
	wire _w20998_ ;
	wire _w20997_ ;
	wire _w20996_ ;
	wire _w20995_ ;
	wire _w20994_ ;
	wire _w20993_ ;
	wire _w20992_ ;
	wire _w20991_ ;
	wire _w20990_ ;
	wire _w20989_ ;
	wire _w20988_ ;
	wire _w20987_ ;
	wire _w20986_ ;
	wire _w20985_ ;
	wire _w20984_ ;
	wire _w20983_ ;
	wire _w20982_ ;
	wire _w20981_ ;
	wire _w20980_ ;
	wire _w20979_ ;
	wire _w20978_ ;
	wire _w20977_ ;
	wire _w20976_ ;
	wire _w20975_ ;
	wire _w20974_ ;
	wire _w20973_ ;
	wire _w20972_ ;
	wire _w20971_ ;
	wire _w20970_ ;
	wire _w20969_ ;
	wire _w20968_ ;
	wire _w20967_ ;
	wire _w20966_ ;
	wire _w20965_ ;
	wire _w20964_ ;
	wire _w20963_ ;
	wire _w20962_ ;
	wire _w20961_ ;
	wire _w20960_ ;
	wire _w20959_ ;
	wire _w20958_ ;
	wire _w20957_ ;
	wire _w20956_ ;
	wire _w20955_ ;
	wire _w20954_ ;
	wire _w20953_ ;
	wire _w20952_ ;
	wire _w20951_ ;
	wire _w20950_ ;
	wire _w20949_ ;
	wire _w20948_ ;
	wire _w20947_ ;
	wire _w20946_ ;
	wire _w20945_ ;
	wire _w20944_ ;
	wire _w20943_ ;
	wire _w20942_ ;
	wire _w20941_ ;
	wire _w20940_ ;
	wire _w20939_ ;
	wire _w20938_ ;
	wire _w20937_ ;
	wire _w20936_ ;
	wire _w20935_ ;
	wire _w20934_ ;
	wire _w20933_ ;
	wire _w20932_ ;
	wire _w20931_ ;
	wire _w20930_ ;
	wire _w20929_ ;
	wire _w20928_ ;
	wire _w20927_ ;
	wire _w20926_ ;
	wire _w20925_ ;
	wire _w20924_ ;
	wire _w20923_ ;
	wire _w20922_ ;
	wire _w20921_ ;
	wire _w20920_ ;
	wire _w20919_ ;
	wire _w20918_ ;
	wire _w20917_ ;
	wire _w20916_ ;
	wire _w20915_ ;
	wire _w20914_ ;
	wire _w20913_ ;
	wire _w20912_ ;
	wire _w20911_ ;
	wire _w20910_ ;
	wire _w20909_ ;
	wire _w20908_ ;
	wire _w20907_ ;
	wire _w20906_ ;
	wire _w20905_ ;
	wire _w20904_ ;
	wire _w20903_ ;
	wire _w20902_ ;
	wire _w20901_ ;
	wire _w20900_ ;
	wire _w20899_ ;
	wire _w20898_ ;
	wire _w20897_ ;
	wire _w20896_ ;
	wire _w20895_ ;
	wire _w20894_ ;
	wire _w20893_ ;
	wire _w20892_ ;
	wire _w20891_ ;
	wire _w20890_ ;
	wire _w20889_ ;
	wire _w20888_ ;
	wire _w20887_ ;
	wire _w20886_ ;
	wire _w20885_ ;
	wire _w20884_ ;
	wire _w20883_ ;
	wire _w20882_ ;
	wire _w20881_ ;
	wire _w20880_ ;
	wire _w20879_ ;
	wire _w20878_ ;
	wire _w20877_ ;
	wire _w20876_ ;
	wire _w20875_ ;
	wire _w20874_ ;
	wire _w20873_ ;
	wire _w20872_ ;
	wire _w20871_ ;
	wire _w20870_ ;
	wire _w20869_ ;
	wire _w20868_ ;
	wire _w20867_ ;
	wire _w20866_ ;
	wire _w20865_ ;
	wire _w20864_ ;
	wire _w20863_ ;
	wire _w20862_ ;
	wire _w20861_ ;
	wire _w20860_ ;
	wire _w20859_ ;
	wire _w20858_ ;
	wire _w20857_ ;
	wire _w20856_ ;
	wire _w20855_ ;
	wire _w20854_ ;
	wire _w20853_ ;
	wire _w20852_ ;
	wire _w20851_ ;
	wire _w20850_ ;
	wire _w20849_ ;
	wire _w20848_ ;
	wire _w20847_ ;
	wire _w20846_ ;
	wire _w20845_ ;
	wire _w20844_ ;
	wire _w20843_ ;
	wire _w20842_ ;
	wire _w20841_ ;
	wire _w20840_ ;
	wire _w20839_ ;
	wire _w20838_ ;
	wire _w20837_ ;
	wire _w20836_ ;
	wire _w20835_ ;
	wire _w20834_ ;
	wire _w20833_ ;
	wire _w20832_ ;
	wire _w20831_ ;
	wire _w20830_ ;
	wire _w20829_ ;
	wire _w20828_ ;
	wire _w20827_ ;
	wire _w20826_ ;
	wire _w20825_ ;
	wire _w20824_ ;
	wire _w20823_ ;
	wire _w20822_ ;
	wire _w20821_ ;
	wire _w20820_ ;
	wire _w20819_ ;
	wire _w20818_ ;
	wire _w20817_ ;
	wire _w20816_ ;
	wire _w20815_ ;
	wire _w20814_ ;
	wire _w20813_ ;
	wire _w20812_ ;
	wire _w20811_ ;
	wire _w20810_ ;
	wire _w20809_ ;
	wire _w20808_ ;
	wire _w20807_ ;
	wire _w20806_ ;
	wire _w20805_ ;
	wire _w20804_ ;
	wire _w20803_ ;
	wire _w20802_ ;
	wire _w20801_ ;
	wire _w20800_ ;
	wire _w20799_ ;
	wire _w20798_ ;
	wire _w20797_ ;
	wire _w20796_ ;
	wire _w20795_ ;
	wire _w20794_ ;
	wire _w20793_ ;
	wire _w20792_ ;
	wire _w20791_ ;
	wire _w20790_ ;
	wire _w20789_ ;
	wire _w20788_ ;
	wire _w20787_ ;
	wire _w20786_ ;
	wire _w15599_ ;
	wire _w15598_ ;
	wire _w15597_ ;
	wire _w15596_ ;
	wire _w15595_ ;
	wire _w15594_ ;
	wire _w15593_ ;
	wire _w15592_ ;
	wire _w15591_ ;
	wire _w15590_ ;
	wire _w15589_ ;
	wire _w15588_ ;
	wire _w15587_ ;
	wire _w15586_ ;
	wire _w15585_ ;
	wire _w15584_ ;
	wire _w15583_ ;
	wire _w15582_ ;
	wire _w15581_ ;
	wire _w15580_ ;
	wire _w15579_ ;
	wire _w15578_ ;
	wire _w15577_ ;
	wire _w15576_ ;
	wire _w15575_ ;
	wire _w15574_ ;
	wire _w15573_ ;
	wire _w15572_ ;
	wire _w15571_ ;
	wire _w15570_ ;
	wire _w15569_ ;
	wire _w15568_ ;
	wire _w15567_ ;
	wire _w15566_ ;
	wire _w15565_ ;
	wire _w15564_ ;
	wire _w15563_ ;
	wire _w15562_ ;
	wire _w15561_ ;
	wire _w15560_ ;
	wire _w15559_ ;
	wire _w15558_ ;
	wire _w15557_ ;
	wire _w15556_ ;
	wire _w15555_ ;
	wire _w15554_ ;
	wire _w15553_ ;
	wire _w15552_ ;
	wire _w15551_ ;
	wire _w15550_ ;
	wire _w15549_ ;
	wire _w15548_ ;
	wire _w15547_ ;
	wire _w15546_ ;
	wire _w15545_ ;
	wire _w15544_ ;
	wire _w15543_ ;
	wire _w15542_ ;
	wire _w15541_ ;
	wire _w15540_ ;
	wire _w15539_ ;
	wire _w15538_ ;
	wire _w15537_ ;
	wire _w15536_ ;
	wire _w15535_ ;
	wire _w15534_ ;
	wire _w15533_ ;
	wire _w15532_ ;
	wire _w15531_ ;
	wire _w15530_ ;
	wire _w15529_ ;
	wire _w15528_ ;
	wire _w15527_ ;
	wire _w15526_ ;
	wire _w15525_ ;
	wire _w15524_ ;
	wire _w15523_ ;
	wire _w15522_ ;
	wire _w15521_ ;
	wire _w15520_ ;
	wire _w15519_ ;
	wire _w15518_ ;
	wire _w15517_ ;
	wire _w15516_ ;
	wire _w15515_ ;
	wire _w15514_ ;
	wire _w15513_ ;
	wire _w15512_ ;
	wire _w15511_ ;
	wire _w15510_ ;
	wire _w15509_ ;
	wire _w15508_ ;
	wire _w15507_ ;
	wire _w15506_ ;
	wire _w15505_ ;
	wire _w15504_ ;
	wire _w15503_ ;
	wire _w15502_ ;
	wire _w15501_ ;
	wire _w15500_ ;
	wire _w15499_ ;
	wire _w15498_ ;
	wire _w15497_ ;
	wire _w15496_ ;
	wire _w15495_ ;
	wire _w15494_ ;
	wire _w15493_ ;
	wire _w15492_ ;
	wire _w15491_ ;
	wire _w15490_ ;
	wire _w15489_ ;
	wire _w15488_ ;
	wire _w15487_ ;
	wire _w15486_ ;
	wire _w15485_ ;
	wire _w15484_ ;
	wire _w15483_ ;
	wire _w15482_ ;
	wire _w15481_ ;
	wire _w15480_ ;
	wire _w15479_ ;
	wire _w15478_ ;
	wire _w15477_ ;
	wire _w15476_ ;
	wire _w15475_ ;
	wire _w15474_ ;
	wire _w15473_ ;
	wire _w15472_ ;
	wire _w15471_ ;
	wire _w15470_ ;
	wire _w15469_ ;
	wire _w15468_ ;
	wire _w15467_ ;
	wire _w15466_ ;
	wire _w15465_ ;
	wire _w15464_ ;
	wire _w15463_ ;
	wire _w15462_ ;
	wire _w15461_ ;
	wire _w15460_ ;
	wire _w15459_ ;
	wire _w15458_ ;
	wire _w15457_ ;
	wire _w15456_ ;
	wire _w15455_ ;
	wire _w15454_ ;
	wire _w15453_ ;
	wire _w15452_ ;
	wire _w15451_ ;
	wire _w15450_ ;
	wire _w15449_ ;
	wire _w15448_ ;
	wire _w15447_ ;
	wire _w15446_ ;
	wire _w15445_ ;
	wire _w15444_ ;
	wire _w15443_ ;
	wire _w15442_ ;
	wire _w15441_ ;
	wire _w15440_ ;
	wire _w15439_ ;
	wire _w15438_ ;
	wire _w15437_ ;
	wire _w15436_ ;
	wire _w15435_ ;
	wire _w15434_ ;
	wire _w15433_ ;
	wire _w15432_ ;
	wire _w15431_ ;
	wire _w15430_ ;
	wire _w15429_ ;
	wire _w15428_ ;
	wire _w15427_ ;
	wire _w15426_ ;
	wire _w15425_ ;
	wire _w15424_ ;
	wire _w15423_ ;
	wire _w15422_ ;
	wire _w15421_ ;
	wire _w15420_ ;
	wire _w15419_ ;
	wire _w15418_ ;
	wire _w15417_ ;
	wire _w15416_ ;
	wire _w15415_ ;
	wire _w15414_ ;
	wire _w15413_ ;
	wire _w15412_ ;
	wire _w15411_ ;
	wire _w15410_ ;
	wire _w15409_ ;
	wire _w15408_ ;
	wire _w15407_ ;
	wire _w15406_ ;
	wire _w15405_ ;
	wire _w15404_ ;
	wire _w15403_ ;
	wire _w15402_ ;
	wire _w15401_ ;
	wire _w15400_ ;
	wire _w15399_ ;
	wire _w15398_ ;
	wire _w15397_ ;
	wire _w15396_ ;
	wire _w15395_ ;
	wire _w15394_ ;
	wire _w15393_ ;
	wire _w15392_ ;
	wire _w15391_ ;
	wire _w15390_ ;
	wire _w15389_ ;
	wire _w15388_ ;
	wire _w15387_ ;
	wire _w15386_ ;
	wire _w15385_ ;
	wire _w15384_ ;
	wire _w15383_ ;
	wire _w15382_ ;
	wire _w15381_ ;
	wire _w15380_ ;
	wire _w15379_ ;
	wire _w15378_ ;
	wire _w15377_ ;
	wire _w15376_ ;
	wire _w15375_ ;
	wire _w15374_ ;
	wire _w15373_ ;
	wire _w15372_ ;
	wire _w15371_ ;
	wire _w15370_ ;
	wire _w15369_ ;
	wire _w15368_ ;
	wire _w15367_ ;
	wire _w15366_ ;
	wire _w15365_ ;
	wire _w15364_ ;
	wire _w15363_ ;
	wire _w15362_ ;
	wire _w15361_ ;
	wire _w15360_ ;
	wire _w15359_ ;
	wire _w15358_ ;
	wire _w15357_ ;
	wire _w15356_ ;
	wire _w15355_ ;
	wire _w15354_ ;
	wire _w15353_ ;
	wire _w15352_ ;
	wire _w15351_ ;
	wire _w15350_ ;
	wire _w15349_ ;
	wire _w15348_ ;
	wire _w15347_ ;
	wire _w15346_ ;
	wire _w15345_ ;
	wire _w15344_ ;
	wire _w15343_ ;
	wire _w15342_ ;
	wire _w15341_ ;
	wire _w15340_ ;
	wire _w15339_ ;
	wire _w15338_ ;
	wire _w15337_ ;
	wire _w15336_ ;
	wire _w15335_ ;
	wire _w15334_ ;
	wire _w15333_ ;
	wire _w15332_ ;
	wire _w15331_ ;
	wire _w15330_ ;
	wire _w15329_ ;
	wire _w15328_ ;
	wire _w15327_ ;
	wire _w15326_ ;
	wire _w15325_ ;
	wire _w15324_ ;
	wire _w15323_ ;
	wire _w15322_ ;
	wire _w15321_ ;
	wire _w15320_ ;
	wire _w15319_ ;
	wire _w15318_ ;
	wire _w15317_ ;
	wire _w15316_ ;
	wire _w15315_ ;
	wire _w15314_ ;
	wire _w15313_ ;
	wire _w15312_ ;
	wire _w15311_ ;
	wire _w15310_ ;
	wire _w15309_ ;
	wire _w15308_ ;
	wire _w15307_ ;
	wire _w15306_ ;
	wire _w15305_ ;
	wire _w15304_ ;
	wire _w15303_ ;
	wire _w15302_ ;
	wire _w15301_ ;
	wire _w15300_ ;
	wire _w15299_ ;
	wire _w15298_ ;
	wire _w15297_ ;
	wire _w15296_ ;
	wire _w15295_ ;
	wire _w15294_ ;
	wire _w15293_ ;
	wire _w15292_ ;
	wire _w15291_ ;
	wire _w15290_ ;
	wire _w15289_ ;
	wire _w15288_ ;
	wire _w15287_ ;
	wire _w15286_ ;
	wire _w15285_ ;
	wire _w15284_ ;
	wire _w15283_ ;
	wire _w15282_ ;
	wire _w15281_ ;
	wire _w15280_ ;
	wire _w15279_ ;
	wire _w15278_ ;
	wire _w15277_ ;
	wire _w15276_ ;
	wire _w15275_ ;
	wire _w15274_ ;
	wire _w15273_ ;
	wire _w15272_ ;
	wire _w15271_ ;
	wire _w15270_ ;
	wire _w15269_ ;
	wire _w15268_ ;
	wire _w15267_ ;
	wire _w15266_ ;
	wire _w15265_ ;
	wire _w15264_ ;
	wire _w15263_ ;
	wire _w15262_ ;
	wire _w15261_ ;
	wire _w15260_ ;
	wire _w15259_ ;
	wire _w15258_ ;
	wire _w15257_ ;
	wire _w15256_ ;
	wire _w15255_ ;
	wire _w15254_ ;
	wire _w15253_ ;
	wire _w15252_ ;
	wire _w15251_ ;
	wire _w15250_ ;
	wire _w15249_ ;
	wire _w15248_ ;
	wire _w15247_ ;
	wire _w15246_ ;
	wire _w15245_ ;
	wire _w15244_ ;
	wire _w15243_ ;
	wire _w15242_ ;
	wire _w15241_ ;
	wire _w15240_ ;
	wire _w15239_ ;
	wire _w15238_ ;
	wire _w15237_ ;
	wire _w15236_ ;
	wire _w15235_ ;
	wire _w15234_ ;
	wire _w15233_ ;
	wire _w15232_ ;
	wire _w15231_ ;
	wire _w15230_ ;
	wire _w15229_ ;
	wire _w15228_ ;
	wire _w15227_ ;
	wire _w15226_ ;
	wire _w15225_ ;
	wire _w15224_ ;
	wire _w15223_ ;
	wire _w15222_ ;
	wire _w15221_ ;
	wire _w15220_ ;
	wire _w15219_ ;
	wire _w15218_ ;
	wire _w15217_ ;
	wire _w15216_ ;
	wire _w15215_ ;
	wire _w15214_ ;
	wire _w15213_ ;
	wire _w15212_ ;
	wire _w15211_ ;
	wire _w15210_ ;
	wire _w15209_ ;
	wire _w15208_ ;
	wire _w15207_ ;
	wire _w15206_ ;
	wire _w15205_ ;
	wire _w15204_ ;
	wire _w15203_ ;
	wire _w15202_ ;
	wire _w15201_ ;
	wire _w15200_ ;
	wire _w15199_ ;
	wire _w15198_ ;
	wire _w15197_ ;
	wire _w15196_ ;
	wire _w15195_ ;
	wire _w15194_ ;
	wire _w15193_ ;
	wire _w15192_ ;
	wire _w15191_ ;
	wire _w15190_ ;
	wire _w15189_ ;
	wire _w15188_ ;
	wire _w15187_ ;
	wire _w15186_ ;
	wire _w15185_ ;
	wire _w15184_ ;
	wire _w15183_ ;
	wire _w15182_ ;
	wire _w15181_ ;
	wire _w15180_ ;
	wire _w15179_ ;
	wire _w15178_ ;
	wire _w15177_ ;
	wire _w15176_ ;
	wire _w15175_ ;
	wire _w15174_ ;
	wire _w15173_ ;
	wire _w15172_ ;
	wire _w15171_ ;
	wire _w15170_ ;
	wire _w15169_ ;
	wire _w15168_ ;
	wire _w15167_ ;
	wire _w15166_ ;
	wire _w15165_ ;
	wire _w15164_ ;
	wire _w15163_ ;
	wire _w15162_ ;
	wire _w15161_ ;
	wire _w15160_ ;
	wire _w15159_ ;
	wire _w15158_ ;
	wire _w15157_ ;
	wire _w15156_ ;
	wire _w15155_ ;
	wire _w15154_ ;
	wire _w15153_ ;
	wire _w15152_ ;
	wire _w15151_ ;
	wire _w15150_ ;
	wire _w15149_ ;
	wire _w15148_ ;
	wire _w15147_ ;
	wire _w15146_ ;
	wire _w15145_ ;
	wire _w15144_ ;
	wire _w15143_ ;
	wire _w15142_ ;
	wire _w15141_ ;
	wire _w15140_ ;
	wire _w15139_ ;
	wire _w15138_ ;
	wire _w15137_ ;
	wire _w15136_ ;
	wire _w15135_ ;
	wire _w15134_ ;
	wire _w15133_ ;
	wire _w15132_ ;
	wire _w15131_ ;
	wire _w15130_ ;
	wire _w15129_ ;
	wire _w15128_ ;
	wire _w15127_ ;
	wire _w15126_ ;
	wire _w15125_ ;
	wire _w15124_ ;
	wire _w15123_ ;
	wire _w15122_ ;
	wire _w15121_ ;
	wire _w15120_ ;
	wire _w15119_ ;
	wire _w15118_ ;
	wire _w15117_ ;
	wire _w15116_ ;
	wire _w15115_ ;
	wire _w15114_ ;
	wire _w15113_ ;
	wire _w15112_ ;
	wire _w15111_ ;
	wire _w15110_ ;
	wire _w15109_ ;
	wire _w15108_ ;
	wire _w15107_ ;
	wire _w15106_ ;
	wire _w15105_ ;
	wire _w15104_ ;
	wire _w15103_ ;
	wire _w15102_ ;
	wire _w15101_ ;
	wire _w15100_ ;
	wire _w15099_ ;
	wire _w15098_ ;
	wire _w15097_ ;
	wire _w15096_ ;
	wire _w15095_ ;
	wire _w15094_ ;
	wire _w15093_ ;
	wire _w15092_ ;
	wire _w15091_ ;
	wire _w15090_ ;
	wire _w15089_ ;
	wire _w15088_ ;
	wire _w15087_ ;
	wire _w15086_ ;
	wire _w15085_ ;
	wire _w15084_ ;
	wire _w15083_ ;
	wire _w15082_ ;
	wire _w15081_ ;
	wire _w15080_ ;
	wire _w15079_ ;
	wire _w15078_ ;
	wire _w15077_ ;
	wire _w15076_ ;
	wire _w15075_ ;
	wire _w15074_ ;
	wire _w15073_ ;
	wire _w15072_ ;
	wire _w15071_ ;
	wire _w15070_ ;
	wire _w15069_ ;
	wire _w15068_ ;
	wire _w15067_ ;
	wire _w15066_ ;
	wire _w15065_ ;
	wire _w15064_ ;
	wire _w15063_ ;
	wire _w15062_ ;
	wire _w15061_ ;
	wire _w15060_ ;
	wire _w15059_ ;
	wire _w15058_ ;
	wire _w15057_ ;
	wire _w15056_ ;
	wire _w15055_ ;
	wire _w15054_ ;
	wire _w15053_ ;
	wire _w15052_ ;
	wire _w15051_ ;
	wire _w15050_ ;
	wire _w15049_ ;
	wire _w15048_ ;
	wire _w15047_ ;
	wire _w15046_ ;
	wire _w15045_ ;
	wire _w15044_ ;
	wire _w15043_ ;
	wire _w15042_ ;
	wire _w15041_ ;
	wire _w15040_ ;
	wire _w15039_ ;
	wire _w15038_ ;
	wire _w15037_ ;
	wire _w15036_ ;
	wire _w15035_ ;
	wire _w15034_ ;
	wire _w15033_ ;
	wire _w15032_ ;
	wire _w15031_ ;
	wire _w15030_ ;
	wire _w15029_ ;
	wire _w15028_ ;
	wire _w15027_ ;
	wire _w15026_ ;
	wire _w15025_ ;
	wire _w15024_ ;
	wire _w15023_ ;
	wire _w15022_ ;
	wire _w15021_ ;
	wire _w15020_ ;
	wire _w15019_ ;
	wire _w15018_ ;
	wire _w15017_ ;
	wire _w15016_ ;
	wire _w15015_ ;
	wire _w15014_ ;
	wire _w15013_ ;
	wire _w15012_ ;
	wire _w15011_ ;
	wire _w15010_ ;
	wire _w15009_ ;
	wire _w15008_ ;
	wire _w15007_ ;
	wire _w15006_ ;
	wire _w15005_ ;
	wire _w15004_ ;
	wire _w15003_ ;
	wire _w15002_ ;
	wire _w15001_ ;
	wire _w15000_ ;
	wire _w14999_ ;
	wire _w14998_ ;
	wire _w14997_ ;
	wire _w14996_ ;
	wire _w14995_ ;
	wire _w14994_ ;
	wire _w14993_ ;
	wire _w14992_ ;
	wire _w14991_ ;
	wire _w14990_ ;
	wire _w14989_ ;
	wire _w14988_ ;
	wire _w14987_ ;
	wire _w14986_ ;
	wire _w14985_ ;
	wire _w14984_ ;
	wire _w14983_ ;
	wire _w14982_ ;
	wire _w14981_ ;
	wire _w14980_ ;
	wire _w14979_ ;
	wire _w14978_ ;
	wire _w14977_ ;
	wire _w14976_ ;
	wire _w14975_ ;
	wire _w14974_ ;
	wire _w14973_ ;
	wire _w14972_ ;
	wire _w14971_ ;
	wire _w14970_ ;
	wire _w14969_ ;
	wire _w14968_ ;
	wire _w14967_ ;
	wire _w14966_ ;
	wire _w14965_ ;
	wire _w14964_ ;
	wire _w14963_ ;
	wire _w14962_ ;
	wire _w14961_ ;
	wire _w14960_ ;
	wire _w14959_ ;
	wire _w14958_ ;
	wire _w14957_ ;
	wire _w14956_ ;
	wire _w14955_ ;
	wire _w14954_ ;
	wire _w14953_ ;
	wire _w14952_ ;
	wire _w14951_ ;
	wire _w14950_ ;
	wire _w14949_ ;
	wire _w14948_ ;
	wire _w14947_ ;
	wire _w14946_ ;
	wire _w14945_ ;
	wire _w14944_ ;
	wire _w14943_ ;
	wire _w14942_ ;
	wire _w14941_ ;
	wire _w14940_ ;
	wire _w14939_ ;
	wire _w14938_ ;
	wire _w14937_ ;
	wire _w14936_ ;
	wire _w14935_ ;
	wire _w14934_ ;
	wire _w14933_ ;
	wire _w14932_ ;
	wire _w14931_ ;
	wire _w14930_ ;
	wire _w14929_ ;
	wire _w14928_ ;
	wire _w14927_ ;
	wire _w14926_ ;
	wire _w14925_ ;
	wire _w14924_ ;
	wire _w14923_ ;
	wire _w14922_ ;
	wire _w14921_ ;
	wire _w14920_ ;
	wire _w14919_ ;
	wire _w14918_ ;
	wire _w14917_ ;
	wire _w14916_ ;
	wire _w14915_ ;
	wire _w14914_ ;
	wire _w14913_ ;
	wire _w14912_ ;
	wire _w14911_ ;
	wire _w14910_ ;
	wire _w14909_ ;
	wire _w14908_ ;
	wire _w14907_ ;
	wire _w14906_ ;
	wire _w14905_ ;
	wire _w14904_ ;
	wire _w14903_ ;
	wire _w14902_ ;
	wire _w14901_ ;
	wire _w14900_ ;
	wire _w14899_ ;
	wire _w14898_ ;
	wire _w14897_ ;
	wire _w14896_ ;
	wire _w14895_ ;
	wire _w14894_ ;
	wire _w14893_ ;
	wire _w14892_ ;
	wire _w14891_ ;
	wire _w14890_ ;
	wire _w14889_ ;
	wire _w14888_ ;
	wire _w14887_ ;
	wire _w14886_ ;
	wire _w14885_ ;
	wire _w14884_ ;
	wire _w14883_ ;
	wire _w14882_ ;
	wire _w14881_ ;
	wire _w14880_ ;
	wire _w14879_ ;
	wire _w14878_ ;
	wire _w14877_ ;
	wire _w14876_ ;
	wire _w14875_ ;
	wire _w14874_ ;
	wire _w14873_ ;
	wire _w14872_ ;
	wire _w14871_ ;
	wire _w14870_ ;
	wire _w14869_ ;
	wire _w14868_ ;
	wire _w14867_ ;
	wire _w14866_ ;
	wire _w14865_ ;
	wire _w14864_ ;
	wire _w14863_ ;
	wire _w14862_ ;
	wire _w14861_ ;
	wire _w14860_ ;
	wire _w14859_ ;
	wire _w14858_ ;
	wire _w14857_ ;
	wire _w14856_ ;
	wire _w14855_ ;
	wire _w14854_ ;
	wire _w14853_ ;
	wire _w14852_ ;
	wire _w14851_ ;
	wire _w14850_ ;
	wire _w14849_ ;
	wire _w14848_ ;
	wire _w14847_ ;
	wire _w14846_ ;
	wire _w14845_ ;
	wire _w14844_ ;
	wire _w14843_ ;
	wire _w14842_ ;
	wire _w14841_ ;
	wire _w14840_ ;
	wire _w14839_ ;
	wire _w14838_ ;
	wire _w14837_ ;
	wire _w14836_ ;
	wire _w14835_ ;
	wire _w14834_ ;
	wire _w14833_ ;
	wire _w14832_ ;
	wire _w14831_ ;
	wire _w14830_ ;
	wire _w14829_ ;
	wire _w14828_ ;
	wire _w14827_ ;
	wire _w14826_ ;
	wire _w14825_ ;
	wire _w14824_ ;
	wire _w14823_ ;
	wire _w14822_ ;
	wire _w14821_ ;
	wire _w14820_ ;
	wire _w14819_ ;
	wire _w14818_ ;
	wire _w14817_ ;
	wire _w14816_ ;
	wire _w14815_ ;
	wire _w14814_ ;
	wire _w14813_ ;
	wire _w14812_ ;
	wire _w14811_ ;
	wire _w14810_ ;
	wire _w14809_ ;
	wire _w14808_ ;
	wire _w14807_ ;
	wire _w14806_ ;
	wire _w14805_ ;
	wire _w14804_ ;
	wire _w14803_ ;
	wire _w14802_ ;
	wire _w14801_ ;
	wire _w14800_ ;
	wire _w14799_ ;
	wire _w14798_ ;
	wire _w14797_ ;
	wire _w14796_ ;
	wire _w14795_ ;
	wire _w14794_ ;
	wire _w14793_ ;
	wire _w14792_ ;
	wire _w14791_ ;
	wire _w14790_ ;
	wire _w14789_ ;
	wire _w14788_ ;
	wire _w14787_ ;
	wire _w14786_ ;
	wire _w14785_ ;
	wire _w14784_ ;
	wire _w14783_ ;
	wire _w14782_ ;
	wire _w14781_ ;
	wire _w14780_ ;
	wire _w14779_ ;
	wire _w14778_ ;
	wire _w14777_ ;
	wire _w14776_ ;
	wire _w14775_ ;
	wire _w14774_ ;
	wire _w14773_ ;
	wire _w14772_ ;
	wire _w14771_ ;
	wire _w14770_ ;
	wire _w14769_ ;
	wire _w14768_ ;
	wire _w14767_ ;
	wire _w14766_ ;
	wire _w14765_ ;
	wire _w14764_ ;
	wire _w14763_ ;
	wire _w14762_ ;
	wire _w14761_ ;
	wire _w14760_ ;
	wire _w14759_ ;
	wire _w14758_ ;
	wire _w14757_ ;
	wire _w14756_ ;
	wire _w14755_ ;
	wire _w14754_ ;
	wire _w14753_ ;
	wire _w14752_ ;
	wire _w14751_ ;
	wire _w14750_ ;
	wire _w14749_ ;
	wire _w14748_ ;
	wire _w14747_ ;
	wire _w14746_ ;
	wire _w14745_ ;
	wire _w14744_ ;
	wire _w14743_ ;
	wire _w14742_ ;
	wire _w14741_ ;
	wire _w14740_ ;
	wire _w14739_ ;
	wire _w14738_ ;
	wire _w14737_ ;
	wire _w14736_ ;
	wire _w14735_ ;
	wire _w14734_ ;
	wire _w14733_ ;
	wire _w14732_ ;
	wire _w14731_ ;
	wire _w14730_ ;
	wire _w14729_ ;
	wire _w14728_ ;
	wire _w14727_ ;
	wire _w14726_ ;
	wire _w14725_ ;
	wire _w14724_ ;
	wire _w14723_ ;
	wire _w14722_ ;
	wire _w14721_ ;
	wire _w14720_ ;
	wire _w14719_ ;
	wire _w14718_ ;
	wire _w14717_ ;
	wire _w14716_ ;
	wire _w14715_ ;
	wire _w14714_ ;
	wire _w14713_ ;
	wire _w14712_ ;
	wire _w14711_ ;
	wire _w14710_ ;
	wire _w14709_ ;
	wire _w14708_ ;
	wire _w14707_ ;
	wire _w14706_ ;
	wire _w14705_ ;
	wire _w14704_ ;
	wire _w14703_ ;
	wire _w14702_ ;
	wire _w14701_ ;
	wire _w14700_ ;
	wire _w14699_ ;
	wire _w14698_ ;
	wire _w14697_ ;
	wire _w14696_ ;
	wire _w14695_ ;
	wire _w14694_ ;
	wire _w14693_ ;
	wire _w14692_ ;
	wire _w14691_ ;
	wire _w14690_ ;
	wire _w14689_ ;
	wire _w14688_ ;
	wire _w14687_ ;
	wire _w14686_ ;
	wire _w14685_ ;
	wire _w14684_ ;
	wire _w14683_ ;
	wire _w14682_ ;
	wire _w14681_ ;
	wire _w14680_ ;
	wire _w14679_ ;
	wire _w14678_ ;
	wire _w14677_ ;
	wire _w14676_ ;
	wire _w14675_ ;
	wire _w14674_ ;
	wire _w14673_ ;
	wire _w14672_ ;
	wire _w14671_ ;
	wire _w14670_ ;
	wire _w14669_ ;
	wire _w14668_ ;
	wire _w14667_ ;
	wire _w14666_ ;
	wire _w14665_ ;
	wire _w14664_ ;
	wire _w14663_ ;
	wire _w14662_ ;
	wire _w14661_ ;
	wire _w14660_ ;
	wire _w14659_ ;
	wire _w14658_ ;
	wire _w14657_ ;
	wire _w14656_ ;
	wire _w14655_ ;
	wire _w14654_ ;
	wire _w14653_ ;
	wire _w14652_ ;
	wire _w14651_ ;
	wire _w14650_ ;
	wire _w14649_ ;
	wire _w14648_ ;
	wire _w14647_ ;
	wire _w14646_ ;
	wire _w14645_ ;
	wire _w14644_ ;
	wire _w14643_ ;
	wire _w14642_ ;
	wire _w14641_ ;
	wire _w14640_ ;
	wire _w14639_ ;
	wire _w14638_ ;
	wire _w14637_ ;
	wire _w14636_ ;
	wire _w14635_ ;
	wire _w14634_ ;
	wire _w14633_ ;
	wire _w14632_ ;
	wire _w14631_ ;
	wire _w14630_ ;
	wire _w14629_ ;
	wire _w14628_ ;
	wire _w14627_ ;
	wire _w14626_ ;
	wire _w14625_ ;
	wire _w14624_ ;
	wire _w14623_ ;
	wire _w14622_ ;
	wire _w14621_ ;
	wire _w14620_ ;
	wire _w14619_ ;
	wire _w14618_ ;
	wire _w14617_ ;
	wire _w14616_ ;
	wire _w14615_ ;
	wire _w14614_ ;
	wire _w14613_ ;
	wire _w14612_ ;
	wire _w14611_ ;
	wire _w14610_ ;
	wire _w14609_ ;
	wire _w14608_ ;
	wire _w14607_ ;
	wire _w14606_ ;
	wire _w14605_ ;
	wire _w14604_ ;
	wire _w14603_ ;
	wire _w14602_ ;
	wire _w14601_ ;
	wire _w14600_ ;
	wire _w14599_ ;
	wire _w14598_ ;
	wire _w14597_ ;
	wire _w14596_ ;
	wire _w14595_ ;
	wire _w14594_ ;
	wire _w14593_ ;
	wire _w14592_ ;
	wire _w14591_ ;
	wire _w14590_ ;
	wire _w14589_ ;
	wire _w14588_ ;
	wire _w14587_ ;
	wire _w14586_ ;
	wire _w14585_ ;
	wire _w14584_ ;
	wire _w14583_ ;
	wire _w14582_ ;
	wire _w14581_ ;
	wire _w14580_ ;
	wire _w14579_ ;
	wire _w14578_ ;
	wire _w14577_ ;
	wire _w14576_ ;
	wire _w14575_ ;
	wire _w14574_ ;
	wire _w14573_ ;
	wire _w14572_ ;
	wire _w14571_ ;
	wire _w14570_ ;
	wire _w14569_ ;
	wire _w14568_ ;
	wire _w14567_ ;
	wire _w14566_ ;
	wire _w14565_ ;
	wire _w14564_ ;
	wire _w14563_ ;
	wire _w14562_ ;
	wire _w14561_ ;
	wire _w14560_ ;
	wire _w14559_ ;
	wire _w14558_ ;
	wire _w14557_ ;
	wire _w14556_ ;
	wire _w14555_ ;
	wire _w14554_ ;
	wire _w14553_ ;
	wire _w14552_ ;
	wire _w14551_ ;
	wire _w14550_ ;
	wire _w14549_ ;
	wire _w14548_ ;
	wire _w14547_ ;
	wire _w14546_ ;
	wire _w14545_ ;
	wire _w14544_ ;
	wire _w14543_ ;
	wire _w14542_ ;
	wire _w14541_ ;
	wire _w14540_ ;
	wire _w14539_ ;
	wire _w14538_ ;
	wire _w14537_ ;
	wire _w14536_ ;
	wire _w14535_ ;
	wire _w14534_ ;
	wire _w14533_ ;
	wire _w14532_ ;
	wire _w14531_ ;
	wire _w14530_ ;
	wire _w14529_ ;
	wire _w14528_ ;
	wire _w14527_ ;
	wire _w14526_ ;
	wire _w14525_ ;
	wire _w14524_ ;
	wire _w14523_ ;
	wire _w14522_ ;
	wire _w14521_ ;
	wire _w14520_ ;
	wire _w14519_ ;
	wire _w14518_ ;
	wire _w14517_ ;
	wire _w14516_ ;
	wire _w14515_ ;
	wire _w14514_ ;
	wire _w14513_ ;
	wire _w14512_ ;
	wire _w14511_ ;
	wire _w14510_ ;
	wire _w14509_ ;
	wire _w14508_ ;
	wire _w14507_ ;
	wire _w14506_ ;
	wire _w14505_ ;
	wire _w14504_ ;
	wire _w14503_ ;
	wire _w14502_ ;
	wire _w14501_ ;
	wire _w14500_ ;
	wire _w14499_ ;
	wire _w14498_ ;
	wire _w14497_ ;
	wire _w14496_ ;
	wire _w14495_ ;
	wire _w14494_ ;
	wire _w14493_ ;
	wire _w14492_ ;
	wire _w14491_ ;
	wire _w14490_ ;
	wire _w14489_ ;
	wire _w14488_ ;
	wire _w14487_ ;
	wire _w14486_ ;
	wire _w14485_ ;
	wire _w14484_ ;
	wire _w14483_ ;
	wire _w14482_ ;
	wire _w14481_ ;
	wire _w14480_ ;
	wire _w14479_ ;
	wire _w14478_ ;
	wire _w14477_ ;
	wire _w14476_ ;
	wire _w14475_ ;
	wire _w14474_ ;
	wire _w14473_ ;
	wire _w14472_ ;
	wire _w14471_ ;
	wire _w14470_ ;
	wire _w14469_ ;
	wire _w14468_ ;
	wire _w14467_ ;
	wire _w14466_ ;
	wire _w14465_ ;
	wire _w14464_ ;
	wire _w14463_ ;
	wire _w14462_ ;
	wire _w14461_ ;
	wire _w14460_ ;
	wire _w14459_ ;
	wire _w14458_ ;
	wire _w14457_ ;
	wire _w14456_ ;
	wire _w14455_ ;
	wire _w14454_ ;
	wire _w14453_ ;
	wire _w14452_ ;
	wire _w14451_ ;
	wire _w14450_ ;
	wire _w14449_ ;
	wire _w14448_ ;
	wire _w14447_ ;
	wire _w14446_ ;
	wire _w14445_ ;
	wire _w14444_ ;
	wire _w14443_ ;
	wire _w14442_ ;
	wire _w14441_ ;
	wire _w14440_ ;
	wire _w14439_ ;
	wire _w14438_ ;
	wire _w14437_ ;
	wire _w14436_ ;
	wire _w14435_ ;
	wire _w14434_ ;
	wire _w14433_ ;
	wire _w14432_ ;
	wire _w14431_ ;
	wire _w14430_ ;
	wire _w14429_ ;
	wire _w14428_ ;
	wire _w14427_ ;
	wire _w14426_ ;
	wire _w14425_ ;
	wire _w14424_ ;
	wire _w14423_ ;
	wire _w14422_ ;
	wire _w14421_ ;
	wire _w14420_ ;
	wire _w14419_ ;
	wire _w14418_ ;
	wire _w14417_ ;
	wire _w14416_ ;
	wire _w14415_ ;
	wire _w14414_ ;
	wire _w14413_ ;
	wire _w14412_ ;
	wire _w14411_ ;
	wire _w14410_ ;
	wire _w14409_ ;
	wire _w14408_ ;
	wire _w14407_ ;
	wire _w14406_ ;
	wire _w14405_ ;
	wire _w14404_ ;
	wire _w14403_ ;
	wire _w14402_ ;
	wire _w14401_ ;
	wire _w14400_ ;
	wire _w14399_ ;
	wire _w14398_ ;
	wire _w14397_ ;
	wire _w14396_ ;
	wire _w14395_ ;
	wire _w14394_ ;
	wire _w14393_ ;
	wire _w14392_ ;
	wire _w14391_ ;
	wire _w14390_ ;
	wire _w14389_ ;
	wire _w14388_ ;
	wire _w14387_ ;
	wire _w14386_ ;
	wire _w14385_ ;
	wire _w14384_ ;
	wire _w14383_ ;
	wire _w14382_ ;
	wire _w14381_ ;
	wire _w14380_ ;
	wire _w14379_ ;
	wire _w14378_ ;
	wire _w14377_ ;
	wire _w14376_ ;
	wire _w14375_ ;
	wire _w14374_ ;
	wire _w14373_ ;
	wire _w14372_ ;
	wire _w14371_ ;
	wire _w14370_ ;
	wire _w14369_ ;
	wire _w14368_ ;
	wire _w14367_ ;
	wire _w14366_ ;
	wire _w14365_ ;
	wire _w14364_ ;
	wire _w14363_ ;
	wire _w14362_ ;
	wire _w14361_ ;
	wire _w14360_ ;
	wire _w14359_ ;
	wire _w14358_ ;
	wire _w14357_ ;
	wire _w14356_ ;
	wire _w14355_ ;
	wire _w14354_ ;
	wire _w14353_ ;
	wire _w14352_ ;
	wire _w14351_ ;
	wire _w14350_ ;
	wire _w14349_ ;
	wire _w14348_ ;
	wire _w14347_ ;
	wire _w14346_ ;
	wire _w14345_ ;
	wire _w14344_ ;
	wire _w14343_ ;
	wire _w14342_ ;
	wire _w14341_ ;
	wire _w14340_ ;
	wire _w14339_ ;
	wire _w14338_ ;
	wire _w14337_ ;
	wire _w14336_ ;
	wire _w14335_ ;
	wire _w14334_ ;
	wire _w14333_ ;
	wire _w14332_ ;
	wire _w14331_ ;
	wire _w14330_ ;
	wire _w14329_ ;
	wire _w14328_ ;
	wire _w14327_ ;
	wire _w14326_ ;
	wire _w14325_ ;
	wire _w14324_ ;
	wire _w14323_ ;
	wire _w14322_ ;
	wire _w14321_ ;
	wire _w14320_ ;
	wire _w14319_ ;
	wire _w14318_ ;
	wire _w14317_ ;
	wire _w14316_ ;
	wire _w14315_ ;
	wire _w14314_ ;
	wire _w14313_ ;
	wire _w14312_ ;
	wire _w14311_ ;
	wire _w14310_ ;
	wire _w14309_ ;
	wire _w14308_ ;
	wire _w14307_ ;
	wire _w14306_ ;
	wire _w14305_ ;
	wire _w14304_ ;
	wire _w14303_ ;
	wire _w14302_ ;
	wire _w14301_ ;
	wire _w14300_ ;
	wire _w14299_ ;
	wire _w14298_ ;
	wire _w14297_ ;
	wire _w14296_ ;
	wire _w14295_ ;
	wire _w14294_ ;
	wire _w14293_ ;
	wire _w14292_ ;
	wire _w14291_ ;
	wire _w14290_ ;
	wire _w14289_ ;
	wire _w14288_ ;
	wire _w14287_ ;
	wire _w14286_ ;
	wire _w14285_ ;
	wire _w14284_ ;
	wire _w14283_ ;
	wire _w14282_ ;
	wire _w14281_ ;
	wire _w14280_ ;
	wire _w14279_ ;
	wire _w14278_ ;
	wire _w14277_ ;
	wire _w14276_ ;
	wire _w14275_ ;
	wire _w14274_ ;
	wire _w14273_ ;
	wire _w14272_ ;
	wire _w14271_ ;
	wire _w14270_ ;
	wire _w14269_ ;
	wire _w14268_ ;
	wire _w14267_ ;
	wire _w14266_ ;
	wire _w14265_ ;
	wire _w14264_ ;
	wire _w14263_ ;
	wire _w14262_ ;
	wire _w14261_ ;
	wire _w14260_ ;
	wire _w14259_ ;
	wire _w14258_ ;
	wire _w14257_ ;
	wire _w14256_ ;
	wire _w14255_ ;
	wire _w14254_ ;
	wire _w14253_ ;
	wire _w14252_ ;
	wire _w14251_ ;
	wire _w14250_ ;
	wire _w14249_ ;
	wire _w14248_ ;
	wire _w14247_ ;
	wire _w14246_ ;
	wire _w14245_ ;
	wire _w14244_ ;
	wire _w14243_ ;
	wire _w14242_ ;
	wire _w14241_ ;
	wire _w14240_ ;
	wire _w14239_ ;
	wire _w14238_ ;
	wire _w14237_ ;
	wire _w14236_ ;
	wire _w14235_ ;
	wire _w14234_ ;
	wire _w14233_ ;
	wire _w14232_ ;
	wire _w14231_ ;
	wire _w14230_ ;
	wire _w14229_ ;
	wire _w14228_ ;
	wire _w14227_ ;
	wire _w14226_ ;
	wire _w14225_ ;
	wire _w14224_ ;
	wire _w14223_ ;
	wire _w14222_ ;
	wire _w14221_ ;
	wire _w14220_ ;
	wire _w14219_ ;
	wire _w14218_ ;
	wire _w14217_ ;
	wire _w14216_ ;
	wire _w14215_ ;
	wire _w14214_ ;
	wire _w14213_ ;
	wire _w14212_ ;
	wire _w14211_ ;
	wire _w14210_ ;
	wire _w14209_ ;
	wire _w14208_ ;
	wire _w14207_ ;
	wire _w14206_ ;
	wire _w14205_ ;
	wire _w14204_ ;
	wire _w14203_ ;
	wire _w14202_ ;
	wire _w14201_ ;
	wire _w14200_ ;
	wire _w14199_ ;
	wire _w14198_ ;
	wire _w14197_ ;
	wire _w14196_ ;
	wire _w14195_ ;
	wire _w14194_ ;
	wire _w14193_ ;
	wire _w14192_ ;
	wire _w14191_ ;
	wire _w14190_ ;
	wire _w14189_ ;
	wire _w14188_ ;
	wire _w14187_ ;
	wire _w14186_ ;
	wire _w14185_ ;
	wire _w14184_ ;
	wire _w14183_ ;
	wire _w14182_ ;
	wire _w14181_ ;
	wire _w14180_ ;
	wire _w14179_ ;
	wire _w14178_ ;
	wire _w14177_ ;
	wire _w14176_ ;
	wire _w14175_ ;
	wire _w14174_ ;
	wire _w14173_ ;
	wire _w14172_ ;
	wire _w14171_ ;
	wire _w14170_ ;
	wire _w14169_ ;
	wire _w14168_ ;
	wire _w14167_ ;
	wire _w14166_ ;
	wire _w14165_ ;
	wire _w14164_ ;
	wire _w14163_ ;
	wire _w14162_ ;
	wire _w14161_ ;
	wire _w14160_ ;
	wire _w14159_ ;
	wire _w14158_ ;
	wire _w14157_ ;
	wire _w14156_ ;
	wire _w14155_ ;
	wire _w14154_ ;
	wire _w14153_ ;
	wire _w14152_ ;
	wire _w14151_ ;
	wire _w14150_ ;
	wire _w14149_ ;
	wire _w14148_ ;
	wire _w14147_ ;
	wire _w14146_ ;
	wire _w14145_ ;
	wire _w14144_ ;
	wire _w14143_ ;
	wire _w14142_ ;
	wire _w14141_ ;
	wire _w14140_ ;
	wire _w14139_ ;
	wire _w14138_ ;
	wire _w14137_ ;
	wire _w14136_ ;
	wire _w14135_ ;
	wire _w14134_ ;
	wire _w14133_ ;
	wire _w14132_ ;
	wire _w14131_ ;
	wire _w14130_ ;
	wire _w14129_ ;
	wire _w14128_ ;
	wire _w14127_ ;
	wire _w14126_ ;
	wire _w14125_ ;
	wire _w14124_ ;
	wire _w14123_ ;
	wire _w14122_ ;
	wire _w14121_ ;
	wire _w14120_ ;
	wire _w14119_ ;
	wire _w14118_ ;
	wire _w14117_ ;
	wire _w14116_ ;
	wire _w14115_ ;
	wire _w14114_ ;
	wire _w14113_ ;
	wire _w14112_ ;
	wire _w14111_ ;
	wire _w14110_ ;
	wire _w14109_ ;
	wire _w14108_ ;
	wire _w14107_ ;
	wire _w14106_ ;
	wire _w14105_ ;
	wire _w14104_ ;
	wire _w14103_ ;
	wire _w14102_ ;
	wire _w14101_ ;
	wire _w14100_ ;
	wire _w14099_ ;
	wire _w14098_ ;
	wire _w14097_ ;
	wire _w14096_ ;
	wire _w14095_ ;
	wire _w14094_ ;
	wire _w14093_ ;
	wire _w14092_ ;
	wire _w14091_ ;
	wire _w14090_ ;
	wire _w14089_ ;
	wire _w14088_ ;
	wire _w14087_ ;
	wire _w14086_ ;
	wire _w14085_ ;
	wire _w14084_ ;
	wire _w14083_ ;
	wire _w14082_ ;
	wire _w14081_ ;
	wire _w14080_ ;
	wire _w14079_ ;
	wire _w14078_ ;
	wire _w14077_ ;
	wire _w14076_ ;
	wire _w14075_ ;
	wire _w14074_ ;
	wire _w14073_ ;
	wire _w14072_ ;
	wire _w14071_ ;
	wire _w14070_ ;
	wire _w14069_ ;
	wire _w14068_ ;
	wire _w14067_ ;
	wire _w14066_ ;
	wire _w14065_ ;
	wire _w14064_ ;
	wire _w14063_ ;
	wire _w14062_ ;
	wire _w14061_ ;
	wire _w14060_ ;
	wire _w14059_ ;
	wire _w14058_ ;
	wire _w14057_ ;
	wire _w14056_ ;
	wire _w14055_ ;
	wire _w14054_ ;
	wire _w14053_ ;
	wire _w14052_ ;
	wire _w14051_ ;
	wire _w14050_ ;
	wire _w14049_ ;
	wire _w14048_ ;
	wire _w14047_ ;
	wire _w14046_ ;
	wire _w14045_ ;
	wire _w14044_ ;
	wire _w14043_ ;
	wire _w14042_ ;
	wire _w14041_ ;
	wire _w14040_ ;
	wire _w14039_ ;
	wire _w14038_ ;
	wire _w14037_ ;
	wire _w14036_ ;
	wire _w14035_ ;
	wire _w14034_ ;
	wire _w14033_ ;
	wire _w14032_ ;
	wire _w14031_ ;
	wire _w14030_ ;
	wire _w14029_ ;
	wire _w14028_ ;
	wire _w14027_ ;
	wire _w14026_ ;
	wire _w14025_ ;
	wire _w14024_ ;
	wire _w14023_ ;
	wire _w14022_ ;
	wire _w14021_ ;
	wire _w14020_ ;
	wire _w14019_ ;
	wire _w14018_ ;
	wire _w14017_ ;
	wire _w14016_ ;
	wire _w14015_ ;
	wire _w14014_ ;
	wire _w14013_ ;
	wire _w14012_ ;
	wire _w14011_ ;
	wire _w14010_ ;
	wire _w14009_ ;
	wire _w14008_ ;
	wire _w14007_ ;
	wire _w14006_ ;
	wire _w14005_ ;
	wire _w14004_ ;
	wire _w14003_ ;
	wire _w14002_ ;
	wire _w14001_ ;
	wire _w14000_ ;
	wire _w13999_ ;
	wire _w13998_ ;
	wire _w13997_ ;
	wire _w13996_ ;
	wire _w13995_ ;
	wire _w13994_ ;
	wire _w13993_ ;
	wire _w13992_ ;
	wire _w13991_ ;
	wire _w13990_ ;
	wire _w13989_ ;
	wire _w13988_ ;
	wire _w13987_ ;
	wire _w13986_ ;
	wire _w13985_ ;
	wire _w13984_ ;
	wire _w13983_ ;
	wire _w13982_ ;
	wire _w13981_ ;
	wire _w13980_ ;
	wire _w13979_ ;
	wire _w13978_ ;
	wire _w13977_ ;
	wire _w13976_ ;
	wire _w13975_ ;
	wire _w13974_ ;
	wire _w13973_ ;
	wire _w13972_ ;
	wire _w13971_ ;
	wire _w13970_ ;
	wire _w13969_ ;
	wire _w13968_ ;
	wire _w13967_ ;
	wire _w13966_ ;
	wire _w13965_ ;
	wire _w13964_ ;
	wire _w13963_ ;
	wire _w13962_ ;
	wire _w13961_ ;
	wire _w13960_ ;
	wire _w13959_ ;
	wire _w13958_ ;
	wire _w13957_ ;
	wire _w13956_ ;
	wire _w13955_ ;
	wire _w13954_ ;
	wire _w13953_ ;
	wire _w13952_ ;
	wire _w13951_ ;
	wire _w13950_ ;
	wire _w13949_ ;
	wire _w13948_ ;
	wire _w13947_ ;
	wire _w13946_ ;
	wire _w13945_ ;
	wire _w13944_ ;
	wire _w13943_ ;
	wire _w13942_ ;
	wire _w13941_ ;
	wire _w13940_ ;
	wire _w13939_ ;
	wire _w13938_ ;
	wire _w13937_ ;
	wire _w13936_ ;
	wire _w13935_ ;
	wire _w13934_ ;
	wire _w13933_ ;
	wire _w13932_ ;
	wire _w13931_ ;
	wire _w13930_ ;
	wire _w13929_ ;
	wire _w13928_ ;
	wire _w13927_ ;
	wire _w13926_ ;
	wire _w13925_ ;
	wire _w13924_ ;
	wire _w13923_ ;
	wire _w13922_ ;
	wire _w13921_ ;
	wire _w13920_ ;
	wire _w13919_ ;
	wire _w13918_ ;
	wire _w13917_ ;
	wire _w13916_ ;
	wire _w13915_ ;
	wire _w13914_ ;
	wire _w13913_ ;
	wire _w13912_ ;
	wire _w13911_ ;
	wire _w13910_ ;
	wire _w13909_ ;
	wire _w13908_ ;
	wire _w13907_ ;
	wire _w13906_ ;
	wire _w13905_ ;
	wire _w13904_ ;
	wire _w13903_ ;
	wire _w13902_ ;
	wire _w13901_ ;
	wire _w13900_ ;
	wire _w13899_ ;
	wire _w13898_ ;
	wire _w13897_ ;
	wire _w13896_ ;
	wire _w13895_ ;
	wire _w13894_ ;
	wire _w13893_ ;
	wire _w13892_ ;
	wire _w13891_ ;
	wire _w13890_ ;
	wire _w13889_ ;
	wire _w13888_ ;
	wire _w13887_ ;
	wire _w13886_ ;
	wire _w13885_ ;
	wire _w13884_ ;
	wire _w13883_ ;
	wire _w13882_ ;
	wire _w13881_ ;
	wire _w13880_ ;
	wire _w13879_ ;
	wire _w13878_ ;
	wire _w13877_ ;
	wire _w13876_ ;
	wire _w13875_ ;
	wire _w13874_ ;
	wire _w13873_ ;
	wire _w13872_ ;
	wire _w13871_ ;
	wire _w13870_ ;
	wire _w13869_ ;
	wire _w13868_ ;
	wire _w13867_ ;
	wire _w13866_ ;
	wire _w13865_ ;
	wire _w13864_ ;
	wire _w13863_ ;
	wire _w13862_ ;
	wire _w13861_ ;
	wire _w13860_ ;
	wire _w13859_ ;
	wire _w13858_ ;
	wire _w13857_ ;
	wire _w13856_ ;
	wire _w13855_ ;
	wire _w13854_ ;
	wire _w13853_ ;
	wire _w13852_ ;
	wire _w13851_ ;
	wire _w13850_ ;
	wire _w13849_ ;
	wire _w13848_ ;
	wire _w13847_ ;
	wire _w13846_ ;
	wire _w13845_ ;
	wire _w13844_ ;
	wire _w13843_ ;
	wire _w13842_ ;
	wire _w13841_ ;
	wire _w13840_ ;
	wire _w13839_ ;
	wire _w13838_ ;
	wire _w13837_ ;
	wire _w13836_ ;
	wire _w13835_ ;
	wire _w13834_ ;
	wire _w13833_ ;
	wire _w13832_ ;
	wire _w13831_ ;
	wire _w13830_ ;
	wire _w13829_ ;
	wire _w13828_ ;
	wire _w13827_ ;
	wire _w13826_ ;
	wire _w13825_ ;
	wire _w13824_ ;
	wire _w13823_ ;
	wire _w13822_ ;
	wire _w13821_ ;
	wire _w13820_ ;
	wire _w13819_ ;
	wire _w13818_ ;
	wire _w13817_ ;
	wire _w13816_ ;
	wire _w13815_ ;
	wire _w13814_ ;
	wire _w13813_ ;
	wire _w13812_ ;
	wire _w13811_ ;
	wire _w13810_ ;
	wire _w13809_ ;
	wire _w13808_ ;
	wire _w13807_ ;
	wire _w13806_ ;
	wire _w13805_ ;
	wire _w13804_ ;
	wire _w13803_ ;
	wire _w13802_ ;
	wire _w13801_ ;
	wire _w13800_ ;
	wire _w13799_ ;
	wire _w13798_ ;
	wire _w13797_ ;
	wire _w13796_ ;
	wire _w13795_ ;
	wire _w13794_ ;
	wire _w13793_ ;
	wire _w13792_ ;
	wire _w13791_ ;
	wire _w13790_ ;
	wire _w13789_ ;
	wire _w13788_ ;
	wire _w13787_ ;
	wire _w13786_ ;
	wire _w13785_ ;
	wire _w13784_ ;
	wire _w13783_ ;
	wire _w13782_ ;
	wire _w13781_ ;
	wire _w13780_ ;
	wire _w13779_ ;
	wire _w13778_ ;
	wire _w13777_ ;
	wire _w13776_ ;
	wire _w13775_ ;
	wire _w13774_ ;
	wire _w13773_ ;
	wire _w13772_ ;
	wire _w13771_ ;
	wire _w13770_ ;
	wire _w13769_ ;
	wire _w13768_ ;
	wire _w13767_ ;
	wire _w13766_ ;
	wire _w13765_ ;
	wire _w13764_ ;
	wire _w13763_ ;
	wire _w13762_ ;
	wire _w13761_ ;
	wire _w13760_ ;
	wire _w13759_ ;
	wire _w13758_ ;
	wire _w13757_ ;
	wire _w13756_ ;
	wire _w13755_ ;
	wire _w13754_ ;
	wire _w13753_ ;
	wire _w13752_ ;
	wire _w13751_ ;
	wire _w13750_ ;
	wire _w13749_ ;
	wire _w13748_ ;
	wire _w13747_ ;
	wire _w13746_ ;
	wire _w13745_ ;
	wire _w13744_ ;
	wire _w13743_ ;
	wire _w13742_ ;
	wire _w13741_ ;
	wire _w13740_ ;
	wire _w13739_ ;
	wire _w13738_ ;
	wire _w13737_ ;
	wire _w13736_ ;
	wire _w13735_ ;
	wire _w13734_ ;
	wire _w13733_ ;
	wire _w13732_ ;
	wire _w13731_ ;
	wire _w13730_ ;
	wire _w13729_ ;
	wire _w13728_ ;
	wire _w13727_ ;
	wire _w13726_ ;
	wire _w13725_ ;
	wire _w13724_ ;
	wire _w13723_ ;
	wire _w13722_ ;
	wire _w13721_ ;
	wire _w13720_ ;
	wire _w13719_ ;
	wire _w13718_ ;
	wire _w13717_ ;
	wire _w13716_ ;
	wire _w13715_ ;
	wire _w13714_ ;
	wire _w13713_ ;
	wire _w13712_ ;
	wire _w13711_ ;
	wire _w13710_ ;
	wire _w13709_ ;
	wire _w13708_ ;
	wire _w13707_ ;
	wire _w13706_ ;
	wire _w13705_ ;
	wire _w13704_ ;
	wire _w13703_ ;
	wire _w13702_ ;
	wire _w13701_ ;
	wire _w13700_ ;
	wire _w13699_ ;
	wire _w13698_ ;
	wire _w13697_ ;
	wire _w13696_ ;
	wire _w13695_ ;
	wire _w13694_ ;
	wire _w13693_ ;
	wire _w13692_ ;
	wire _w13691_ ;
	wire _w13690_ ;
	wire _w13689_ ;
	wire _w13688_ ;
	wire _w13687_ ;
	wire _w13686_ ;
	wire _w13685_ ;
	wire _w13684_ ;
	wire _w13683_ ;
	wire _w13682_ ;
	wire _w13681_ ;
	wire _w13680_ ;
	wire _w13679_ ;
	wire _w13678_ ;
	wire _w13677_ ;
	wire _w13676_ ;
	wire _w13675_ ;
	wire _w13674_ ;
	wire _w13673_ ;
	wire _w13672_ ;
	wire _w13671_ ;
	wire _w13670_ ;
	wire _w13669_ ;
	wire _w13668_ ;
	wire _w13667_ ;
	wire _w13666_ ;
	wire _w13665_ ;
	wire _w13664_ ;
	wire _w13663_ ;
	wire _w13662_ ;
	wire _w13661_ ;
	wire _w13660_ ;
	wire _w13659_ ;
	wire _w13658_ ;
	wire _w13657_ ;
	wire _w13656_ ;
	wire _w13655_ ;
	wire _w13654_ ;
	wire _w13653_ ;
	wire _w13652_ ;
	wire _w13651_ ;
	wire _w13650_ ;
	wire _w13649_ ;
	wire _w13648_ ;
	wire _w13647_ ;
	wire _w13646_ ;
	wire _w13645_ ;
	wire _w13644_ ;
	wire _w13643_ ;
	wire _w13642_ ;
	wire _w13641_ ;
	wire _w13640_ ;
	wire _w13639_ ;
	wire _w13638_ ;
	wire _w13637_ ;
	wire _w13636_ ;
	wire _w13635_ ;
	wire _w13634_ ;
	wire _w13633_ ;
	wire _w13632_ ;
	wire _w13631_ ;
	wire _w13630_ ;
	wire _w13629_ ;
	wire _w13628_ ;
	wire _w13627_ ;
	wire _w13626_ ;
	wire _w13625_ ;
	wire _w13624_ ;
	wire _w13623_ ;
	wire _w13622_ ;
	wire _w13621_ ;
	wire _w13620_ ;
	wire _w13619_ ;
	wire _w13618_ ;
	wire _w13617_ ;
	wire _w13616_ ;
	wire _w13615_ ;
	wire _w13614_ ;
	wire _w13613_ ;
	wire _w13612_ ;
	wire _w13611_ ;
	wire _w13610_ ;
	wire _w13609_ ;
	wire _w13608_ ;
	wire _w13607_ ;
	wire _w13606_ ;
	wire _w13605_ ;
	wire _w13604_ ;
	wire _w13603_ ;
	wire _w13602_ ;
	wire _w13601_ ;
	wire _w13600_ ;
	wire _w13599_ ;
	wire _w13598_ ;
	wire _w13597_ ;
	wire _w13596_ ;
	wire _w13595_ ;
	wire _w13594_ ;
	wire _w13593_ ;
	wire _w13592_ ;
	wire _w13591_ ;
	wire _w13590_ ;
	wire _w13589_ ;
	wire _w13588_ ;
	wire _w13587_ ;
	wire _w13586_ ;
	wire _w13585_ ;
	wire _w13584_ ;
	wire _w13583_ ;
	wire _w13582_ ;
	wire _w13581_ ;
	wire _w13580_ ;
	wire _w13579_ ;
	wire _w13578_ ;
	wire _w13577_ ;
	wire _w13576_ ;
	wire _w13575_ ;
	wire _w13574_ ;
	wire _w13573_ ;
	wire _w13572_ ;
	wire _w13571_ ;
	wire _w13570_ ;
	wire _w13569_ ;
	wire _w13568_ ;
	wire _w13567_ ;
	wire _w13566_ ;
	wire _w13565_ ;
	wire _w13564_ ;
	wire _w13563_ ;
	wire _w13562_ ;
	wire _w13561_ ;
	wire _w13560_ ;
	wire _w13559_ ;
	wire _w13558_ ;
	wire _w13557_ ;
	wire _w13556_ ;
	wire _w13555_ ;
	wire _w13554_ ;
	wire _w13553_ ;
	wire _w13552_ ;
	wire _w13551_ ;
	wire _w13550_ ;
	wire _w13549_ ;
	wire _w13548_ ;
	wire _w13547_ ;
	wire _w13546_ ;
	wire _w13545_ ;
	wire _w13544_ ;
	wire _w13543_ ;
	wire _w13542_ ;
	wire _w13541_ ;
	wire _w13540_ ;
	wire _w13539_ ;
	wire _w13538_ ;
	wire _w13537_ ;
	wire _w13536_ ;
	wire _w13535_ ;
	wire _w13534_ ;
	wire _w13533_ ;
	wire _w13532_ ;
	wire _w13531_ ;
	wire _w13530_ ;
	wire _w13529_ ;
	wire _w13528_ ;
	wire _w13527_ ;
	wire _w13526_ ;
	wire _w13525_ ;
	wire _w13524_ ;
	wire _w13523_ ;
	wire _w13522_ ;
	wire _w13521_ ;
	wire _w13520_ ;
	wire _w13519_ ;
	wire _w13518_ ;
	wire _w13517_ ;
	wire _w13516_ ;
	wire _w13515_ ;
	wire _w13514_ ;
	wire _w13513_ ;
	wire _w13512_ ;
	wire _w13511_ ;
	wire _w13510_ ;
	wire _w13509_ ;
	wire _w13508_ ;
	wire _w13507_ ;
	wire _w13506_ ;
	wire _w13505_ ;
	wire _w13504_ ;
	wire _w13503_ ;
	wire _w13502_ ;
	wire _w13501_ ;
	wire _w13500_ ;
	wire _w13499_ ;
	wire _w13498_ ;
	wire _w13497_ ;
	wire _w13496_ ;
	wire _w13495_ ;
	wire _w13494_ ;
	wire _w13493_ ;
	wire _w13492_ ;
	wire _w13491_ ;
	wire _w13490_ ;
	wire _w13489_ ;
	wire _w13488_ ;
	wire _w13487_ ;
	wire _w13486_ ;
	wire _w13485_ ;
	wire _w13484_ ;
	wire _w13483_ ;
	wire _w13482_ ;
	wire _w13481_ ;
	wire _w13480_ ;
	wire _w13479_ ;
	wire _w13478_ ;
	wire _w13477_ ;
	wire _w13476_ ;
	wire _w13475_ ;
	wire _w13474_ ;
	wire _w13473_ ;
	wire _w13472_ ;
	wire _w13471_ ;
	wire _w13470_ ;
	wire _w13469_ ;
	wire _w13468_ ;
	wire _w13467_ ;
	wire _w13466_ ;
	wire _w13465_ ;
	wire _w13464_ ;
	wire _w13463_ ;
	wire _w13462_ ;
	wire _w13461_ ;
	wire _w13460_ ;
	wire _w13459_ ;
	wire _w13458_ ;
	wire _w13457_ ;
	wire _w13456_ ;
	wire _w13455_ ;
	wire _w13454_ ;
	wire _w13453_ ;
	wire _w13452_ ;
	wire _w13451_ ;
	wire _w13450_ ;
	wire _w13449_ ;
	wire _w13448_ ;
	wire _w13447_ ;
	wire _w13446_ ;
	wire _w13445_ ;
	wire _w13444_ ;
	wire _w13443_ ;
	wire _w13442_ ;
	wire _w13441_ ;
	wire _w13440_ ;
	wire _w13439_ ;
	wire _w13438_ ;
	wire _w13437_ ;
	wire _w13436_ ;
	wire _w13435_ ;
	wire _w13434_ ;
	wire _w13433_ ;
	wire _w13432_ ;
	wire _w13431_ ;
	wire _w13430_ ;
	wire _w13429_ ;
	wire _w13428_ ;
	wire _w13427_ ;
	wire _w13426_ ;
	wire _w13425_ ;
	wire _w13424_ ;
	wire _w13423_ ;
	wire _w13422_ ;
	wire _w13421_ ;
	wire _w13420_ ;
	wire _w13419_ ;
	wire _w13418_ ;
	wire _w13417_ ;
	wire _w13416_ ;
	wire _w13415_ ;
	wire _w13414_ ;
	wire _w13413_ ;
	wire _w13412_ ;
	wire _w13411_ ;
	wire _w13410_ ;
	wire _w13409_ ;
	wire _w13408_ ;
	wire _w13407_ ;
	wire _w13406_ ;
	wire _w13405_ ;
	wire _w13404_ ;
	wire _w13403_ ;
	wire _w13402_ ;
	wire _w13401_ ;
	wire _w13400_ ;
	wire _w13399_ ;
	wire _w13398_ ;
	wire _w13397_ ;
	wire _w13396_ ;
	wire _w13395_ ;
	wire _w13394_ ;
	wire _w13393_ ;
	wire _w13392_ ;
	wire _w13391_ ;
	wire _w13390_ ;
	wire _w13389_ ;
	wire _w13388_ ;
	wire _w13387_ ;
	wire _w13386_ ;
	wire _w13385_ ;
	wire _w13384_ ;
	wire _w13383_ ;
	wire _w13382_ ;
	wire _w13381_ ;
	wire _w13380_ ;
	wire _w13379_ ;
	wire _w13378_ ;
	wire _w13377_ ;
	wire _w13376_ ;
	wire _w13375_ ;
	wire _w13374_ ;
	wire _w13373_ ;
	wire _w13372_ ;
	wire _w13371_ ;
	wire _w13370_ ;
	wire _w13369_ ;
	wire _w13368_ ;
	wire _w13367_ ;
	wire _w13366_ ;
	wire _w13365_ ;
	wire _w13364_ ;
	wire _w13363_ ;
	wire _w13362_ ;
	wire _w13361_ ;
	wire _w13360_ ;
	wire _w13359_ ;
	wire _w13358_ ;
	wire _w13357_ ;
	wire _w13356_ ;
	wire _w13355_ ;
	wire _w13354_ ;
	wire _w13353_ ;
	wire _w13352_ ;
	wire _w13351_ ;
	wire _w13350_ ;
	wire _w13349_ ;
	wire _w13348_ ;
	wire _w13347_ ;
	wire _w13346_ ;
	wire _w13345_ ;
	wire _w13344_ ;
	wire _w13343_ ;
	wire _w13342_ ;
	wire _w13341_ ;
	wire _w13340_ ;
	wire _w13339_ ;
	wire _w13338_ ;
	wire _w13337_ ;
	wire _w13336_ ;
	wire _w13335_ ;
	wire _w13334_ ;
	wire _w13333_ ;
	wire _w13332_ ;
	wire _w13331_ ;
	wire _w13330_ ;
	wire _w13329_ ;
	wire _w13328_ ;
	wire _w13327_ ;
	wire _w13326_ ;
	wire _w13325_ ;
	wire _w13324_ ;
	wire _w13323_ ;
	wire _w13322_ ;
	wire _w13321_ ;
	wire _w13320_ ;
	wire _w13319_ ;
	wire _w13318_ ;
	wire _w13317_ ;
	wire _w13316_ ;
	wire _w13315_ ;
	wire _w13314_ ;
	wire _w13313_ ;
	wire _w13312_ ;
	wire _w13311_ ;
	wire _w13310_ ;
	wire _w13309_ ;
	wire _w13308_ ;
	wire _w13307_ ;
	wire _w13306_ ;
	wire _w13305_ ;
	wire _w13304_ ;
	wire _w13303_ ;
	wire _w13302_ ;
	wire _w13301_ ;
	wire _w13300_ ;
	wire _w13299_ ;
	wire _w13298_ ;
	wire _w13297_ ;
	wire _w13296_ ;
	wire _w13295_ ;
	wire _w13294_ ;
	wire _w13293_ ;
	wire _w13292_ ;
	wire _w13291_ ;
	wire _w13290_ ;
	wire _w13289_ ;
	wire _w13288_ ;
	wire _w13287_ ;
	wire _w13286_ ;
	wire _w13285_ ;
	wire _w13284_ ;
	wire _w13283_ ;
	wire _w13282_ ;
	wire _w13281_ ;
	wire _w13280_ ;
	wire _w13279_ ;
	wire _w13278_ ;
	wire _w13277_ ;
	wire _w13276_ ;
	wire _w13275_ ;
	wire _w13274_ ;
	wire _w13273_ ;
	wire _w13272_ ;
	wire _w13271_ ;
	wire _w13270_ ;
	wire _w13269_ ;
	wire _w13268_ ;
	wire _w13267_ ;
	wire _w13266_ ;
	wire _w13265_ ;
	wire _w13264_ ;
	wire _w13263_ ;
	wire _w13262_ ;
	wire _w13261_ ;
	wire _w13260_ ;
	wire _w13259_ ;
	wire _w13258_ ;
	wire _w13257_ ;
	wire _w13256_ ;
	wire _w13255_ ;
	wire _w13254_ ;
	wire _w13253_ ;
	wire _w13252_ ;
	wire _w13251_ ;
	wire _w13250_ ;
	wire _w13249_ ;
	wire _w13248_ ;
	wire _w13247_ ;
	wire _w13246_ ;
	wire _w13245_ ;
	wire _w13244_ ;
	wire _w13243_ ;
	wire _w13242_ ;
	wire _w13241_ ;
	wire _w13240_ ;
	wire _w13239_ ;
	wire _w13238_ ;
	wire _w13237_ ;
	wire _w13236_ ;
	wire _w13235_ ;
	wire _w13234_ ;
	wire _w13233_ ;
	wire _w13232_ ;
	wire _w13231_ ;
	wire _w13230_ ;
	wire _w13229_ ;
	wire _w13228_ ;
	wire _w13227_ ;
	wire _w13226_ ;
	wire _w13225_ ;
	wire _w13224_ ;
	wire _w13223_ ;
	wire _w13222_ ;
	wire _w13221_ ;
	wire _w13220_ ;
	wire _w13219_ ;
	wire _w13218_ ;
	wire _w13217_ ;
	wire _w13216_ ;
	wire _w13215_ ;
	wire _w13214_ ;
	wire _w13213_ ;
	wire _w13212_ ;
	wire _w13211_ ;
	wire _w13210_ ;
	wire _w13209_ ;
	wire _w13208_ ;
	wire _w13207_ ;
	wire _w13206_ ;
	wire _w13205_ ;
	wire _w13204_ ;
	wire _w13203_ ;
	wire _w13202_ ;
	wire _w13201_ ;
	wire _w13200_ ;
	wire _w13199_ ;
	wire _w13198_ ;
	wire _w13197_ ;
	wire _w13196_ ;
	wire _w13195_ ;
	wire _w13194_ ;
	wire _w13193_ ;
	wire _w13192_ ;
	wire _w13191_ ;
	wire _w13190_ ;
	wire _w13189_ ;
	wire _w13188_ ;
	wire _w13187_ ;
	wire _w13186_ ;
	wire _w13185_ ;
	wire _w13184_ ;
	wire _w13183_ ;
	wire _w13182_ ;
	wire _w13181_ ;
	wire _w13180_ ;
	wire _w13179_ ;
	wire _w13178_ ;
	wire _w13177_ ;
	wire _w13176_ ;
	wire _w13175_ ;
	wire _w13174_ ;
	wire _w13173_ ;
	wire _w13172_ ;
	wire _w13171_ ;
	wire _w13170_ ;
	wire _w13169_ ;
	wire _w13168_ ;
	wire _w13167_ ;
	wire _w13166_ ;
	wire _w13165_ ;
	wire _w13164_ ;
	wire _w13163_ ;
	wire _w13162_ ;
	wire _w13161_ ;
	wire _w13160_ ;
	wire _w13159_ ;
	wire _w13158_ ;
	wire _w13157_ ;
	wire _w13156_ ;
	wire _w13155_ ;
	wire _w13154_ ;
	wire _w13153_ ;
	wire _w13152_ ;
	wire _w13151_ ;
	wire _w13150_ ;
	wire _w13149_ ;
	wire _w13148_ ;
	wire _w13147_ ;
	wire _w13146_ ;
	wire _w13145_ ;
	wire _w13144_ ;
	wire _w13143_ ;
	wire _w13142_ ;
	wire _w13141_ ;
	wire _w13140_ ;
	wire _w13139_ ;
	wire _w13138_ ;
	wire _w13137_ ;
	wire _w13136_ ;
	wire _w13135_ ;
	wire _w13134_ ;
	wire _w13133_ ;
	wire _w13132_ ;
	wire _w13131_ ;
	wire _w13130_ ;
	wire _w13129_ ;
	wire _w13128_ ;
	wire _w13127_ ;
	wire _w13126_ ;
	wire _w13125_ ;
	wire _w13124_ ;
	wire _w13123_ ;
	wire _w13122_ ;
	wire _w13121_ ;
	wire _w13120_ ;
	wire _w13119_ ;
	wire _w13118_ ;
	wire _w13117_ ;
	wire _w13116_ ;
	wire _w13115_ ;
	wire _w13114_ ;
	wire _w13113_ ;
	wire _w13112_ ;
	wire _w13111_ ;
	wire _w13110_ ;
	wire _w13109_ ;
	wire _w13108_ ;
	wire _w13107_ ;
	wire _w13106_ ;
	wire _w13105_ ;
	wire _w13104_ ;
	wire _w13103_ ;
	wire _w13102_ ;
	wire _w13101_ ;
	wire _w13100_ ;
	wire _w13099_ ;
	wire _w13098_ ;
	wire _w13097_ ;
	wire _w13096_ ;
	wire _w13095_ ;
	wire _w13094_ ;
	wire _w13093_ ;
	wire _w13092_ ;
	wire _w13091_ ;
	wire _w13090_ ;
	wire _w13089_ ;
	wire _w13088_ ;
	wire _w13087_ ;
	wire _w13086_ ;
	wire _w13085_ ;
	wire _w13084_ ;
	wire _w13083_ ;
	wire _w13082_ ;
	wire _w13081_ ;
	wire _w13080_ ;
	wire _w13079_ ;
	wire _w13078_ ;
	wire _w13077_ ;
	wire _w13076_ ;
	wire _w13075_ ;
	wire _w13074_ ;
	wire _w13073_ ;
	wire _w13072_ ;
	wire _w13071_ ;
	wire _w13070_ ;
	wire _w13069_ ;
	wire _w13068_ ;
	wire _w13067_ ;
	wire _w13066_ ;
	wire _w13065_ ;
	wire _w13064_ ;
	wire _w13063_ ;
	wire _w13062_ ;
	wire _w13061_ ;
	wire _w13060_ ;
	wire _w13059_ ;
	wire _w13058_ ;
	wire _w13057_ ;
	wire _w13056_ ;
	wire _w13055_ ;
	wire _w13054_ ;
	wire _w13053_ ;
	wire _w13052_ ;
	wire _w13051_ ;
	wire _w13050_ ;
	wire _w13049_ ;
	wire _w13048_ ;
	wire _w13047_ ;
	wire _w13046_ ;
	wire _w13045_ ;
	wire _w13044_ ;
	wire _w13043_ ;
	wire _w13042_ ;
	wire _w13041_ ;
	wire _w13040_ ;
	wire _w13039_ ;
	wire _w13038_ ;
	wire _w13037_ ;
	wire _w13036_ ;
	wire _w13035_ ;
	wire _w13034_ ;
	wire _w13033_ ;
	wire _w13032_ ;
	wire _w13031_ ;
	wire _w13030_ ;
	wire _w13029_ ;
	wire _w13028_ ;
	wire _w13027_ ;
	wire _w13026_ ;
	wire _w13025_ ;
	wire _w13024_ ;
	wire _w13023_ ;
	wire _w13022_ ;
	wire _w13021_ ;
	wire _w13020_ ;
	wire _w13019_ ;
	wire _w13018_ ;
	wire _w13017_ ;
	wire _w13016_ ;
	wire _w13015_ ;
	wire _w13014_ ;
	wire _w13013_ ;
	wire _w13012_ ;
	wire _w13011_ ;
	wire _w13010_ ;
	wire _w13009_ ;
	wire _w13008_ ;
	wire _w13007_ ;
	wire _w13006_ ;
	wire _w13005_ ;
	wire _w13004_ ;
	wire _w13003_ ;
	wire _w13002_ ;
	wire _w13001_ ;
	wire _w13000_ ;
	wire _w12999_ ;
	wire _w12998_ ;
	wire _w12997_ ;
	wire _w12996_ ;
	wire _w12995_ ;
	wire _w12994_ ;
	wire _w12993_ ;
	wire _w12992_ ;
	wire _w12991_ ;
	wire _w12990_ ;
	wire _w12989_ ;
	wire _w12988_ ;
	wire _w12987_ ;
	wire _w12986_ ;
	wire _w12985_ ;
	wire _w12984_ ;
	wire _w12983_ ;
	wire _w12982_ ;
	wire _w12981_ ;
	wire _w12980_ ;
	wire _w12979_ ;
	wire _w12978_ ;
	wire _w12977_ ;
	wire _w12976_ ;
	wire _w12975_ ;
	wire _w12974_ ;
	wire _w12973_ ;
	wire _w12972_ ;
	wire _w12971_ ;
	wire _w12970_ ;
	wire _w12969_ ;
	wire _w12968_ ;
	wire _w12967_ ;
	wire _w12966_ ;
	wire _w12965_ ;
	wire _w12964_ ;
	wire _w12963_ ;
	wire _w12962_ ;
	wire _w12961_ ;
	wire _w12960_ ;
	wire _w12959_ ;
	wire _w12958_ ;
	wire _w12957_ ;
	wire _w12956_ ;
	wire _w12955_ ;
	wire _w12954_ ;
	wire _w12953_ ;
	wire _w12952_ ;
	wire _w12951_ ;
	wire _w12950_ ;
	wire _w12949_ ;
	wire _w12948_ ;
	wire _w12947_ ;
	wire _w12946_ ;
	wire _w12945_ ;
	wire _w12944_ ;
	wire _w12943_ ;
	wire _w12942_ ;
	wire _w12941_ ;
	wire _w12940_ ;
	wire _w12939_ ;
	wire _w12938_ ;
	wire _w12937_ ;
	wire _w12936_ ;
	wire _w12935_ ;
	wire _w12934_ ;
	wire _w12933_ ;
	wire _w12932_ ;
	wire _w12931_ ;
	wire _w12930_ ;
	wire _w12929_ ;
	wire _w12928_ ;
	wire _w12927_ ;
	wire _w12926_ ;
	wire _w12925_ ;
	wire _w12924_ ;
	wire _w12923_ ;
	wire _w12922_ ;
	wire _w12921_ ;
	wire _w12920_ ;
	wire _w12919_ ;
	wire _w12918_ ;
	wire _w12917_ ;
	wire _w12916_ ;
	wire _w12915_ ;
	wire _w12914_ ;
	wire _w12913_ ;
	wire _w12912_ ;
	wire _w12911_ ;
	wire _w12910_ ;
	wire _w12909_ ;
	wire _w12908_ ;
	wire _w12907_ ;
	wire _w12906_ ;
	wire _w12905_ ;
	wire _w12904_ ;
	wire _w12903_ ;
	wire _w12902_ ;
	wire _w12901_ ;
	wire _w12900_ ;
	wire _w12899_ ;
	wire _w12898_ ;
	wire _w12897_ ;
	wire _w12896_ ;
	wire _w12895_ ;
	wire _w12894_ ;
	wire _w12893_ ;
	wire _w12892_ ;
	wire _w12891_ ;
	wire _w12890_ ;
	wire _w12889_ ;
	wire _w12888_ ;
	wire _w12887_ ;
	wire _w12886_ ;
	wire _w12885_ ;
	wire _w12884_ ;
	wire _w12883_ ;
	wire _w12882_ ;
	wire _w12881_ ;
	wire _w12880_ ;
	wire _w12879_ ;
	wire _w12878_ ;
	wire _w12877_ ;
	wire _w12876_ ;
	wire _w12875_ ;
	wire _w12874_ ;
	wire _w12873_ ;
	wire _w12872_ ;
	wire _w12871_ ;
	wire _w12870_ ;
	wire _w11621_ ;
	wire _w11620_ ;
	wire _w11619_ ;
	wire _w11618_ ;
	wire _w11617_ ;
	wire _w11616_ ;
	wire _w11615_ ;
	wire _w11614_ ;
	wire _w11613_ ;
	wire _w11612_ ;
	wire _w11611_ ;
	wire _w11610_ ;
	wire _w11609_ ;
	wire _w11608_ ;
	wire _w11607_ ;
	wire _w11606_ ;
	wire _w11605_ ;
	wire _w11604_ ;
	wire _w11603_ ;
	wire _w11602_ ;
	wire _w11601_ ;
	wire _w11600_ ;
	wire _w11599_ ;
	wire _w11598_ ;
	wire _w11597_ ;
	wire _w11596_ ;
	wire _w11595_ ;
	wire _w11594_ ;
	wire _w11593_ ;
	wire _w11592_ ;
	wire _w11591_ ;
	wire _w11590_ ;
	wire _w11589_ ;
	wire _w11588_ ;
	wire _w11587_ ;
	wire _w11586_ ;
	wire _w11585_ ;
	wire _w11584_ ;
	wire _w11583_ ;
	wire _w11582_ ;
	wire _w11581_ ;
	wire _w11580_ ;
	wire _w11579_ ;
	wire _w11578_ ;
	wire _w11577_ ;
	wire _w11576_ ;
	wire _w11575_ ;
	wire _w11574_ ;
	wire _w11573_ ;
	wire _w11572_ ;
	wire _w11571_ ;
	wire _w11570_ ;
	wire _w11569_ ;
	wire _w11568_ ;
	wire _w11567_ ;
	wire _w11566_ ;
	wire _w11565_ ;
	wire _w11564_ ;
	wire _w11563_ ;
	wire _w11562_ ;
	wire _w11561_ ;
	wire _w11560_ ;
	wire _w11559_ ;
	wire _w11558_ ;
	wire _w11557_ ;
	wire _w11556_ ;
	wire _w11555_ ;
	wire _w11554_ ;
	wire _w11553_ ;
	wire _w11552_ ;
	wire _w11551_ ;
	wire _w11549_ ;
	wire _w11548_ ;
	wire _w11547_ ;
	wire _w11546_ ;
	wire _w11545_ ;
	wire _w11544_ ;
	wire _w11543_ ;
	wire _w11542_ ;
	wire _w11541_ ;
	wire _w11540_ ;
	wire _w11539_ ;
	wire _w11538_ ;
	wire _w11537_ ;
	wire _w11536_ ;
	wire _w11535_ ;
	wire _w11534_ ;
	wire _w11533_ ;
	wire _w11532_ ;
	wire _w11531_ ;
	wire _w11530_ ;
	wire _w11529_ ;
	wire _w11528_ ;
	wire _w11527_ ;
	wire _w11526_ ;
	wire _w11525_ ;
	wire _w11524_ ;
	wire _w11523_ ;
	wire _w11522_ ;
	wire _w11521_ ;
	wire _w11520_ ;
	wire _w11519_ ;
	wire _w11518_ ;
	wire _w11517_ ;
	wire _w11516_ ;
	wire _w11515_ ;
	wire _w11514_ ;
	wire _w11513_ ;
	wire _w11512_ ;
	wire _w11511_ ;
	wire _w11510_ ;
	wire _w11509_ ;
	wire _w11508_ ;
	wire _w11507_ ;
	wire _w11506_ ;
	wire _w11505_ ;
	wire _w11504_ ;
	wire _w11503_ ;
	wire _w11502_ ;
	wire _w11501_ ;
	wire _w11500_ ;
	wire _w11499_ ;
	wire _w11498_ ;
	wire _w11497_ ;
	wire _w11496_ ;
	wire _w11495_ ;
	wire _w11494_ ;
	wire _w11493_ ;
	wire _w11492_ ;
	wire _w11491_ ;
	wire _w11490_ ;
	wire _w11489_ ;
	wire _w11488_ ;
	wire _w11487_ ;
	wire _w11486_ ;
	wire _w11485_ ;
	wire _w11484_ ;
	wire _w11483_ ;
	wire _w11482_ ;
	wire _w11481_ ;
	wire _w11480_ ;
	wire _w11479_ ;
	wire _w11478_ ;
	wire _w11477_ ;
	wire _w11476_ ;
	wire _w11475_ ;
	wire _w11474_ ;
	wire _w11473_ ;
	wire _w11472_ ;
	wire _w11471_ ;
	wire _w11470_ ;
	wire _w11469_ ;
	wire _w11468_ ;
	wire _w11467_ ;
	wire _w11466_ ;
	wire _w11465_ ;
	wire _w11464_ ;
	wire _w11463_ ;
	wire _w11462_ ;
	wire _w11461_ ;
	wire _w11460_ ;
	wire _w11459_ ;
	wire _w11458_ ;
	wire _w11457_ ;
	wire _w11456_ ;
	wire _w11455_ ;
	wire _w11454_ ;
	wire _w11453_ ;
	wire _w11452_ ;
	wire _w11451_ ;
	wire _w11450_ ;
	wire _w11449_ ;
	wire _w11448_ ;
	wire _w11447_ ;
	wire _w11446_ ;
	wire _w11445_ ;
	wire _w11444_ ;
	wire _w11443_ ;
	wire _w11442_ ;
	wire _w11441_ ;
	wire _w11440_ ;
	wire _w11439_ ;
	wire _w11438_ ;
	wire _w11437_ ;
	wire _w11436_ ;
	wire _w11435_ ;
	wire _w11434_ ;
	wire _w11433_ ;
	wire _w11432_ ;
	wire _w11431_ ;
	wire _w11430_ ;
	wire _w11429_ ;
	wire _w11428_ ;
	wire _w11427_ ;
	wire _w11426_ ;
	wire _w11425_ ;
	wire _w11424_ ;
	wire _w11423_ ;
	wire _w11422_ ;
	wire _w11421_ ;
	wire _w11420_ ;
	wire _w11419_ ;
	wire _w11418_ ;
	wire _w11417_ ;
	wire _w11416_ ;
	wire _w11415_ ;
	wire _w11414_ ;
	wire _w11413_ ;
	wire _w11412_ ;
	wire _w11411_ ;
	wire _w11410_ ;
	wire _w11409_ ;
	wire _w11408_ ;
	wire _w11407_ ;
	wire _w11406_ ;
	wire _w11405_ ;
	wire _w11404_ ;
	wire _w11403_ ;
	wire _w11402_ ;
	wire _w11401_ ;
	wire _w11400_ ;
	wire _w11399_ ;
	wire _w11398_ ;
	wire _w11397_ ;
	wire _w11396_ ;
	wire _w11395_ ;
	wire _w11394_ ;
	wire _w11393_ ;
	wire _w11392_ ;
	wire _w11391_ ;
	wire _w11390_ ;
	wire _w11389_ ;
	wire _w11388_ ;
	wire _w11387_ ;
	wire _w11386_ ;
	wire _w11385_ ;
	wire _w11384_ ;
	wire _w11383_ ;
	wire _w11382_ ;
	wire _w11381_ ;
	wire _w11380_ ;
	wire _w11379_ ;
	wire _w11378_ ;
	wire _w11377_ ;
	wire _w11376_ ;
	wire _w11375_ ;
	wire _w11374_ ;
	wire _w11373_ ;
	wire _w11372_ ;
	wire _w11371_ ;
	wire _w11370_ ;
	wire _w11369_ ;
	wire _w11368_ ;
	wire _w11367_ ;
	wire _w11366_ ;
	wire _w11365_ ;
	wire _w11364_ ;
	wire _w11363_ ;
	wire _w11362_ ;
	wire _w11361_ ;
	wire _w11360_ ;
	wire _w11359_ ;
	wire _w11358_ ;
	wire _w11357_ ;
	wire _w11356_ ;
	wire _w11355_ ;
	wire _w11354_ ;
	wire _w11353_ ;
	wire _w11352_ ;
	wire _w11351_ ;
	wire _w11350_ ;
	wire _w11349_ ;
	wire _w11348_ ;
	wire _w11347_ ;
	wire _w11346_ ;
	wire _w11345_ ;
	wire _w11344_ ;
	wire _w11343_ ;
	wire _w11342_ ;
	wire _w11341_ ;
	wire _w11340_ ;
	wire _w11339_ ;
	wire _w11338_ ;
	wire _w11337_ ;
	wire _w11336_ ;
	wire _w11335_ ;
	wire _w11334_ ;
	wire _w11333_ ;
	wire _w11332_ ;
	wire _w11331_ ;
	wire _w11330_ ;
	wire _w11329_ ;
	wire _w11328_ ;
	wire _w11327_ ;
	wire _w11326_ ;
	wire _w11325_ ;
	wire _w11324_ ;
	wire _w11323_ ;
	wire _w11322_ ;
	wire _w11321_ ;
	wire _w11320_ ;
	wire _w11319_ ;
	wire _w11318_ ;
	wire _w11317_ ;
	wire _w11316_ ;
	wire _w11315_ ;
	wire _w11314_ ;
	wire _w11313_ ;
	wire _w11312_ ;
	wire _w11311_ ;
	wire _w11310_ ;
	wire _w11309_ ;
	wire _w11308_ ;
	wire _w11307_ ;
	wire _w11306_ ;
	wire _w11305_ ;
	wire _w11304_ ;
	wire _w11303_ ;
	wire _w11302_ ;
	wire _w11301_ ;
	wire _w11300_ ;
	wire _w11299_ ;
	wire _w11298_ ;
	wire _w11297_ ;
	wire _w11296_ ;
	wire _w11295_ ;
	wire _w11294_ ;
	wire _w11293_ ;
	wire _w11292_ ;
	wire _w11291_ ;
	wire _w11290_ ;
	wire _w11289_ ;
	wire _w11288_ ;
	wire _w11287_ ;
	wire _w11286_ ;
	wire _w11285_ ;
	wire _w11284_ ;
	wire _w11283_ ;
	wire _w11282_ ;
	wire _w11281_ ;
	wire _w11280_ ;
	wire _w11279_ ;
	wire _w11278_ ;
	wire _w11277_ ;
	wire _w11276_ ;
	wire _w11275_ ;
	wire _w11274_ ;
	wire _w11273_ ;
	wire _w11272_ ;
	wire _w11271_ ;
	wire _w11270_ ;
	wire _w11269_ ;
	wire _w11268_ ;
	wire _w11267_ ;
	wire _w11266_ ;
	wire _w11265_ ;
	wire _w11264_ ;
	wire _w11263_ ;
	wire _w11262_ ;
	wire _w11261_ ;
	wire _w11260_ ;
	wire _w11259_ ;
	wire _w11258_ ;
	wire _w11257_ ;
	wire _w11256_ ;
	wire _w11255_ ;
	wire _w11254_ ;
	wire _w11253_ ;
	wire _w11252_ ;
	wire _w11251_ ;
	wire _w11250_ ;
	wire _w11249_ ;
	wire _w11248_ ;
	wire _w11247_ ;
	wire _w11246_ ;
	wire _w11245_ ;
	wire _w11244_ ;
	wire _w11243_ ;
	wire _w11242_ ;
	wire _w11241_ ;
	wire _w11240_ ;
	wire _w11239_ ;
	wire _w11238_ ;
	wire _w11237_ ;
	wire _w11236_ ;
	wire _w11235_ ;
	wire _w11234_ ;
	wire _w11233_ ;
	wire _w11232_ ;
	wire _w11231_ ;
	wire _w11230_ ;
	wire _w11229_ ;
	wire _w11228_ ;
	wire _w11227_ ;
	wire _w11226_ ;
	wire _w11225_ ;
	wire _w11224_ ;
	wire _w11223_ ;
	wire _w11222_ ;
	wire _w11221_ ;
	wire _w11220_ ;
	wire _w11219_ ;
	wire _w11218_ ;
	wire _w11217_ ;
	wire _w11216_ ;
	wire _w11215_ ;
	wire _w11214_ ;
	wire _w11213_ ;
	wire _w11212_ ;
	wire _w11211_ ;
	wire _w11210_ ;
	wire _w11209_ ;
	wire _w11208_ ;
	wire _w11207_ ;
	wire _w11206_ ;
	wire _w11205_ ;
	wire _w11204_ ;
	wire _w11203_ ;
	wire _w11202_ ;
	wire _w11201_ ;
	wire _w11200_ ;
	wire _w11199_ ;
	wire _w11198_ ;
	wire _w11197_ ;
	wire _w11196_ ;
	wire _w11195_ ;
	wire _w11194_ ;
	wire _w11193_ ;
	wire _w11192_ ;
	wire _w11191_ ;
	wire _w11190_ ;
	wire _w11189_ ;
	wire _w11188_ ;
	wire _w11187_ ;
	wire _w11186_ ;
	wire _w11185_ ;
	wire _w11184_ ;
	wire _w11183_ ;
	wire _w11182_ ;
	wire _w11181_ ;
	wire _w11180_ ;
	wire _w11179_ ;
	wire _w11178_ ;
	wire _w11177_ ;
	wire _w11176_ ;
	wire _w11175_ ;
	wire _w11174_ ;
	wire _w11173_ ;
	wire _w11172_ ;
	wire _w11171_ ;
	wire _w11170_ ;
	wire _w11169_ ;
	wire _w11168_ ;
	wire _w11167_ ;
	wire _w11166_ ;
	wire _w11165_ ;
	wire _w11164_ ;
	wire _w11163_ ;
	wire _w11162_ ;
	wire _w11161_ ;
	wire _w11160_ ;
	wire _w11159_ ;
	wire _w11158_ ;
	wire _w11157_ ;
	wire _w11156_ ;
	wire _w11155_ ;
	wire _w11154_ ;
	wire _w11153_ ;
	wire _w11152_ ;
	wire _w11151_ ;
	wire _w11150_ ;
	wire _w11149_ ;
	wire _w11148_ ;
	wire _w11147_ ;
	wire _w11146_ ;
	wire _w11145_ ;
	wire _w11144_ ;
	wire _w11143_ ;
	wire _w11142_ ;
	wire _w11141_ ;
	wire _w11140_ ;
	wire _w11139_ ;
	wire _w11138_ ;
	wire _w11137_ ;
	wire _w11136_ ;
	wire _w11135_ ;
	wire _w11134_ ;
	wire _w11133_ ;
	wire _w11132_ ;
	wire _w11131_ ;
	wire _w11130_ ;
	wire _w11129_ ;
	wire _w11128_ ;
	wire _w11127_ ;
	wire _w11126_ ;
	wire _w11125_ ;
	wire _w11124_ ;
	wire _w11123_ ;
	wire _w11122_ ;
	wire _w11121_ ;
	wire _w11120_ ;
	wire _w11119_ ;
	wire _w11118_ ;
	wire _w11117_ ;
	wire _w11116_ ;
	wire _w11115_ ;
	wire _w11114_ ;
	wire _w11113_ ;
	wire _w11112_ ;
	wire _w11111_ ;
	wire _w11110_ ;
	wire _w11109_ ;
	wire _w11108_ ;
	wire _w11107_ ;
	wire _w11106_ ;
	wire _w11105_ ;
	wire _w11104_ ;
	wire _w11103_ ;
	wire _w11102_ ;
	wire _w11101_ ;
	wire _w11100_ ;
	wire _w11099_ ;
	wire _w11098_ ;
	wire _w11097_ ;
	wire _w11096_ ;
	wire _w11095_ ;
	wire _w11094_ ;
	wire _w11093_ ;
	wire _w11092_ ;
	wire _w11091_ ;
	wire _w11090_ ;
	wire _w11089_ ;
	wire _w11088_ ;
	wire _w11087_ ;
	wire _w11086_ ;
	wire _w11085_ ;
	wire _w11084_ ;
	wire _w11083_ ;
	wire _w11082_ ;
	wire _w11081_ ;
	wire _w11080_ ;
	wire _w11079_ ;
	wire _w11078_ ;
	wire _w11077_ ;
	wire _w11076_ ;
	wire _w11075_ ;
	wire _w11074_ ;
	wire _w11073_ ;
	wire _w11072_ ;
	wire _w11071_ ;
	wire _w11070_ ;
	wire _w11069_ ;
	wire _w11068_ ;
	wire _w11067_ ;
	wire _w11066_ ;
	wire _w11065_ ;
	wire _w11064_ ;
	wire _w11063_ ;
	wire _w11062_ ;
	wire _w11061_ ;
	wire _w11060_ ;
	wire _w11059_ ;
	wire _w11058_ ;
	wire _w11057_ ;
	wire _w11056_ ;
	wire _w11055_ ;
	wire _w11054_ ;
	wire _w10769_ ;
	wire _w10768_ ;
	wire _w10767_ ;
	wire _w10766_ ;
	wire _w10765_ ;
	wire _w10764_ ;
	wire _w10763_ ;
	wire _w10762_ ;
	wire _w10761_ ;
	wire _w10760_ ;
	wire _w10759_ ;
	wire _w10758_ ;
	wire _w10757_ ;
	wire _w10756_ ;
	wire _w10755_ ;
	wire _w10754_ ;
	wire _w10753_ ;
	wire _w10752_ ;
	wire _w10751_ ;
	wire _w10750_ ;
	wire _w10749_ ;
	wire _w10748_ ;
	wire _w10747_ ;
	wire _w10746_ ;
	wire _w10745_ ;
	wire _w10744_ ;
	wire _w10743_ ;
	wire _w10742_ ;
	wire _w10741_ ;
	wire _w10739_ ;
	wire _w11550_ ;
	wire _w12245_ ;
	wire _w10738_ ;
	wire _w10737_ ;
	wire _w10736_ ;
	wire _w10735_ ;
	wire _w10734_ ;
	wire _w10733_ ;
	wire _w21213_ ;
	wire _w460_ ;
	wire _w10732_ ;
	wire _w10731_ ;
	wire _w10730_ ;
	wire _w10729_ ;
	wire _w10728_ ;
	wire _w10727_ ;
	wire _w10726_ ;
	wire _w10725_ ;
	wire _w10724_ ;
	wire _w10723_ ;
	wire _w10722_ ;
	wire _w10721_ ;
	wire _w10720_ ;
	wire _w10719_ ;
	wire _w10718_ ;
	wire _w10717_ ;
	wire _w10716_ ;
	wire _w10715_ ;
	wire _w10714_ ;
	wire _w10713_ ;
	wire _w10712_ ;
	wire _w10711_ ;
	wire _w10710_ ;
	wire _w10709_ ;
	wire _w10708_ ;
	wire _w10707_ ;
	wire _w10706_ ;
	wire _w10705_ ;
	wire _w10704_ ;
	wire _w10703_ ;
	wire _w10702_ ;
	wire _w10701_ ;
	wire _w10700_ ;
	wire _w10699_ ;
	wire _w10698_ ;
	wire _w10697_ ;
	wire _w10696_ ;
	wire _w10695_ ;
	wire _w10694_ ;
	wire _w10693_ ;
	wire _w10692_ ;
	wire _w10691_ ;
	wire _w10690_ ;
	wire _w10689_ ;
	wire _w10688_ ;
	wire _w10687_ ;
	wire _w10686_ ;
	wire _w10685_ ;
	wire _w10684_ ;
	wire _w10683_ ;
	wire _w10682_ ;
	wire _w10681_ ;
	wire _w10680_ ;
	wire _w10679_ ;
	wire _w10678_ ;
	wire _w10677_ ;
	wire _w10676_ ;
	wire _w10675_ ;
	wire _w10674_ ;
	wire _w10673_ ;
	wire _w10672_ ;
	wire _w10671_ ;
	wire _w10670_ ;
	wire _w10669_ ;
	wire _w10668_ ;
	wire _w10667_ ;
	wire _w10666_ ;
	wire _w10665_ ;
	wire _w10664_ ;
	wire _w10663_ ;
	wire _w10662_ ;
	wire _w10661_ ;
	wire _w10660_ ;
	wire _w10659_ ;
	wire _w10658_ ;
	wire _w10657_ ;
	wire _w10656_ ;
	wire _w10655_ ;
	wire _w10654_ ;
	wire _w10653_ ;
	wire _w10652_ ;
	wire _w10651_ ;
	wire _w10650_ ;
	wire _w10649_ ;
	wire _w10648_ ;
	wire _w10647_ ;
	wire _w10646_ ;
	wire _w10645_ ;
	wire _w10644_ ;
	wire _w10643_ ;
	wire _w10642_ ;
	wire _w10641_ ;
	wire _w10640_ ;
	wire _w10571_ ;
	wire _w10570_ ;
	wire _w10569_ ;
	wire _w10568_ ;
	wire _w10567_ ;
	wire _w10566_ ;
	wire _w10565_ ;
	wire _w10564_ ;
	wire _w10563_ ;
	wire _w10562_ ;
	wire _w10561_ ;
	wire _w10560_ ;
	wire _w10559_ ;
	wire _w10558_ ;
	wire _w10557_ ;
	wire _w10556_ ;
	wire _w10555_ ;
	wire _w10554_ ;
	wire _w10553_ ;
	wire _w10552_ ;
	wire _w10551_ ;
	wire _w10550_ ;
	wire _w10548_ ;
	wire _w10547_ ;
	wire _w10546_ ;
	wire _w10545_ ;
	wire _w10544_ ;
	wire _w10543_ ;
	wire _w10542_ ;
	wire _w10525_ ;
	wire _w10524_ ;
	wire _w10523_ ;
	wire _w10549_ ;
	wire _w10740_ ;
	wire _w10620_ ;
	wire _w10521_ ;
	wire _w10520_ ;
	wire _w10519_ ;
	wire _w10518_ ;
	wire _w10517_ ;
	wire _w10516_ ;
	wire _w10515_ ;
	wire _w10514_ ;
	wire _w10522_ ;
	wire _w10526_ ;
	wire _w10527_ ;
	wire _w10528_ ;
	wire _w10529_ ;
	wire _w10530_ ;
	wire _w10531_ ;
	wire _w10532_ ;
	wire _w10533_ ;
	wire _w10534_ ;
	wire _w10535_ ;
	wire _w10536_ ;
	wire _w10537_ ;
	wire _w10538_ ;
	wire _w10539_ ;
	wire _w10540_ ;
	wire _w10541_ ;
	wire _w10572_ ;
	wire _w10573_ ;
	wire _w10574_ ;
	wire _w10575_ ;
	wire _w10576_ ;
	wire _w10577_ ;
	wire _w10578_ ;
	wire _w10579_ ;
	wire _w10580_ ;
	wire _w10581_ ;
	wire _w10582_ ;
	wire _w10583_ ;
	wire _w10584_ ;
	wire _w10585_ ;
	wire _w10586_ ;
	wire _w10587_ ;
	wire _w10588_ ;
	wire _w10589_ ;
	wire _w10590_ ;
	wire _w10591_ ;
	wire _w10592_ ;
	wire _w10593_ ;
	wire _w10594_ ;
	wire _w10595_ ;
	wire _w10596_ ;
	wire _w10597_ ;
	wire _w10598_ ;
	wire _w10599_ ;
	wire _w10600_ ;
	wire _w10601_ ;
	wire _w10602_ ;
	wire _w10603_ ;
	wire _w10604_ ;
	wire _w10605_ ;
	wire _w10606_ ;
	wire _w10607_ ;
	wire _w10608_ ;
	wire _w10609_ ;
	wire _w10610_ ;
	wire _w10611_ ;
	wire _w10612_ ;
	wire _w10613_ ;
	wire _w10614_ ;
	wire _w10615_ ;
	wire _w10616_ ;
	wire _w10617_ ;
	wire _w10618_ ;
	wire _w10619_ ;
	wire _w10621_ ;
	wire _w10622_ ;
	wire _w10623_ ;
	wire _w10624_ ;
	wire _w10625_ ;
	wire _w10626_ ;
	wire _w10627_ ;
	wire _w10628_ ;
	wire _w10629_ ;
	wire _w10630_ ;
	wire _w10631_ ;
	wire _w10632_ ;
	wire _w10633_ ;
	wire _w10634_ ;
	wire _w10635_ ;
	wire _w10636_ ;
	wire _w10637_ ;
	wire _w10638_ ;
	wire _w10639_ ;
	wire _w10770_ ;
	wire _w10771_ ;
	wire _w10772_ ;
	wire _w10773_ ;
	wire _w10774_ ;
	wire _w10775_ ;
	wire _w10776_ ;
	wire _w10777_ ;
	wire _w10778_ ;
	wire _w10779_ ;
	wire _w10780_ ;
	wire _w10781_ ;
	wire _w10782_ ;
	wire _w10783_ ;
	wire _w10784_ ;
	wire _w10785_ ;
	wire _w10786_ ;
	wire _w10787_ ;
	wire _w10788_ ;
	wire _w10789_ ;
	wire _w10790_ ;
	wire _w10791_ ;
	wire _w10792_ ;
	wire _w10793_ ;
	wire _w10794_ ;
	wire _w10795_ ;
	wire _w10796_ ;
	wire _w10797_ ;
	wire _w10798_ ;
	wire _w10799_ ;
	wire _w10800_ ;
	wire _w10801_ ;
	wire _w10802_ ;
	wire _w10803_ ;
	wire _w10804_ ;
	wire _w10805_ ;
	wire _w10806_ ;
	wire _w10807_ ;
	wire _w10808_ ;
	wire _w10809_ ;
	wire _w10810_ ;
	wire _w10811_ ;
	wire _w10812_ ;
	wire _w10813_ ;
	wire _w10814_ ;
	wire _w10815_ ;
	wire _w10816_ ;
	wire _w10817_ ;
	wire _w10818_ ;
	wire _w10819_ ;
	wire _w10820_ ;
	wire _w10821_ ;
	wire _w10822_ ;
	wire _w10823_ ;
	wire _w10824_ ;
	wire _w10825_ ;
	wire _w10826_ ;
	wire _w10827_ ;
	wire _w10828_ ;
	wire _w10829_ ;
	wire _w10830_ ;
	wire _w10831_ ;
	wire _w10832_ ;
	wire _w10833_ ;
	wire _w10834_ ;
	wire _w10835_ ;
	wire _w10836_ ;
	wire _w10837_ ;
	wire _w10838_ ;
	wire _w10839_ ;
	wire _w10840_ ;
	wire _w10841_ ;
	wire _w10842_ ;
	wire _w10843_ ;
	wire _w10844_ ;
	wire _w10845_ ;
	wire _w10846_ ;
	wire _w10847_ ;
	wire _w10848_ ;
	wire _w10849_ ;
	wire _w10850_ ;
	wire _w10851_ ;
	wire _w10852_ ;
	wire _w10853_ ;
	wire _w10854_ ;
	wire _w10855_ ;
	wire _w10856_ ;
	wire _w10857_ ;
	wire _w10858_ ;
	wire _w10859_ ;
	wire _w10860_ ;
	wire _w10861_ ;
	wire _w10862_ ;
	wire _w10863_ ;
	wire _w10864_ ;
	wire _w10865_ ;
	wire _w10866_ ;
	wire _w10867_ ;
	wire _w10868_ ;
	wire _w10869_ ;
	wire _w10870_ ;
	wire _w10871_ ;
	wire _w10872_ ;
	wire _w10873_ ;
	wire _w10874_ ;
	wire _w10875_ ;
	wire _w10876_ ;
	wire _w10877_ ;
	wire _w10878_ ;
	wire _w10879_ ;
	wire _w10880_ ;
	wire _w10881_ ;
	wire _w10882_ ;
	wire _w10883_ ;
	wire _w10884_ ;
	wire _w10885_ ;
	wire _w10886_ ;
	wire _w10887_ ;
	wire _w10888_ ;
	wire _w10889_ ;
	wire _w10890_ ;
	wire _w10891_ ;
	wire _w10892_ ;
	wire _w10893_ ;
	wire _w10894_ ;
	wire _w10895_ ;
	wire _w10896_ ;
	wire _w10897_ ;
	wire _w10898_ ;
	wire _w10899_ ;
	wire _w10900_ ;
	wire _w10901_ ;
	wire _w10902_ ;
	wire _w10903_ ;
	wire _w10904_ ;
	wire _w10905_ ;
	wire _w10906_ ;
	wire _w10907_ ;
	wire _w10908_ ;
	wire _w10909_ ;
	wire _w10910_ ;
	wire _w10911_ ;
	wire _w10912_ ;
	wire _w10913_ ;
	wire _w10914_ ;
	wire _w10915_ ;
	wire _w10916_ ;
	wire _w10917_ ;
	wire _w10918_ ;
	wire _w10919_ ;
	wire _w10920_ ;
	wire _w10921_ ;
	wire _w10922_ ;
	wire _w10923_ ;
	wire _w10924_ ;
	wire _w10925_ ;
	wire _w10926_ ;
	wire _w10927_ ;
	wire _w10928_ ;
	wire _w10929_ ;
	wire _w10930_ ;
	wire _w10931_ ;
	wire _w10932_ ;
	wire _w10933_ ;
	wire _w10934_ ;
	wire _w10935_ ;
	wire _w10936_ ;
	wire _w10937_ ;
	wire _w10938_ ;
	wire _w10939_ ;
	wire _w10940_ ;
	wire _w10941_ ;
	wire _w10942_ ;
	wire _w10943_ ;
	wire _w10944_ ;
	wire _w10945_ ;
	wire _w10946_ ;
	wire _w10947_ ;
	wire _w10948_ ;
	wire _w10949_ ;
	wire _w10950_ ;
	wire _w10951_ ;
	wire _w10952_ ;
	wire _w10953_ ;
	wire _w10954_ ;
	wire _w10955_ ;
	wire _w10956_ ;
	wire _w10957_ ;
	wire _w10958_ ;
	wire _w10959_ ;
	wire _w10960_ ;
	wire _w10961_ ;
	wire _w10962_ ;
	wire _w10963_ ;
	wire _w10964_ ;
	wire _w10965_ ;
	wire _w10966_ ;
	wire _w10967_ ;
	wire _w10968_ ;
	wire _w10969_ ;
	wire _w10970_ ;
	wire _w10971_ ;
	wire _w10972_ ;
	wire _w10973_ ;
	wire _w10974_ ;
	wire _w10975_ ;
	wire _w10976_ ;
	wire _w10977_ ;
	wire _w10978_ ;
	wire _w10979_ ;
	wire _w10980_ ;
	wire _w10981_ ;
	wire _w10982_ ;
	wire _w10983_ ;
	wire _w10984_ ;
	wire _w10985_ ;
	wire _w10986_ ;
	wire _w10987_ ;
	wire _w10988_ ;
	wire _w10989_ ;
	wire _w10990_ ;
	wire _w10991_ ;
	wire _w10992_ ;
	wire _w10993_ ;
	wire _w10994_ ;
	wire _w10995_ ;
	wire _w10996_ ;
	wire _w10997_ ;
	wire _w10998_ ;
	wire _w10999_ ;
	wire _w11000_ ;
	wire _w11001_ ;
	wire _w11002_ ;
	wire _w11003_ ;
	wire _w11004_ ;
	wire _w11005_ ;
	wire _w11006_ ;
	wire _w11007_ ;
	wire _w11008_ ;
	wire _w11009_ ;
	wire _w11010_ ;
	wire _w11011_ ;
	wire _w11012_ ;
	wire _w11013_ ;
	wire _w11014_ ;
	wire _w11015_ ;
	wire _w11016_ ;
	wire _w11017_ ;
	wire _w11018_ ;
	wire _w11019_ ;
	wire _w11020_ ;
	wire _w11021_ ;
	wire _w11022_ ;
	wire _w11023_ ;
	wire _w11024_ ;
	wire _w11025_ ;
	wire _w11026_ ;
	wire _w11027_ ;
	wire _w11028_ ;
	wire _w11029_ ;
	wire _w11030_ ;
	wire _w11031_ ;
	wire _w11032_ ;
	wire _w11033_ ;
	wire _w11034_ ;
	wire _w11035_ ;
	wire _w11036_ ;
	wire _w11037_ ;
	wire _w11038_ ;
	wire _w11039_ ;
	wire _w11040_ ;
	wire _w11041_ ;
	wire _w11042_ ;
	wire _w11043_ ;
	wire _w11044_ ;
	wire _w11045_ ;
	wire _w11046_ ;
	wire _w11047_ ;
	wire _w11048_ ;
	wire _w11049_ ;
	wire _w11050_ ;
	wire _w11051_ ;
	wire _w11052_ ;
	wire _w11053_ ;
	wire _w11622_ ;
	wire _w11623_ ;
	wire _w11624_ ;
	wire _w11625_ ;
	wire _w11626_ ;
	wire _w11627_ ;
	wire _w11628_ ;
	wire _w11629_ ;
	wire _w11630_ ;
	wire _w11631_ ;
	wire _w11632_ ;
	wire _w11633_ ;
	wire _w11634_ ;
	wire _w11635_ ;
	wire _w11636_ ;
	wire _w11637_ ;
	wire _w11638_ ;
	wire _w11639_ ;
	wire _w11640_ ;
	wire _w11641_ ;
	wire _w11642_ ;
	wire _w11643_ ;
	wire _w11644_ ;
	wire _w11645_ ;
	wire _w11646_ ;
	wire _w11647_ ;
	wire _w11648_ ;
	wire _w11649_ ;
	wire _w11650_ ;
	wire _w11651_ ;
	wire _w11652_ ;
	wire _w11653_ ;
	wire _w11654_ ;
	wire _w11655_ ;
	wire _w11656_ ;
	wire _w11657_ ;
	wire _w11658_ ;
	wire _w11659_ ;
	wire _w11660_ ;
	wire _w11661_ ;
	wire _w11662_ ;
	wire _w11663_ ;
	wire _w11664_ ;
	wire _w11665_ ;
	wire _w11666_ ;
	wire _w11667_ ;
	wire _w11668_ ;
	wire _w11669_ ;
	wire _w11670_ ;
	wire _w11671_ ;
	wire _w11672_ ;
	wire _w11673_ ;
	wire _w11674_ ;
	wire _w11675_ ;
	wire _w11676_ ;
	wire _w11677_ ;
	wire _w11678_ ;
	wire _w11679_ ;
	wire _w11680_ ;
	wire _w11681_ ;
	wire _w11682_ ;
	wire _w11683_ ;
	wire _w11684_ ;
	wire _w11685_ ;
	wire _w11686_ ;
	wire _w11687_ ;
	wire _w11688_ ;
	wire _w11689_ ;
	wire _w11690_ ;
	wire _w11691_ ;
	wire _w11692_ ;
	wire _w11693_ ;
	wire _w11694_ ;
	wire _w11695_ ;
	wire _w11696_ ;
	wire _w11697_ ;
	wire _w11698_ ;
	wire _w11699_ ;
	wire _w11700_ ;
	wire _w11701_ ;
	wire _w11702_ ;
	wire _w11703_ ;
	wire _w11704_ ;
	wire _w11705_ ;
	wire _w11706_ ;
	wire _w11707_ ;
	wire _w11708_ ;
	wire _w11709_ ;
	wire _w11710_ ;
	wire _w11711_ ;
	wire _w11712_ ;
	wire _w11713_ ;
	wire _w11714_ ;
	wire _w11715_ ;
	wire _w11716_ ;
	wire _w11717_ ;
	wire _w11718_ ;
	wire _w11719_ ;
	wire _w11720_ ;
	wire _w11721_ ;
	wire _w11722_ ;
	wire _w11723_ ;
	wire _w11724_ ;
	wire _w11725_ ;
	wire _w11726_ ;
	wire _w11727_ ;
	wire _w11728_ ;
	wire _w11729_ ;
	wire _w11730_ ;
	wire _w11731_ ;
	wire _w11732_ ;
	wire _w11733_ ;
	wire _w11734_ ;
	wire _w11735_ ;
	wire _w11736_ ;
	wire _w11737_ ;
	wire _w11738_ ;
	wire _w11739_ ;
	wire _w11740_ ;
	wire _w11741_ ;
	wire _w11742_ ;
	wire _w11743_ ;
	wire _w11744_ ;
	wire _w11745_ ;
	wire _w11746_ ;
	wire _w11747_ ;
	wire _w11748_ ;
	wire _w11749_ ;
	wire _w11750_ ;
	wire _w11751_ ;
	wire _w11752_ ;
	wire _w11753_ ;
	wire _w11754_ ;
	wire _w11755_ ;
	wire _w11756_ ;
	wire _w11757_ ;
	wire _w11758_ ;
	wire _w11759_ ;
	wire _w11760_ ;
	wire _w11761_ ;
	wire _w11762_ ;
	wire _w11763_ ;
	wire _w11764_ ;
	wire _w11765_ ;
	wire _w11766_ ;
	wire _w11767_ ;
	wire _w11768_ ;
	wire _w11769_ ;
	wire _w11770_ ;
	wire _w11771_ ;
	wire _w11772_ ;
	wire _w11773_ ;
	wire _w11774_ ;
	wire _w11775_ ;
	wire _w11776_ ;
	wire _w11777_ ;
	wire _w11778_ ;
	wire _w11779_ ;
	wire _w11780_ ;
	wire _w11781_ ;
	wire _w11782_ ;
	wire _w11783_ ;
	wire _w11784_ ;
	wire _w11785_ ;
	wire _w11786_ ;
	wire _w11787_ ;
	wire _w11788_ ;
	wire _w11789_ ;
	wire _w11790_ ;
	wire _w11791_ ;
	wire _w11792_ ;
	wire _w11793_ ;
	wire _w11794_ ;
	wire _w11795_ ;
	wire _w11796_ ;
	wire _w11797_ ;
	wire _w11798_ ;
	wire _w11799_ ;
	wire _w11800_ ;
	wire _w11801_ ;
	wire _w11802_ ;
	wire _w11803_ ;
	wire _w11804_ ;
	wire _w11805_ ;
	wire _w11806_ ;
	wire _w11807_ ;
	wire _w11808_ ;
	wire _w11809_ ;
	wire _w11810_ ;
	wire _w11811_ ;
	wire _w11812_ ;
	wire _w11813_ ;
	wire _w11814_ ;
	wire _w11815_ ;
	wire _w11816_ ;
	wire _w11817_ ;
	wire _w11818_ ;
	wire _w11819_ ;
	wire _w11820_ ;
	wire _w11821_ ;
	wire _w11822_ ;
	wire _w11823_ ;
	wire _w11824_ ;
	wire _w11825_ ;
	wire _w11826_ ;
	wire _w11827_ ;
	wire _w11828_ ;
	wire _w11829_ ;
	wire _w11830_ ;
	wire _w11831_ ;
	wire _w11832_ ;
	wire _w11833_ ;
	wire _w11834_ ;
	wire _w11835_ ;
	wire _w11836_ ;
	wire _w11837_ ;
	wire _w11838_ ;
	wire _w11839_ ;
	wire _w11840_ ;
	wire _w11841_ ;
	wire _w11842_ ;
	wire _w11843_ ;
	wire _w11844_ ;
	wire _w11845_ ;
	wire _w11846_ ;
	wire _w11847_ ;
	wire _w11848_ ;
	wire _w11849_ ;
	wire _w11850_ ;
	wire _w11851_ ;
	wire _w11852_ ;
	wire _w11853_ ;
	wire _w11854_ ;
	wire _w11855_ ;
	wire _w11856_ ;
	wire _w11857_ ;
	wire _w11858_ ;
	wire _w11859_ ;
	wire _w11860_ ;
	wire _w11861_ ;
	wire _w11862_ ;
	wire _w11863_ ;
	wire _w11864_ ;
	wire _w11865_ ;
	wire _w11866_ ;
	wire _w11867_ ;
	wire _w11868_ ;
	wire _w11869_ ;
	wire _w11870_ ;
	wire _w11871_ ;
	wire _w11872_ ;
	wire _w11873_ ;
	wire _w11874_ ;
	wire _w11875_ ;
	wire _w11876_ ;
	wire _w11877_ ;
	wire _w11878_ ;
	wire _w11879_ ;
	wire _w11880_ ;
	wire _w11881_ ;
	wire _w11882_ ;
	wire _w11883_ ;
	wire _w11884_ ;
	wire _w11885_ ;
	wire _w11886_ ;
	wire _w11887_ ;
	wire _w11888_ ;
	wire _w11889_ ;
	wire _w11890_ ;
	wire _w11891_ ;
	wire _w11892_ ;
	wire _w11893_ ;
	wire _w11894_ ;
	wire _w11895_ ;
	wire _w11896_ ;
	wire _w11897_ ;
	wire _w11898_ ;
	wire _w11899_ ;
	wire _w11900_ ;
	wire _w11901_ ;
	wire _w11902_ ;
	wire _w11903_ ;
	wire _w11904_ ;
	wire _w11905_ ;
	wire _w11906_ ;
	wire _w11907_ ;
	wire _w11908_ ;
	wire _w11909_ ;
	wire _w11910_ ;
	wire _w11911_ ;
	wire _w11912_ ;
	wire _w11913_ ;
	wire _w11914_ ;
	wire _w11915_ ;
	wire _w11916_ ;
	wire _w11917_ ;
	wire _w11918_ ;
	wire _w11919_ ;
	wire _w11920_ ;
	wire _w11921_ ;
	wire _w11922_ ;
	wire _w11923_ ;
	wire _w11924_ ;
	wire _w11925_ ;
	wire _w11926_ ;
	wire _w11927_ ;
	wire _w11928_ ;
	wire _w11929_ ;
	wire _w11930_ ;
	wire _w11931_ ;
	wire _w11932_ ;
	wire _w11933_ ;
	wire _w11934_ ;
	wire _w11935_ ;
	wire _w11936_ ;
	wire _w11937_ ;
	wire _w11938_ ;
	wire _w11939_ ;
	wire _w11940_ ;
	wire _w11941_ ;
	wire _w11942_ ;
	wire _w11943_ ;
	wire _w11944_ ;
	wire _w11945_ ;
	wire _w11946_ ;
	wire _w11947_ ;
	wire _w11948_ ;
	wire _w11949_ ;
	wire _w11950_ ;
	wire _w11951_ ;
	wire _w11952_ ;
	wire _w11953_ ;
	wire _w11954_ ;
	wire _w11955_ ;
	wire _w11956_ ;
	wire _w11957_ ;
	wire _w11958_ ;
	wire _w11959_ ;
	wire _w11960_ ;
	wire _w11961_ ;
	wire _w11962_ ;
	wire _w11963_ ;
	wire _w11964_ ;
	wire _w11965_ ;
	wire _w11966_ ;
	wire _w11967_ ;
	wire _w11968_ ;
	wire _w11969_ ;
	wire _w11970_ ;
	wire _w11971_ ;
	wire _w11972_ ;
	wire _w11973_ ;
	wire _w11974_ ;
	wire _w11975_ ;
	wire _w11976_ ;
	wire _w11977_ ;
	wire _w11978_ ;
	wire _w11979_ ;
	wire _w11980_ ;
	wire _w11981_ ;
	wire _w11982_ ;
	wire _w11983_ ;
	wire _w11984_ ;
	wire _w11985_ ;
	wire _w11986_ ;
	wire _w11987_ ;
	wire _w11988_ ;
	wire _w11989_ ;
	wire _w11990_ ;
	wire _w11991_ ;
	wire _w11992_ ;
	wire _w11993_ ;
	wire _w11994_ ;
	wire _w11995_ ;
	wire _w11996_ ;
	wire _w11997_ ;
	wire _w11998_ ;
	wire _w11999_ ;
	wire _w12000_ ;
	wire _w12001_ ;
	wire _w12002_ ;
	wire _w12003_ ;
	wire _w12004_ ;
	wire _w12005_ ;
	wire _w12006_ ;
	wire _w12007_ ;
	wire _w12008_ ;
	wire _w12009_ ;
	wire _w12010_ ;
	wire _w12011_ ;
	wire _w12012_ ;
	wire _w12013_ ;
	wire _w12014_ ;
	wire _w12015_ ;
	wire _w12016_ ;
	wire _w12017_ ;
	wire _w12018_ ;
	wire _w12019_ ;
	wire _w12020_ ;
	wire _w12021_ ;
	wire _w12022_ ;
	wire _w12023_ ;
	wire _w12024_ ;
	wire _w12025_ ;
	wire _w12026_ ;
	wire _w12027_ ;
	wire _w12028_ ;
	wire _w12029_ ;
	wire _w12030_ ;
	wire _w12031_ ;
	wire _w12032_ ;
	wire _w12033_ ;
	wire _w12034_ ;
	wire _w12035_ ;
	wire _w12036_ ;
	wire _w12037_ ;
	wire _w12038_ ;
	wire _w12039_ ;
	wire _w12040_ ;
	wire _w12041_ ;
	wire _w12042_ ;
	wire _w12043_ ;
	wire _w12044_ ;
	wire _w12045_ ;
	wire _w12046_ ;
	wire _w12047_ ;
	wire _w12048_ ;
	wire _w12049_ ;
	wire _w12050_ ;
	wire _w12051_ ;
	wire _w12052_ ;
	wire _w12053_ ;
	wire _w12054_ ;
	wire _w12055_ ;
	wire _w12056_ ;
	wire _w12057_ ;
	wire _w12058_ ;
	wire _w12059_ ;
	wire _w12060_ ;
	wire _w12061_ ;
	wire _w12062_ ;
	wire _w12063_ ;
	wire _w12064_ ;
	wire _w12065_ ;
	wire _w12066_ ;
	wire _w12067_ ;
	wire _w12068_ ;
	wire _w12069_ ;
	wire _w12070_ ;
	wire _w12071_ ;
	wire _w12072_ ;
	wire _w12073_ ;
	wire _w12074_ ;
	wire _w12075_ ;
	wire _w12076_ ;
	wire _w12077_ ;
	wire _w12078_ ;
	wire _w12079_ ;
	wire _w12080_ ;
	wire _w12081_ ;
	wire _w12082_ ;
	wire _w12083_ ;
	wire _w12084_ ;
	wire _w12085_ ;
	wire _w12086_ ;
	wire _w12087_ ;
	wire _w12088_ ;
	wire _w12089_ ;
	wire _w12090_ ;
	wire _w12091_ ;
	wire _w12092_ ;
	wire _w12093_ ;
	wire _w12094_ ;
	wire _w12095_ ;
	wire _w12096_ ;
	wire _w12097_ ;
	wire _w12098_ ;
	wire _w12099_ ;
	wire _w12100_ ;
	wire _w12101_ ;
	wire _w12102_ ;
	wire _w12103_ ;
	wire _w12104_ ;
	wire _w12105_ ;
	wire _w12106_ ;
	wire _w12107_ ;
	wire _w12108_ ;
	wire _w12109_ ;
	wire _w12110_ ;
	wire _w12111_ ;
	wire _w12112_ ;
	wire _w12113_ ;
	wire _w12114_ ;
	wire _w12115_ ;
	wire _w12116_ ;
	wire _w12117_ ;
	wire _w12118_ ;
	wire _w12119_ ;
	wire _w12120_ ;
	wire _w12121_ ;
	wire _w12122_ ;
	wire _w12123_ ;
	wire _w12124_ ;
	wire _w12125_ ;
	wire _w12126_ ;
	wire _w12127_ ;
	wire _w12128_ ;
	wire _w12129_ ;
	wire _w12130_ ;
	wire _w12131_ ;
	wire _w12132_ ;
	wire _w12133_ ;
	wire _w12134_ ;
	wire _w12135_ ;
	wire _w12136_ ;
	wire _w12137_ ;
	wire _w12138_ ;
	wire _w12139_ ;
	wire _w12140_ ;
	wire _w12141_ ;
	wire _w12142_ ;
	wire _w12143_ ;
	wire _w12144_ ;
	wire _w12145_ ;
	wire _w12146_ ;
	wire _w12147_ ;
	wire _w12148_ ;
	wire _w12149_ ;
	wire _w12150_ ;
	wire _w12151_ ;
	wire _w12152_ ;
	wire _w12153_ ;
	wire _w12154_ ;
	wire _w12155_ ;
	wire _w12156_ ;
	wire _w12157_ ;
	wire _w12158_ ;
	wire _w12159_ ;
	wire _w12160_ ;
	wire _w12161_ ;
	wire _w12162_ ;
	wire _w12163_ ;
	wire _w12164_ ;
	wire _w12165_ ;
	wire _w12166_ ;
	wire _w12167_ ;
	wire _w12168_ ;
	wire _w12169_ ;
	wire _w12170_ ;
	wire _w12171_ ;
	wire _w12172_ ;
	wire _w12173_ ;
	wire _w12174_ ;
	wire _w12175_ ;
	wire _w12176_ ;
	wire _w12177_ ;
	wire _w12178_ ;
	wire _w12179_ ;
	wire _w12180_ ;
	wire _w12181_ ;
	wire _w12182_ ;
	wire _w12183_ ;
	wire _w12184_ ;
	wire _w12185_ ;
	wire _w12186_ ;
	wire _w12187_ ;
	wire _w12188_ ;
	wire _w12189_ ;
	wire _w12190_ ;
	wire _w12191_ ;
	wire _w12192_ ;
	wire _w12193_ ;
	wire _w12194_ ;
	wire _w12195_ ;
	wire _w12196_ ;
	wire _w12197_ ;
	wire _w12198_ ;
	wire _w12199_ ;
	wire _w12200_ ;
	wire _w12201_ ;
	wire _w12202_ ;
	wire _w12203_ ;
	wire _w12204_ ;
	wire _w12205_ ;
	wire _w12206_ ;
	wire _w12207_ ;
	wire _w12208_ ;
	wire _w12209_ ;
	wire _w12210_ ;
	wire _w12211_ ;
	wire _w12212_ ;
	wire _w12213_ ;
	wire _w12214_ ;
	wire _w12215_ ;
	wire _w12216_ ;
	wire _w12217_ ;
	wire _w12218_ ;
	wire _w12219_ ;
	wire _w12220_ ;
	wire _w12221_ ;
	wire _w12222_ ;
	wire _w12223_ ;
	wire _w12224_ ;
	wire _w12225_ ;
	wire _w12226_ ;
	wire _w12227_ ;
	wire _w12228_ ;
	wire _w12229_ ;
	wire _w12230_ ;
	wire _w12231_ ;
	wire _w12232_ ;
	wire _w12233_ ;
	wire _w12234_ ;
	wire _w12235_ ;
	wire _w12236_ ;
	wire _w12237_ ;
	wire _w12238_ ;
	wire _w12239_ ;
	wire _w12240_ ;
	wire _w12241_ ;
	wire _w12242_ ;
	wire _w12243_ ;
	wire _w12244_ ;
	wire _w12246_ ;
	wire _w12247_ ;
	wire _w12248_ ;
	wire _w12249_ ;
	wire _w12250_ ;
	wire _w12251_ ;
	wire _w12252_ ;
	wire _w12253_ ;
	wire _w12254_ ;
	wire _w12255_ ;
	wire _w12256_ ;
	wire _w12257_ ;
	wire _w12258_ ;
	wire _w12259_ ;
	wire _w12260_ ;
	wire _w12261_ ;
	wire _w12262_ ;
	wire _w12263_ ;
	wire _w12264_ ;
	wire _w12265_ ;
	wire _w12266_ ;
	wire _w12267_ ;
	wire _w12268_ ;
	wire _w12269_ ;
	wire _w12270_ ;
	wire _w12271_ ;
	wire _w12272_ ;
	wire _w12273_ ;
	wire _w12274_ ;
	wire _w12275_ ;
	wire _w12276_ ;
	wire _w12277_ ;
	wire _w12278_ ;
	wire _w12279_ ;
	wire _w12280_ ;
	wire _w12281_ ;
	wire _w12282_ ;
	wire _w12283_ ;
	wire _w12284_ ;
	wire _w12285_ ;
	wire _w12286_ ;
	wire _w12287_ ;
	wire _w12288_ ;
	wire _w12289_ ;
	wire _w12290_ ;
	wire _w12291_ ;
	wire _w12292_ ;
	wire _w12293_ ;
	wire _w12294_ ;
	wire _w12295_ ;
	wire _w12296_ ;
	wire _w12297_ ;
	wire _w12298_ ;
	wire _w12299_ ;
	wire _w12300_ ;
	wire _w12301_ ;
	wire _w12302_ ;
	wire _w12303_ ;
	wire _w12304_ ;
	wire _w12305_ ;
	wire _w12306_ ;
	wire _w12307_ ;
	wire _w12308_ ;
	wire _w12309_ ;
	wire _w12310_ ;
	wire _w12311_ ;
	wire _w12312_ ;
	wire _w12313_ ;
	wire _w12314_ ;
	wire _w12315_ ;
	wire _w12316_ ;
	wire _w12317_ ;
	wire _w12318_ ;
	wire _w12319_ ;
	wire _w12320_ ;
	wire _w12321_ ;
	wire _w12322_ ;
	wire _w12323_ ;
	wire _w12324_ ;
	wire _w12325_ ;
	wire _w12326_ ;
	wire _w12327_ ;
	wire _w12328_ ;
	wire _w12329_ ;
	wire _w12330_ ;
	wire _w12331_ ;
	wire _w12332_ ;
	wire _w12333_ ;
	wire _w12334_ ;
	wire _w12335_ ;
	wire _w12336_ ;
	wire _w12337_ ;
	wire _w12338_ ;
	wire _w12339_ ;
	wire _w12340_ ;
	wire _w12341_ ;
	wire _w12342_ ;
	wire _w12343_ ;
	wire _w12344_ ;
	wire _w12345_ ;
	wire _w12346_ ;
	wire _w12347_ ;
	wire _w12348_ ;
	wire _w12349_ ;
	wire _w12350_ ;
	wire _w12351_ ;
	wire _w12352_ ;
	wire _w12353_ ;
	wire _w12354_ ;
	wire _w12355_ ;
	wire _w12356_ ;
	wire _w12357_ ;
	wire _w12358_ ;
	wire _w12359_ ;
	wire _w12360_ ;
	wire _w12361_ ;
	wire _w12362_ ;
	wire _w12363_ ;
	wire _w12364_ ;
	wire _w12365_ ;
	wire _w12366_ ;
	wire _w12367_ ;
	wire _w12368_ ;
	wire _w12369_ ;
	wire _w12370_ ;
	wire _w12371_ ;
	wire _w12372_ ;
	wire _w12373_ ;
	wire _w12374_ ;
	wire _w12375_ ;
	wire _w12376_ ;
	wire _w12377_ ;
	wire _w12378_ ;
	wire _w12379_ ;
	wire _w12380_ ;
	wire _w12381_ ;
	wire _w12382_ ;
	wire _w12383_ ;
	wire _w12384_ ;
	wire _w12385_ ;
	wire _w12386_ ;
	wire _w12387_ ;
	wire _w12388_ ;
	wire _w12389_ ;
	wire _w12390_ ;
	wire _w12391_ ;
	wire _w12392_ ;
	wire _w12393_ ;
	wire _w12394_ ;
	wire _w12395_ ;
	wire _w12396_ ;
	wire _w12397_ ;
	wire _w12398_ ;
	wire _w12399_ ;
	wire _w12400_ ;
	wire _w12401_ ;
	wire _w12402_ ;
	wire _w12403_ ;
	wire _w12404_ ;
	wire _w12405_ ;
	wire _w12406_ ;
	wire _w12407_ ;
	wire _w12408_ ;
	wire _w12409_ ;
	wire _w12410_ ;
	wire _w12411_ ;
	wire _w12412_ ;
	wire _w12413_ ;
	wire _w12414_ ;
	wire _w12415_ ;
	wire _w12416_ ;
	wire _w12417_ ;
	wire _w12418_ ;
	wire _w12419_ ;
	wire _w12420_ ;
	wire _w12421_ ;
	wire _w12422_ ;
	wire _w12423_ ;
	wire _w12424_ ;
	wire _w12425_ ;
	wire _w12426_ ;
	wire _w12427_ ;
	wire _w12428_ ;
	wire _w12429_ ;
	wire _w12430_ ;
	wire _w12431_ ;
	wire _w12432_ ;
	wire _w12433_ ;
	wire _w12434_ ;
	wire _w12435_ ;
	wire _w12436_ ;
	wire _w12437_ ;
	wire _w12438_ ;
	wire _w12439_ ;
	wire _w12440_ ;
	wire _w12441_ ;
	wire _w12442_ ;
	wire _w12443_ ;
	wire _w12444_ ;
	wire _w12445_ ;
	wire _w12446_ ;
	wire _w12447_ ;
	wire _w12448_ ;
	wire _w12449_ ;
	wire _w12450_ ;
	wire _w12451_ ;
	wire _w12452_ ;
	wire _w12453_ ;
	wire _w12454_ ;
	wire _w12455_ ;
	wire _w12456_ ;
	wire _w12457_ ;
	wire _w12458_ ;
	wire _w12459_ ;
	wire _w12460_ ;
	wire _w12461_ ;
	wire _w12462_ ;
	wire _w12463_ ;
	wire _w12464_ ;
	wire _w12465_ ;
	wire _w12466_ ;
	wire _w12467_ ;
	wire _w12468_ ;
	wire _w12469_ ;
	wire _w12470_ ;
	wire _w12471_ ;
	wire _w12472_ ;
	wire _w12473_ ;
	wire _w12474_ ;
	wire _w12475_ ;
	wire _w12476_ ;
	wire _w12477_ ;
	wire _w12478_ ;
	wire _w12479_ ;
	wire _w12480_ ;
	wire _w12481_ ;
	wire _w12482_ ;
	wire _w12483_ ;
	wire _w12484_ ;
	wire _w12485_ ;
	wire _w12486_ ;
	wire _w12487_ ;
	wire _w12488_ ;
	wire _w12489_ ;
	wire _w12490_ ;
	wire _w12491_ ;
	wire _w12492_ ;
	wire _w12493_ ;
	wire _w12494_ ;
	wire _w12495_ ;
	wire _w12496_ ;
	wire _w12497_ ;
	wire _w12498_ ;
	wire _w12499_ ;
	wire _w12500_ ;
	wire _w12501_ ;
	wire _w12502_ ;
	wire _w12503_ ;
	wire _w12504_ ;
	wire _w12505_ ;
	wire _w12506_ ;
	wire _w12507_ ;
	wire _w12508_ ;
	wire _w12509_ ;
	wire _w12510_ ;
	wire _w12511_ ;
	wire _w12512_ ;
	wire _w12513_ ;
	wire _w12514_ ;
	wire _w12515_ ;
	wire _w12516_ ;
	wire _w12517_ ;
	wire _w12518_ ;
	wire _w12519_ ;
	wire _w12520_ ;
	wire _w12521_ ;
	wire _w12522_ ;
	wire _w12523_ ;
	wire _w12524_ ;
	wire _w12525_ ;
	wire _w12526_ ;
	wire _w12527_ ;
	wire _w12528_ ;
	wire _w12529_ ;
	wire _w12530_ ;
	wire _w12531_ ;
	wire _w12532_ ;
	wire _w12533_ ;
	wire _w12534_ ;
	wire _w12535_ ;
	wire _w12536_ ;
	wire _w12537_ ;
	wire _w12538_ ;
	wire _w12539_ ;
	wire _w12540_ ;
	wire _w12541_ ;
	wire _w12542_ ;
	wire _w12543_ ;
	wire _w12544_ ;
	wire _w12545_ ;
	wire _w12546_ ;
	wire _w12547_ ;
	wire _w12548_ ;
	wire _w12549_ ;
	wire _w12550_ ;
	wire _w12551_ ;
	wire _w12552_ ;
	wire _w12553_ ;
	wire _w12554_ ;
	wire _w12555_ ;
	wire _w12556_ ;
	wire _w12557_ ;
	wire _w12558_ ;
	wire _w12559_ ;
	wire _w12560_ ;
	wire _w12561_ ;
	wire _w12562_ ;
	wire _w12563_ ;
	wire _w12564_ ;
	wire _w12565_ ;
	wire _w12566_ ;
	wire _w12567_ ;
	wire _w12568_ ;
	wire _w12569_ ;
	wire _w12570_ ;
	wire _w12571_ ;
	wire _w12572_ ;
	wire _w12573_ ;
	wire _w12574_ ;
	wire _w12575_ ;
	wire _w12576_ ;
	wire _w12577_ ;
	wire _w12578_ ;
	wire _w12579_ ;
	wire _w12580_ ;
	wire _w12581_ ;
	wire _w12582_ ;
	wire _w12583_ ;
	wire _w12584_ ;
	wire _w12585_ ;
	wire _w12586_ ;
	wire _w12587_ ;
	wire _w12588_ ;
	wire _w12589_ ;
	wire _w12590_ ;
	wire _w12591_ ;
	wire _w12592_ ;
	wire _w12593_ ;
	wire _w12594_ ;
	wire _w12595_ ;
	wire _w12596_ ;
	wire _w12597_ ;
	wire _w12598_ ;
	wire _w12599_ ;
	wire _w12600_ ;
	wire _w12601_ ;
	wire _w12602_ ;
	wire _w12603_ ;
	wire _w12604_ ;
	wire _w12605_ ;
	wire _w12606_ ;
	wire _w12607_ ;
	wire _w12608_ ;
	wire _w12609_ ;
	wire _w12610_ ;
	wire _w12611_ ;
	wire _w12612_ ;
	wire _w12613_ ;
	wire _w12614_ ;
	wire _w12615_ ;
	wire _w12616_ ;
	wire _w12617_ ;
	wire _w12618_ ;
	wire _w12619_ ;
	wire _w12620_ ;
	wire _w12621_ ;
	wire _w12622_ ;
	wire _w12623_ ;
	wire _w12624_ ;
	wire _w12625_ ;
	wire _w12626_ ;
	wire _w12627_ ;
	wire _w12628_ ;
	wire _w12629_ ;
	wire _w12630_ ;
	wire _w12631_ ;
	wire _w12632_ ;
	wire _w12633_ ;
	wire _w12634_ ;
	wire _w12635_ ;
	wire _w12636_ ;
	wire _w12637_ ;
	wire _w12638_ ;
	wire _w12639_ ;
	wire _w12640_ ;
	wire _w12641_ ;
	wire _w12642_ ;
	wire _w12643_ ;
	wire _w12644_ ;
	wire _w12645_ ;
	wire _w12646_ ;
	wire _w12647_ ;
	wire _w12648_ ;
	wire _w12649_ ;
	wire _w12650_ ;
	wire _w12651_ ;
	wire _w12652_ ;
	wire _w12653_ ;
	wire _w12654_ ;
	wire _w12655_ ;
	wire _w12656_ ;
	wire _w12657_ ;
	wire _w12658_ ;
	wire _w12659_ ;
	wire _w12660_ ;
	wire _w12661_ ;
	wire _w12662_ ;
	wire _w12663_ ;
	wire _w12664_ ;
	wire _w12665_ ;
	wire _w12666_ ;
	wire _w12667_ ;
	wire _w12668_ ;
	wire _w12669_ ;
	wire _w12670_ ;
	wire _w12671_ ;
	wire _w12672_ ;
	wire _w12673_ ;
	wire _w12674_ ;
	wire _w12675_ ;
	wire _w12676_ ;
	wire _w12677_ ;
	wire _w12678_ ;
	wire _w12679_ ;
	wire _w12680_ ;
	wire _w12681_ ;
	wire _w12682_ ;
	wire _w12683_ ;
	wire _w12684_ ;
	wire _w12685_ ;
	wire _w12686_ ;
	wire _w12687_ ;
	wire _w12688_ ;
	wire _w12689_ ;
	wire _w12690_ ;
	wire _w12691_ ;
	wire _w12692_ ;
	wire _w12693_ ;
	wire _w12694_ ;
	wire _w12695_ ;
	wire _w12696_ ;
	wire _w12697_ ;
	wire _w12698_ ;
	wire _w12699_ ;
	wire _w12700_ ;
	wire _w12701_ ;
	wire _w12702_ ;
	wire _w12703_ ;
	wire _w12704_ ;
	wire _w12705_ ;
	wire _w12706_ ;
	wire _w12707_ ;
	wire _w12708_ ;
	wire _w12709_ ;
	wire _w12710_ ;
	wire _w12711_ ;
	wire _w12712_ ;
	wire _w12713_ ;
	wire _w12714_ ;
	wire _w12715_ ;
	wire _w12716_ ;
	wire _w12717_ ;
	wire _w12718_ ;
	wire _w12719_ ;
	wire _w12720_ ;
	wire _w12721_ ;
	wire _w12722_ ;
	wire _w12723_ ;
	wire _w12724_ ;
	wire _w12725_ ;
	wire _w12726_ ;
	wire _w12727_ ;
	wire _w12728_ ;
	wire _w12729_ ;
	wire _w12730_ ;
	wire _w12731_ ;
	wire _w12732_ ;
	wire _w12733_ ;
	wire _w12734_ ;
	wire _w12735_ ;
	wire _w12736_ ;
	wire _w12737_ ;
	wire _w12738_ ;
	wire _w12739_ ;
	wire _w12740_ ;
	wire _w12741_ ;
	wire _w12742_ ;
	wire _w12743_ ;
	wire _w12744_ ;
	wire _w12745_ ;
	wire _w12746_ ;
	wire _w12747_ ;
	wire _w12748_ ;
	wire _w12749_ ;
	wire _w12750_ ;
	wire _w12751_ ;
	wire _w12752_ ;
	wire _w12753_ ;
	wire _w12754_ ;
	wire _w12755_ ;
	wire _w12756_ ;
	wire _w12757_ ;
	wire _w12758_ ;
	wire _w12759_ ;
	wire _w12760_ ;
	wire _w12761_ ;
	wire _w12762_ ;
	wire _w12763_ ;
	wire _w12764_ ;
	wire _w12765_ ;
	wire _w12766_ ;
	wire _w12767_ ;
	wire _w12768_ ;
	wire _w12769_ ;
	wire _w12770_ ;
	wire _w12771_ ;
	wire _w12772_ ;
	wire _w12773_ ;
	wire _w12774_ ;
	wire _w12775_ ;
	wire _w12776_ ;
	wire _w12777_ ;
	wire _w12778_ ;
	wire _w12779_ ;
	wire _w12780_ ;
	wire _w12781_ ;
	wire _w12782_ ;
	wire _w12783_ ;
	wire _w12784_ ;
	wire _w12785_ ;
	wire _w12786_ ;
	wire _w12787_ ;
	wire _w12788_ ;
	wire _w12789_ ;
	wire _w12790_ ;
	wire _w12791_ ;
	wire _w12792_ ;
	wire _w12793_ ;
	wire _w12794_ ;
	wire _w12795_ ;
	wire _w12796_ ;
	wire _w12797_ ;
	wire _w12798_ ;
	wire _w12799_ ;
	wire _w12800_ ;
	wire _w12801_ ;
	wire _w12802_ ;
	wire _w12803_ ;
	wire _w12804_ ;
	wire _w12805_ ;
	wire _w12806_ ;
	wire _w12807_ ;
	wire _w12808_ ;
	wire _w12809_ ;
	wire _w12810_ ;
	wire _w12811_ ;
	wire _w12812_ ;
	wire _w12813_ ;
	wire _w12814_ ;
	wire _w12815_ ;
	wire _w12816_ ;
	wire _w12817_ ;
	wire _w12818_ ;
	wire _w12819_ ;
	wire _w12820_ ;
	wire _w12821_ ;
	wire _w12822_ ;
	wire _w12823_ ;
	wire _w12824_ ;
	wire _w12825_ ;
	wire _w12826_ ;
	wire _w12827_ ;
	wire _w12828_ ;
	wire _w12829_ ;
	wire _w12830_ ;
	wire _w12831_ ;
	wire _w12832_ ;
	wire _w12833_ ;
	wire _w12834_ ;
	wire _w12835_ ;
	wire _w12836_ ;
	wire _w12837_ ;
	wire _w12838_ ;
	wire _w12839_ ;
	wire _w12840_ ;
	wire _w12841_ ;
	wire _w12842_ ;
	wire _w12843_ ;
	wire _w12844_ ;
	wire _w12845_ ;
	wire _w12846_ ;
	wire _w12847_ ;
	wire _w12848_ ;
	wire _w12849_ ;
	wire _w12850_ ;
	wire _w12851_ ;
	wire _w12852_ ;
	wire _w12853_ ;
	wire _w12854_ ;
	wire _w12855_ ;
	wire _w12856_ ;
	wire _w12857_ ;
	wire _w12858_ ;
	wire _w12859_ ;
	wire _w12860_ ;
	wire _w12861_ ;
	wire _w12862_ ;
	wire _w12863_ ;
	wire _w12864_ ;
	wire _w12865_ ;
	wire _w12866_ ;
	wire _w12867_ ;
	wire _w12868_ ;
	wire _w12869_ ;
	wire _w15600_ ;
	wire _w15601_ ;
	wire _w15602_ ;
	wire _w15603_ ;
	wire _w15604_ ;
	wire _w15605_ ;
	wire _w15606_ ;
	wire _w15607_ ;
	wire _w15608_ ;
	wire _w15609_ ;
	wire _w15610_ ;
	wire _w15611_ ;
	wire _w15612_ ;
	wire _w15613_ ;
	wire _w15614_ ;
	wire _w15615_ ;
	wire _w15616_ ;
	wire _w15617_ ;
	wire _w15618_ ;
	wire _w15619_ ;
	wire _w15620_ ;
	wire _w15621_ ;
	wire _w15622_ ;
	wire _w15623_ ;
	wire _w15624_ ;
	wire _w15625_ ;
	wire _w15626_ ;
	wire _w15627_ ;
	wire _w15628_ ;
	wire _w15629_ ;
	wire _w15630_ ;
	wire _w15631_ ;
	wire _w15632_ ;
	wire _w15633_ ;
	wire _w15634_ ;
	wire _w15635_ ;
	wire _w15636_ ;
	wire _w15637_ ;
	wire _w15638_ ;
	wire _w15639_ ;
	wire _w15640_ ;
	wire _w15641_ ;
	wire _w15642_ ;
	wire _w15643_ ;
	wire _w15644_ ;
	wire _w15645_ ;
	wire _w15646_ ;
	wire _w15647_ ;
	wire _w15648_ ;
	wire _w15649_ ;
	wire _w15650_ ;
	wire _w15651_ ;
	wire _w15652_ ;
	wire _w15653_ ;
	wire _w15654_ ;
	wire _w15655_ ;
	wire _w15656_ ;
	wire _w15657_ ;
	wire _w15658_ ;
	wire _w15659_ ;
	wire _w15660_ ;
	wire _w15661_ ;
	wire _w15662_ ;
	wire _w15663_ ;
	wire _w15664_ ;
	wire _w15665_ ;
	wire _w15666_ ;
	wire _w15667_ ;
	wire _w15668_ ;
	wire _w15669_ ;
	wire _w15670_ ;
	wire _w15671_ ;
	wire _w15672_ ;
	wire _w15673_ ;
	wire _w15674_ ;
	wire _w15675_ ;
	wire _w15676_ ;
	wire _w15677_ ;
	wire _w15678_ ;
	wire _w15679_ ;
	wire _w15680_ ;
	wire _w15681_ ;
	wire _w15682_ ;
	wire _w15683_ ;
	wire _w15684_ ;
	wire _w15685_ ;
	wire _w15686_ ;
	wire _w15687_ ;
	wire _w15688_ ;
	wire _w15689_ ;
	wire _w15690_ ;
	wire _w15691_ ;
	wire _w15692_ ;
	wire _w15693_ ;
	wire _w15694_ ;
	wire _w15695_ ;
	wire _w15696_ ;
	wire _w15697_ ;
	wire _w15698_ ;
	wire _w15699_ ;
	wire _w15700_ ;
	wire _w15701_ ;
	wire _w15702_ ;
	wire _w15703_ ;
	wire _w15704_ ;
	wire _w15705_ ;
	wire _w15706_ ;
	wire _w15707_ ;
	wire _w15708_ ;
	wire _w15709_ ;
	wire _w15710_ ;
	wire _w15711_ ;
	wire _w15712_ ;
	wire _w15713_ ;
	wire _w15714_ ;
	wire _w15715_ ;
	wire _w15716_ ;
	wire _w15717_ ;
	wire _w15718_ ;
	wire _w15719_ ;
	wire _w15720_ ;
	wire _w15721_ ;
	wire _w15722_ ;
	wire _w15723_ ;
	wire _w15724_ ;
	wire _w15725_ ;
	wire _w15726_ ;
	wire _w15727_ ;
	wire _w15728_ ;
	wire _w15729_ ;
	wire _w15730_ ;
	wire _w15731_ ;
	wire _w15732_ ;
	wire _w15733_ ;
	wire _w15734_ ;
	wire _w15735_ ;
	wire _w15736_ ;
	wire _w15737_ ;
	wire _w15738_ ;
	wire _w15739_ ;
	wire _w15740_ ;
	wire _w15741_ ;
	wire _w15742_ ;
	wire _w15743_ ;
	wire _w15744_ ;
	wire _w15745_ ;
	wire _w15746_ ;
	wire _w15747_ ;
	wire _w15748_ ;
	wire _w15749_ ;
	wire _w15750_ ;
	wire _w15751_ ;
	wire _w15752_ ;
	wire _w15753_ ;
	wire _w15754_ ;
	wire _w15755_ ;
	wire _w15756_ ;
	wire _w15757_ ;
	wire _w15758_ ;
	wire _w15759_ ;
	wire _w15760_ ;
	wire _w15761_ ;
	wire _w15762_ ;
	wire _w15763_ ;
	wire _w15764_ ;
	wire _w15765_ ;
	wire _w15766_ ;
	wire _w15767_ ;
	wire _w15768_ ;
	wire _w15769_ ;
	wire _w15770_ ;
	wire _w15771_ ;
	wire _w15772_ ;
	wire _w15773_ ;
	wire _w15774_ ;
	wire _w15775_ ;
	wire _w15776_ ;
	wire _w15777_ ;
	wire _w15778_ ;
	wire _w15779_ ;
	wire _w15780_ ;
	wire _w15781_ ;
	wire _w15782_ ;
	wire _w15783_ ;
	wire _w15784_ ;
	wire _w15785_ ;
	wire _w15786_ ;
	wire _w15787_ ;
	wire _w15788_ ;
	wire _w15789_ ;
	wire _w15790_ ;
	wire _w15791_ ;
	wire _w15792_ ;
	wire _w15793_ ;
	wire _w15794_ ;
	wire _w15795_ ;
	wire _w15796_ ;
	wire _w15797_ ;
	wire _w15798_ ;
	wire _w15799_ ;
	wire _w15800_ ;
	wire _w15801_ ;
	wire _w15802_ ;
	wire _w15803_ ;
	wire _w15804_ ;
	wire _w15805_ ;
	wire _w15806_ ;
	wire _w15807_ ;
	wire _w15808_ ;
	wire _w15809_ ;
	wire _w15810_ ;
	wire _w15811_ ;
	wire _w15812_ ;
	wire _w15813_ ;
	wire _w15814_ ;
	wire _w15815_ ;
	wire _w15816_ ;
	wire _w15817_ ;
	wire _w15818_ ;
	wire _w15819_ ;
	wire _w15820_ ;
	wire _w15821_ ;
	wire _w15822_ ;
	wire _w15823_ ;
	wire _w15824_ ;
	wire _w15825_ ;
	wire _w15826_ ;
	wire _w15827_ ;
	wire _w15828_ ;
	wire _w15829_ ;
	wire _w15830_ ;
	wire _w15831_ ;
	wire _w15832_ ;
	wire _w15833_ ;
	wire _w15834_ ;
	wire _w15835_ ;
	wire _w15836_ ;
	wire _w15837_ ;
	wire _w15838_ ;
	wire _w15839_ ;
	wire _w15840_ ;
	wire _w15841_ ;
	wire _w15842_ ;
	wire _w15843_ ;
	wire _w15844_ ;
	wire _w15845_ ;
	wire _w15846_ ;
	wire _w15847_ ;
	wire _w15848_ ;
	wire _w15849_ ;
	wire _w15850_ ;
	wire _w15851_ ;
	wire _w15852_ ;
	wire _w15853_ ;
	wire _w15854_ ;
	wire _w15855_ ;
	wire _w15856_ ;
	wire _w15857_ ;
	wire _w15858_ ;
	wire _w15859_ ;
	wire _w15860_ ;
	wire _w15861_ ;
	wire _w15862_ ;
	wire _w15863_ ;
	wire _w15864_ ;
	wire _w15865_ ;
	wire _w15866_ ;
	wire _w15867_ ;
	wire _w15868_ ;
	wire _w15869_ ;
	wire _w15870_ ;
	wire _w15871_ ;
	wire _w15872_ ;
	wire _w15873_ ;
	wire _w15874_ ;
	wire _w15875_ ;
	wire _w15876_ ;
	wire _w15877_ ;
	wire _w15878_ ;
	wire _w15879_ ;
	wire _w15880_ ;
	wire _w15881_ ;
	wire _w15882_ ;
	wire _w15883_ ;
	wire _w15884_ ;
	wire _w15885_ ;
	wire _w15886_ ;
	wire _w15887_ ;
	wire _w15888_ ;
	wire _w15889_ ;
	wire _w15890_ ;
	wire _w15891_ ;
	wire _w15892_ ;
	wire _w15893_ ;
	wire _w15894_ ;
	wire _w15895_ ;
	wire _w15896_ ;
	wire _w15897_ ;
	wire _w15898_ ;
	wire _w15899_ ;
	wire _w15900_ ;
	wire _w15901_ ;
	wire _w15902_ ;
	wire _w15903_ ;
	wire _w15904_ ;
	wire _w15905_ ;
	wire _w15906_ ;
	wire _w15907_ ;
	wire _w15908_ ;
	wire _w15909_ ;
	wire _w15910_ ;
	wire _w15911_ ;
	wire _w15912_ ;
	wire _w15913_ ;
	wire _w15914_ ;
	wire _w15915_ ;
	wire _w15916_ ;
	wire _w15917_ ;
	wire _w15918_ ;
	wire _w15919_ ;
	wire _w15920_ ;
	wire _w15921_ ;
	wire _w15922_ ;
	wire _w15923_ ;
	wire _w15924_ ;
	wire _w15925_ ;
	wire _w15926_ ;
	wire _w15927_ ;
	wire _w15928_ ;
	wire _w15929_ ;
	wire _w15930_ ;
	wire _w15931_ ;
	wire _w15932_ ;
	wire _w15933_ ;
	wire _w15934_ ;
	wire _w15935_ ;
	wire _w15936_ ;
	wire _w15937_ ;
	wire _w15938_ ;
	wire _w15939_ ;
	wire _w15940_ ;
	wire _w15941_ ;
	wire _w15942_ ;
	wire _w15943_ ;
	wire _w15944_ ;
	wire _w15945_ ;
	wire _w15946_ ;
	wire _w15947_ ;
	wire _w15948_ ;
	wire _w15949_ ;
	wire _w15950_ ;
	wire _w15951_ ;
	wire _w15952_ ;
	wire _w15953_ ;
	wire _w15954_ ;
	wire _w15955_ ;
	wire _w15956_ ;
	wire _w15957_ ;
	wire _w15958_ ;
	wire _w15959_ ;
	wire _w15960_ ;
	wire _w15961_ ;
	wire _w15962_ ;
	wire _w15963_ ;
	wire _w15964_ ;
	wire _w15965_ ;
	wire _w15966_ ;
	wire _w15967_ ;
	wire _w15968_ ;
	wire _w15969_ ;
	wire _w15970_ ;
	wire _w15971_ ;
	wire _w15972_ ;
	wire _w15973_ ;
	wire _w15974_ ;
	wire _w15975_ ;
	wire _w15976_ ;
	wire _w15977_ ;
	wire _w15978_ ;
	wire _w15979_ ;
	wire _w15980_ ;
	wire _w15981_ ;
	wire _w15982_ ;
	wire _w15983_ ;
	wire _w15984_ ;
	wire _w15985_ ;
	wire _w15986_ ;
	wire _w15987_ ;
	wire _w15988_ ;
	wire _w15989_ ;
	wire _w15990_ ;
	wire _w15991_ ;
	wire _w15992_ ;
	wire _w15993_ ;
	wire _w15994_ ;
	wire _w15995_ ;
	wire _w15996_ ;
	wire _w15997_ ;
	wire _w15998_ ;
	wire _w15999_ ;
	wire _w16000_ ;
	wire _w16001_ ;
	wire _w16002_ ;
	wire _w16003_ ;
	wire _w16004_ ;
	wire _w16005_ ;
	wire _w16006_ ;
	wire _w16007_ ;
	wire _w16008_ ;
	wire _w16009_ ;
	wire _w16010_ ;
	wire _w16011_ ;
	wire _w16012_ ;
	wire _w16013_ ;
	wire _w16014_ ;
	wire _w16015_ ;
	wire _w16016_ ;
	wire _w16017_ ;
	wire _w16018_ ;
	wire _w16019_ ;
	wire _w16020_ ;
	wire _w16021_ ;
	wire _w16022_ ;
	wire _w16023_ ;
	wire _w16024_ ;
	wire _w16025_ ;
	wire _w16026_ ;
	wire _w16027_ ;
	wire _w16028_ ;
	wire _w16029_ ;
	wire _w16030_ ;
	wire _w16031_ ;
	wire _w16032_ ;
	wire _w16033_ ;
	wire _w16034_ ;
	wire _w16035_ ;
	wire _w16036_ ;
	wire _w16037_ ;
	wire _w16038_ ;
	wire _w16039_ ;
	wire _w16040_ ;
	wire _w16041_ ;
	wire _w16042_ ;
	wire _w16043_ ;
	wire _w16044_ ;
	wire _w16045_ ;
	wire _w16046_ ;
	wire _w16047_ ;
	wire _w16048_ ;
	wire _w16049_ ;
	wire _w16050_ ;
	wire _w16051_ ;
	wire _w16052_ ;
	wire _w16053_ ;
	wire _w16054_ ;
	wire _w16055_ ;
	wire _w16056_ ;
	wire _w16057_ ;
	wire _w16058_ ;
	wire _w16059_ ;
	wire _w16060_ ;
	wire _w16061_ ;
	wire _w16062_ ;
	wire _w16063_ ;
	wire _w16064_ ;
	wire _w16065_ ;
	wire _w16066_ ;
	wire _w16067_ ;
	wire _w16068_ ;
	wire _w16069_ ;
	wire _w16070_ ;
	wire _w16071_ ;
	wire _w16072_ ;
	wire _w16073_ ;
	wire _w16074_ ;
	wire _w16075_ ;
	wire _w16076_ ;
	wire _w16077_ ;
	wire _w16078_ ;
	wire _w16079_ ;
	wire _w16080_ ;
	wire _w16081_ ;
	wire _w16082_ ;
	wire _w16083_ ;
	wire _w16084_ ;
	wire _w16085_ ;
	wire _w16086_ ;
	wire _w16087_ ;
	wire _w16088_ ;
	wire _w16089_ ;
	wire _w16090_ ;
	wire _w16091_ ;
	wire _w16092_ ;
	wire _w16093_ ;
	wire _w16094_ ;
	wire _w16095_ ;
	wire _w16096_ ;
	wire _w16097_ ;
	wire _w16098_ ;
	wire _w16099_ ;
	wire _w16100_ ;
	wire _w16101_ ;
	wire _w16102_ ;
	wire _w16103_ ;
	wire _w16104_ ;
	wire _w16105_ ;
	wire _w16106_ ;
	wire _w16107_ ;
	wire _w16108_ ;
	wire _w16109_ ;
	wire _w16110_ ;
	wire _w16111_ ;
	wire _w16112_ ;
	wire _w16113_ ;
	wire _w16114_ ;
	wire _w16115_ ;
	wire _w16116_ ;
	wire _w16117_ ;
	wire _w16118_ ;
	wire _w16119_ ;
	wire _w16120_ ;
	wire _w16121_ ;
	wire _w16122_ ;
	wire _w16123_ ;
	wire _w16124_ ;
	wire _w16125_ ;
	wire _w16126_ ;
	wire _w16127_ ;
	wire _w16128_ ;
	wire _w16129_ ;
	wire _w16130_ ;
	wire _w16131_ ;
	wire _w16132_ ;
	wire _w16133_ ;
	wire _w16134_ ;
	wire _w16135_ ;
	wire _w16136_ ;
	wire _w16137_ ;
	wire _w16138_ ;
	wire _w16139_ ;
	wire _w16140_ ;
	wire _w16141_ ;
	wire _w16142_ ;
	wire _w16143_ ;
	wire _w16144_ ;
	wire _w16145_ ;
	wire _w16146_ ;
	wire _w16147_ ;
	wire _w16148_ ;
	wire _w16149_ ;
	wire _w16150_ ;
	wire _w16151_ ;
	wire _w16152_ ;
	wire _w16153_ ;
	wire _w16154_ ;
	wire _w16155_ ;
	wire _w16156_ ;
	wire _w16157_ ;
	wire _w16158_ ;
	wire _w16159_ ;
	wire _w16160_ ;
	wire _w16161_ ;
	wire _w16162_ ;
	wire _w16163_ ;
	wire _w16164_ ;
	wire _w16165_ ;
	wire _w16166_ ;
	wire _w16167_ ;
	wire _w16168_ ;
	wire _w16169_ ;
	wire _w16170_ ;
	wire _w16171_ ;
	wire _w16172_ ;
	wire _w16173_ ;
	wire _w16174_ ;
	wire _w16175_ ;
	wire _w16176_ ;
	wire _w16177_ ;
	wire _w16178_ ;
	wire _w16179_ ;
	wire _w16180_ ;
	wire _w16181_ ;
	wire _w16182_ ;
	wire _w16183_ ;
	wire _w16184_ ;
	wire _w16185_ ;
	wire _w16186_ ;
	wire _w16187_ ;
	wire _w16188_ ;
	wire _w16189_ ;
	wire _w16190_ ;
	wire _w16191_ ;
	wire _w16192_ ;
	wire _w16193_ ;
	wire _w16194_ ;
	wire _w16195_ ;
	wire _w16196_ ;
	wire _w16197_ ;
	wire _w16198_ ;
	wire _w16199_ ;
	wire _w16200_ ;
	wire _w16201_ ;
	wire _w16202_ ;
	wire _w16203_ ;
	wire _w16204_ ;
	wire _w16205_ ;
	wire _w16206_ ;
	wire _w16207_ ;
	wire _w16208_ ;
	wire _w16209_ ;
	wire _w16210_ ;
	wire _w16211_ ;
	wire _w16212_ ;
	wire _w16213_ ;
	wire _w16214_ ;
	wire _w16215_ ;
	wire _w16216_ ;
	wire _w16217_ ;
	wire _w16218_ ;
	wire _w16219_ ;
	wire _w16220_ ;
	wire _w16221_ ;
	wire _w16222_ ;
	wire _w16223_ ;
	wire _w16224_ ;
	wire _w16225_ ;
	wire _w16226_ ;
	wire _w16227_ ;
	wire _w16228_ ;
	wire _w16229_ ;
	wire _w16230_ ;
	wire _w16231_ ;
	wire _w16232_ ;
	wire _w16233_ ;
	wire _w16234_ ;
	wire _w16235_ ;
	wire _w16236_ ;
	wire _w16237_ ;
	wire _w16238_ ;
	wire _w16239_ ;
	wire _w16240_ ;
	wire _w16241_ ;
	wire _w16242_ ;
	wire _w16243_ ;
	wire _w16244_ ;
	wire _w16245_ ;
	wire _w16246_ ;
	wire _w16247_ ;
	wire _w16248_ ;
	wire _w16249_ ;
	wire _w16250_ ;
	wire _w16251_ ;
	wire _w16252_ ;
	wire _w16253_ ;
	wire _w16254_ ;
	wire _w16255_ ;
	wire _w16256_ ;
	wire _w16257_ ;
	wire _w16258_ ;
	wire _w16259_ ;
	wire _w16260_ ;
	wire _w16261_ ;
	wire _w16262_ ;
	wire _w16263_ ;
	wire _w16264_ ;
	wire _w16265_ ;
	wire _w16266_ ;
	wire _w16267_ ;
	wire _w16268_ ;
	wire _w16269_ ;
	wire _w16270_ ;
	wire _w16271_ ;
	wire _w16272_ ;
	wire _w16273_ ;
	wire _w16274_ ;
	wire _w16275_ ;
	wire _w16276_ ;
	wire _w16277_ ;
	wire _w16278_ ;
	wire _w16279_ ;
	wire _w16280_ ;
	wire _w16281_ ;
	wire _w16282_ ;
	wire _w16283_ ;
	wire _w16284_ ;
	wire _w16285_ ;
	wire _w16286_ ;
	wire _w16287_ ;
	wire _w16288_ ;
	wire _w16289_ ;
	wire _w16290_ ;
	wire _w16291_ ;
	wire _w16292_ ;
	wire _w16293_ ;
	wire _w16294_ ;
	wire _w16295_ ;
	wire _w16296_ ;
	wire _w16297_ ;
	wire _w16298_ ;
	wire _w16299_ ;
	wire _w16300_ ;
	wire _w16301_ ;
	wire _w16302_ ;
	wire _w16303_ ;
	wire _w16304_ ;
	wire _w16305_ ;
	wire _w16306_ ;
	wire _w16307_ ;
	wire _w16308_ ;
	wire _w16309_ ;
	wire _w16310_ ;
	wire _w16311_ ;
	wire _w16312_ ;
	wire _w16313_ ;
	wire _w16314_ ;
	wire _w16315_ ;
	wire _w16316_ ;
	wire _w16317_ ;
	wire _w16318_ ;
	wire _w16319_ ;
	wire _w16320_ ;
	wire _w16321_ ;
	wire _w16322_ ;
	wire _w16323_ ;
	wire _w16324_ ;
	wire _w16325_ ;
	wire _w16326_ ;
	wire _w16327_ ;
	wire _w16328_ ;
	wire _w16329_ ;
	wire _w16330_ ;
	wire _w16331_ ;
	wire _w16332_ ;
	wire _w16333_ ;
	wire _w16334_ ;
	wire _w16335_ ;
	wire _w16336_ ;
	wire _w16337_ ;
	wire _w16338_ ;
	wire _w16339_ ;
	wire _w16340_ ;
	wire _w16341_ ;
	wire _w16342_ ;
	wire _w16343_ ;
	wire _w16344_ ;
	wire _w16345_ ;
	wire _w16346_ ;
	wire _w16347_ ;
	wire _w16348_ ;
	wire _w16349_ ;
	wire _w16350_ ;
	wire _w16351_ ;
	wire _w16352_ ;
	wire _w16353_ ;
	wire _w16354_ ;
	wire _w16355_ ;
	wire _w16356_ ;
	wire _w16357_ ;
	wire _w16358_ ;
	wire _w16359_ ;
	wire _w16360_ ;
	wire _w16361_ ;
	wire _w16362_ ;
	wire _w16363_ ;
	wire _w16364_ ;
	wire _w16365_ ;
	wire _w16366_ ;
	wire _w16367_ ;
	wire _w16368_ ;
	wire _w16369_ ;
	wire _w16370_ ;
	wire _w16371_ ;
	wire _w16372_ ;
	wire _w16373_ ;
	wire _w16374_ ;
	wire _w16375_ ;
	wire _w16376_ ;
	wire _w16377_ ;
	wire _w16378_ ;
	wire _w16379_ ;
	wire _w16380_ ;
	wire _w16381_ ;
	wire _w16382_ ;
	wire _w16383_ ;
	wire _w16384_ ;
	wire _w16385_ ;
	wire _w16386_ ;
	wire _w16387_ ;
	wire _w16388_ ;
	wire _w16389_ ;
	wire _w16390_ ;
	wire _w16391_ ;
	wire _w16392_ ;
	wire _w16393_ ;
	wire _w16394_ ;
	wire _w16395_ ;
	wire _w16396_ ;
	wire _w16397_ ;
	wire _w16398_ ;
	wire _w16399_ ;
	wire _w16400_ ;
	wire _w16401_ ;
	wire _w16402_ ;
	wire _w16403_ ;
	wire _w16404_ ;
	wire _w16405_ ;
	wire _w16406_ ;
	wire _w16407_ ;
	wire _w16408_ ;
	wire _w16409_ ;
	wire _w16410_ ;
	wire _w16411_ ;
	wire _w16412_ ;
	wire _w16413_ ;
	wire _w16414_ ;
	wire _w16415_ ;
	wire _w16416_ ;
	wire _w16417_ ;
	wire _w16418_ ;
	wire _w16419_ ;
	wire _w16420_ ;
	wire _w16421_ ;
	wire _w16422_ ;
	wire _w16423_ ;
	wire _w16424_ ;
	wire _w16425_ ;
	wire _w16426_ ;
	wire _w16427_ ;
	wire _w16428_ ;
	wire _w16429_ ;
	wire _w16430_ ;
	wire _w16431_ ;
	wire _w16432_ ;
	wire _w16433_ ;
	wire _w16434_ ;
	wire _w16435_ ;
	wire _w16436_ ;
	wire _w16437_ ;
	wire _w16438_ ;
	wire _w16439_ ;
	wire _w16440_ ;
	wire _w16441_ ;
	wire _w16442_ ;
	wire _w16443_ ;
	wire _w16444_ ;
	wire _w16445_ ;
	wire _w16446_ ;
	wire _w16447_ ;
	wire _w16448_ ;
	wire _w16449_ ;
	wire _w16450_ ;
	wire _w16451_ ;
	wire _w16452_ ;
	wire _w16453_ ;
	wire _w16454_ ;
	wire _w16455_ ;
	wire _w16456_ ;
	wire _w16457_ ;
	wire _w16458_ ;
	wire _w16459_ ;
	wire _w16460_ ;
	wire _w16461_ ;
	wire _w16462_ ;
	wire _w16463_ ;
	wire _w16464_ ;
	wire _w16465_ ;
	wire _w16466_ ;
	wire _w16467_ ;
	wire _w16468_ ;
	wire _w16469_ ;
	wire _w16470_ ;
	wire _w16471_ ;
	wire _w16472_ ;
	wire _w16473_ ;
	wire _w16474_ ;
	wire _w16475_ ;
	wire _w16476_ ;
	wire _w16477_ ;
	wire _w16478_ ;
	wire _w16479_ ;
	wire _w16480_ ;
	wire _w16481_ ;
	wire _w16482_ ;
	wire _w16483_ ;
	wire _w16484_ ;
	wire _w16485_ ;
	wire _w16486_ ;
	wire _w16487_ ;
	wire _w16488_ ;
	wire _w16489_ ;
	wire _w16490_ ;
	wire _w16491_ ;
	wire _w16492_ ;
	wire _w16493_ ;
	wire _w16494_ ;
	wire _w16495_ ;
	wire _w16496_ ;
	wire _w16497_ ;
	wire _w16498_ ;
	wire _w16499_ ;
	wire _w16500_ ;
	wire _w16501_ ;
	wire _w16502_ ;
	wire _w16503_ ;
	wire _w16504_ ;
	wire _w16505_ ;
	wire _w16506_ ;
	wire _w16507_ ;
	wire _w16508_ ;
	wire _w16509_ ;
	wire _w16510_ ;
	wire _w16511_ ;
	wire _w16512_ ;
	wire _w16513_ ;
	wire _w16514_ ;
	wire _w16515_ ;
	wire _w16516_ ;
	wire _w16517_ ;
	wire _w16518_ ;
	wire _w16519_ ;
	wire _w16520_ ;
	wire _w16521_ ;
	wire _w16522_ ;
	wire _w16523_ ;
	wire _w16524_ ;
	wire _w16525_ ;
	wire _w16526_ ;
	wire _w16527_ ;
	wire _w16528_ ;
	wire _w16529_ ;
	wire _w16530_ ;
	wire _w16531_ ;
	wire _w16532_ ;
	wire _w16533_ ;
	wire _w16534_ ;
	wire _w16535_ ;
	wire _w16536_ ;
	wire _w16537_ ;
	wire _w16538_ ;
	wire _w16539_ ;
	wire _w16540_ ;
	wire _w16541_ ;
	wire _w16542_ ;
	wire _w16543_ ;
	wire _w16544_ ;
	wire _w16545_ ;
	wire _w16546_ ;
	wire _w16547_ ;
	wire _w16548_ ;
	wire _w16549_ ;
	wire _w16550_ ;
	wire _w16551_ ;
	wire _w16552_ ;
	wire _w16553_ ;
	wire _w16554_ ;
	wire _w16555_ ;
	wire _w16556_ ;
	wire _w16557_ ;
	wire _w16558_ ;
	wire _w16559_ ;
	wire _w16560_ ;
	wire _w16561_ ;
	wire _w16562_ ;
	wire _w16563_ ;
	wire _w16564_ ;
	wire _w16565_ ;
	wire _w16566_ ;
	wire _w16567_ ;
	wire _w16568_ ;
	wire _w16569_ ;
	wire _w16570_ ;
	wire _w16571_ ;
	wire _w16572_ ;
	wire _w16573_ ;
	wire _w16574_ ;
	wire _w16575_ ;
	wire _w16576_ ;
	wire _w16577_ ;
	wire _w16578_ ;
	wire _w16579_ ;
	wire _w16580_ ;
	wire _w16581_ ;
	wire _w16582_ ;
	wire _w16583_ ;
	wire _w16584_ ;
	wire _w16585_ ;
	wire _w16586_ ;
	wire _w16587_ ;
	wire _w16588_ ;
	wire _w16589_ ;
	wire _w16590_ ;
	wire _w16591_ ;
	wire _w16592_ ;
	wire _w16593_ ;
	wire _w16594_ ;
	wire _w16595_ ;
	wire _w16596_ ;
	wire _w16597_ ;
	wire _w16598_ ;
	wire _w16599_ ;
	wire _w16600_ ;
	wire _w16601_ ;
	wire _w16602_ ;
	wire _w16603_ ;
	wire _w16604_ ;
	wire _w16605_ ;
	wire _w16606_ ;
	wire _w16607_ ;
	wire _w16608_ ;
	wire _w16609_ ;
	wire _w16610_ ;
	wire _w16611_ ;
	wire _w16612_ ;
	wire _w16613_ ;
	wire _w16614_ ;
	wire _w16615_ ;
	wire _w16616_ ;
	wire _w16617_ ;
	wire _w16618_ ;
	wire _w16619_ ;
	wire _w16620_ ;
	wire _w16621_ ;
	wire _w16622_ ;
	wire _w16623_ ;
	wire _w16624_ ;
	wire _w16625_ ;
	wire _w16626_ ;
	wire _w16627_ ;
	wire _w16628_ ;
	wire _w16629_ ;
	wire _w16630_ ;
	wire _w16631_ ;
	wire _w16632_ ;
	wire _w16633_ ;
	wire _w16634_ ;
	wire _w16635_ ;
	wire _w16636_ ;
	wire _w16637_ ;
	wire _w16638_ ;
	wire _w16639_ ;
	wire _w16640_ ;
	wire _w16641_ ;
	wire _w16642_ ;
	wire _w16643_ ;
	wire _w16644_ ;
	wire _w16645_ ;
	wire _w16646_ ;
	wire _w16647_ ;
	wire _w16648_ ;
	wire _w16649_ ;
	wire _w16650_ ;
	wire _w16651_ ;
	wire _w16652_ ;
	wire _w16653_ ;
	wire _w16654_ ;
	wire _w16655_ ;
	wire _w16656_ ;
	wire _w16657_ ;
	wire _w16658_ ;
	wire _w16659_ ;
	wire _w16660_ ;
	wire _w16661_ ;
	wire _w16662_ ;
	wire _w16663_ ;
	wire _w16664_ ;
	wire _w16665_ ;
	wire _w16666_ ;
	wire _w16667_ ;
	wire _w16668_ ;
	wire _w16669_ ;
	wire _w16670_ ;
	wire _w16671_ ;
	wire _w16672_ ;
	wire _w16673_ ;
	wire _w16674_ ;
	wire _w16675_ ;
	wire _w16676_ ;
	wire _w16677_ ;
	wire _w16678_ ;
	wire _w16679_ ;
	wire _w16680_ ;
	wire _w16681_ ;
	wire _w16682_ ;
	wire _w16683_ ;
	wire _w16684_ ;
	wire _w16685_ ;
	wire _w16686_ ;
	wire _w16687_ ;
	wire _w16688_ ;
	wire _w16689_ ;
	wire _w16690_ ;
	wire _w16691_ ;
	wire _w16692_ ;
	wire _w16693_ ;
	wire _w16694_ ;
	wire _w16695_ ;
	wire _w16696_ ;
	wire _w16697_ ;
	wire _w16698_ ;
	wire _w16699_ ;
	wire _w16700_ ;
	wire _w16701_ ;
	wire _w16702_ ;
	wire _w16703_ ;
	wire _w16704_ ;
	wire _w16705_ ;
	wire _w16706_ ;
	wire _w16707_ ;
	wire _w16708_ ;
	wire _w16709_ ;
	wire _w16710_ ;
	wire _w16711_ ;
	wire _w16712_ ;
	wire _w16713_ ;
	wire _w16714_ ;
	wire _w16715_ ;
	wire _w16716_ ;
	wire _w16717_ ;
	wire _w16718_ ;
	wire _w16719_ ;
	wire _w16720_ ;
	wire _w16721_ ;
	wire _w16722_ ;
	wire _w16723_ ;
	wire _w16724_ ;
	wire _w16725_ ;
	wire _w16726_ ;
	wire _w16727_ ;
	wire _w16728_ ;
	wire _w16729_ ;
	wire _w16730_ ;
	wire _w16731_ ;
	wire _w16732_ ;
	wire _w16733_ ;
	wire _w16734_ ;
	wire _w16735_ ;
	wire _w16736_ ;
	wire _w16737_ ;
	wire _w16738_ ;
	wire _w16739_ ;
	wire _w16740_ ;
	wire _w16741_ ;
	wire _w16742_ ;
	wire _w16743_ ;
	wire _w16744_ ;
	wire _w16745_ ;
	wire _w16746_ ;
	wire _w16747_ ;
	wire _w16748_ ;
	wire _w16749_ ;
	wire _w16750_ ;
	wire _w16751_ ;
	wire _w16752_ ;
	wire _w16753_ ;
	wire _w16754_ ;
	wire _w16755_ ;
	wire _w16756_ ;
	wire _w16757_ ;
	wire _w16758_ ;
	wire _w16759_ ;
	wire _w16760_ ;
	wire _w16761_ ;
	wire _w16762_ ;
	wire _w16763_ ;
	wire _w16764_ ;
	wire _w16765_ ;
	wire _w16766_ ;
	wire _w16767_ ;
	wire _w16768_ ;
	wire _w16769_ ;
	wire _w16770_ ;
	wire _w16771_ ;
	wire _w16772_ ;
	wire _w16773_ ;
	wire _w16774_ ;
	wire _w16775_ ;
	wire _w16776_ ;
	wire _w16777_ ;
	wire _w16778_ ;
	wire _w16779_ ;
	wire _w16780_ ;
	wire _w16781_ ;
	wire _w16782_ ;
	wire _w16783_ ;
	wire _w16784_ ;
	wire _w16785_ ;
	wire _w16786_ ;
	wire _w16787_ ;
	wire _w16788_ ;
	wire _w16789_ ;
	wire _w16790_ ;
	wire _w16791_ ;
	wire _w16792_ ;
	wire _w16793_ ;
	wire _w16794_ ;
	wire _w16795_ ;
	wire _w16796_ ;
	wire _w16797_ ;
	wire _w16798_ ;
	wire _w16799_ ;
	wire _w16800_ ;
	wire _w16801_ ;
	wire _w16802_ ;
	wire _w16803_ ;
	wire _w16804_ ;
	wire _w16805_ ;
	wire _w16806_ ;
	wire _w16807_ ;
	wire _w16808_ ;
	wire _w16809_ ;
	wire _w16810_ ;
	wire _w16811_ ;
	wire _w16812_ ;
	wire _w16813_ ;
	wire _w16814_ ;
	wire _w16815_ ;
	wire _w16816_ ;
	wire _w16817_ ;
	wire _w16818_ ;
	wire _w16819_ ;
	wire _w16820_ ;
	wire _w16821_ ;
	wire _w16822_ ;
	wire _w16823_ ;
	wire _w16824_ ;
	wire _w16825_ ;
	wire _w16826_ ;
	wire _w16827_ ;
	wire _w16828_ ;
	wire _w16829_ ;
	wire _w16830_ ;
	wire _w16831_ ;
	wire _w16832_ ;
	wire _w16833_ ;
	wire _w16834_ ;
	wire _w16835_ ;
	wire _w16836_ ;
	wire _w16837_ ;
	wire _w16838_ ;
	wire _w16839_ ;
	wire _w16840_ ;
	wire _w16841_ ;
	wire _w16842_ ;
	wire _w16843_ ;
	wire _w16844_ ;
	wire _w16845_ ;
	wire _w16846_ ;
	wire _w16847_ ;
	wire _w16848_ ;
	wire _w16849_ ;
	wire _w16850_ ;
	wire _w16851_ ;
	wire _w16852_ ;
	wire _w16853_ ;
	wire _w16854_ ;
	wire _w16855_ ;
	wire _w16856_ ;
	wire _w16857_ ;
	wire _w16858_ ;
	wire _w16859_ ;
	wire _w16860_ ;
	wire _w16861_ ;
	wire _w16862_ ;
	wire _w16863_ ;
	wire _w16864_ ;
	wire _w16865_ ;
	wire _w16866_ ;
	wire _w16867_ ;
	wire _w16868_ ;
	wire _w16869_ ;
	wire _w16870_ ;
	wire _w16871_ ;
	wire _w16872_ ;
	wire _w16873_ ;
	wire _w16874_ ;
	wire _w16875_ ;
	wire _w16876_ ;
	wire _w16877_ ;
	wire _w16878_ ;
	wire _w16879_ ;
	wire _w16880_ ;
	wire _w16881_ ;
	wire _w16882_ ;
	wire _w16883_ ;
	wire _w16884_ ;
	wire _w16885_ ;
	wire _w16886_ ;
	wire _w16887_ ;
	wire _w16888_ ;
	wire _w16889_ ;
	wire _w16890_ ;
	wire _w16891_ ;
	wire _w16892_ ;
	wire _w16893_ ;
	wire _w16894_ ;
	wire _w16895_ ;
	wire _w16896_ ;
	wire _w16897_ ;
	wire _w16898_ ;
	wire _w16899_ ;
	wire _w16900_ ;
	wire _w16901_ ;
	wire _w16902_ ;
	wire _w16903_ ;
	wire _w16904_ ;
	wire _w16905_ ;
	wire _w16906_ ;
	wire _w16907_ ;
	wire _w16908_ ;
	wire _w16909_ ;
	wire _w16910_ ;
	wire _w16911_ ;
	wire _w16912_ ;
	wire _w16913_ ;
	wire _w16914_ ;
	wire _w16915_ ;
	wire _w16916_ ;
	wire _w16917_ ;
	wire _w16918_ ;
	wire _w16919_ ;
	wire _w16920_ ;
	wire _w16921_ ;
	wire _w16922_ ;
	wire _w16923_ ;
	wire _w16924_ ;
	wire _w16925_ ;
	wire _w16926_ ;
	wire _w16927_ ;
	wire _w16928_ ;
	wire _w16929_ ;
	wire _w16930_ ;
	wire _w16931_ ;
	wire _w16932_ ;
	wire _w16933_ ;
	wire _w16934_ ;
	wire _w16935_ ;
	wire _w16936_ ;
	wire _w16937_ ;
	wire _w16938_ ;
	wire _w16939_ ;
	wire _w16940_ ;
	wire _w16941_ ;
	wire _w16942_ ;
	wire _w16943_ ;
	wire _w16944_ ;
	wire _w16945_ ;
	wire _w16946_ ;
	wire _w16947_ ;
	wire _w16948_ ;
	wire _w16949_ ;
	wire _w16950_ ;
	wire _w16951_ ;
	wire _w16952_ ;
	wire _w16953_ ;
	wire _w16954_ ;
	wire _w16955_ ;
	wire _w16956_ ;
	wire _w16957_ ;
	wire _w16958_ ;
	wire _w16959_ ;
	wire _w16960_ ;
	wire _w16961_ ;
	wire _w16962_ ;
	wire _w16963_ ;
	wire _w16964_ ;
	wire _w16965_ ;
	wire _w16966_ ;
	wire _w16967_ ;
	wire _w16968_ ;
	wire _w16969_ ;
	wire _w16970_ ;
	wire _w16971_ ;
	wire _w16972_ ;
	wire _w16973_ ;
	wire _w16974_ ;
	wire _w16975_ ;
	wire _w16976_ ;
	wire _w16977_ ;
	wire _w16978_ ;
	wire _w16979_ ;
	wire _w16980_ ;
	wire _w16981_ ;
	wire _w16982_ ;
	wire _w16983_ ;
	wire _w16984_ ;
	wire _w16985_ ;
	wire _w16986_ ;
	wire _w16987_ ;
	wire _w16988_ ;
	wire _w16989_ ;
	wire _w16990_ ;
	wire _w16991_ ;
	wire _w16992_ ;
	wire _w16993_ ;
	wire _w16994_ ;
	wire _w16995_ ;
	wire _w16996_ ;
	wire _w16997_ ;
	wire _w16998_ ;
	wire _w16999_ ;
	wire _w17000_ ;
	wire _w17001_ ;
	wire _w17002_ ;
	wire _w17003_ ;
	wire _w17004_ ;
	wire _w17005_ ;
	wire _w17006_ ;
	wire _w17007_ ;
	wire _w17008_ ;
	wire _w17009_ ;
	wire _w17010_ ;
	wire _w17011_ ;
	wire _w17012_ ;
	wire _w17013_ ;
	wire _w17014_ ;
	wire _w17015_ ;
	wire _w17016_ ;
	wire _w17017_ ;
	wire _w17018_ ;
	wire _w17019_ ;
	wire _w17020_ ;
	wire _w17021_ ;
	wire _w17022_ ;
	wire _w17023_ ;
	wire _w17024_ ;
	wire _w17025_ ;
	wire _w17026_ ;
	wire _w17027_ ;
	wire _w17028_ ;
	wire _w17029_ ;
	wire _w17030_ ;
	wire _w17031_ ;
	wire _w17032_ ;
	wire _w17033_ ;
	wire _w17034_ ;
	wire _w17035_ ;
	wire _w17036_ ;
	wire _w17037_ ;
	wire _w17038_ ;
	wire _w17039_ ;
	wire _w17040_ ;
	wire _w17041_ ;
	wire _w17042_ ;
	wire _w17043_ ;
	wire _w17044_ ;
	wire _w17045_ ;
	wire _w17046_ ;
	wire _w17047_ ;
	wire _w17048_ ;
	wire _w17049_ ;
	wire _w17050_ ;
	wire _w17051_ ;
	wire _w17052_ ;
	wire _w17053_ ;
	wire _w17054_ ;
	wire _w17055_ ;
	wire _w17056_ ;
	wire _w17057_ ;
	wire _w17058_ ;
	wire _w17059_ ;
	wire _w17060_ ;
	wire _w17061_ ;
	wire _w17062_ ;
	wire _w17063_ ;
	wire _w17064_ ;
	wire _w17065_ ;
	wire _w17066_ ;
	wire _w17067_ ;
	wire _w17068_ ;
	wire _w17069_ ;
	wire _w17070_ ;
	wire _w17071_ ;
	wire _w17072_ ;
	wire _w17073_ ;
	wire _w17074_ ;
	wire _w17075_ ;
	wire _w17076_ ;
	wire _w17077_ ;
	wire _w17078_ ;
	wire _w17079_ ;
	wire _w17080_ ;
	wire _w17081_ ;
	wire _w17082_ ;
	wire _w17083_ ;
	wire _w17084_ ;
	wire _w17085_ ;
	wire _w17086_ ;
	wire _w17087_ ;
	wire _w17088_ ;
	wire _w17089_ ;
	wire _w17090_ ;
	wire _w17091_ ;
	wire _w17092_ ;
	wire _w17093_ ;
	wire _w17094_ ;
	wire _w17095_ ;
	wire _w17096_ ;
	wire _w17097_ ;
	wire _w17098_ ;
	wire _w17099_ ;
	wire _w17100_ ;
	wire _w17101_ ;
	wire _w17102_ ;
	wire _w17103_ ;
	wire _w17104_ ;
	wire _w17105_ ;
	wire _w17106_ ;
	wire _w17107_ ;
	wire _w17108_ ;
	wire _w17109_ ;
	wire _w17110_ ;
	wire _w17111_ ;
	wire _w17112_ ;
	wire _w17113_ ;
	wire _w17114_ ;
	wire _w17115_ ;
	wire _w17116_ ;
	wire _w17117_ ;
	wire _w17118_ ;
	wire _w17119_ ;
	wire _w17120_ ;
	wire _w17121_ ;
	wire _w17122_ ;
	wire _w17123_ ;
	wire _w17124_ ;
	wire _w17125_ ;
	wire _w17126_ ;
	wire _w17127_ ;
	wire _w17128_ ;
	wire _w17129_ ;
	wire _w17130_ ;
	wire _w17131_ ;
	wire _w17132_ ;
	wire _w17133_ ;
	wire _w17134_ ;
	wire _w17135_ ;
	wire _w17136_ ;
	wire _w17137_ ;
	wire _w17138_ ;
	wire _w17139_ ;
	wire _w17140_ ;
	wire _w17141_ ;
	wire _w17142_ ;
	wire _w17143_ ;
	wire _w17144_ ;
	wire _w17145_ ;
	wire _w17146_ ;
	wire _w17147_ ;
	wire _w17148_ ;
	wire _w17149_ ;
	wire _w17150_ ;
	wire _w17151_ ;
	wire _w17152_ ;
	wire _w17153_ ;
	wire _w17154_ ;
	wire _w17155_ ;
	wire _w17156_ ;
	wire _w17157_ ;
	wire _w17158_ ;
	wire _w17159_ ;
	wire _w17160_ ;
	wire _w17161_ ;
	wire _w17162_ ;
	wire _w17163_ ;
	wire _w17164_ ;
	wire _w17165_ ;
	wire _w17166_ ;
	wire _w17167_ ;
	wire _w17168_ ;
	wire _w17169_ ;
	wire _w17170_ ;
	wire _w17171_ ;
	wire _w17172_ ;
	wire _w17173_ ;
	wire _w17174_ ;
	wire _w17175_ ;
	wire _w17176_ ;
	wire _w17177_ ;
	wire _w17178_ ;
	wire _w17179_ ;
	wire _w17180_ ;
	wire _w17181_ ;
	wire _w17182_ ;
	wire _w17183_ ;
	wire _w17184_ ;
	wire _w17185_ ;
	wire _w17186_ ;
	wire _w17187_ ;
	wire _w17188_ ;
	wire _w17189_ ;
	wire _w17190_ ;
	wire _w17191_ ;
	wire _w17192_ ;
	wire _w17193_ ;
	wire _w17194_ ;
	wire _w17195_ ;
	wire _w17196_ ;
	wire _w17197_ ;
	wire _w17198_ ;
	wire _w17199_ ;
	wire _w17200_ ;
	wire _w17201_ ;
	wire _w17202_ ;
	wire _w17203_ ;
	wire _w17204_ ;
	wire _w17205_ ;
	wire _w17206_ ;
	wire _w17207_ ;
	wire _w17208_ ;
	wire _w17209_ ;
	wire _w17210_ ;
	wire _w17211_ ;
	wire _w17212_ ;
	wire _w17213_ ;
	wire _w17214_ ;
	wire _w17215_ ;
	wire _w17216_ ;
	wire _w17217_ ;
	wire _w17218_ ;
	wire _w17219_ ;
	wire _w17220_ ;
	wire _w17221_ ;
	wire _w17222_ ;
	wire _w17223_ ;
	wire _w17224_ ;
	wire _w17225_ ;
	wire _w17226_ ;
	wire _w17227_ ;
	wire _w17228_ ;
	wire _w17229_ ;
	wire _w17230_ ;
	wire _w17231_ ;
	wire _w17232_ ;
	wire _w17233_ ;
	wire _w17234_ ;
	wire _w17235_ ;
	wire _w17236_ ;
	wire _w17237_ ;
	wire _w17238_ ;
	wire _w17239_ ;
	wire _w17240_ ;
	wire _w17241_ ;
	wire _w17242_ ;
	wire _w17243_ ;
	wire _w17244_ ;
	wire _w17245_ ;
	wire _w17246_ ;
	wire _w17247_ ;
	wire _w17248_ ;
	wire _w17249_ ;
	wire _w17250_ ;
	wire _w17251_ ;
	wire _w17252_ ;
	wire _w17253_ ;
	wire _w17254_ ;
	wire _w17255_ ;
	wire _w17256_ ;
	wire _w17257_ ;
	wire _w17258_ ;
	wire _w17259_ ;
	wire _w17260_ ;
	wire _w17261_ ;
	wire _w17262_ ;
	wire _w17263_ ;
	wire _w17264_ ;
	wire _w17265_ ;
	wire _w17266_ ;
	wire _w17267_ ;
	wire _w17268_ ;
	wire _w17269_ ;
	wire _w17270_ ;
	wire _w17271_ ;
	wire _w17272_ ;
	wire _w17273_ ;
	wire _w17274_ ;
	wire _w17275_ ;
	wire _w17276_ ;
	wire _w17277_ ;
	wire _w17278_ ;
	wire _w17279_ ;
	wire _w17280_ ;
	wire _w17281_ ;
	wire _w17282_ ;
	wire _w17283_ ;
	wire _w17284_ ;
	wire _w17285_ ;
	wire _w17286_ ;
	wire _w17287_ ;
	wire _w17288_ ;
	wire _w17289_ ;
	wire _w17290_ ;
	wire _w17291_ ;
	wire _w17292_ ;
	wire _w17293_ ;
	wire _w17294_ ;
	wire _w17295_ ;
	wire _w17296_ ;
	wire _w17297_ ;
	wire _w17298_ ;
	wire _w17299_ ;
	wire _w17300_ ;
	wire _w17301_ ;
	wire _w17302_ ;
	wire _w17303_ ;
	wire _w17304_ ;
	wire _w17305_ ;
	wire _w17306_ ;
	wire _w17307_ ;
	wire _w17308_ ;
	wire _w17309_ ;
	wire _w17310_ ;
	wire _w17311_ ;
	wire _w17312_ ;
	wire _w17313_ ;
	wire _w17314_ ;
	wire _w17315_ ;
	wire _w17316_ ;
	wire _w17317_ ;
	wire _w17318_ ;
	wire _w17319_ ;
	wire _w17320_ ;
	wire _w17321_ ;
	wire _w17322_ ;
	wire _w17323_ ;
	wire _w17324_ ;
	wire _w17325_ ;
	wire _w17326_ ;
	wire _w17327_ ;
	wire _w17328_ ;
	wire _w17329_ ;
	wire _w17330_ ;
	wire _w17331_ ;
	wire _w17332_ ;
	wire _w17333_ ;
	wire _w17334_ ;
	wire _w17335_ ;
	wire _w17336_ ;
	wire _w17337_ ;
	wire _w17338_ ;
	wire _w17339_ ;
	wire _w17340_ ;
	wire _w17341_ ;
	wire _w17342_ ;
	wire _w17343_ ;
	wire _w17344_ ;
	wire _w17345_ ;
	wire _w17346_ ;
	wire _w17347_ ;
	wire _w17348_ ;
	wire _w17349_ ;
	wire _w17350_ ;
	wire _w17351_ ;
	wire _w17352_ ;
	wire _w17353_ ;
	wire _w17354_ ;
	wire _w17355_ ;
	wire _w17356_ ;
	wire _w17357_ ;
	wire _w17358_ ;
	wire _w17359_ ;
	wire _w17360_ ;
	wire _w17361_ ;
	wire _w17362_ ;
	wire _w17363_ ;
	wire _w17364_ ;
	wire _w17365_ ;
	wire _w17366_ ;
	wire _w17367_ ;
	wire _w17368_ ;
	wire _w17369_ ;
	wire _w17370_ ;
	wire _w17371_ ;
	wire _w17372_ ;
	wire _w17373_ ;
	wire _w17374_ ;
	wire _w17375_ ;
	wire _w17376_ ;
	wire _w17377_ ;
	wire _w17378_ ;
	wire _w17379_ ;
	wire _w17380_ ;
	wire _w17381_ ;
	wire _w17382_ ;
	wire _w17383_ ;
	wire _w17384_ ;
	wire _w17385_ ;
	wire _w17386_ ;
	wire _w17387_ ;
	wire _w17388_ ;
	wire _w17389_ ;
	wire _w17390_ ;
	wire _w17391_ ;
	wire _w17392_ ;
	wire _w17393_ ;
	wire _w17394_ ;
	wire _w17395_ ;
	wire _w17396_ ;
	wire _w17397_ ;
	wire _w17398_ ;
	wire _w17399_ ;
	wire _w17400_ ;
	wire _w17401_ ;
	wire _w17402_ ;
	wire _w17403_ ;
	wire _w17404_ ;
	wire _w17405_ ;
	wire _w17406_ ;
	wire _w17407_ ;
	wire _w17408_ ;
	wire _w17409_ ;
	wire _w17410_ ;
	wire _w17411_ ;
	wire _w17412_ ;
	wire _w17413_ ;
	wire _w17414_ ;
	wire _w17415_ ;
	wire _w17416_ ;
	wire _w17417_ ;
	wire _w17418_ ;
	wire _w17419_ ;
	wire _w17420_ ;
	wire _w17421_ ;
	wire _w17422_ ;
	wire _w17423_ ;
	wire _w17424_ ;
	wire _w17425_ ;
	wire _w17426_ ;
	wire _w17427_ ;
	wire _w17428_ ;
	wire _w17429_ ;
	wire _w17430_ ;
	wire _w17431_ ;
	wire _w17432_ ;
	wire _w17433_ ;
	wire _w17434_ ;
	wire _w17435_ ;
	wire _w17436_ ;
	wire _w17437_ ;
	wire _w17438_ ;
	wire _w17439_ ;
	wire _w17440_ ;
	wire _w17441_ ;
	wire _w17442_ ;
	wire _w17443_ ;
	wire _w17444_ ;
	wire _w17445_ ;
	wire _w17446_ ;
	wire _w17447_ ;
	wire _w17448_ ;
	wire _w17449_ ;
	wire _w17450_ ;
	wire _w17451_ ;
	wire _w17452_ ;
	wire _w17453_ ;
	wire _w17454_ ;
	wire _w17455_ ;
	wire _w17456_ ;
	wire _w17457_ ;
	wire _w17458_ ;
	wire _w17459_ ;
	wire _w17460_ ;
	wire _w17461_ ;
	wire _w17462_ ;
	wire _w17463_ ;
	wire _w17464_ ;
	wire _w17465_ ;
	wire _w17466_ ;
	wire _w17467_ ;
	wire _w17468_ ;
	wire _w17469_ ;
	wire _w17470_ ;
	wire _w17471_ ;
	wire _w17472_ ;
	wire _w17473_ ;
	wire _w17474_ ;
	wire _w17475_ ;
	wire _w17476_ ;
	wire _w17477_ ;
	wire _w17478_ ;
	wire _w17479_ ;
	wire _w17480_ ;
	wire _w17481_ ;
	wire _w17482_ ;
	wire _w17483_ ;
	wire _w17484_ ;
	wire _w17485_ ;
	wire _w17486_ ;
	wire _w17487_ ;
	wire _w17488_ ;
	wire _w17489_ ;
	wire _w17490_ ;
	wire _w17491_ ;
	wire _w17492_ ;
	wire _w17493_ ;
	wire _w17494_ ;
	wire _w17495_ ;
	wire _w17496_ ;
	wire _w17497_ ;
	wire _w17498_ ;
	wire _w17499_ ;
	wire _w17500_ ;
	wire _w17501_ ;
	wire _w17502_ ;
	wire _w17503_ ;
	wire _w17504_ ;
	wire _w17505_ ;
	wire _w17506_ ;
	wire _w17507_ ;
	wire _w17508_ ;
	wire _w17509_ ;
	wire _w17510_ ;
	wire _w17511_ ;
	wire _w17512_ ;
	wire _w17513_ ;
	wire _w17514_ ;
	wire _w17515_ ;
	wire _w17516_ ;
	wire _w17517_ ;
	wire _w17518_ ;
	wire _w17519_ ;
	wire _w17520_ ;
	wire _w17521_ ;
	wire _w17522_ ;
	wire _w17523_ ;
	wire _w17524_ ;
	wire _w17525_ ;
	wire _w17526_ ;
	wire _w17527_ ;
	wire _w17528_ ;
	wire _w17529_ ;
	wire _w17530_ ;
	wire _w17531_ ;
	wire _w17532_ ;
	wire _w17533_ ;
	wire _w17534_ ;
	wire _w17535_ ;
	wire _w17536_ ;
	wire _w17537_ ;
	wire _w17538_ ;
	wire _w17539_ ;
	wire _w17540_ ;
	wire _w17541_ ;
	wire _w17542_ ;
	wire _w17543_ ;
	wire _w17544_ ;
	wire _w17545_ ;
	wire _w17546_ ;
	wire _w17547_ ;
	wire _w17548_ ;
	wire _w17549_ ;
	wire _w17550_ ;
	wire _w17551_ ;
	wire _w17552_ ;
	wire _w17553_ ;
	wire _w17554_ ;
	wire _w17555_ ;
	wire _w17556_ ;
	wire _w17557_ ;
	wire _w17558_ ;
	wire _w17559_ ;
	wire _w17560_ ;
	wire _w17561_ ;
	wire _w17562_ ;
	wire _w17563_ ;
	wire _w17564_ ;
	wire _w17565_ ;
	wire _w17566_ ;
	wire _w17567_ ;
	wire _w17568_ ;
	wire _w17569_ ;
	wire _w17570_ ;
	wire _w17571_ ;
	wire _w17572_ ;
	wire _w17573_ ;
	wire _w17574_ ;
	wire _w17575_ ;
	wire _w17576_ ;
	wire _w17577_ ;
	wire _w17578_ ;
	wire _w17579_ ;
	wire _w17580_ ;
	wire _w17581_ ;
	wire _w17582_ ;
	wire _w17583_ ;
	wire _w17584_ ;
	wire _w17585_ ;
	wire _w17586_ ;
	wire _w17587_ ;
	wire _w17588_ ;
	wire _w17589_ ;
	wire _w17590_ ;
	wire _w17591_ ;
	wire _w17592_ ;
	wire _w17593_ ;
	wire _w17594_ ;
	wire _w17595_ ;
	wire _w17596_ ;
	wire _w17597_ ;
	wire _w17598_ ;
	wire _w17599_ ;
	wire _w17600_ ;
	wire _w17601_ ;
	wire _w17602_ ;
	wire _w17603_ ;
	wire _w17604_ ;
	wire _w17605_ ;
	wire _w17606_ ;
	wire _w17607_ ;
	wire _w17608_ ;
	wire _w17609_ ;
	wire _w17610_ ;
	wire _w17611_ ;
	wire _w17612_ ;
	wire _w17613_ ;
	wire _w17614_ ;
	wire _w17615_ ;
	wire _w17616_ ;
	wire _w17617_ ;
	wire _w17618_ ;
	wire _w17619_ ;
	wire _w17620_ ;
	wire _w17621_ ;
	wire _w17622_ ;
	wire _w17623_ ;
	wire _w17624_ ;
	wire _w17625_ ;
	wire _w17626_ ;
	wire _w17627_ ;
	wire _w17628_ ;
	wire _w17629_ ;
	wire _w17630_ ;
	wire _w17631_ ;
	wire _w17632_ ;
	wire _w17633_ ;
	wire _w17634_ ;
	wire _w17635_ ;
	wire _w17636_ ;
	wire _w17637_ ;
	wire _w17638_ ;
	wire _w17639_ ;
	wire _w17640_ ;
	wire _w17641_ ;
	wire _w17642_ ;
	wire _w17643_ ;
	wire _w17644_ ;
	wire _w17645_ ;
	wire _w17646_ ;
	wire _w17647_ ;
	wire _w17648_ ;
	wire _w17649_ ;
	wire _w17650_ ;
	wire _w17651_ ;
	wire _w17652_ ;
	wire _w17653_ ;
	wire _w17654_ ;
	wire _w17655_ ;
	wire _w17656_ ;
	wire _w17657_ ;
	wire _w17658_ ;
	wire _w17659_ ;
	wire _w17660_ ;
	wire _w17661_ ;
	wire _w17662_ ;
	wire _w17663_ ;
	wire _w17664_ ;
	wire _w17665_ ;
	wire _w17666_ ;
	wire _w17667_ ;
	wire _w17668_ ;
	wire _w17669_ ;
	wire _w17670_ ;
	wire _w17671_ ;
	wire _w17672_ ;
	wire _w17673_ ;
	wire _w17674_ ;
	wire _w17675_ ;
	wire _w17676_ ;
	wire _w17677_ ;
	wire _w17678_ ;
	wire _w17679_ ;
	wire _w17680_ ;
	wire _w17681_ ;
	wire _w17682_ ;
	wire _w17683_ ;
	wire _w17684_ ;
	wire _w17685_ ;
	wire _w17686_ ;
	wire _w17687_ ;
	wire _w17688_ ;
	wire _w17689_ ;
	wire _w17690_ ;
	wire _w17691_ ;
	wire _w17692_ ;
	wire _w17693_ ;
	wire _w17694_ ;
	wire _w17695_ ;
	wire _w17696_ ;
	wire _w17697_ ;
	wire _w17698_ ;
	wire _w17699_ ;
	wire _w17700_ ;
	wire _w17701_ ;
	wire _w17702_ ;
	wire _w17703_ ;
	wire _w17704_ ;
	wire _w17705_ ;
	wire _w17706_ ;
	wire _w17707_ ;
	wire _w17708_ ;
	wire _w17709_ ;
	wire _w17710_ ;
	wire _w17711_ ;
	wire _w17712_ ;
	wire _w17713_ ;
	wire _w17714_ ;
	wire _w17715_ ;
	wire _w17716_ ;
	wire _w17717_ ;
	wire _w17718_ ;
	wire _w17719_ ;
	wire _w17720_ ;
	wire _w17721_ ;
	wire _w17722_ ;
	wire _w17723_ ;
	wire _w17724_ ;
	wire _w17725_ ;
	wire _w17726_ ;
	wire _w17727_ ;
	wire _w17728_ ;
	wire _w17729_ ;
	wire _w17730_ ;
	wire _w17731_ ;
	wire _w17732_ ;
	wire _w17733_ ;
	wire _w17734_ ;
	wire _w17735_ ;
	wire _w17736_ ;
	wire _w17737_ ;
	wire _w17738_ ;
	wire _w17739_ ;
	wire _w17740_ ;
	wire _w17741_ ;
	wire _w17742_ ;
	wire _w17743_ ;
	wire _w17744_ ;
	wire _w17745_ ;
	wire _w17746_ ;
	wire _w17747_ ;
	wire _w17748_ ;
	wire _w17749_ ;
	wire _w17750_ ;
	wire _w17751_ ;
	wire _w17752_ ;
	wire _w17753_ ;
	wire _w17754_ ;
	wire _w17755_ ;
	wire _w17756_ ;
	wire _w17757_ ;
	wire _w17758_ ;
	wire _w17759_ ;
	wire _w17760_ ;
	wire _w17761_ ;
	wire _w17762_ ;
	wire _w17763_ ;
	wire _w17764_ ;
	wire _w17765_ ;
	wire _w17766_ ;
	wire _w17767_ ;
	wire _w17768_ ;
	wire _w17769_ ;
	wire _w17770_ ;
	wire _w17771_ ;
	wire _w17772_ ;
	wire _w17773_ ;
	wire _w17774_ ;
	wire _w17775_ ;
	wire _w17776_ ;
	wire _w17777_ ;
	wire _w17778_ ;
	wire _w17779_ ;
	wire _w17780_ ;
	wire _w17781_ ;
	wire _w17782_ ;
	wire _w17783_ ;
	wire _w17784_ ;
	wire _w17785_ ;
	wire _w17786_ ;
	wire _w17787_ ;
	wire _w17788_ ;
	wire _w17789_ ;
	wire _w17790_ ;
	wire _w17791_ ;
	wire _w17792_ ;
	wire _w17793_ ;
	wire _w17794_ ;
	wire _w17795_ ;
	wire _w17796_ ;
	wire _w17797_ ;
	wire _w17798_ ;
	wire _w17799_ ;
	wire _w17800_ ;
	wire _w17801_ ;
	wire _w17802_ ;
	wire _w17803_ ;
	wire _w17804_ ;
	wire _w17805_ ;
	wire _w17806_ ;
	wire _w17807_ ;
	wire _w17808_ ;
	wire _w17809_ ;
	wire _w17810_ ;
	wire _w17811_ ;
	wire _w17812_ ;
	wire _w17813_ ;
	wire _w17814_ ;
	wire _w17815_ ;
	wire _w17816_ ;
	wire _w17817_ ;
	wire _w17818_ ;
	wire _w17819_ ;
	wire _w17820_ ;
	wire _w17821_ ;
	wire _w17822_ ;
	wire _w17823_ ;
	wire _w17824_ ;
	wire _w17825_ ;
	wire _w17826_ ;
	wire _w17827_ ;
	wire _w17828_ ;
	wire _w17829_ ;
	wire _w17830_ ;
	wire _w17831_ ;
	wire _w17832_ ;
	wire _w17833_ ;
	wire _w17834_ ;
	wire _w17835_ ;
	wire _w17836_ ;
	wire _w17837_ ;
	wire _w17838_ ;
	wire _w17839_ ;
	wire _w17840_ ;
	wire _w17841_ ;
	wire _w17842_ ;
	wire _w17843_ ;
	wire _w17844_ ;
	wire _w17845_ ;
	wire _w17846_ ;
	wire _w17847_ ;
	wire _w17848_ ;
	wire _w17849_ ;
	wire _w17850_ ;
	wire _w17851_ ;
	wire _w17852_ ;
	wire _w17853_ ;
	wire _w17854_ ;
	wire _w17855_ ;
	wire _w17856_ ;
	wire _w17857_ ;
	wire _w17858_ ;
	wire _w17859_ ;
	wire _w17860_ ;
	wire _w17861_ ;
	wire _w17862_ ;
	wire _w17863_ ;
	wire _w17864_ ;
	wire _w17865_ ;
	wire _w17866_ ;
	wire _w17867_ ;
	wire _w17868_ ;
	wire _w17869_ ;
	wire _w17870_ ;
	wire _w17871_ ;
	wire _w17872_ ;
	wire _w17873_ ;
	wire _w17874_ ;
	wire _w17875_ ;
	wire _w17876_ ;
	wire _w17877_ ;
	wire _w17878_ ;
	wire _w17879_ ;
	wire _w17880_ ;
	wire _w17881_ ;
	wire _w17882_ ;
	wire _w17883_ ;
	wire _w17884_ ;
	wire _w17885_ ;
	wire _w17886_ ;
	wire _w17887_ ;
	wire _w17888_ ;
	wire _w17889_ ;
	wire _w17890_ ;
	wire _w17891_ ;
	wire _w17892_ ;
	wire _w17893_ ;
	wire _w17894_ ;
	wire _w17895_ ;
	wire _w17896_ ;
	wire _w17897_ ;
	wire _w17898_ ;
	wire _w17899_ ;
	wire _w17900_ ;
	wire _w17901_ ;
	wire _w17902_ ;
	wire _w17903_ ;
	wire _w17904_ ;
	wire _w17905_ ;
	wire _w17906_ ;
	wire _w17907_ ;
	wire _w17908_ ;
	wire _w17909_ ;
	wire _w17910_ ;
	wire _w17911_ ;
	wire _w17912_ ;
	wire _w17913_ ;
	wire _w17914_ ;
	wire _w17915_ ;
	wire _w17916_ ;
	wire _w17917_ ;
	wire _w17918_ ;
	wire _w17919_ ;
	wire _w17920_ ;
	wire _w17921_ ;
	wire _w17922_ ;
	wire _w17923_ ;
	wire _w17924_ ;
	wire _w17925_ ;
	wire _w17926_ ;
	wire _w17927_ ;
	wire _w17928_ ;
	wire _w17929_ ;
	wire _w17930_ ;
	wire _w17931_ ;
	wire _w17932_ ;
	wire _w17933_ ;
	wire _w17934_ ;
	wire _w17935_ ;
	wire _w17936_ ;
	wire _w17937_ ;
	wire _w17938_ ;
	wire _w17939_ ;
	wire _w17940_ ;
	wire _w17941_ ;
	wire _w17942_ ;
	wire _w17943_ ;
	wire _w17944_ ;
	wire _w17945_ ;
	wire _w17946_ ;
	wire _w17947_ ;
	wire _w17948_ ;
	wire _w17949_ ;
	wire _w17950_ ;
	wire _w17951_ ;
	wire _w17952_ ;
	wire _w17953_ ;
	wire _w17954_ ;
	wire _w17955_ ;
	wire _w17956_ ;
	wire _w17957_ ;
	wire _w17958_ ;
	wire _w17959_ ;
	wire _w17960_ ;
	wire _w17961_ ;
	wire _w17962_ ;
	wire _w17963_ ;
	wire _w17964_ ;
	wire _w17965_ ;
	wire _w17966_ ;
	wire _w17967_ ;
	wire _w17968_ ;
	wire _w17969_ ;
	wire _w17970_ ;
	wire _w17971_ ;
	wire _w17972_ ;
	wire _w17973_ ;
	wire _w17974_ ;
	wire _w17975_ ;
	wire _w17976_ ;
	wire _w17977_ ;
	wire _w17978_ ;
	wire _w17979_ ;
	wire _w17980_ ;
	wire _w17981_ ;
	wire _w17982_ ;
	wire _w17983_ ;
	wire _w17984_ ;
	wire _w17985_ ;
	wire _w17986_ ;
	wire _w17987_ ;
	wire _w17988_ ;
	wire _w17989_ ;
	wire _w17990_ ;
	wire _w17991_ ;
	wire _w17992_ ;
	wire _w17993_ ;
	wire _w17994_ ;
	wire _w17995_ ;
	wire _w17996_ ;
	wire _w17997_ ;
	wire _w17998_ ;
	wire _w17999_ ;
	wire _w18000_ ;
	wire _w18001_ ;
	wire _w18002_ ;
	wire _w18003_ ;
	wire _w18004_ ;
	wire _w18005_ ;
	wire _w18006_ ;
	wire _w18007_ ;
	wire _w18008_ ;
	wire _w18009_ ;
	wire _w18010_ ;
	wire _w18011_ ;
	wire _w18012_ ;
	wire _w18013_ ;
	wire _w18014_ ;
	wire _w18015_ ;
	wire _w18016_ ;
	wire _w18017_ ;
	wire _w18018_ ;
	wire _w18019_ ;
	wire _w18020_ ;
	wire _w18021_ ;
	wire _w18022_ ;
	wire _w18023_ ;
	wire _w18024_ ;
	wire _w18025_ ;
	wire _w18026_ ;
	wire _w18027_ ;
	wire _w18028_ ;
	wire _w18029_ ;
	wire _w18030_ ;
	wire _w18031_ ;
	wire _w18032_ ;
	wire _w18033_ ;
	wire _w18034_ ;
	wire _w18035_ ;
	wire _w18036_ ;
	wire _w18037_ ;
	wire _w18038_ ;
	wire _w18039_ ;
	wire _w18040_ ;
	wire _w18041_ ;
	wire _w18042_ ;
	wire _w18043_ ;
	wire _w18044_ ;
	wire _w18045_ ;
	wire _w18046_ ;
	wire _w18047_ ;
	wire _w18048_ ;
	wire _w18049_ ;
	wire _w18050_ ;
	wire _w18051_ ;
	wire _w18052_ ;
	wire _w18053_ ;
	wire _w18054_ ;
	wire _w18055_ ;
	wire _w18056_ ;
	wire _w18057_ ;
	wire _w18058_ ;
	wire _w18059_ ;
	wire _w18060_ ;
	wire _w18061_ ;
	wire _w18062_ ;
	wire _w18063_ ;
	wire _w18064_ ;
	wire _w18065_ ;
	wire _w18066_ ;
	wire _w18067_ ;
	wire _w18068_ ;
	wire _w18069_ ;
	wire _w18070_ ;
	wire _w18071_ ;
	wire _w18072_ ;
	wire _w18073_ ;
	wire _w18074_ ;
	wire _w18075_ ;
	wire _w18076_ ;
	wire _w18077_ ;
	wire _w18078_ ;
	wire _w18079_ ;
	wire _w18080_ ;
	wire _w18081_ ;
	wire _w18082_ ;
	wire _w18083_ ;
	wire _w18084_ ;
	wire _w18085_ ;
	wire _w18086_ ;
	wire _w18087_ ;
	wire _w18088_ ;
	wire _w18089_ ;
	wire _w18090_ ;
	wire _w18091_ ;
	wire _w18092_ ;
	wire _w18093_ ;
	wire _w18094_ ;
	wire _w18095_ ;
	wire _w18096_ ;
	wire _w18097_ ;
	wire _w18098_ ;
	wire _w18099_ ;
	wire _w18100_ ;
	wire _w18101_ ;
	wire _w18102_ ;
	wire _w18103_ ;
	wire _w18104_ ;
	wire _w18105_ ;
	wire _w18106_ ;
	wire _w18107_ ;
	wire _w18108_ ;
	wire _w18109_ ;
	wire _w18110_ ;
	wire _w18111_ ;
	wire _w18112_ ;
	wire _w18113_ ;
	wire _w18114_ ;
	wire _w18115_ ;
	wire _w18116_ ;
	wire _w18117_ ;
	wire _w18118_ ;
	wire _w18119_ ;
	wire _w18120_ ;
	wire _w18121_ ;
	wire _w18122_ ;
	wire _w18123_ ;
	wire _w18124_ ;
	wire _w18125_ ;
	wire _w18126_ ;
	wire _w18127_ ;
	wire _w18128_ ;
	wire _w18129_ ;
	wire _w18130_ ;
	wire _w18131_ ;
	wire _w18132_ ;
	wire _w18133_ ;
	wire _w18134_ ;
	wire _w18135_ ;
	wire _w18136_ ;
	wire _w18137_ ;
	wire _w18138_ ;
	wire _w18139_ ;
	wire _w18140_ ;
	wire _w18141_ ;
	wire _w18142_ ;
	wire _w18143_ ;
	wire _w18144_ ;
	wire _w18145_ ;
	wire _w18146_ ;
	wire _w18147_ ;
	wire _w18148_ ;
	wire _w18149_ ;
	wire _w18150_ ;
	wire _w18151_ ;
	wire _w18152_ ;
	wire _w18153_ ;
	wire _w18154_ ;
	wire _w18155_ ;
	wire _w18156_ ;
	wire _w18157_ ;
	wire _w18158_ ;
	wire _w18159_ ;
	wire _w18160_ ;
	wire _w18161_ ;
	wire _w18162_ ;
	wire _w18163_ ;
	wire _w18164_ ;
	wire _w18165_ ;
	wire _w18166_ ;
	wire _w18167_ ;
	wire _w18168_ ;
	wire _w18169_ ;
	wire _w18170_ ;
	wire _w18171_ ;
	wire _w18172_ ;
	wire _w18173_ ;
	wire _w18174_ ;
	wire _w18175_ ;
	wire _w18176_ ;
	wire _w18177_ ;
	wire _w18178_ ;
	wire _w18179_ ;
	wire _w18180_ ;
	wire _w18181_ ;
	wire _w18182_ ;
	wire _w18183_ ;
	wire _w18184_ ;
	wire _w18185_ ;
	wire _w18186_ ;
	wire _w18187_ ;
	wire _w18188_ ;
	wire _w18189_ ;
	wire _w18190_ ;
	wire _w18191_ ;
	wire _w18192_ ;
	wire _w18193_ ;
	wire _w18194_ ;
	wire _w18195_ ;
	wire _w18196_ ;
	wire _w18197_ ;
	wire _w18198_ ;
	wire _w18199_ ;
	wire _w18200_ ;
	wire _w18201_ ;
	wire _w18202_ ;
	wire _w18203_ ;
	wire _w18204_ ;
	wire _w18205_ ;
	wire _w18206_ ;
	wire _w18207_ ;
	wire _w18208_ ;
	wire _w18209_ ;
	wire _w18210_ ;
	wire _w18211_ ;
	wire _w18212_ ;
	wire _w18213_ ;
	wire _w18214_ ;
	wire _w18215_ ;
	wire _w18216_ ;
	wire _w18217_ ;
	wire _w18218_ ;
	wire _w18219_ ;
	wire _w18220_ ;
	wire _w18221_ ;
	wire _w18222_ ;
	wire _w18223_ ;
	wire _w18224_ ;
	wire _w18225_ ;
	wire _w18226_ ;
	wire _w18227_ ;
	wire _w18228_ ;
	wire _w18229_ ;
	wire _w18230_ ;
	wire _w18231_ ;
	wire _w18232_ ;
	wire _w18233_ ;
	wire _w18234_ ;
	wire _w18235_ ;
	wire _w18236_ ;
	wire _w18237_ ;
	wire _w18238_ ;
	wire _w18239_ ;
	wire _w18240_ ;
	wire _w18241_ ;
	wire _w18242_ ;
	wire _w18243_ ;
	wire _w18244_ ;
	wire _w18245_ ;
	wire _w18246_ ;
	wire _w18247_ ;
	wire _w18248_ ;
	wire _w18249_ ;
	wire _w18250_ ;
	wire _w18251_ ;
	wire _w18252_ ;
	wire _w18253_ ;
	wire _w18254_ ;
	wire _w18255_ ;
	wire _w18256_ ;
	wire _w18257_ ;
	wire _w18258_ ;
	wire _w18259_ ;
	wire _w18260_ ;
	wire _w18261_ ;
	wire _w18262_ ;
	wire _w18263_ ;
	wire _w18264_ ;
	wire _w18265_ ;
	wire _w18266_ ;
	wire _w18267_ ;
	wire _w18268_ ;
	wire _w18269_ ;
	wire _w18270_ ;
	wire _w18271_ ;
	wire _w18272_ ;
	wire _w18273_ ;
	wire _w18274_ ;
	wire _w18275_ ;
	wire _w18276_ ;
	wire _w18277_ ;
	wire _w18278_ ;
	wire _w18279_ ;
	wire _w18280_ ;
	wire _w18281_ ;
	wire _w18282_ ;
	wire _w18283_ ;
	wire _w18284_ ;
	wire _w18285_ ;
	wire _w18286_ ;
	wire _w18287_ ;
	wire _w18288_ ;
	wire _w18289_ ;
	wire _w18290_ ;
	wire _w18291_ ;
	wire _w18292_ ;
	wire _w18293_ ;
	wire _w18294_ ;
	wire _w18295_ ;
	wire _w18296_ ;
	wire _w18297_ ;
	wire _w18298_ ;
	wire _w18299_ ;
	wire _w18300_ ;
	wire _w18301_ ;
	wire _w18302_ ;
	wire _w18303_ ;
	wire _w18304_ ;
	wire _w18305_ ;
	wire _w18306_ ;
	wire _w18307_ ;
	wire _w18308_ ;
	wire _w18309_ ;
	wire _w18310_ ;
	wire _w18311_ ;
	wire _w18312_ ;
	wire _w18313_ ;
	wire _w18314_ ;
	wire _w18315_ ;
	wire _w18316_ ;
	wire _w18317_ ;
	wire _w18318_ ;
	wire _w18319_ ;
	wire _w18320_ ;
	wire _w18321_ ;
	wire _w18322_ ;
	wire _w18323_ ;
	wire _w18324_ ;
	wire _w18325_ ;
	wire _w18326_ ;
	wire _w18327_ ;
	wire _w18328_ ;
	wire _w18329_ ;
	wire _w18330_ ;
	wire _w18331_ ;
	wire _w18332_ ;
	wire _w18333_ ;
	wire _w18334_ ;
	wire _w18335_ ;
	wire _w18336_ ;
	wire _w18337_ ;
	wire _w18338_ ;
	wire _w18339_ ;
	wire _w18340_ ;
	wire _w18341_ ;
	wire _w18342_ ;
	wire _w18343_ ;
	wire _w18344_ ;
	wire _w18345_ ;
	wire _w18346_ ;
	wire _w18347_ ;
	wire _w18348_ ;
	wire _w18349_ ;
	wire _w18350_ ;
	wire _w18351_ ;
	wire _w18352_ ;
	wire _w18353_ ;
	wire _w18354_ ;
	wire _w18355_ ;
	wire _w18356_ ;
	wire _w18357_ ;
	wire _w18358_ ;
	wire _w18359_ ;
	wire _w18360_ ;
	wire _w18361_ ;
	wire _w18362_ ;
	wire _w18363_ ;
	wire _w18364_ ;
	wire _w18365_ ;
	wire _w18366_ ;
	wire _w18367_ ;
	wire _w18368_ ;
	wire _w18369_ ;
	wire _w18370_ ;
	wire _w18371_ ;
	wire _w18372_ ;
	wire _w18373_ ;
	wire _w18374_ ;
	wire _w18375_ ;
	wire _w18376_ ;
	wire _w18377_ ;
	wire _w18378_ ;
	wire _w18379_ ;
	wire _w18380_ ;
	wire _w18381_ ;
	wire _w18382_ ;
	wire _w18383_ ;
	wire _w18384_ ;
	wire _w18385_ ;
	wire _w18386_ ;
	wire _w18387_ ;
	wire _w18388_ ;
	wire _w18389_ ;
	wire _w18390_ ;
	wire _w18391_ ;
	wire _w18392_ ;
	wire _w18393_ ;
	wire _w18394_ ;
	wire _w18395_ ;
	wire _w18396_ ;
	wire _w18397_ ;
	wire _w18398_ ;
	wire _w18399_ ;
	wire _w18400_ ;
	wire _w18401_ ;
	wire _w18402_ ;
	wire _w18403_ ;
	wire _w18404_ ;
	wire _w18405_ ;
	wire _w18406_ ;
	wire _w18407_ ;
	wire _w18408_ ;
	wire _w18409_ ;
	wire _w18410_ ;
	wire _w18411_ ;
	wire _w18412_ ;
	wire _w18413_ ;
	wire _w18414_ ;
	wire _w18415_ ;
	wire _w18416_ ;
	wire _w18417_ ;
	wire _w18418_ ;
	wire _w18419_ ;
	wire _w18420_ ;
	wire _w18421_ ;
	wire _w18422_ ;
	wire _w18423_ ;
	wire _w18424_ ;
	wire _w18425_ ;
	wire _w18426_ ;
	wire _w18427_ ;
	wire _w18428_ ;
	wire _w18429_ ;
	wire _w18430_ ;
	wire _w18431_ ;
	wire _w18432_ ;
	wire _w18433_ ;
	wire _w18434_ ;
	wire _w18435_ ;
	wire _w18436_ ;
	wire _w18437_ ;
	wire _w18438_ ;
	wire _w18439_ ;
	wire _w18440_ ;
	wire _w18441_ ;
	wire _w18442_ ;
	wire _w18443_ ;
	wire _w18444_ ;
	wire _w18445_ ;
	wire _w18446_ ;
	wire _w18447_ ;
	wire _w18448_ ;
	wire _w18449_ ;
	wire _w18450_ ;
	wire _w18451_ ;
	wire _w18452_ ;
	wire _w18453_ ;
	wire _w18454_ ;
	wire _w18455_ ;
	wire _w18456_ ;
	wire _w18457_ ;
	wire _w18458_ ;
	wire _w18459_ ;
	wire _w18460_ ;
	wire _w18461_ ;
	wire _w18462_ ;
	wire _w18463_ ;
	wire _w18464_ ;
	wire _w18465_ ;
	wire _w18466_ ;
	wire _w18467_ ;
	wire _w18468_ ;
	wire _w18469_ ;
	wire _w18470_ ;
	wire _w18471_ ;
	wire _w18472_ ;
	wire _w18473_ ;
	wire _w18474_ ;
	wire _w18475_ ;
	wire _w18476_ ;
	wire _w18477_ ;
	wire _w18478_ ;
	wire _w18479_ ;
	wire _w18480_ ;
	wire _w18481_ ;
	wire _w18482_ ;
	wire _w18483_ ;
	wire _w18484_ ;
	wire _w18485_ ;
	wire _w18486_ ;
	wire _w18487_ ;
	wire _w18488_ ;
	wire _w18489_ ;
	wire _w18490_ ;
	wire _w18491_ ;
	wire _w18492_ ;
	wire _w18493_ ;
	wire _w18494_ ;
	wire _w18495_ ;
	wire _w18496_ ;
	wire _w18497_ ;
	wire _w18498_ ;
	wire _w18499_ ;
	wire _w18500_ ;
	wire _w18501_ ;
	wire _w18502_ ;
	wire _w18503_ ;
	wire _w18504_ ;
	wire _w18505_ ;
	wire _w18506_ ;
	wire _w18507_ ;
	wire _w18508_ ;
	wire _w18509_ ;
	wire _w18510_ ;
	wire _w18511_ ;
	wire _w18512_ ;
	wire _w18513_ ;
	wire _w18514_ ;
	wire _w18515_ ;
	wire _w18516_ ;
	wire _w18517_ ;
	wire _w18518_ ;
	wire _w18519_ ;
	wire _w18520_ ;
	wire _w18521_ ;
	wire _w18522_ ;
	wire _w18523_ ;
	wire _w18524_ ;
	wire _w18525_ ;
	wire _w18526_ ;
	wire _w18527_ ;
	wire _w18528_ ;
	wire _w18529_ ;
	wire _w18530_ ;
	wire _w18531_ ;
	wire _w18532_ ;
	wire _w18533_ ;
	wire _w18534_ ;
	wire _w18535_ ;
	wire _w18536_ ;
	wire _w18537_ ;
	wire _w18538_ ;
	wire _w18539_ ;
	wire _w18540_ ;
	wire _w18541_ ;
	wire _w18542_ ;
	wire _w18543_ ;
	wire _w18544_ ;
	wire _w18545_ ;
	wire _w18546_ ;
	wire _w18547_ ;
	wire _w18548_ ;
	wire _w18549_ ;
	wire _w18550_ ;
	wire _w18551_ ;
	wire _w18552_ ;
	wire _w18553_ ;
	wire _w18554_ ;
	wire _w18555_ ;
	wire _w18556_ ;
	wire _w18557_ ;
	wire _w18558_ ;
	wire _w18559_ ;
	wire _w18560_ ;
	wire _w18561_ ;
	wire _w18562_ ;
	wire _w18563_ ;
	wire _w18564_ ;
	wire _w18565_ ;
	wire _w18566_ ;
	wire _w18567_ ;
	wire _w18568_ ;
	wire _w18569_ ;
	wire _w18570_ ;
	wire _w18571_ ;
	wire _w18572_ ;
	wire _w18573_ ;
	wire _w18574_ ;
	wire _w18575_ ;
	wire _w18576_ ;
	wire _w18577_ ;
	wire _w18578_ ;
	wire _w18579_ ;
	wire _w18580_ ;
	wire _w18581_ ;
	wire _w18582_ ;
	wire _w18583_ ;
	wire _w18584_ ;
	wire _w18585_ ;
	wire _w18586_ ;
	wire _w18587_ ;
	wire _w18588_ ;
	wire _w18589_ ;
	wire _w18590_ ;
	wire _w18591_ ;
	wire _w18592_ ;
	wire _w18593_ ;
	wire _w18594_ ;
	wire _w18595_ ;
	wire _w18596_ ;
	wire _w18597_ ;
	wire _w18598_ ;
	wire _w18599_ ;
	wire _w18600_ ;
	wire _w18601_ ;
	wire _w18602_ ;
	wire _w18603_ ;
	wire _w18604_ ;
	wire _w18605_ ;
	wire _w18606_ ;
	wire _w18607_ ;
	wire _w18608_ ;
	wire _w18609_ ;
	wire _w18610_ ;
	wire _w18611_ ;
	wire _w18612_ ;
	wire _w18613_ ;
	wire _w18614_ ;
	wire _w18615_ ;
	wire _w18616_ ;
	wire _w18617_ ;
	wire _w18618_ ;
	wire _w18619_ ;
	wire _w18620_ ;
	wire _w18621_ ;
	wire _w18622_ ;
	wire _w18623_ ;
	wire _w18624_ ;
	wire _w18625_ ;
	wire _w18626_ ;
	wire _w18627_ ;
	wire _w18628_ ;
	wire _w18629_ ;
	wire _w18630_ ;
	wire _w18631_ ;
	wire _w18632_ ;
	wire _w18633_ ;
	wire _w18634_ ;
	wire _w18635_ ;
	wire _w18636_ ;
	wire _w18637_ ;
	wire _w18638_ ;
	wire _w18639_ ;
	wire _w18640_ ;
	wire _w18641_ ;
	wire _w18642_ ;
	wire _w18643_ ;
	wire _w18644_ ;
	wire _w18645_ ;
	wire _w18646_ ;
	wire _w18647_ ;
	wire _w18648_ ;
	wire _w18649_ ;
	wire _w18650_ ;
	wire _w18651_ ;
	wire _w18652_ ;
	wire _w18653_ ;
	wire _w18654_ ;
	wire _w18655_ ;
	wire _w18656_ ;
	wire _w18657_ ;
	wire _w18658_ ;
	wire _w18659_ ;
	wire _w18660_ ;
	wire _w18661_ ;
	wire _w18662_ ;
	wire _w18663_ ;
	wire _w18664_ ;
	wire _w18665_ ;
	wire _w18666_ ;
	wire _w18667_ ;
	wire _w18668_ ;
	wire _w18669_ ;
	wire _w18670_ ;
	wire _w18671_ ;
	wire _w18672_ ;
	wire _w18673_ ;
	wire _w18674_ ;
	wire _w18675_ ;
	wire _w18676_ ;
	wire _w18677_ ;
	wire _w18678_ ;
	wire _w18679_ ;
	wire _w18680_ ;
	wire _w18681_ ;
	wire _w18682_ ;
	wire _w18683_ ;
	wire _w18684_ ;
	wire _w18685_ ;
	wire _w18686_ ;
	wire _w18687_ ;
	wire _w18688_ ;
	wire _w18689_ ;
	wire _w18690_ ;
	wire _w18691_ ;
	wire _w18692_ ;
	wire _w18693_ ;
	wire _w18694_ ;
	wire _w18695_ ;
	wire _w18696_ ;
	wire _w18697_ ;
	wire _w18698_ ;
	wire _w18699_ ;
	wire _w18700_ ;
	wire _w18701_ ;
	wire _w18702_ ;
	wire _w18703_ ;
	wire _w18704_ ;
	wire _w18705_ ;
	wire _w18706_ ;
	wire _w18707_ ;
	wire _w18708_ ;
	wire _w18709_ ;
	wire _w18710_ ;
	wire _w18711_ ;
	wire _w18712_ ;
	wire _w18713_ ;
	wire _w18714_ ;
	wire _w18715_ ;
	wire _w18716_ ;
	wire _w18717_ ;
	wire _w18718_ ;
	wire _w18719_ ;
	wire _w18720_ ;
	wire _w18721_ ;
	wire _w18722_ ;
	wire _w18723_ ;
	wire _w18724_ ;
	wire _w18725_ ;
	wire _w18726_ ;
	wire _w18727_ ;
	wire _w18728_ ;
	wire _w18729_ ;
	wire _w18730_ ;
	wire _w18731_ ;
	wire _w18732_ ;
	wire _w18733_ ;
	wire _w18734_ ;
	wire _w18735_ ;
	wire _w18736_ ;
	wire _w18737_ ;
	wire _w18738_ ;
	wire _w18739_ ;
	wire _w18740_ ;
	wire _w18741_ ;
	wire _w18742_ ;
	wire _w18743_ ;
	wire _w18744_ ;
	wire _w18745_ ;
	wire _w18746_ ;
	wire _w18747_ ;
	wire _w18748_ ;
	wire _w18749_ ;
	wire _w18750_ ;
	wire _w18751_ ;
	wire _w18752_ ;
	wire _w18753_ ;
	wire _w18754_ ;
	wire _w18755_ ;
	wire _w18756_ ;
	wire _w18757_ ;
	wire _w18758_ ;
	wire _w18759_ ;
	wire _w18760_ ;
	wire _w18761_ ;
	wire _w18762_ ;
	wire _w18763_ ;
	wire _w18764_ ;
	wire _w18765_ ;
	wire _w18766_ ;
	wire _w18767_ ;
	wire _w18768_ ;
	wire _w18769_ ;
	wire _w18770_ ;
	wire _w18771_ ;
	wire _w18772_ ;
	wire _w18773_ ;
	wire _w18774_ ;
	wire _w18775_ ;
	wire _w18776_ ;
	wire _w18777_ ;
	wire _w18778_ ;
	wire _w18779_ ;
	wire _w18780_ ;
	wire _w18781_ ;
	wire _w18782_ ;
	wire _w18783_ ;
	wire _w18784_ ;
	wire _w18785_ ;
	wire _w18786_ ;
	wire _w18787_ ;
	wire _w18788_ ;
	wire _w18789_ ;
	wire _w18790_ ;
	wire _w18791_ ;
	wire _w18792_ ;
	wire _w18793_ ;
	wire _w18794_ ;
	wire _w18795_ ;
	wire _w18796_ ;
	wire _w18797_ ;
	wire _w18798_ ;
	wire _w18799_ ;
	wire _w18800_ ;
	wire _w18801_ ;
	wire _w18802_ ;
	wire _w18803_ ;
	wire _w18804_ ;
	wire _w18805_ ;
	wire _w18806_ ;
	wire _w18807_ ;
	wire _w18808_ ;
	wire _w18809_ ;
	wire _w18810_ ;
	wire _w18811_ ;
	wire _w18812_ ;
	wire _w18813_ ;
	wire _w18814_ ;
	wire _w18815_ ;
	wire _w18816_ ;
	wire _w18817_ ;
	wire _w18818_ ;
	wire _w18819_ ;
	wire _w18820_ ;
	wire _w18821_ ;
	wire _w18822_ ;
	wire _w18823_ ;
	wire _w18824_ ;
	wire _w18825_ ;
	wire _w18826_ ;
	wire _w18827_ ;
	wire _w18828_ ;
	wire _w18829_ ;
	wire _w18830_ ;
	wire _w18831_ ;
	wire _w18832_ ;
	wire _w18833_ ;
	wire _w18834_ ;
	wire _w18835_ ;
	wire _w18836_ ;
	wire _w18837_ ;
	wire _w18838_ ;
	wire _w18839_ ;
	wire _w18840_ ;
	wire _w18841_ ;
	wire _w18842_ ;
	wire _w18843_ ;
	wire _w18844_ ;
	wire _w18845_ ;
	wire _w18846_ ;
	wire _w18847_ ;
	wire _w18848_ ;
	wire _w18849_ ;
	wire _w18850_ ;
	wire _w18851_ ;
	wire _w18852_ ;
	wire _w18853_ ;
	wire _w18854_ ;
	wire _w18855_ ;
	wire _w18856_ ;
	wire _w18857_ ;
	wire _w18858_ ;
	wire _w18859_ ;
	wire _w18860_ ;
	wire _w18861_ ;
	wire _w18862_ ;
	wire _w18863_ ;
	wire _w18864_ ;
	wire _w18865_ ;
	wire _w18866_ ;
	wire _w18867_ ;
	wire _w18868_ ;
	wire _w18869_ ;
	wire _w18870_ ;
	wire _w18871_ ;
	wire _w18872_ ;
	wire _w18873_ ;
	wire _w18874_ ;
	wire _w18875_ ;
	wire _w18876_ ;
	wire _w18877_ ;
	wire _w18878_ ;
	wire _w18879_ ;
	wire _w18880_ ;
	wire _w18881_ ;
	wire _w18882_ ;
	wire _w18883_ ;
	wire _w18884_ ;
	wire _w18885_ ;
	wire _w18886_ ;
	wire _w18887_ ;
	wire _w18888_ ;
	wire _w18889_ ;
	wire _w18890_ ;
	wire _w18891_ ;
	wire _w18892_ ;
	wire _w18893_ ;
	wire _w18894_ ;
	wire _w18895_ ;
	wire _w18896_ ;
	wire _w18897_ ;
	wire _w18898_ ;
	wire _w18899_ ;
	wire _w18900_ ;
	wire _w18901_ ;
	wire _w18902_ ;
	wire _w18903_ ;
	wire _w18904_ ;
	wire _w18905_ ;
	wire _w18906_ ;
	wire _w18907_ ;
	wire _w18908_ ;
	wire _w18909_ ;
	wire _w18910_ ;
	wire _w18911_ ;
	wire _w18912_ ;
	wire _w18913_ ;
	wire _w18914_ ;
	wire _w18915_ ;
	wire _w18916_ ;
	wire _w18917_ ;
	wire _w18918_ ;
	wire _w18919_ ;
	wire _w18920_ ;
	wire _w18921_ ;
	wire _w18922_ ;
	wire _w18923_ ;
	wire _w18924_ ;
	wire _w18925_ ;
	wire _w18926_ ;
	wire _w18927_ ;
	wire _w18928_ ;
	wire _w18929_ ;
	wire _w18930_ ;
	wire _w18931_ ;
	wire _w18932_ ;
	wire _w18933_ ;
	wire _w18934_ ;
	wire _w18935_ ;
	wire _w18936_ ;
	wire _w18937_ ;
	wire _w18938_ ;
	wire _w18939_ ;
	wire _w18940_ ;
	wire _w18941_ ;
	wire _w18942_ ;
	wire _w18943_ ;
	wire _w18944_ ;
	wire _w18945_ ;
	wire _w18946_ ;
	wire _w18947_ ;
	wire _w18948_ ;
	wire _w18949_ ;
	wire _w18950_ ;
	wire _w18951_ ;
	wire _w18952_ ;
	wire _w18953_ ;
	wire _w18954_ ;
	wire _w18955_ ;
	wire _w18956_ ;
	wire _w18957_ ;
	wire _w18958_ ;
	wire _w18959_ ;
	wire _w18960_ ;
	wire _w18961_ ;
	wire _w18962_ ;
	wire _w18963_ ;
	wire _w18964_ ;
	wire _w18965_ ;
	wire _w18966_ ;
	wire _w18967_ ;
	wire _w18968_ ;
	wire _w18969_ ;
	wire _w18970_ ;
	wire _w18971_ ;
	wire _w18972_ ;
	wire _w18973_ ;
	wire _w18974_ ;
	wire _w18975_ ;
	wire _w18976_ ;
	wire _w18977_ ;
	wire _w18978_ ;
	wire _w18979_ ;
	wire _w18980_ ;
	wire _w18981_ ;
	wire _w18982_ ;
	wire _w18983_ ;
	wire _w18984_ ;
	wire _w18985_ ;
	wire _w18986_ ;
	wire _w18987_ ;
	wire _w18988_ ;
	wire _w18989_ ;
	wire _w18990_ ;
	wire _w18991_ ;
	wire _w18992_ ;
	wire _w18993_ ;
	wire _w18994_ ;
	wire _w18995_ ;
	wire _w18996_ ;
	wire _w18997_ ;
	wire _w18998_ ;
	wire _w18999_ ;
	wire _w19000_ ;
	wire _w19001_ ;
	wire _w19002_ ;
	wire _w19003_ ;
	wire _w19004_ ;
	wire _w19005_ ;
	wire _w19006_ ;
	wire _w19007_ ;
	wire _w19008_ ;
	wire _w19009_ ;
	wire _w19010_ ;
	wire _w19011_ ;
	wire _w19012_ ;
	wire _w19013_ ;
	wire _w19014_ ;
	wire _w19015_ ;
	wire _w19016_ ;
	wire _w19017_ ;
	wire _w19018_ ;
	wire _w19019_ ;
	wire _w19020_ ;
	wire _w19021_ ;
	wire _w19022_ ;
	wire _w19023_ ;
	wire _w19024_ ;
	wire _w19025_ ;
	wire _w19026_ ;
	wire _w19027_ ;
	wire _w19028_ ;
	wire _w19029_ ;
	wire _w19030_ ;
	wire _w19031_ ;
	wire _w19032_ ;
	wire _w19033_ ;
	wire _w19034_ ;
	wire _w19035_ ;
	wire _w19036_ ;
	wire _w19037_ ;
	wire _w19038_ ;
	wire _w19039_ ;
	wire _w19040_ ;
	wire _w19041_ ;
	wire _w19042_ ;
	wire _w19043_ ;
	wire _w19044_ ;
	wire _w19045_ ;
	wire _w19046_ ;
	wire _w19047_ ;
	wire _w19048_ ;
	wire _w19049_ ;
	wire _w19050_ ;
	wire _w19051_ ;
	wire _w19052_ ;
	wire _w19053_ ;
	wire _w19054_ ;
	wire _w19055_ ;
	wire _w19056_ ;
	wire _w19057_ ;
	wire _w19058_ ;
	wire _w19059_ ;
	wire _w19060_ ;
	wire _w19061_ ;
	wire _w19062_ ;
	wire _w19063_ ;
	wire _w19064_ ;
	wire _w19065_ ;
	wire _w19066_ ;
	wire _w19067_ ;
	wire _w19068_ ;
	wire _w19069_ ;
	wire _w19070_ ;
	wire _w19071_ ;
	wire _w19072_ ;
	wire _w19073_ ;
	wire _w19074_ ;
	wire _w19075_ ;
	wire _w19076_ ;
	wire _w19077_ ;
	wire _w19078_ ;
	wire _w19079_ ;
	wire _w19080_ ;
	wire _w19081_ ;
	wire _w19082_ ;
	wire _w19083_ ;
	wire _w19084_ ;
	wire _w19085_ ;
	wire _w19086_ ;
	wire _w19087_ ;
	wire _w19088_ ;
	wire _w19089_ ;
	wire _w19090_ ;
	wire _w19091_ ;
	wire _w19092_ ;
	wire _w19093_ ;
	wire _w19094_ ;
	wire _w19095_ ;
	wire _w19096_ ;
	wire _w19097_ ;
	wire _w19098_ ;
	wire _w19099_ ;
	wire _w19100_ ;
	wire _w19101_ ;
	wire _w19102_ ;
	wire _w19103_ ;
	wire _w19104_ ;
	wire _w19105_ ;
	wire _w19106_ ;
	wire _w19107_ ;
	wire _w19108_ ;
	wire _w19109_ ;
	wire _w19110_ ;
	wire _w19111_ ;
	wire _w19112_ ;
	wire _w19113_ ;
	wire _w19114_ ;
	wire _w19115_ ;
	wire _w19116_ ;
	wire _w19117_ ;
	wire _w19118_ ;
	wire _w19119_ ;
	wire _w19120_ ;
	wire _w19121_ ;
	wire _w19122_ ;
	wire _w19123_ ;
	wire _w19124_ ;
	wire _w19125_ ;
	wire _w19126_ ;
	wire _w19127_ ;
	wire _w19128_ ;
	wire _w19129_ ;
	wire _w19130_ ;
	wire _w19131_ ;
	wire _w19132_ ;
	wire _w19133_ ;
	wire _w19134_ ;
	wire _w19135_ ;
	wire _w19136_ ;
	wire _w19137_ ;
	wire _w19138_ ;
	wire _w19139_ ;
	wire _w19140_ ;
	wire _w19141_ ;
	wire _w19142_ ;
	wire _w19143_ ;
	wire _w19144_ ;
	wire _w19145_ ;
	wire _w19146_ ;
	wire _w19147_ ;
	wire _w19148_ ;
	wire _w19149_ ;
	wire _w19150_ ;
	wire _w19151_ ;
	wire _w19152_ ;
	wire _w19153_ ;
	wire _w19154_ ;
	wire _w19155_ ;
	wire _w19156_ ;
	wire _w19157_ ;
	wire _w19158_ ;
	wire _w19159_ ;
	wire _w19160_ ;
	wire _w19161_ ;
	wire _w19162_ ;
	wire _w19163_ ;
	wire _w19164_ ;
	wire _w19165_ ;
	wire _w19166_ ;
	wire _w19167_ ;
	wire _w19168_ ;
	wire _w19169_ ;
	wire _w19170_ ;
	wire _w19171_ ;
	wire _w19172_ ;
	wire _w19173_ ;
	wire _w19174_ ;
	wire _w19175_ ;
	wire _w19176_ ;
	wire _w19177_ ;
	wire _w19178_ ;
	wire _w19179_ ;
	wire _w19180_ ;
	wire _w19181_ ;
	wire _w19182_ ;
	wire _w19183_ ;
	wire _w19184_ ;
	wire _w19185_ ;
	wire _w19186_ ;
	wire _w19187_ ;
	wire _w19188_ ;
	wire _w19189_ ;
	wire _w19190_ ;
	wire _w19191_ ;
	wire _w19192_ ;
	wire _w19193_ ;
	wire _w19194_ ;
	wire _w19195_ ;
	wire _w19196_ ;
	wire _w19197_ ;
	wire _w19198_ ;
	wire _w19199_ ;
	wire _w19200_ ;
	wire _w19201_ ;
	wire _w19202_ ;
	wire _w19203_ ;
	wire _w19204_ ;
	wire _w19205_ ;
	wire _w19206_ ;
	wire _w19207_ ;
	wire _w19208_ ;
	wire _w19209_ ;
	wire _w19210_ ;
	wire _w19211_ ;
	wire _w19212_ ;
	wire _w19213_ ;
	wire _w19214_ ;
	wire _w19215_ ;
	wire _w19216_ ;
	wire _w19217_ ;
	wire _w19218_ ;
	wire _w19219_ ;
	wire _w19220_ ;
	wire _w19221_ ;
	wire _w19222_ ;
	wire _w19223_ ;
	wire _w19224_ ;
	wire _w19225_ ;
	wire _w19226_ ;
	wire _w19227_ ;
	wire _w19228_ ;
	wire _w19229_ ;
	wire _w19230_ ;
	wire _w19231_ ;
	wire _w19232_ ;
	wire _w19233_ ;
	wire _w19234_ ;
	wire _w19235_ ;
	wire _w19236_ ;
	wire _w19237_ ;
	wire _w19238_ ;
	wire _w19239_ ;
	wire _w19240_ ;
	wire _w19241_ ;
	wire _w19242_ ;
	wire _w19243_ ;
	wire _w19244_ ;
	wire _w19245_ ;
	wire _w19246_ ;
	wire _w19247_ ;
	wire _w19248_ ;
	wire _w19249_ ;
	wire _w19250_ ;
	wire _w19251_ ;
	wire _w19252_ ;
	wire _w19253_ ;
	wire _w19254_ ;
	wire _w19255_ ;
	wire _w19256_ ;
	wire _w19257_ ;
	wire _w19258_ ;
	wire _w19259_ ;
	wire _w19260_ ;
	wire _w19261_ ;
	wire _w19262_ ;
	wire _w19263_ ;
	wire _w19264_ ;
	wire _w19265_ ;
	wire _w19266_ ;
	wire _w19267_ ;
	wire _w19268_ ;
	wire _w19269_ ;
	wire _w19270_ ;
	wire _w19271_ ;
	wire _w19272_ ;
	wire _w19273_ ;
	wire _w19274_ ;
	wire _w19275_ ;
	wire _w19276_ ;
	wire _w19277_ ;
	wire _w19278_ ;
	wire _w19279_ ;
	wire _w19280_ ;
	wire _w19281_ ;
	wire _w19282_ ;
	wire _w19283_ ;
	wire _w19284_ ;
	wire _w19285_ ;
	wire _w19286_ ;
	wire _w19287_ ;
	wire _w19288_ ;
	wire _w19289_ ;
	wire _w19290_ ;
	wire _w19291_ ;
	wire _w19292_ ;
	wire _w19293_ ;
	wire _w19294_ ;
	wire _w19295_ ;
	wire _w19296_ ;
	wire _w19297_ ;
	wire _w19298_ ;
	wire _w19299_ ;
	wire _w19300_ ;
	wire _w19301_ ;
	wire _w19302_ ;
	wire _w19303_ ;
	wire _w19304_ ;
	wire _w19305_ ;
	wire _w19306_ ;
	wire _w19307_ ;
	wire _w19308_ ;
	wire _w19309_ ;
	wire _w19310_ ;
	wire _w19311_ ;
	wire _w19312_ ;
	wire _w19313_ ;
	wire _w19314_ ;
	wire _w19315_ ;
	wire _w19316_ ;
	wire _w19317_ ;
	wire _w19318_ ;
	wire _w19319_ ;
	wire _w19320_ ;
	wire _w19321_ ;
	wire _w19322_ ;
	wire _w19323_ ;
	wire _w19324_ ;
	wire _w19325_ ;
	wire _w19326_ ;
	wire _w19327_ ;
	wire _w19328_ ;
	wire _w19329_ ;
	wire _w19330_ ;
	wire _w19331_ ;
	wire _w19332_ ;
	wire _w19333_ ;
	wire _w19334_ ;
	wire _w19335_ ;
	wire _w19336_ ;
	wire _w19337_ ;
	wire _w19338_ ;
	wire _w19339_ ;
	wire _w19340_ ;
	wire _w19341_ ;
	wire _w19342_ ;
	wire _w19343_ ;
	wire _w19344_ ;
	wire _w19345_ ;
	wire _w19346_ ;
	wire _w19347_ ;
	wire _w19348_ ;
	wire _w19349_ ;
	wire _w19350_ ;
	wire _w19351_ ;
	wire _w19352_ ;
	wire _w19353_ ;
	wire _w19354_ ;
	wire _w19355_ ;
	wire _w19356_ ;
	wire _w19357_ ;
	wire _w19358_ ;
	wire _w19359_ ;
	wire _w19360_ ;
	wire _w19361_ ;
	wire _w19362_ ;
	wire _w19363_ ;
	wire _w19364_ ;
	wire _w19365_ ;
	wire _w19366_ ;
	wire _w19367_ ;
	wire _w19368_ ;
	wire _w19369_ ;
	wire _w19370_ ;
	wire _w19371_ ;
	wire _w19372_ ;
	wire _w19373_ ;
	wire _w19374_ ;
	wire _w19375_ ;
	wire _w19376_ ;
	wire _w19377_ ;
	wire _w19378_ ;
	wire _w19379_ ;
	wire _w19380_ ;
	wire _w19381_ ;
	wire _w19382_ ;
	wire _w19383_ ;
	wire _w19384_ ;
	wire _w19385_ ;
	wire _w19386_ ;
	wire _w19387_ ;
	wire _w19388_ ;
	wire _w19389_ ;
	wire _w19390_ ;
	wire _w19391_ ;
	wire _w19392_ ;
	wire _w19393_ ;
	wire _w19394_ ;
	wire _w19395_ ;
	wire _w19396_ ;
	wire _w19397_ ;
	wire _w19398_ ;
	wire _w19399_ ;
	wire _w19400_ ;
	wire _w19401_ ;
	wire _w19402_ ;
	wire _w19403_ ;
	wire _w19404_ ;
	wire _w19405_ ;
	wire _w19406_ ;
	wire _w19407_ ;
	wire _w19408_ ;
	wire _w19409_ ;
	wire _w19410_ ;
	wire _w19411_ ;
	wire _w19412_ ;
	wire _w19413_ ;
	wire _w19414_ ;
	wire _w19415_ ;
	wire _w19416_ ;
	wire _w19417_ ;
	wire _w19418_ ;
	wire _w19419_ ;
	wire _w19420_ ;
	wire _w19421_ ;
	wire _w19422_ ;
	wire _w19423_ ;
	wire _w19424_ ;
	wire _w19425_ ;
	wire _w19426_ ;
	wire _w19427_ ;
	wire _w19428_ ;
	wire _w19429_ ;
	wire _w19430_ ;
	wire _w19431_ ;
	wire _w19432_ ;
	wire _w19433_ ;
	wire _w19434_ ;
	wire _w19435_ ;
	wire _w19436_ ;
	wire _w19437_ ;
	wire _w19438_ ;
	wire _w19439_ ;
	wire _w19440_ ;
	wire _w19441_ ;
	wire _w19442_ ;
	wire _w19443_ ;
	wire _w19444_ ;
	wire _w19445_ ;
	wire _w19446_ ;
	wire _w19447_ ;
	wire _w19448_ ;
	wire _w19449_ ;
	wire _w19450_ ;
	wire _w19451_ ;
	wire _w19452_ ;
	wire _w19453_ ;
	wire _w19454_ ;
	wire _w19455_ ;
	wire _w19456_ ;
	wire _w19457_ ;
	wire _w19458_ ;
	wire _w19459_ ;
	wire _w19460_ ;
	wire _w19461_ ;
	wire _w19462_ ;
	wire _w19463_ ;
	wire _w19464_ ;
	wire _w19465_ ;
	wire _w19466_ ;
	wire _w19467_ ;
	wire _w19468_ ;
	wire _w19469_ ;
	wire _w19470_ ;
	wire _w19471_ ;
	wire _w19472_ ;
	wire _w19473_ ;
	wire _w19474_ ;
	wire _w19475_ ;
	wire _w19476_ ;
	wire _w19477_ ;
	wire _w19478_ ;
	wire _w19479_ ;
	wire _w19480_ ;
	wire _w19481_ ;
	wire _w19482_ ;
	wire _w19483_ ;
	wire _w19484_ ;
	wire _w19485_ ;
	wire _w19486_ ;
	wire _w19487_ ;
	wire _w19488_ ;
	wire _w19489_ ;
	wire _w19490_ ;
	wire _w19491_ ;
	wire _w19492_ ;
	wire _w19493_ ;
	wire _w19494_ ;
	wire _w19495_ ;
	wire _w19496_ ;
	wire _w19497_ ;
	wire _w19498_ ;
	wire _w19499_ ;
	wire _w19500_ ;
	wire _w19501_ ;
	wire _w19502_ ;
	wire _w19503_ ;
	wire _w19504_ ;
	wire _w19505_ ;
	wire _w19506_ ;
	wire _w19507_ ;
	wire _w19508_ ;
	wire _w19509_ ;
	wire _w19510_ ;
	wire _w19511_ ;
	wire _w19512_ ;
	wire _w19513_ ;
	wire _w19514_ ;
	wire _w19515_ ;
	wire _w19516_ ;
	wire _w19517_ ;
	wire _w19518_ ;
	wire _w19519_ ;
	wire _w19520_ ;
	wire _w19521_ ;
	wire _w19522_ ;
	wire _w19523_ ;
	wire _w19524_ ;
	wire _w19525_ ;
	wire _w19526_ ;
	wire _w19527_ ;
	wire _w19528_ ;
	wire _w19529_ ;
	wire _w19530_ ;
	wire _w19531_ ;
	wire _w19532_ ;
	wire _w19533_ ;
	wire _w19534_ ;
	wire _w19535_ ;
	wire _w19536_ ;
	wire _w19537_ ;
	wire _w19538_ ;
	wire _w19539_ ;
	wire _w19540_ ;
	wire _w19541_ ;
	wire _w19542_ ;
	wire _w19543_ ;
	wire _w19544_ ;
	wire _w19545_ ;
	wire _w19546_ ;
	wire _w19547_ ;
	wire _w19548_ ;
	wire _w19549_ ;
	wire _w19550_ ;
	wire _w19551_ ;
	wire _w19552_ ;
	wire _w19553_ ;
	wire _w19554_ ;
	wire _w19555_ ;
	wire _w19556_ ;
	wire _w19557_ ;
	wire _w19558_ ;
	wire _w19559_ ;
	wire _w19560_ ;
	wire _w19561_ ;
	wire _w19562_ ;
	wire _w19563_ ;
	wire _w19564_ ;
	wire _w19565_ ;
	wire _w19566_ ;
	wire _w19567_ ;
	wire _w19568_ ;
	wire _w19569_ ;
	wire _w19570_ ;
	wire _w19571_ ;
	wire _w19572_ ;
	wire _w19573_ ;
	wire _w19574_ ;
	wire _w19575_ ;
	wire _w19576_ ;
	wire _w19577_ ;
	wire _w19578_ ;
	wire _w19579_ ;
	wire _w19580_ ;
	wire _w19581_ ;
	wire _w19582_ ;
	wire _w19583_ ;
	wire _w19584_ ;
	wire _w19585_ ;
	wire _w19586_ ;
	wire _w19587_ ;
	wire _w19588_ ;
	wire _w19589_ ;
	wire _w19590_ ;
	wire _w19591_ ;
	wire _w19592_ ;
	wire _w19593_ ;
	wire _w19594_ ;
	wire _w19595_ ;
	wire _w19596_ ;
	wire _w19597_ ;
	wire _w19598_ ;
	wire _w19599_ ;
	wire _w19600_ ;
	wire _w19601_ ;
	wire _w19602_ ;
	wire _w19603_ ;
	wire _w19604_ ;
	wire _w19605_ ;
	wire _w19606_ ;
	wire _w19607_ ;
	wire _w19608_ ;
	wire _w19609_ ;
	wire _w19610_ ;
	wire _w19611_ ;
	wire _w19612_ ;
	wire _w19613_ ;
	wire _w19614_ ;
	wire _w19615_ ;
	wire _w19616_ ;
	wire _w19617_ ;
	wire _w19618_ ;
	wire _w19619_ ;
	wire _w19620_ ;
	wire _w19621_ ;
	wire _w19622_ ;
	wire _w19623_ ;
	wire _w19624_ ;
	wire _w19625_ ;
	wire _w19626_ ;
	wire _w19627_ ;
	wire _w19628_ ;
	wire _w19629_ ;
	wire _w19630_ ;
	wire _w19631_ ;
	wire _w19632_ ;
	wire _w19633_ ;
	wire _w19634_ ;
	wire _w19635_ ;
	wire _w19636_ ;
	wire _w19637_ ;
	wire _w19638_ ;
	wire _w19639_ ;
	wire _w19640_ ;
	wire _w19641_ ;
	wire _w19642_ ;
	wire _w19643_ ;
	wire _w19644_ ;
	wire _w19645_ ;
	wire _w19646_ ;
	wire _w19647_ ;
	wire _w19648_ ;
	wire _w19649_ ;
	wire _w19650_ ;
	wire _w19651_ ;
	wire _w19652_ ;
	wire _w19653_ ;
	wire _w19654_ ;
	wire _w19655_ ;
	wire _w19656_ ;
	wire _w19657_ ;
	wire _w19658_ ;
	wire _w19659_ ;
	wire _w19660_ ;
	wire _w19661_ ;
	wire _w19662_ ;
	wire _w19663_ ;
	wire _w19664_ ;
	wire _w19665_ ;
	wire _w19666_ ;
	wire _w19667_ ;
	wire _w19668_ ;
	wire _w19669_ ;
	wire _w19670_ ;
	wire _w19671_ ;
	wire _w19672_ ;
	wire _w19673_ ;
	wire _w19674_ ;
	wire _w19675_ ;
	wire _w19676_ ;
	wire _w19677_ ;
	wire _w19678_ ;
	wire _w19679_ ;
	wire _w19680_ ;
	wire _w19681_ ;
	wire _w19682_ ;
	wire _w19683_ ;
	wire _w19684_ ;
	wire _w19685_ ;
	wire _w19686_ ;
	wire _w19687_ ;
	wire _w19688_ ;
	wire _w19689_ ;
	wire _w19690_ ;
	wire _w19691_ ;
	wire _w19692_ ;
	wire _w19693_ ;
	wire _w19694_ ;
	wire _w19695_ ;
	wire _w19696_ ;
	wire _w19697_ ;
	wire _w19698_ ;
	wire _w19699_ ;
	wire _w19700_ ;
	wire _w19701_ ;
	wire _w19702_ ;
	wire _w19703_ ;
	wire _w19704_ ;
	wire _w19705_ ;
	wire _w19706_ ;
	wire _w19707_ ;
	wire _w19708_ ;
	wire _w19709_ ;
	wire _w19710_ ;
	wire _w19711_ ;
	wire _w19712_ ;
	wire _w19713_ ;
	wire _w19714_ ;
	wire _w19715_ ;
	wire _w19716_ ;
	wire _w19717_ ;
	wire _w19718_ ;
	wire _w19719_ ;
	wire _w19720_ ;
	wire _w19721_ ;
	wire _w19722_ ;
	wire _w19723_ ;
	wire _w19724_ ;
	wire _w19725_ ;
	wire _w19726_ ;
	wire _w19727_ ;
	wire _w19728_ ;
	wire _w19729_ ;
	wire _w19730_ ;
	wire _w19731_ ;
	wire _w19732_ ;
	wire _w19733_ ;
	wire _w19734_ ;
	wire _w19735_ ;
	wire _w19736_ ;
	wire _w19737_ ;
	wire _w19738_ ;
	wire _w19739_ ;
	wire _w19740_ ;
	wire _w19741_ ;
	wire _w19742_ ;
	wire _w19743_ ;
	wire _w19744_ ;
	wire _w19745_ ;
	wire _w19746_ ;
	wire _w19747_ ;
	wire _w19748_ ;
	wire _w19749_ ;
	wire _w19750_ ;
	wire _w19751_ ;
	wire _w19752_ ;
	wire _w19753_ ;
	wire _w19754_ ;
	wire _w19755_ ;
	wire _w19756_ ;
	wire _w19757_ ;
	wire _w19758_ ;
	wire _w19759_ ;
	wire _w19760_ ;
	wire _w19761_ ;
	wire _w19762_ ;
	wire _w19763_ ;
	wire _w19764_ ;
	wire _w19765_ ;
	wire _w19766_ ;
	wire _w19767_ ;
	wire _w19768_ ;
	wire _w19769_ ;
	wire _w19770_ ;
	wire _w19771_ ;
	wire _w19772_ ;
	wire _w19773_ ;
	wire _w19774_ ;
	wire _w19775_ ;
	wire _w19776_ ;
	wire _w19777_ ;
	wire _w19778_ ;
	wire _w19779_ ;
	wire _w19780_ ;
	wire _w19781_ ;
	wire _w19782_ ;
	wire _w19783_ ;
	wire _w19784_ ;
	wire _w19785_ ;
	wire _w19786_ ;
	wire _w19787_ ;
	wire _w19788_ ;
	wire _w19789_ ;
	wire _w19790_ ;
	wire _w19791_ ;
	wire _w19792_ ;
	wire _w19793_ ;
	wire _w19794_ ;
	wire _w19795_ ;
	wire _w19796_ ;
	wire _w19797_ ;
	wire _w19798_ ;
	wire _w19799_ ;
	wire _w19800_ ;
	wire _w19801_ ;
	wire _w19802_ ;
	wire _w19803_ ;
	wire _w19804_ ;
	wire _w19805_ ;
	wire _w19806_ ;
	wire _w19807_ ;
	wire _w19808_ ;
	wire _w19809_ ;
	wire _w19810_ ;
	wire _w19811_ ;
	wire _w19812_ ;
	wire _w19813_ ;
	wire _w19814_ ;
	wire _w19815_ ;
	wire _w19816_ ;
	wire _w19817_ ;
	wire _w19818_ ;
	wire _w19819_ ;
	wire _w19820_ ;
	wire _w19821_ ;
	wire _w19822_ ;
	wire _w19823_ ;
	wire _w19824_ ;
	wire _w19825_ ;
	wire _w19826_ ;
	wire _w19827_ ;
	wire _w19828_ ;
	wire _w19829_ ;
	wire _w19830_ ;
	wire _w19831_ ;
	wire _w19832_ ;
	wire _w19833_ ;
	wire _w19834_ ;
	wire _w19835_ ;
	wire _w19836_ ;
	wire _w19837_ ;
	wire _w19838_ ;
	wire _w19839_ ;
	wire _w19840_ ;
	wire _w19841_ ;
	wire _w19842_ ;
	wire _w19843_ ;
	wire _w19844_ ;
	wire _w19845_ ;
	wire _w19846_ ;
	wire _w19847_ ;
	wire _w19848_ ;
	wire _w19849_ ;
	wire _w19850_ ;
	wire _w19851_ ;
	wire _w19852_ ;
	wire _w19853_ ;
	wire _w19854_ ;
	wire _w19855_ ;
	wire _w19856_ ;
	wire _w19857_ ;
	wire _w19858_ ;
	wire _w19859_ ;
	wire _w19860_ ;
	wire _w19861_ ;
	wire _w19862_ ;
	wire _w19863_ ;
	wire _w19864_ ;
	wire _w19865_ ;
	wire _w19866_ ;
	wire _w19867_ ;
	wire _w19868_ ;
	wire _w19869_ ;
	wire _w19870_ ;
	wire _w19871_ ;
	wire _w19872_ ;
	wire _w19873_ ;
	wire _w19874_ ;
	wire _w19875_ ;
	wire _w19876_ ;
	wire _w19877_ ;
	wire _w19878_ ;
	wire _w19879_ ;
	wire _w19880_ ;
	wire _w19881_ ;
	wire _w19882_ ;
	wire _w19883_ ;
	wire _w19884_ ;
	wire _w19885_ ;
	wire _w19886_ ;
	wire _w19887_ ;
	wire _w19888_ ;
	wire _w19889_ ;
	wire _w19890_ ;
	wire _w19891_ ;
	wire _w19892_ ;
	wire _w19893_ ;
	wire _w19894_ ;
	wire _w19895_ ;
	wire _w19896_ ;
	wire _w19897_ ;
	wire _w19898_ ;
	wire _w19899_ ;
	wire _w19900_ ;
	wire _w19901_ ;
	wire _w19902_ ;
	wire _w19903_ ;
	wire _w19904_ ;
	wire _w19905_ ;
	wire _w19906_ ;
	wire _w19907_ ;
	wire _w19908_ ;
	wire _w19909_ ;
	wire _w19910_ ;
	wire _w19911_ ;
	wire _w19912_ ;
	wire _w19913_ ;
	wire _w19914_ ;
	wire _w19915_ ;
	wire _w19916_ ;
	wire _w19917_ ;
	wire _w19918_ ;
	wire _w19919_ ;
	wire _w19920_ ;
	wire _w19921_ ;
	wire _w19922_ ;
	wire _w19923_ ;
	wire _w19924_ ;
	wire _w19925_ ;
	wire _w19926_ ;
	wire _w19927_ ;
	wire _w19928_ ;
	wire _w19929_ ;
	wire _w19930_ ;
	wire _w19931_ ;
	wire _w19932_ ;
	wire _w19933_ ;
	wire _w19934_ ;
	wire _w19935_ ;
	wire _w19936_ ;
	wire _w19937_ ;
	wire _w19938_ ;
	wire _w19939_ ;
	wire _w19940_ ;
	wire _w19941_ ;
	wire _w19942_ ;
	wire _w19943_ ;
	wire _w19944_ ;
	wire _w19945_ ;
	wire _w19946_ ;
	wire _w19947_ ;
	wire _w19948_ ;
	wire _w19949_ ;
	wire _w19950_ ;
	wire _w19951_ ;
	wire _w19952_ ;
	wire _w19953_ ;
	wire _w19954_ ;
	wire _w19955_ ;
	wire _w19956_ ;
	wire _w19957_ ;
	wire _w19958_ ;
	wire _w19959_ ;
	wire _w19960_ ;
	wire _w19961_ ;
	wire _w19962_ ;
	wire _w19963_ ;
	wire _w19964_ ;
	wire _w19965_ ;
	wire _w19966_ ;
	wire _w19967_ ;
	wire _w19968_ ;
	wire _w19969_ ;
	wire _w19970_ ;
	wire _w19971_ ;
	wire _w19972_ ;
	wire _w19973_ ;
	wire _w19974_ ;
	wire _w19975_ ;
	wire _w19976_ ;
	wire _w19977_ ;
	wire _w19978_ ;
	wire _w19979_ ;
	wire _w19980_ ;
	wire _w19981_ ;
	wire _w19982_ ;
	wire _w19983_ ;
	wire _w19984_ ;
	wire _w19985_ ;
	wire _w19986_ ;
	wire _w19987_ ;
	wire _w19988_ ;
	wire _w19989_ ;
	wire _w19990_ ;
	wire _w19991_ ;
	wire _w19992_ ;
	wire _w19993_ ;
	wire _w19994_ ;
	wire _w19995_ ;
	wire _w19996_ ;
	wire _w19997_ ;
	wire _w19998_ ;
	wire _w19999_ ;
	wire _w20000_ ;
	wire _w20001_ ;
	wire _w20002_ ;
	wire _w20003_ ;
	wire _w20004_ ;
	wire _w20005_ ;
	wire _w20006_ ;
	wire _w20007_ ;
	wire _w20008_ ;
	wire _w20009_ ;
	wire _w20010_ ;
	wire _w20011_ ;
	wire _w20012_ ;
	wire _w20013_ ;
	wire _w20014_ ;
	wire _w20015_ ;
	wire _w20016_ ;
	wire _w20017_ ;
	wire _w20018_ ;
	wire _w20019_ ;
	wire _w20020_ ;
	wire _w20021_ ;
	wire _w20022_ ;
	wire _w20023_ ;
	wire _w20024_ ;
	wire _w20025_ ;
	wire _w20026_ ;
	wire _w20027_ ;
	wire _w20028_ ;
	wire _w20029_ ;
	wire _w20030_ ;
	wire _w20031_ ;
	wire _w20032_ ;
	wire _w20033_ ;
	wire _w20034_ ;
	wire _w20035_ ;
	wire _w20036_ ;
	wire _w20037_ ;
	wire _w20038_ ;
	wire _w20039_ ;
	wire _w20040_ ;
	wire _w20041_ ;
	wire _w20042_ ;
	wire _w20043_ ;
	wire _w20044_ ;
	wire _w20045_ ;
	wire _w20046_ ;
	wire _w20047_ ;
	wire _w20048_ ;
	wire _w20049_ ;
	wire _w20050_ ;
	wire _w20051_ ;
	wire _w20052_ ;
	wire _w20053_ ;
	wire _w20054_ ;
	wire _w20055_ ;
	wire _w20056_ ;
	wire _w20057_ ;
	wire _w20058_ ;
	wire _w20059_ ;
	wire _w20060_ ;
	wire _w20061_ ;
	wire _w20062_ ;
	wire _w20063_ ;
	wire _w20064_ ;
	wire _w20065_ ;
	wire _w20066_ ;
	wire _w20067_ ;
	wire _w20068_ ;
	wire _w20069_ ;
	wire _w20070_ ;
	wire _w20071_ ;
	wire _w20072_ ;
	wire _w20073_ ;
	wire _w20074_ ;
	wire _w20075_ ;
	wire _w20076_ ;
	wire _w20077_ ;
	wire _w20078_ ;
	wire _w20079_ ;
	wire _w20080_ ;
	wire _w20081_ ;
	wire _w20082_ ;
	wire _w20083_ ;
	wire _w20084_ ;
	wire _w20085_ ;
	wire _w20086_ ;
	wire _w20087_ ;
	wire _w20088_ ;
	wire _w20089_ ;
	wire _w20090_ ;
	wire _w20091_ ;
	wire _w20092_ ;
	wire _w20093_ ;
	wire _w20094_ ;
	wire _w20095_ ;
	wire _w20096_ ;
	wire _w20097_ ;
	wire _w20098_ ;
	wire _w20099_ ;
	wire _w20100_ ;
	wire _w20101_ ;
	wire _w20102_ ;
	wire _w20103_ ;
	wire _w20104_ ;
	wire _w20105_ ;
	wire _w20106_ ;
	wire _w20107_ ;
	wire _w20108_ ;
	wire _w20109_ ;
	wire _w20110_ ;
	wire _w20111_ ;
	wire _w20112_ ;
	wire _w20113_ ;
	wire _w20114_ ;
	wire _w20115_ ;
	wire _w20116_ ;
	wire _w20117_ ;
	wire _w20118_ ;
	wire _w20119_ ;
	wire _w20120_ ;
	wire _w20121_ ;
	wire _w20122_ ;
	wire _w20123_ ;
	wire _w20124_ ;
	wire _w20125_ ;
	wire _w20126_ ;
	wire _w20127_ ;
	wire _w20128_ ;
	wire _w20129_ ;
	wire _w20130_ ;
	wire _w20131_ ;
	wire _w20132_ ;
	wire _w20133_ ;
	wire _w20134_ ;
	wire _w20135_ ;
	wire _w20136_ ;
	wire _w20137_ ;
	wire _w20138_ ;
	wire _w20139_ ;
	wire _w20140_ ;
	wire _w20141_ ;
	wire _w20142_ ;
	wire _w20143_ ;
	wire _w20144_ ;
	wire _w20145_ ;
	wire _w20146_ ;
	wire _w20147_ ;
	wire _w20148_ ;
	wire _w20149_ ;
	wire _w20150_ ;
	wire _w20151_ ;
	wire _w20152_ ;
	wire _w20153_ ;
	wire _w20154_ ;
	wire _w20155_ ;
	wire _w20156_ ;
	wire _w20157_ ;
	wire _w20158_ ;
	wire _w20159_ ;
	wire _w20160_ ;
	wire _w20161_ ;
	wire _w20162_ ;
	wire _w20163_ ;
	wire _w20164_ ;
	wire _w20165_ ;
	wire _w20166_ ;
	wire _w20167_ ;
	wire _w20168_ ;
	wire _w20169_ ;
	wire _w20170_ ;
	wire _w20171_ ;
	wire _w20172_ ;
	wire _w20173_ ;
	wire _w20174_ ;
	wire _w20175_ ;
	wire _w20176_ ;
	wire _w20177_ ;
	wire _w20178_ ;
	wire _w20179_ ;
	wire _w20180_ ;
	wire _w20181_ ;
	wire _w20182_ ;
	wire _w20183_ ;
	wire _w20184_ ;
	wire _w20185_ ;
	wire _w20186_ ;
	wire _w20187_ ;
	wire _w20188_ ;
	wire _w20189_ ;
	wire _w20190_ ;
	wire _w20191_ ;
	wire _w20192_ ;
	wire _w20193_ ;
	wire _w20194_ ;
	wire _w20195_ ;
	wire _w20196_ ;
	wire _w20197_ ;
	wire _w20198_ ;
	wire _w20199_ ;
	wire _w20200_ ;
	wire _w20201_ ;
	wire _w20202_ ;
	wire _w20203_ ;
	wire _w20204_ ;
	wire _w20205_ ;
	wire _w20206_ ;
	wire _w20207_ ;
	wire _w20208_ ;
	wire _w20209_ ;
	wire _w20210_ ;
	wire _w20211_ ;
	wire _w20212_ ;
	wire _w20213_ ;
	wire _w20214_ ;
	wire _w20215_ ;
	wire _w20216_ ;
	wire _w20217_ ;
	wire _w20218_ ;
	wire _w20219_ ;
	wire _w20220_ ;
	wire _w20221_ ;
	wire _w20222_ ;
	wire _w20223_ ;
	wire _w20224_ ;
	wire _w20225_ ;
	wire _w20226_ ;
	wire _w20227_ ;
	wire _w20228_ ;
	wire _w20229_ ;
	wire _w20230_ ;
	wire _w20231_ ;
	wire _w20232_ ;
	wire _w20233_ ;
	wire _w20234_ ;
	wire _w20235_ ;
	wire _w20236_ ;
	wire _w20237_ ;
	wire _w20238_ ;
	wire _w20239_ ;
	wire _w20240_ ;
	wire _w20241_ ;
	wire _w20242_ ;
	wire _w20243_ ;
	wire _w20244_ ;
	wire _w20245_ ;
	wire _w20246_ ;
	wire _w20247_ ;
	wire _w20248_ ;
	wire _w20249_ ;
	wire _w20250_ ;
	wire _w20251_ ;
	wire _w20252_ ;
	wire _w20253_ ;
	wire _w20254_ ;
	wire _w20255_ ;
	wire _w20256_ ;
	wire _w20257_ ;
	wire _w20258_ ;
	wire _w20259_ ;
	wire _w20260_ ;
	wire _w20261_ ;
	wire _w20262_ ;
	wire _w20263_ ;
	wire _w20264_ ;
	wire _w20265_ ;
	wire _w20266_ ;
	wire _w20267_ ;
	wire _w20268_ ;
	wire _w20269_ ;
	wire _w20270_ ;
	wire _w20271_ ;
	wire _w20272_ ;
	wire _w20273_ ;
	wire _w20274_ ;
	wire _w20275_ ;
	wire _w20276_ ;
	wire _w20277_ ;
	wire _w20278_ ;
	wire _w20279_ ;
	wire _w20280_ ;
	wire _w20281_ ;
	wire _w20282_ ;
	wire _w20283_ ;
	wire _w20284_ ;
	wire _w20285_ ;
	wire _w20286_ ;
	wire _w20287_ ;
	wire _w20288_ ;
	wire _w20289_ ;
	wire _w20290_ ;
	wire _w20291_ ;
	wire _w20292_ ;
	wire _w20293_ ;
	wire _w20294_ ;
	wire _w20295_ ;
	wire _w20296_ ;
	wire _w20297_ ;
	wire _w20298_ ;
	wire _w20299_ ;
	wire _w20300_ ;
	wire _w20301_ ;
	wire _w20302_ ;
	wire _w20303_ ;
	wire _w20304_ ;
	wire _w20305_ ;
	wire _w20306_ ;
	wire _w20307_ ;
	wire _w20308_ ;
	wire _w20309_ ;
	wire _w20310_ ;
	wire _w20311_ ;
	wire _w20312_ ;
	wire _w20313_ ;
	wire _w20314_ ;
	wire _w20315_ ;
	wire _w20316_ ;
	wire _w20317_ ;
	wire _w20318_ ;
	wire _w20319_ ;
	wire _w20320_ ;
	wire _w20321_ ;
	wire _w20322_ ;
	wire _w20323_ ;
	wire _w20324_ ;
	wire _w20325_ ;
	wire _w20326_ ;
	wire _w20327_ ;
	wire _w20328_ ;
	wire _w20329_ ;
	wire _w20330_ ;
	wire _w20331_ ;
	wire _w20332_ ;
	wire _w20333_ ;
	wire _w20334_ ;
	wire _w20335_ ;
	wire _w20336_ ;
	wire _w20337_ ;
	wire _w20338_ ;
	wire _w20339_ ;
	wire _w20340_ ;
	wire _w20341_ ;
	wire _w20342_ ;
	wire _w20343_ ;
	wire _w20344_ ;
	wire _w20345_ ;
	wire _w20346_ ;
	wire _w20347_ ;
	wire _w20348_ ;
	wire _w20349_ ;
	wire _w20350_ ;
	wire _w20351_ ;
	wire _w20352_ ;
	wire _w20353_ ;
	wire _w20354_ ;
	wire _w20355_ ;
	wire _w20356_ ;
	wire _w20357_ ;
	wire _w20358_ ;
	wire _w20359_ ;
	wire _w20360_ ;
	wire _w20361_ ;
	wire _w20362_ ;
	wire _w20363_ ;
	wire _w20364_ ;
	wire _w20365_ ;
	wire _w20366_ ;
	wire _w20367_ ;
	wire _w20368_ ;
	wire _w20369_ ;
	wire _w20370_ ;
	wire _w20371_ ;
	wire _w20372_ ;
	wire _w20373_ ;
	wire _w20374_ ;
	wire _w20375_ ;
	wire _w20376_ ;
	wire _w20377_ ;
	wire _w20378_ ;
	wire _w20379_ ;
	wire _w20380_ ;
	wire _w20381_ ;
	wire _w20382_ ;
	wire _w20383_ ;
	wire _w20384_ ;
	wire _w20385_ ;
	wire _w20386_ ;
	wire _w20387_ ;
	wire _w20388_ ;
	wire _w20389_ ;
	wire _w20390_ ;
	wire _w20391_ ;
	wire _w20392_ ;
	wire _w20393_ ;
	wire _w20394_ ;
	wire _w20395_ ;
	wire _w20396_ ;
	wire _w20397_ ;
	wire _w20398_ ;
	wire _w20399_ ;
	wire _w20400_ ;
	wire _w20401_ ;
	wire _w20402_ ;
	wire _w20403_ ;
	wire _w20404_ ;
	wire _w20405_ ;
	wire _w20406_ ;
	wire _w20407_ ;
	wire _w20408_ ;
	wire _w20409_ ;
	wire _w20410_ ;
	wire _w20411_ ;
	wire _w20412_ ;
	wire _w20413_ ;
	wire _w20414_ ;
	wire _w20415_ ;
	wire _w20416_ ;
	wire _w20417_ ;
	wire _w20418_ ;
	wire _w20419_ ;
	wire _w20420_ ;
	wire _w20421_ ;
	wire _w20422_ ;
	wire _w20423_ ;
	wire _w20424_ ;
	wire _w20425_ ;
	wire _w20426_ ;
	wire _w20427_ ;
	wire _w20428_ ;
	wire _w20429_ ;
	wire _w20430_ ;
	wire _w20431_ ;
	wire _w20432_ ;
	wire _w20433_ ;
	wire _w20434_ ;
	wire _w20435_ ;
	wire _w20436_ ;
	wire _w20437_ ;
	wire _w20438_ ;
	wire _w20439_ ;
	wire _w20440_ ;
	wire _w20441_ ;
	wire _w20442_ ;
	wire _w20443_ ;
	wire _w20444_ ;
	wire _w20445_ ;
	wire _w20446_ ;
	wire _w20447_ ;
	wire _w20448_ ;
	wire _w20449_ ;
	wire _w20450_ ;
	wire _w20451_ ;
	wire _w20452_ ;
	wire _w20453_ ;
	wire _w20454_ ;
	wire _w20455_ ;
	wire _w20456_ ;
	wire _w20457_ ;
	wire _w20458_ ;
	wire _w20459_ ;
	wire _w20460_ ;
	wire _w20461_ ;
	wire _w20462_ ;
	wire _w20463_ ;
	wire _w20464_ ;
	wire _w20465_ ;
	wire _w20466_ ;
	wire _w20467_ ;
	wire _w20468_ ;
	wire _w20469_ ;
	wire _w20470_ ;
	wire _w20471_ ;
	wire _w20472_ ;
	wire _w20473_ ;
	wire _w20474_ ;
	wire _w20475_ ;
	wire _w20476_ ;
	wire _w20477_ ;
	wire _w20478_ ;
	wire _w20479_ ;
	wire _w20480_ ;
	wire _w20481_ ;
	wire _w20482_ ;
	wire _w20483_ ;
	wire _w20484_ ;
	wire _w20485_ ;
	wire _w20486_ ;
	wire _w20487_ ;
	wire _w20488_ ;
	wire _w20489_ ;
	wire _w20490_ ;
	wire _w20491_ ;
	wire _w20492_ ;
	wire _w20493_ ;
	wire _w20494_ ;
	wire _w20495_ ;
	wire _w20496_ ;
	wire _w20497_ ;
	wire _w20498_ ;
	wire _w20499_ ;
	wire _w20500_ ;
	wire _w20501_ ;
	wire _w20502_ ;
	wire _w20503_ ;
	wire _w20504_ ;
	wire _w20505_ ;
	wire _w20506_ ;
	wire _w20507_ ;
	wire _w20508_ ;
	wire _w20509_ ;
	wire _w20510_ ;
	wire _w20511_ ;
	wire _w20512_ ;
	wire _w20513_ ;
	wire _w20514_ ;
	wire _w20515_ ;
	wire _w20516_ ;
	wire _w20517_ ;
	wire _w20518_ ;
	wire _w20519_ ;
	wire _w20520_ ;
	wire _w20521_ ;
	wire _w20522_ ;
	wire _w20523_ ;
	wire _w20524_ ;
	wire _w20525_ ;
	wire _w20526_ ;
	wire _w20527_ ;
	wire _w20528_ ;
	wire _w20529_ ;
	wire _w20530_ ;
	wire _w20531_ ;
	wire _w20532_ ;
	wire _w20533_ ;
	wire _w20534_ ;
	wire _w20535_ ;
	wire _w20536_ ;
	wire _w20537_ ;
	wire _w20538_ ;
	wire _w20539_ ;
	wire _w20540_ ;
	wire _w20541_ ;
	wire _w20542_ ;
	wire _w20543_ ;
	wire _w20544_ ;
	wire _w20545_ ;
	wire _w20546_ ;
	wire _w20547_ ;
	wire _w20548_ ;
	wire _w20549_ ;
	wire _w20550_ ;
	wire _w20551_ ;
	wire _w20552_ ;
	wire _w20553_ ;
	wire _w20554_ ;
	wire _w20555_ ;
	wire _w20556_ ;
	wire _w20557_ ;
	wire _w20558_ ;
	wire _w20559_ ;
	wire _w20560_ ;
	wire _w20561_ ;
	wire _w20562_ ;
	wire _w20563_ ;
	wire _w20564_ ;
	wire _w20565_ ;
	wire _w20566_ ;
	wire _w20567_ ;
	wire _w20568_ ;
	wire _w20569_ ;
	wire _w20570_ ;
	wire _w20571_ ;
	wire _w20572_ ;
	wire _w20573_ ;
	wire _w20574_ ;
	wire _w20575_ ;
	wire _w20576_ ;
	wire _w20577_ ;
	wire _w20578_ ;
	wire _w20579_ ;
	wire _w20580_ ;
	wire _w20581_ ;
	wire _w20582_ ;
	wire _w20583_ ;
	wire _w20584_ ;
	wire _w20585_ ;
	wire _w20586_ ;
	wire _w20587_ ;
	wire _w20588_ ;
	wire _w20589_ ;
	wire _w20590_ ;
	wire _w20591_ ;
	wire _w20592_ ;
	wire _w20593_ ;
	wire _w20594_ ;
	wire _w20595_ ;
	wire _w20596_ ;
	wire _w20597_ ;
	wire _w20598_ ;
	wire _w20599_ ;
	wire _w20600_ ;
	wire _w20601_ ;
	wire _w20602_ ;
	wire _w20603_ ;
	wire _w20604_ ;
	wire _w20605_ ;
	wire _w20606_ ;
	wire _w20607_ ;
	wire _w20608_ ;
	wire _w20609_ ;
	wire _w20610_ ;
	wire _w20611_ ;
	wire _w20612_ ;
	wire _w20613_ ;
	wire _w20614_ ;
	wire _w20615_ ;
	wire _w20616_ ;
	wire _w20617_ ;
	wire _w20618_ ;
	wire _w20619_ ;
	wire _w20620_ ;
	wire _w20621_ ;
	wire _w20622_ ;
	wire _w20623_ ;
	wire _w20624_ ;
	wire _w20625_ ;
	wire _w20626_ ;
	wire _w20627_ ;
	wire _w20628_ ;
	wire _w20629_ ;
	wire _w20630_ ;
	wire _w20631_ ;
	wire _w20632_ ;
	wire _w20633_ ;
	wire _w20634_ ;
	wire _w20635_ ;
	wire _w20636_ ;
	wire _w20637_ ;
	wire _w20638_ ;
	wire _w20639_ ;
	wire _w20640_ ;
	wire _w20641_ ;
	wire _w20642_ ;
	wire _w20643_ ;
	wire _w20644_ ;
	wire _w20645_ ;
	wire _w20646_ ;
	wire _w20647_ ;
	wire _w20648_ ;
	wire _w20649_ ;
	wire _w20650_ ;
	wire _w20651_ ;
	wire _w20652_ ;
	wire _w20653_ ;
	wire _w20654_ ;
	wire _w20655_ ;
	wire _w20656_ ;
	wire _w20657_ ;
	wire _w20658_ ;
	wire _w20659_ ;
	wire _w20660_ ;
	wire _w20661_ ;
	wire _w20662_ ;
	wire _w20663_ ;
	wire _w20664_ ;
	wire _w20665_ ;
	wire _w20666_ ;
	wire _w20667_ ;
	wire _w20668_ ;
	wire _w20669_ ;
	wire _w20670_ ;
	wire _w20671_ ;
	wire _w20672_ ;
	wire _w20673_ ;
	wire _w20674_ ;
	wire _w20675_ ;
	wire _w20676_ ;
	wire _w20677_ ;
	wire _w20678_ ;
	wire _w20679_ ;
	wire _w20680_ ;
	wire _w20681_ ;
	wire _w20682_ ;
	wire _w20683_ ;
	wire _w20684_ ;
	wire _w20685_ ;
	wire _w20686_ ;
	wire _w20687_ ;
	wire _w20688_ ;
	wire _w20689_ ;
	wire _w20690_ ;
	wire _w20691_ ;
	wire _w20692_ ;
	wire _w20693_ ;
	wire _w20694_ ;
	wire _w20695_ ;
	wire _w20696_ ;
	wire _w20697_ ;
	wire _w20698_ ;
	wire _w20699_ ;
	wire _w20700_ ;
	wire _w20701_ ;
	wire _w20702_ ;
	wire _w20703_ ;
	wire _w20704_ ;
	wire _w20705_ ;
	wire _w20706_ ;
	wire _w20707_ ;
	wire _w20708_ ;
	wire _w20709_ ;
	wire _w20710_ ;
	wire _w20711_ ;
	wire _w20712_ ;
	wire _w20713_ ;
	wire _w20714_ ;
	wire _w20715_ ;
	wire _w20716_ ;
	wire _w20717_ ;
	wire _w20718_ ;
	wire _w20719_ ;
	wire _w20720_ ;
	wire _w20721_ ;
	wire _w20722_ ;
	wire _w20723_ ;
	wire _w20724_ ;
	wire _w20725_ ;
	wire _w20726_ ;
	wire _w20727_ ;
	wire _w20728_ ;
	wire _w20729_ ;
	wire _w20730_ ;
	wire _w20731_ ;
	wire _w20732_ ;
	wire _w20733_ ;
	wire _w20734_ ;
	wire _w20735_ ;
	wire _w20736_ ;
	wire _w20737_ ;
	wire _w20738_ ;
	wire _w20739_ ;
	wire _w20740_ ;
	wire _w20741_ ;
	wire _w20742_ ;
	wire _w20743_ ;
	wire _w20744_ ;
	wire _w20745_ ;
	wire _w20746_ ;
	wire _w20747_ ;
	wire _w20748_ ;
	wire _w20749_ ;
	wire _w20750_ ;
	wire _w20751_ ;
	wire _w20752_ ;
	wire _w20753_ ;
	wire _w20754_ ;
	wire _w20755_ ;
	wire _w20756_ ;
	wire _w20757_ ;
	wire _w20758_ ;
	wire _w20759_ ;
	wire _w20760_ ;
	wire _w20761_ ;
	wire _w20762_ ;
	wire _w20763_ ;
	wire _w20764_ ;
	wire _w20765_ ;
	wire _w20766_ ;
	wire _w20767_ ;
	wire _w20768_ ;
	wire _w20769_ ;
	wire _w20770_ ;
	wire _w20771_ ;
	wire _w20772_ ;
	wire _w20773_ ;
	wire _w20774_ ;
	wire _w20775_ ;
	wire _w20776_ ;
	wire _w20777_ ;
	wire _w20778_ ;
	wire _w20779_ ;
	wire _w20780_ ;
	wire _w20781_ ;
	wire _w20782_ ;
	wire _w20783_ ;
	wire _w20784_ ;
	wire _w20785_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		_w460_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w10514_
	);
	LUT4 #(
		.INIT('h0001)
	) name2 (
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w10515_
	);
	LUT4 #(
		.INIT('h0001)
	) name3 (
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		_w10516_
	);
	LUT4 #(
		.INIT('h0001)
	) name4 (
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w10517_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w10518_
	);
	LUT4 #(
		.INIT('h8000)
	) name6 (
		_w10515_,
		_w10516_,
		_w10517_,
		_w10518_,
		_w10519_
	);
	LUT4 #(
		.INIT('h0002)
	) name7 (
		\rxethmac1_crcrx_Crc_reg[26]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[27]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[28]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[2]/NET0131 ,
		_w10520_
	);
	LUT4 #(
		.INIT('h1000)
	) name8 (
		\rxethmac1_crcrx_Crc_reg[22]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[23]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[24]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[25]/NET0131 ,
		_w10521_
	);
	LUT4 #(
		.INIT('h0020)
	) name9 (
		\rxethmac1_crcrx_Crc_reg[6]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[7]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[8]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[9]/NET0131 ,
		_w10522_
	);
	LUT4 #(
		.INIT('h8000)
	) name10 (
		\rxethmac1_crcrx_Crc_reg[30]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[3]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[4]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[5]/NET0131 ,
		_w10523_
	);
	LUT4 #(
		.INIT('h8000)
	) name11 (
		_w10520_,
		_w10521_,
		_w10522_,
		_w10523_,
		_w10524_
	);
	LUT4 #(
		.INIT('h0800)
	) name12 (
		\rxethmac1_crcrx_Crc_reg[11]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[12]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[13]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[14]/NET0131 ,
		_w10525_
	);
	LUT4 #(
		.INIT('h0800)
	) name13 (
		\rxethmac1_crcrx_Crc_reg[0]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[10]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[29]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[31]/NET0131 ,
		_w10526_
	);
	LUT4 #(
		.INIT('h0004)
	) name14 (
		\rxethmac1_crcrx_Crc_reg[19]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[1]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[20]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[21]/NET0131 ,
		_w10527_
	);
	LUT4 #(
		.INIT('h0200)
	) name15 (
		\rxethmac1_crcrx_Crc_reg[15]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[16]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[17]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[18]/NET0131 ,
		_w10528_
	);
	LUT4 #(
		.INIT('h8000)
	) name16 (
		_w10525_,
		_w10526_,
		_w10527_,
		_w10528_,
		_w10529_
	);
	LUT4 #(
		.INIT('h0777)
	) name17 (
		_w10514_,
		_w10519_,
		_w10524_,
		_w10529_,
		_w10530_
	);
	LUT3 #(
		.INIT('h0e)
	) name18 (
		\macstatus1_LatchedCrcError_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w10531_
	);
	LUT3 #(
		.INIT('hd0)
	) name19 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10530_,
		_w10531_,
		_w10532_
	);
	LUT4 #(
		.INIT('h8000)
	) name20 (
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		_w10515_,
		_w10516_,
		_w10517_,
		_w10533_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10534_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w10535_
	);
	LUT4 #(
		.INIT('h0400)
	) name23 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10536_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		\rxethmac1_crcrx_Crc_reg[27]/NET0131 ,
		_w10536_,
		_w10537_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		wb_rst_i_pad,
		_w10538_
	);
	LUT3 #(
		.INIT('h02)
	) name26 (
		\rxethmac1_CrcHash_reg[1]/P0001 ,
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		wb_rst_i_pad,
		_w10539_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		_w10536_,
		_w10538_,
		_w10540_
	);
	LUT4 #(
		.INIT('h7270)
	) name28 (
		_w10533_,
		_w10537_,
		_w10539_,
		_w10540_,
		_w10541_
	);
	LUT4 #(
		.INIT('hfe00)
	) name29 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131 ,
		_w10542_
	);
	LUT4 #(
		.INIT('h0001)
	) name30 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131 ,
		_w10543_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		\rxethmac1_crcrx_Crc_reg[27]/NET0131 ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w10544_
	);
	LUT4 #(
		.INIT('h02ff)
	) name32 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		_w10542_,
		_w10543_,
		_w10544_,
		_w10545_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		_w10546_
	);
	LUT4 #(
		.INIT('hf531)
	) name34 (
		\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 ,
		\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		_w10547_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		_w10546_,
		_w10547_,
		_w10548_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name36 (
		\ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		_w10549_
	);
	LUT4 #(
		.INIT('h8caf)
	) name37 (
		\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		_w10550_
	);
	LUT4 #(
		.INIT('hf351)
	) name38 (
		\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w10551_
	);
	LUT4 #(
		.INIT('h8caf)
	) name39 (
		\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w10552_
	);
	LUT4 #(
		.INIT('h8000)
	) name40 (
		_w10549_,
		_w10550_,
		_w10551_,
		_w10552_,
		_w10553_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		_w10548_,
		_w10553_,
		_w10554_
	);
	LUT4 #(
		.INIT('h8caf)
	) name42 (
		\ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w10555_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		_w10556_
	);
	LUT3 #(
		.INIT('h51)
	) name44 (
		\ethreg1_MODER_1_DataOut_reg[6]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		_w10557_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name45 (
		\ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w10558_
	);
	LUT3 #(
		.INIT('h80)
	) name46 (
		_w10555_,
		_w10557_,
		_w10558_,
		_w10559_
	);
	LUT4 #(
		.INIT('hf351)
	) name47 (
		\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		_w10560_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w10561_
	);
	LUT4 #(
		.INIT('haf23)
	) name49 (
		\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w10562_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w10563_
	);
	LUT4 #(
		.INIT('hcf45)
	) name51 (
		\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		_w10564_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w10565_
	);
	LUT4 #(
		.INIT('hf351)
	) name53 (
		\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w10566_
	);
	LUT4 #(
		.INIT('h8000)
	) name54 (
		_w10560_,
		_w10562_,
		_w10564_,
		_w10566_,
		_w10567_
	);
	LUT4 #(
		.INIT('h8caf)
	) name55 (
		\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w10568_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name56 (
		\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		_w10569_
	);
	LUT2 #(
		.INIT('h9)
	) name57 (
		\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		_w10570_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name58 (
		\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w10571_
	);
	LUT4 #(
		.INIT('h8000)
	) name59 (
		_w10568_,
		_w10569_,
		_w10570_,
		_w10571_,
		_w10572_
	);
	LUT3 #(
		.INIT('h80)
	) name60 (
		_w10559_,
		_w10567_,
		_w10572_,
		_w10573_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		_w10574_
	);
	LUT3 #(
		.INIT('h20)
	) name62 (
		\RxEnSync_reg/NET0131 ,
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		mrxdv_pad_i_pad,
		_w10575_
	);
	LUT4 #(
		.INIT('h13df)
	) name63 (
		\RxEnSync_reg/NET0131 ,
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		mrxdv_pad_i_pad,
		mtxen_pad_o_pad,
		_w10576_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		_w10574_,
		_w10576_,
		_w10577_
	);
	LUT3 #(
		.INIT('h1b)
	) name65 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[2]_pad ,
		\mtxd_pad_o[2]_pad ,
		_w10578_
	);
	LUT3 #(
		.INIT('he4)
	) name66 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[2]_pad ,
		\mtxd_pad_o[2]_pad ,
		_w10579_
	);
	LUT4 #(
		.INIT('h1be4)
	) name67 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[2]_pad ,
		\mtxd_pad_o[2]_pad ,
		\rxethmac1_crcrx_Crc_reg[29]/NET0131 ,
		_w10580_
	);
	LUT3 #(
		.INIT('h10)
	) name68 (
		_w10574_,
		_w10576_,
		_w10580_,
		_w10581_
	);
	LUT4 #(
		.INIT('h3331)
	) name69 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w10542_,
		_w10543_,
		_w10582_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		\rxethmac1_crcrx_Crc_reg[23]/NET0131 ,
		_w10582_,
		_w10583_
	);
	LUT4 #(
		.INIT('h8f00)
	) name71 (
		_w10554_,
		_w10573_,
		_w10581_,
		_w10583_,
		_w10584_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		\rxethmac1_crcrx_Crc_reg[23]/NET0131 ,
		_w10582_,
		_w10585_
	);
	LUT4 #(
		.INIT('h7000)
	) name73 (
		_w10554_,
		_w10573_,
		_w10581_,
		_w10585_,
		_w10586_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w10584_,
		_w10586_,
		_w10587_
	);
	LUT3 #(
		.INIT('h1b)
	) name75 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[1]_pad ,
		\mtxd_pad_o[1]_pad ,
		_w10588_
	);
	LUT3 #(
		.INIT('he4)
	) name76 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[1]_pad ,
		\mtxd_pad_o[1]_pad ,
		_w10589_
	);
	LUT4 #(
		.INIT('h1be4)
	) name77 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[1]_pad ,
		\mtxd_pad_o[1]_pad ,
		\rxethmac1_crcrx_Crc_reg[30]/NET0131 ,
		_w10590_
	);
	LUT3 #(
		.INIT('h10)
	) name78 (
		_w10574_,
		_w10576_,
		_w10590_,
		_w10591_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		\rxethmac1_crcrx_Crc_reg[24]/NET0131 ,
		_w10582_,
		_w10592_
	);
	LUT4 #(
		.INIT('h8f00)
	) name80 (
		_w10554_,
		_w10573_,
		_w10591_,
		_w10592_,
		_w10593_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		\rxethmac1_crcrx_Crc_reg[24]/NET0131 ,
		_w10582_,
		_w10594_
	);
	LUT4 #(
		.INIT('h7000)
	) name82 (
		_w10554_,
		_w10573_,
		_w10591_,
		_w10594_,
		_w10595_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w10593_,
		_w10595_,
		_w10596_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		\rxethmac1_crcrx_Crc_reg[26]/NET0131 ,
		_w10536_,
		_w10597_
	);
	LUT3 #(
		.INIT('h02)
	) name85 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		wb_rst_i_pad,
		_w10598_
	);
	LUT4 #(
		.INIT('h5f08)
	) name86 (
		_w10533_,
		_w10540_,
		_w10597_,
		_w10598_,
		_w10599_
	);
	LUT3 #(
		.INIT('h01)
	) name87 (
		\ethreg1_MODER_1_DataOut_reg[7]/NET0131 ,
		\maccontrol1_transmitcontrol1_SendingCtrlFrm_reg/NET0131 ,
		\wishbone_TxStatus_reg[12]/NET0131 ,
		_w10600_
	);
	LUT3 #(
		.INIT('h01)
	) name88 (
		\ethreg1_MODER_1_DataOut_reg[5]/NET0131 ,
		\maccontrol1_transmitcontrol1_SendingCtrlFrm_reg/NET0131 ,
		\wishbone_TxStatus_reg[11]/NET0131 ,
		_w10601_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_TxCtrlEndFrm_reg/NET0131 ,
		_w10602_
	);
	LUT3 #(
		.INIT('h27)
	) name90 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_TxCtrlEndFrm_reg/NET0131 ,
		\wishbone_TxEndFrm_reg/NET0131 ,
		_w10603_
	);
	LUT2 #(
		.INIT('h2)
	) name91 (
		\Collision_Tx2_reg/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		_w10604_
	);
	LUT3 #(
		.INIT('hd0)
	) name92 (
		\Collision_Tx2_reg/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		_w10605_
	);
	LUT3 #(
		.INIT('h20)
	) name93 (
		_w10601_,
		_w10603_,
		_w10605_,
		_w10606_
	);
	LUT4 #(
		.INIT('h0800)
	) name94 (
		_w10600_,
		_w10601_,
		_w10603_,
		_w10605_,
		_w10607_
	);
	LUT4 #(
		.INIT('h0001)
	) name95 (
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 ,
		_w10608_
	);
	LUT2 #(
		.INIT('h9)
	) name96 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		_w10608_,
		_w10609_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 ,
		_w10610_
	);
	LUT4 #(
		.INIT('h0002)
	) name98 (
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 ,
		_w10611_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w10610_,
		_w10611_,
		_w10612_
	);
	LUT3 #(
		.INIT('h40)
	) name100 (
		\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 ,
		_w10610_,
		_w10611_,
		_w10613_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 ,
		_w10614_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		_w10608_,
		_w10614_,
		_w10615_
	);
	LUT3 #(
		.INIT('h01)
	) name103 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		_w10616_
	);
	LUT4 #(
		.INIT('h2111)
	) name104 (
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 ,
		_w10608_,
		_w10614_,
		_w10617_
	);
	LUT4 #(
		.INIT('h0001)
	) name105 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 ,
		_w10618_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		_w10619_
	);
	LUT4 #(
		.INIT('hdeee)
	) name107 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10620_
	);
	LUT4 #(
		.INIT('h0080)
	) name108 (
		_w10609_,
		_w10613_,
		_w10617_,
		_w10620_,
		_w10621_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name109 (
		\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10619_,
		_w10622_
	);
	LUT3 #(
		.INIT('h01)
	) name110 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 ,
		_w10623_
	);
	LUT4 #(
		.INIT('h1555)
	) name111 (
		\ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10623_,
		_w10624_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		_w10622_,
		_w10624_,
		_w10625_
	);
	LUT4 #(
		.INIT('h0001)
	) name113 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131 ,
		_w10626_
	);
	LUT3 #(
		.INIT('h80)
	) name114 (
		_w10608_,
		_w10618_,
		_w10626_,
		_w10627_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name115 (
		\ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10626_,
		_w10628_
	);
	LUT4 #(
		.INIT('h4000)
	) name116 (
		\ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10626_,
		_w10629_
	);
	LUT4 #(
		.INIT('h9555)
	) name117 (
		\ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10626_,
		_w10630_
	);
	LUT4 #(
		.INIT('hbfea)
	) name118 (
		\txethmac1_txcounters1_NibCnt_reg[15]/NET0131 ,
		_w10621_,
		_w10625_,
		_w10630_,
		_w10631_
	);
	LUT3 #(
		.INIT('h8c)
	) name119 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 ,
		_w10608_,
		_w10632_
	);
	LUT3 #(
		.INIT('h01)
	) name120 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		_w10633_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		_w10611_,
		_w10633_,
		_w10634_
	);
	LUT4 #(
		.INIT('h4c00)
	) name122 (
		_w10608_,
		_w10611_,
		_w10614_,
		_w10633_,
		_w10635_
	);
	LUT3 #(
		.INIT('h10)
	) name123 (
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		_w10632_,
		_w10635_,
		_w10636_
	);
	LUT3 #(
		.INIT('h2a)
	) name124 (
		\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 ,
		_w10608_,
		_w10616_,
		_w10637_
	);
	LUT3 #(
		.INIT('h15)
	) name125 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10638_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		_w10637_,
		_w10638_,
		_w10639_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name127 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10640_
	);
	LUT4 #(
		.INIT('h1555)
	) name128 (
		\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10619_,
		_w10641_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		_w10640_,
		_w10641_,
		_w10642_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name130 (
		\ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10623_,
		_w10643_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w10627_,
		_w10643_,
		_w10644_
	);
	LUT3 #(
		.INIT('h54)
	) name132 (
		\txethmac1_txcounters1_NibCnt_reg[14]/NET0131 ,
		_w10627_,
		_w10643_,
		_w10645_
	);
	LUT4 #(
		.INIT('h7f00)
	) name133 (
		_w10636_,
		_w10639_,
		_w10642_,
		_w10645_,
		_w10646_
	);
	LUT3 #(
		.INIT('h01)
	) name134 (
		\txethmac1_txcounters1_NibCnt_reg[14]/NET0131 ,
		_w10627_,
		_w10643_,
		_w10647_
	);
	LUT4 #(
		.INIT('h8000)
	) name135 (
		_w10636_,
		_w10639_,
		_w10642_,
		_w10647_,
		_w10648_
	);
	LUT3 #(
		.INIT('h02)
	) name136 (
		_w10631_,
		_w10646_,
		_w10648_,
		_w10649_
	);
	LUT4 #(
		.INIT('h9555)
	) name137 (
		\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10619_,
		_w10650_
	);
	LUT3 #(
		.INIT('hd7)
	) name138 (
		\txethmac1_txcounters1_NibCnt_reg[13]/NET0131 ,
		_w10621_,
		_w10650_,
		_w10651_
	);
	LUT4 #(
		.INIT('h0002)
	) name139 (
		_w10631_,
		_w10646_,
		_w10648_,
		_w10651_,
		_w10652_
	);
	LUT3 #(
		.INIT('hbe)
	) name140 (
		\txethmac1_txcounters1_NibCnt_reg[13]/NET0131 ,
		_w10621_,
		_w10650_,
		_w10653_
	);
	LUT4 #(
		.INIT('h6333)
	) name141 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10654_
	);
	LUT4 #(
		.INIT('hd57f)
	) name142 (
		\txethmac1_txcounters1_NibCnt_reg[12]/NET0131 ,
		_w10636_,
		_w10639_,
		_w10654_,
		_w10655_
	);
	LUT2 #(
		.INIT('h2)
	) name143 (
		_w10653_,
		_w10655_,
		_w10656_
	);
	LUT3 #(
		.INIT('h40)
	) name144 (
		_w10622_,
		_w10624_,
		_w10630_,
		_w10657_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		_w10621_,
		_w10657_,
		_w10658_
	);
	LUT4 #(
		.INIT('h2a80)
	) name146 (
		\txethmac1_txcounters1_NibCnt_reg[15]/NET0131 ,
		_w10621_,
		_w10625_,
		_w10630_,
		_w10659_
	);
	LUT4 #(
		.INIT('h007f)
	) name147 (
		_w10636_,
		_w10639_,
		_w10642_,
		_w10644_,
		_w10660_
	);
	LUT4 #(
		.INIT('h0010)
	) name148 (
		_w10627_,
		_w10640_,
		_w10641_,
		_w10643_,
		_w10661_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name149 (
		\txethmac1_txcounters1_NibCnt_reg[14]/NET0131 ,
		_w10636_,
		_w10639_,
		_w10661_,
		_w10662_
	);
	LUT4 #(
		.INIT('h3133)
	) name150 (
		_w10631_,
		_w10659_,
		_w10660_,
		_w10662_,
		_w10663_
	);
	LUT4 #(
		.INIT('h1300)
	) name151 (
		_w10649_,
		_w10652_,
		_w10656_,
		_w10663_,
		_w10664_
	);
	LUT4 #(
		.INIT('h1222)
	) name152 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[11]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10665_
	);
	LUT4 #(
		.INIT('h7f00)
	) name153 (
		_w10609_,
		_w10613_,
		_w10617_,
		_w10665_,
		_w10666_
	);
	LUT4 #(
		.INIT('h2111)
	) name154 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[11]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10667_
	);
	LUT4 #(
		.INIT('h8000)
	) name155 (
		_w10609_,
		_w10613_,
		_w10617_,
		_w10667_,
		_w10668_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		_w10666_,
		_w10668_,
		_w10669_
	);
	LUT4 #(
		.INIT('h4000)
	) name157 (
		\txethmac1_txcounters1_NibCnt_reg[10]/NET0131 ,
		_w10609_,
		_w10613_,
		_w10617_,
		_w10670_
	);
	LUT4 #(
		.INIT('h6333)
	) name158 (
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 ,
		_w10608_,
		_w10614_,
		_w10671_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		\txethmac1_txcounters1_NibCnt_reg[10]/NET0131 ,
		_w10671_,
		_w10672_
	);
	LUT3 #(
		.INIT('h23)
	) name160 (
		_w10636_,
		_w10670_,
		_w10672_,
		_w10673_
	);
	LUT3 #(
		.INIT('h95)
	) name161 (
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		_w10608_,
		_w10614_,
		_w10674_
	);
	LUT3 #(
		.INIT('h07)
	) name162 (
		_w10609_,
		_w10613_,
		_w10674_,
		_w10675_
	);
	LUT3 #(
		.INIT('h63)
	) name163 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 ,
		_w10608_,
		_w10676_
	);
	LUT4 #(
		.INIT('ha802)
	) name164 (
		\txethmac1_txcounters1_NibCnt_reg[8]/NET0131 ,
		_w10615_,
		_w10632_,
		_w10634_,
		_w10677_
	);
	LUT4 #(
		.INIT('h54fd)
	) name165 (
		\txethmac1_txcounters1_NibCnt_reg[9]/NET0131 ,
		_w10636_,
		_w10675_,
		_w10677_,
		_w10678_
	);
	LUT3 #(
		.INIT('h08)
	) name166 (
		_w10669_,
		_w10673_,
		_w10678_,
		_w10679_
	);
	LUT4 #(
		.INIT('h4888)
	) name167 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[11]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10680_
	);
	LUT4 #(
		.INIT('h8000)
	) name168 (
		_w10609_,
		_w10613_,
		_w10617_,
		_w10680_,
		_w10681_
	);
	LUT4 #(
		.INIT('h8444)
	) name169 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[11]/NET0131 ,
		_w10608_,
		_w10618_,
		_w10682_
	);
	LUT4 #(
		.INIT('h7f00)
	) name170 (
		_w10609_,
		_w10613_,
		_w10617_,
		_w10682_,
		_w10683_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		_w10681_,
		_w10683_,
		_w10684_
	);
	LUT4 #(
		.INIT('h00ef)
	) name172 (
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		_w10632_,
		_w10635_,
		_w10671_,
		_w10685_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name173 (
		\txethmac1_txcounters1_NibCnt_reg[10]/NET0131 ,
		_w10609_,
		_w10613_,
		_w10617_,
		_w10686_
	);
	LUT4 #(
		.INIT('h0100)
	) name174 (
		_w10666_,
		_w10668_,
		_w10685_,
		_w10686_,
		_w10687_
	);
	LUT2 #(
		.INIT('h2)
	) name175 (
		_w10684_,
		_w10687_,
		_w10688_
	);
	LUT4 #(
		.INIT('hbfea)
	) name176 (
		\txethmac1_txcounters1_NibCnt_reg[12]/NET0131 ,
		_w10636_,
		_w10639_,
		_w10654_,
		_w10689_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		_w10653_,
		_w10689_,
		_w10690_
	);
	LUT4 #(
		.INIT('h8a00)
	) name178 (
		_w10649_,
		_w10679_,
		_w10688_,
		_w10690_,
		_w10691_
	);
	LUT3 #(
		.INIT('hd7)
	) name179 (
		\txethmac1_txcounters1_NibCnt_reg[7]/NET0131 ,
		_w10609_,
		_w10612_,
		_w10692_
	);
	LUT3 #(
		.INIT('hbe)
	) name180 (
		\txethmac1_txcounters1_NibCnt_reg[7]/NET0131 ,
		_w10609_,
		_w10612_,
		_w10693_
	);
	LUT3 #(
		.INIT('he0)
	) name181 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		_w10694_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 ,
		_w10695_
	);
	LUT3 #(
		.INIT('h45)
	) name183 (
		\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 ,
		_w10694_,
		_w10695_,
		_w10696_
	);
	LUT3 #(
		.INIT('h10)
	) name184 (
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 ,
		_w10697_
	);
	LUT3 #(
		.INIT('h45)
	) name185 (
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w10694_,
		_w10697_,
		_w10698_
	);
	LUT2 #(
		.INIT('h4)
	) name186 (
		_w10696_,
		_w10698_,
		_w10699_
	);
	LUT3 #(
		.INIT('ha2)
	) name187 (
		_w10692_,
		_w10693_,
		_w10699_,
		_w10700_
	);
	LUT2 #(
		.INIT('h6)
	) name188 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 ,
		_w10701_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w10702_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w10703_
	);
	LUT3 #(
		.INIT('h17)
	) name191 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w10704_
	);
	LUT4 #(
		.INIT('hffe1)
	) name192 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10705_
	);
	LUT4 #(
		.INIT('h8e00)
	) name193 (
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w10701_,
		_w10704_,
		_w10705_,
		_w10706_
	);
	LUT4 #(
		.INIT('h001f)
	) name194 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		_w10707_
	);
	LUT4 #(
		.INIT('he000)
	) name195 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		_w10708_
	);
	LUT4 #(
		.INIT('h1eff)
	) name196 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10709_
	);
	LUT4 #(
		.INIT('hfd00)
	) name197 (
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10707_,
		_w10708_,
		_w10709_,
		_w10710_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		_w10706_,
		_w10710_,
		_w10711_
	);
	LUT4 #(
		.INIT('h3c1e)
	) name199 (
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 ,
		_w10610_,
		_w10712_
	);
	LUT3 #(
		.INIT('hde)
	) name200 (
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10694_,
		_w10713_
	);
	LUT3 #(
		.INIT('he0)
	) name201 (
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w10712_,
		_w10713_,
		_w10714_
	);
	LUT4 #(
		.INIT('hb7bb)
	) name202 (
		\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w10694_,
		_w10695_,
		_w10715_
	);
	LUT3 #(
		.INIT('h70)
	) name203 (
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w10712_,
		_w10715_,
		_w10716_
	);
	LUT4 #(
		.INIT('h8a00)
	) name204 (
		_w10692_,
		_w10711_,
		_w10714_,
		_w10716_,
		_w10717_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		_w10700_,
		_w10717_,
		_w10718_
	);
	LUT3 #(
		.INIT('hbe)
	) name206 (
		\txethmac1_txcounters1_NibCnt_reg[8]/NET0131 ,
		_w10634_,
		_w10676_,
		_w10719_
	);
	LUT4 #(
		.INIT('hab00)
	) name207 (
		\txethmac1_txcounters1_NibCnt_reg[9]/NET0131 ,
		_w10636_,
		_w10675_,
		_w10719_,
		_w10720_
	);
	LUT3 #(
		.INIT('h80)
	) name208 (
		_w10669_,
		_w10673_,
		_w10720_,
		_w10721_
	);
	LUT4 #(
		.INIT('h8000)
	) name209 (
		_w10649_,
		_w10690_,
		_w10718_,
		_w10721_,
		_w10722_
	);
	LUT4 #(
		.INIT('h1555)
	) name210 (
		_w10629_,
		_w10636_,
		_w10639_,
		_w10661_,
		_w10723_
	);
	LUT4 #(
		.INIT('h0526)
	) name211 (
		\ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131 ,
		_w10628_,
		_w10658_,
		_w10723_,
		_w10724_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		_w10606_,
		_w10724_,
		_w10725_
	);
	LUT4 #(
		.INIT('hfd00)
	) name213 (
		_w10664_,
		_w10691_,
		_w10722_,
		_w10725_,
		_w10726_
	);
	LUT3 #(
		.INIT('h80)
	) name214 (
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w10727_
	);
	LUT3 #(
		.INIT('hd0)
	) name215 (
		\Collision_Tx2_reg/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w10728_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		_w10727_,
		_w10728_,
		_w10729_
	);
	LUT3 #(
		.INIT('h51)
	) name217 (
		\ethreg1_MODER_1_DataOut_reg[6]/NET0131 ,
		\ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		_w10730_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name218 (
		\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[13]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[15]/NET0131 ,
		_w10731_
	);
	LUT4 #(
		.INIT('hf351)
	) name219 (
		\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		_w10732_
	);
	LUT3 #(
		.INIT('h80)
	) name220 (
		_w10730_,
		_w10731_,
		_w10732_,
		_w10733_
	);
	LUT4 #(
		.INIT('h8acf)
	) name221 (
		\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[13]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		_w10734_
	);
	LUT4 #(
		.INIT('hcf45)
	) name222 (
		\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[10]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[8]/NET0131 ,
		_w10735_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name223 (
		\ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 ,
		_w10736_
	);
	LUT4 #(
		.INIT('haf23)
	) name224 (
		\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 ,
		\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[7]/NET0131 ,
		_w10737_
	);
	LUT4 #(
		.INIT('h8000)
	) name225 (
		_w10734_,
		_w10735_,
		_w10736_,
		_w10737_,
		_w10738_
	);
	LUT4 #(
		.INIT('haf23)
	) name226 (
		\ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w10739_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name227 (
		\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[11]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 ,
		_w10740_
	);
	LUT4 #(
		.INIT('hf531)
	) name228 (
		\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 ,
		_w10741_
	);
	LUT4 #(
		.INIT('hf531)
	) name229 (
		\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[10]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[15]/NET0131 ,
		_w10742_
	);
	LUT4 #(
		.INIT('h8000)
	) name230 (
		_w10739_,
		_w10740_,
		_w10741_,
		_w10742_,
		_w10743_
	);
	LUT3 #(
		.INIT('h80)
	) name231 (
		_w10733_,
		_w10738_,
		_w10743_,
		_w10744_
	);
	LUT4 #(
		.INIT('h00d0)
	) name232 (
		\Collision_Tx2_reg/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		\wishbone_TxUnderRun_reg/NET0131 ,
		_w10745_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		_w10728_,
		_w10745_,
		_w10746_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[8]/NET0131 ,
		_w10747_
	);
	LUT4 #(
		.INIT('h8acf)
	) name235 (
		\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[7]/NET0131 ,
		_w10748_
	);
	LUT2 #(
		.INIT('h4)
	) name236 (
		_w10747_,
		_w10748_,
		_w10749_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name237 (
		\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[14]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w10750_
	);
	LUT4 #(
		.INIT('h8acf)
	) name238 (
		\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[14]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		_w10751_
	);
	LUT4 #(
		.INIT('hf531)
	) name239 (
		\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 ,
		_w10752_
	);
	LUT4 #(
		.INIT('h8caf)
	) name240 (
		\ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[11]/NET0131 ,
		_w10753_
	);
	LUT4 #(
		.INIT('h8000)
	) name241 (
		_w10750_,
		_w10751_,
		_w10752_,
		_w10753_,
		_w10754_
	);
	LUT2 #(
		.INIT('h8)
	) name242 (
		_w10749_,
		_w10754_,
		_w10755_
	);
	LUT3 #(
		.INIT('h40)
	) name243 (
		_w10746_,
		_w10749_,
		_w10754_,
		_w10756_
	);
	LUT3 #(
		.INIT('h15)
	) name244 (
		_w10729_,
		_w10744_,
		_w10756_,
		_w10757_
	);
	LUT4 #(
		.INIT('hf531)
	) name245 (
		\ethreg1_IPGR1_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_IPGR1_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10758_
	);
	LUT4 #(
		.INIT('h8caf)
	) name246 (
		\ethreg1_IPGR1_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_IPGR1_0_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w10759_
	);
	LUT2 #(
		.INIT('h4)
	) name247 (
		_w10758_,
		_w10759_,
		_w10760_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name248 (
		\ethreg1_IPGR1_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_IPGR1_0_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w10761_
	);
	LUT3 #(
		.INIT('h0b)
	) name249 (
		\ethreg1_IPGR1_0_DataOut_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w10762_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		\ethreg1_IPGR1_0_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w10763_
	);
	LUT3 #(
		.INIT('h01)
	) name251 (
		_w10761_,
		_w10762_,
		_w10763_,
		_w10764_
	);
	LUT4 #(
		.INIT('h8caf)
	) name252 (
		\ethreg1_IPGR1_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_IPGR1_0_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10765_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		_w10759_,
		_w10765_,
		_w10766_
	);
	LUT4 #(
		.INIT('hf531)
	) name254 (
		\ethreg1_IPGR1_0_DataOut_reg[5]/NET0131 ,
		\ethreg1_IPGR1_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w10767_
	);
	LUT4 #(
		.INIT('h4500)
	) name255 (
		_w10760_,
		_w10764_,
		_w10766_,
		_w10767_,
		_w10768_
	);
	LUT4 #(
		.INIT('h8caf)
	) name256 (
		\ethreg1_IPGR2_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_IPGR2_0_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w10769_
	);
	LUT4 #(
		.INIT('hf531)
	) name257 (
		\ethreg1_IPGR2_0_DataOut_reg[5]/NET0131 ,
		\ethreg1_IPGR2_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w10770_
	);
	LUT4 #(
		.INIT('hf531)
	) name258 (
		\ethreg1_IPGR2_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_IPGR2_0_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10771_
	);
	LUT3 #(
		.INIT('h80)
	) name259 (
		_w10769_,
		_w10770_,
		_w10771_,
		_w10772_
	);
	LUT4 #(
		.INIT('h8caf)
	) name260 (
		\ethreg1_IPGR2_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_IPGR2_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w10773_
	);
	LUT2 #(
		.INIT('h2)
	) name261 (
		\ethreg1_IPGR2_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10774_
	);
	LUT4 #(
		.INIT('haf23)
	) name262 (
		\ethreg1_IPGR2_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_IPGR2_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10775_
	);
	LUT4 #(
		.INIT('h8caf)
	) name263 (
		\ethreg1_IPGR2_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_IPGR2_0_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w10776_
	);
	LUT4 #(
		.INIT('hf531)
	) name264 (
		\ethreg1_IPGR2_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_IPGR2_0_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w10777_
	);
	LUT4 #(
		.INIT('h8000)
	) name265 (
		_w10773_,
		_w10775_,
		_w10776_,
		_w10777_,
		_w10778_
	);
	LUT2 #(
		.INIT('h2)
	) name266 (
		\CarrierSense_Tx2_reg/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		_w10779_
	);
	LUT4 #(
		.INIT('h0b00)
	) name267 (
		\ethreg1_IPGR1_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		\txethmac1_txstatem1_Rule1_reg/NET0131 ,
		\txethmac1_txstatem1_StateIPG_reg/NET0131 ,
		_w10780_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		_w10779_,
		_w10780_,
		_w10781_
	);
	LUT3 #(
		.INIT('h70)
	) name269 (
		_w10772_,
		_w10778_,
		_w10781_,
		_w10782_
	);
	LUT2 #(
		.INIT('h4)
	) name270 (
		_w10768_,
		_w10782_,
		_w10783_
	);
	LUT4 #(
		.INIT('h8000)
	) name271 (
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w10784_
	);
	LUT4 #(
		.INIT('h8421)
	) name272 (
		\ethreg1_COLLCONF_2_DataOut_reg[2]/NET0131 ,
		\ethreg1_COLLCONF_2_DataOut_reg[3]/NET0131 ,
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w10785_
	);
	LUT4 #(
		.INIT('h8421)
	) name273 (
		\ethreg1_COLLCONF_2_DataOut_reg[0]/NET0131 ,
		\ethreg1_COLLCONF_2_DataOut_reg[1]/NET0131 ,
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		_w10786_
	);
	LUT3 #(
		.INIT('h2a)
	) name274 (
		\txethmac1_ColWindow_reg/NET0131 ,
		_w10785_,
		_w10786_,
		_w10787_
	);
	LUT4 #(
		.INIT('h0001)
	) name275 (
		\txethmac1_random1_RandomLatched_reg[6]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[7]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[8]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[9]/NET0131 ,
		_w10788_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		\txethmac1_random1_RandomLatched_reg[0]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[1]/NET0131 ,
		_w10789_
	);
	LUT4 #(
		.INIT('h0001)
	) name277 (
		\txethmac1_random1_RandomLatched_reg[2]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[3]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[4]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[5]/NET0131 ,
		_w10790_
	);
	LUT4 #(
		.INIT('h1555)
	) name278 (
		\ethreg1_MODER_1_DataOut_reg[0]/NET0131 ,
		_w10788_,
		_w10789_,
		_w10790_,
		_w10791_
	);
	LUT3 #(
		.INIT('h2a)
	) name279 (
		_w10784_,
		_w10787_,
		_w10791_,
		_w10792_
	);
	LUT4 #(
		.INIT('hf531)
	) name280 (
		\txethmac1_random1_RandomLatched_reg[1]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w10793_
	);
	LUT4 #(
		.INIT('h8caf)
	) name281 (
		\txethmac1_random1_RandomLatched_reg[1]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[6]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 ,
		_w10794_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		_w10793_,
		_w10794_,
		_w10795_
	);
	LUT4 #(
		.INIT('haf23)
	) name283 (
		\txethmac1_random1_RandomLatched_reg[8]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[9]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[8]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 ,
		_w10796_
	);
	LUT4 #(
		.INIT('haf23)
	) name284 (
		\txethmac1_random1_RandomLatched_reg[3]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[8]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[8]/NET0131 ,
		_w10797_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name285 (
		\txethmac1_random1_RandomLatched_reg[3]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w10798_
	);
	LUT4 #(
		.INIT('hf531)
	) name286 (
		\txethmac1_random1_RandomLatched_reg[6]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[7]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[7]/NET0131 ,
		_w10799_
	);
	LUT4 #(
		.INIT('h8000)
	) name287 (
		_w10796_,
		_w10797_,
		_w10798_,
		_w10799_,
		_w10800_
	);
	LUT4 #(
		.INIT('h8000)
	) name288 (
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10801_
	);
	LUT2 #(
		.INIT('h8)
	) name289 (
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w10802_
	);
	LUT4 #(
		.INIT('h8000)
	) name290 (
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		\txethmac1_txstatem1_StateBackOff_reg/NET0131 ,
		_w10803_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		_w10801_,
		_w10803_,
		_w10804_
	);
	LUT4 #(
		.INIT('hf531)
	) name292 (
		\txethmac1_random1_RandomLatched_reg[0]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		_w10805_
	);
	LUT4 #(
		.INIT('h8caf)
	) name293 (
		\txethmac1_random1_RandomLatched_reg[2]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[9]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 ,
		_w10806_
	);
	LUT2 #(
		.INIT('h6)
	) name294 (
		\txethmac1_random1_RandomLatched_reg[5]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		_w10807_
	);
	LUT4 #(
		.INIT('h8caf)
	) name295 (
		\txethmac1_random1_RandomLatched_reg[0]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[7]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[7]/NET0131 ,
		_w10808_
	);
	LUT4 #(
		.INIT('h0800)
	) name296 (
		_w10805_,
		_w10806_,
		_w10807_,
		_w10808_,
		_w10809_
	);
	LUT4 #(
		.INIT('h8000)
	) name297 (
		_w10795_,
		_w10800_,
		_w10804_,
		_w10809_,
		_w10810_
	);
	LUT3 #(
		.INIT('h20)
	) name298 (
		\CarrierSense_Tx2_reg/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		_w10811_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		\txethmac1_txstatem1_StateBackOff_reg/NET0131 ,
		\wishbone_TxUnderRun_reg/NET0131 ,
		_w10812_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		_w10811_,
		_w10812_,
		_w10813_
	);
	LUT3 #(
		.INIT('h10)
	) name301 (
		_w10792_,
		_w10810_,
		_w10813_,
		_w10814_
	);
	LUT3 #(
		.INIT('h20)
	) name302 (
		_w10757_,
		_w10783_,
		_w10814_,
		_w10815_
	);
	LUT3 #(
		.INIT('h10)
	) name303 (
		_w10607_,
		_w10726_,
		_w10815_,
		_w10816_
	);
	LUT3 #(
		.INIT('h10)
	) name304 (
		_w10601_,
		_w10603_,
		_w10605_,
		_w10817_
	);
	LUT4 #(
		.INIT('h0200)
	) name305 (
		_w10600_,
		_w10601_,
		_w10603_,
		_w10605_,
		_w10818_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		_w10724_,
		_w10817_,
		_w10819_
	);
	LUT4 #(
		.INIT('hfd00)
	) name307 (
		_w10664_,
		_w10691_,
		_w10722_,
		_w10819_,
		_w10820_
	);
	LUT3 #(
		.INIT('hd0)
	) name308 (
		\Collision_Tx2_reg/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\txethmac1_txstatem1_StatePAD_reg/NET0131 ,
		_w10821_
	);
	LUT2 #(
		.INIT('h4)
	) name309 (
		_w10601_,
		_w10821_,
		_w10822_
	);
	LUT2 #(
		.INIT('h8)
	) name310 (
		_w10724_,
		_w10822_,
		_w10823_
	);
	LUT4 #(
		.INIT('hfd00)
	) name311 (
		_w10664_,
		_w10691_,
		_w10722_,
		_w10823_,
		_w10824_
	);
	LUT4 #(
		.INIT('hd000)
	) name312 (
		\Collision_Tx2_reg/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		\wishbone_TxUnderRun_reg/NET0131 ,
		_w10825_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name313 (
		\Collision_Tx2_reg/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		\wishbone_TxUnderRun_reg/NET0131 ,
		_w10826_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		\txethmac1_txstatem1_StatePAD_reg/NET0131 ,
		_w10827_
	);
	LUT4 #(
		.INIT('h0001)
	) name315 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		\txethmac1_txstatem1_StatePAD_reg/NET0131 ,
		_w10828_
	);
	LUT3 #(
		.INIT('h70)
	) name316 (
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w10801_,
		_w10828_,
		_w10829_
	);
	LUT4 #(
		.INIT('h080f)
	) name317 (
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w10801_,
		_w10826_,
		_w10828_,
		_w10830_
	);
	LUT4 #(
		.INIT('h0004)
	) name318 (
		\txethmac1_txcounters1_NibCnt_reg[11]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[12]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[13]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10831_
	);
	LUT4 #(
		.INIT('h4000)
	) name319 (
		\ethreg1_MODER_1_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[10]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w10832_
	);
	LUT4 #(
		.INIT('h4000)
	) name320 (
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[7]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[8]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[9]/NET0131 ,
		_w10833_
	);
	LUT4 #(
		.INIT('h8000)
	) name321 (
		_w10727_,
		_w10831_,
		_w10832_,
		_w10833_,
		_w10834_
	);
	LUT3 #(
		.INIT('h10)
	) name322 (
		\maccontrol1_receivecontrol1_Pause_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w10835_
	);
	LUT4 #(
		.INIT('h2e3f)
	) name323 (
		\maccontrol1_receivecontrol1_Pause_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w10836_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		\txethmac1_txstatem1_StateDefer_reg/NET0131 ,
		_w10836_,
		_w10837_
	);
	LUT3 #(
		.INIT('hd0)
	) name325 (
		\CarrierSense_Tx2_reg/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\txethmac1_txstatem1_StateDefer_reg/NET0131 ,
		_w10838_
	);
	LUT2 #(
		.INIT('h4)
	) name326 (
		_w10834_,
		_w10838_,
		_w10839_
	);
	LUT4 #(
		.INIT('h0105)
	) name327 (
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w10784_,
		_w10801_,
		_w10840_
	);
	LUT4 #(
		.INIT('h2700)
	) name328 (
		_w10834_,
		_w10837_,
		_w10838_,
		_w10840_,
		_w10841_
	);
	LUT2 #(
		.INIT('h4)
	) name329 (
		_w10830_,
		_w10841_,
		_w10842_
	);
	LUT4 #(
		.INIT('h0100)
	) name330 (
		_w10818_,
		_w10820_,
		_w10824_,
		_w10842_,
		_w10843_
	);
	LUT2 #(
		.INIT('h2)
	) name331 (
		\txethmac1_txstatem1_StateDefer_reg/NET0131 ,
		_w10836_,
		_w10844_
	);
	LUT3 #(
		.INIT('h01)
	) name332 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w10845_
	);
	LUT3 #(
		.INIT('h01)
	) name333 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		\txethmac1_txstatem1_StatePAD_reg/NET0131 ,
		_w10846_
	);
	LUT2 #(
		.INIT('h8)
	) name334 (
		_w10845_,
		_w10846_,
		_w10847_
	);
	LUT2 #(
		.INIT('h7)
	) name335 (
		_w10845_,
		_w10846_,
		_w10848_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		\txethmac1_txstatem1_StateBackOff_reg/NET0131 ,
		\txethmac1_txstatem1_StateIPG_reg/NET0131 ,
		_w10849_
	);
	LUT3 #(
		.INIT('h80)
	) name337 (
		_w10845_,
		_w10846_,
		_w10849_,
		_w10850_
	);
	LUT4 #(
		.INIT('h9a55)
	) name338 (
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		_w10834_,
		_w10844_,
		_w10850_,
		_w10851_
	);
	LUT3 #(
		.INIT('h80)
	) name339 (
		_w10816_,
		_w10843_,
		_w10851_,
		_w10852_
	);
	LUT3 #(
		.INIT('h80)
	) name340 (
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w10853_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		_w10801_,
		_w10853_,
		_w10854_
	);
	LUT4 #(
		.INIT('h4f00)
	) name342 (
		_w10834_,
		_w10844_,
		_w10850_,
		_w10854_,
		_w10855_
	);
	LUT3 #(
		.INIT('h80)
	) name343 (
		\txethmac1_txcounters1_NibCnt_reg[7]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[8]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[9]/NET0131 ,
		_w10856_
	);
	LUT2 #(
		.INIT('h8)
	) name344 (
		\txethmac1_txcounters1_NibCnt_reg[10]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[11]/NET0131 ,
		_w10857_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name345 (
		\txethmac1_txcounters1_NibCnt_reg[10]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[11]/NET0131 ,
		_w10855_,
		_w10856_,
		_w10858_
	);
	LUT3 #(
		.INIT('h80)
	) name346 (
		_w10816_,
		_w10843_,
		_w10858_,
		_w10859_
	);
	LUT4 #(
		.INIT('h1555)
	) name347 (
		\txethmac1_txcounters1_NibCnt_reg[12]/NET0131 ,
		_w10855_,
		_w10856_,
		_w10857_,
		_w10860_
	);
	LUT3 #(
		.INIT('h80)
	) name348 (
		\txethmac1_txcounters1_NibCnt_reg[10]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[11]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[12]/NET0131 ,
		_w10861_
	);
	LUT3 #(
		.INIT('h80)
	) name349 (
		_w10855_,
		_w10856_,
		_w10861_,
		_w10862_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		_w10860_,
		_w10862_,
		_w10863_
	);
	LUT3 #(
		.INIT('h80)
	) name351 (
		_w10816_,
		_w10843_,
		_w10863_,
		_w10864_
	);
	LUT3 #(
		.INIT('h6a)
	) name352 (
		\txethmac1_txcounters1_NibCnt_reg[10]/NET0131 ,
		_w10855_,
		_w10856_,
		_w10865_
	);
	LUT3 #(
		.INIT('h80)
	) name353 (
		_w10816_,
		_w10843_,
		_w10865_,
		_w10866_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name354 (
		\txethmac1_txcounters1_NibCnt_reg[13]/NET0131 ,
		_w10855_,
		_w10856_,
		_w10861_,
		_w10867_
	);
	LUT3 #(
		.INIT('h80)
	) name355 (
		_w10816_,
		_w10843_,
		_w10867_,
		_w10868_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		\txethmac1_txcounters1_NibCnt_reg[13]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[14]/NET0131 ,
		_w10869_
	);
	LUT4 #(
		.INIT('h8000)
	) name357 (
		_w10855_,
		_w10856_,
		_w10861_,
		_w10869_,
		_w10870_
	);
	LUT3 #(
		.INIT('h6c)
	) name358 (
		\txethmac1_txcounters1_NibCnt_reg[13]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[14]/NET0131 ,
		_w10862_,
		_w10871_
	);
	LUT3 #(
		.INIT('h80)
	) name359 (
		_w10816_,
		_w10843_,
		_w10871_,
		_w10872_
	);
	LUT3 #(
		.INIT('h80)
	) name360 (
		\txethmac1_txcounters1_NibCnt_reg[13]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[14]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[15]/NET0131 ,
		_w10873_
	);
	LUT4 #(
		.INIT('h8000)
	) name361 (
		_w10855_,
		_w10856_,
		_w10861_,
		_w10873_,
		_w10874_
	);
	LUT3 #(
		.INIT('h0e)
	) name362 (
		\txethmac1_txcounters1_NibCnt_reg[15]/NET0131 ,
		_w10870_,
		_w10874_,
		_w10875_
	);
	LUT3 #(
		.INIT('h80)
	) name363 (
		_w10816_,
		_w10843_,
		_w10875_,
		_w10876_
	);
	LUT4 #(
		.INIT('h4000)
	) name364 (
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w10845_,
		_w10846_,
		_w10849_,
		_w10877_
	);
	LUT4 #(
		.INIT('h1055)
	) name365 (
		_w10703_,
		_w10834_,
		_w10844_,
		_w10877_,
		_w10878_
	);
	LUT4 #(
		.INIT('h20aa)
	) name366 (
		_w10702_,
		_w10834_,
		_w10844_,
		_w10850_,
		_w10879_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		_w10878_,
		_w10879_,
		_w10880_
	);
	LUT3 #(
		.INIT('h80)
	) name368 (
		_w10816_,
		_w10843_,
		_w10880_,
		_w10881_
	);
	LUT3 #(
		.INIT('h07)
	) name369 (
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w10882_
	);
	LUT4 #(
		.INIT('h4000)
	) name370 (
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w10845_,
		_w10846_,
		_w10849_,
		_w10883_
	);
	LUT4 #(
		.INIT('h040f)
	) name371 (
		_w10834_,
		_w10844_,
		_w10882_,
		_w10883_,
		_w10884_
	);
	LUT4 #(
		.INIT('h20aa)
	) name372 (
		_w10727_,
		_w10834_,
		_w10844_,
		_w10850_,
		_w10885_
	);
	LUT2 #(
		.INIT('h2)
	) name373 (
		_w10884_,
		_w10885_,
		_w10886_
	);
	LUT3 #(
		.INIT('h80)
	) name374 (
		_w10816_,
		_w10843_,
		_w10886_,
		_w10887_
	);
	LUT4 #(
		.INIT('h20aa)
	) name375 (
		_w10801_,
		_w10834_,
		_w10844_,
		_w10850_,
		_w10888_
	);
	LUT4 #(
		.INIT('h007f)
	) name376 (
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10889_
	);
	LUT4 #(
		.INIT('h4000)
	) name377 (
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10845_,
		_w10846_,
		_w10849_,
		_w10890_
	);
	LUT4 #(
		.INIT('h040f)
	) name378 (
		_w10834_,
		_w10844_,
		_w10889_,
		_w10890_,
		_w10891_
	);
	LUT2 #(
		.INIT('h4)
	) name379 (
		_w10888_,
		_w10891_,
		_w10892_
	);
	LUT3 #(
		.INIT('h80)
	) name380 (
		_w10816_,
		_w10843_,
		_w10892_,
		_w10893_
	);
	LUT2 #(
		.INIT('h8)
	) name381 (
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10801_,
		_w10894_
	);
	LUT4 #(
		.INIT('h4f00)
	) name382 (
		_w10834_,
		_w10844_,
		_w10850_,
		_w10894_,
		_w10895_
	);
	LUT2 #(
		.INIT('h1)
	) name383 (
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10801_,
		_w10896_
	);
	LUT4 #(
		.INIT('h4000)
	) name384 (
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10845_,
		_w10846_,
		_w10849_,
		_w10897_
	);
	LUT4 #(
		.INIT('h040f)
	) name385 (
		_w10834_,
		_w10844_,
		_w10896_,
		_w10897_,
		_w10898_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		_w10895_,
		_w10898_,
		_w10899_
	);
	LUT3 #(
		.INIT('h80)
	) name387 (
		_w10816_,
		_w10843_,
		_w10899_,
		_w10900_
	);
	LUT2 #(
		.INIT('h8)
	) name388 (
		_w10801_,
		_w10802_,
		_w10901_
	);
	LUT4 #(
		.INIT('h4f00)
	) name389 (
		_w10834_,
		_w10844_,
		_w10850_,
		_w10901_,
		_w10902_
	);
	LUT3 #(
		.INIT('h0e)
	) name390 (
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w10895_,
		_w10902_,
		_w10903_
	);
	LUT3 #(
		.INIT('h80)
	) name391 (
		_w10816_,
		_w10843_,
		_w10903_,
		_w10904_
	);
	LUT3 #(
		.INIT('h32)
	) name392 (
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w10855_,
		_w10902_,
		_w10905_
	);
	LUT3 #(
		.INIT('h80)
	) name393 (
		_w10816_,
		_w10843_,
		_w10905_,
		_w10906_
	);
	LUT2 #(
		.INIT('h6)
	) name394 (
		\txethmac1_txcounters1_NibCnt_reg[7]/NET0131 ,
		_w10855_,
		_w10907_
	);
	LUT3 #(
		.INIT('h80)
	) name395 (
		_w10816_,
		_w10843_,
		_w10907_,
		_w10908_
	);
	LUT3 #(
		.INIT('h6c)
	) name396 (
		\txethmac1_txcounters1_NibCnt_reg[7]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[8]/NET0131 ,
		_w10855_,
		_w10909_
	);
	LUT3 #(
		.INIT('h80)
	) name397 (
		_w10816_,
		_w10843_,
		_w10909_,
		_w10910_
	);
	LUT4 #(
		.INIT('h78f0)
	) name398 (
		\txethmac1_txcounters1_NibCnt_reg[7]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[8]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[9]/NET0131 ,
		_w10855_,
		_w10911_
	);
	LUT3 #(
		.INIT('h80)
	) name399 (
		_w10816_,
		_w10843_,
		_w10911_,
		_w10912_
	);
	LUT3 #(
		.INIT('h01)
	) name400 (
		\txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		_w10913_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w10914_
	);
	LUT3 #(
		.INIT('h01)
	) name402 (
		\txethmac1_txcrc_Crc_reg[26]/NET0131 ,
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w10915_
	);
	LUT2 #(
		.INIT('h7)
	) name403 (
		_w10913_,
		_w10915_,
		_w10916_
	);
	LUT3 #(
		.INIT('h01)
	) name404 (
		\txethmac1_txcrc_Crc_reg[27]/NET0131 ,
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w10917_
	);
	LUT2 #(
		.INIT('h7)
	) name405 (
		_w10913_,
		_w10917_,
		_w10918_
	);
	LUT3 #(
		.INIT('h0b)
	) name406 (
		\ethreg1_IPGR2_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		\txethmac1_txstatem1_Rule1_reg/NET0131 ,
		_w10919_
	);
	LUT2 #(
		.INIT('h4)
	) name407 (
		_w10770_,
		_w10919_,
		_w10920_
	);
	LUT4 #(
		.INIT('h5010)
	) name408 (
		\ethreg1_IPGR2_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_IPGR2_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10921_
	);
	LUT4 #(
		.INIT('h0c04)
	) name409 (
		_w10769_,
		_w10771_,
		_w10774_,
		_w10777_,
		_w10922_
	);
	LUT2 #(
		.INIT('h8)
	) name410 (
		_w10776_,
		_w10919_,
		_w10923_
	);
	LUT4 #(
		.INIT('h5455)
	) name411 (
		_w10920_,
		_w10921_,
		_w10922_,
		_w10923_,
		_w10924_
	);
	LUT4 #(
		.INIT('h4f00)
	) name412 (
		\ethreg1_IPGT_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		\txethmac1_txstatem1_Rule1_reg/NET0131 ,
		\txethmac1_txstatem1_StateIPG_reg/NET0131 ,
		_w10925_
	);
	LUT4 #(
		.INIT('hf531)
	) name413 (
		\ethreg1_IPGT_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_IPGT_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10926_
	);
	LUT4 #(
		.INIT('h8caf)
	) name414 (
		\ethreg1_IPGT_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_IPGT_0_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w10927_
	);
	LUT2 #(
		.INIT('h4)
	) name415 (
		_w10926_,
		_w10927_,
		_w10928_
	);
	LUT4 #(
		.INIT('h080a)
	) name416 (
		\ethreg1_IPGT_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_IPGT_0_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w10929_
	);
	LUT4 #(
		.INIT('hf531)
	) name417 (
		\ethreg1_IPGT_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_IPGT_0_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w10930_
	);
	LUT4 #(
		.INIT('h8caf)
	) name418 (
		\ethreg1_IPGT_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_IPGT_0_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10931_
	);
	LUT4 #(
		.INIT('h8a00)
	) name419 (
		_w10927_,
		_w10929_,
		_w10930_,
		_w10931_,
		_w10932_
	);
	LUT4 #(
		.INIT('hf531)
	) name420 (
		\ethreg1_IPGT_0_DataOut_reg[5]/NET0131 ,
		\ethreg1_IPGT_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w10933_
	);
	LUT2 #(
		.INIT('h8)
	) name421 (
		\txethmac1_txstatem1_StateIPG_reg/NET0131 ,
		_w10933_,
		_w10934_
	);
	LUT4 #(
		.INIT('h5455)
	) name422 (
		_w10925_,
		_w10928_,
		_w10932_,
		_w10934_,
		_w10935_
	);
	LUT3 #(
		.INIT('h80)
	) name423 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		_w10936_
	);
	LUT4 #(
		.INIT('h1000)
	) name424 (
		\maccontrol1_receivecontrol1_Pause_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w10937_
	);
	LUT3 #(
		.INIT('h54)
	) name425 (
		_w10779_,
		_w10936_,
		_w10937_,
		_w10938_
	);
	LUT4 #(
		.INIT('h00ae)
	) name426 (
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		_w10924_,
		_w10935_,
		_w10938_,
		_w10939_
	);
	LUT4 #(
		.INIT('h1000)
	) name427 (
		_w10607_,
		_w10726_,
		_w10815_,
		_w10939_,
		_w10940_
	);
	LUT4 #(
		.INIT('h0100)
	) name428 (
		\txethmac1_txstatem1_StateDefer_reg/NET0131 ,
		_w10607_,
		_w10726_,
		_w10815_,
		_w10941_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		_w10839_,
		_w10941_,
		_w10942_
	);
	LUT3 #(
		.INIT('h1b)
	) name430 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[3]_pad ,
		\mtxd_pad_o[3]_pad ,
		_w10943_
	);
	LUT3 #(
		.INIT('he4)
	) name431 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[3]_pad ,
		\mtxd_pad_o[3]_pad ,
		_w10944_
	);
	LUT4 #(
		.INIT('h1be4)
	) name432 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[3]_pad ,
		\mtxd_pad_o[3]_pad ,
		\rxethmac1_crcrx_Crc_reg[28]/NET0131 ,
		_w10945_
	);
	LUT2 #(
		.INIT('h6)
	) name433 (
		_w10580_,
		_w10945_,
		_w10946_
	);
	LUT3 #(
		.INIT('h14)
	) name434 (
		\rxethmac1_crcrx_Crc_reg[19]/NET0131 ,
		_w10580_,
		_w10945_,
		_w10947_
	);
	LUT4 #(
		.INIT('h7000)
	) name435 (
		_w10554_,
		_w10573_,
		_w10577_,
		_w10947_,
		_w10948_
	);
	LUT2 #(
		.INIT('h4)
	) name436 (
		\rxethmac1_crcrx_Crc_reg[19]/NET0131 ,
		_w10582_,
		_w10949_
	);
	LUT2 #(
		.INIT('h8)
	) name437 (
		_w10582_,
		_w10946_,
		_w10950_
	);
	LUT4 #(
		.INIT('h7000)
	) name438 (
		_w10554_,
		_w10573_,
		_w10577_,
		_w10950_,
		_w10951_
	);
	LUT3 #(
		.INIT('hab)
	) name439 (
		_w10948_,
		_w10949_,
		_w10951_,
		_w10952_
	);
	LUT2 #(
		.INIT('h9)
	) name440 (
		_w10580_,
		_w10590_,
		_w10953_
	);
	LUT3 #(
		.INIT('h14)
	) name441 (
		\rxethmac1_crcrx_Crc_reg[20]/NET0131 ,
		_w10580_,
		_w10590_,
		_w10954_
	);
	LUT4 #(
		.INIT('h7000)
	) name442 (
		_w10554_,
		_w10573_,
		_w10577_,
		_w10954_,
		_w10955_
	);
	LUT2 #(
		.INIT('h4)
	) name443 (
		\rxethmac1_crcrx_Crc_reg[20]/NET0131 ,
		_w10582_,
		_w10956_
	);
	LUT2 #(
		.INIT('h2)
	) name444 (
		_w10582_,
		_w10953_,
		_w10957_
	);
	LUT4 #(
		.INIT('h7000)
	) name445 (
		_w10554_,
		_w10573_,
		_w10577_,
		_w10957_,
		_w10958_
	);
	LUT3 #(
		.INIT('hab)
	) name446 (
		_w10955_,
		_w10956_,
		_w10958_,
		_w10959_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		\rxethmac1_crcrx_Crc_reg[26]/NET0131 ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w10960_
	);
	LUT4 #(
		.INIT('h02ff)
	) name448 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		_w10542_,
		_w10543_,
		_w10960_,
		_w10961_
	);
	LUT4 #(
		.INIT('h0001)
	) name449 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w10818_,
		_w10820_,
		_w10824_,
		_w10962_
	);
	LUT3 #(
		.INIT('h02)
	) name450 (
		_w10816_,
		_w10830_,
		_w10962_,
		_w10963_
	);
	LUT2 #(
		.INIT('h4)
	) name451 (
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w10826_,
		_w10964_
	);
	LUT4 #(
		.INIT('h1500)
	) name452 (
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w10801_,
		_w10828_,
		_w10965_
	);
	LUT2 #(
		.INIT('h8)
	) name453 (
		\txethmac1_ColWindow_reg/NET0131 ,
		_w10784_,
		_w10966_
	);
	LUT4 #(
		.INIT('h0888)
	) name454 (
		\txethmac1_ColWindow_reg/NET0131 ,
		_w10784_,
		_w10785_,
		_w10786_,
		_w10967_
	);
	LUT4 #(
		.INIT('h0103)
	) name455 (
		_w10791_,
		_w10964_,
		_w10965_,
		_w10967_,
		_w10968_
	);
	LUT4 #(
		.INIT('h1000)
	) name456 (
		_w10607_,
		_w10726_,
		_w10815_,
		_w10968_,
		_w10969_
	);
	LUT4 #(
		.INIT('h0001)
	) name457 (
		_w10818_,
		_w10820_,
		_w10824_,
		_w10830_,
		_w10970_
	);
	LUT4 #(
		.INIT('hfd00)
	) name458 (
		_w10664_,
		_w10691_,
		_w10722_,
		_w10724_,
		_w10971_
	);
	LUT3 #(
		.INIT('h10)
	) name459 (
		_w10600_,
		_w10603_,
		_w10605_,
		_w10972_
	);
	LUT3 #(
		.INIT('h45)
	) name460 (
		\txethmac1_txstatem1_StatePAD_reg/NET0131 ,
		_w10971_,
		_w10972_,
		_w10973_
	);
	LUT2 #(
		.INIT('h2)
	) name461 (
		_w10970_,
		_w10973_,
		_w10974_
	);
	LUT2 #(
		.INIT('h4)
	) name462 (
		\txethmac1_StopExcessiveDeferOccured_reg/NET0131 ,
		\txethmac1_txstatem1_StateDefer_reg/NET0131 ,
		_w10975_
	);
	LUT2 #(
		.INIT('h4)
	) name463 (
		_w10836_,
		_w10975_,
		_w10976_
	);
	LUT2 #(
		.INIT('h1)
	) name464 (
		\wishbone_TxUnderRun_reg/NET0131 ,
		_w10784_,
		_w10977_
	);
	LUT2 #(
		.INIT('h2)
	) name465 (
		\txethmac1_ColWindow_reg/NET0131 ,
		\wishbone_TxUnderRun_reg/NET0131 ,
		_w10978_
	);
	LUT3 #(
		.INIT('h70)
	) name466 (
		_w10785_,
		_w10786_,
		_w10978_,
		_w10979_
	);
	LUT4 #(
		.INIT('h7770)
	) name467 (
		_w10834_,
		_w10976_,
		_w10977_,
		_w10979_,
		_w10980_
	);
	LUT4 #(
		.INIT('h1500)
	) name468 (
		_w10729_,
		_w10744_,
		_w10756_,
		_w10980_,
		_w10981_
	);
	LUT2 #(
		.INIT('h4)
	) name469 (
		_w10791_,
		_w10966_,
		_w10982_
	);
	LUT3 #(
		.INIT('h56)
	) name470 (
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		_w10810_,
		_w10982_,
		_w10983_
	);
	LUT4 #(
		.INIT('h1000)
	) name471 (
		_w10607_,
		_w10726_,
		_w10981_,
		_w10983_,
		_w10984_
	);
	LUT2 #(
		.INIT('h8)
	) name472 (
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		_w10985_
	);
	LUT3 #(
		.INIT('h80)
	) name473 (
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		_w10986_
	);
	LUT4 #(
		.INIT('h56aa)
	) name474 (
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		_w10810_,
		_w10982_,
		_w10985_,
		_w10987_
	);
	LUT4 #(
		.INIT('h1000)
	) name475 (
		_w10607_,
		_w10726_,
		_w10981_,
		_w10987_,
		_w10988_
	);
	LUT4 #(
		.INIT('h0155)
	) name476 (
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w10810_,
		_w10982_,
		_w10986_,
		_w10989_
	);
	LUT4 #(
		.INIT('h8000)
	) name477 (
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w10990_
	);
	LUT3 #(
		.INIT('he0)
	) name478 (
		_w10810_,
		_w10982_,
		_w10990_,
		_w10991_
	);
	LUT2 #(
		.INIT('h1)
	) name479 (
		_w10989_,
		_w10991_,
		_w10992_
	);
	LUT4 #(
		.INIT('h1000)
	) name480 (
		_w10607_,
		_w10726_,
		_w10981_,
		_w10992_,
		_w10993_
	);
	LUT4 #(
		.INIT('h666c)
	) name481 (
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		_w10810_,
		_w10982_,
		_w10994_
	);
	LUT4 #(
		.INIT('h1000)
	) name482 (
		_w10607_,
		_w10726_,
		_w10981_,
		_w10994_,
		_w10995_
	);
	LUT2 #(
		.INIT('h4)
	) name483 (
		\maccontrol1_transmitcontrol1_ControlData_reg[7]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w10996_
	);
	LUT4 #(
		.INIT('h3020)
	) name484 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\wishbone_TxData_reg[7]/NET0131 ,
		_w10997_
	);
	LUT4 #(
		.INIT('hb080)
	) name485 (
		\maccontrol1_transmitcontrol1_ControlData_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		\wishbone_TxData_reg[3]/NET0131 ,
		_w10998_
	);
	LUT3 #(
		.INIT('h0b)
	) name486 (
		_w10996_,
		_w10997_,
		_w10998_,
		_w10999_
	);
	LUT4 #(
		.INIT('haa65)
	) name487 (
		\txethmac1_txcrc_Crc_reg[28]/NET0131 ,
		_w10996_,
		_w10997_,
		_w10998_,
		_w11000_
	);
	LUT2 #(
		.INIT('h4)
	) name488 (
		\maccontrol1_transmitcontrol1_ControlData_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w11001_
	);
	LUT4 #(
		.INIT('h3020)
	) name489 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\wishbone_TxData_reg[4]/NET0131 ,
		_w11002_
	);
	LUT4 #(
		.INIT('hb080)
	) name490 (
		\maccontrol1_transmitcontrol1_ControlData_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		\wishbone_TxData_reg[0]/NET0131 ,
		_w11003_
	);
	LUT3 #(
		.INIT('h0b)
	) name491 (
		_w11001_,
		_w11002_,
		_w11003_,
		_w11004_
	);
	LUT4 #(
		.INIT('h559a)
	) name492 (
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		_w11001_,
		_w11002_,
		_w11003_,
		_w11005_
	);
	LUT4 #(
		.INIT('h1001)
	) name493 (
		\txethmac1_txcrc_Crc_reg[22]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11000_,
		_w11005_,
		_w11006_
	);
	LUT2 #(
		.INIT('h8)
	) name494 (
		_w10913_,
		_w10914_,
		_w11007_
	);
	LUT3 #(
		.INIT('h40)
	) name495 (
		\txethmac1_txcrc_Crc_reg[22]/NET0131 ,
		_w10913_,
		_w10914_,
		_w11008_
	);
	LUT4 #(
		.INIT('h4100)
	) name496 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11000_,
		_w11005_,
		_w11007_,
		_w11009_
	);
	LUT3 #(
		.INIT('hab)
	) name497 (
		_w11006_,
		_w11008_,
		_w11009_,
		_w11010_
	);
	LUT4 #(
		.INIT('hb080)
	) name498 (
		\maccontrol1_transmitcontrol1_ControlData_reg[2]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		\wishbone_TxData_reg[2]/NET0131 ,
		_w11011_
	);
	LUT2 #(
		.INIT('h4)
	) name499 (
		\maccontrol1_transmitcontrol1_ControlData_reg[6]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w11012_
	);
	LUT4 #(
		.INIT('h3020)
	) name500 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\wishbone_TxData_reg[6]/NET0131 ,
		_w11013_
	);
	LUT3 #(
		.INIT('h45)
	) name501 (
		_w11011_,
		_w11012_,
		_w11013_,
		_w11014_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11015_
	);
	LUT4 #(
		.INIT('hba00)
	) name503 (
		_w11011_,
		_w11012_,
		_w11013_,
		_w11015_,
		_w11016_
	);
	LUT2 #(
		.INIT('h2)
	) name504 (
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11017_
	);
	LUT4 #(
		.INIT('h4500)
	) name505 (
		_w11011_,
		_w11012_,
		_w11013_,
		_w11017_,
		_w11018_
	);
	LUT3 #(
		.INIT('h02)
	) name506 (
		\txethmac1_txcrc_Crc_reg[23]/NET0131 ,
		_w11016_,
		_w11018_,
		_w11019_
	);
	LUT3 #(
		.INIT('h01)
	) name507 (
		\txethmac1_txcrc_Crc_reg[23]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11020_
	);
	LUT4 #(
		.INIT('hba00)
	) name508 (
		_w11011_,
		_w11012_,
		_w11013_,
		_w11020_,
		_w11021_
	);
	LUT3 #(
		.INIT('h04)
	) name509 (
		\txethmac1_txcrc_Crc_reg[23]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11022_
	);
	LUT4 #(
		.INIT('h4500)
	) name510 (
		_w11011_,
		_w11012_,
		_w11013_,
		_w11022_,
		_w11023_
	);
	LUT3 #(
		.INIT('h02)
	) name511 (
		_w11007_,
		_w11021_,
		_w11023_,
		_w11024_
	);
	LUT2 #(
		.INIT('hb)
	) name512 (
		_w11019_,
		_w11024_,
		_w11025_
	);
	LUT3 #(
		.INIT('hc8)
	) name513 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\wishbone_TxData_reg[5]/NET0131 ,
		_w11026_
	);
	LUT3 #(
		.INIT('h0b)
	) name514 (
		\maccontrol1_transmitcontrol1_ControlData_reg[5]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		_w11027_
	);
	LUT4 #(
		.INIT('hb080)
	) name515 (
		\maccontrol1_transmitcontrol1_ControlData_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		\wishbone_TxData_reg[1]/NET0131 ,
		_w11028_
	);
	LUT2 #(
		.INIT('h1)
	) name516 (
		\txethmac1_txcrc_Crc_reg[30]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11029_
	);
	LUT4 #(
		.INIT('hf800)
	) name517 (
		_w11026_,
		_w11027_,
		_w11028_,
		_w11029_,
		_w11030_
	);
	LUT2 #(
		.INIT('h2)
	) name518 (
		\txethmac1_txcrc_Crc_reg[30]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11031_
	);
	LUT4 #(
		.INIT('h0700)
	) name519 (
		_w11026_,
		_w11027_,
		_w11028_,
		_w11031_,
		_w11032_
	);
	LUT3 #(
		.INIT('h02)
	) name520 (
		\txethmac1_txcrc_Crc_reg[24]/NET0131 ,
		_w11030_,
		_w11032_,
		_w11033_
	);
	LUT3 #(
		.INIT('h01)
	) name521 (
		\txethmac1_txcrc_Crc_reg[24]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[30]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11034_
	);
	LUT4 #(
		.INIT('hf800)
	) name522 (
		_w11026_,
		_w11027_,
		_w11028_,
		_w11034_,
		_w11035_
	);
	LUT3 #(
		.INIT('h04)
	) name523 (
		\txethmac1_txcrc_Crc_reg[24]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[30]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11036_
	);
	LUT4 #(
		.INIT('h0700)
	) name524 (
		_w11026_,
		_w11027_,
		_w11028_,
		_w11036_,
		_w11037_
	);
	LUT3 #(
		.INIT('h02)
	) name525 (
		_w11007_,
		_w11035_,
		_w11037_,
		_w11038_
	);
	LUT2 #(
		.INIT('hb)
	) name526 (
		_w11033_,
		_w11038_,
		_w11039_
	);
	LUT3 #(
		.INIT('h45)
	) name527 (
		\txethmac1_txstatem1_StateIPG_reg/NET0131 ,
		_w10834_,
		_w10838_,
		_w11040_
	);
	LUT3 #(
		.INIT('h0d)
	) name528 (
		_w10924_,
		_w10935_,
		_w11040_,
		_w11041_
	);
	LUT4 #(
		.INIT('h1000)
	) name529 (
		_w10607_,
		_w10726_,
		_w10815_,
		_w11041_,
		_w11042_
	);
	LUT3 #(
		.INIT('h15)
	) name530 (
		\txethmac1_txstatem1_StateBackOff_reg/NET0131 ,
		_w10791_,
		_w10967_,
		_w11043_
	);
	LUT4 #(
		.INIT('h0010)
	) name531 (
		_w10607_,
		_w10726_,
		_w10815_,
		_w11043_,
		_w11044_
	);
	LUT3 #(
		.INIT('h1b)
	) name532 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[0]_pad ,
		\mtxd_pad_o[0]_pad ,
		_w11045_
	);
	LUT3 #(
		.INIT('he4)
	) name533 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[0]_pad ,
		\mtxd_pad_o[0]_pad ,
		_w11046_
	);
	LUT4 #(
		.INIT('h1be4)
	) name534 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[0]_pad ,
		\mtxd_pad_o[0]_pad ,
		\rxethmac1_crcrx_Crc_reg[31]/NET0131 ,
		_w11047_
	);
	LUT2 #(
		.INIT('h9)
	) name535 (
		_w10945_,
		_w11047_,
		_w11048_
	);
	LUT4 #(
		.INIT('h0070)
	) name536 (
		_w10554_,
		_w10573_,
		_w10577_,
		_w11048_,
		_w11049_
	);
	LUT3 #(
		.INIT('h7b)
	) name537 (
		\rxethmac1_crcrx_Crc_reg[22]/NET0131 ,
		_w10582_,
		_w11049_,
		_w11050_
	);
	LUT2 #(
		.INIT('h2)
	) name538 (
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11051_
	);
	LUT4 #(
		.INIT('h0b00)
	) name539 (
		_w11001_,
		_w11002_,
		_w11003_,
		_w11051_,
		_w11052_
	);
	LUT2 #(
		.INIT('h1)
	) name540 (
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11053_
	);
	LUT4 #(
		.INIT('hf400)
	) name541 (
		_w11001_,
		_w11002_,
		_w11003_,
		_w11053_,
		_w11054_
	);
	LUT3 #(
		.INIT('h02)
	) name542 (
		\txethmac1_txcrc_Crc_reg[25]/NET0131 ,
		_w11052_,
		_w11054_,
		_w11055_
	);
	LUT3 #(
		.INIT('h01)
	) name543 (
		\txethmac1_txcrc_Crc_reg[25]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11056_
	);
	LUT4 #(
		.INIT('hf400)
	) name544 (
		_w11001_,
		_w11002_,
		_w11003_,
		_w11056_,
		_w11057_
	);
	LUT3 #(
		.INIT('h04)
	) name545 (
		\txethmac1_txcrc_Crc_reg[25]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11058_
	);
	LUT4 #(
		.INIT('h0b00)
	) name546 (
		_w11001_,
		_w11002_,
		_w11003_,
		_w11058_,
		_w11059_
	);
	LUT3 #(
		.INIT('h02)
	) name547 (
		_w11007_,
		_w11057_,
		_w11059_,
		_w11060_
	);
	LUT2 #(
		.INIT('hb)
	) name548 (
		_w11055_,
		_w11060_,
		_w11061_
	);
	LUT3 #(
		.INIT('h07)
	) name549 (
		_w10744_,
		_w10756_,
		_w10825_,
		_w11062_
	);
	LUT3 #(
		.INIT('hf8)
	) name550 (
		_w10744_,
		_w10756_,
		_w10825_,
		_w11063_
	);
	LUT3 #(
		.INIT('h80)
	) name551 (
		\txethmac1_ColWindow_reg/NET0131 ,
		_w10785_,
		_w10786_,
		_w11064_
	);
	LUT2 #(
		.INIT('h8)
	) name552 (
		_w10830_,
		_w11064_,
		_w11065_
	);
	LUT3 #(
		.INIT('h01)
	) name553 (
		\txethmac1_ColWindow_reg/NET0131 ,
		_w10825_,
		_w10826_,
		_w11066_
	);
	LUT2 #(
		.INIT('h4)
	) name554 (
		_w10829_,
		_w11066_,
		_w11067_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name555 (
		_w10829_,
		_w10834_,
		_w10976_,
		_w11066_,
		_w11068_
	);
	LUT2 #(
		.INIT('h4)
	) name556 (
		_w11065_,
		_w11068_,
		_w11069_
	);
	LUT3 #(
		.INIT('h40)
	) name557 (
		_w10729_,
		_w11062_,
		_w11069_,
		_w11070_
	);
	LUT3 #(
		.INIT('hef)
	) name558 (
		_w10607_,
		_w10726_,
		_w11070_,
		_w11071_
	);
	LUT3 #(
		.INIT('h15)
	) name559 (
		\txethmac1_TxDone_reg/NET0131 ,
		_w10727_,
		_w10728_,
		_w11072_
	);
	LUT3 #(
		.INIT('h08)
	) name560 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		\txethmac1_StatusLatch_reg/NET0131 ,
		_w11073_
	);
	LUT4 #(
		.INIT('h0100)
	) name561 (
		\maccontrol1_receivecontrol1_Pause_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_StatusLatch_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w11074_
	);
	LUT2 #(
		.INIT('h1)
	) name562 (
		_w11073_,
		_w11074_,
		_w11075_
	);
	LUT4 #(
		.INIT('hef00)
	) name563 (
		_w10607_,
		_w10726_,
		_w11072_,
		_w11075_,
		_w11076_
	);
	LUT2 #(
		.INIT('h4)
	) name564 (
		\ethreg1_ResetTxCIrq_sync2_reg/NET0131 ,
		\ethreg1_SetTxCIrq_txclk_reg/NET0131 ,
		_w11077_
	);
	LUT4 #(
		.INIT('h45cf)
	) name565 (
		\ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_ResetTxCIrq_sync2_reg/NET0131 ,
		\ethreg1_SetTxCIrq_txclk_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_TxCtrlEndFrm_reg/NET0131 ,
		_w11078_
	);
	LUT3 #(
		.INIT('h07)
	) name566 (
		_w10727_,
		_w10728_,
		_w11077_,
		_w11079_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name567 (
		_w10607_,
		_w10726_,
		_w11078_,
		_w11079_,
		_w11080_
	);
	LUT3 #(
		.INIT('h10)
	) name568 (
		_w10574_,
		_w10576_,
		_w11047_,
		_w11081_
	);
	LUT2 #(
		.INIT('h4)
	) name569 (
		\rxethmac1_crcrx_Crc_reg[15]/NET0131 ,
		_w10582_,
		_w11082_
	);
	LUT4 #(
		.INIT('h8f00)
	) name570 (
		_w10554_,
		_w10573_,
		_w11081_,
		_w11082_,
		_w11083_
	);
	LUT2 #(
		.INIT('h8)
	) name571 (
		\rxethmac1_crcrx_Crc_reg[15]/NET0131 ,
		_w10582_,
		_w11084_
	);
	LUT4 #(
		.INIT('h7000)
	) name572 (
		_w10554_,
		_w10573_,
		_w11081_,
		_w11084_,
		_w11085_
	);
	LUT2 #(
		.INIT('h1)
	) name573 (
		_w11083_,
		_w11085_,
		_w11086_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		\rxethmac1_crcrx_Crc_reg[16]/NET0131 ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w11087_
	);
	LUT4 #(
		.INIT('h02ff)
	) name575 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		_w10542_,
		_w10543_,
		_w11087_,
		_w11088_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		\txethmac1_txcrc_Crc_reg[28]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11089_
	);
	LUT4 #(
		.INIT('hf400)
	) name577 (
		_w10996_,
		_w10997_,
		_w10998_,
		_w11089_,
		_w11090_
	);
	LUT2 #(
		.INIT('h2)
	) name578 (
		\txethmac1_txcrc_Crc_reg[28]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11091_
	);
	LUT4 #(
		.INIT('h0b00)
	) name579 (
		_w10996_,
		_w10997_,
		_w10998_,
		_w11091_,
		_w11092_
	);
	LUT3 #(
		.INIT('h02)
	) name580 (
		\txethmac1_txcrc_Crc_reg[18]/NET0131 ,
		_w11090_,
		_w11092_,
		_w11093_
	);
	LUT3 #(
		.INIT('h01)
	) name581 (
		\txethmac1_txcrc_Crc_reg[18]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[28]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11094_
	);
	LUT4 #(
		.INIT('hf400)
	) name582 (
		_w10996_,
		_w10997_,
		_w10998_,
		_w11094_,
		_w11095_
	);
	LUT3 #(
		.INIT('h04)
	) name583 (
		\txethmac1_txcrc_Crc_reg[18]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[28]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11096_
	);
	LUT4 #(
		.INIT('h0b00)
	) name584 (
		_w10996_,
		_w10997_,
		_w10998_,
		_w11096_,
		_w11097_
	);
	LUT3 #(
		.INIT('h02)
	) name585 (
		_w11007_,
		_w11095_,
		_w11097_,
		_w11098_
	);
	LUT2 #(
		.INIT('hb)
	) name586 (
		_w11093_,
		_w11098_,
		_w11099_
	);
	LUT2 #(
		.INIT('h9)
	) name587 (
		\txethmac1_txcrc_Crc_reg[28]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		_w11100_
	);
	LUT4 #(
		.INIT('hebbe)
	) name588 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w10999_,
		_w11014_,
		_w11100_,
		_w11101_
	);
	LUT2 #(
		.INIT('h1)
	) name589 (
		\txethmac1_txcrc_Crc_reg[19]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11102_
	);
	LUT4 #(
		.INIT('h96ff)
	) name590 (
		_w10999_,
		_w11014_,
		_w11100_,
		_w11102_,
		_w11103_
	);
	LUT4 #(
		.INIT('hb3ff)
	) name591 (
		\txethmac1_txcrc_Crc_reg[19]/NET0131 ,
		_w11007_,
		_w11101_,
		_w11103_,
		_w11104_
	);
	LUT4 #(
		.INIT('h6566)
	) name592 (
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		_w11011_,
		_w11012_,
		_w11013_,
		_w11105_
	);
	LUT4 #(
		.INIT('h556a)
	) name593 (
		\txethmac1_txcrc_Crc_reg[30]/NET0131 ,
		_w11026_,
		_w11027_,
		_w11028_,
		_w11106_
	);
	LUT2 #(
		.INIT('h1)
	) name594 (
		\txethmac1_txcrc_Crc_reg[20]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11107_
	);
	LUT3 #(
		.INIT('h60)
	) name595 (
		_w11105_,
		_w11106_,
		_w11107_,
		_w11108_
	);
	LUT3 #(
		.INIT('h40)
	) name596 (
		\txethmac1_txcrc_Crc_reg[20]/NET0131 ,
		_w10913_,
		_w10914_,
		_w11109_
	);
	LUT3 #(
		.INIT('h40)
	) name597 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w10913_,
		_w10914_,
		_w11110_
	);
	LUT4 #(
		.INIT('h090f)
	) name598 (
		_w11105_,
		_w11106_,
		_w11109_,
		_w11110_,
		_w11111_
	);
	LUT2 #(
		.INIT('he)
	) name599 (
		_w11108_,
		_w11111_,
		_w11112_
	);
	LUT3 #(
		.INIT('h10)
	) name600 (
		_w10574_,
		_w10576_,
		_w10945_,
		_w11113_
	);
	LUT2 #(
		.INIT('h4)
	) name601 (
		\rxethmac1_crcrx_Crc_reg[12]/NET0131 ,
		_w10582_,
		_w11114_
	);
	LUT4 #(
		.INIT('h8f00)
	) name602 (
		_w10554_,
		_w10573_,
		_w11113_,
		_w11114_,
		_w11115_
	);
	LUT2 #(
		.INIT('h8)
	) name603 (
		\rxethmac1_crcrx_Crc_reg[12]/NET0131 ,
		_w10582_,
		_w11116_
	);
	LUT4 #(
		.INIT('h7000)
	) name604 (
		_w10554_,
		_w10573_,
		_w11113_,
		_w11116_,
		_w11117_
	);
	LUT2 #(
		.INIT('h1)
	) name605 (
		_w11115_,
		_w11117_,
		_w11118_
	);
	LUT2 #(
		.INIT('h4)
	) name606 (
		\rxethmac1_crcrx_Crc_reg[18]/NET0131 ,
		_w10582_,
		_w11119_
	);
	LUT4 #(
		.INIT('h8f00)
	) name607 (
		_w10554_,
		_w10573_,
		_w11113_,
		_w11119_,
		_w11120_
	);
	LUT2 #(
		.INIT('h8)
	) name608 (
		\rxethmac1_crcrx_Crc_reg[18]/NET0131 ,
		_w10582_,
		_w11121_
	);
	LUT4 #(
		.INIT('h7000)
	) name609 (
		_w10554_,
		_w10573_,
		_w11113_,
		_w11121_,
		_w11122_
	);
	LUT2 #(
		.INIT('h1)
	) name610 (
		_w11120_,
		_w11122_,
		_w11123_
	);
	LUT4 #(
		.INIT('h0110)
	) name611 (
		\txethmac1_txcrc_Crc_reg[21]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11005_,
		_w11106_,
		_w11124_
	);
	LUT3 #(
		.INIT('h40)
	) name612 (
		\txethmac1_txcrc_Crc_reg[21]/NET0131 ,
		_w10913_,
		_w10914_,
		_w11125_
	);
	LUT4 #(
		.INIT('h1040)
	) name613 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11005_,
		_w11007_,
		_w11106_,
		_w11126_
	);
	LUT3 #(
		.INIT('hab)
	) name614 (
		_w11124_,
		_w11125_,
		_w11126_,
		_w11127_
	);
	LUT2 #(
		.INIT('h4)
	) name615 (
		\rxethmac1_crcrx_Crc_reg[11]/NET0131 ,
		_w10582_,
		_w11128_
	);
	LUT4 #(
		.INIT('h8f00)
	) name616 (
		_w10554_,
		_w10573_,
		_w11081_,
		_w11128_,
		_w11129_
	);
	LUT2 #(
		.INIT('h8)
	) name617 (
		\rxethmac1_crcrx_Crc_reg[11]/NET0131 ,
		_w10582_,
		_w11130_
	);
	LUT4 #(
		.INIT('h7000)
	) name618 (
		_w10554_,
		_w10573_,
		_w11081_,
		_w11130_,
		_w11131_
	);
	LUT2 #(
		.INIT('h1)
	) name619 (
		_w11129_,
		_w11131_,
		_w11132_
	);
	LUT3 #(
		.INIT('hd0)
	) name620 (
		\ethreg1_ResetRxCIrq_sync2_reg/NET0131 ,
		\ethreg1_ResetRxCIrq_sync3_reg/NET0131 ,
		\ethreg1_SetRxCIrq_rxclk_reg/NET0131 ,
		_w11133_
	);
	LUT2 #(
		.INIT('h8)
	) name621 (
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w11134_
	);
	LUT4 #(
		.INIT('h8000)
	) name622 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		_w11135_
	);
	LUT3 #(
		.INIT('h80)
	) name623 (
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		_w11136_
	);
	LUT3 #(
		.INIT('h80)
	) name624 (
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w11137_
	);
	LUT3 #(
		.INIT('h80)
	) name625 (
		_w11135_,
		_w11136_,
		_w11137_,
		_w11138_
	);
	LUT3 #(
		.INIT('h80)
	) name626 (
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		_w11139_
	);
	LUT4 #(
		.INIT('h8000)
	) name627 (
		_w11135_,
		_w11136_,
		_w11137_,
		_w11139_,
		_w11140_
	);
	LUT4 #(
		.INIT('h7df5)
	) name628 (
		\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		_w11140_,
		_w11141_
	);
	LUT4 #(
		.INIT('h1450)
	) name629 (
		\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		_w11140_,
		_w11142_
	);
	LUT3 #(
		.INIT('h7d)
	) name630 (
		\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		_w11140_,
		_w11143_
	);
	LUT2 #(
		.INIT('h1)
	) name631 (
		_w11142_,
		_w11143_,
		_w11144_
	);
	LUT4 #(
		.INIT('h8000)
	) name632 (
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11137_,
		_w11145_
	);
	LUT2 #(
		.INIT('h8)
	) name633 (
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		_w11146_
	);
	LUT4 #(
		.INIT('h8000)
	) name634 (
		_w11135_,
		_w11136_,
		_w11137_,
		_w11146_,
		_w11147_
	);
	LUT4 #(
		.INIT('h1450)
	) name635 (
		\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		_w11138_,
		_w11148_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name636 (
		_w10563_,
		_w11135_,
		_w11136_,
		_w11137_,
		_w11149_
	);
	LUT2 #(
		.INIT('h1)
	) name637 (
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w11150_
	);
	LUT4 #(
		.INIT('h8000)
	) name638 (
		_w11135_,
		_w11136_,
		_w11137_,
		_w11150_,
		_w11151_
	);
	LUT2 #(
		.INIT('h1)
	) name639 (
		_w11149_,
		_w11151_,
		_w11152_
	);
	LUT3 #(
		.INIT('h7d)
	) name640 (
		\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		_w11147_,
		_w11153_
	);
	LUT3 #(
		.INIT('h7d)
	) name641 (
		\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		_w11145_,
		_w11154_
	);
	LUT4 #(
		.INIT('hb000)
	) name642 (
		_w11148_,
		_w11152_,
		_w11153_,
		_w11154_,
		_w11155_
	);
	LUT4 #(
		.INIT('h7ddd)
	) name643 (
		\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11156_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name644 (
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w10561_,
		_w11135_,
		_w11136_,
		_w11157_
	);
	LUT2 #(
		.INIT('h8)
	) name645 (
		\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w11158_
	);
	LUT4 #(
		.INIT('h8000)
	) name646 (
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11158_,
		_w11159_
	);
	LUT3 #(
		.INIT('h02)
	) name647 (
		_w11156_,
		_w11157_,
		_w11159_,
		_w11160_
	);
	LUT2 #(
		.INIT('h8)
	) name648 (
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w11161_
	);
	LUT4 #(
		.INIT('h1555)
	) name649 (
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11161_,
		_w11162_
	);
	LUT4 #(
		.INIT('h1555)
	) name650 (
		\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11137_,
		_w11163_
	);
	LUT4 #(
		.INIT('h1333)
	) name651 (
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11164_
	);
	LUT4 #(
		.INIT('h1555)
	) name652 (
		\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11161_,
		_w11165_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name653 (
		_w11162_,
		_w11163_,
		_w11164_,
		_w11165_,
		_w11166_
	);
	LUT2 #(
		.INIT('h4)
	) name654 (
		_w11160_,
		_w11166_,
		_w11167_
	);
	LUT2 #(
		.INIT('h8)
	) name655 (
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		_w11168_
	);
	LUT4 #(
		.INIT('h1450)
	) name656 (
		\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		_w11135_,
		_w11169_
	);
	LUT3 #(
		.INIT('heb)
	) name657 (
		\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w11135_,
		_w11170_
	);
	LUT4 #(
		.INIT('h7ddd)
	) name658 (
		\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		_w11135_,
		_w11168_,
		_w11171_
	);
	LUT4 #(
		.INIT('h7df5)
	) name659 (
		\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		_w11135_,
		_w11172_
	);
	LUT4 #(
		.INIT('hb000)
	) name660 (
		_w11169_,
		_w11170_,
		_w11171_,
		_w11172_,
		_w11173_
	);
	LUT2 #(
		.INIT('h6)
	) name661 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		_w11174_
	);
	LUT3 #(
		.INIT('h31)
	) name662 (
		\ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w11175_
	);
	LUT3 #(
		.INIT('h23)
	) name663 (
		_w10555_,
		_w11174_,
		_w11175_,
		_w11176_
	);
	LUT3 #(
		.INIT('h80)
	) name664 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w11177_
	);
	LUT3 #(
		.INIT('h78)
	) name665 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w11178_
	);
	LUT4 #(
		.INIT('h804c)
	) name666 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w11179_
	);
	LUT4 #(
		.INIT('h7310)
	) name667 (
		\ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w11180_
	);
	LUT3 #(
		.INIT('h31)
	) name668 (
		\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 ,
		_w11179_,
		_w11180_,
		_w11181_
	);
	LUT4 #(
		.INIT('h007f)
	) name669 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		_w11182_
	);
	LUT4 #(
		.INIT('h1320)
	) name670 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w11183_
	);
	LUT4 #(
		.INIT('h00fe)
	) name671 (
		\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 ,
		_w11135_,
		_w11182_,
		_w11183_,
		_w11184_
	);
	LUT3 #(
		.INIT('hb0)
	) name672 (
		_w11176_,
		_w11181_,
		_w11184_,
		_w11185_
	);
	LUT3 #(
		.INIT('h7d)
	) name673 (
		\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w11135_,
		_w11186_
	);
	LUT3 #(
		.INIT('h7d)
	) name674 (
		\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		_w11177_,
		_w11187_
	);
	LUT4 #(
		.INIT('h8000)
	) name675 (
		_w11171_,
		_w11172_,
		_w11186_,
		_w11187_,
		_w11188_
	);
	LUT3 #(
		.INIT('h45)
	) name676 (
		_w11173_,
		_w11185_,
		_w11188_,
		_w11189_
	);
	LUT3 #(
		.INIT('h15)
	) name677 (
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		_w11135_,
		_w11168_,
		_w11190_
	);
	LUT3 #(
		.INIT('h15)
	) name678 (
		\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11191_
	);
	LUT4 #(
		.INIT('hebbb)
	) name679 (
		\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11192_
	);
	LUT3 #(
		.INIT('hb0)
	) name680 (
		_w11190_,
		_w11191_,
		_w11192_,
		_w11193_
	);
	LUT2 #(
		.INIT('h8)
	) name681 (
		_w11166_,
		_w11193_,
		_w11194_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name682 (
		_w10556_,
		_w11135_,
		_w11136_,
		_w11161_,
		_w11195_
	);
	LUT2 #(
		.INIT('h8)
	) name683 (
		\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		_w11196_
	);
	LUT4 #(
		.INIT('h8000)
	) name684 (
		_w11135_,
		_w11136_,
		_w11161_,
		_w11196_,
		_w11197_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name685 (
		_w10565_,
		_w11135_,
		_w11136_,
		_w11137_,
		_w11198_
	);
	LUT2 #(
		.INIT('h8)
	) name686 (
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w11199_
	);
	LUT4 #(
		.INIT('h8000)
	) name687 (
		_w11135_,
		_w11136_,
		_w11137_,
		_w11199_,
		_w11200_
	);
	LUT4 #(
		.INIT('h0001)
	) name688 (
		_w11195_,
		_w11197_,
		_w11198_,
		_w11200_,
		_w11201_
	);
	LUT3 #(
		.INIT('h80)
	) name689 (
		_w11153_,
		_w11154_,
		_w11201_,
		_w11202_
	);
	LUT4 #(
		.INIT('h1500)
	) name690 (
		_w11167_,
		_w11189_,
		_w11194_,
		_w11202_,
		_w11203_
	);
	LUT4 #(
		.INIT('h0504)
	) name691 (
		\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		_w11140_,
		_w11147_,
		_w11204_
	);
	LUT3 #(
		.INIT('heb)
	) name692 (
		\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		_w11140_,
		_w11205_
	);
	LUT3 #(
		.INIT('h10)
	) name693 (
		_w11142_,
		_w11204_,
		_w11205_,
		_w11206_
	);
	LUT4 #(
		.INIT('h5455)
	) name694 (
		_w11144_,
		_w11155_,
		_w11203_,
		_w11206_,
		_w11207_
	);
	LUT4 #(
		.INIT('h7df5)
	) name695 (
		\ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		_w11140_,
		_w11208_
	);
	LUT3 #(
		.INIT('h7d)
	) name696 (
		\ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		_w11140_,
		_w11209_
	);
	LUT3 #(
		.INIT('h7d)
	) name697 (
		\ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		_w11147_,
		_w11210_
	);
	LUT3 #(
		.INIT('h80)
	) name698 (
		_w11208_,
		_w11209_,
		_w11210_,
		_w11211_
	);
	LUT4 #(
		.INIT('h1450)
	) name699 (
		\ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		_w11140_,
		_w11212_
	);
	LUT3 #(
		.INIT('heb)
	) name700 (
		\ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		_w11140_,
		_w11213_
	);
	LUT3 #(
		.INIT('h31)
	) name701 (
		_w11208_,
		_w11212_,
		_w11213_,
		_w11214_
	);
	LUT2 #(
		.INIT('h4)
	) name702 (
		_w11211_,
		_w11214_,
		_w11215_
	);
	LUT2 #(
		.INIT('h4)
	) name703 (
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w11216_
	);
	LUT4 #(
		.INIT('h7f00)
	) name704 (
		_w11135_,
		_w11136_,
		_w11137_,
		_w11216_,
		_w11217_
	);
	LUT2 #(
		.INIT('h1)
	) name705 (
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w11218_
	);
	LUT4 #(
		.INIT('h8000)
	) name706 (
		_w11135_,
		_w11136_,
		_w11137_,
		_w11218_,
		_w11219_
	);
	LUT4 #(
		.INIT('h1555)
	) name707 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11137_,
		_w11220_
	);
	LUT4 #(
		.INIT('h0203)
	) name708 (
		_w11162_,
		_w11217_,
		_w11219_,
		_w11220_,
		_w11221_
	);
	LUT2 #(
		.INIT('h2)
	) name709 (
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w11222_
	);
	LUT4 #(
		.INIT('h7f00)
	) name710 (
		_w11135_,
		_w11136_,
		_w11137_,
		_w11222_,
		_w11223_
	);
	LUT2 #(
		.INIT('h8)
	) name711 (
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w11224_
	);
	LUT4 #(
		.INIT('h8000)
	) name712 (
		_w11135_,
		_w11136_,
		_w11137_,
		_w11224_,
		_w11225_
	);
	LUT2 #(
		.INIT('h1)
	) name713 (
		_w11223_,
		_w11225_,
		_w11226_
	);
	LUT3 #(
		.INIT('h7d)
	) name714 (
		\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		_w11145_,
		_w11227_
	);
	LUT3 #(
		.INIT('h40)
	) name715 (
		_w11221_,
		_w11226_,
		_w11227_,
		_w11228_
	);
	LUT4 #(
		.INIT('h7ddd)
	) name716 (
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11229_
	);
	LUT4 #(
		.INIT('hebbb)
	) name717 (
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11230_
	);
	LUT4 #(
		.INIT('h1555)
	) name718 (
		\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11161_,
		_w11231_
	);
	LUT3 #(
		.INIT('h8c)
	) name719 (
		_w11164_,
		_w11230_,
		_w11231_,
		_w11232_
	);
	LUT4 #(
		.INIT('h2030)
	) name720 (
		_w11164_,
		_w11229_,
		_w11230_,
		_w11231_,
		_w11233_
	);
	LUT3 #(
		.INIT('heb)
	) name721 (
		\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w11135_,
		_w11234_
	);
	LUT4 #(
		.INIT('h1450)
	) name722 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		_w11135_,
		_w11235_
	);
	LUT4 #(
		.INIT('h7ddd)
	) name723 (
		\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		_w11135_,
		_w11168_,
		_w11236_
	);
	LUT4 #(
		.INIT('h7df5)
	) name724 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		_w11135_,
		_w11237_
	);
	LUT4 #(
		.INIT('hd000)
	) name725 (
		_w11234_,
		_w11235_,
		_w11236_,
		_w11237_,
		_w11238_
	);
	LUT4 #(
		.INIT('h08ce)
	) name726 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w11239_
	);
	LUT4 #(
		.INIT('h804c)
	) name727 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w11240_
	);
	LUT4 #(
		.INIT('h004d)
	) name728 (
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		_w11174_,
		_w11239_,
		_w11240_,
		_w11241_
	);
	LUT4 #(
		.INIT('h1320)
	) name729 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w11242_
	);
	LUT4 #(
		.INIT('h00fe)
	) name730 (
		\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 ,
		_w11135_,
		_w11182_,
		_w11242_,
		_w11243_
	);
	LUT2 #(
		.INIT('h4)
	) name731 (
		_w11241_,
		_w11243_,
		_w11244_
	);
	LUT3 #(
		.INIT('h7d)
	) name732 (
		\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w11135_,
		_w11245_
	);
	LUT3 #(
		.INIT('h7d)
	) name733 (
		\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		_w11177_,
		_w11246_
	);
	LUT4 #(
		.INIT('h8000)
	) name734 (
		_w11236_,
		_w11237_,
		_w11245_,
		_w11246_,
		_w11247_
	);
	LUT3 #(
		.INIT('h45)
	) name735 (
		_w11238_,
		_w11244_,
		_w11247_,
		_w11248_
	);
	LUT3 #(
		.INIT('h15)
	) name736 (
		\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11249_
	);
	LUT2 #(
		.INIT('h4)
	) name737 (
		_w11190_,
		_w11249_,
		_w11250_
	);
	LUT2 #(
		.INIT('h2)
	) name738 (
		_w11232_,
		_w11250_,
		_w11251_
	);
	LUT2 #(
		.INIT('h2)
	) name739 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		_w11252_
	);
	LUT4 #(
		.INIT('h7f00)
	) name740 (
		_w11135_,
		_w11136_,
		_w11161_,
		_w11252_,
		_w11253_
	);
	LUT2 #(
		.INIT('h8)
	) name741 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		_w11254_
	);
	LUT4 #(
		.INIT('h8000)
	) name742 (
		_w11135_,
		_w11136_,
		_w11161_,
		_w11254_,
		_w11255_
	);
	LUT2 #(
		.INIT('h2)
	) name743 (
		\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w11256_
	);
	LUT4 #(
		.INIT('h7f00)
	) name744 (
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11256_,
		_w11257_
	);
	LUT2 #(
		.INIT('h8)
	) name745 (
		\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w11258_
	);
	LUT4 #(
		.INIT('h8000)
	) name746 (
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w11135_,
		_w11136_,
		_w11258_,
		_w11259_
	);
	LUT4 #(
		.INIT('h0001)
	) name747 (
		_w11253_,
		_w11255_,
		_w11257_,
		_w11259_,
		_w11260_
	);
	LUT3 #(
		.INIT('h80)
	) name748 (
		_w11226_,
		_w11227_,
		_w11260_,
		_w11261_
	);
	LUT4 #(
		.INIT('h1500)
	) name749 (
		_w11233_,
		_w11248_,
		_w11251_,
		_w11261_,
		_w11262_
	);
	LUT4 #(
		.INIT('h0504)
	) name750 (
		\ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		_w11140_,
		_w11147_,
		_w11263_
	);
	LUT4 #(
		.INIT('h1450)
	) name751 (
		\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		_w11138_,
		_w11264_
	);
	LUT2 #(
		.INIT('h1)
	) name752 (
		_w11263_,
		_w11264_,
		_w11265_
	);
	LUT2 #(
		.INIT('h8)
	) name753 (
		_w11214_,
		_w11265_,
		_w11266_
	);
	LUT4 #(
		.INIT('h5455)
	) name754 (
		_w11215_,
		_w11228_,
		_w11262_,
		_w11266_,
		_w11267_
	);
	LUT4 #(
		.INIT('h0800)
	) name755 (
		\ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		\macstatus1_LatchedCrcError_reg/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w11268_
	);
	LUT4 #(
		.INIT('h7000)
	) name756 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11268_,
		_w11269_
	);
	LUT2 #(
		.INIT('he)
	) name757 (
		_w11133_,
		_w11269_,
		_w11270_
	);
	LUT2 #(
		.INIT('h1)
	) name758 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[11]/NET0131 ,
		_w11271_
	);
	LUT4 #(
		.INIT('h0001)
	) name759 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[12]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[14]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131 ,
		_w11272_
	);
	LUT2 #(
		.INIT('h8)
	) name760 (
		_w11271_,
		_w11272_,
		_w11273_
	);
	LUT4 #(
		.INIT('h0001)
	) name761 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[8]/NET0131 ,
		_w11274_
	);
	LUT2 #(
		.INIT('h1)
	) name762 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[5]/NET0131 ,
		_w11275_
	);
	LUT4 #(
		.INIT('h0001)
	) name763 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[15]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131 ,
		_w11276_
	);
	LUT3 #(
		.INIT('h80)
	) name764 (
		_w11274_,
		_w11275_,
		_w11276_,
		_w11277_
	);
	LUT2 #(
		.INIT('h8)
	) name765 (
		_w11273_,
		_w11277_,
		_w11278_
	);
	LUT4 #(
		.INIT('h8000)
	) name766 (
		\ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_Divider2_reg/NET0131 ,
		\maccontrol1_receivecontrol1_Pause_reg/NET0131 ,
		\maccontrol1_receivecontrol1_SlotTimer_reg[0]/NET0131 ,
		_w11279_
	);
	LUT3 #(
		.INIT('h80)
	) name767 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_SlotTimer_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_SlotTimer_reg[3]/NET0131 ,
		_w11280_
	);
	LUT2 #(
		.INIT('h8)
	) name768 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[4]/NET0131 ,
		\maccontrol1_receivecontrol1_SlotTimer_reg[5]/NET0131 ,
		_w11281_
	);
	LUT3 #(
		.INIT('h80)
	) name769 (
		_w11279_,
		_w11280_,
		_w11281_,
		_w11282_
	);
	LUT2 #(
		.INIT('h1)
	) name770 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[1]/NET0131 ,
		_w11283_
	);
	LUT4 #(
		.INIT('h8000)
	) name771 (
		_w11279_,
		_w11280_,
		_w11281_,
		_w11283_,
		_w11284_
	);
	LUT3 #(
		.INIT('h70)
	) name772 (
		_w11273_,
		_w11277_,
		_w11284_,
		_w11285_
	);
	LUT2 #(
		.INIT('h1)
	) name773 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131 ,
		_w11286_
	);
	LUT4 #(
		.INIT('h7000)
	) name774 (
		_w11273_,
		_w11277_,
		_w11284_,
		_w11286_,
		_w11287_
	);
	LUT3 #(
		.INIT('h63)
	) name775 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131 ,
		_w11285_,
		_w11288_
	);
	LUT2 #(
		.INIT('h4)
	) name776 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[3]/NET0131 ,
		_w11268_,
		_w11289_
	);
	LUT4 #(
		.INIT('h7000)
	) name777 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11289_,
		_w11290_
	);
	LUT3 #(
		.INIT('h0b)
	) name778 (
		_w11269_,
		_w11288_,
		_w11290_,
		_w11291_
	);
	LUT4 #(
		.INIT('h4000)
	) name779 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131 ,
		_w11279_,
		_w11280_,
		_w11281_,
		_w11292_
	);
	LUT4 #(
		.INIT('h6a55)
	) name780 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131 ,
		_w11273_,
		_w11277_,
		_w11282_,
		_w11293_
	);
	LUT2 #(
		.INIT('h4)
	) name781 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[0]/NET0131 ,
		_w11268_,
		_w11294_
	);
	LUT4 #(
		.INIT('h7000)
	) name782 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11294_,
		_w11295_
	);
	LUT3 #(
		.INIT('h0b)
	) name783 (
		_w11269_,
		_w11293_,
		_w11295_,
		_w11296_
	);
	LUT4 #(
		.INIT('h0001)
	) name784 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[5]/NET0131 ,
		_w11297_
	);
	LUT4 #(
		.INIT('h7000)
	) name785 (
		_w11273_,
		_w11277_,
		_w11284_,
		_w11297_,
		_w11298_
	);
	LUT3 #(
		.INIT('h01)
	) name786 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[8]/NET0131 ,
		_w11299_
	);
	LUT2 #(
		.INIT('h1)
	) name787 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131 ,
		_w11300_
	);
	LUT4 #(
		.INIT('h6555)
	) name788 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131 ,
		_w11298_,
		_w11299_,
		_w11301_
	);
	LUT2 #(
		.INIT('h4)
	) name789 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[10]/NET0131 ,
		_w11268_,
		_w11302_
	);
	LUT4 #(
		.INIT('h7000)
	) name790 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11302_,
		_w11303_
	);
	LUT3 #(
		.INIT('h0b)
	) name791 (
		_w11269_,
		_w11301_,
		_w11303_,
		_w11304_
	);
	LUT4 #(
		.INIT('h0001)
	) name792 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[11]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[12]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131 ,
		_w11305_
	);
	LUT3 #(
		.INIT('h80)
	) name793 (
		_w11298_,
		_w11299_,
		_w11305_,
		_w11306_
	);
	LUT4 #(
		.INIT('h9555)
	) name794 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131 ,
		_w11298_,
		_w11299_,
		_w11305_,
		_w11307_
	);
	LUT2 #(
		.INIT('h4)
	) name795 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[13]/NET0131 ,
		_w11268_,
		_w11308_
	);
	LUT4 #(
		.INIT('h7000)
	) name796 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11308_,
		_w11309_
	);
	LUT3 #(
		.INIT('h0b)
	) name797 (
		_w11269_,
		_w11307_,
		_w11309_,
		_w11310_
	);
	LUT3 #(
		.INIT('h01)
	) name798 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[11]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131 ,
		_w11311_
	);
	LUT3 #(
		.INIT('h80)
	) name799 (
		_w11298_,
		_w11299_,
		_w11311_,
		_w11312_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name800 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[11]/NET0131 ,
		_w11298_,
		_w11299_,
		_w11300_,
		_w11313_
	);
	LUT2 #(
		.INIT('h1)
	) name801 (
		_w11312_,
		_w11313_,
		_w11314_
	);
	LUT2 #(
		.INIT('h4)
	) name802 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[11]/NET0131 ,
		_w11268_,
		_w11315_
	);
	LUT4 #(
		.INIT('h7000)
	) name803 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11315_,
		_w11316_
	);
	LUT3 #(
		.INIT('h0b)
	) name804 (
		_w11269_,
		_w11314_,
		_w11316_,
		_w11317_
	);
	LUT4 #(
		.INIT('h80aa)
	) name805 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[1]/NET0131 ,
		_w11273_,
		_w11277_,
		_w11292_,
		_w11318_
	);
	LUT2 #(
		.INIT('h1)
	) name806 (
		_w11285_,
		_w11318_,
		_w11319_
	);
	LUT2 #(
		.INIT('h4)
	) name807 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[1]/NET0131 ,
		_w11268_,
		_w11320_
	);
	LUT4 #(
		.INIT('h7000)
	) name808 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11320_,
		_w11321_
	);
	LUT3 #(
		.INIT('h0b)
	) name809 (
		_w11269_,
		_w11319_,
		_w11321_,
		_w11322_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name810 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[15]/NET0131 ,
		_w11273_,
		_w11298_,
		_w11299_,
		_w11323_
	);
	LUT2 #(
		.INIT('h8)
	) name811 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[15]/NET0131 ,
		_w11268_,
		_w11324_
	);
	LUT4 #(
		.INIT('h7000)
	) name812 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11324_,
		_w11325_
	);
	LUT3 #(
		.INIT('hf4)
	) name813 (
		_w11269_,
		_w11323_,
		_w11325_,
		_w11326_
	);
	LUT4 #(
		.INIT('h6a55)
	) name814 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131 ,
		_w11273_,
		_w11277_,
		_w11284_,
		_w11327_
	);
	LUT2 #(
		.INIT('h4)
	) name815 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[2]/NET0131 ,
		_w11268_,
		_w11328_
	);
	LUT4 #(
		.INIT('h7000)
	) name816 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11328_,
		_w11329_
	);
	LUT3 #(
		.INIT('h0b)
	) name817 (
		_w11269_,
		_w11327_,
		_w11329_,
		_w11330_
	);
	LUT3 #(
		.INIT('h63)
	) name818 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131 ,
		_w11298_,
		_w11331_
	);
	LUT2 #(
		.INIT('h4)
	) name819 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[7]/NET0131 ,
		_w11268_,
		_w11332_
	);
	LUT4 #(
		.INIT('h7000)
	) name820 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11332_,
		_w11333_
	);
	LUT3 #(
		.INIT('h0b)
	) name821 (
		_w11269_,
		_w11331_,
		_w11333_,
		_w11334_
	);
	LUT3 #(
		.INIT('h95)
	) name822 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131 ,
		_w11298_,
		_w11299_,
		_w11335_
	);
	LUT2 #(
		.INIT('h4)
	) name823 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[9]/NET0131 ,
		_w11268_,
		_w11336_
	);
	LUT4 #(
		.INIT('h7000)
	) name824 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11336_,
		_w11337_
	);
	LUT3 #(
		.INIT('h0b)
	) name825 (
		_w11269_,
		_w11335_,
		_w11337_,
		_w11338_
	);
	LUT3 #(
		.INIT('h01)
	) name826 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131 ,
		_w11339_
	);
	LUT4 #(
		.INIT('h7000)
	) name827 (
		_w11273_,
		_w11277_,
		_w11284_,
		_w11339_,
		_w11340_
	);
	LUT3 #(
		.INIT('h0d)
	) name828 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131 ,
		_w11287_,
		_w11340_,
		_w11341_
	);
	LUT2 #(
		.INIT('h4)
	) name829 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[4]/NET0131 ,
		_w11268_,
		_w11342_
	);
	LUT4 #(
		.INIT('h7000)
	) name830 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11342_,
		_w11343_
	);
	LUT3 #(
		.INIT('h0b)
	) name831 (
		_w11269_,
		_w11341_,
		_w11343_,
		_w11344_
	);
	LUT3 #(
		.INIT('h31)
	) name832 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[5]/NET0131 ,
		_w11298_,
		_w11340_,
		_w11345_
	);
	LUT2 #(
		.INIT('h4)
	) name833 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[5]/NET0131 ,
		_w11268_,
		_w11346_
	);
	LUT4 #(
		.INIT('h7000)
	) name834 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11346_,
		_w11347_
	);
	LUT3 #(
		.INIT('h0b)
	) name835 (
		_w11269_,
		_w11345_,
		_w11347_,
		_w11348_
	);
	LUT3 #(
		.INIT('h9c)
	) name836 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[14]/NET0131 ,
		_w11306_,
		_w11349_
	);
	LUT2 #(
		.INIT('h4)
	) name837 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[14]/NET0131 ,
		_w11268_,
		_w11350_
	);
	LUT4 #(
		.INIT('h7000)
	) name838 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11350_,
		_w11351_
	);
	LUT3 #(
		.INIT('h0e)
	) name839 (
		_w11269_,
		_w11349_,
		_w11351_,
		_w11352_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name840 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[8]/NET0131 ,
		_w11298_,
		_w11353_
	);
	LUT2 #(
		.INIT('h4)
	) name841 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[8]/NET0131 ,
		_w11268_,
		_w11354_
	);
	LUT4 #(
		.INIT('h7000)
	) name842 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11354_,
		_w11355_
	);
	LUT3 #(
		.INIT('h0b)
	) name843 (
		_w11269_,
		_w11353_,
		_w11355_,
		_w11356_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name844 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[12]/NET0131 ,
		_w11298_,
		_w11299_,
		_w11311_,
		_w11357_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		_w11306_,
		_w11357_,
		_w11358_
	);
	LUT2 #(
		.INIT('h4)
	) name846 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[12]/NET0131 ,
		_w11268_,
		_w11359_
	);
	LUT4 #(
		.INIT('h7000)
	) name847 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11359_,
		_w11360_
	);
	LUT3 #(
		.INIT('h0b)
	) name848 (
		_w11269_,
		_w11358_,
		_w11360_,
		_w11361_
	);
	LUT2 #(
		.INIT('h9)
	) name849 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131 ,
		_w11298_,
		_w11362_
	);
	LUT2 #(
		.INIT('h4)
	) name850 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[6]/NET0131 ,
		_w11268_,
		_w11363_
	);
	LUT4 #(
		.INIT('h7000)
	) name851 (
		_w11141_,
		_w11207_,
		_w11267_,
		_w11363_,
		_w11364_
	);
	LUT3 #(
		.INIT('h0b)
	) name852 (
		_w11269_,
		_w11362_,
		_w11364_,
		_w11365_
	);
	LUT2 #(
		.INIT('h6)
	) name853 (
		_w10590_,
		_w11047_,
		_w11366_
	);
	LUT3 #(
		.INIT('h96)
	) name854 (
		_w10580_,
		_w10590_,
		_w11047_,
		_w11367_
	);
	LUT4 #(
		.INIT('h7000)
	) name855 (
		_w10554_,
		_w10573_,
		_w10577_,
		_w11367_,
		_w11368_
	);
	LUT3 #(
		.INIT('h7b)
	) name856 (
		\rxethmac1_crcrx_Crc_reg[9]/NET0131 ,
		_w10582_,
		_w11368_,
		_w11369_
	);
	LUT3 #(
		.INIT('h02)
	) name857 (
		\txethmac1_txcrc_Crc_reg[14]/NET0131 ,
		_w11030_,
		_w11032_,
		_w11370_
	);
	LUT3 #(
		.INIT('h01)
	) name858 (
		\txethmac1_txcrc_Crc_reg[14]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[30]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11371_
	);
	LUT4 #(
		.INIT('hf800)
	) name859 (
		_w11026_,
		_w11027_,
		_w11028_,
		_w11371_,
		_w11372_
	);
	LUT3 #(
		.INIT('h04)
	) name860 (
		\txethmac1_txcrc_Crc_reg[14]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[30]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11373_
	);
	LUT4 #(
		.INIT('h0700)
	) name861 (
		_w11026_,
		_w11027_,
		_w11028_,
		_w11373_,
		_w11374_
	);
	LUT3 #(
		.INIT('h02)
	) name862 (
		_w11007_,
		_w11372_,
		_w11374_,
		_w11375_
	);
	LUT2 #(
		.INIT('hb)
	) name863 (
		_w11370_,
		_w11375_,
		_w11376_
	);
	LUT3 #(
		.INIT('h02)
	) name864 (
		\txethmac1_txcrc_Crc_reg[15]/NET0131 ,
		_w11052_,
		_w11054_,
		_w11377_
	);
	LUT3 #(
		.INIT('h01)
	) name865 (
		\txethmac1_txcrc_Crc_reg[15]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11378_
	);
	LUT4 #(
		.INIT('hf400)
	) name866 (
		_w11001_,
		_w11002_,
		_w11003_,
		_w11378_,
		_w11379_
	);
	LUT3 #(
		.INIT('h04)
	) name867 (
		\txethmac1_txcrc_Crc_reg[15]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11380_
	);
	LUT4 #(
		.INIT('h0b00)
	) name868 (
		_w11001_,
		_w11002_,
		_w11003_,
		_w11380_,
		_w11381_
	);
	LUT3 #(
		.INIT('h02)
	) name869 (
		_w11007_,
		_w11379_,
		_w11381_,
		_w11382_
	);
	LUT2 #(
		.INIT('hb)
	) name870 (
		_w11377_,
		_w11382_,
		_w11383_
	);
	LUT3 #(
		.INIT('h01)
	) name871 (
		\txethmac1_txcrc_Crc_reg[16]/NET0131 ,
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w11384_
	);
	LUT2 #(
		.INIT('h7)
	) name872 (
		_w10913_,
		_w11384_,
		_w11385_
	);
	LUT3 #(
		.INIT('h70)
	) name873 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		mtxen_pad_o_pad,
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		_w11386_
	);
	LUT2 #(
		.INIT('h4)
	) name874 (
		_w10575_,
		_w11386_,
		_w11387_
	);
	LUT2 #(
		.INIT('h8)
	) name875 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10576_,
		_w11388_
	);
	LUT3 #(
		.INIT('h80)
	) name876 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10548_,
		_w10553_,
		_w11389_
	);
	LUT3 #(
		.INIT('h13)
	) name877 (
		_w10573_,
		_w11388_,
		_w11389_,
		_w11390_
	);
	LUT4 #(
		.INIT('h0103)
	) name878 (
		_w10573_,
		_w11387_,
		_w11388_,
		_w11389_,
		_w11391_
	);
	LUT4 #(
		.INIT('hfefc)
	) name879 (
		_w10573_,
		_w11387_,
		_w11388_,
		_w11389_,
		_w11392_
	);
	LUT3 #(
		.INIT('h45)
	) name880 (
		\macstatus1_ShortFrame_reg/NET0131 ,
		_w10575_,
		_w11386_,
		_w11393_
	);
	LUT4 #(
		.INIT('h1300)
	) name881 (
		_w10573_,
		_w11388_,
		_w11389_,
		_w11393_,
		_w11394_
	);
	LUT2 #(
		.INIT('h1)
	) name882 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		_w11394_,
		_w11395_
	);
	LUT3 #(
		.INIT('hd0)
	) name883 (
		_w11267_,
		_w11391_,
		_w11395_,
		_w11396_
	);
	LUT3 #(
		.INIT('h96)
	) name884 (
		_w10580_,
		_w10590_,
		_w10945_,
		_w11397_
	);
	LUT4 #(
		.INIT('h7000)
	) name885 (
		_w10554_,
		_w10573_,
		_w10577_,
		_w11397_,
		_w11398_
	);
	LUT3 #(
		.INIT('h7b)
	) name886 (
		\rxethmac1_crcrx_Crc_reg[8]/NET0131 ,
		_w10582_,
		_w11398_,
		_w11399_
	);
	LUT2 #(
		.INIT('h4)
	) name887 (
		\rxethmac1_crcrx_Crc_reg[14]/NET0131 ,
		_w10582_,
		_w11400_
	);
	LUT4 #(
		.INIT('h8f00)
	) name888 (
		_w10554_,
		_w10573_,
		_w10591_,
		_w11400_,
		_w11401_
	);
	LUT2 #(
		.INIT('h8)
	) name889 (
		\rxethmac1_crcrx_Crc_reg[14]/NET0131 ,
		_w10582_,
		_w11402_
	);
	LUT4 #(
		.INIT('h7000)
	) name890 (
		_w10554_,
		_w10573_,
		_w10591_,
		_w11402_,
		_w11403_
	);
	LUT2 #(
		.INIT('h1)
	) name891 (
		_w11401_,
		_w11403_,
		_w11404_
	);
	LUT3 #(
		.INIT('h01)
	) name892 (
		\txethmac1_txcrc_Crc_reg[17]/NET0131 ,
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w11405_
	);
	LUT2 #(
		.INIT('h7)
	) name893 (
		_w10913_,
		_w11405_,
		_w11406_
	);
	LUT3 #(
		.INIT('h8a)
	) name894 (
		\macstatus1_ReceivedPacketTooBig_reg/NET0131 ,
		_w10575_,
		_w11386_,
		_w11407_
	);
	LUT4 #(
		.INIT('h1300)
	) name895 (
		_w10573_,
		_w11388_,
		_w11389_,
		_w11407_,
		_w11408_
	);
	LUT3 #(
		.INIT('h04)
	) name896 (
		\ethreg1_MODER_1_DataOut_reg[6]/NET0131 ,
		_w11141_,
		_w11391_,
		_w11409_
	);
	LUT4 #(
		.INIT('h5450)
	) name897 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		_w11207_,
		_w11408_,
		_w11409_,
		_w11410_
	);
	LUT3 #(
		.INIT('h02)
	) name898 (
		\txethmac1_txcrc_Crc_reg[12]/NET0131 ,
		_w11090_,
		_w11092_,
		_w11411_
	);
	LUT3 #(
		.INIT('h01)
	) name899 (
		\txethmac1_txcrc_Crc_reg[12]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[28]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11412_
	);
	LUT4 #(
		.INIT('hf400)
	) name900 (
		_w10996_,
		_w10997_,
		_w10998_,
		_w11412_,
		_w11413_
	);
	LUT3 #(
		.INIT('h04)
	) name901 (
		\txethmac1_txcrc_Crc_reg[12]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[28]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11414_
	);
	LUT4 #(
		.INIT('h0b00)
	) name902 (
		_w10996_,
		_w10997_,
		_w10998_,
		_w11414_,
		_w11415_
	);
	LUT3 #(
		.INIT('h02)
	) name903 (
		_w11007_,
		_w11413_,
		_w11415_,
		_w11416_
	);
	LUT2 #(
		.INIT('hb)
	) name904 (
		_w11411_,
		_w11416_,
		_w11417_
	);
	LUT2 #(
		.INIT('h9)
	) name905 (
		\rxethmac1_crcrx_Crc_reg[29]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[31]/NET0131 ,
		_w11418_
	);
	LUT4 #(
		.INIT('h9669)
	) name906 (
		_w10578_,
		_w10945_,
		_w11045_,
		_w11418_,
		_w11419_
	);
	LUT4 #(
		.INIT('h7000)
	) name907 (
		_w10554_,
		_w10573_,
		_w10577_,
		_w11419_,
		_w11420_
	);
	LUT3 #(
		.INIT('h7b)
	) name908 (
		\rxethmac1_crcrx_Crc_reg[7]/NET0131 ,
		_w10582_,
		_w11420_,
		_w11421_
	);
	LUT3 #(
		.INIT('h02)
	) name909 (
		\txethmac1_txcrc_Crc_reg[13]/NET0131 ,
		_w11016_,
		_w11018_,
		_w11422_
	);
	LUT3 #(
		.INIT('h01)
	) name910 (
		\txethmac1_txcrc_Crc_reg[13]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11423_
	);
	LUT4 #(
		.INIT('hba00)
	) name911 (
		_w11011_,
		_w11012_,
		_w11013_,
		_w11423_,
		_w11424_
	);
	LUT3 #(
		.INIT('h04)
	) name912 (
		\txethmac1_txcrc_Crc_reg[13]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11425_
	);
	LUT4 #(
		.INIT('h4500)
	) name913 (
		_w11011_,
		_w11012_,
		_w11013_,
		_w11425_,
		_w11426_
	);
	LUT3 #(
		.INIT('h02)
	) name914 (
		_w11007_,
		_w11424_,
		_w11426_,
		_w11427_
	);
	LUT2 #(
		.INIT('hb)
	) name915 (
		_w11422_,
		_w11427_,
		_w11428_
	);
	LUT3 #(
		.INIT('h14)
	) name916 (
		\rxethmac1_crcrx_Crc_reg[5]/NET0131 ,
		_w10580_,
		_w10590_,
		_w11429_
	);
	LUT4 #(
		.INIT('h7000)
	) name917 (
		_w10554_,
		_w10573_,
		_w10577_,
		_w11429_,
		_w11430_
	);
	LUT2 #(
		.INIT('h4)
	) name918 (
		\rxethmac1_crcrx_Crc_reg[5]/NET0131 ,
		_w10582_,
		_w11431_
	);
	LUT3 #(
		.INIT('hcd)
	) name919 (
		_w10958_,
		_w11430_,
		_w11431_,
		_w11432_
	);
	LUT4 #(
		.INIT('h0110)
	) name920 (
		\txethmac1_txcrc_Crc_reg[10]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11005_,
		_w11106_,
		_w11433_
	);
	LUT3 #(
		.INIT('h40)
	) name921 (
		\txethmac1_txcrc_Crc_reg[10]/NET0131 ,
		_w10913_,
		_w10914_,
		_w11434_
	);
	LUT3 #(
		.INIT('hab)
	) name922 (
		_w11433_,
		_w11434_,
		_w11126_,
		_w11435_
	);
	LUT3 #(
		.INIT('h02)
	) name923 (
		\txethmac1_txcrc_Crc_reg[11]/NET0131 ,
		_w11052_,
		_w11054_,
		_w11436_
	);
	LUT3 #(
		.INIT('h01)
	) name924 (
		\txethmac1_txcrc_Crc_reg[11]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11437_
	);
	LUT4 #(
		.INIT('hf400)
	) name925 (
		_w11001_,
		_w11002_,
		_w11003_,
		_w11437_,
		_w11438_
	);
	LUT3 #(
		.INIT('h04)
	) name926 (
		\txethmac1_txcrc_Crc_reg[11]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11439_
	);
	LUT4 #(
		.INIT('h0b00)
	) name927 (
		_w11001_,
		_w11002_,
		_w11003_,
		_w11439_,
		_w11440_
	);
	LUT3 #(
		.INIT('h02)
	) name928 (
		_w11007_,
		_w11438_,
		_w11440_,
		_w11441_
	);
	LUT2 #(
		.INIT('hb)
	) name929 (
		_w11436_,
		_w11441_,
		_w11442_
	);
	LUT3 #(
		.INIT('h14)
	) name930 (
		\rxethmac1_crcrx_Crc_reg[10]/NET0131 ,
		_w10590_,
		_w11047_,
		_w11443_
	);
	LUT4 #(
		.INIT('h7000)
	) name931 (
		_w10554_,
		_w10573_,
		_w10577_,
		_w11443_,
		_w11444_
	);
	LUT2 #(
		.INIT('h4)
	) name932 (
		\rxethmac1_crcrx_Crc_reg[10]/NET0131 ,
		_w10582_,
		_w11445_
	);
	LUT2 #(
		.INIT('h8)
	) name933 (
		_w10582_,
		_w11366_,
		_w11446_
	);
	LUT4 #(
		.INIT('h7000)
	) name934 (
		_w10554_,
		_w10573_,
		_w10577_,
		_w11446_,
		_w11447_
	);
	LUT3 #(
		.INIT('hab)
	) name935 (
		_w11444_,
		_w11445_,
		_w11447_,
		_w11448_
	);
	LUT3 #(
		.INIT('h7b)
	) name936 (
		\rxethmac1_crcrx_Crc_reg[4]/NET0131 ,
		_w10582_,
		_w11420_,
		_w11449_
	);
	LUT2 #(
		.INIT('h1)
	) name937 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		_w11450_
	);
	LUT2 #(
		.INIT('h8)
	) name938 (
		\maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w11451_
	);
	LUT3 #(
		.INIT('h40)
	) name939 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w11452_
	);
	LUT2 #(
		.INIT('h8)
	) name940 (
		_w11450_,
		_w11452_,
		_w11453_
	);
	LUT2 #(
		.INIT('h1)
	) name941 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		_w11454_
	);
	LUT3 #(
		.INIT('h01)
	) name942 (
		\rxethmac1_RxData_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11455_
	);
	LUT3 #(
		.INIT('h01)
	) name943 (
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11456_
	);
	LUT2 #(
		.INIT('h2)
	) name944 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11457_
	);
	LUT3 #(
		.INIT('h80)
	) name945 (
		_w11455_,
		_w11456_,
		_w11457_,
		_w11458_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name946 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131 ,
		\ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11459_
	);
	LUT4 #(
		.INIT('h8caf)
	) name947 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131 ,
		\ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11460_
	);
	LUT4 #(
		.INIT('h8421)
	) name948 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131 ,
		\ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11461_
	);
	LUT3 #(
		.INIT('h80)
	) name949 (
		_w11459_,
		_w11460_,
		_w11461_,
		_w11462_
	);
	LUT4 #(
		.INIT('hf531)
	) name950 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131 ,
		\ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11463_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name951 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131 ,
		\ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11464_
	);
	LUT4 #(
		.INIT('hf531)
	) name952 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131 ,
		\ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11465_
	);
	LUT4 #(
		.INIT('h8caf)
	) name953 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131 ,
		\ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11466_
	);
	LUT4 #(
		.INIT('h8000)
	) name954 (
		_w11463_,
		_w11464_,
		_w11465_,
		_w11466_,
		_w11467_
	);
	LUT4 #(
		.INIT('ha888)
	) name955 (
		_w11454_,
		_w11458_,
		_w11462_,
		_w11467_,
		_w11468_
	);
	LUT4 #(
		.INIT('h0100)
	) name956 (
		\rxethmac1_RxData_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11469_
	);
	LUT2 #(
		.INIT('h1)
	) name957 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11470_
	);
	LUT4 #(
		.INIT('h0001)
	) name958 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11471_
	);
	LUT2 #(
		.INIT('h8)
	) name959 (
		_w11469_,
		_w11471_,
		_w11472_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name960 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131 ,
		\ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11473_
	);
	LUT4 #(
		.INIT('h8caf)
	) name961 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11474_
	);
	LUT4 #(
		.INIT('h8421)
	) name962 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w11475_
	);
	LUT3 #(
		.INIT('h80)
	) name963 (
		_w11473_,
		_w11474_,
		_w11475_,
		_w11476_
	);
	LUT4 #(
		.INIT('hf531)
	) name964 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11477_
	);
	LUT4 #(
		.INIT('haf23)
	) name965 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11478_
	);
	LUT4 #(
		.INIT('hf531)
	) name966 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11479_
	);
	LUT4 #(
		.INIT('h8caf)
	) name967 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11480_
	);
	LUT4 #(
		.INIT('h8000)
	) name968 (
		_w11477_,
		_w11478_,
		_w11479_,
		_w11480_,
		_w11481_
	);
	LUT2 #(
		.INIT('h2)
	) name969 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		_w11482_
	);
	LUT3 #(
		.INIT('h08)
	) name970 (
		\maccontrol1_receivecontrol1_AddressOK_reg/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		_w11483_
	);
	LUT4 #(
		.INIT('hea00)
	) name971 (
		_w11472_,
		_w11476_,
		_w11481_,
		_w11483_,
		_w11484_
	);
	LUT3 #(
		.INIT('ha8)
	) name972 (
		_w11453_,
		_w11468_,
		_w11484_,
		_w11485_
	);
	LUT4 #(
		.INIT('h2000)
	) name973 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w11486_
	);
	LUT2 #(
		.INIT('h1)
	) name974 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		_w11487_
	);
	LUT3 #(
		.INIT('h15)
	) name975 (
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w11486_,
		_w11487_,
		_w11488_
	);
	LUT2 #(
		.INIT('h4)
	) name976 (
		_w11453_,
		_w11488_,
		_w11489_
	);
	LUT4 #(
		.INIT('haf23)
	) name977 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w11490_
	);
	LUT4 #(
		.INIT('h8caf)
	) name978 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11491_
	);
	LUT4 #(
		.INIT('h8421)
	) name979 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131 ,
		\ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11492_
	);
	LUT3 #(
		.INIT('h80)
	) name980 (
		_w11490_,
		_w11491_,
		_w11492_,
		_w11493_
	);
	LUT4 #(
		.INIT('hf531)
	) name981 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11494_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name982 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w11495_
	);
	LUT4 #(
		.INIT('hf531)
	) name983 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11496_
	);
	LUT4 #(
		.INIT('h8caf)
	) name984 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11497_
	);
	LUT4 #(
		.INIT('h8000)
	) name985 (
		_w11494_,
		_w11495_,
		_w11496_,
		_w11497_,
		_w11498_
	);
	LUT4 #(
		.INIT('hc888)
	) name986 (
		_w11458_,
		_w11482_,
		_w11493_,
		_w11498_,
		_w11499_
	);
	LUT3 #(
		.INIT('h80)
	) name987 (
		_w11455_,
		_w11456_,
		_w11470_,
		_w11500_
	);
	LUT4 #(
		.INIT('haf23)
	) name988 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131 ,
		\ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11501_
	);
	LUT4 #(
		.INIT('h8caf)
	) name989 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131 ,
		\ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11502_
	);
	LUT4 #(
		.INIT('h8421)
	) name990 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131 ,
		\ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11503_
	);
	LUT3 #(
		.INIT('h80)
	) name991 (
		_w11501_,
		_w11502_,
		_w11503_,
		_w11504_
	);
	LUT4 #(
		.INIT('hf531)
	) name992 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131 ,
		\ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11505_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name993 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131 ,
		\ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11506_
	);
	LUT4 #(
		.INIT('hf531)
	) name994 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131 ,
		\ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11507_
	);
	LUT4 #(
		.INIT('h8caf)
	) name995 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131 ,
		\ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11508_
	);
	LUT4 #(
		.INIT('h8000)
	) name996 (
		_w11505_,
		_w11506_,
		_w11507_,
		_w11508_,
		_w11509_
	);
	LUT4 #(
		.INIT('ha888)
	) name997 (
		_w11454_,
		_w11500_,
		_w11504_,
		_w11509_,
		_w11510_
	);
	LUT4 #(
		.INIT('h0200)
	) name998 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131 ,
		_w11451_,
		_w11511_
	);
	LUT4 #(
		.INIT('h0155)
	) name999 (
		_w11489_,
		_w11499_,
		_w11510_,
		_w11511_,
		_w11512_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name1000 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131 ,
		\ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11513_
	);
	LUT4 #(
		.INIT('h8caf)
	) name1001 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131 ,
		\ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11514_
	);
	LUT4 #(
		.INIT('h8421)
	) name1002 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131 ,
		\ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11515_
	);
	LUT3 #(
		.INIT('h80)
	) name1003 (
		_w11513_,
		_w11514_,
		_w11515_,
		_w11516_
	);
	LUT4 #(
		.INIT('hf531)
	) name1004 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131 ,
		\ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11517_
	);
	LUT4 #(
		.INIT('haf23)
	) name1005 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131 ,
		\ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11518_
	);
	LUT4 #(
		.INIT('hf531)
	) name1006 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131 ,
		\ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11519_
	);
	LUT4 #(
		.INIT('h8caf)
	) name1007 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131 ,
		\ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11520_
	);
	LUT4 #(
		.INIT('h8000)
	) name1008 (
		_w11517_,
		_w11518_,
		_w11519_,
		_w11520_,
		_w11521_
	);
	LUT2 #(
		.INIT('h8)
	) name1009 (
		_w11516_,
		_w11521_,
		_w11522_
	);
	LUT4 #(
		.INIT('h2000)
	) name1010 (
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11523_
	);
	LUT4 #(
		.INIT('h0001)
	) name1011 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11524_
	);
	LUT3 #(
		.INIT('h15)
	) name1012 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		_w11523_,
		_w11524_,
		_w11525_
	);
	LUT3 #(
		.INIT('h70)
	) name1013 (
		_w11516_,
		_w11521_,
		_w11525_,
		_w11526_
	);
	LUT4 #(
		.INIT('haf23)
	) name1014 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131 ,
		\ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11527_
	);
	LUT4 #(
		.INIT('h8caf)
	) name1015 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131 ,
		\ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11528_
	);
	LUT4 #(
		.INIT('h8421)
	) name1016 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131 ,
		\ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11529_
	);
	LUT3 #(
		.INIT('h80)
	) name1017 (
		_w11527_,
		_w11528_,
		_w11529_,
		_w11530_
	);
	LUT4 #(
		.INIT('hf531)
	) name1018 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131 ,
		\ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11531_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name1019 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131 ,
		\ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11532_
	);
	LUT4 #(
		.INIT('hf531)
	) name1020 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131 ,
		\ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11533_
	);
	LUT4 #(
		.INIT('h8caf)
	) name1021 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131 ,
		\ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11534_
	);
	LUT4 #(
		.INIT('h8000)
	) name1022 (
		_w11531_,
		_w11532_,
		_w11533_,
		_w11534_,
		_w11535_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1023 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		_w11455_,
		_w11456_,
		_w11470_,
		_w11536_
	);
	LUT3 #(
		.INIT('h02)
	) name1024 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		_w11537_
	);
	LUT2 #(
		.INIT('h8)
	) name1025 (
		_w11452_,
		_w11537_,
		_w11538_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1026 (
		_w11530_,
		_w11535_,
		_w11536_,
		_w11538_,
		_w11539_
	);
	LUT2 #(
		.INIT('h4)
	) name1027 (
		_w11526_,
		_w11539_,
		_w11540_
	);
	LUT4 #(
		.INIT('heece)
	) name1028 (
		\maccontrol1_receivecontrol1_AddressOK_reg/NET0131 ,
		_w11485_,
		_w11512_,
		_w11540_,
		_w11541_
	);
	LUT2 #(
		.INIT('h4)
	) name1029 (
		\rxethmac1_crcrx_Crc_reg[25]/NET0131 ,
		_w10582_,
		_w11542_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1030 (
		_w10554_,
		_w10573_,
		_w11081_,
		_w11542_,
		_w11543_
	);
	LUT2 #(
		.INIT('h8)
	) name1031 (
		\rxethmac1_crcrx_Crc_reg[25]/NET0131 ,
		_w10582_,
		_w11544_
	);
	LUT4 #(
		.INIT('h7000)
	) name1032 (
		_w10554_,
		_w10573_,
		_w11081_,
		_w11544_,
		_w11545_
	);
	LUT2 #(
		.INIT('h1)
	) name1033 (
		_w11543_,
		_w11545_,
		_w11546_
	);
	LUT3 #(
		.INIT('h20)
	) name1034 (
		\WillTransmit_q2_reg/P0001 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		_w11547_
	);
	LUT3 #(
		.INIT('h04)
	) name1035 (
		_w10578_,
		_w10588_,
		_w11045_,
		_w11548_
	);
	LUT4 #(
		.INIT('he400)
	) name1036 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[3]_pad ,
		\mtxd_pad_o[3]_pad ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w11549_
	);
	LUT4 #(
		.INIT('h0400)
	) name1037 (
		_w10578_,
		_w10588_,
		_w11045_,
		_w11549_,
		_w11550_
	);
	LUT2 #(
		.INIT('h1)
	) name1038 (
		\rxethmac1_rxcounters1_IFGCounter_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131 ,
		_w11551_
	);
	LUT3 #(
		.INIT('h40)
	) name1039 (
		\rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_IFGCounter_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_IFGCounter_reg[4]/NET0131 ,
		_w11552_
	);
	LUT3 #(
		.INIT('h15)
	) name1040 (
		\ethreg1_MODER_0_DataOut_reg[6]/NET0131 ,
		_w11551_,
		_w11552_,
		_w11553_
	);
	LUT3 #(
		.INIT('h15)
	) name1041 (
		_w11547_,
		_w11550_,
		_w11553_,
		_w11554_
	);
	LUT4 #(
		.INIT('h2033)
	) name1042 (
		_w10573_,
		_w10576_,
		_w11389_,
		_w11554_,
		_w11555_
	);
	LUT2 #(
		.INIT('h2)
	) name1043 (
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		_w10576_,
		_w11556_
	);
	LUT4 #(
		.INIT('h3222)
	) name1044 (
		\ethreg1_MODER_0_DataOut_reg[6]/NET0131 ,
		_w10576_,
		_w11551_,
		_w11552_,
		_w11557_
	);
	LUT3 #(
		.INIT('h01)
	) name1045 (
		\rxethmac1_rxstatem1_StateDrop_reg/NET0131 ,
		\rxethmac1_rxstatem1_StatePreamble_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w11558_
	);
	LUT3 #(
		.INIT('h4c)
	) name1046 (
		_w10574_,
		_w10576_,
		_w11558_,
		_w11559_
	);
	LUT4 #(
		.INIT('h0013)
	) name1047 (
		_w11550_,
		_w11556_,
		_w11557_,
		_w11559_,
		_w11560_
	);
	LUT4 #(
		.INIT('h0040)
	) name1048 (
		_w10578_,
		_w10588_,
		_w10943_,
		_w11045_,
		_w11561_
	);
	LUT3 #(
		.INIT('hd0)
	) name1049 (
		\WillTransmit_q2_reg/P0001 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		_w11562_
	);
	LUT2 #(
		.INIT('h4)
	) name1050 (
		_w10576_,
		_w11562_,
		_w11563_
	);
	LUT4 #(
		.INIT('h002f)
	) name1051 (
		\WillTransmit_q2_reg/P0001 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		\rxethmac1_rxstatem1_StatePreamble_reg/NET0131 ,
		_w11564_
	);
	LUT2 #(
		.INIT('h1)
	) name1052 (
		_w10576_,
		_w11564_,
		_w11565_
	);
	LUT4 #(
		.INIT('hce8a)
	) name1053 (
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w11561_,
		_w11563_,
		_w11565_,
		_w11566_
	);
	LUT2 #(
		.INIT('h8)
	) name1054 (
		_w11560_,
		_w11566_,
		_w11567_
	);
	LUT2 #(
		.INIT('h4)
	) name1055 (
		_w11555_,
		_w11567_,
		_w11568_
	);
	LUT4 #(
		.INIT('hebbe)
	) name1056 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11000_,
		_w11105_,
		_w11106_,
		_w11569_
	);
	LUT2 #(
		.INIT('h1)
	) name1057 (
		\txethmac1_txcrc_Crc_reg[8]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11570_
	);
	LUT4 #(
		.INIT('h96ff)
	) name1058 (
		_w11000_,
		_w11105_,
		_w11106_,
		_w11570_,
		_w11571_
	);
	LUT4 #(
		.INIT('hb3ff)
	) name1059 (
		\txethmac1_txcrc_Crc_reg[8]/NET0131 ,
		_w11007_,
		_w11569_,
		_w11571_,
		_w11572_
	);
	LUT3 #(
		.INIT('h96)
	) name1060 (
		_w10590_,
		_w10945_,
		_w11047_,
		_w11573_
	);
	LUT4 #(
		.INIT('h7000)
	) name1061 (
		_w10554_,
		_w10573_,
		_w10577_,
		_w11573_,
		_w11574_
	);
	LUT3 #(
		.INIT('h7b)
	) name1062 (
		\rxethmac1_crcrx_Crc_reg[3]/NET0131 ,
		_w10582_,
		_w11574_,
		_w11575_
	);
	LUT2 #(
		.INIT('h1)
	) name1063 (
		\rxethmac1_rxstatem1_StatePreamble_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w11576_
	);
	LUT2 #(
		.INIT('h4)
	) name1064 (
		_w11562_,
		_w11576_,
		_w11577_
	);
	LUT3 #(
		.INIT('hc4)
	) name1065 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		_w10543_,
		_w11578_
	);
	LUT3 #(
		.INIT('h80)
	) name1066 (
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		_w11579_
	);
	LUT2 #(
		.INIT('h8)
	) name1067 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w11580_
	);
	LUT3 #(
		.INIT('h80)
	) name1068 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w11581_
	);
	LUT3 #(
		.INIT('h80)
	) name1069 (
		_w11579_,
		_w11136_,
		_w11581_,
		_w11582_
	);
	LUT4 #(
		.INIT('h8000)
	) name1070 (
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w11583_
	);
	LUT2 #(
		.INIT('h8)
	) name1071 (
		_w11139_,
		_w11583_,
		_w11584_
	);
	LUT4 #(
		.INIT('h5ddd)
	) name1072 (
		_w11577_,
		_w11578_,
		_w11582_,
		_w11584_,
		_w11585_
	);
	LUT2 #(
		.INIT('h1)
	) name1073 (
		_w10576_,
		_w11550_,
		_w11586_
	);
	LUT4 #(
		.INIT('h7000)
	) name1074 (
		_w10573_,
		_w11389_,
		_w11585_,
		_w11586_,
		_w11587_
	);
	LUT4 #(
		.INIT('h3320)
	) name1075 (
		_w10573_,
		_w10576_,
		_w11389_,
		_w11550_,
		_w11588_
	);
	LUT3 #(
		.INIT('h06)
	) name1076 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		_w11587_,
		_w11588_,
		_w11589_
	);
	LUT3 #(
		.INIT('h80)
	) name1077 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w11590_
	);
	LUT3 #(
		.INIT('h80)
	) name1078 (
		_w11579_,
		_w11136_,
		_w11590_,
		_w11591_
	);
	LUT4 #(
		.INIT('h1555)
	) name1079 (
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w11587_,
		_w11591_,
		_w11592_
	);
	LUT4 #(
		.INIT('h8000)
	) name1080 (
		_w11579_,
		_w11136_,
		_w11580_,
		_w11137_,
		_w11593_
	);
	LUT3 #(
		.INIT('h13)
	) name1081 (
		_w11587_,
		_w11588_,
		_w11593_,
		_w11594_
	);
	LUT2 #(
		.INIT('h4)
	) name1082 (
		_w11592_,
		_w11594_,
		_w11595_
	);
	LUT4 #(
		.INIT('h060a)
	) name1083 (
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w11587_,
		_w11588_,
		_w11593_,
		_w11596_
	);
	LUT4 #(
		.INIT('h1555)
	) name1084 (
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		_w11146_,
		_w11587_,
		_w11593_,
		_w11597_
	);
	LUT4 #(
		.INIT('h070f)
	) name1085 (
		_w11139_,
		_w11587_,
		_w11588_,
		_w11593_,
		_w11598_
	);
	LUT2 #(
		.INIT('h4)
	) name1086 (
		_w11597_,
		_w11598_,
		_w11599_
	);
	LUT4 #(
		.INIT('h1333)
	) name1087 (
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		_w11587_,
		_w11593_,
		_w11600_
	);
	LUT4 #(
		.INIT('h070f)
	) name1088 (
		_w11146_,
		_w11587_,
		_w11588_,
		_w11593_,
		_w11601_
	);
	LUT2 #(
		.INIT('h4)
	) name1089 (
		_w11600_,
		_w11601_,
		_w11602_
	);
	LUT4 #(
		.INIT('h1555)
	) name1090 (
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		_w11139_,
		_w11587_,
		_w11593_,
		_w11603_
	);
	LUT3 #(
		.INIT('h80)
	) name1091 (
		_w11579_,
		_w11136_,
		_w11580_,
		_w11604_
	);
	LUT2 #(
		.INIT('h8)
	) name1092 (
		_w11584_,
		_w11604_,
		_w11605_
	);
	LUT3 #(
		.INIT('h13)
	) name1093 (
		_w11587_,
		_w11588_,
		_w11605_,
		_w11606_
	);
	LUT2 #(
		.INIT('h4)
	) name1094 (
		_w11603_,
		_w11606_,
		_w11607_
	);
	LUT4 #(
		.INIT('h060a)
	) name1095 (
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		_w11587_,
		_w11588_,
		_w11605_,
		_w11608_
	);
	LUT4 #(
		.INIT('h006c)
	) name1096 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w11587_,
		_w11588_,
		_w11609_
	);
	LUT3 #(
		.INIT('h80)
	) name1097 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		_w11610_
	);
	LUT4 #(
		.INIT('h006a)
	) name1098 (
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		_w11580_,
		_w11587_,
		_w11588_,
		_w11611_
	);
	LUT4 #(
		.INIT('h8000)
	) name1099 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w11612_
	);
	LUT4 #(
		.INIT('h060a)
	) name1100 (
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w11587_,
		_w11588_,
		_w11610_,
		_w11613_
	);
	LUT3 #(
		.INIT('h15)
	) name1101 (
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		_w11587_,
		_w11612_,
		_w11614_
	);
	LUT2 #(
		.INIT('h8)
	) name1102 (
		_w11579_,
		_w11580_,
		_w11615_
	);
	LUT3 #(
		.INIT('h13)
	) name1103 (
		_w11587_,
		_w11588_,
		_w11615_,
		_w11616_
	);
	LUT2 #(
		.INIT('h4)
	) name1104 (
		_w11614_,
		_w11616_,
		_w11617_
	);
	LUT3 #(
		.INIT('h15)
	) name1105 (
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w11587_,
		_w11615_,
		_w11618_
	);
	LUT3 #(
		.INIT('h80)
	) name1106 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w11619_
	);
	LUT2 #(
		.INIT('h8)
	) name1107 (
		_w11579_,
		_w11619_,
		_w11620_
	);
	LUT3 #(
		.INIT('h13)
	) name1108 (
		_w11587_,
		_w11588_,
		_w11620_,
		_w11621_
	);
	LUT2 #(
		.INIT('h4)
	) name1109 (
		_w11618_,
		_w11621_,
		_w11622_
	);
	LUT4 #(
		.INIT('h060a)
	) name1110 (
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		_w11587_,
		_w11588_,
		_w11620_,
		_w11623_
	);
	LUT4 #(
		.INIT('h1333)
	) name1111 (
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		_w11587_,
		_w11620_,
		_w11624_
	);
	LUT3 #(
		.INIT('h13)
	) name1112 (
		_w11587_,
		_w11588_,
		_w11604_,
		_w11625_
	);
	LUT2 #(
		.INIT('h4)
	) name1113 (
		_w11624_,
		_w11625_,
		_w11626_
	);
	LUT3 #(
		.INIT('h15)
	) name1114 (
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w11587_,
		_w11604_,
		_w11627_
	);
	LUT3 #(
		.INIT('h13)
	) name1115 (
		_w11587_,
		_w11588_,
		_w11591_,
		_w11628_
	);
	LUT2 #(
		.INIT('h4)
	) name1116 (
		_w11627_,
		_w11628_,
		_w11629_
	);
	LUT4 #(
		.INIT('h060a)
	) name1117 (
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w11587_,
		_w11588_,
		_w11591_,
		_w11630_
	);
	LUT4 #(
		.INIT('hbeeb)
	) name1118 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11005_,
		_w11105_,
		_w11106_,
		_w11631_
	);
	LUT2 #(
		.INIT('h1)
	) name1119 (
		\txethmac1_txcrc_Crc_reg[9]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11632_
	);
	LUT4 #(
		.INIT('h69ff)
	) name1120 (
		_w11005_,
		_w11105_,
		_w11106_,
		_w11632_,
		_w11633_
	);
	LUT4 #(
		.INIT('hb3ff)
	) name1121 (
		\txethmac1_txcrc_Crc_reg[9]/NET0131 ,
		_w11007_,
		_w11631_,
		_w11633_,
		_w11634_
	);
	LUT2 #(
		.INIT('h2)
	) name1122 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10576_,
		_w11635_
	);
	LUT4 #(
		.INIT('h4055)
	) name1123 (
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		_w10554_,
		_w10573_,
		_w11635_,
		_w11636_
	);
	LUT3 #(
		.INIT('h04)
	) name1124 (
		_w11555_,
		_w11560_,
		_w11636_,
		_w11637_
	);
	LUT2 #(
		.INIT('h4)
	) name1125 (
		_w10576_,
		_w11549_,
		_w11638_
	);
	LUT4 #(
		.INIT('h0001)
	) name1126 (
		\rxethmac1_rxstatem1_StateDrop_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		\rxethmac1_rxstatem1_StatePreamble_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w11639_
	);
	LUT4 #(
		.INIT('h0015)
	) name1127 (
		\ethreg1_MODER_0_DataOut_reg[6]/NET0131 ,
		_w11551_,
		_w11552_,
		_w11639_,
		_w11640_
	);
	LUT2 #(
		.INIT('h2)
	) name1128 (
		\rxethmac1_rxcounters1_IFGCounter_reg[0]/NET0131 ,
		\rxethmac1_rxstatem1_StateDrop_reg/NET0131 ,
		_w11641_
	);
	LUT4 #(
		.INIT('h7000)
	) name1129 (
		_w11548_,
		_w11638_,
		_w11640_,
		_w11641_,
		_w11642_
	);
	LUT3 #(
		.INIT('h80)
	) name1130 (
		\rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_IFGCounter_reg[3]/NET0131 ,
		_w11643_
	);
	LUT3 #(
		.INIT('h15)
	) name1131 (
		\rxethmac1_rxstatem1_StateDrop_reg/NET0131 ,
		_w11548_,
		_w11638_,
		_w11644_
	);
	LUT4 #(
		.INIT('h6a00)
	) name1132 (
		\rxethmac1_rxcounters1_IFGCounter_reg[4]/NET0131 ,
		_w11642_,
		_w11643_,
		_w11644_,
		_w11645_
	);
	LUT2 #(
		.INIT('h8)
	) name1133 (
		\rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131 ,
		_w11646_
	);
	LUT4 #(
		.INIT('h6c00)
	) name1134 (
		\rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131 ,
		_w11642_,
		_w11644_,
		_w11647_
	);
	LUT3 #(
		.INIT('h15)
	) name1135 (
		\rxethmac1_rxcounters1_IFGCounter_reg[3]/NET0131 ,
		_w11642_,
		_w11646_,
		_w11648_
	);
	LUT3 #(
		.INIT('h70)
	) name1136 (
		_w11642_,
		_w11643_,
		_w11644_,
		_w11649_
	);
	LUT2 #(
		.INIT('h4)
	) name1137 (
		_w11648_,
		_w11649_,
		_w11650_
	);
	LUT4 #(
		.INIT('h0700)
	) name1138 (
		_w11548_,
		_w11638_,
		_w11640_,
		_w11641_,
		_w11651_
	);
	LUT2 #(
		.INIT('h1)
	) name1139 (
		\rxethmac1_rxcounters1_IFGCounter_reg[0]/NET0131 ,
		\rxethmac1_rxstatem1_StateDrop_reg/NET0131 ,
		_w11652_
	);
	LUT4 #(
		.INIT('h7000)
	) name1140 (
		_w11548_,
		_w11638_,
		_w11640_,
		_w11652_,
		_w11653_
	);
	LUT2 #(
		.INIT('he)
	) name1141 (
		_w11651_,
		_w11653_,
		_w11654_
	);
	LUT2 #(
		.INIT('h8)
	) name1142 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		_w11655_
	);
	LUT2 #(
		.INIT('h4)
	) name1143 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w11656_
	);
	LUT3 #(
		.INIT('h40)
	) name1144 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w11657_
	);
	LUT3 #(
		.INIT('h40)
	) name1145 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_Flop_reg/NET0131 ,
		_w11658_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1146 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_Flop_reg/NET0131 ,
		\wishbone_TxData_reg[1]/NET0131 ,
		_w11659_
	);
	LUT3 #(
		.INIT('h70)
	) name1147 (
		_w11655_,
		_w11657_,
		_w11659_,
		_w11660_
	);
	LUT4 #(
		.INIT('h57df)
	) name1148 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[17]/NET0131 ,
		\wishbone_TxDataLatched_reg[1]/NET0131 ,
		_w11661_
	);
	LUT4 #(
		.INIT('habef)
	) name1149 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[25]/NET0131 ,
		\wishbone_TxDataLatched_reg[9]/NET0131 ,
		_w11662_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		_w11661_,
		_w11662_,
		_w11663_
	);
	LUT3 #(
		.INIT('h70)
	) name1151 (
		_w11655_,
		_w11657_,
		_w11658_,
		_w11664_
	);
	LUT3 #(
		.INIT('h80)
	) name1152 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[25]/P0001 ,
		_w11665_
	);
	LUT2 #(
		.INIT('h4)
	) name1153 (
		\wishbone_TxStartFrm_reg/NET0131 ,
		\wishbone_TxStartFrm_sync2_reg/NET0131 ,
		_w11666_
	);
	LUT3 #(
		.INIT('h07)
	) name1154 (
		_w11657_,
		_w11665_,
		_w11666_,
		_w11667_
	);
	LUT4 #(
		.INIT('h4500)
	) name1155 (
		_w11660_,
		_w11663_,
		_w11664_,
		_w11667_,
		_w11668_
	);
	LUT3 #(
		.INIT('h10)
	) name1156 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[25]/P0001 ,
		_w11669_
	);
	LUT3 #(
		.INIT('h40)
	) name1157 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[9]/P0001 ,
		_w11670_
	);
	LUT4 #(
		.INIT('h57df)
	) name1158 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[17]/P0001 ,
		\wishbone_tx_fifo_data_out_reg[1]/P0001 ,
		_w11671_
	);
	LUT4 #(
		.INIT('h0200)
	) name1159 (
		_w11666_,
		_w11669_,
		_w11670_,
		_w11671_,
		_w11672_
	);
	LUT2 #(
		.INIT('h1)
	) name1160 (
		_w11668_,
		_w11672_,
		_w11673_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1161 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_Flop_reg/NET0131 ,
		\wishbone_TxData_reg[2]/NET0131 ,
		_w11674_
	);
	LUT3 #(
		.INIT('h70)
	) name1162 (
		_w11655_,
		_w11657_,
		_w11674_,
		_w11675_
	);
	LUT4 #(
		.INIT('haebf)
	) name1163 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[10]/NET0131 ,
		\wishbone_TxDataLatched_reg[26]/NET0131 ,
		_w11676_
	);
	LUT4 #(
		.INIT('h57df)
	) name1164 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[18]/NET0131 ,
		\wishbone_TxDataLatched_reg[2]/NET0131 ,
		_w11677_
	);
	LUT2 #(
		.INIT('h8)
	) name1165 (
		_w11676_,
		_w11677_,
		_w11678_
	);
	LUT3 #(
		.INIT('h80)
	) name1166 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[26]/P0001 ,
		_w11679_
	);
	LUT3 #(
		.INIT('h13)
	) name1167 (
		_w11657_,
		_w11666_,
		_w11679_,
		_w11680_
	);
	LUT4 #(
		.INIT('h3100)
	) name1168 (
		_w11664_,
		_w11675_,
		_w11678_,
		_w11680_,
		_w11681_
	);
	LUT3 #(
		.INIT('h10)
	) name1169 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[26]/P0001 ,
		_w11682_
	);
	LUT3 #(
		.INIT('h40)
	) name1170 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[10]/P0001 ,
		_w11683_
	);
	LUT4 #(
		.INIT('h57df)
	) name1171 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[18]/P0001 ,
		\wishbone_tx_fifo_data_out_reg[2]/P0001 ,
		_w11684_
	);
	LUT4 #(
		.INIT('h0200)
	) name1172 (
		_w11666_,
		_w11682_,
		_w11683_,
		_w11684_,
		_w11685_
	);
	LUT2 #(
		.INIT('h1)
	) name1173 (
		_w11681_,
		_w11685_,
		_w11686_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1174 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_Flop_reg/NET0131 ,
		\wishbone_TxData_reg[3]/NET0131 ,
		_w11687_
	);
	LUT3 #(
		.INIT('h70)
	) name1175 (
		_w11655_,
		_w11657_,
		_w11687_,
		_w11688_
	);
	LUT4 #(
		.INIT('h57df)
	) name1176 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[19]/NET0131 ,
		\wishbone_TxDataLatched_reg[3]/NET0131 ,
		_w11689_
	);
	LUT4 #(
		.INIT('haebf)
	) name1177 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[11]/NET0131 ,
		\wishbone_TxDataLatched_reg[27]/NET0131 ,
		_w11690_
	);
	LUT2 #(
		.INIT('h8)
	) name1178 (
		_w11689_,
		_w11690_,
		_w11691_
	);
	LUT3 #(
		.INIT('h80)
	) name1179 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[27]/P0001 ,
		_w11692_
	);
	LUT3 #(
		.INIT('h13)
	) name1180 (
		_w11657_,
		_w11666_,
		_w11692_,
		_w11693_
	);
	LUT4 #(
		.INIT('h3100)
	) name1181 (
		_w11664_,
		_w11688_,
		_w11691_,
		_w11693_,
		_w11694_
	);
	LUT3 #(
		.INIT('h10)
	) name1182 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[27]/P0001 ,
		_w11695_
	);
	LUT3 #(
		.INIT('h40)
	) name1183 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[11]/P0001 ,
		_w11696_
	);
	LUT4 #(
		.INIT('h57df)
	) name1184 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[19]/P0001 ,
		\wishbone_tx_fifo_data_out_reg[3]/P0001 ,
		_w11697_
	);
	LUT4 #(
		.INIT('h0200)
	) name1185 (
		_w11666_,
		_w11695_,
		_w11696_,
		_w11697_,
		_w11698_
	);
	LUT2 #(
		.INIT('h1)
	) name1186 (
		_w11694_,
		_w11698_,
		_w11699_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1187 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_Flop_reg/NET0131 ,
		\wishbone_TxData_reg[4]/NET0131 ,
		_w11700_
	);
	LUT3 #(
		.INIT('h70)
	) name1188 (
		_w11655_,
		_w11657_,
		_w11700_,
		_w11701_
	);
	LUT4 #(
		.INIT('h57df)
	) name1189 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[20]/NET0131 ,
		\wishbone_TxDataLatched_reg[4]/NET0131 ,
		_w11702_
	);
	LUT4 #(
		.INIT('haebf)
	) name1190 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[12]/NET0131 ,
		\wishbone_TxDataLatched_reg[28]/NET0131 ,
		_w11703_
	);
	LUT2 #(
		.INIT('h8)
	) name1191 (
		_w11702_,
		_w11703_,
		_w11704_
	);
	LUT3 #(
		.INIT('h80)
	) name1192 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[28]/P0001 ,
		_w11705_
	);
	LUT3 #(
		.INIT('h13)
	) name1193 (
		_w11657_,
		_w11666_,
		_w11705_,
		_w11706_
	);
	LUT4 #(
		.INIT('h3100)
	) name1194 (
		_w11664_,
		_w11701_,
		_w11704_,
		_w11706_,
		_w11707_
	);
	LUT3 #(
		.INIT('h10)
	) name1195 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[28]/P0001 ,
		_w11708_
	);
	LUT3 #(
		.INIT('h40)
	) name1196 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[12]/P0001 ,
		_w11709_
	);
	LUT4 #(
		.INIT('h57df)
	) name1197 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[20]/P0001 ,
		\wishbone_tx_fifo_data_out_reg[4]/P0001 ,
		_w11710_
	);
	LUT4 #(
		.INIT('h0200)
	) name1198 (
		_w11666_,
		_w11708_,
		_w11709_,
		_w11710_,
		_w11711_
	);
	LUT2 #(
		.INIT('h1)
	) name1199 (
		_w11707_,
		_w11711_,
		_w11712_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1200 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_Flop_reg/NET0131 ,
		\wishbone_TxData_reg[0]/NET0131 ,
		_w11713_
	);
	LUT3 #(
		.INIT('h70)
	) name1201 (
		_w11655_,
		_w11657_,
		_w11713_,
		_w11714_
	);
	LUT4 #(
		.INIT('habef)
	) name1202 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[24]/NET0131 ,
		\wishbone_TxDataLatched_reg[8]/NET0131 ,
		_w11715_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name1203 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[0]/NET0131 ,
		\wishbone_TxDataLatched_reg[16]/NET0131 ,
		_w11716_
	);
	LUT2 #(
		.INIT('h8)
	) name1204 (
		_w11715_,
		_w11716_,
		_w11717_
	);
	LUT3 #(
		.INIT('h80)
	) name1205 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[24]/P0001 ,
		_w11718_
	);
	LUT3 #(
		.INIT('h13)
	) name1206 (
		_w11657_,
		_w11666_,
		_w11718_,
		_w11719_
	);
	LUT4 #(
		.INIT('h3100)
	) name1207 (
		_w11664_,
		_w11714_,
		_w11717_,
		_w11719_,
		_w11720_
	);
	LUT3 #(
		.INIT('h10)
	) name1208 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[24]/P0001 ,
		_w11721_
	);
	LUT3 #(
		.INIT('h40)
	) name1209 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[8]/P0001 ,
		_w11722_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name1210 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[0]/P0001 ,
		\wishbone_tx_fifo_data_out_reg[16]/P0001 ,
		_w11723_
	);
	LUT4 #(
		.INIT('h0200)
	) name1211 (
		_w11666_,
		_w11721_,
		_w11722_,
		_w11723_,
		_w11724_
	);
	LUT2 #(
		.INIT('h1)
	) name1212 (
		_w11720_,
		_w11724_,
		_w11725_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1213 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_Flop_reg/NET0131 ,
		\wishbone_TxData_reg[6]/NET0131 ,
		_w11726_
	);
	LUT3 #(
		.INIT('h70)
	) name1214 (
		_w11655_,
		_w11657_,
		_w11726_,
		_w11727_
	);
	LUT4 #(
		.INIT('h57df)
	) name1215 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[22]/NET0131 ,
		\wishbone_TxDataLatched_reg[6]/NET0131 ,
		_w11728_
	);
	LUT4 #(
		.INIT('haebf)
	) name1216 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[14]/NET0131 ,
		\wishbone_TxDataLatched_reg[30]/NET0131 ,
		_w11729_
	);
	LUT2 #(
		.INIT('h8)
	) name1217 (
		_w11728_,
		_w11729_,
		_w11730_
	);
	LUT3 #(
		.INIT('h80)
	) name1218 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[30]/P0001 ,
		_w11731_
	);
	LUT3 #(
		.INIT('h13)
	) name1219 (
		_w11657_,
		_w11666_,
		_w11731_,
		_w11732_
	);
	LUT4 #(
		.INIT('h3100)
	) name1220 (
		_w11664_,
		_w11727_,
		_w11730_,
		_w11732_,
		_w11733_
	);
	LUT3 #(
		.INIT('h10)
	) name1221 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[30]/P0001 ,
		_w11734_
	);
	LUT3 #(
		.INIT('h40)
	) name1222 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[14]/P0001 ,
		_w11735_
	);
	LUT4 #(
		.INIT('h57df)
	) name1223 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[22]/P0001 ,
		\wishbone_tx_fifo_data_out_reg[6]/P0001 ,
		_w11736_
	);
	LUT4 #(
		.INIT('h0200)
	) name1224 (
		_w11666_,
		_w11734_,
		_w11735_,
		_w11736_,
		_w11737_
	);
	LUT2 #(
		.INIT('h1)
	) name1225 (
		_w11733_,
		_w11737_,
		_w11738_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1226 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_Flop_reg/NET0131 ,
		\wishbone_TxData_reg[5]/NET0131 ,
		_w11739_
	);
	LUT3 #(
		.INIT('h70)
	) name1227 (
		_w11655_,
		_w11657_,
		_w11739_,
		_w11740_
	);
	LUT4 #(
		.INIT('h57df)
	) name1228 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[21]/NET0131 ,
		\wishbone_TxDataLatched_reg[5]/NET0131 ,
		_w11741_
	);
	LUT4 #(
		.INIT('haebf)
	) name1229 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[13]/NET0131 ,
		\wishbone_TxDataLatched_reg[29]/NET0131 ,
		_w11742_
	);
	LUT2 #(
		.INIT('h8)
	) name1230 (
		_w11741_,
		_w11742_,
		_w11743_
	);
	LUT3 #(
		.INIT('h80)
	) name1231 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[29]/P0001 ,
		_w11744_
	);
	LUT3 #(
		.INIT('h13)
	) name1232 (
		_w11657_,
		_w11666_,
		_w11744_,
		_w11745_
	);
	LUT4 #(
		.INIT('h3100)
	) name1233 (
		_w11664_,
		_w11740_,
		_w11743_,
		_w11745_,
		_w11746_
	);
	LUT3 #(
		.INIT('h10)
	) name1234 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[29]/P0001 ,
		_w11747_
	);
	LUT3 #(
		.INIT('h40)
	) name1235 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[13]/P0001 ,
		_w11748_
	);
	LUT4 #(
		.INIT('h57df)
	) name1236 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[21]/P0001 ,
		\wishbone_tx_fifo_data_out_reg[5]/P0001 ,
		_w11749_
	);
	LUT4 #(
		.INIT('h0200)
	) name1237 (
		_w11666_,
		_w11747_,
		_w11748_,
		_w11749_,
		_w11750_
	);
	LUT2 #(
		.INIT('h1)
	) name1238 (
		_w11746_,
		_w11750_,
		_w11751_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1239 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_Flop_reg/NET0131 ,
		\wishbone_TxData_reg[7]/NET0131 ,
		_w11752_
	);
	LUT3 #(
		.INIT('h70)
	) name1240 (
		_w11655_,
		_w11657_,
		_w11752_,
		_w11753_
	);
	LUT4 #(
		.INIT('h57df)
	) name1241 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[23]/NET0131 ,
		\wishbone_TxDataLatched_reg[7]/NET0131 ,
		_w11754_
	);
	LUT4 #(
		.INIT('haebf)
	) name1242 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxDataLatched_reg[15]/NET0131 ,
		\wishbone_TxDataLatched_reg[31]/NET0131 ,
		_w11755_
	);
	LUT2 #(
		.INIT('h8)
	) name1243 (
		_w11754_,
		_w11755_,
		_w11756_
	);
	LUT3 #(
		.INIT('h80)
	) name1244 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[31]/P0001 ,
		_w11757_
	);
	LUT3 #(
		.INIT('h13)
	) name1245 (
		_w11657_,
		_w11666_,
		_w11757_,
		_w11758_
	);
	LUT4 #(
		.INIT('h3100)
	) name1246 (
		_w11664_,
		_w11753_,
		_w11756_,
		_w11758_,
		_w11759_
	);
	LUT3 #(
		.INIT('h10)
	) name1247 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[31]/P0001 ,
		_w11760_
	);
	LUT3 #(
		.INIT('h40)
	) name1248 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[15]/P0001 ,
		_w11761_
	);
	LUT4 #(
		.INIT('h57df)
	) name1249 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_tx_fifo_data_out_reg[23]/P0001 ,
		\wishbone_tx_fifo_data_out_reg[7]/P0001 ,
		_w11762_
	);
	LUT4 #(
		.INIT('h0200)
	) name1250 (
		_w11666_,
		_w11760_,
		_w11761_,
		_w11762_,
		_w11763_
	);
	LUT2 #(
		.INIT('h1)
	) name1251 (
		_w11759_,
		_w11763_,
		_w11764_
	);
	LUT3 #(
		.INIT('h7b)
	) name1252 (
		\rxethmac1_crcrx_Crc_reg[1]/NET0131 ,
		_w10582_,
		_w11420_,
		_w11765_
	);
	LUT2 #(
		.INIT('h2)
	) name1253 (
		\rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131 ,
		\rxethmac1_rxstatem1_StateDrop_reg/NET0131 ,
		_w11766_
	);
	LUT3 #(
		.INIT('h70)
	) name1254 (
		_w11548_,
		_w11638_,
		_w11766_,
		_w11767_
	);
	LUT2 #(
		.INIT('h1)
	) name1255 (
		\rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131 ,
		\rxethmac1_rxstatem1_StateDrop_reg/NET0131 ,
		_w11768_
	);
	LUT3 #(
		.INIT('h70)
	) name1256 (
		_w11548_,
		_w11638_,
		_w11768_,
		_w11769_
	);
	LUT3 #(
		.INIT('he4)
	) name1257 (
		_w11642_,
		_w11767_,
		_w11769_,
		_w11770_
	);
	LUT3 #(
		.INIT('h01)
	) name1258 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		_w11771_
	);
	LUT3 #(
		.INIT('h2a)
	) name1259 (
		_w10576_,
		_w11558_,
		_w11771_,
		_w11772_
	);
	LUT2 #(
		.INIT('h9)
	) name1260 (
		\txethmac1_txcrc_Crc_reg[30]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		_w11773_
	);
	LUT4 #(
		.INIT('h00f8)
	) name1261 (
		_w11026_,
		_w11027_,
		_w11028_,
		_w11773_,
		_w11774_
	);
	LUT4 #(
		.INIT('h0007)
	) name1262 (
		_w11026_,
		_w11027_,
		_w11028_,
		_w11773_,
		_w11775_
	);
	LUT4 #(
		.INIT('h096f)
	) name1263 (
		_w11000_,
		_w11004_,
		_w11774_,
		_w11775_,
		_w11776_
	);
	LUT4 #(
		.INIT('hf800)
	) name1264 (
		_w11026_,
		_w11027_,
		_w11028_,
		_w11773_,
		_w11777_
	);
	LUT4 #(
		.INIT('h0700)
	) name1265 (
		_w11026_,
		_w11027_,
		_w11028_,
		_w11773_,
		_w11778_
	);
	LUT4 #(
		.INIT('h069f)
	) name1266 (
		_w11000_,
		_w11004_,
		_w11777_,
		_w11778_,
		_w11779_
	);
	LUT4 #(
		.INIT('h1000)
	) name1267 (
		\txethmac1_txcrc_Crc_reg[6]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11776_,
		_w11779_,
		_w11780_
	);
	LUT3 #(
		.INIT('h40)
	) name1268 (
		\txethmac1_txcrc_Crc_reg[6]/NET0131 ,
		_w10913_,
		_w10914_,
		_w11781_
	);
	LUT4 #(
		.INIT('h4000)
	) name1269 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11007_,
		_w11776_,
		_w11779_,
		_w11782_
	);
	LUT3 #(
		.INIT('hab)
	) name1270 (
		_w11780_,
		_w11781_,
		_w11782_,
		_w11783_
	);
	LUT2 #(
		.INIT('h9)
	) name1271 (
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		_w11784_
	);
	LUT4 #(
		.INIT('h00ba)
	) name1272 (
		_w11011_,
		_w11012_,
		_w11013_,
		_w11784_,
		_w11785_
	);
	LUT4 #(
		.INIT('h0045)
	) name1273 (
		_w11011_,
		_w11012_,
		_w11013_,
		_w11784_,
		_w11786_
	);
	LUT4 #(
		.INIT('h096f)
	) name1274 (
		_w11000_,
		_w11004_,
		_w11785_,
		_w11786_,
		_w11787_
	);
	LUT4 #(
		.INIT('hba00)
	) name1275 (
		_w11011_,
		_w11012_,
		_w11013_,
		_w11784_,
		_w11788_
	);
	LUT4 #(
		.INIT('h4500)
	) name1276 (
		_w11011_,
		_w11012_,
		_w11013_,
		_w11784_,
		_w11789_
	);
	LUT4 #(
		.INIT('h069f)
	) name1277 (
		_w11000_,
		_w11004_,
		_w11788_,
		_w11789_,
		_w11790_
	);
	LUT4 #(
		.INIT('h1000)
	) name1278 (
		\txethmac1_txcrc_Crc_reg[7]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11787_,
		_w11790_,
		_w11791_
	);
	LUT3 #(
		.INIT('h40)
	) name1279 (
		\txethmac1_txcrc_Crc_reg[7]/NET0131 ,
		_w10913_,
		_w10914_,
		_w11792_
	);
	LUT4 #(
		.INIT('h4000)
	) name1280 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11007_,
		_w11787_,
		_w11790_,
		_w11793_
	);
	LUT3 #(
		.INIT('hab)
	) name1281 (
		_w11791_,
		_w11792_,
		_w11793_,
		_w11794_
	);
	LUT2 #(
		.INIT('h1)
	) name1282 (
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		\rxethmac1_rxaddrcheck1_RxAbort_reg/NET0131 ,
		_w11795_
	);
	LUT3 #(
		.INIT('h02)
	) name1283 (
		\rxethmac1_Broadcast_reg/NET0131 ,
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		\rxethmac1_rxaddrcheck1_RxAbort_reg/NET0131 ,
		_w11796_
	);
	LUT4 #(
		.INIT('h4000)
	) name1284 (
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		_w10515_,
		_w10516_,
		_w10517_,
		_w11797_
	);
	LUT4 #(
		.INIT('h8000)
	) name1285 (
		\rxethmac1_LatchedByte_reg[4]/NET0131 ,
		\rxethmac1_LatchedByte_reg[5]/NET0131 ,
		\rxethmac1_LatchedByte_reg[6]/NET0131 ,
		\rxethmac1_LatchedByte_reg[7]/NET0131 ,
		_w11798_
	);
	LUT2 #(
		.INIT('h2)
	) name1286 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w11799_
	);
	LUT4 #(
		.INIT('h0200)
	) name1287 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w11800_
	);
	LUT2 #(
		.INIT('h8)
	) name1288 (
		_w11798_,
		_w11800_,
		_w11801_
	);
	LUT3 #(
		.INIT('h15)
	) name1289 (
		_w11796_,
		_w11797_,
		_w11801_,
		_w11802_
	);
	LUT3 #(
		.INIT('h80)
	) name1290 (
		_w10515_,
		_w10516_,
		_w10517_,
		_w11803_
	);
	LUT4 #(
		.INIT('h8000)
	) name1291 (
		\rxethmac1_LatchedByte_reg[0]/NET0131 ,
		\rxethmac1_LatchedByte_reg[1]/NET0131 ,
		\rxethmac1_LatchedByte_reg[2]/NET0131 ,
		\rxethmac1_LatchedByte_reg[3]/NET0131 ,
		_w11804_
	);
	LUT4 #(
		.INIT('h0222)
	) name1292 (
		_w10534_,
		_w11610_,
		_w11798_,
		_w11804_,
		_w11805_
	);
	LUT2 #(
		.INIT('h8)
	) name1293 (
		_w11803_,
		_w11805_,
		_w11806_
	);
	LUT2 #(
		.INIT('h1)
	) name1294 (
		_w11802_,
		_w11806_,
		_w11807_
	);
	LUT4 #(
		.INIT('h0105)
	) name1295 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w11550_,
		_w11556_,
		_w11557_,
		_w11808_
	);
	LUT4 #(
		.INIT('h008f)
	) name1296 (
		_w10554_,
		_w10573_,
		_w11635_,
		_w11808_,
		_w11809_
	);
	LUT3 #(
		.INIT('h10)
	) name1297 (
		_w11555_,
		_w11559_,
		_w11809_,
		_w11810_
	);
	LUT4 #(
		.INIT('h8b8a)
	) name1298 (
		\rxethmac1_rxstatem1_StatePreamble_reg/NET0131 ,
		_w10576_,
		_w11561_,
		_w11562_,
		_w11811_
	);
	LUT2 #(
		.INIT('h4)
	) name1299 (
		_w11559_,
		_w11811_,
		_w11812_
	);
	LUT2 #(
		.INIT('h4)
	) name1300 (
		_w11555_,
		_w11812_,
		_w11813_
	);
	LUT4 #(
		.INIT('h4440)
	) name1301 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		_w11814_
	);
	LUT2 #(
		.INIT('h8)
	) name1302 (
		_w10519_,
		_w11814_,
		_w11815_
	);
	LUT3 #(
		.INIT('h54)
	) name1303 (
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		_w11816_
	);
	LUT2 #(
		.INIT('h8)
	) name1304 (
		_w10514_,
		_w11816_,
		_w11817_
	);
	LUT2 #(
		.INIT('h8)
	) name1305 (
		_w10533_,
		_w11817_,
		_w11818_
	);
	LUT4 #(
		.INIT('h8880)
	) name1306 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		_w11819_
	);
	LUT2 #(
		.INIT('h8)
	) name1307 (
		_w10519_,
		_w11819_,
		_w11820_
	);
	LUT4 #(
		.INIT('h8000)
	) name1308 (
		_w10533_,
		_w11516_,
		_w11521_,
		_w11817_,
		_w11821_
	);
	LUT3 #(
		.INIT('h04)
	) name1309 (
		_w11522_,
		_w11818_,
		_w11820_,
		_w11822_
	);
	LUT2 #(
		.INIT('h8)
	) name1310 (
		_w11799_,
		_w11816_,
		_w11823_
	);
	LUT2 #(
		.INIT('h8)
	) name1311 (
		_w10533_,
		_w11823_,
		_w11824_
	);
	LUT2 #(
		.INIT('h8)
	) name1312 (
		_w10535_,
		_w11816_,
		_w11825_
	);
	LUT4 #(
		.INIT('h8000)
	) name1313 (
		_w10533_,
		_w11504_,
		_w11509_,
		_w11825_,
		_w11826_
	);
	LUT2 #(
		.INIT('h8)
	) name1314 (
		_w11580_,
		_w11816_,
		_w11827_
	);
	LUT4 #(
		.INIT('h4e4c)
	) name1315 (
		_w10533_,
		_w11795_,
		_w11825_,
		_w11827_,
		_w11828_
	);
	LUT4 #(
		.INIT('h2a00)
	) name1316 (
		_w10533_,
		_w11493_,
		_w11498_,
		_w11827_,
		_w11829_
	);
	LUT4 #(
		.INIT('hbbab)
	) name1317 (
		_w11824_,
		_w11826_,
		_w11828_,
		_w11829_,
		_w11830_
	);
	LUT4 #(
		.INIT('h8000)
	) name1318 (
		_w10533_,
		_w11530_,
		_w11535_,
		_w11823_,
		_w11831_
	);
	LUT3 #(
		.INIT('h01)
	) name1319 (
		_w11820_,
		_w11821_,
		_w11831_,
		_w11832_
	);
	LUT4 #(
		.INIT('h2a00)
	) name1320 (
		_w10519_,
		_w11476_,
		_w11481_,
		_w11819_,
		_w11833_
	);
	LUT2 #(
		.INIT('h2)
	) name1321 (
		\rxethmac1_rxaddrcheck1_UnicastOK_reg/NET0131 ,
		_w11833_,
		_w11834_
	);
	LUT4 #(
		.INIT('h1500)
	) name1322 (
		_w11822_,
		_w11830_,
		_w11832_,
		_w11834_,
		_w11835_
	);
	LUT4 #(
		.INIT('h2a00)
	) name1323 (
		_w10519_,
		_w11462_,
		_w11467_,
		_w11814_,
		_w11836_
	);
	LUT3 #(
		.INIT('h0e)
	) name1324 (
		_w11815_,
		_w11835_,
		_w11836_,
		_w11837_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name1325 (
		\WillTransmit_q2_reg/P0001 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_rxstatem1_StateDrop_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		_w11838_
	);
	LUT3 #(
		.INIT('h70)
	) name1326 (
		_w11550_,
		_w11553_,
		_w11838_,
		_w11839_
	);
	LUT4 #(
		.INIT('h2033)
	) name1327 (
		_w10573_,
		_w10576_,
		_w11389_,
		_w11839_,
		_w11840_
	);
	LUT3 #(
		.INIT('h0b)
	) name1328 (
		\ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131 ,
		\rxethmac1_rxaddrcheck1_RxAbort_reg/NET0131 ,
		_w11841_
	);
	LUT2 #(
		.INIT('h4)
	) name1329 (
		\macstatus1_InvalidSymbol_reg/NET0131 ,
		\macstatus1_LatchedMRxErr_reg/NET0131 ,
		_w11842_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1330 (
		\RxAbortRst_reg/NET0131 ,
		\RxAbort_latch_reg/NET0131 ,
		\ethreg1_MODER_2_DataOut_reg[0]/NET0131 ,
		\macstatus1_ShortFrame_reg/NET0131 ,
		_w11843_
	);
	LUT3 #(
		.INIT('hdf)
	) name1331 (
		_w11841_,
		_w11842_,
		_w11843_,
		_w11844_
	);
	LUT4 #(
		.INIT('h8000)
	) name1332 (
		\m_wb_adr_o[2]_pad ,
		\m_wb_adr_o[3]_pad ,
		\m_wb_adr_o[4]_pad ,
		\m_wb_adr_o[5]_pad ,
		_w11845_
	);
	LUT3 #(
		.INIT('h80)
	) name1333 (
		\m_wb_adr_o[6]_pad ,
		\m_wb_adr_o[7]_pad ,
		\m_wb_adr_o[8]_pad ,
		_w11846_
	);
	LUT2 #(
		.INIT('h8)
	) name1334 (
		\m_wb_adr_o[10]_pad ,
		\m_wb_adr_o[9]_pad ,
		_w11847_
	);
	LUT3 #(
		.INIT('h80)
	) name1335 (
		\m_wb_adr_o[10]_pad ,
		\m_wb_adr_o[11]_pad ,
		\m_wb_adr_o[9]_pad ,
		_w11848_
	);
	LUT3 #(
		.INIT('h80)
	) name1336 (
		_w11845_,
		_w11846_,
		_w11848_,
		_w11849_
	);
	LUT4 #(
		.INIT('h8000)
	) name1337 (
		\m_wb_adr_o[12]_pad ,
		\m_wb_adr_o[13]_pad ,
		\m_wb_adr_o[14]_pad ,
		\m_wb_adr_o[15]_pad ,
		_w11850_
	);
	LUT4 #(
		.INIT('h8000)
	) name1338 (
		_w11845_,
		_w11846_,
		_w11848_,
		_w11850_,
		_w11851_
	);
	LUT4 #(
		.INIT('h8000)
	) name1339 (
		\m_wb_adr_o[16]_pad ,
		\m_wb_adr_o[17]_pad ,
		\m_wb_adr_o[18]_pad ,
		\m_wb_adr_o[19]_pad ,
		_w11852_
	);
	LUT2 #(
		.INIT('h8)
	) name1340 (
		_w11851_,
		_w11852_,
		_w11853_
	);
	LUT2 #(
		.INIT('h8)
	) name1341 (
		\m_wb_adr_o[20]_pad ,
		\m_wb_adr_o[21]_pad ,
		_w11854_
	);
	LUT3 #(
		.INIT('h80)
	) name1342 (
		\m_wb_adr_o[22]_pad ,
		\m_wb_adr_o[23]_pad ,
		\m_wb_adr_o[24]_pad ,
		_w11855_
	);
	LUT2 #(
		.INIT('h8)
	) name1343 (
		\m_wb_adr_o[25]_pad ,
		\m_wb_adr_o[26]_pad ,
		_w11856_
	);
	LUT3 #(
		.INIT('h80)
	) name1344 (
		_w11854_,
		_w11855_,
		_w11856_,
		_w11857_
	);
	LUT3 #(
		.INIT('h80)
	) name1345 (
		_w11851_,
		_w11852_,
		_w11857_,
		_w11858_
	);
	LUT2 #(
		.INIT('h8)
	) name1346 (
		\m_wb_adr_o[27]_pad ,
		\m_wb_adr_o[28]_pad ,
		_w11859_
	);
	LUT3 #(
		.INIT('h80)
	) name1347 (
		\m_wb_adr_o[27]_pad ,
		\m_wb_adr_o[28]_pad ,
		\m_wb_adr_o[29]_pad ,
		_w11860_
	);
	LUT4 #(
		.INIT('h8000)
	) name1348 (
		_w11851_,
		_w11852_,
		_w11857_,
		_w11860_,
		_w11861_
	);
	LUT2 #(
		.INIT('h1)
	) name1349 (
		\m_wb_adr_o[30]_pad ,
		_w11861_,
		_w11862_
	);
	LUT4 #(
		.INIT('h8000)
	) name1350 (
		\m_wb_adr_o[27]_pad ,
		\m_wb_adr_o[28]_pad ,
		\m_wb_adr_o[29]_pad ,
		\m_wb_adr_o[30]_pad ,
		_w11863_
	);
	LUT4 #(
		.INIT('h8000)
	) name1351 (
		_w11851_,
		_w11852_,
		_w11857_,
		_w11863_,
		_w11864_
	);
	LUT2 #(
		.INIT('h1)
	) name1352 (
		\wishbone_rx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[1]/NET0131 ,
		_w11865_
	);
	LUT3 #(
		.INIT('h01)
	) name1353 (
		\wishbone_rx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[1]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[2]/NET0131 ,
		_w11866_
	);
	LUT2 #(
		.INIT('h1)
	) name1354 (
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[4]/NET0131 ,
		_w11867_
	);
	LUT2 #(
		.INIT('h1)
	) name1355 (
		m_wb_ack_i_pad,
		m_wb_err_i_pad,
		_w11868_
	);
	LUT4 #(
		.INIT('h1fef)
	) name1356 (
		m_wb_ack_i_pad,
		m_wb_err_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w11869_
	);
	LUT4 #(
		.INIT('h2a00)
	) name1357 (
		\wishbone_rx_burst_en_reg/NET0131 ,
		_w11866_,
		_w11867_,
		_w11869_,
		_w11870_
	);
	LUT2 #(
		.INIT('h4)
	) name1358 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w11871_
	);
	LUT3 #(
		.INIT('h0e)
	) name1359 (
		m_wb_ack_i_pad,
		m_wb_err_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		_w11872_
	);
	LUT3 #(
		.INIT('h09)
	) name1360 (
		\wishbone_MasterWbTX_reg/NET0131 ,
		_w11871_,
		_w11872_,
		_w11873_
	);
	LUT4 #(
		.INIT('h0001)
	) name1361 (
		\wishbone_RxPointerMSB_reg[30]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w11874_
	);
	LUT3 #(
		.INIT('h40)
	) name1362 (
		\wishbone_BlockReadTxDataFromMemory_reg/NET0131 ,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_ReadTxDataFromMemory_reg/NET0131 ,
		_w11875_
	);
	LUT2 #(
		.INIT('h8)
	) name1363 (
		_w11868_,
		_w11875_,
		_w11876_
	);
	LUT3 #(
		.INIT('h13)
	) name1364 (
		_w11868_,
		_w11874_,
		_w11875_,
		_w11877_
	);
	LUT3 #(
		.INIT('h80)
	) name1365 (
		_w11870_,
		_w11873_,
		_w11877_,
		_w11878_
	);
	LUT4 #(
		.INIT('h1001)
	) name1366 (
		m_wb_ack_i_pad,
		m_wb_err_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w11879_
	);
	LUT3 #(
		.INIT('h40)
	) name1367 (
		\wishbone_BlockReadTxDataFromMemory_reg/NET0131 ,
		\wishbone_ReadTxDataFromMemory_reg/NET0131 ,
		\wishbone_tx_burst_en_reg/NET0131 ,
		_w11880_
	);
	LUT4 #(
		.INIT('hfef1)
	) name1368 (
		m_wb_ack_i_pad,
		m_wb_err_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w11881_
	);
	LUT4 #(
		.INIT('hbf1f)
	) name1369 (
		\wishbone_MasterWbTX_reg/NET0131 ,
		_w11879_,
		_w11880_,
		_w11881_,
		_w11882_
	);
	LUT3 #(
		.INIT('h01)
	) name1370 (
		m_wb_ack_i_pad,
		m_wb_err_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		_w11883_
	);
	LUT3 #(
		.INIT('h70)
	) name1371 (
		_w11866_,
		_w11867_,
		_w11883_,
		_w11884_
	);
	LUT3 #(
		.INIT('h01)
	) name1372 (
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w11885_
	);
	LUT4 #(
		.INIT('h008f)
	) name1373 (
		_w11866_,
		_w11867_,
		_w11883_,
		_w11885_,
		_w11886_
	);
	LUT2 #(
		.INIT('h4)
	) name1374 (
		_w11882_,
		_w11886_,
		_w11887_
	);
	LUT3 #(
		.INIT('h54)
	) name1375 (
		_w11864_,
		_w11878_,
		_w11887_,
		_w11888_
	);
	LUT2 #(
		.INIT('h4)
	) name1376 (
		_w11862_,
		_w11888_,
		_w11889_
	);
	LUT2 #(
		.INIT('h1)
	) name1377 (
		_w11882_,
		_w11884_,
		_w11890_
	);
	LUT3 #(
		.INIT('h04)
	) name1378 (
		\wishbone_BlockReadTxDataFromMemory_reg/NET0131 ,
		\wishbone_ReadTxDataFromMemory_reg/NET0131 ,
		\wishbone_tx_burst_en_reg/NET0131 ,
		_w11891_
	);
	LUT2 #(
		.INIT('h1)
	) name1379 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_MasterWbTX_reg/NET0131 ,
		_w11892_
	);
	LUT3 #(
		.INIT('h01)
	) name1380 (
		m_wb_ack_i_pad,
		m_wb_err_i_pad,
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w11893_
	);
	LUT2 #(
		.INIT('h8)
	) name1381 (
		_w11892_,
		_w11893_,
		_w11894_
	);
	LUT4 #(
		.INIT('h8000)
	) name1382 (
		_w11866_,
		_w11867_,
		_w11892_,
		_w11893_,
		_w11895_
	);
	LUT3 #(
		.INIT('h15)
	) name1383 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		_w11866_,
		_w11867_,
		_w11896_
	);
	LUT3 #(
		.INIT('h10)
	) name1384 (
		m_wb_ack_i_pad,
		m_wb_err_i_pad,
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w11897_
	);
	LUT2 #(
		.INIT('h6)
	) name1385 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_MasterWbTX_reg/NET0131 ,
		_w11898_
	);
	LUT2 #(
		.INIT('h8)
	) name1386 (
		_w11897_,
		_w11898_,
		_w11899_
	);
	LUT4 #(
		.INIT('h7577)
	) name1387 (
		_w11891_,
		_w11895_,
		_w11896_,
		_w11899_,
		_w11900_
	);
	LUT2 #(
		.INIT('h4)
	) name1388 (
		_w11890_,
		_w11900_,
		_w11901_
	);
	LUT3 #(
		.INIT('h08)
	) name1389 (
		_w11870_,
		_w11873_,
		_w11876_,
		_w11902_
	);
	LUT3 #(
		.INIT('h15)
	) name1390 (
		\wishbone_rx_burst_en_reg/NET0131 ,
		_w11866_,
		_w11867_,
		_w11903_
	);
	LUT3 #(
		.INIT('h40)
	) name1391 (
		_w11875_,
		_w11897_,
		_w11898_,
		_w11904_
	);
	LUT3 #(
		.INIT('hc8)
	) name1392 (
		_w11894_,
		_w11903_,
		_w11904_,
		_w11905_
	);
	LUT2 #(
		.INIT('h1)
	) name1393 (
		_w11902_,
		_w11905_,
		_w11906_
	);
	LUT4 #(
		.INIT('h0004)
	) name1394 (
		_w11890_,
		_w11900_,
		_w11902_,
		_w11905_,
		_w11907_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1395 (
		_w11866_,
		_w11867_,
		_w11883_,
		_w11885_,
		_w11908_
	);
	LUT2 #(
		.INIT('h4)
	) name1396 (
		_w11882_,
		_w11908_,
		_w11909_
	);
	LUT3 #(
		.INIT('ha2)
	) name1397 (
		\wishbone_TxPointerMSB_reg[30]/NET0131 ,
		_w11900_,
		_w11909_,
		_w11910_
	);
	LUT3 #(
		.INIT('h01)
	) name1398 (
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w11911_
	);
	LUT4 #(
		.INIT('h00ea)
	) name1399 (
		\wishbone_rx_burst_en_reg/NET0131 ,
		_w11866_,
		_w11867_,
		_w11911_,
		_w11912_
	);
	LUT3 #(
		.INIT('h07)
	) name1400 (
		_w11892_,
		_w11893_,
		_w11911_,
		_w11913_
	);
	LUT3 #(
		.INIT('h23)
	) name1401 (
		_w11904_,
		_w11912_,
		_w11913_,
		_w11914_
	);
	LUT4 #(
		.INIT('h080a)
	) name1402 (
		\wishbone_RxPointerMSB_reg[30]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w11915_
	);
	LUT3 #(
		.INIT('he0)
	) name1403 (
		_w11902_,
		_w11905_,
		_w11915_,
		_w11916_
	);
	LUT4 #(
		.INIT('h0007)
	) name1404 (
		\m_wb_adr_o[30]_pad ,
		_w11907_,
		_w11910_,
		_w11916_,
		_w11917_
	);
	LUT2 #(
		.INIT('hb)
	) name1405 (
		_w11889_,
		_w11917_,
		_w11918_
	);
	LUT3 #(
		.INIT('h08)
	) name1406 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11919_
	);
	LUT4 #(
		.INIT('h070f)
	) name1407 (
		_w11455_,
		_w11456_,
		_w11482_,
		_w11919_,
		_w11920_
	);
	LUT4 #(
		.INIT('h1000)
	) name1408 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w11921_
	);
	LUT4 #(
		.INIT('h2a7f)
	) name1409 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		_w11486_,
		_w11921_,
		_w11922_
	);
	LUT3 #(
		.INIT('ha2)
	) name1410 (
		\maccontrol1_receivecontrol1_OpCodeOK_reg/NET0131 ,
		_w11920_,
		_w11922_,
		_w11923_
	);
	LUT2 #(
		.INIT('h8)
	) name1411 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		_w11486_,
		_w11924_
	);
	LUT4 #(
		.INIT('h0004)
	) name1412 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11925_
	);
	LUT3 #(
		.INIT('h80)
	) name1413 (
		_w11455_,
		_w11456_,
		_w11925_,
		_w11926_
	);
	LUT2 #(
		.INIT('h8)
	) name1414 (
		_w11924_,
		_w11926_,
		_w11927_
	);
	LUT2 #(
		.INIT('he)
	) name1415 (
		_w11923_,
		_w11927_,
		_w11928_
	);
	LUT4 #(
		.INIT('h0010)
	) name1416 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11929_
	);
	LUT4 #(
		.INIT('h0400)
	) name1417 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w11930_
	);
	LUT3 #(
		.INIT('h80)
	) name1418 (
		\wishbone_bd_ram_mem3_reg[164][28]/P0001 ,
		_w11929_,
		_w11930_,
		_w11931_
	);
	LUT4 #(
		.INIT('h0001)
	) name1419 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w11932_
	);
	LUT4 #(
		.INIT('h0020)
	) name1420 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11933_
	);
	LUT3 #(
		.INIT('h80)
	) name1421 (
		\wishbone_bd_ram_mem3_reg[5][28]/P0001 ,
		_w11932_,
		_w11933_,
		_w11934_
	);
	LUT4 #(
		.INIT('h0002)
	) name1422 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w11935_
	);
	LUT4 #(
		.INIT('h0800)
	) name1423 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11936_
	);
	LUT3 #(
		.INIT('h80)
	) name1424 (
		\wishbone_bd_ram_mem3_reg[27][28]/P0001 ,
		_w11935_,
		_w11936_,
		_w11937_
	);
	LUT4 #(
		.INIT('h0008)
	) name1425 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11938_
	);
	LUT3 #(
		.INIT('h80)
	) name1426 (
		\wishbone_bd_ram_mem3_reg[163][28]/P0001 ,
		_w11930_,
		_w11938_,
		_w11939_
	);
	LUT4 #(
		.INIT('h0001)
	) name1427 (
		_w11931_,
		_w11934_,
		_w11937_,
		_w11939_,
		_w11940_
	);
	LUT4 #(
		.INIT('h0001)
	) name1428 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11941_
	);
	LUT4 #(
		.INIT('h0800)
	) name1429 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w11942_
	);
	LUT3 #(
		.INIT('h80)
	) name1430 (
		\wishbone_bd_ram_mem3_reg[176][28]/P0001 ,
		_w11941_,
		_w11942_,
		_w11943_
	);
	LUT4 #(
		.INIT('h0400)
	) name1431 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11944_
	);
	LUT4 #(
		.INIT('h1000)
	) name1432 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w11945_
	);
	LUT3 #(
		.INIT('h80)
	) name1433 (
		\wishbone_bd_ram_mem3_reg[202][28]/P0001 ,
		_w11944_,
		_w11945_,
		_w11946_
	);
	LUT3 #(
		.INIT('h80)
	) name1434 (
		\wishbone_bd_ram_mem3_reg[160][28]/P0001 ,
		_w11930_,
		_w11941_,
		_w11947_
	);
	LUT4 #(
		.INIT('h4000)
	) name1435 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11948_
	);
	LUT4 #(
		.INIT('h0010)
	) name1436 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w11949_
	);
	LUT3 #(
		.INIT('h80)
	) name1437 (
		\wishbone_bd_ram_mem3_reg[78][28]/P0001 ,
		_w11948_,
		_w11949_,
		_w11950_
	);
	LUT4 #(
		.INIT('h0001)
	) name1438 (
		_w11943_,
		_w11946_,
		_w11947_,
		_w11950_,
		_w11951_
	);
	LUT4 #(
		.INIT('h8000)
	) name1439 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w11952_
	);
	LUT3 #(
		.INIT('h80)
	) name1440 (
		\wishbone_bd_ram_mem3_reg[254][28]/P0001 ,
		_w11948_,
		_w11952_,
		_w11953_
	);
	LUT4 #(
		.INIT('h1000)
	) name1441 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11954_
	);
	LUT4 #(
		.INIT('h0100)
	) name1442 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w11955_
	);
	LUT3 #(
		.INIT('h80)
	) name1443 (
		\wishbone_bd_ram_mem3_reg[140][28]/P0001 ,
		_w11954_,
		_w11955_,
		_w11956_
	);
	LUT4 #(
		.INIT('h0004)
	) name1444 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w11957_
	);
	LUT3 #(
		.INIT('h80)
	) name1445 (
		\wishbone_bd_ram_mem3_reg[44][28]/P0001 ,
		_w11954_,
		_w11957_,
		_w11958_
	);
	LUT4 #(
		.INIT('h0200)
	) name1446 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w11959_
	);
	LUT3 #(
		.INIT('h80)
	) name1447 (
		\wishbone_bd_ram_mem3_reg[158][28]/P0001 ,
		_w11948_,
		_w11959_,
		_w11960_
	);
	LUT4 #(
		.INIT('h0001)
	) name1448 (
		_w11953_,
		_w11956_,
		_w11958_,
		_w11960_,
		_w11961_
	);
	LUT3 #(
		.INIT('h80)
	) name1449 (
		\wishbone_bd_ram_mem3_reg[46][28]/P0001 ,
		_w11948_,
		_w11957_,
		_w11962_
	);
	LUT4 #(
		.INIT('h0004)
	) name1450 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11963_
	);
	LUT3 #(
		.INIT('h80)
	) name1451 (
		\wishbone_bd_ram_mem3_reg[178][28]/P0001 ,
		_w11942_,
		_w11963_,
		_w11964_
	);
	LUT4 #(
		.INIT('h0040)
	) name1452 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w11965_
	);
	LUT4 #(
		.INIT('h2000)
	) name1453 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11966_
	);
	LUT3 #(
		.INIT('h80)
	) name1454 (
		\wishbone_bd_ram_mem3_reg[109][28]/P0001 ,
		_w11965_,
		_w11966_,
		_w11967_
	);
	LUT4 #(
		.INIT('h0200)
	) name1455 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11968_
	);
	LUT3 #(
		.INIT('h80)
	) name1456 (
		\wishbone_bd_ram_mem3_reg[153][28]/P0001 ,
		_w11959_,
		_w11968_,
		_w11969_
	);
	LUT4 #(
		.INIT('h0001)
	) name1457 (
		_w11962_,
		_w11964_,
		_w11967_,
		_w11969_,
		_w11970_
	);
	LUT4 #(
		.INIT('h8000)
	) name1458 (
		_w11940_,
		_w11951_,
		_w11961_,
		_w11970_,
		_w11971_
	);
	LUT4 #(
		.INIT('h0020)
	) name1459 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w11972_
	);
	LUT4 #(
		.INIT('h8000)
	) name1460 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11973_
	);
	LUT3 #(
		.INIT('h80)
	) name1461 (
		\wishbone_bd_ram_mem3_reg[95][28]/P0001 ,
		_w11972_,
		_w11973_,
		_w11974_
	);
	LUT4 #(
		.INIT('h0080)
	) name1462 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11975_
	);
	LUT3 #(
		.INIT('h80)
	) name1463 (
		\wishbone_bd_ram_mem3_reg[103][28]/P0001 ,
		_w11965_,
		_w11975_,
		_w11976_
	);
	LUT4 #(
		.INIT('h0002)
	) name1464 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11977_
	);
	LUT3 #(
		.INIT('h80)
	) name1465 (
		\wishbone_bd_ram_mem3_reg[17][28]/P0001 ,
		_w11935_,
		_w11977_,
		_w11978_
	);
	LUT4 #(
		.INIT('h0008)
	) name1466 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w11979_
	);
	LUT3 #(
		.INIT('h80)
	) name1467 (
		\wishbone_bd_ram_mem3_reg[63][28]/P0001 ,
		_w11973_,
		_w11979_,
		_w11980_
	);
	LUT4 #(
		.INIT('h0001)
	) name1468 (
		_w11974_,
		_w11976_,
		_w11978_,
		_w11980_,
		_w11981_
	);
	LUT4 #(
		.INIT('h4000)
	) name1469 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w11982_
	);
	LUT3 #(
		.INIT('h80)
	) name1470 (
		\wishbone_bd_ram_mem3_reg[233][28]/P0001 ,
		_w11968_,
		_w11982_,
		_w11983_
	);
	LUT4 #(
		.INIT('h2000)
	) name1471 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w11984_
	);
	LUT3 #(
		.INIT('h80)
	) name1472 (
		\wishbone_bd_ram_mem3_reg[223][28]/P0001 ,
		_w11973_,
		_w11984_,
		_w11985_
	);
	LUT4 #(
		.INIT('h0040)
	) name1473 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11986_
	);
	LUT3 #(
		.INIT('h80)
	) name1474 (
		\wishbone_bd_ram_mem3_reg[70][28]/P0001 ,
		_w11949_,
		_w11986_,
		_w11987_
	);
	LUT3 #(
		.INIT('h80)
	) name1475 (
		\wishbone_bd_ram_mem3_reg[42][28]/P0001 ,
		_w11944_,
		_w11957_,
		_w11988_
	);
	LUT4 #(
		.INIT('h0001)
	) name1476 (
		_w11983_,
		_w11985_,
		_w11987_,
		_w11988_,
		_w11989_
	);
	LUT4 #(
		.INIT('h0100)
	) name1477 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w11990_
	);
	LUT3 #(
		.INIT('h80)
	) name1478 (
		\wishbone_bd_ram_mem3_reg[88][28]/P0001 ,
		_w11972_,
		_w11990_,
		_w11991_
	);
	LUT3 #(
		.INIT('h80)
	) name1479 (
		\wishbone_bd_ram_mem3_reg[239][28]/P0001 ,
		_w11973_,
		_w11982_,
		_w11992_
	);
	LUT3 #(
		.INIT('h80)
	) name1480 (
		\wishbone_bd_ram_mem3_reg[240][28]/P0001 ,
		_w11941_,
		_w11952_,
		_w11993_
	);
	LUT3 #(
		.INIT('h80)
	) name1481 (
		\wishbone_bd_ram_mem3_reg[3][28]/P0001 ,
		_w11932_,
		_w11938_,
		_w11994_
	);
	LUT4 #(
		.INIT('h0001)
	) name1482 (
		_w11991_,
		_w11992_,
		_w11993_,
		_w11994_,
		_w11995_
	);
	LUT3 #(
		.INIT('h80)
	) name1483 (
		\wishbone_bd_ram_mem3_reg[131][28]/P0001 ,
		_w11938_,
		_w11955_,
		_w11996_
	);
	LUT3 #(
		.INIT('h80)
	) name1484 (
		\wishbone_bd_ram_mem3_reg[173][28]/P0001 ,
		_w11930_,
		_w11966_,
		_w11997_
	);
	LUT3 #(
		.INIT('h80)
	) name1485 (
		\wishbone_bd_ram_mem3_reg[231][28]/P0001 ,
		_w11975_,
		_w11982_,
		_w11998_
	);
	LUT3 #(
		.INIT('h80)
	) name1486 (
		\wishbone_bd_ram_mem3_reg[190][28]/P0001 ,
		_w11942_,
		_w11948_,
		_w11999_
	);
	LUT4 #(
		.INIT('h0001)
	) name1487 (
		_w11996_,
		_w11997_,
		_w11998_,
		_w11999_,
		_w12000_
	);
	LUT4 #(
		.INIT('h8000)
	) name1488 (
		_w11981_,
		_w11989_,
		_w11995_,
		_w12000_,
		_w12001_
	);
	LUT3 #(
		.INIT('h80)
	) name1489 (
		\wishbone_bd_ram_mem3_reg[185][28]/P0001 ,
		_w11942_,
		_w11968_,
		_w12002_
	);
	LUT3 #(
		.INIT('h80)
	) name1490 (
		\wishbone_bd_ram_mem3_reg[82][28]/P0001 ,
		_w11963_,
		_w11972_,
		_w12003_
	);
	LUT3 #(
		.INIT('h80)
	) name1491 (
		\wishbone_bd_ram_mem3_reg[172][28]/P0001 ,
		_w11930_,
		_w11954_,
		_w12004_
	);
	LUT3 #(
		.INIT('h80)
	) name1492 (
		\wishbone_bd_ram_mem3_reg[68][28]/P0001 ,
		_w11929_,
		_w11949_,
		_w12005_
	);
	LUT4 #(
		.INIT('h0001)
	) name1493 (
		_w12002_,
		_w12003_,
		_w12004_,
		_w12005_,
		_w12006_
	);
	LUT3 #(
		.INIT('h80)
	) name1494 (
		\wishbone_bd_ram_mem3_reg[242][28]/P0001 ,
		_w11952_,
		_w11963_,
		_w12007_
	);
	LUT3 #(
		.INIT('h80)
	) name1495 (
		\wishbone_bd_ram_mem3_reg[84][28]/P0001 ,
		_w11929_,
		_w11972_,
		_w12008_
	);
	LUT3 #(
		.INIT('h80)
	) name1496 (
		\wishbone_bd_ram_mem3_reg[227][28]/P0001 ,
		_w11938_,
		_w11982_,
		_w12009_
	);
	LUT3 #(
		.INIT('h80)
	) name1497 (
		\wishbone_bd_ram_mem3_reg[192][28]/P0001 ,
		_w11941_,
		_w11945_,
		_w12010_
	);
	LUT4 #(
		.INIT('h0001)
	) name1498 (
		_w12007_,
		_w12008_,
		_w12009_,
		_w12010_,
		_w12011_
	);
	LUT4 #(
		.INIT('h0080)
	) name1499 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w12012_
	);
	LUT3 #(
		.INIT('h80)
	) name1500 (
		\wishbone_bd_ram_mem3_reg[125][28]/P0001 ,
		_w11966_,
		_w12012_,
		_w12013_
	);
	LUT3 #(
		.INIT('h80)
	) name1501 (
		\wishbone_bd_ram_mem3_reg[138][28]/P0001 ,
		_w11944_,
		_w11955_,
		_w12014_
	);
	LUT3 #(
		.INIT('h80)
	) name1502 (
		\wishbone_bd_ram_mem3_reg[100][28]/P0001 ,
		_w11929_,
		_w11965_,
		_w12015_
	);
	LUT3 #(
		.INIT('h80)
	) name1503 (
		\wishbone_bd_ram_mem3_reg[154][28]/P0001 ,
		_w11944_,
		_w11959_,
		_w12016_
	);
	LUT4 #(
		.INIT('h0001)
	) name1504 (
		_w12013_,
		_w12014_,
		_w12015_,
		_w12016_,
		_w12017_
	);
	LUT3 #(
		.INIT('h80)
	) name1505 (
		\wishbone_bd_ram_mem3_reg[188][28]/P0001 ,
		_w11942_,
		_w11954_,
		_w12018_
	);
	LUT3 #(
		.INIT('h80)
	) name1506 (
		\wishbone_bd_ram_mem3_reg[81][28]/P0001 ,
		_w11972_,
		_w11977_,
		_w12019_
	);
	LUT3 #(
		.INIT('h80)
	) name1507 (
		\wishbone_bd_ram_mem3_reg[29][28]/P0001 ,
		_w11935_,
		_w11966_,
		_w12020_
	);
	LUT3 #(
		.INIT('h80)
	) name1508 (
		\wishbone_bd_ram_mem3_reg[206][28]/P0001 ,
		_w11945_,
		_w11948_,
		_w12021_
	);
	LUT4 #(
		.INIT('h0001)
	) name1509 (
		_w12018_,
		_w12019_,
		_w12020_,
		_w12021_,
		_w12022_
	);
	LUT4 #(
		.INIT('h8000)
	) name1510 (
		_w12006_,
		_w12011_,
		_w12017_,
		_w12022_,
		_w12023_
	);
	LUT3 #(
		.INIT('h80)
	) name1511 (
		\wishbone_bd_ram_mem3_reg[45][28]/P0001 ,
		_w11957_,
		_w11966_,
		_w12024_
	);
	LUT3 #(
		.INIT('h80)
	) name1512 (
		\wishbone_bd_ram_mem3_reg[171][28]/P0001 ,
		_w11930_,
		_w11936_,
		_w12025_
	);
	LUT3 #(
		.INIT('h80)
	) name1513 (
		\wishbone_bd_ram_mem3_reg[96][28]/P0001 ,
		_w11941_,
		_w11965_,
		_w12026_
	);
	LUT3 #(
		.INIT('h80)
	) name1514 (
		\wishbone_bd_ram_mem3_reg[130][28]/P0001 ,
		_w11955_,
		_w11963_,
		_w12027_
	);
	LUT4 #(
		.INIT('h0001)
	) name1515 (
		_w12024_,
		_w12025_,
		_w12026_,
		_w12027_,
		_w12028_
	);
	LUT3 #(
		.INIT('h80)
	) name1516 (
		\wishbone_bd_ram_mem3_reg[249][28]/P0001 ,
		_w11952_,
		_w11968_,
		_w12029_
	);
	LUT3 #(
		.INIT('h80)
	) name1517 (
		\wishbone_bd_ram_mem3_reg[224][28]/P0001 ,
		_w11941_,
		_w11982_,
		_w12030_
	);
	LUT3 #(
		.INIT('h80)
	) name1518 (
		\wishbone_bd_ram_mem3_reg[47][28]/P0001 ,
		_w11957_,
		_w11973_,
		_w12031_
	);
	LUT3 #(
		.INIT('h80)
	) name1519 (
		\wishbone_bd_ram_mem3_reg[21][28]/P0001 ,
		_w11933_,
		_w11935_,
		_w12032_
	);
	LUT4 #(
		.INIT('h0001)
	) name1520 (
		_w12029_,
		_w12030_,
		_w12031_,
		_w12032_,
		_w12033_
	);
	LUT3 #(
		.INIT('h80)
	) name1521 (
		\wishbone_bd_ram_mem3_reg[210][28]/P0001 ,
		_w11963_,
		_w11984_,
		_w12034_
	);
	LUT3 #(
		.INIT('h80)
	) name1522 (
		\wishbone_bd_ram_mem3_reg[157][28]/P0001 ,
		_w11959_,
		_w11966_,
		_w12035_
	);
	LUT3 #(
		.INIT('h80)
	) name1523 (
		\wishbone_bd_ram_mem3_reg[142][28]/P0001 ,
		_w11948_,
		_w11955_,
		_w12036_
	);
	LUT3 #(
		.INIT('h80)
	) name1524 (
		\wishbone_bd_ram_mem3_reg[34][28]/P0001 ,
		_w11957_,
		_w11963_,
		_w12037_
	);
	LUT4 #(
		.INIT('h0001)
	) name1525 (
		_w12034_,
		_w12035_,
		_w12036_,
		_w12037_,
		_w12038_
	);
	LUT3 #(
		.INIT('h80)
	) name1526 (
		\wishbone_bd_ram_mem3_reg[83][28]/P0001 ,
		_w11938_,
		_w11972_,
		_w12039_
	);
	LUT3 #(
		.INIT('h80)
	) name1527 (
		\wishbone_bd_ram_mem3_reg[73][28]/P0001 ,
		_w11949_,
		_w11968_,
		_w12040_
	);
	LUT3 #(
		.INIT('h80)
	) name1528 (
		\wishbone_bd_ram_mem3_reg[8][28]/P0001 ,
		_w11932_,
		_w11990_,
		_w12041_
	);
	LUT3 #(
		.INIT('h80)
	) name1529 (
		\wishbone_bd_ram_mem3_reg[143][28]/P0001 ,
		_w11955_,
		_w11973_,
		_w12042_
	);
	LUT4 #(
		.INIT('h0001)
	) name1530 (
		_w12039_,
		_w12040_,
		_w12041_,
		_w12042_,
		_w12043_
	);
	LUT4 #(
		.INIT('h8000)
	) name1531 (
		_w12028_,
		_w12033_,
		_w12038_,
		_w12043_,
		_w12044_
	);
	LUT4 #(
		.INIT('h8000)
	) name1532 (
		_w11971_,
		_w12001_,
		_w12023_,
		_w12044_,
		_w12045_
	);
	LUT3 #(
		.INIT('h80)
	) name1533 (
		\wishbone_bd_ram_mem3_reg[149][28]/P0001 ,
		_w11933_,
		_w11959_,
		_w12046_
	);
	LUT3 #(
		.INIT('h80)
	) name1534 (
		\wishbone_bd_ram_mem3_reg[111][28]/P0001 ,
		_w11965_,
		_w11973_,
		_w12047_
	);
	LUT3 #(
		.INIT('h80)
	) name1535 (
		\wishbone_bd_ram_mem3_reg[244][28]/P0001 ,
		_w11929_,
		_w11952_,
		_w12048_
	);
	LUT3 #(
		.INIT('h80)
	) name1536 (
		\wishbone_bd_ram_mem3_reg[107][28]/P0001 ,
		_w11936_,
		_w11965_,
		_w12049_
	);
	LUT4 #(
		.INIT('h0001)
	) name1537 (
		_w12046_,
		_w12047_,
		_w12048_,
		_w12049_,
		_w12050_
	);
	LUT3 #(
		.INIT('h80)
	) name1538 (
		\wishbone_bd_ram_mem3_reg[236][28]/P0001 ,
		_w11954_,
		_w11982_,
		_w12051_
	);
	LUT3 #(
		.INIT('h80)
	) name1539 (
		\wishbone_bd_ram_mem3_reg[112][28]/P0001 ,
		_w11941_,
		_w12012_,
		_w12052_
	);
	LUT3 #(
		.INIT('h80)
	) name1540 (
		\wishbone_bd_ram_mem3_reg[86][28]/P0001 ,
		_w11972_,
		_w11986_,
		_w12053_
	);
	LUT3 #(
		.INIT('h80)
	) name1541 (
		\wishbone_bd_ram_mem3_reg[69][28]/P0001 ,
		_w11933_,
		_w11949_,
		_w12054_
	);
	LUT4 #(
		.INIT('h0001)
	) name1542 (
		_w12051_,
		_w12052_,
		_w12053_,
		_w12054_,
		_w12055_
	);
	LUT3 #(
		.INIT('h80)
	) name1543 (
		\wishbone_bd_ram_mem3_reg[133][28]/P0001 ,
		_w11933_,
		_w11955_,
		_w12056_
	);
	LUT3 #(
		.INIT('h80)
	) name1544 (
		\wishbone_bd_ram_mem3_reg[134][28]/P0001 ,
		_w11955_,
		_w11986_,
		_w12057_
	);
	LUT3 #(
		.INIT('h80)
	) name1545 (
		\wishbone_bd_ram_mem3_reg[228][28]/P0001 ,
		_w11929_,
		_w11982_,
		_w12058_
	);
	LUT3 #(
		.INIT('h80)
	) name1546 (
		\wishbone_bd_ram_mem3_reg[199][28]/P0001 ,
		_w11945_,
		_w11975_,
		_w12059_
	);
	LUT4 #(
		.INIT('h0001)
	) name1547 (
		_w12056_,
		_w12057_,
		_w12058_,
		_w12059_,
		_w12060_
	);
	LUT3 #(
		.INIT('h80)
	) name1548 (
		\wishbone_bd_ram_mem3_reg[105][28]/P0001 ,
		_w11965_,
		_w11968_,
		_w12061_
	);
	LUT3 #(
		.INIT('h80)
	) name1549 (
		\wishbone_bd_ram_mem3_reg[161][28]/P0001 ,
		_w11930_,
		_w11977_,
		_w12062_
	);
	LUT3 #(
		.INIT('h80)
	) name1550 (
		\wishbone_bd_ram_mem3_reg[144][28]/P0001 ,
		_w11941_,
		_w11959_,
		_w12063_
	);
	LUT3 #(
		.INIT('h80)
	) name1551 (
		\wishbone_bd_ram_mem3_reg[232][28]/P0001 ,
		_w11982_,
		_w11990_,
		_w12064_
	);
	LUT4 #(
		.INIT('h0001)
	) name1552 (
		_w12061_,
		_w12062_,
		_w12063_,
		_w12064_,
		_w12065_
	);
	LUT4 #(
		.INIT('h8000)
	) name1553 (
		_w12050_,
		_w12055_,
		_w12060_,
		_w12065_,
		_w12066_
	);
	LUT3 #(
		.INIT('h80)
	) name1554 (
		\wishbone_bd_ram_mem3_reg[80][28]/P0001 ,
		_w11941_,
		_w11972_,
		_w12067_
	);
	LUT3 #(
		.INIT('h80)
	) name1555 (
		\wishbone_bd_ram_mem3_reg[235][28]/P0001 ,
		_w11936_,
		_w11982_,
		_w12068_
	);
	LUT3 #(
		.INIT('h80)
	) name1556 (
		\wishbone_bd_ram_mem3_reg[26][28]/P0001 ,
		_w11935_,
		_w11944_,
		_w12069_
	);
	LUT3 #(
		.INIT('h80)
	) name1557 (
		\wishbone_bd_ram_mem3_reg[35][28]/P0001 ,
		_w11938_,
		_w11957_,
		_w12070_
	);
	LUT4 #(
		.INIT('h0001)
	) name1558 (
		_w12067_,
		_w12068_,
		_w12069_,
		_w12070_,
		_w12071_
	);
	LUT3 #(
		.INIT('h80)
	) name1559 (
		\wishbone_bd_ram_mem3_reg[4][28]/P0001 ,
		_w11929_,
		_w11932_,
		_w12072_
	);
	LUT3 #(
		.INIT('h80)
	) name1560 (
		\wishbone_bd_ram_mem3_reg[62][28]/P0001 ,
		_w11948_,
		_w11979_,
		_w12073_
	);
	LUT3 #(
		.INIT('h80)
	) name1561 (
		\wishbone_bd_ram_mem3_reg[18][28]/P0001 ,
		_w11935_,
		_w11963_,
		_w12074_
	);
	LUT3 #(
		.INIT('h80)
	) name1562 (
		\wishbone_bd_ram_mem3_reg[102][28]/P0001 ,
		_w11965_,
		_w11986_,
		_w12075_
	);
	LUT4 #(
		.INIT('h0001)
	) name1563 (
		_w12072_,
		_w12073_,
		_w12074_,
		_w12075_,
		_w12076_
	);
	LUT3 #(
		.INIT('h80)
	) name1564 (
		\wishbone_bd_ram_mem3_reg[0][28]/P0001 ,
		_w11932_,
		_w11941_,
		_w12077_
	);
	LUT3 #(
		.INIT('h80)
	) name1565 (
		\wishbone_bd_ram_mem3_reg[169][28]/P0001 ,
		_w11930_,
		_w11968_,
		_w12078_
	);
	LUT3 #(
		.INIT('h80)
	) name1566 (
		\wishbone_bd_ram_mem3_reg[61][28]/P0001 ,
		_w11966_,
		_w11979_,
		_w12079_
	);
	LUT3 #(
		.INIT('h80)
	) name1567 (
		\wishbone_bd_ram_mem3_reg[7][28]/P0001 ,
		_w11932_,
		_w11975_,
		_w12080_
	);
	LUT4 #(
		.INIT('h0001)
	) name1568 (
		_w12077_,
		_w12078_,
		_w12079_,
		_w12080_,
		_w12081_
	);
	LUT3 #(
		.INIT('h80)
	) name1569 (
		\wishbone_bd_ram_mem3_reg[120][28]/P0001 ,
		_w11990_,
		_w12012_,
		_w12082_
	);
	LUT3 #(
		.INIT('h80)
	) name1570 (
		\wishbone_bd_ram_mem3_reg[229][28]/P0001 ,
		_w11933_,
		_w11982_,
		_w12083_
	);
	LUT3 #(
		.INIT('h80)
	) name1571 (
		\wishbone_bd_ram_mem3_reg[106][28]/P0001 ,
		_w11944_,
		_w11965_,
		_w12084_
	);
	LUT3 #(
		.INIT('h80)
	) name1572 (
		\wishbone_bd_ram_mem3_reg[117][28]/P0001 ,
		_w11933_,
		_w12012_,
		_w12085_
	);
	LUT4 #(
		.INIT('h0001)
	) name1573 (
		_w12082_,
		_w12083_,
		_w12084_,
		_w12085_,
		_w12086_
	);
	LUT4 #(
		.INIT('h8000)
	) name1574 (
		_w12071_,
		_w12076_,
		_w12081_,
		_w12086_,
		_w12087_
	);
	LUT3 #(
		.INIT('h80)
	) name1575 (
		\wishbone_bd_ram_mem3_reg[74][28]/P0001 ,
		_w11944_,
		_w11949_,
		_w12088_
	);
	LUT3 #(
		.INIT('h80)
	) name1576 (
		\wishbone_bd_ram_mem3_reg[139][28]/P0001 ,
		_w11936_,
		_w11955_,
		_w12089_
	);
	LUT3 #(
		.INIT('h80)
	) name1577 (
		\wishbone_bd_ram_mem3_reg[98][28]/P0001 ,
		_w11963_,
		_w11965_,
		_w12090_
	);
	LUT3 #(
		.INIT('h80)
	) name1578 (
		\wishbone_bd_ram_mem3_reg[247][28]/P0001 ,
		_w11952_,
		_w11975_,
		_w12091_
	);
	LUT4 #(
		.INIT('h0001)
	) name1579 (
		_w12088_,
		_w12089_,
		_w12090_,
		_w12091_,
		_w12092_
	);
	LUT3 #(
		.INIT('h80)
	) name1580 (
		\wishbone_bd_ram_mem3_reg[243][28]/P0001 ,
		_w11938_,
		_w11952_,
		_w12093_
	);
	LUT3 #(
		.INIT('h80)
	) name1581 (
		\wishbone_bd_ram_mem3_reg[219][28]/P0001 ,
		_w11936_,
		_w11984_,
		_w12094_
	);
	LUT3 #(
		.INIT('h80)
	) name1582 (
		\wishbone_bd_ram_mem3_reg[9][28]/P0001 ,
		_w11932_,
		_w11968_,
		_w12095_
	);
	LUT3 #(
		.INIT('h80)
	) name1583 (
		\wishbone_bd_ram_mem3_reg[72][28]/P0001 ,
		_w11949_,
		_w11990_,
		_w12096_
	);
	LUT4 #(
		.INIT('h0001)
	) name1584 (
		_w12093_,
		_w12094_,
		_w12095_,
		_w12096_,
		_w12097_
	);
	LUT3 #(
		.INIT('h80)
	) name1585 (
		\wishbone_bd_ram_mem3_reg[181][28]/P0001 ,
		_w11933_,
		_w11942_,
		_w12098_
	);
	LUT3 #(
		.INIT('h80)
	) name1586 (
		\wishbone_bd_ram_mem3_reg[118][28]/P0001 ,
		_w11986_,
		_w12012_,
		_w12099_
	);
	LUT3 #(
		.INIT('h80)
	) name1587 (
		\wishbone_bd_ram_mem3_reg[198][28]/P0001 ,
		_w11945_,
		_w11986_,
		_w12100_
	);
	LUT3 #(
		.INIT('h80)
	) name1588 (
		\wishbone_bd_ram_mem3_reg[197][28]/P0001 ,
		_w11933_,
		_w11945_,
		_w12101_
	);
	LUT4 #(
		.INIT('h0001)
	) name1589 (
		_w12098_,
		_w12099_,
		_w12100_,
		_w12101_,
		_w12102_
	);
	LUT3 #(
		.INIT('h80)
	) name1590 (
		\wishbone_bd_ram_mem3_reg[182][28]/P0001 ,
		_w11942_,
		_w11986_,
		_w12103_
	);
	LUT3 #(
		.INIT('h80)
	) name1591 (
		\wishbone_bd_ram_mem3_reg[201][28]/P0001 ,
		_w11945_,
		_w11968_,
		_w12104_
	);
	LUT3 #(
		.INIT('h80)
	) name1592 (
		\wishbone_bd_ram_mem3_reg[66][28]/P0001 ,
		_w11949_,
		_w11963_,
		_w12105_
	);
	LUT3 #(
		.INIT('h80)
	) name1593 (
		\wishbone_bd_ram_mem3_reg[75][28]/P0001 ,
		_w11936_,
		_w11949_,
		_w12106_
	);
	LUT4 #(
		.INIT('h0001)
	) name1594 (
		_w12103_,
		_w12104_,
		_w12105_,
		_w12106_,
		_w12107_
	);
	LUT4 #(
		.INIT('h8000)
	) name1595 (
		_w12092_,
		_w12097_,
		_w12102_,
		_w12107_,
		_w12108_
	);
	LUT3 #(
		.INIT('h80)
	) name1596 (
		\wishbone_bd_ram_mem3_reg[56][28]/P0001 ,
		_w11979_,
		_w11990_,
		_w12109_
	);
	LUT3 #(
		.INIT('h80)
	) name1597 (
		\wishbone_bd_ram_mem3_reg[59][28]/P0001 ,
		_w11936_,
		_w11979_,
		_w12110_
	);
	LUT3 #(
		.INIT('h80)
	) name1598 (
		\wishbone_bd_ram_mem3_reg[186][28]/P0001 ,
		_w11942_,
		_w11944_,
		_w12111_
	);
	LUT3 #(
		.INIT('h80)
	) name1599 (
		\wishbone_bd_ram_mem3_reg[55][28]/P0001 ,
		_w11975_,
		_w11979_,
		_w12112_
	);
	LUT4 #(
		.INIT('h0001)
	) name1600 (
		_w12109_,
		_w12110_,
		_w12111_,
		_w12112_,
		_w12113_
	);
	LUT3 #(
		.INIT('h80)
	) name1601 (
		\wishbone_bd_ram_mem3_reg[54][28]/P0001 ,
		_w11979_,
		_w11986_,
		_w12114_
	);
	LUT3 #(
		.INIT('h80)
	) name1602 (
		\wishbone_bd_ram_mem3_reg[194][28]/P0001 ,
		_w11945_,
		_w11963_,
		_w12115_
	);
	LUT3 #(
		.INIT('h80)
	) name1603 (
		\wishbone_bd_ram_mem3_reg[159][28]/P0001 ,
		_w11959_,
		_w11973_,
		_w12116_
	);
	LUT3 #(
		.INIT('h80)
	) name1604 (
		\wishbone_bd_ram_mem3_reg[129][28]/P0001 ,
		_w11955_,
		_w11977_,
		_w12117_
	);
	LUT4 #(
		.INIT('h0001)
	) name1605 (
		_w12114_,
		_w12115_,
		_w12116_,
		_w12117_,
		_w12118_
	);
	LUT3 #(
		.INIT('h80)
	) name1606 (
		\wishbone_bd_ram_mem3_reg[212][28]/P0001 ,
		_w11929_,
		_w11984_,
		_w12119_
	);
	LUT3 #(
		.INIT('h80)
	) name1607 (
		\wishbone_bd_ram_mem3_reg[71][28]/P0001 ,
		_w11949_,
		_w11975_,
		_w12120_
	);
	LUT3 #(
		.INIT('h80)
	) name1608 (
		\wishbone_bd_ram_mem3_reg[36][28]/P0001 ,
		_w11929_,
		_w11957_,
		_w12121_
	);
	LUT3 #(
		.INIT('h80)
	) name1609 (
		\wishbone_bd_ram_mem3_reg[221][28]/P0001 ,
		_w11966_,
		_w11984_,
		_w12122_
	);
	LUT4 #(
		.INIT('h0001)
	) name1610 (
		_w12119_,
		_w12120_,
		_w12121_,
		_w12122_,
		_w12123_
	);
	LUT3 #(
		.INIT('h80)
	) name1611 (
		\wishbone_bd_ram_mem3_reg[183][28]/P0001 ,
		_w11942_,
		_w11975_,
		_w12124_
	);
	LUT3 #(
		.INIT('h80)
	) name1612 (
		\wishbone_bd_ram_mem3_reg[248][28]/P0001 ,
		_w11952_,
		_w11990_,
		_w12125_
	);
	LUT3 #(
		.INIT('h80)
	) name1613 (
		\wishbone_bd_ram_mem3_reg[180][28]/P0001 ,
		_w11929_,
		_w11942_,
		_w12126_
	);
	LUT3 #(
		.INIT('h80)
	) name1614 (
		\wishbone_bd_ram_mem3_reg[128][28]/P0001 ,
		_w11941_,
		_w11955_,
		_w12127_
	);
	LUT4 #(
		.INIT('h0001)
	) name1615 (
		_w12124_,
		_w12125_,
		_w12126_,
		_w12127_,
		_w12128_
	);
	LUT4 #(
		.INIT('h8000)
	) name1616 (
		_w12113_,
		_w12118_,
		_w12123_,
		_w12128_,
		_w12129_
	);
	LUT4 #(
		.INIT('h8000)
	) name1617 (
		_w12066_,
		_w12087_,
		_w12108_,
		_w12129_,
		_w12130_
	);
	LUT3 #(
		.INIT('h80)
	) name1618 (
		\wishbone_bd_ram_mem3_reg[40][28]/P0001 ,
		_w11957_,
		_w11990_,
		_w12131_
	);
	LUT3 #(
		.INIT('h80)
	) name1619 (
		\wishbone_bd_ram_mem3_reg[67][28]/P0001 ,
		_w11938_,
		_w11949_,
		_w12132_
	);
	LUT3 #(
		.INIT('h80)
	) name1620 (
		\wishbone_bd_ram_mem3_reg[150][28]/P0001 ,
		_w11959_,
		_w11986_,
		_w12133_
	);
	LUT3 #(
		.INIT('h80)
	) name1621 (
		\wishbone_bd_ram_mem3_reg[226][28]/P0001 ,
		_w11963_,
		_w11982_,
		_w12134_
	);
	LUT4 #(
		.INIT('h0001)
	) name1622 (
		_w12131_,
		_w12132_,
		_w12133_,
		_w12134_,
		_w12135_
	);
	LUT3 #(
		.INIT('h80)
	) name1623 (
		\wishbone_bd_ram_mem3_reg[135][28]/P0001 ,
		_w11955_,
		_w11975_,
		_w12136_
	);
	LUT3 #(
		.INIT('h80)
	) name1624 (
		\wishbone_bd_ram_mem3_reg[175][28]/P0001 ,
		_w11930_,
		_w11973_,
		_w12137_
	);
	LUT3 #(
		.INIT('h80)
	) name1625 (
		\wishbone_bd_ram_mem3_reg[250][28]/P0001 ,
		_w11944_,
		_w11952_,
		_w12138_
	);
	LUT3 #(
		.INIT('h80)
	) name1626 (
		\wishbone_bd_ram_mem3_reg[122][28]/P0001 ,
		_w11944_,
		_w12012_,
		_w12139_
	);
	LUT4 #(
		.INIT('h0001)
	) name1627 (
		_w12136_,
		_w12137_,
		_w12138_,
		_w12139_,
		_w12140_
	);
	LUT3 #(
		.INIT('h80)
	) name1628 (
		\wishbone_bd_ram_mem3_reg[104][28]/P0001 ,
		_w11965_,
		_w11990_,
		_w12141_
	);
	LUT3 #(
		.INIT('h80)
	) name1629 (
		\wishbone_bd_ram_mem3_reg[50][28]/P0001 ,
		_w11963_,
		_w11979_,
		_w12142_
	);
	LUT3 #(
		.INIT('h80)
	) name1630 (
		\wishbone_bd_ram_mem3_reg[209][28]/P0001 ,
		_w11977_,
		_w11984_,
		_w12143_
	);
	LUT3 #(
		.INIT('h80)
	) name1631 (
		\wishbone_bd_ram_mem3_reg[87][28]/P0001 ,
		_w11972_,
		_w11975_,
		_w12144_
	);
	LUT4 #(
		.INIT('h0001)
	) name1632 (
		_w12141_,
		_w12142_,
		_w12143_,
		_w12144_,
		_w12145_
	);
	LUT3 #(
		.INIT('h80)
	) name1633 (
		\wishbone_bd_ram_mem3_reg[16][28]/P0001 ,
		_w11935_,
		_w11941_,
		_w12146_
	);
	LUT3 #(
		.INIT('h80)
	) name1634 (
		\wishbone_bd_ram_mem3_reg[151][28]/P0001 ,
		_w11959_,
		_w11975_,
		_w12147_
	);
	LUT3 #(
		.INIT('h80)
	) name1635 (
		\wishbone_bd_ram_mem3_reg[195][28]/P0001 ,
		_w11938_,
		_w11945_,
		_w12148_
	);
	LUT3 #(
		.INIT('h80)
	) name1636 (
		\wishbone_bd_ram_mem3_reg[147][28]/P0001 ,
		_w11938_,
		_w11959_,
		_w12149_
	);
	LUT4 #(
		.INIT('h0001)
	) name1637 (
		_w12146_,
		_w12147_,
		_w12148_,
		_w12149_,
		_w12150_
	);
	LUT4 #(
		.INIT('h8000)
	) name1638 (
		_w12135_,
		_w12140_,
		_w12145_,
		_w12150_,
		_w12151_
	);
	LUT3 #(
		.INIT('h80)
	) name1639 (
		\wishbone_bd_ram_mem3_reg[253][28]/P0001 ,
		_w11952_,
		_w11966_,
		_w12152_
	);
	LUT3 #(
		.INIT('h80)
	) name1640 (
		\wishbone_bd_ram_mem3_reg[37][28]/P0001 ,
		_w11933_,
		_w11957_,
		_w12153_
	);
	LUT3 #(
		.INIT('h80)
	) name1641 (
		\wishbone_bd_ram_mem3_reg[30][28]/P0001 ,
		_w11935_,
		_w11948_,
		_w12154_
	);
	LUT3 #(
		.INIT('h80)
	) name1642 (
		\wishbone_bd_ram_mem3_reg[145][28]/P0001 ,
		_w11959_,
		_w11977_,
		_w12155_
	);
	LUT4 #(
		.INIT('h0001)
	) name1643 (
		_w12152_,
		_w12153_,
		_w12154_,
		_w12155_,
		_w12156_
	);
	LUT3 #(
		.INIT('h80)
	) name1644 (
		\wishbone_bd_ram_mem3_reg[225][28]/P0001 ,
		_w11977_,
		_w11982_,
		_w12157_
	);
	LUT3 #(
		.INIT('h80)
	) name1645 (
		\wishbone_bd_ram_mem3_reg[222][28]/P0001 ,
		_w11948_,
		_w11984_,
		_w12158_
	);
	LUT3 #(
		.INIT('h80)
	) name1646 (
		\wishbone_bd_ram_mem3_reg[97][28]/P0001 ,
		_w11965_,
		_w11977_,
		_w12159_
	);
	LUT3 #(
		.INIT('h80)
	) name1647 (
		\wishbone_bd_ram_mem3_reg[162][28]/P0001 ,
		_w11930_,
		_w11963_,
		_w12160_
	);
	LUT4 #(
		.INIT('h0001)
	) name1648 (
		_w12157_,
		_w12158_,
		_w12159_,
		_w12160_,
		_w12161_
	);
	LUT3 #(
		.INIT('h80)
	) name1649 (
		\wishbone_bd_ram_mem3_reg[57][28]/P0001 ,
		_w11968_,
		_w11979_,
		_w12162_
	);
	LUT3 #(
		.INIT('h80)
	) name1650 (
		\wishbone_bd_ram_mem3_reg[12][28]/P0001 ,
		_w11932_,
		_w11954_,
		_w12163_
	);
	LUT3 #(
		.INIT('h80)
	) name1651 (
		\wishbone_bd_ram_mem3_reg[32][28]/P0001 ,
		_w11941_,
		_w11957_,
		_w12164_
	);
	LUT3 #(
		.INIT('h80)
	) name1652 (
		\wishbone_bd_ram_mem3_reg[155][28]/P0001 ,
		_w11936_,
		_w11959_,
		_w12165_
	);
	LUT4 #(
		.INIT('h0001)
	) name1653 (
		_w12162_,
		_w12163_,
		_w12164_,
		_w12165_,
		_w12166_
	);
	LUT3 #(
		.INIT('h80)
	) name1654 (
		\wishbone_bd_ram_mem3_reg[25][28]/P0001 ,
		_w11935_,
		_w11968_,
		_w12167_
	);
	LUT3 #(
		.INIT('h80)
	) name1655 (
		\wishbone_bd_ram_mem3_reg[22][28]/P0001 ,
		_w11935_,
		_w11986_,
		_w12168_
	);
	LUT3 #(
		.INIT('h80)
	) name1656 (
		\wishbone_bd_ram_mem3_reg[115][28]/P0001 ,
		_w11938_,
		_w12012_,
		_w12169_
	);
	LUT3 #(
		.INIT('h80)
	) name1657 (
		\wishbone_bd_ram_mem3_reg[123][28]/P0001 ,
		_w11936_,
		_w12012_,
		_w12170_
	);
	LUT4 #(
		.INIT('h0001)
	) name1658 (
		_w12167_,
		_w12168_,
		_w12169_,
		_w12170_,
		_w12171_
	);
	LUT4 #(
		.INIT('h8000)
	) name1659 (
		_w12156_,
		_w12161_,
		_w12166_,
		_w12171_,
		_w12172_
	);
	LUT3 #(
		.INIT('h80)
	) name1660 (
		\wishbone_bd_ram_mem3_reg[187][28]/P0001 ,
		_w11936_,
		_w11942_,
		_w12173_
	);
	LUT3 #(
		.INIT('h80)
	) name1661 (
		\wishbone_bd_ram_mem3_reg[31][28]/P0001 ,
		_w11935_,
		_w11973_,
		_w12174_
	);
	LUT3 #(
		.INIT('h80)
	) name1662 (
		\wishbone_bd_ram_mem3_reg[43][28]/P0001 ,
		_w11936_,
		_w11957_,
		_w12175_
	);
	LUT3 #(
		.INIT('h80)
	) name1663 (
		\wishbone_bd_ram_mem3_reg[114][28]/P0001 ,
		_w11963_,
		_w12012_,
		_w12176_
	);
	LUT4 #(
		.INIT('h0001)
	) name1664 (
		_w12173_,
		_w12174_,
		_w12175_,
		_w12176_,
		_w12177_
	);
	LUT3 #(
		.INIT('h80)
	) name1665 (
		\wishbone_bd_ram_mem3_reg[217][28]/P0001 ,
		_w11968_,
		_w11984_,
		_w12178_
	);
	LUT3 #(
		.INIT('h80)
	) name1666 (
		\wishbone_bd_ram_mem3_reg[156][28]/P0001 ,
		_w11954_,
		_w11959_,
		_w12179_
	);
	LUT3 #(
		.INIT('h80)
	) name1667 (
		\wishbone_bd_ram_mem3_reg[101][28]/P0001 ,
		_w11933_,
		_w11965_,
		_w12180_
	);
	LUT3 #(
		.INIT('h80)
	) name1668 (
		\wishbone_bd_ram_mem3_reg[11][28]/P0001 ,
		_w11932_,
		_w11936_,
		_w12181_
	);
	LUT4 #(
		.INIT('h0001)
	) name1669 (
		_w12178_,
		_w12179_,
		_w12180_,
		_w12181_,
		_w12182_
	);
	LUT3 #(
		.INIT('h80)
	) name1670 (
		\wishbone_bd_ram_mem3_reg[79][28]/P0001 ,
		_w11949_,
		_w11973_,
		_w12183_
	);
	LUT3 #(
		.INIT('h80)
	) name1671 (
		\wishbone_bd_ram_mem3_reg[234][28]/P0001 ,
		_w11944_,
		_w11982_,
		_w12184_
	);
	LUT3 #(
		.INIT('h80)
	) name1672 (
		\wishbone_bd_ram_mem3_reg[85][28]/P0001 ,
		_w11933_,
		_w11972_,
		_w12185_
	);
	LUT3 #(
		.INIT('h80)
	) name1673 (
		\wishbone_bd_ram_mem3_reg[126][28]/P0001 ,
		_w11948_,
		_w12012_,
		_w12186_
	);
	LUT4 #(
		.INIT('h0001)
	) name1674 (
		_w12183_,
		_w12184_,
		_w12185_,
		_w12186_,
		_w12187_
	);
	LUT3 #(
		.INIT('h80)
	) name1675 (
		\wishbone_bd_ram_mem3_reg[60][28]/P0001 ,
		_w11954_,
		_w11979_,
		_w12188_
	);
	LUT3 #(
		.INIT('h80)
	) name1676 (
		\wishbone_bd_ram_mem3_reg[218][28]/P0001 ,
		_w11944_,
		_w11984_,
		_w12189_
	);
	LUT3 #(
		.INIT('h80)
	) name1677 (
		\wishbone_bd_ram_mem3_reg[168][28]/P0001 ,
		_w11930_,
		_w11990_,
		_w12190_
	);
	LUT3 #(
		.INIT('h80)
	) name1678 (
		\wishbone_bd_ram_mem3_reg[15][28]/P0001 ,
		_w11932_,
		_w11973_,
		_w12191_
	);
	LUT4 #(
		.INIT('h0001)
	) name1679 (
		_w12188_,
		_w12189_,
		_w12190_,
		_w12191_,
		_w12192_
	);
	LUT4 #(
		.INIT('h8000)
	) name1680 (
		_w12177_,
		_w12182_,
		_w12187_,
		_w12192_,
		_w12193_
	);
	LUT3 #(
		.INIT('h80)
	) name1681 (
		\wishbone_bd_ram_mem3_reg[127][28]/P0001 ,
		_w11973_,
		_w12012_,
		_w12194_
	);
	LUT3 #(
		.INIT('h80)
	) name1682 (
		\wishbone_bd_ram_mem3_reg[211][28]/P0001 ,
		_w11938_,
		_w11984_,
		_w12195_
	);
	LUT3 #(
		.INIT('h80)
	) name1683 (
		\wishbone_bd_ram_mem3_reg[137][28]/P0001 ,
		_w11955_,
		_w11968_,
		_w12196_
	);
	LUT3 #(
		.INIT('h80)
	) name1684 (
		\wishbone_bd_ram_mem3_reg[28][28]/P0001 ,
		_w11935_,
		_w11954_,
		_w12197_
	);
	LUT4 #(
		.INIT('h0001)
	) name1685 (
		_w12194_,
		_w12195_,
		_w12196_,
		_w12197_,
		_w12198_
	);
	LUT3 #(
		.INIT('h80)
	) name1686 (
		\wishbone_bd_ram_mem3_reg[108][28]/P0001 ,
		_w11954_,
		_w11965_,
		_w12199_
	);
	LUT3 #(
		.INIT('h80)
	) name1687 (
		\wishbone_bd_ram_mem3_reg[203][28]/P0001 ,
		_w11936_,
		_w11945_,
		_w12200_
	);
	LUT3 #(
		.INIT('h80)
	) name1688 (
		\wishbone_bd_ram_mem3_reg[238][28]/P0001 ,
		_w11948_,
		_w11982_,
		_w12201_
	);
	LUT3 #(
		.INIT('h80)
	) name1689 (
		\wishbone_bd_ram_mem3_reg[204][28]/P0001 ,
		_w11945_,
		_w11954_,
		_w12202_
	);
	LUT4 #(
		.INIT('h0001)
	) name1690 (
		_w12199_,
		_w12200_,
		_w12201_,
		_w12202_,
		_w12203_
	);
	LUT3 #(
		.INIT('h80)
	) name1691 (
		\wishbone_bd_ram_mem3_reg[207][28]/P0001 ,
		_w11945_,
		_w11973_,
		_w12204_
	);
	LUT3 #(
		.INIT('h80)
	) name1692 (
		\wishbone_bd_ram_mem3_reg[38][28]/P0001 ,
		_w11957_,
		_w11986_,
		_w12205_
	);
	LUT3 #(
		.INIT('h80)
	) name1693 (
		\wishbone_bd_ram_mem3_reg[76][28]/P0001 ,
		_w11949_,
		_w11954_,
		_w12206_
	);
	LUT3 #(
		.INIT('h80)
	) name1694 (
		\wishbone_bd_ram_mem3_reg[94][28]/P0001 ,
		_w11948_,
		_w11972_,
		_w12207_
	);
	LUT4 #(
		.INIT('h0001)
	) name1695 (
		_w12204_,
		_w12205_,
		_w12206_,
		_w12207_,
		_w12208_
	);
	LUT3 #(
		.INIT('h80)
	) name1696 (
		\wishbone_bd_ram_mem3_reg[10][28]/P0001 ,
		_w11932_,
		_w11944_,
		_w12209_
	);
	LUT3 #(
		.INIT('h80)
	) name1697 (
		\wishbone_bd_ram_mem3_reg[20][28]/P0001 ,
		_w11929_,
		_w11935_,
		_w12210_
	);
	LUT3 #(
		.INIT('h80)
	) name1698 (
		\wishbone_bd_ram_mem3_reg[65][28]/P0001 ,
		_w11949_,
		_w11977_,
		_w12211_
	);
	LUT3 #(
		.INIT('h80)
	) name1699 (
		\wishbone_bd_ram_mem3_reg[13][28]/P0001 ,
		_w11932_,
		_w11966_,
		_w12212_
	);
	LUT4 #(
		.INIT('h0001)
	) name1700 (
		_w12209_,
		_w12210_,
		_w12211_,
		_w12212_,
		_w12213_
	);
	LUT4 #(
		.INIT('h8000)
	) name1701 (
		_w12198_,
		_w12203_,
		_w12208_,
		_w12213_,
		_w12214_
	);
	LUT4 #(
		.INIT('h8000)
	) name1702 (
		_w12151_,
		_w12172_,
		_w12193_,
		_w12214_,
		_w12215_
	);
	LUT3 #(
		.INIT('h80)
	) name1703 (
		\wishbone_bd_ram_mem3_reg[141][28]/P0001 ,
		_w11955_,
		_w11966_,
		_w12216_
	);
	LUT3 #(
		.INIT('h80)
	) name1704 (
		\wishbone_bd_ram_mem3_reg[241][28]/P0001 ,
		_w11952_,
		_w11977_,
		_w12217_
	);
	LUT3 #(
		.INIT('h80)
	) name1705 (
		\wishbone_bd_ram_mem3_reg[23][28]/P0001 ,
		_w11935_,
		_w11975_,
		_w12218_
	);
	LUT3 #(
		.INIT('h80)
	) name1706 (
		\wishbone_bd_ram_mem3_reg[92][28]/P0001 ,
		_w11954_,
		_w11972_,
		_w12219_
	);
	LUT4 #(
		.INIT('h0001)
	) name1707 (
		_w12216_,
		_w12217_,
		_w12218_,
		_w12219_,
		_w12220_
	);
	LUT3 #(
		.INIT('h80)
	) name1708 (
		\wishbone_bd_ram_mem3_reg[177][28]/P0001 ,
		_w11942_,
		_w11977_,
		_w12221_
	);
	LUT3 #(
		.INIT('h80)
	) name1709 (
		\wishbone_bd_ram_mem3_reg[116][28]/P0001 ,
		_w11929_,
		_w12012_,
		_w12222_
	);
	LUT3 #(
		.INIT('h80)
	) name1710 (
		\wishbone_bd_ram_mem3_reg[148][28]/P0001 ,
		_w11929_,
		_w11959_,
		_w12223_
	);
	LUT3 #(
		.INIT('h80)
	) name1711 (
		\wishbone_bd_ram_mem3_reg[213][28]/P0001 ,
		_w11933_,
		_w11984_,
		_w12224_
	);
	LUT4 #(
		.INIT('h0001)
	) name1712 (
		_w12221_,
		_w12222_,
		_w12223_,
		_w12224_,
		_w12225_
	);
	LUT3 #(
		.INIT('h80)
	) name1713 (
		\wishbone_bd_ram_mem3_reg[53][28]/P0001 ,
		_w11933_,
		_w11979_,
		_w12226_
	);
	LUT3 #(
		.INIT('h80)
	) name1714 (
		\wishbone_bd_ram_mem3_reg[245][28]/P0001 ,
		_w11933_,
		_w11952_,
		_w12227_
	);
	LUT3 #(
		.INIT('h80)
	) name1715 (
		\wishbone_bd_ram_mem3_reg[51][28]/P0001 ,
		_w11938_,
		_w11979_,
		_w12228_
	);
	LUT3 #(
		.INIT('h80)
	) name1716 (
		\wishbone_bd_ram_mem3_reg[113][28]/P0001 ,
		_w11977_,
		_w12012_,
		_w12229_
	);
	LUT4 #(
		.INIT('h0001)
	) name1717 (
		_w12226_,
		_w12227_,
		_w12228_,
		_w12229_,
		_w12230_
	);
	LUT3 #(
		.INIT('h80)
	) name1718 (
		\wishbone_bd_ram_mem3_reg[19][28]/P0001 ,
		_w11935_,
		_w11938_,
		_w12231_
	);
	LUT3 #(
		.INIT('h80)
	) name1719 (
		\wishbone_bd_ram_mem3_reg[1][28]/P0001 ,
		_w11932_,
		_w11977_,
		_w12232_
	);
	LUT3 #(
		.INIT('h80)
	) name1720 (
		\wishbone_bd_ram_mem3_reg[93][28]/P0001 ,
		_w11966_,
		_w11972_,
		_w12233_
	);
	LUT3 #(
		.INIT('h80)
	) name1721 (
		\wishbone_bd_ram_mem3_reg[39][28]/P0001 ,
		_w11957_,
		_w11975_,
		_w12234_
	);
	LUT4 #(
		.INIT('h0001)
	) name1722 (
		_w12231_,
		_w12232_,
		_w12233_,
		_w12234_,
		_w12235_
	);
	LUT4 #(
		.INIT('h8000)
	) name1723 (
		_w12220_,
		_w12225_,
		_w12230_,
		_w12235_,
		_w12236_
	);
	LUT3 #(
		.INIT('h80)
	) name1724 (
		\wishbone_bd_ram_mem3_reg[174][28]/P0001 ,
		_w11930_,
		_w11948_,
		_w12237_
	);
	LUT3 #(
		.INIT('h80)
	) name1725 (
		\wishbone_bd_ram_mem3_reg[215][28]/P0001 ,
		_w11975_,
		_w11984_,
		_w12238_
	);
	LUT3 #(
		.INIT('h80)
	) name1726 (
		\wishbone_bd_ram_mem3_reg[64][28]/P0001 ,
		_w11941_,
		_w11949_,
		_w12239_
	);
	LUT3 #(
		.INIT('h80)
	) name1727 (
		\wishbone_bd_ram_mem3_reg[90][28]/P0001 ,
		_w11944_,
		_w11972_,
		_w12240_
	);
	LUT4 #(
		.INIT('h0001)
	) name1728 (
		_w12237_,
		_w12238_,
		_w12239_,
		_w12240_,
		_w12241_
	);
	LUT3 #(
		.INIT('h80)
	) name1729 (
		\wishbone_bd_ram_mem3_reg[89][28]/P0001 ,
		_w11968_,
		_w11972_,
		_w12242_
	);
	LUT3 #(
		.INIT('h80)
	) name1730 (
		\wishbone_bd_ram_mem3_reg[152][28]/P0001 ,
		_w11959_,
		_w11990_,
		_w12243_
	);
	LUT3 #(
		.INIT('h80)
	) name1731 (
		\wishbone_bd_ram_mem3_reg[6][28]/P0001 ,
		_w11932_,
		_w11986_,
		_w12244_
	);
	LUT3 #(
		.INIT('h80)
	) name1732 (
		\wishbone_bd_ram_mem3_reg[48][28]/P0001 ,
		_w11941_,
		_w11979_,
		_w12245_
	);
	LUT4 #(
		.INIT('h0001)
	) name1733 (
		_w12242_,
		_w12243_,
		_w12244_,
		_w12245_,
		_w12246_
	);
	LUT3 #(
		.INIT('h80)
	) name1734 (
		\wishbone_bd_ram_mem3_reg[200][28]/P0001 ,
		_w11945_,
		_w11990_,
		_w12247_
	);
	LUT3 #(
		.INIT('h80)
	) name1735 (
		\wishbone_bd_ram_mem3_reg[237][28]/P0001 ,
		_w11966_,
		_w11982_,
		_w12248_
	);
	LUT3 #(
		.INIT('h80)
	) name1736 (
		\wishbone_bd_ram_mem3_reg[132][28]/P0001 ,
		_w11929_,
		_w11955_,
		_w12249_
	);
	LUT3 #(
		.INIT('h80)
	) name1737 (
		\wishbone_bd_ram_mem3_reg[49][28]/P0001 ,
		_w11977_,
		_w11979_,
		_w12250_
	);
	LUT4 #(
		.INIT('h0001)
	) name1738 (
		_w12247_,
		_w12248_,
		_w12249_,
		_w12250_,
		_w12251_
	);
	LUT3 #(
		.INIT('h80)
	) name1739 (
		\wishbone_bd_ram_mem3_reg[33][28]/P0001 ,
		_w11957_,
		_w11977_,
		_w12252_
	);
	LUT3 #(
		.INIT('h80)
	) name1740 (
		\wishbone_bd_ram_mem3_reg[77][28]/P0001 ,
		_w11949_,
		_w11966_,
		_w12253_
	);
	LUT3 #(
		.INIT('h80)
	) name1741 (
		\wishbone_bd_ram_mem3_reg[214][28]/P0001 ,
		_w11984_,
		_w11986_,
		_w12254_
	);
	LUT3 #(
		.INIT('h80)
	) name1742 (
		\wishbone_bd_ram_mem3_reg[167][28]/P0001 ,
		_w11930_,
		_w11975_,
		_w12255_
	);
	LUT4 #(
		.INIT('h0001)
	) name1743 (
		_w12252_,
		_w12253_,
		_w12254_,
		_w12255_,
		_w12256_
	);
	LUT4 #(
		.INIT('h8000)
	) name1744 (
		_w12241_,
		_w12246_,
		_w12251_,
		_w12256_,
		_w12257_
	);
	LUT3 #(
		.INIT('h80)
	) name1745 (
		\wishbone_bd_ram_mem3_reg[205][28]/P0001 ,
		_w11945_,
		_w11966_,
		_w12258_
	);
	LUT3 #(
		.INIT('h80)
	) name1746 (
		\wishbone_bd_ram_mem3_reg[58][28]/P0001 ,
		_w11944_,
		_w11979_,
		_w12259_
	);
	LUT3 #(
		.INIT('h80)
	) name1747 (
		\wishbone_bd_ram_mem3_reg[255][28]/P0001 ,
		_w11952_,
		_w11973_,
		_w12260_
	);
	LUT3 #(
		.INIT('h80)
	) name1748 (
		\wishbone_bd_ram_mem3_reg[91][28]/P0001 ,
		_w11936_,
		_w11972_,
		_w12261_
	);
	LUT4 #(
		.INIT('h0001)
	) name1749 (
		_w12258_,
		_w12259_,
		_w12260_,
		_w12261_,
		_w12262_
	);
	LUT3 #(
		.INIT('h80)
	) name1750 (
		\wishbone_bd_ram_mem3_reg[146][28]/P0001 ,
		_w11959_,
		_w11963_,
		_w12263_
	);
	LUT3 #(
		.INIT('h80)
	) name1751 (
		\wishbone_bd_ram_mem3_reg[184][28]/P0001 ,
		_w11942_,
		_w11990_,
		_w12264_
	);
	LUT3 #(
		.INIT('h80)
	) name1752 (
		\wishbone_bd_ram_mem3_reg[136][28]/P0001 ,
		_w11955_,
		_w11990_,
		_w12265_
	);
	LUT3 #(
		.INIT('h80)
	) name1753 (
		\wishbone_bd_ram_mem3_reg[220][28]/P0001 ,
		_w11954_,
		_w11984_,
		_w12266_
	);
	LUT4 #(
		.INIT('h0001)
	) name1754 (
		_w12263_,
		_w12264_,
		_w12265_,
		_w12266_,
		_w12267_
	);
	LUT3 #(
		.INIT('h80)
	) name1755 (
		\wishbone_bd_ram_mem3_reg[24][28]/P0001 ,
		_w11935_,
		_w11990_,
		_w12268_
	);
	LUT3 #(
		.INIT('h80)
	) name1756 (
		\wishbone_bd_ram_mem3_reg[14][28]/P0001 ,
		_w11932_,
		_w11948_,
		_w12269_
	);
	LUT3 #(
		.INIT('h80)
	) name1757 (
		\wishbone_bd_ram_mem3_reg[2][28]/P0001 ,
		_w11932_,
		_w11963_,
		_w12270_
	);
	LUT3 #(
		.INIT('h80)
	) name1758 (
		\wishbone_bd_ram_mem3_reg[196][28]/P0001 ,
		_w11929_,
		_w11945_,
		_w12271_
	);
	LUT4 #(
		.INIT('h0001)
	) name1759 (
		_w12268_,
		_w12269_,
		_w12270_,
		_w12271_,
		_w12272_
	);
	LUT3 #(
		.INIT('h80)
	) name1760 (
		\wishbone_bd_ram_mem3_reg[246][28]/P0001 ,
		_w11952_,
		_w11986_,
		_w12273_
	);
	LUT3 #(
		.INIT('h80)
	) name1761 (
		\wishbone_bd_ram_mem3_reg[121][28]/P0001 ,
		_w11968_,
		_w12012_,
		_w12274_
	);
	LUT3 #(
		.INIT('h80)
	) name1762 (
		\wishbone_bd_ram_mem3_reg[252][28]/P0001 ,
		_w11952_,
		_w11954_,
		_w12275_
	);
	LUT3 #(
		.INIT('h80)
	) name1763 (
		\wishbone_bd_ram_mem3_reg[52][28]/P0001 ,
		_w11929_,
		_w11979_,
		_w12276_
	);
	LUT4 #(
		.INIT('h0001)
	) name1764 (
		_w12273_,
		_w12274_,
		_w12275_,
		_w12276_,
		_w12277_
	);
	LUT4 #(
		.INIT('h8000)
	) name1765 (
		_w12262_,
		_w12267_,
		_w12272_,
		_w12277_,
		_w12278_
	);
	LUT3 #(
		.INIT('h80)
	) name1766 (
		\wishbone_bd_ram_mem3_reg[230][28]/P0001 ,
		_w11982_,
		_w11986_,
		_w12279_
	);
	LUT3 #(
		.INIT('h80)
	) name1767 (
		\wishbone_bd_ram_mem3_reg[99][28]/P0001 ,
		_w11938_,
		_w11965_,
		_w12280_
	);
	LUT3 #(
		.INIT('h80)
	) name1768 (
		\wishbone_bd_ram_mem3_reg[166][28]/P0001 ,
		_w11930_,
		_w11986_,
		_w12281_
	);
	LUT3 #(
		.INIT('h80)
	) name1769 (
		\wishbone_bd_ram_mem3_reg[189][28]/P0001 ,
		_w11942_,
		_w11966_,
		_w12282_
	);
	LUT4 #(
		.INIT('h0001)
	) name1770 (
		_w12279_,
		_w12280_,
		_w12281_,
		_w12282_,
		_w12283_
	);
	LUT3 #(
		.INIT('h80)
	) name1771 (
		\wishbone_bd_ram_mem3_reg[216][28]/P0001 ,
		_w11984_,
		_w11990_,
		_w12284_
	);
	LUT3 #(
		.INIT('h80)
	) name1772 (
		\wishbone_bd_ram_mem3_reg[170][28]/P0001 ,
		_w11930_,
		_w11944_,
		_w12285_
	);
	LUT3 #(
		.INIT('h80)
	) name1773 (
		\wishbone_bd_ram_mem3_reg[208][28]/P0001 ,
		_w11941_,
		_w11984_,
		_w12286_
	);
	LUT3 #(
		.INIT('h80)
	) name1774 (
		\wishbone_bd_ram_mem3_reg[191][28]/P0001 ,
		_w11942_,
		_w11973_,
		_w12287_
	);
	LUT4 #(
		.INIT('h0001)
	) name1775 (
		_w12284_,
		_w12285_,
		_w12286_,
		_w12287_,
		_w12288_
	);
	LUT3 #(
		.INIT('h80)
	) name1776 (
		\wishbone_bd_ram_mem3_reg[41][28]/P0001 ,
		_w11957_,
		_w11968_,
		_w12289_
	);
	LUT3 #(
		.INIT('h80)
	) name1777 (
		\wishbone_bd_ram_mem3_reg[251][28]/P0001 ,
		_w11936_,
		_w11952_,
		_w12290_
	);
	LUT3 #(
		.INIT('h80)
	) name1778 (
		\wishbone_bd_ram_mem3_reg[193][28]/P0001 ,
		_w11945_,
		_w11977_,
		_w12291_
	);
	LUT3 #(
		.INIT('h80)
	) name1779 (
		\wishbone_bd_ram_mem3_reg[124][28]/P0001 ,
		_w11954_,
		_w12012_,
		_w12292_
	);
	LUT4 #(
		.INIT('h0001)
	) name1780 (
		_w12289_,
		_w12290_,
		_w12291_,
		_w12292_,
		_w12293_
	);
	LUT3 #(
		.INIT('h80)
	) name1781 (
		\wishbone_bd_ram_mem3_reg[165][28]/P0001 ,
		_w11930_,
		_w11933_,
		_w12294_
	);
	LUT3 #(
		.INIT('h80)
	) name1782 (
		\wishbone_bd_ram_mem3_reg[110][28]/P0001 ,
		_w11948_,
		_w11965_,
		_w12295_
	);
	LUT3 #(
		.INIT('h80)
	) name1783 (
		\wishbone_bd_ram_mem3_reg[119][28]/P0001 ,
		_w11975_,
		_w12012_,
		_w12296_
	);
	LUT3 #(
		.INIT('h80)
	) name1784 (
		\wishbone_bd_ram_mem3_reg[179][28]/P0001 ,
		_w11938_,
		_w11942_,
		_w12297_
	);
	LUT4 #(
		.INIT('h0001)
	) name1785 (
		_w12294_,
		_w12295_,
		_w12296_,
		_w12297_,
		_w12298_
	);
	LUT4 #(
		.INIT('h8000)
	) name1786 (
		_w12283_,
		_w12288_,
		_w12293_,
		_w12298_,
		_w12299_
	);
	LUT4 #(
		.INIT('h8000)
	) name1787 (
		_w12236_,
		_w12257_,
		_w12278_,
		_w12299_,
		_w12300_
	);
	LUT4 #(
		.INIT('h8000)
	) name1788 (
		_w12045_,
		_w12130_,
		_w12215_,
		_w12300_,
		_w12301_
	);
	LUT3 #(
		.INIT('h80)
	) name1789 (
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w12302_
	);
	LUT4 #(
		.INIT('h4000)
	) name1790 (
		wb_rst_i_pad,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w12303_
	);
	LUT2 #(
		.INIT('h8)
	) name1791 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		_w12304_
	);
	LUT3 #(
		.INIT('h70)
	) name1792 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_TxLength_reg[12]/NET0131 ,
		_w12305_
	);
	LUT2 #(
		.INIT('h4)
	) name1793 (
		_w12302_,
		_w12305_,
		_w12306_
	);
	LUT3 #(
		.INIT('h01)
	) name1794 (
		\wishbone_TxLength_reg[7]/NET0131 ,
		\wishbone_TxLength_reg[8]/NET0131 ,
		\wishbone_TxLength_reg[9]/NET0131 ,
		_w12307_
	);
	LUT2 #(
		.INIT('h1)
	) name1795 (
		\wishbone_TxLength_reg[2]/NET0131 ,
		\wishbone_TxLength_reg[3]/NET0131 ,
		_w12308_
	);
	LUT3 #(
		.INIT('h01)
	) name1796 (
		\wishbone_TxLength_reg[2]/NET0131 ,
		\wishbone_TxLength_reg[3]/NET0131 ,
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w12309_
	);
	LUT2 #(
		.INIT('h1)
	) name1797 (
		\wishbone_TxLength_reg[5]/NET0131 ,
		\wishbone_TxLength_reg[6]/NET0131 ,
		_w12310_
	);
	LUT2 #(
		.INIT('h8)
	) name1798 (
		_w12309_,
		_w12310_,
		_w12311_
	);
	LUT3 #(
		.INIT('h80)
	) name1799 (
		_w12307_,
		_w12309_,
		_w12310_,
		_w12312_
	);
	LUT2 #(
		.INIT('h1)
	) name1800 (
		\wishbone_TxLength_reg[10]/NET0131 ,
		\wishbone_TxLength_reg[11]/NET0131 ,
		_w12313_
	);
	LUT3 #(
		.INIT('h01)
	) name1801 (
		\wishbone_TxLength_reg[10]/NET0131 ,
		\wishbone_TxLength_reg[11]/NET0131 ,
		\wishbone_TxLength_reg[14]/NET0131 ,
		_w12314_
	);
	LUT2 #(
		.INIT('h1)
	) name1802 (
		\wishbone_TxLength_reg[12]/NET0131 ,
		\wishbone_TxLength_reg[13]/NET0131 ,
		_w12315_
	);
	LUT3 #(
		.INIT('h01)
	) name1803 (
		\wishbone_TxLength_reg[12]/NET0131 ,
		\wishbone_TxLength_reg[13]/NET0131 ,
		\wishbone_TxLength_reg[15]/NET0131 ,
		_w12316_
	);
	LUT2 #(
		.INIT('h8)
	) name1804 (
		_w12314_,
		_w12316_,
		_w12317_
	);
	LUT2 #(
		.INIT('h4)
	) name1805 (
		_w12302_,
		_w12304_,
		_w12318_
	);
	LUT3 #(
		.INIT('h70)
	) name1806 (
		_w12312_,
		_w12317_,
		_w12318_,
		_w12319_
	);
	LUT4 #(
		.INIT('h4055)
	) name1807 (
		_w12306_,
		_w12312_,
		_w12317_,
		_w12318_,
		_w12320_
	);
	LUT2 #(
		.INIT('h8)
	) name1808 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		_w12321_
	);
	LUT3 #(
		.INIT('h80)
	) name1809 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		_w12322_
	);
	LUT4 #(
		.INIT('hec80)
	) name1810 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w12323_
	);
	LUT4 #(
		.INIT('h8000)
	) name1811 (
		_w12307_,
		_w12309_,
		_w12310_,
		_w12313_,
		_w12324_
	);
	LUT4 #(
		.INIT('hedee)
	) name1812 (
		\wishbone_TxLength_reg[12]/NET0131 ,
		_w12306_,
		_w12323_,
		_w12324_,
		_w12325_
	);
	LUT2 #(
		.INIT('h4)
	) name1813 (
		_w12320_,
		_w12325_,
		_w12326_
	);
	LUT3 #(
		.INIT('hf4)
	) name1814 (
		_w12301_,
		_w12303_,
		_w12326_,
		_w12327_
	);
	LUT3 #(
		.INIT('h80)
	) name1815 (
		\wishbone_bd_ram_mem3_reg[77][29]/P0001 ,
		_w11949_,
		_w11966_,
		_w12328_
	);
	LUT3 #(
		.INIT('h80)
	) name1816 (
		\wishbone_bd_ram_mem3_reg[42][29]/P0001 ,
		_w11944_,
		_w11957_,
		_w12329_
	);
	LUT3 #(
		.INIT('h80)
	) name1817 (
		\wishbone_bd_ram_mem3_reg[65][29]/P0001 ,
		_w11949_,
		_w11977_,
		_w12330_
	);
	LUT3 #(
		.INIT('h80)
	) name1818 (
		\wishbone_bd_ram_mem3_reg[70][29]/P0001 ,
		_w11949_,
		_w11986_,
		_w12331_
	);
	LUT4 #(
		.INIT('h0001)
	) name1819 (
		_w12328_,
		_w12329_,
		_w12330_,
		_w12331_,
		_w12332_
	);
	LUT3 #(
		.INIT('h80)
	) name1820 (
		\wishbone_bd_ram_mem3_reg[202][29]/P0001 ,
		_w11944_,
		_w11945_,
		_w12333_
	);
	LUT3 #(
		.INIT('h80)
	) name1821 (
		\wishbone_bd_ram_mem3_reg[111][29]/P0001 ,
		_w11965_,
		_w11973_,
		_w12334_
	);
	LUT3 #(
		.INIT('h80)
	) name1822 (
		\wishbone_bd_ram_mem3_reg[160][29]/P0001 ,
		_w11930_,
		_w11941_,
		_w12335_
	);
	LUT3 #(
		.INIT('h80)
	) name1823 (
		\wishbone_bd_ram_mem3_reg[127][29]/P0001 ,
		_w11973_,
		_w12012_,
		_w12336_
	);
	LUT4 #(
		.INIT('h0001)
	) name1824 (
		_w12333_,
		_w12334_,
		_w12335_,
		_w12336_,
		_w12337_
	);
	LUT3 #(
		.INIT('h80)
	) name1825 (
		\wishbone_bd_ram_mem3_reg[71][29]/P0001 ,
		_w11949_,
		_w11975_,
		_w12338_
	);
	LUT3 #(
		.INIT('h80)
	) name1826 (
		\wishbone_bd_ram_mem3_reg[113][29]/P0001 ,
		_w11977_,
		_w12012_,
		_w12339_
	);
	LUT3 #(
		.INIT('h80)
	) name1827 (
		\wishbone_bd_ram_mem3_reg[86][29]/P0001 ,
		_w11972_,
		_w11986_,
		_w12340_
	);
	LUT3 #(
		.INIT('h80)
	) name1828 (
		\wishbone_bd_ram_mem3_reg[158][29]/P0001 ,
		_w11948_,
		_w11959_,
		_w12341_
	);
	LUT4 #(
		.INIT('h0001)
	) name1829 (
		_w12338_,
		_w12339_,
		_w12340_,
		_w12341_,
		_w12342_
	);
	LUT3 #(
		.INIT('h80)
	) name1830 (
		\wishbone_bd_ram_mem3_reg[46][29]/P0001 ,
		_w11948_,
		_w11957_,
		_w12343_
	);
	LUT3 #(
		.INIT('h80)
	) name1831 (
		\wishbone_bd_ram_mem3_reg[112][29]/P0001 ,
		_w11941_,
		_w12012_,
		_w12344_
	);
	LUT3 #(
		.INIT('h80)
	) name1832 (
		\wishbone_bd_ram_mem3_reg[36][29]/P0001 ,
		_w11929_,
		_w11957_,
		_w12345_
	);
	LUT3 #(
		.INIT('h80)
	) name1833 (
		\wishbone_bd_ram_mem3_reg[90][29]/P0001 ,
		_w11944_,
		_w11972_,
		_w12346_
	);
	LUT4 #(
		.INIT('h0001)
	) name1834 (
		_w12343_,
		_w12344_,
		_w12345_,
		_w12346_,
		_w12347_
	);
	LUT4 #(
		.INIT('h8000)
	) name1835 (
		_w12332_,
		_w12337_,
		_w12342_,
		_w12347_,
		_w12348_
	);
	LUT3 #(
		.INIT('h80)
	) name1836 (
		\wishbone_bd_ram_mem3_reg[125][29]/P0001 ,
		_w11966_,
		_w12012_,
		_w12349_
	);
	LUT3 #(
		.INIT('h80)
	) name1837 (
		\wishbone_bd_ram_mem3_reg[121][29]/P0001 ,
		_w11968_,
		_w12012_,
		_w12350_
	);
	LUT3 #(
		.INIT('h80)
	) name1838 (
		\wishbone_bd_ram_mem3_reg[4][29]/P0001 ,
		_w11929_,
		_w11932_,
		_w12351_
	);
	LUT3 #(
		.INIT('h80)
	) name1839 (
		\wishbone_bd_ram_mem3_reg[81][29]/P0001 ,
		_w11972_,
		_w11977_,
		_w12352_
	);
	LUT4 #(
		.INIT('h0001)
	) name1840 (
		_w12349_,
		_w12350_,
		_w12351_,
		_w12352_,
		_w12353_
	);
	LUT3 #(
		.INIT('h80)
	) name1841 (
		\wishbone_bd_ram_mem3_reg[233][29]/P0001 ,
		_w11968_,
		_w11982_,
		_w12354_
	);
	LUT3 #(
		.INIT('h80)
	) name1842 (
		\wishbone_bd_ram_mem3_reg[191][29]/P0001 ,
		_w11942_,
		_w11973_,
		_w12355_
	);
	LUT3 #(
		.INIT('h80)
	) name1843 (
		\wishbone_bd_ram_mem3_reg[83][29]/P0001 ,
		_w11938_,
		_w11972_,
		_w12356_
	);
	LUT3 #(
		.INIT('h80)
	) name1844 (
		\wishbone_bd_ram_mem3_reg[27][29]/P0001 ,
		_w11935_,
		_w11936_,
		_w12357_
	);
	LUT4 #(
		.INIT('h0001)
	) name1845 (
		_w12354_,
		_w12355_,
		_w12356_,
		_w12357_,
		_w12358_
	);
	LUT3 #(
		.INIT('h80)
	) name1846 (
		\wishbone_bd_ram_mem3_reg[104][29]/P0001 ,
		_w11965_,
		_w11990_,
		_w12359_
	);
	LUT3 #(
		.INIT('h80)
	) name1847 (
		\wishbone_bd_ram_mem3_reg[201][29]/P0001 ,
		_w11945_,
		_w11968_,
		_w12360_
	);
	LUT3 #(
		.INIT('h80)
	) name1848 (
		\wishbone_bd_ram_mem3_reg[75][29]/P0001 ,
		_w11936_,
		_w11949_,
		_w12361_
	);
	LUT3 #(
		.INIT('h80)
	) name1849 (
		\wishbone_bd_ram_mem3_reg[2][29]/P0001 ,
		_w11932_,
		_w11963_,
		_w12362_
	);
	LUT4 #(
		.INIT('h0001)
	) name1850 (
		_w12359_,
		_w12360_,
		_w12361_,
		_w12362_,
		_w12363_
	);
	LUT3 #(
		.INIT('h80)
	) name1851 (
		\wishbone_bd_ram_mem3_reg[67][29]/P0001 ,
		_w11938_,
		_w11949_,
		_w12364_
	);
	LUT3 #(
		.INIT('h80)
	) name1852 (
		\wishbone_bd_ram_mem3_reg[106][29]/P0001 ,
		_w11944_,
		_w11965_,
		_w12365_
	);
	LUT3 #(
		.INIT('h80)
	) name1853 (
		\wishbone_bd_ram_mem3_reg[174][29]/P0001 ,
		_w11930_,
		_w11948_,
		_w12366_
	);
	LUT3 #(
		.INIT('h80)
	) name1854 (
		\wishbone_bd_ram_mem3_reg[181][29]/P0001 ,
		_w11933_,
		_w11942_,
		_w12367_
	);
	LUT4 #(
		.INIT('h0001)
	) name1855 (
		_w12364_,
		_w12365_,
		_w12366_,
		_w12367_,
		_w12368_
	);
	LUT4 #(
		.INIT('h8000)
	) name1856 (
		_w12353_,
		_w12358_,
		_w12363_,
		_w12368_,
		_w12369_
	);
	LUT3 #(
		.INIT('h80)
	) name1857 (
		\wishbone_bd_ram_mem3_reg[224][29]/P0001 ,
		_w11941_,
		_w11982_,
		_w12370_
	);
	LUT3 #(
		.INIT('h80)
	) name1858 (
		\wishbone_bd_ram_mem3_reg[188][29]/P0001 ,
		_w11942_,
		_w11954_,
		_w12371_
	);
	LUT3 #(
		.INIT('h80)
	) name1859 (
		\wishbone_bd_ram_mem3_reg[105][29]/P0001 ,
		_w11965_,
		_w11968_,
		_w12372_
	);
	LUT3 #(
		.INIT('h80)
	) name1860 (
		\wishbone_bd_ram_mem3_reg[58][29]/P0001 ,
		_w11944_,
		_w11979_,
		_w12373_
	);
	LUT4 #(
		.INIT('h0001)
	) name1861 (
		_w12370_,
		_w12371_,
		_w12372_,
		_w12373_,
		_w12374_
	);
	LUT3 #(
		.INIT('h80)
	) name1862 (
		\wishbone_bd_ram_mem3_reg[199][29]/P0001 ,
		_w11945_,
		_w11975_,
		_w12375_
	);
	LUT3 #(
		.INIT('h80)
	) name1863 (
		\wishbone_bd_ram_mem3_reg[49][29]/P0001 ,
		_w11977_,
		_w11979_,
		_w12376_
	);
	LUT3 #(
		.INIT('h80)
	) name1864 (
		\wishbone_bd_ram_mem3_reg[250][29]/P0001 ,
		_w11944_,
		_w11952_,
		_w12377_
	);
	LUT3 #(
		.INIT('h80)
	) name1865 (
		\wishbone_bd_ram_mem3_reg[126][29]/P0001 ,
		_w11948_,
		_w12012_,
		_w12378_
	);
	LUT4 #(
		.INIT('h0001)
	) name1866 (
		_w12375_,
		_w12376_,
		_w12377_,
		_w12378_,
		_w12379_
	);
	LUT3 #(
		.INIT('h80)
	) name1867 (
		\wishbone_bd_ram_mem3_reg[143][29]/P0001 ,
		_w11955_,
		_w11973_,
		_w12380_
	);
	LUT3 #(
		.INIT('h80)
	) name1868 (
		\wishbone_bd_ram_mem3_reg[147][29]/P0001 ,
		_w11938_,
		_w11959_,
		_w12381_
	);
	LUT3 #(
		.INIT('h80)
	) name1869 (
		\wishbone_bd_ram_mem3_reg[100][29]/P0001 ,
		_w11929_,
		_w11965_,
		_w12382_
	);
	LUT3 #(
		.INIT('h80)
	) name1870 (
		\wishbone_bd_ram_mem3_reg[94][29]/P0001 ,
		_w11948_,
		_w11972_,
		_w12383_
	);
	LUT4 #(
		.INIT('h0001)
	) name1871 (
		_w12380_,
		_w12381_,
		_w12382_,
		_w12383_,
		_w12384_
	);
	LUT3 #(
		.INIT('h80)
	) name1872 (
		\wishbone_bd_ram_mem3_reg[193][29]/P0001 ,
		_w11945_,
		_w11977_,
		_w12385_
	);
	LUT3 #(
		.INIT('h80)
	) name1873 (
		\wishbone_bd_ram_mem3_reg[178][29]/P0001 ,
		_w11942_,
		_w11963_,
		_w12386_
	);
	LUT3 #(
		.INIT('h80)
	) name1874 (
		\wishbone_bd_ram_mem3_reg[47][29]/P0001 ,
		_w11957_,
		_w11973_,
		_w12387_
	);
	LUT3 #(
		.INIT('h80)
	) name1875 (
		\wishbone_bd_ram_mem3_reg[225][29]/P0001 ,
		_w11977_,
		_w11982_,
		_w12388_
	);
	LUT4 #(
		.INIT('h0001)
	) name1876 (
		_w12385_,
		_w12386_,
		_w12387_,
		_w12388_,
		_w12389_
	);
	LUT4 #(
		.INIT('h8000)
	) name1877 (
		_w12374_,
		_w12379_,
		_w12384_,
		_w12389_,
		_w12390_
	);
	LUT3 #(
		.INIT('h80)
	) name1878 (
		\wishbone_bd_ram_mem3_reg[123][29]/P0001 ,
		_w11936_,
		_w12012_,
		_w12391_
	);
	LUT3 #(
		.INIT('h80)
	) name1879 (
		\wishbone_bd_ram_mem3_reg[192][29]/P0001 ,
		_w11941_,
		_w11945_,
		_w12392_
	);
	LUT3 #(
		.INIT('h80)
	) name1880 (
		\wishbone_bd_ram_mem3_reg[173][29]/P0001 ,
		_w11930_,
		_w11966_,
		_w12393_
	);
	LUT3 #(
		.INIT('h80)
	) name1881 (
		\wishbone_bd_ram_mem3_reg[120][29]/P0001 ,
		_w11990_,
		_w12012_,
		_w12394_
	);
	LUT4 #(
		.INIT('h0001)
	) name1882 (
		_w12391_,
		_w12392_,
		_w12393_,
		_w12394_,
		_w12395_
	);
	LUT3 #(
		.INIT('h80)
	) name1883 (
		\wishbone_bd_ram_mem3_reg[253][29]/P0001 ,
		_w11952_,
		_w11966_,
		_w12396_
	);
	LUT3 #(
		.INIT('h80)
	) name1884 (
		\wishbone_bd_ram_mem3_reg[243][29]/P0001 ,
		_w11938_,
		_w11952_,
		_w12397_
	);
	LUT3 #(
		.INIT('h80)
	) name1885 (
		\wishbone_bd_ram_mem3_reg[57][29]/P0001 ,
		_w11968_,
		_w11979_,
		_w12398_
	);
	LUT3 #(
		.INIT('h80)
	) name1886 (
		\wishbone_bd_ram_mem3_reg[44][29]/P0001 ,
		_w11954_,
		_w11957_,
		_w12399_
	);
	LUT4 #(
		.INIT('h0001)
	) name1887 (
		_w12396_,
		_w12397_,
		_w12398_,
		_w12399_,
		_w12400_
	);
	LUT3 #(
		.INIT('h80)
	) name1888 (
		\wishbone_bd_ram_mem3_reg[210][29]/P0001 ,
		_w11963_,
		_w11984_,
		_w12401_
	);
	LUT3 #(
		.INIT('h80)
	) name1889 (
		\wishbone_bd_ram_mem3_reg[85][29]/P0001 ,
		_w11933_,
		_w11972_,
		_w12402_
	);
	LUT3 #(
		.INIT('h80)
	) name1890 (
		\wishbone_bd_ram_mem3_reg[134][29]/P0001 ,
		_w11955_,
		_w11986_,
		_w12403_
	);
	LUT3 #(
		.INIT('h80)
	) name1891 (
		\wishbone_bd_ram_mem3_reg[95][29]/P0001 ,
		_w11972_,
		_w11973_,
		_w12404_
	);
	LUT4 #(
		.INIT('h0001)
	) name1892 (
		_w12401_,
		_w12402_,
		_w12403_,
		_w12404_,
		_w12405_
	);
	LUT3 #(
		.INIT('h80)
	) name1893 (
		\wishbone_bd_ram_mem3_reg[48][29]/P0001 ,
		_w11941_,
		_w11979_,
		_w12406_
	);
	LUT3 #(
		.INIT('h80)
	) name1894 (
		\wishbone_bd_ram_mem3_reg[35][29]/P0001 ,
		_w11938_,
		_w11957_,
		_w12407_
	);
	LUT3 #(
		.INIT('h80)
	) name1895 (
		\wishbone_bd_ram_mem3_reg[24][29]/P0001 ,
		_w11935_,
		_w11990_,
		_w12408_
	);
	LUT3 #(
		.INIT('h80)
	) name1896 (
		\wishbone_bd_ram_mem3_reg[231][29]/P0001 ,
		_w11975_,
		_w11982_,
		_w12409_
	);
	LUT4 #(
		.INIT('h0001)
	) name1897 (
		_w12406_,
		_w12407_,
		_w12408_,
		_w12409_,
		_w12410_
	);
	LUT4 #(
		.INIT('h8000)
	) name1898 (
		_w12395_,
		_w12400_,
		_w12405_,
		_w12410_,
		_w12411_
	);
	LUT4 #(
		.INIT('h8000)
	) name1899 (
		_w12348_,
		_w12369_,
		_w12390_,
		_w12411_,
		_w12412_
	);
	LUT3 #(
		.INIT('h80)
	) name1900 (
		\wishbone_bd_ram_mem3_reg[80][29]/P0001 ,
		_w11941_,
		_w11972_,
		_w12413_
	);
	LUT3 #(
		.INIT('h80)
	) name1901 (
		\wishbone_bd_ram_mem3_reg[91][29]/P0001 ,
		_w11936_,
		_w11972_,
		_w12414_
	);
	LUT3 #(
		.INIT('h80)
	) name1902 (
		\wishbone_bd_ram_mem3_reg[212][29]/P0001 ,
		_w11929_,
		_w11984_,
		_w12415_
	);
	LUT3 #(
		.INIT('h80)
	) name1903 (
		\wishbone_bd_ram_mem3_reg[107][29]/P0001 ,
		_w11936_,
		_w11965_,
		_w12416_
	);
	LUT4 #(
		.INIT('h0001)
	) name1904 (
		_w12413_,
		_w12414_,
		_w12415_,
		_w12416_,
		_w12417_
	);
	LUT3 #(
		.INIT('h80)
	) name1905 (
		\wishbone_bd_ram_mem3_reg[247][29]/P0001 ,
		_w11952_,
		_w11975_,
		_w12418_
	);
	LUT3 #(
		.INIT('h80)
	) name1906 (
		\wishbone_bd_ram_mem3_reg[222][29]/P0001 ,
		_w11948_,
		_w11984_,
		_w12419_
	);
	LUT3 #(
		.INIT('h80)
	) name1907 (
		\wishbone_bd_ram_mem3_reg[34][29]/P0001 ,
		_w11957_,
		_w11963_,
		_w12420_
	);
	LUT3 #(
		.INIT('h80)
	) name1908 (
		\wishbone_bd_ram_mem3_reg[17][29]/P0001 ,
		_w11935_,
		_w11977_,
		_w12421_
	);
	LUT4 #(
		.INIT('h0001)
	) name1909 (
		_w12418_,
		_w12419_,
		_w12420_,
		_w12421_,
		_w12422_
	);
	LUT3 #(
		.INIT('h80)
	) name1910 (
		\wishbone_bd_ram_mem3_reg[139][29]/P0001 ,
		_w11936_,
		_w11955_,
		_w12423_
	);
	LUT3 #(
		.INIT('h80)
	) name1911 (
		\wishbone_bd_ram_mem3_reg[142][29]/P0001 ,
		_w11948_,
		_w11955_,
		_w12424_
	);
	LUT3 #(
		.INIT('h80)
	) name1912 (
		\wishbone_bd_ram_mem3_reg[198][29]/P0001 ,
		_w11945_,
		_w11986_,
		_w12425_
	);
	LUT3 #(
		.INIT('h80)
	) name1913 (
		\wishbone_bd_ram_mem3_reg[244][29]/P0001 ,
		_w11929_,
		_w11952_,
		_w12426_
	);
	LUT4 #(
		.INIT('h0001)
	) name1914 (
		_w12423_,
		_w12424_,
		_w12425_,
		_w12426_,
		_w12427_
	);
	LUT3 #(
		.INIT('h80)
	) name1915 (
		\wishbone_bd_ram_mem3_reg[169][29]/P0001 ,
		_w11930_,
		_w11968_,
		_w12428_
	);
	LUT3 #(
		.INIT('h80)
	) name1916 (
		\wishbone_bd_ram_mem3_reg[149][29]/P0001 ,
		_w11933_,
		_w11959_,
		_w12429_
	);
	LUT3 #(
		.INIT('h80)
	) name1917 (
		\wishbone_bd_ram_mem3_reg[182][29]/P0001 ,
		_w11942_,
		_w11986_,
		_w12430_
	);
	LUT3 #(
		.INIT('h80)
	) name1918 (
		\wishbone_bd_ram_mem3_reg[154][29]/P0001 ,
		_w11944_,
		_w11959_,
		_w12431_
	);
	LUT4 #(
		.INIT('h0001)
	) name1919 (
		_w12428_,
		_w12429_,
		_w12430_,
		_w12431_,
		_w12432_
	);
	LUT4 #(
		.INIT('h8000)
	) name1920 (
		_w12417_,
		_w12422_,
		_w12427_,
		_w12432_,
		_w12433_
	);
	LUT3 #(
		.INIT('h80)
	) name1921 (
		\wishbone_bd_ram_mem3_reg[144][29]/P0001 ,
		_w11941_,
		_w11959_,
		_w12434_
	);
	LUT3 #(
		.INIT('h80)
	) name1922 (
		\wishbone_bd_ram_mem3_reg[61][29]/P0001 ,
		_w11966_,
		_w11979_,
		_w12435_
	);
	LUT3 #(
		.INIT('h80)
	) name1923 (
		\wishbone_bd_ram_mem3_reg[135][29]/P0001 ,
		_w11955_,
		_w11975_,
		_w12436_
	);
	LUT3 #(
		.INIT('h80)
	) name1924 (
		\wishbone_bd_ram_mem3_reg[66][29]/P0001 ,
		_w11949_,
		_w11963_,
		_w12437_
	);
	LUT4 #(
		.INIT('h0001)
	) name1925 (
		_w12434_,
		_w12435_,
		_w12436_,
		_w12437_,
		_w12438_
	);
	LUT3 #(
		.INIT('h80)
	) name1926 (
		\wishbone_bd_ram_mem3_reg[175][29]/P0001 ,
		_w11930_,
		_w11973_,
		_w12439_
	);
	LUT3 #(
		.INIT('h80)
	) name1927 (
		\wishbone_bd_ram_mem3_reg[141][29]/P0001 ,
		_w11955_,
		_w11966_,
		_w12440_
	);
	LUT3 #(
		.INIT('h80)
	) name1928 (
		\wishbone_bd_ram_mem3_reg[189][29]/P0001 ,
		_w11942_,
		_w11966_,
		_w12441_
	);
	LUT3 #(
		.INIT('h80)
	) name1929 (
		\wishbone_bd_ram_mem3_reg[185][29]/P0001 ,
		_w11942_,
		_w11968_,
		_w12442_
	);
	LUT4 #(
		.INIT('h0001)
	) name1930 (
		_w12439_,
		_w12440_,
		_w12441_,
		_w12442_,
		_w12443_
	);
	LUT3 #(
		.INIT('h80)
	) name1931 (
		\wishbone_bd_ram_mem3_reg[13][29]/P0001 ,
		_w11932_,
		_w11966_,
		_w12444_
	);
	LUT3 #(
		.INIT('h80)
	) name1932 (
		\wishbone_bd_ram_mem3_reg[162][29]/P0001 ,
		_w11930_,
		_w11963_,
		_w12445_
	);
	LUT3 #(
		.INIT('h80)
	) name1933 (
		\wishbone_bd_ram_mem3_reg[131][29]/P0001 ,
		_w11938_,
		_w11955_,
		_w12446_
	);
	LUT3 #(
		.INIT('h80)
	) name1934 (
		\wishbone_bd_ram_mem3_reg[22][29]/P0001 ,
		_w11935_,
		_w11986_,
		_w12447_
	);
	LUT4 #(
		.INIT('h0001)
	) name1935 (
		_w12444_,
		_w12445_,
		_w12446_,
		_w12447_,
		_w12448_
	);
	LUT3 #(
		.INIT('h80)
	) name1936 (
		\wishbone_bd_ram_mem3_reg[103][29]/P0001 ,
		_w11965_,
		_w11975_,
		_w12449_
	);
	LUT3 #(
		.INIT('h80)
	) name1937 (
		\wishbone_bd_ram_mem3_reg[240][29]/P0001 ,
		_w11941_,
		_w11952_,
		_w12450_
	);
	LUT3 #(
		.INIT('h80)
	) name1938 (
		\wishbone_bd_ram_mem3_reg[170][29]/P0001 ,
		_w11930_,
		_w11944_,
		_w12451_
	);
	LUT3 #(
		.INIT('h80)
	) name1939 (
		\wishbone_bd_ram_mem3_reg[136][29]/P0001 ,
		_w11955_,
		_w11990_,
		_w12452_
	);
	LUT4 #(
		.INIT('h0001)
	) name1940 (
		_w12449_,
		_w12450_,
		_w12451_,
		_w12452_,
		_w12453_
	);
	LUT4 #(
		.INIT('h8000)
	) name1941 (
		_w12438_,
		_w12443_,
		_w12448_,
		_w12453_,
		_w12454_
	);
	LUT3 #(
		.INIT('h80)
	) name1942 (
		\wishbone_bd_ram_mem3_reg[6][29]/P0001 ,
		_w11932_,
		_w11986_,
		_w12455_
	);
	LUT3 #(
		.INIT('h80)
	) name1943 (
		\wishbone_bd_ram_mem3_reg[110][29]/P0001 ,
		_w11948_,
		_w11965_,
		_w12456_
	);
	LUT3 #(
		.INIT('h80)
	) name1944 (
		\wishbone_bd_ram_mem3_reg[89][29]/P0001 ,
		_w11968_,
		_w11972_,
		_w12457_
	);
	LUT3 #(
		.INIT('h80)
	) name1945 (
		\wishbone_bd_ram_mem3_reg[64][29]/P0001 ,
		_w11941_,
		_w11949_,
		_w12458_
	);
	LUT4 #(
		.INIT('h0001)
	) name1946 (
		_w12455_,
		_w12456_,
		_w12457_,
		_w12458_,
		_w12459_
	);
	LUT3 #(
		.INIT('h80)
	) name1947 (
		\wishbone_bd_ram_mem3_reg[220][29]/P0001 ,
		_w11954_,
		_w11984_,
		_w12460_
	);
	LUT3 #(
		.INIT('h80)
	) name1948 (
		\wishbone_bd_ram_mem3_reg[216][29]/P0001 ,
		_w11984_,
		_w11990_,
		_w12461_
	);
	LUT3 #(
		.INIT('h80)
	) name1949 (
		\wishbone_bd_ram_mem3_reg[12][29]/P0001 ,
		_w11932_,
		_w11954_,
		_w12462_
	);
	LUT3 #(
		.INIT('h80)
	) name1950 (
		\wishbone_bd_ram_mem3_reg[56][29]/P0001 ,
		_w11979_,
		_w11990_,
		_w12463_
	);
	LUT4 #(
		.INIT('h0001)
	) name1951 (
		_w12460_,
		_w12461_,
		_w12462_,
		_w12463_,
		_w12464_
	);
	LUT3 #(
		.INIT('h80)
	) name1952 (
		\wishbone_bd_ram_mem3_reg[194][29]/P0001 ,
		_w11945_,
		_w11963_,
		_w12465_
	);
	LUT3 #(
		.INIT('h80)
	) name1953 (
		\wishbone_bd_ram_mem3_reg[39][29]/P0001 ,
		_w11957_,
		_w11975_,
		_w12466_
	);
	LUT3 #(
		.INIT('h80)
	) name1954 (
		\wishbone_bd_ram_mem3_reg[237][29]/P0001 ,
		_w11966_,
		_w11982_,
		_w12467_
	);
	LUT3 #(
		.INIT('h80)
	) name1955 (
		\wishbone_bd_ram_mem3_reg[204][29]/P0001 ,
		_w11945_,
		_w11954_,
		_w12468_
	);
	LUT4 #(
		.INIT('h0001)
	) name1956 (
		_w12465_,
		_w12466_,
		_w12467_,
		_w12468_,
		_w12469_
	);
	LUT3 #(
		.INIT('h80)
	) name1957 (
		\wishbone_bd_ram_mem3_reg[171][29]/P0001 ,
		_w11930_,
		_w11936_,
		_w12470_
	);
	LUT3 #(
		.INIT('h80)
	) name1958 (
		\wishbone_bd_ram_mem3_reg[239][29]/P0001 ,
		_w11973_,
		_w11982_,
		_w12471_
	);
	LUT3 #(
		.INIT('h80)
	) name1959 (
		\wishbone_bd_ram_mem3_reg[93][29]/P0001 ,
		_w11966_,
		_w11972_,
		_w12472_
	);
	LUT3 #(
		.INIT('h80)
	) name1960 (
		\wishbone_bd_ram_mem3_reg[59][29]/P0001 ,
		_w11936_,
		_w11979_,
		_w12473_
	);
	LUT4 #(
		.INIT('h0001)
	) name1961 (
		_w12470_,
		_w12471_,
		_w12472_,
		_w12473_,
		_w12474_
	);
	LUT4 #(
		.INIT('h8000)
	) name1962 (
		_w12459_,
		_w12464_,
		_w12469_,
		_w12474_,
		_w12475_
	);
	LUT3 #(
		.INIT('h80)
	) name1963 (
		\wishbone_bd_ram_mem3_reg[38][29]/P0001 ,
		_w11957_,
		_w11986_,
		_w12476_
	);
	LUT3 #(
		.INIT('h80)
	) name1964 (
		\wishbone_bd_ram_mem3_reg[45][29]/P0001 ,
		_w11957_,
		_w11966_,
		_w12477_
	);
	LUT3 #(
		.INIT('h80)
	) name1965 (
		\wishbone_bd_ram_mem3_reg[195][29]/P0001 ,
		_w11938_,
		_w11945_,
		_w12478_
	);
	LUT3 #(
		.INIT('h80)
	) name1966 (
		\wishbone_bd_ram_mem3_reg[196][29]/P0001 ,
		_w11929_,
		_w11945_,
		_w12479_
	);
	LUT4 #(
		.INIT('h0001)
	) name1967 (
		_w12476_,
		_w12477_,
		_w12478_,
		_w12479_,
		_w12480_
	);
	LUT3 #(
		.INIT('h80)
	) name1968 (
		\wishbone_bd_ram_mem3_reg[101][29]/P0001 ,
		_w11933_,
		_w11965_,
		_w12481_
	);
	LUT3 #(
		.INIT('h80)
	) name1969 (
		\wishbone_bd_ram_mem3_reg[226][29]/P0001 ,
		_w11963_,
		_w11982_,
		_w12482_
	);
	LUT3 #(
		.INIT('h80)
	) name1970 (
		\wishbone_bd_ram_mem3_reg[159][29]/P0001 ,
		_w11959_,
		_w11973_,
		_w12483_
	);
	LUT3 #(
		.INIT('h80)
	) name1971 (
		\wishbone_bd_ram_mem3_reg[116][29]/P0001 ,
		_w11929_,
		_w12012_,
		_w12484_
	);
	LUT4 #(
		.INIT('h0001)
	) name1972 (
		_w12481_,
		_w12482_,
		_w12483_,
		_w12484_,
		_w12485_
	);
	LUT3 #(
		.INIT('h80)
	) name1973 (
		\wishbone_bd_ram_mem3_reg[203][29]/P0001 ,
		_w11936_,
		_w11945_,
		_w12486_
	);
	LUT3 #(
		.INIT('h80)
	) name1974 (
		\wishbone_bd_ram_mem3_reg[117][29]/P0001 ,
		_w11933_,
		_w12012_,
		_w12487_
	);
	LUT3 #(
		.INIT('h80)
	) name1975 (
		\wishbone_bd_ram_mem3_reg[73][29]/P0001 ,
		_w11949_,
		_w11968_,
		_w12488_
	);
	LUT3 #(
		.INIT('h80)
	) name1976 (
		\wishbone_bd_ram_mem3_reg[251][29]/P0001 ,
		_w11936_,
		_w11952_,
		_w12489_
	);
	LUT4 #(
		.INIT('h0001)
	) name1977 (
		_w12486_,
		_w12487_,
		_w12488_,
		_w12489_,
		_w12490_
	);
	LUT3 #(
		.INIT('h80)
	) name1978 (
		\wishbone_bd_ram_mem3_reg[183][29]/P0001 ,
		_w11942_,
		_w11975_,
		_w12491_
	);
	LUT3 #(
		.INIT('h80)
	) name1979 (
		\wishbone_bd_ram_mem3_reg[252][29]/P0001 ,
		_w11952_,
		_w11954_,
		_w12492_
	);
	LUT3 #(
		.INIT('h80)
	) name1980 (
		\wishbone_bd_ram_mem3_reg[180][29]/P0001 ,
		_w11929_,
		_w11942_,
		_w12493_
	);
	LUT3 #(
		.INIT('h80)
	) name1981 (
		\wishbone_bd_ram_mem3_reg[29][29]/P0001 ,
		_w11935_,
		_w11966_,
		_w12494_
	);
	LUT4 #(
		.INIT('h0001)
	) name1982 (
		_w12491_,
		_w12492_,
		_w12493_,
		_w12494_,
		_w12495_
	);
	LUT4 #(
		.INIT('h8000)
	) name1983 (
		_w12480_,
		_w12485_,
		_w12490_,
		_w12495_,
		_w12496_
	);
	LUT4 #(
		.INIT('h8000)
	) name1984 (
		_w12433_,
		_w12454_,
		_w12475_,
		_w12496_,
		_w12497_
	);
	LUT3 #(
		.INIT('h80)
	) name1985 (
		\wishbone_bd_ram_mem3_reg[40][29]/P0001 ,
		_w11957_,
		_w11990_,
		_w12498_
	);
	LUT3 #(
		.INIT('h80)
	) name1986 (
		\wishbone_bd_ram_mem3_reg[1][29]/P0001 ,
		_w11932_,
		_w11977_,
		_w12499_
	);
	LUT3 #(
		.INIT('h80)
	) name1987 (
		\wishbone_bd_ram_mem3_reg[82][29]/P0001 ,
		_w11963_,
		_w11972_,
		_w12500_
	);
	LUT3 #(
		.INIT('h80)
	) name1988 (
		\wishbone_bd_ram_mem3_reg[206][29]/P0001 ,
		_w11945_,
		_w11948_,
		_w12501_
	);
	LUT4 #(
		.INIT('h0001)
	) name1989 (
		_w12498_,
		_w12499_,
		_w12500_,
		_w12501_,
		_w12502_
	);
	LUT3 #(
		.INIT('h80)
	) name1990 (
		\wishbone_bd_ram_mem3_reg[157][29]/P0001 ,
		_w11959_,
		_w11966_,
		_w12503_
	);
	LUT3 #(
		.INIT('h80)
	) name1991 (
		\wishbone_bd_ram_mem3_reg[8][29]/P0001 ,
		_w11932_,
		_w11990_,
		_w12504_
	);
	LUT3 #(
		.INIT('h80)
	) name1992 (
		\wishbone_bd_ram_mem3_reg[213][29]/P0001 ,
		_w11933_,
		_w11984_,
		_w12505_
	);
	LUT3 #(
		.INIT('h80)
	) name1993 (
		\wishbone_bd_ram_mem3_reg[63][29]/P0001 ,
		_w11973_,
		_w11979_,
		_w12506_
	);
	LUT4 #(
		.INIT('h0001)
	) name1994 (
		_w12503_,
		_w12504_,
		_w12505_,
		_w12506_,
		_w12507_
	);
	LUT3 #(
		.INIT('h80)
	) name1995 (
		\wishbone_bd_ram_mem3_reg[166][29]/P0001 ,
		_w11930_,
		_w11986_,
		_w12508_
	);
	LUT3 #(
		.INIT('h80)
	) name1996 (
		\wishbone_bd_ram_mem3_reg[69][29]/P0001 ,
		_w11933_,
		_w11949_,
		_w12509_
	);
	LUT3 #(
		.INIT('h80)
	) name1997 (
		\wishbone_bd_ram_mem3_reg[84][29]/P0001 ,
		_w11929_,
		_w11972_,
		_w12510_
	);
	LUT3 #(
		.INIT('h80)
	) name1998 (
		\wishbone_bd_ram_mem3_reg[53][29]/P0001 ,
		_w11933_,
		_w11979_,
		_w12511_
	);
	LUT4 #(
		.INIT('h0001)
	) name1999 (
		_w12508_,
		_w12509_,
		_w12510_,
		_w12511_,
		_w12512_
	);
	LUT3 #(
		.INIT('h80)
	) name2000 (
		\wishbone_bd_ram_mem3_reg[148][29]/P0001 ,
		_w11929_,
		_w11959_,
		_w12513_
	);
	LUT3 #(
		.INIT('h80)
	) name2001 (
		\wishbone_bd_ram_mem3_reg[98][29]/P0001 ,
		_w11963_,
		_w11965_,
		_w12514_
	);
	LUT3 #(
		.INIT('h80)
	) name2002 (
		\wishbone_bd_ram_mem3_reg[186][29]/P0001 ,
		_w11942_,
		_w11944_,
		_w12515_
	);
	LUT3 #(
		.INIT('h80)
	) name2003 (
		\wishbone_bd_ram_mem3_reg[7][29]/P0001 ,
		_w11932_,
		_w11975_,
		_w12516_
	);
	LUT4 #(
		.INIT('h0001)
	) name2004 (
		_w12513_,
		_w12514_,
		_w12515_,
		_w12516_,
		_w12517_
	);
	LUT4 #(
		.INIT('h8000)
	) name2005 (
		_w12502_,
		_w12507_,
		_w12512_,
		_w12517_,
		_w12518_
	);
	LUT3 #(
		.INIT('h80)
	) name2006 (
		\wishbone_bd_ram_mem3_reg[221][29]/P0001 ,
		_w11966_,
		_w11984_,
		_w12519_
	);
	LUT3 #(
		.INIT('h80)
	) name2007 (
		\wishbone_bd_ram_mem3_reg[0][29]/P0001 ,
		_w11932_,
		_w11941_,
		_w12520_
	);
	LUT3 #(
		.INIT('h80)
	) name2008 (
		\wishbone_bd_ram_mem3_reg[50][29]/P0001 ,
		_w11963_,
		_w11979_,
		_w12521_
	);
	LUT3 #(
		.INIT('h80)
	) name2009 (
		\wishbone_bd_ram_mem3_reg[230][29]/P0001 ,
		_w11982_,
		_w11986_,
		_w12522_
	);
	LUT4 #(
		.INIT('h0001)
	) name2010 (
		_w12519_,
		_w12520_,
		_w12521_,
		_w12522_,
		_w12523_
	);
	LUT3 #(
		.INIT('h80)
	) name2011 (
		\wishbone_bd_ram_mem3_reg[190][29]/P0001 ,
		_w11942_,
		_w11948_,
		_w12524_
	);
	LUT3 #(
		.INIT('h80)
	) name2012 (
		\wishbone_bd_ram_mem3_reg[232][29]/P0001 ,
		_w11982_,
		_w11990_,
		_w12525_
	);
	LUT3 #(
		.INIT('h80)
	) name2013 (
		\wishbone_bd_ram_mem3_reg[228][29]/P0001 ,
		_w11929_,
		_w11982_,
		_w12526_
	);
	LUT3 #(
		.INIT('h80)
	) name2014 (
		\wishbone_bd_ram_mem3_reg[214][29]/P0001 ,
		_w11984_,
		_w11986_,
		_w12527_
	);
	LUT4 #(
		.INIT('h0001)
	) name2015 (
		_w12524_,
		_w12525_,
		_w12526_,
		_w12527_,
		_w12528_
	);
	LUT3 #(
		.INIT('h80)
	) name2016 (
		\wishbone_bd_ram_mem3_reg[119][29]/P0001 ,
		_w11975_,
		_w12012_,
		_w12529_
	);
	LUT3 #(
		.INIT('h80)
	) name2017 (
		\wishbone_bd_ram_mem3_reg[9][29]/P0001 ,
		_w11932_,
		_w11968_,
		_w12530_
	);
	LUT3 #(
		.INIT('h80)
	) name2018 (
		\wishbone_bd_ram_mem3_reg[215][29]/P0001 ,
		_w11975_,
		_w11984_,
		_w12531_
	);
	LUT3 #(
		.INIT('h80)
	) name2019 (
		\wishbone_bd_ram_mem3_reg[74][29]/P0001 ,
		_w11944_,
		_w11949_,
		_w12532_
	);
	LUT4 #(
		.INIT('h0001)
	) name2020 (
		_w12529_,
		_w12530_,
		_w12531_,
		_w12532_,
		_w12533_
	);
	LUT3 #(
		.INIT('h80)
	) name2021 (
		\wishbone_bd_ram_mem3_reg[32][29]/P0001 ,
		_w11941_,
		_w11957_,
		_w12534_
	);
	LUT3 #(
		.INIT('h80)
	) name2022 (
		\wishbone_bd_ram_mem3_reg[41][29]/P0001 ,
		_w11957_,
		_w11968_,
		_w12535_
	);
	LUT3 #(
		.INIT('h80)
	) name2023 (
		\wishbone_bd_ram_mem3_reg[51][29]/P0001 ,
		_w11938_,
		_w11979_,
		_w12536_
	);
	LUT3 #(
		.INIT('h80)
	) name2024 (
		\wishbone_bd_ram_mem3_reg[208][29]/P0001 ,
		_w11941_,
		_w11984_,
		_w12537_
	);
	LUT4 #(
		.INIT('h0001)
	) name2025 (
		_w12534_,
		_w12535_,
		_w12536_,
		_w12537_,
		_w12538_
	);
	LUT4 #(
		.INIT('h8000)
	) name2026 (
		_w12523_,
		_w12528_,
		_w12533_,
		_w12538_,
		_w12539_
	);
	LUT3 #(
		.INIT('h80)
	) name2027 (
		\wishbone_bd_ram_mem3_reg[249][29]/P0001 ,
		_w11952_,
		_w11968_,
		_w12540_
	);
	LUT3 #(
		.INIT('h80)
	) name2028 (
		\wishbone_bd_ram_mem3_reg[15][29]/P0001 ,
		_w11932_,
		_w11973_,
		_w12541_
	);
	LUT3 #(
		.INIT('h80)
	) name2029 (
		\wishbone_bd_ram_mem3_reg[68][29]/P0001 ,
		_w11929_,
		_w11949_,
		_w12542_
	);
	LUT3 #(
		.INIT('h80)
	) name2030 (
		\wishbone_bd_ram_mem3_reg[72][29]/P0001 ,
		_w11949_,
		_w11990_,
		_w12543_
	);
	LUT4 #(
		.INIT('h0001)
	) name2031 (
		_w12540_,
		_w12541_,
		_w12542_,
		_w12543_,
		_w12544_
	);
	LUT3 #(
		.INIT('h80)
	) name2032 (
		\wishbone_bd_ram_mem3_reg[87][29]/P0001 ,
		_w11972_,
		_w11975_,
		_w12545_
	);
	LUT3 #(
		.INIT('h80)
	) name2033 (
		\wishbone_bd_ram_mem3_reg[130][29]/P0001 ,
		_w11955_,
		_w11963_,
		_w12546_
	);
	LUT3 #(
		.INIT('h80)
	) name2034 (
		\wishbone_bd_ram_mem3_reg[138][29]/P0001 ,
		_w11944_,
		_w11955_,
		_w12547_
	);
	LUT3 #(
		.INIT('h80)
	) name2035 (
		\wishbone_bd_ram_mem3_reg[115][29]/P0001 ,
		_w11938_,
		_w12012_,
		_w12548_
	);
	LUT4 #(
		.INIT('h0001)
	) name2036 (
		_w12545_,
		_w12546_,
		_w12547_,
		_w12548_,
		_w12549_
	);
	LUT3 #(
		.INIT('h80)
	) name2037 (
		\wishbone_bd_ram_mem3_reg[43][29]/P0001 ,
		_w11936_,
		_w11957_,
		_w12550_
	);
	LUT3 #(
		.INIT('h80)
	) name2038 (
		\wishbone_bd_ram_mem3_reg[241][29]/P0001 ,
		_w11952_,
		_w11977_,
		_w12551_
	);
	LUT3 #(
		.INIT('h80)
	) name2039 (
		\wishbone_bd_ram_mem3_reg[118][29]/P0001 ,
		_w11986_,
		_w12012_,
		_w12552_
	);
	LUT3 #(
		.INIT('h80)
	) name2040 (
		\wishbone_bd_ram_mem3_reg[242][29]/P0001 ,
		_w11952_,
		_w11963_,
		_w12553_
	);
	LUT4 #(
		.INIT('h0001)
	) name2041 (
		_w12550_,
		_w12551_,
		_w12552_,
		_w12553_,
		_w12554_
	);
	LUT3 #(
		.INIT('h80)
	) name2042 (
		\wishbone_bd_ram_mem3_reg[60][29]/P0001 ,
		_w11954_,
		_w11979_,
		_w12555_
	);
	LUT3 #(
		.INIT('h80)
	) name2043 (
		\wishbone_bd_ram_mem3_reg[168][29]/P0001 ,
		_w11930_,
		_w11990_,
		_w12556_
	);
	LUT3 #(
		.INIT('h80)
	) name2044 (
		\wishbone_bd_ram_mem3_reg[122][29]/P0001 ,
		_w11944_,
		_w12012_,
		_w12557_
	);
	LUT3 #(
		.INIT('h80)
	) name2045 (
		\wishbone_bd_ram_mem3_reg[109][29]/P0001 ,
		_w11965_,
		_w11966_,
		_w12558_
	);
	LUT4 #(
		.INIT('h0001)
	) name2046 (
		_w12555_,
		_w12556_,
		_w12557_,
		_w12558_,
		_w12559_
	);
	LUT4 #(
		.INIT('h8000)
	) name2047 (
		_w12544_,
		_w12549_,
		_w12554_,
		_w12559_,
		_w12560_
	);
	LUT3 #(
		.INIT('h80)
	) name2048 (
		\wishbone_bd_ram_mem3_reg[108][29]/P0001 ,
		_w11954_,
		_w11965_,
		_w12561_
	);
	LUT3 #(
		.INIT('h80)
	) name2049 (
		\wishbone_bd_ram_mem3_reg[211][29]/P0001 ,
		_w11938_,
		_w11984_,
		_w12562_
	);
	LUT3 #(
		.INIT('h80)
	) name2050 (
		\wishbone_bd_ram_mem3_reg[97][29]/P0001 ,
		_w11965_,
		_w11977_,
		_w12563_
	);
	LUT3 #(
		.INIT('h80)
	) name2051 (
		\wishbone_bd_ram_mem3_reg[19][29]/P0001 ,
		_w11935_,
		_w11938_,
		_w12564_
	);
	LUT4 #(
		.INIT('h0001)
	) name2052 (
		_w12561_,
		_w12562_,
		_w12563_,
		_w12564_,
		_w12565_
	);
	LUT3 #(
		.INIT('h80)
	) name2053 (
		\wishbone_bd_ram_mem3_reg[145][29]/P0001 ,
		_w11959_,
		_w11977_,
		_w12566_
	);
	LUT3 #(
		.INIT('h80)
	) name2054 (
		\wishbone_bd_ram_mem3_reg[114][29]/P0001 ,
		_w11963_,
		_w12012_,
		_w12567_
	);
	LUT3 #(
		.INIT('h80)
	) name2055 (
		\wishbone_bd_ram_mem3_reg[246][29]/P0001 ,
		_w11952_,
		_w11986_,
		_w12568_
	);
	LUT3 #(
		.INIT('h80)
	) name2056 (
		\wishbone_bd_ram_mem3_reg[255][29]/P0001 ,
		_w11952_,
		_w11973_,
		_w12569_
	);
	LUT4 #(
		.INIT('h0001)
	) name2057 (
		_w12566_,
		_w12567_,
		_w12568_,
		_w12569_,
		_w12570_
	);
	LUT3 #(
		.INIT('h80)
	) name2058 (
		\wishbone_bd_ram_mem3_reg[207][29]/P0001 ,
		_w11945_,
		_w11973_,
		_w12571_
	);
	LUT3 #(
		.INIT('h80)
	) name2059 (
		\wishbone_bd_ram_mem3_reg[20][29]/P0001 ,
		_w11929_,
		_w11935_,
		_w12572_
	);
	LUT3 #(
		.INIT('h80)
	) name2060 (
		\wishbone_bd_ram_mem3_reg[25][29]/P0001 ,
		_w11935_,
		_w11968_,
		_w12573_
	);
	LUT3 #(
		.INIT('h80)
	) name2061 (
		\wishbone_bd_ram_mem3_reg[238][29]/P0001 ,
		_w11948_,
		_w11982_,
		_w12574_
	);
	LUT4 #(
		.INIT('h0001)
	) name2062 (
		_w12571_,
		_w12572_,
		_w12573_,
		_w12574_,
		_w12575_
	);
	LUT3 #(
		.INIT('h80)
	) name2063 (
		\wishbone_bd_ram_mem3_reg[11][29]/P0001 ,
		_w11932_,
		_w11936_,
		_w12576_
	);
	LUT3 #(
		.INIT('h80)
	) name2064 (
		\wishbone_bd_ram_mem3_reg[161][29]/P0001 ,
		_w11930_,
		_w11977_,
		_w12577_
	);
	LUT3 #(
		.INIT('h80)
	) name2065 (
		\wishbone_bd_ram_mem3_reg[21][29]/P0001 ,
		_w11933_,
		_w11935_,
		_w12578_
	);
	LUT3 #(
		.INIT('h80)
	) name2066 (
		\wishbone_bd_ram_mem3_reg[33][29]/P0001 ,
		_w11957_,
		_w11977_,
		_w12579_
	);
	LUT4 #(
		.INIT('h0001)
	) name2067 (
		_w12576_,
		_w12577_,
		_w12578_,
		_w12579_,
		_w12580_
	);
	LUT4 #(
		.INIT('h8000)
	) name2068 (
		_w12565_,
		_w12570_,
		_w12575_,
		_w12580_,
		_w12581_
	);
	LUT4 #(
		.INIT('h8000)
	) name2069 (
		_w12518_,
		_w12539_,
		_w12560_,
		_w12581_,
		_w12582_
	);
	LUT3 #(
		.INIT('h80)
	) name2070 (
		\wishbone_bd_ram_mem3_reg[62][29]/P0001 ,
		_w11948_,
		_w11979_,
		_w12583_
	);
	LUT3 #(
		.INIT('h80)
	) name2071 (
		\wishbone_bd_ram_mem3_reg[248][29]/P0001 ,
		_w11952_,
		_w11990_,
		_w12584_
	);
	LUT3 #(
		.INIT('h80)
	) name2072 (
		\wishbone_bd_ram_mem3_reg[152][29]/P0001 ,
		_w11959_,
		_w11990_,
		_w12585_
	);
	LUT3 #(
		.INIT('h80)
	) name2073 (
		\wishbone_bd_ram_mem3_reg[172][29]/P0001 ,
		_w11930_,
		_w11954_,
		_w12586_
	);
	LUT4 #(
		.INIT('h0001)
	) name2074 (
		_w12583_,
		_w12584_,
		_w12585_,
		_w12586_,
		_w12587_
	);
	LUT3 #(
		.INIT('h80)
	) name2075 (
		\wishbone_bd_ram_mem3_reg[146][29]/P0001 ,
		_w11959_,
		_w11963_,
		_w12588_
	);
	LUT3 #(
		.INIT('h80)
	) name2076 (
		\wishbone_bd_ram_mem3_reg[54][29]/P0001 ,
		_w11979_,
		_w11986_,
		_w12589_
	);
	LUT3 #(
		.INIT('h80)
	) name2077 (
		\wishbone_bd_ram_mem3_reg[128][29]/P0001 ,
		_w11941_,
		_w11955_,
		_w12590_
	);
	LUT3 #(
		.INIT('h80)
	) name2078 (
		\wishbone_bd_ram_mem3_reg[229][29]/P0001 ,
		_w11933_,
		_w11982_,
		_w12591_
	);
	LUT4 #(
		.INIT('h0001)
	) name2079 (
		_w12588_,
		_w12589_,
		_w12590_,
		_w12591_,
		_w12592_
	);
	LUT3 #(
		.INIT('h80)
	) name2080 (
		\wishbone_bd_ram_mem3_reg[165][29]/P0001 ,
		_w11930_,
		_w11933_,
		_w12593_
	);
	LUT3 #(
		.INIT('h80)
	) name2081 (
		\wishbone_bd_ram_mem3_reg[254][29]/P0001 ,
		_w11948_,
		_w11952_,
		_w12594_
	);
	LUT3 #(
		.INIT('h80)
	) name2082 (
		\wishbone_bd_ram_mem3_reg[76][29]/P0001 ,
		_w11949_,
		_w11954_,
		_w12595_
	);
	LUT3 #(
		.INIT('h80)
	) name2083 (
		\wishbone_bd_ram_mem3_reg[179][29]/P0001 ,
		_w11938_,
		_w11942_,
		_w12596_
	);
	LUT4 #(
		.INIT('h0001)
	) name2084 (
		_w12593_,
		_w12594_,
		_w12595_,
		_w12596_,
		_w12597_
	);
	LUT3 #(
		.INIT('h80)
	) name2085 (
		\wishbone_bd_ram_mem3_reg[28][29]/P0001 ,
		_w11935_,
		_w11954_,
		_w12598_
	);
	LUT3 #(
		.INIT('h80)
	) name2086 (
		\wishbone_bd_ram_mem3_reg[3][29]/P0001 ,
		_w11932_,
		_w11938_,
		_w12599_
	);
	LUT3 #(
		.INIT('h80)
	) name2087 (
		\wishbone_bd_ram_mem3_reg[137][29]/P0001 ,
		_w11955_,
		_w11968_,
		_w12600_
	);
	LUT3 #(
		.INIT('h80)
	) name2088 (
		\wishbone_bd_ram_mem3_reg[78][29]/P0001 ,
		_w11948_,
		_w11949_,
		_w12601_
	);
	LUT4 #(
		.INIT('h0001)
	) name2089 (
		_w12598_,
		_w12599_,
		_w12600_,
		_w12601_,
		_w12602_
	);
	LUT4 #(
		.INIT('h8000)
	) name2090 (
		_w12587_,
		_w12592_,
		_w12597_,
		_w12602_,
		_w12603_
	);
	LUT3 #(
		.INIT('h80)
	) name2091 (
		\wishbone_bd_ram_mem3_reg[151][29]/P0001 ,
		_w11959_,
		_w11975_,
		_w12604_
	);
	LUT3 #(
		.INIT('h80)
	) name2092 (
		\wishbone_bd_ram_mem3_reg[14][29]/P0001 ,
		_w11932_,
		_w11948_,
		_w12605_
	);
	LUT3 #(
		.INIT('h80)
	) name2093 (
		\wishbone_bd_ram_mem3_reg[26][29]/P0001 ,
		_w11935_,
		_w11944_,
		_w12606_
	);
	LUT3 #(
		.INIT('h80)
	) name2094 (
		\wishbone_bd_ram_mem3_reg[200][29]/P0001 ,
		_w11945_,
		_w11990_,
		_w12607_
	);
	LUT4 #(
		.INIT('h0001)
	) name2095 (
		_w12604_,
		_w12605_,
		_w12606_,
		_w12607_,
		_w12608_
	);
	LUT3 #(
		.INIT('h80)
	) name2096 (
		\wishbone_bd_ram_mem3_reg[102][29]/P0001 ,
		_w11965_,
		_w11986_,
		_w12609_
	);
	LUT3 #(
		.INIT('h80)
	) name2097 (
		\wishbone_bd_ram_mem3_reg[129][29]/P0001 ,
		_w11955_,
		_w11977_,
		_w12610_
	);
	LUT3 #(
		.INIT('h80)
	) name2098 (
		\wishbone_bd_ram_mem3_reg[10][29]/P0001 ,
		_w11932_,
		_w11944_,
		_w12611_
	);
	LUT3 #(
		.INIT('h80)
	) name2099 (
		\wishbone_bd_ram_mem3_reg[163][29]/P0001 ,
		_w11930_,
		_w11938_,
		_w12612_
	);
	LUT4 #(
		.INIT('h0001)
	) name2100 (
		_w12609_,
		_w12610_,
		_w12611_,
		_w12612_,
		_w12613_
	);
	LUT3 #(
		.INIT('h80)
	) name2101 (
		\wishbone_bd_ram_mem3_reg[205][29]/P0001 ,
		_w11945_,
		_w11966_,
		_w12614_
	);
	LUT3 #(
		.INIT('h80)
	) name2102 (
		\wishbone_bd_ram_mem3_reg[176][29]/P0001 ,
		_w11941_,
		_w11942_,
		_w12615_
	);
	LUT3 #(
		.INIT('h80)
	) name2103 (
		\wishbone_bd_ram_mem3_reg[23][29]/P0001 ,
		_w11935_,
		_w11975_,
		_w12616_
	);
	LUT3 #(
		.INIT('h80)
	) name2104 (
		\wishbone_bd_ram_mem3_reg[164][29]/P0001 ,
		_w11929_,
		_w11930_,
		_w12617_
	);
	LUT4 #(
		.INIT('h0001)
	) name2105 (
		_w12614_,
		_w12615_,
		_w12616_,
		_w12617_,
		_w12618_
	);
	LUT3 #(
		.INIT('h80)
	) name2106 (
		\wishbone_bd_ram_mem3_reg[18][29]/P0001 ,
		_w11935_,
		_w11963_,
		_w12619_
	);
	LUT3 #(
		.INIT('h80)
	) name2107 (
		\wishbone_bd_ram_mem3_reg[88][29]/P0001 ,
		_w11972_,
		_w11990_,
		_w12620_
	);
	LUT3 #(
		.INIT('h80)
	) name2108 (
		\wishbone_bd_ram_mem3_reg[219][29]/P0001 ,
		_w11936_,
		_w11984_,
		_w12621_
	);
	LUT3 #(
		.INIT('h80)
	) name2109 (
		\wishbone_bd_ram_mem3_reg[167][29]/P0001 ,
		_w11930_,
		_w11975_,
		_w12622_
	);
	LUT4 #(
		.INIT('h0001)
	) name2110 (
		_w12619_,
		_w12620_,
		_w12621_,
		_w12622_,
		_w12623_
	);
	LUT4 #(
		.INIT('h8000)
	) name2111 (
		_w12608_,
		_w12613_,
		_w12618_,
		_w12623_,
		_w12624_
	);
	LUT3 #(
		.INIT('h80)
	) name2112 (
		\wishbone_bd_ram_mem3_reg[236][29]/P0001 ,
		_w11954_,
		_w11982_,
		_w12625_
	);
	LUT3 #(
		.INIT('h80)
	) name2113 (
		\wishbone_bd_ram_mem3_reg[79][29]/P0001 ,
		_w11949_,
		_w11973_,
		_w12626_
	);
	LUT3 #(
		.INIT('h80)
	) name2114 (
		\wishbone_bd_ram_mem3_reg[140][29]/P0001 ,
		_w11954_,
		_w11955_,
		_w12627_
	);
	LUT3 #(
		.INIT('h80)
	) name2115 (
		\wishbone_bd_ram_mem3_reg[124][29]/P0001 ,
		_w11954_,
		_w12012_,
		_w12628_
	);
	LUT4 #(
		.INIT('h0001)
	) name2116 (
		_w12625_,
		_w12626_,
		_w12627_,
		_w12628_,
		_w12629_
	);
	LUT3 #(
		.INIT('h80)
	) name2117 (
		\wishbone_bd_ram_mem3_reg[177][29]/P0001 ,
		_w11942_,
		_w11977_,
		_w12630_
	);
	LUT3 #(
		.INIT('h80)
	) name2118 (
		\wishbone_bd_ram_mem3_reg[133][29]/P0001 ,
		_w11933_,
		_w11955_,
		_w12631_
	);
	LUT3 #(
		.INIT('h80)
	) name2119 (
		\wishbone_bd_ram_mem3_reg[218][29]/P0001 ,
		_w11944_,
		_w11984_,
		_w12632_
	);
	LUT3 #(
		.INIT('h80)
	) name2120 (
		\wishbone_bd_ram_mem3_reg[235][29]/P0001 ,
		_w11936_,
		_w11982_,
		_w12633_
	);
	LUT4 #(
		.INIT('h0001)
	) name2121 (
		_w12630_,
		_w12631_,
		_w12632_,
		_w12633_,
		_w12634_
	);
	LUT3 #(
		.INIT('h80)
	) name2122 (
		\wishbone_bd_ram_mem3_reg[5][29]/P0001 ,
		_w11932_,
		_w11933_,
		_w12635_
	);
	LUT3 #(
		.INIT('h80)
	) name2123 (
		\wishbone_bd_ram_mem3_reg[31][29]/P0001 ,
		_w11935_,
		_w11973_,
		_w12636_
	);
	LUT3 #(
		.INIT('h80)
	) name2124 (
		\wishbone_bd_ram_mem3_reg[30][29]/P0001 ,
		_w11935_,
		_w11948_,
		_w12637_
	);
	LUT3 #(
		.INIT('h80)
	) name2125 (
		\wishbone_bd_ram_mem3_reg[184][29]/P0001 ,
		_w11942_,
		_w11990_,
		_w12638_
	);
	LUT4 #(
		.INIT('h0001)
	) name2126 (
		_w12635_,
		_w12636_,
		_w12637_,
		_w12638_,
		_w12639_
	);
	LUT3 #(
		.INIT('h80)
	) name2127 (
		\wishbone_bd_ram_mem3_reg[245][29]/P0001 ,
		_w11933_,
		_w11952_,
		_w12640_
	);
	LUT3 #(
		.INIT('h80)
	) name2128 (
		\wishbone_bd_ram_mem3_reg[16][29]/P0001 ,
		_w11935_,
		_w11941_,
		_w12641_
	);
	LUT3 #(
		.INIT('h80)
	) name2129 (
		\wishbone_bd_ram_mem3_reg[227][29]/P0001 ,
		_w11938_,
		_w11982_,
		_w12642_
	);
	LUT3 #(
		.INIT('h80)
	) name2130 (
		\wishbone_bd_ram_mem3_reg[52][29]/P0001 ,
		_w11929_,
		_w11979_,
		_w12643_
	);
	LUT4 #(
		.INIT('h0001)
	) name2131 (
		_w12640_,
		_w12641_,
		_w12642_,
		_w12643_,
		_w12644_
	);
	LUT4 #(
		.INIT('h8000)
	) name2132 (
		_w12629_,
		_w12634_,
		_w12639_,
		_w12644_,
		_w12645_
	);
	LUT3 #(
		.INIT('h80)
	) name2133 (
		\wishbone_bd_ram_mem3_reg[153][29]/P0001 ,
		_w11959_,
		_w11968_,
		_w12646_
	);
	LUT3 #(
		.INIT('h80)
	) name2134 (
		\wishbone_bd_ram_mem3_reg[155][29]/P0001 ,
		_w11936_,
		_w11959_,
		_w12647_
	);
	LUT3 #(
		.INIT('h80)
	) name2135 (
		\wishbone_bd_ram_mem3_reg[96][29]/P0001 ,
		_w11941_,
		_w11965_,
		_w12648_
	);
	LUT3 #(
		.INIT('h80)
	) name2136 (
		\wishbone_bd_ram_mem3_reg[156][29]/P0001 ,
		_w11954_,
		_w11959_,
		_w12649_
	);
	LUT4 #(
		.INIT('h0001)
	) name2137 (
		_w12646_,
		_w12647_,
		_w12648_,
		_w12649_,
		_w12650_
	);
	LUT3 #(
		.INIT('h80)
	) name2138 (
		\wishbone_bd_ram_mem3_reg[217][29]/P0001 ,
		_w11968_,
		_w11984_,
		_w12651_
	);
	LUT3 #(
		.INIT('h80)
	) name2139 (
		\wishbone_bd_ram_mem3_reg[209][29]/P0001 ,
		_w11977_,
		_w11984_,
		_w12652_
	);
	LUT3 #(
		.INIT('h80)
	) name2140 (
		\wishbone_bd_ram_mem3_reg[150][29]/P0001 ,
		_w11959_,
		_w11986_,
		_w12653_
	);
	LUT3 #(
		.INIT('h80)
	) name2141 (
		\wishbone_bd_ram_mem3_reg[223][29]/P0001 ,
		_w11973_,
		_w11984_,
		_w12654_
	);
	LUT4 #(
		.INIT('h0001)
	) name2142 (
		_w12651_,
		_w12652_,
		_w12653_,
		_w12654_,
		_w12655_
	);
	LUT3 #(
		.INIT('h80)
	) name2143 (
		\wishbone_bd_ram_mem3_reg[55][29]/P0001 ,
		_w11975_,
		_w11979_,
		_w12656_
	);
	LUT3 #(
		.INIT('h80)
	) name2144 (
		\wishbone_bd_ram_mem3_reg[99][29]/P0001 ,
		_w11938_,
		_w11965_,
		_w12657_
	);
	LUT3 #(
		.INIT('h80)
	) name2145 (
		\wishbone_bd_ram_mem3_reg[234][29]/P0001 ,
		_w11944_,
		_w11982_,
		_w12658_
	);
	LUT3 #(
		.INIT('h80)
	) name2146 (
		\wishbone_bd_ram_mem3_reg[187][29]/P0001 ,
		_w11936_,
		_w11942_,
		_w12659_
	);
	LUT4 #(
		.INIT('h0001)
	) name2147 (
		_w12656_,
		_w12657_,
		_w12658_,
		_w12659_,
		_w12660_
	);
	LUT3 #(
		.INIT('h80)
	) name2148 (
		\wishbone_bd_ram_mem3_reg[92][29]/P0001 ,
		_w11954_,
		_w11972_,
		_w12661_
	);
	LUT3 #(
		.INIT('h80)
	) name2149 (
		\wishbone_bd_ram_mem3_reg[132][29]/P0001 ,
		_w11929_,
		_w11955_,
		_w12662_
	);
	LUT3 #(
		.INIT('h80)
	) name2150 (
		\wishbone_bd_ram_mem3_reg[37][29]/P0001 ,
		_w11933_,
		_w11957_,
		_w12663_
	);
	LUT3 #(
		.INIT('h80)
	) name2151 (
		\wishbone_bd_ram_mem3_reg[197][29]/P0001 ,
		_w11933_,
		_w11945_,
		_w12664_
	);
	LUT4 #(
		.INIT('h0001)
	) name2152 (
		_w12661_,
		_w12662_,
		_w12663_,
		_w12664_,
		_w12665_
	);
	LUT4 #(
		.INIT('h8000)
	) name2153 (
		_w12650_,
		_w12655_,
		_w12660_,
		_w12665_,
		_w12666_
	);
	LUT4 #(
		.INIT('h8000)
	) name2154 (
		_w12603_,
		_w12624_,
		_w12645_,
		_w12666_,
		_w12667_
	);
	LUT4 #(
		.INIT('h8000)
	) name2155 (
		_w12412_,
		_w12497_,
		_w12582_,
		_w12667_,
		_w12668_
	);
	LUT2 #(
		.INIT('h1)
	) name2156 (
		_w12302_,
		_w12304_,
		_w12669_
	);
	LUT3 #(
		.INIT('h10)
	) name2157 (
		\wishbone_TxLength_reg[12]/NET0131 ,
		_w12323_,
		_w12324_,
		_w12670_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2158 (
		\wishbone_TxLength_reg[13]/NET0131 ,
		_w12319_,
		_w12669_,
		_w12670_,
		_w12671_
	);
	LUT3 #(
		.INIT('h20)
	) name2159 (
		_w12315_,
		_w12323_,
		_w12324_,
		_w12672_
	);
	LUT2 #(
		.INIT('h8)
	) name2160 (
		_w12319_,
		_w12672_,
		_w12673_
	);
	LUT2 #(
		.INIT('h1)
	) name2161 (
		_w12671_,
		_w12673_,
		_w12674_
	);
	LUT3 #(
		.INIT('h2f)
	) name2162 (
		_w12303_,
		_w12668_,
		_w12674_,
		_w12675_
	);
	LUT3 #(
		.INIT('h80)
	) name2163 (
		\wishbone_bd_ram_mem3_reg[64][30]/P0001 ,
		_w11941_,
		_w11949_,
		_w12676_
	);
	LUT3 #(
		.INIT('h80)
	) name2164 (
		\wishbone_bd_ram_mem3_reg[211][30]/P0001 ,
		_w11938_,
		_w11984_,
		_w12677_
	);
	LUT3 #(
		.INIT('h80)
	) name2165 (
		\wishbone_bd_ram_mem3_reg[1][30]/P0001 ,
		_w11932_,
		_w11977_,
		_w12678_
	);
	LUT3 #(
		.INIT('h80)
	) name2166 (
		\wishbone_bd_ram_mem3_reg[10][30]/P0001 ,
		_w11932_,
		_w11944_,
		_w12679_
	);
	LUT4 #(
		.INIT('h0001)
	) name2167 (
		_w12676_,
		_w12677_,
		_w12678_,
		_w12679_,
		_w12680_
	);
	LUT3 #(
		.INIT('h80)
	) name2168 (
		\wishbone_bd_ram_mem3_reg[132][30]/P0001 ,
		_w11929_,
		_w11955_,
		_w12681_
	);
	LUT3 #(
		.INIT('h80)
	) name2169 (
		\wishbone_bd_ram_mem3_reg[237][30]/P0001 ,
		_w11966_,
		_w11982_,
		_w12682_
	);
	LUT3 #(
		.INIT('h80)
	) name2170 (
		\wishbone_bd_ram_mem3_reg[119][30]/P0001 ,
		_w11975_,
		_w12012_,
		_w12683_
	);
	LUT3 #(
		.INIT('h80)
	) name2171 (
		\wishbone_bd_ram_mem3_reg[242][30]/P0001 ,
		_w11952_,
		_w11963_,
		_w12684_
	);
	LUT4 #(
		.INIT('h0001)
	) name2172 (
		_w12681_,
		_w12682_,
		_w12683_,
		_w12684_,
		_w12685_
	);
	LUT3 #(
		.INIT('h80)
	) name2173 (
		\wishbone_bd_ram_mem3_reg[206][30]/P0001 ,
		_w11945_,
		_w11948_,
		_w12686_
	);
	LUT3 #(
		.INIT('h80)
	) name2174 (
		\wishbone_bd_ram_mem3_reg[175][30]/P0001 ,
		_w11930_,
		_w11973_,
		_w12687_
	);
	LUT3 #(
		.INIT('h80)
	) name2175 (
		\wishbone_bd_ram_mem3_reg[77][30]/P0001 ,
		_w11949_,
		_w11966_,
		_w12688_
	);
	LUT3 #(
		.INIT('h80)
	) name2176 (
		\wishbone_bd_ram_mem3_reg[232][30]/P0001 ,
		_w11982_,
		_w11990_,
		_w12689_
	);
	LUT4 #(
		.INIT('h0001)
	) name2177 (
		_w12686_,
		_w12687_,
		_w12688_,
		_w12689_,
		_w12690_
	);
	LUT3 #(
		.INIT('h80)
	) name2178 (
		\wishbone_bd_ram_mem3_reg[109][30]/P0001 ,
		_w11965_,
		_w11966_,
		_w12691_
	);
	LUT3 #(
		.INIT('h80)
	) name2179 (
		\wishbone_bd_ram_mem3_reg[181][30]/P0001 ,
		_w11933_,
		_w11942_,
		_w12692_
	);
	LUT3 #(
		.INIT('h80)
	) name2180 (
		\wishbone_bd_ram_mem3_reg[74][30]/P0001 ,
		_w11944_,
		_w11949_,
		_w12693_
	);
	LUT3 #(
		.INIT('h80)
	) name2181 (
		\wishbone_bd_ram_mem3_reg[192][30]/P0001 ,
		_w11941_,
		_w11945_,
		_w12694_
	);
	LUT4 #(
		.INIT('h0001)
	) name2182 (
		_w12691_,
		_w12692_,
		_w12693_,
		_w12694_,
		_w12695_
	);
	LUT4 #(
		.INIT('h8000)
	) name2183 (
		_w12680_,
		_w12685_,
		_w12690_,
		_w12695_,
		_w12696_
	);
	LUT3 #(
		.INIT('h80)
	) name2184 (
		\wishbone_bd_ram_mem3_reg[104][30]/P0001 ,
		_w11965_,
		_w11990_,
		_w12697_
	);
	LUT3 #(
		.INIT('h80)
	) name2185 (
		\wishbone_bd_ram_mem3_reg[102][30]/P0001 ,
		_w11965_,
		_w11986_,
		_w12698_
	);
	LUT3 #(
		.INIT('h80)
	) name2186 (
		\wishbone_bd_ram_mem3_reg[50][30]/P0001 ,
		_w11963_,
		_w11979_,
		_w12699_
	);
	LUT3 #(
		.INIT('h80)
	) name2187 (
		\wishbone_bd_ram_mem3_reg[163][30]/P0001 ,
		_w11930_,
		_w11938_,
		_w12700_
	);
	LUT4 #(
		.INIT('h0001)
	) name2188 (
		_w12697_,
		_w12698_,
		_w12699_,
		_w12700_,
		_w12701_
	);
	LUT3 #(
		.INIT('h80)
	) name2189 (
		\wishbone_bd_ram_mem3_reg[226][30]/P0001 ,
		_w11963_,
		_w11982_,
		_w12702_
	);
	LUT3 #(
		.INIT('h80)
	) name2190 (
		\wishbone_bd_ram_mem3_reg[199][30]/P0001 ,
		_w11945_,
		_w11975_,
		_w12703_
	);
	LUT3 #(
		.INIT('h80)
	) name2191 (
		\wishbone_bd_ram_mem3_reg[32][30]/P0001 ,
		_w11941_,
		_w11957_,
		_w12704_
	);
	LUT3 #(
		.INIT('h80)
	) name2192 (
		\wishbone_bd_ram_mem3_reg[67][30]/P0001 ,
		_w11938_,
		_w11949_,
		_w12705_
	);
	LUT4 #(
		.INIT('h0001)
	) name2193 (
		_w12702_,
		_w12703_,
		_w12704_,
		_w12705_,
		_w12706_
	);
	LUT3 #(
		.INIT('h80)
	) name2194 (
		\wishbone_bd_ram_mem3_reg[182][30]/P0001 ,
		_w11942_,
		_w11986_,
		_w12707_
	);
	LUT3 #(
		.INIT('h80)
	) name2195 (
		\wishbone_bd_ram_mem3_reg[227][30]/P0001 ,
		_w11938_,
		_w11982_,
		_w12708_
	);
	LUT3 #(
		.INIT('h80)
	) name2196 (
		\wishbone_bd_ram_mem3_reg[216][30]/P0001 ,
		_w11984_,
		_w11990_,
		_w12709_
	);
	LUT3 #(
		.INIT('h80)
	) name2197 (
		\wishbone_bd_ram_mem3_reg[43][30]/P0001 ,
		_w11936_,
		_w11957_,
		_w12710_
	);
	LUT4 #(
		.INIT('h0001)
	) name2198 (
		_w12707_,
		_w12708_,
		_w12709_,
		_w12710_,
		_w12711_
	);
	LUT3 #(
		.INIT('h80)
	) name2199 (
		\wishbone_bd_ram_mem3_reg[58][30]/P0001 ,
		_w11944_,
		_w11979_,
		_w12712_
	);
	LUT3 #(
		.INIT('h80)
	) name2200 (
		\wishbone_bd_ram_mem3_reg[205][30]/P0001 ,
		_w11945_,
		_w11966_,
		_w12713_
	);
	LUT3 #(
		.INIT('h80)
	) name2201 (
		\wishbone_bd_ram_mem3_reg[144][30]/P0001 ,
		_w11941_,
		_w11959_,
		_w12714_
	);
	LUT3 #(
		.INIT('h80)
	) name2202 (
		\wishbone_bd_ram_mem3_reg[215][30]/P0001 ,
		_w11975_,
		_w11984_,
		_w12715_
	);
	LUT4 #(
		.INIT('h0001)
	) name2203 (
		_w12712_,
		_w12713_,
		_w12714_,
		_w12715_,
		_w12716_
	);
	LUT4 #(
		.INIT('h8000)
	) name2204 (
		_w12701_,
		_w12706_,
		_w12711_,
		_w12716_,
		_w12717_
	);
	LUT3 #(
		.INIT('h80)
	) name2205 (
		\wishbone_bd_ram_mem3_reg[173][30]/P0001 ,
		_w11930_,
		_w11966_,
		_w12718_
	);
	LUT3 #(
		.INIT('h80)
	) name2206 (
		\wishbone_bd_ram_mem3_reg[123][30]/P0001 ,
		_w11936_,
		_w12012_,
		_w12719_
	);
	LUT3 #(
		.INIT('h80)
	) name2207 (
		\wishbone_bd_ram_mem3_reg[193][30]/P0001 ,
		_w11945_,
		_w11977_,
		_w12720_
	);
	LUT3 #(
		.INIT('h80)
	) name2208 (
		\wishbone_bd_ram_mem3_reg[3][30]/P0001 ,
		_w11932_,
		_w11938_,
		_w12721_
	);
	LUT4 #(
		.INIT('h0001)
	) name2209 (
		_w12718_,
		_w12719_,
		_w12720_,
		_w12721_,
		_w12722_
	);
	LUT3 #(
		.INIT('h80)
	) name2210 (
		\wishbone_bd_ram_mem3_reg[183][30]/P0001 ,
		_w11942_,
		_w11975_,
		_w12723_
	);
	LUT3 #(
		.INIT('h80)
	) name2211 (
		\wishbone_bd_ram_mem3_reg[131][30]/P0001 ,
		_w11938_,
		_w11955_,
		_w12724_
	);
	LUT3 #(
		.INIT('h80)
	) name2212 (
		\wishbone_bd_ram_mem3_reg[213][30]/P0001 ,
		_w11933_,
		_w11984_,
		_w12725_
	);
	LUT3 #(
		.INIT('h80)
	) name2213 (
		\wishbone_bd_ram_mem3_reg[156][30]/P0001 ,
		_w11954_,
		_w11959_,
		_w12726_
	);
	LUT4 #(
		.INIT('h0001)
	) name2214 (
		_w12723_,
		_w12724_,
		_w12725_,
		_w12726_,
		_w12727_
	);
	LUT3 #(
		.INIT('h80)
	) name2215 (
		\wishbone_bd_ram_mem3_reg[107][30]/P0001 ,
		_w11936_,
		_w11965_,
		_w12728_
	);
	LUT3 #(
		.INIT('h80)
	) name2216 (
		\wishbone_bd_ram_mem3_reg[73][30]/P0001 ,
		_w11949_,
		_w11968_,
		_w12729_
	);
	LUT3 #(
		.INIT('h80)
	) name2217 (
		\wishbone_bd_ram_mem3_reg[208][30]/P0001 ,
		_w11941_,
		_w11984_,
		_w12730_
	);
	LUT3 #(
		.INIT('h80)
	) name2218 (
		\wishbone_bd_ram_mem3_reg[241][30]/P0001 ,
		_w11952_,
		_w11977_,
		_w12731_
	);
	LUT4 #(
		.INIT('h0001)
	) name2219 (
		_w12728_,
		_w12729_,
		_w12730_,
		_w12731_,
		_w12732_
	);
	LUT3 #(
		.INIT('h80)
	) name2220 (
		\wishbone_bd_ram_mem3_reg[154][30]/P0001 ,
		_w11944_,
		_w11959_,
		_w12733_
	);
	LUT3 #(
		.INIT('h80)
	) name2221 (
		\wishbone_bd_ram_mem3_reg[252][30]/P0001 ,
		_w11952_,
		_w11954_,
		_w12734_
	);
	LUT3 #(
		.INIT('h80)
	) name2222 (
		\wishbone_bd_ram_mem3_reg[72][30]/P0001 ,
		_w11949_,
		_w11990_,
		_w12735_
	);
	LUT3 #(
		.INIT('h80)
	) name2223 (
		\wishbone_bd_ram_mem3_reg[229][30]/P0001 ,
		_w11933_,
		_w11982_,
		_w12736_
	);
	LUT4 #(
		.INIT('h0001)
	) name2224 (
		_w12733_,
		_w12734_,
		_w12735_,
		_w12736_,
		_w12737_
	);
	LUT4 #(
		.INIT('h8000)
	) name2225 (
		_w12722_,
		_w12727_,
		_w12732_,
		_w12737_,
		_w12738_
	);
	LUT3 #(
		.INIT('h80)
	) name2226 (
		\wishbone_bd_ram_mem3_reg[83][30]/P0001 ,
		_w11938_,
		_w11972_,
		_w12739_
	);
	LUT3 #(
		.INIT('h80)
	) name2227 (
		\wishbone_bd_ram_mem3_reg[130][30]/P0001 ,
		_w11955_,
		_w11963_,
		_w12740_
	);
	LUT3 #(
		.INIT('h80)
	) name2228 (
		\wishbone_bd_ram_mem3_reg[98][30]/P0001 ,
		_w11963_,
		_w11965_,
		_w12741_
	);
	LUT3 #(
		.INIT('h80)
	) name2229 (
		\wishbone_bd_ram_mem3_reg[146][30]/P0001 ,
		_w11959_,
		_w11963_,
		_w12742_
	);
	LUT4 #(
		.INIT('h0001)
	) name2230 (
		_w12739_,
		_w12740_,
		_w12741_,
		_w12742_,
		_w12743_
	);
	LUT3 #(
		.INIT('h80)
	) name2231 (
		\wishbone_bd_ram_mem3_reg[210][30]/P0001 ,
		_w11963_,
		_w11984_,
		_w12744_
	);
	LUT3 #(
		.INIT('h80)
	) name2232 (
		\wishbone_bd_ram_mem3_reg[180][30]/P0001 ,
		_w11929_,
		_w11942_,
		_w12745_
	);
	LUT3 #(
		.INIT('h80)
	) name2233 (
		\wishbone_bd_ram_mem3_reg[56][30]/P0001 ,
		_w11979_,
		_w11990_,
		_w12746_
	);
	LUT3 #(
		.INIT('h80)
	) name2234 (
		\wishbone_bd_ram_mem3_reg[27][30]/P0001 ,
		_w11935_,
		_w11936_,
		_w12747_
	);
	LUT4 #(
		.INIT('h0001)
	) name2235 (
		_w12744_,
		_w12745_,
		_w12746_,
		_w12747_,
		_w12748_
	);
	LUT3 #(
		.INIT('h80)
	) name2236 (
		\wishbone_bd_ram_mem3_reg[196][30]/P0001 ,
		_w11929_,
		_w11945_,
		_w12749_
	);
	LUT3 #(
		.INIT('h80)
	) name2237 (
		\wishbone_bd_ram_mem3_reg[61][30]/P0001 ,
		_w11966_,
		_w11979_,
		_w12750_
	);
	LUT3 #(
		.INIT('h80)
	) name2238 (
		\wishbone_bd_ram_mem3_reg[116][30]/P0001 ,
		_w11929_,
		_w12012_,
		_w12751_
	);
	LUT3 #(
		.INIT('h80)
	) name2239 (
		\wishbone_bd_ram_mem3_reg[148][30]/P0001 ,
		_w11929_,
		_w11959_,
		_w12752_
	);
	LUT4 #(
		.INIT('h0001)
	) name2240 (
		_w12749_,
		_w12750_,
		_w12751_,
		_w12752_,
		_w12753_
	);
	LUT3 #(
		.INIT('h80)
	) name2241 (
		\wishbone_bd_ram_mem3_reg[66][30]/P0001 ,
		_w11949_,
		_w11963_,
		_w12754_
	);
	LUT3 #(
		.INIT('h80)
	) name2242 (
		\wishbone_bd_ram_mem3_reg[15][30]/P0001 ,
		_w11932_,
		_w11973_,
		_w12755_
	);
	LUT3 #(
		.INIT('h80)
	) name2243 (
		\wishbone_bd_ram_mem3_reg[33][30]/P0001 ,
		_w11957_,
		_w11977_,
		_w12756_
	);
	LUT3 #(
		.INIT('h80)
	) name2244 (
		\wishbone_bd_ram_mem3_reg[174][30]/P0001 ,
		_w11930_,
		_w11948_,
		_w12757_
	);
	LUT4 #(
		.INIT('h0001)
	) name2245 (
		_w12754_,
		_w12755_,
		_w12756_,
		_w12757_,
		_w12758_
	);
	LUT4 #(
		.INIT('h8000)
	) name2246 (
		_w12743_,
		_w12748_,
		_w12753_,
		_w12758_,
		_w12759_
	);
	LUT4 #(
		.INIT('h8000)
	) name2247 (
		_w12696_,
		_w12717_,
		_w12738_,
		_w12759_,
		_w12760_
	);
	LUT3 #(
		.INIT('h80)
	) name2248 (
		\wishbone_bd_ram_mem3_reg[34][30]/P0001 ,
		_w11957_,
		_w11963_,
		_w12761_
	);
	LUT3 #(
		.INIT('h80)
	) name2249 (
		\wishbone_bd_ram_mem3_reg[169][30]/P0001 ,
		_w11930_,
		_w11968_,
		_w12762_
	);
	LUT3 #(
		.INIT('h80)
	) name2250 (
		\wishbone_bd_ram_mem3_reg[200][30]/P0001 ,
		_w11945_,
		_w11990_,
		_w12763_
	);
	LUT3 #(
		.INIT('h80)
	) name2251 (
		\wishbone_bd_ram_mem3_reg[230][30]/P0001 ,
		_w11982_,
		_w11986_,
		_w12764_
	);
	LUT4 #(
		.INIT('h0001)
	) name2252 (
		_w12761_,
		_w12762_,
		_w12763_,
		_w12764_,
		_w12765_
	);
	LUT3 #(
		.INIT('h80)
	) name2253 (
		\wishbone_bd_ram_mem3_reg[255][30]/P0001 ,
		_w11952_,
		_w11973_,
		_w12766_
	);
	LUT3 #(
		.INIT('h80)
	) name2254 (
		\wishbone_bd_ram_mem3_reg[87][30]/P0001 ,
		_w11972_,
		_w11975_,
		_w12767_
	);
	LUT3 #(
		.INIT('h80)
	) name2255 (
		\wishbone_bd_ram_mem3_reg[0][30]/P0001 ,
		_w11932_,
		_w11941_,
		_w12768_
	);
	LUT3 #(
		.INIT('h80)
	) name2256 (
		\wishbone_bd_ram_mem3_reg[18][30]/P0001 ,
		_w11935_,
		_w11963_,
		_w12769_
	);
	LUT4 #(
		.INIT('h0001)
	) name2257 (
		_w12766_,
		_w12767_,
		_w12768_,
		_w12769_,
		_w12770_
	);
	LUT3 #(
		.INIT('h80)
	) name2258 (
		\wishbone_bd_ram_mem3_reg[186][30]/P0001 ,
		_w11942_,
		_w11944_,
		_w12771_
	);
	LUT3 #(
		.INIT('h80)
	) name2259 (
		\wishbone_bd_ram_mem3_reg[136][30]/P0001 ,
		_w11955_,
		_w11990_,
		_w12772_
	);
	LUT3 #(
		.INIT('h80)
	) name2260 (
		\wishbone_bd_ram_mem3_reg[158][30]/P0001 ,
		_w11948_,
		_w11959_,
		_w12773_
	);
	LUT3 #(
		.INIT('h80)
	) name2261 (
		\wishbone_bd_ram_mem3_reg[212][30]/P0001 ,
		_w11929_,
		_w11984_,
		_w12774_
	);
	LUT4 #(
		.INIT('h0001)
	) name2262 (
		_w12771_,
		_w12772_,
		_w12773_,
		_w12774_,
		_w12775_
	);
	LUT3 #(
		.INIT('h80)
	) name2263 (
		\wishbone_bd_ram_mem3_reg[112][30]/P0001 ,
		_w11941_,
		_w12012_,
		_w12776_
	);
	LUT3 #(
		.INIT('h80)
	) name2264 (
		\wishbone_bd_ram_mem3_reg[86][30]/P0001 ,
		_w11972_,
		_w11986_,
		_w12777_
	);
	LUT3 #(
		.INIT('h80)
	) name2265 (
		\wishbone_bd_ram_mem3_reg[153][30]/P0001 ,
		_w11959_,
		_w11968_,
		_w12778_
	);
	LUT3 #(
		.INIT('h80)
	) name2266 (
		\wishbone_bd_ram_mem3_reg[234][30]/P0001 ,
		_w11944_,
		_w11982_,
		_w12779_
	);
	LUT4 #(
		.INIT('h0001)
	) name2267 (
		_w12776_,
		_w12777_,
		_w12778_,
		_w12779_,
		_w12780_
	);
	LUT4 #(
		.INIT('h8000)
	) name2268 (
		_w12765_,
		_w12770_,
		_w12775_,
		_w12780_,
		_w12781_
	);
	LUT3 #(
		.INIT('h80)
	) name2269 (
		\wishbone_bd_ram_mem3_reg[20][30]/P0001 ,
		_w11929_,
		_w11935_,
		_w12782_
	);
	LUT3 #(
		.INIT('h80)
	) name2270 (
		\wishbone_bd_ram_mem3_reg[224][30]/P0001 ,
		_w11941_,
		_w11982_,
		_w12783_
	);
	LUT3 #(
		.INIT('h80)
	) name2271 (
		\wishbone_bd_ram_mem3_reg[60][30]/P0001 ,
		_w11954_,
		_w11979_,
		_w12784_
	);
	LUT3 #(
		.INIT('h80)
	) name2272 (
		\wishbone_bd_ram_mem3_reg[36][30]/P0001 ,
		_w11929_,
		_w11957_,
		_w12785_
	);
	LUT4 #(
		.INIT('h0001)
	) name2273 (
		_w12782_,
		_w12783_,
		_w12784_,
		_w12785_,
		_w12786_
	);
	LUT3 #(
		.INIT('h80)
	) name2274 (
		\wishbone_bd_ram_mem3_reg[164][30]/P0001 ,
		_w11929_,
		_w11930_,
		_w12787_
	);
	LUT3 #(
		.INIT('h80)
	) name2275 (
		\wishbone_bd_ram_mem3_reg[135][30]/P0001 ,
		_w11955_,
		_w11975_,
		_w12788_
	);
	LUT3 #(
		.INIT('h80)
	) name2276 (
		\wishbone_bd_ram_mem3_reg[19][30]/P0001 ,
		_w11935_,
		_w11938_,
		_w12789_
	);
	LUT3 #(
		.INIT('h80)
	) name2277 (
		\wishbone_bd_ram_mem3_reg[103][30]/P0001 ,
		_w11965_,
		_w11975_,
		_w12790_
	);
	LUT4 #(
		.INIT('h0001)
	) name2278 (
		_w12787_,
		_w12788_,
		_w12789_,
		_w12790_,
		_w12791_
	);
	LUT3 #(
		.INIT('h80)
	) name2279 (
		\wishbone_bd_ram_mem3_reg[9][30]/P0001 ,
		_w11932_,
		_w11968_,
		_w12792_
	);
	LUT3 #(
		.INIT('h80)
	) name2280 (
		\wishbone_bd_ram_mem3_reg[97][30]/P0001 ,
		_w11965_,
		_w11977_,
		_w12793_
	);
	LUT3 #(
		.INIT('h80)
	) name2281 (
		\wishbone_bd_ram_mem3_reg[149][30]/P0001 ,
		_w11933_,
		_w11959_,
		_w12794_
	);
	LUT3 #(
		.INIT('h80)
	) name2282 (
		\wishbone_bd_ram_mem3_reg[28][30]/P0001 ,
		_w11935_,
		_w11954_,
		_w12795_
	);
	LUT4 #(
		.INIT('h0001)
	) name2283 (
		_w12792_,
		_w12793_,
		_w12794_,
		_w12795_,
		_w12796_
	);
	LUT3 #(
		.INIT('h80)
	) name2284 (
		\wishbone_bd_ram_mem3_reg[89][30]/P0001 ,
		_w11968_,
		_w11972_,
		_w12797_
	);
	LUT3 #(
		.INIT('h80)
	) name2285 (
		\wishbone_bd_ram_mem3_reg[250][30]/P0001 ,
		_w11944_,
		_w11952_,
		_w12798_
	);
	LUT3 #(
		.INIT('h80)
	) name2286 (
		\wishbone_bd_ram_mem3_reg[185][30]/P0001 ,
		_w11942_,
		_w11968_,
		_w12799_
	);
	LUT3 #(
		.INIT('h80)
	) name2287 (
		\wishbone_bd_ram_mem3_reg[100][30]/P0001 ,
		_w11929_,
		_w11965_,
		_w12800_
	);
	LUT4 #(
		.INIT('h0001)
	) name2288 (
		_w12797_,
		_w12798_,
		_w12799_,
		_w12800_,
		_w12801_
	);
	LUT4 #(
		.INIT('h8000)
	) name2289 (
		_w12786_,
		_w12791_,
		_w12796_,
		_w12801_,
		_w12802_
	);
	LUT3 #(
		.INIT('h80)
	) name2290 (
		\wishbone_bd_ram_mem3_reg[129][30]/P0001 ,
		_w11955_,
		_w11977_,
		_w12803_
	);
	LUT3 #(
		.INIT('h80)
	) name2291 (
		\wishbone_bd_ram_mem3_reg[91][30]/P0001 ,
		_w11936_,
		_w11972_,
		_w12804_
	);
	LUT3 #(
		.INIT('h80)
	) name2292 (
		\wishbone_bd_ram_mem3_reg[166][30]/P0001 ,
		_w11930_,
		_w11986_,
		_w12805_
	);
	LUT3 #(
		.INIT('h80)
	) name2293 (
		\wishbone_bd_ram_mem3_reg[204][30]/P0001 ,
		_w11945_,
		_w11954_,
		_w12806_
	);
	LUT4 #(
		.INIT('h0001)
	) name2294 (
		_w12803_,
		_w12804_,
		_w12805_,
		_w12806_,
		_w12807_
	);
	LUT3 #(
		.INIT('h80)
	) name2295 (
		\wishbone_bd_ram_mem3_reg[236][30]/P0001 ,
		_w11954_,
		_w11982_,
		_w12808_
	);
	LUT3 #(
		.INIT('h80)
	) name2296 (
		\wishbone_bd_ram_mem3_reg[187][30]/P0001 ,
		_w11936_,
		_w11942_,
		_w12809_
	);
	LUT3 #(
		.INIT('h80)
	) name2297 (
		\wishbone_bd_ram_mem3_reg[13][30]/P0001 ,
		_w11932_,
		_w11966_,
		_w12810_
	);
	LUT3 #(
		.INIT('h80)
	) name2298 (
		\wishbone_bd_ram_mem3_reg[26][30]/P0001 ,
		_w11935_,
		_w11944_,
		_w12811_
	);
	LUT4 #(
		.INIT('h0001)
	) name2299 (
		_w12808_,
		_w12809_,
		_w12810_,
		_w12811_,
		_w12812_
	);
	LUT3 #(
		.INIT('h80)
	) name2300 (
		\wishbone_bd_ram_mem3_reg[178][30]/P0001 ,
		_w11942_,
		_w11963_,
		_w12813_
	);
	LUT3 #(
		.INIT('h80)
	) name2301 (
		\wishbone_bd_ram_mem3_reg[157][30]/P0001 ,
		_w11959_,
		_w11966_,
		_w12814_
	);
	LUT3 #(
		.INIT('h80)
	) name2302 (
		\wishbone_bd_ram_mem3_reg[176][30]/P0001 ,
		_w11941_,
		_w11942_,
		_w12815_
	);
	LUT3 #(
		.INIT('h80)
	) name2303 (
		\wishbone_bd_ram_mem3_reg[235][30]/P0001 ,
		_w11936_,
		_w11982_,
		_w12816_
	);
	LUT4 #(
		.INIT('h0001)
	) name2304 (
		_w12813_,
		_w12814_,
		_w12815_,
		_w12816_,
		_w12817_
	);
	LUT3 #(
		.INIT('h80)
	) name2305 (
		\wishbone_bd_ram_mem3_reg[96][30]/P0001 ,
		_w11941_,
		_w11965_,
		_w12818_
	);
	LUT3 #(
		.INIT('h80)
	) name2306 (
		\wishbone_bd_ram_mem3_reg[190][30]/P0001 ,
		_w11942_,
		_w11948_,
		_w12819_
	);
	LUT3 #(
		.INIT('h80)
	) name2307 (
		\wishbone_bd_ram_mem3_reg[92][30]/P0001 ,
		_w11954_,
		_w11972_,
		_w12820_
	);
	LUT3 #(
		.INIT('h80)
	) name2308 (
		\wishbone_bd_ram_mem3_reg[117][30]/P0001 ,
		_w11933_,
		_w12012_,
		_w12821_
	);
	LUT4 #(
		.INIT('h0001)
	) name2309 (
		_w12818_,
		_w12819_,
		_w12820_,
		_w12821_,
		_w12822_
	);
	LUT4 #(
		.INIT('h8000)
	) name2310 (
		_w12807_,
		_w12812_,
		_w12817_,
		_w12822_,
		_w12823_
	);
	LUT3 #(
		.INIT('h80)
	) name2311 (
		\wishbone_bd_ram_mem3_reg[47][30]/P0001 ,
		_w11957_,
		_w11973_,
		_w12824_
	);
	LUT3 #(
		.INIT('h80)
	) name2312 (
		\wishbone_bd_ram_mem3_reg[54][30]/P0001 ,
		_w11979_,
		_w11986_,
		_w12825_
	);
	LUT3 #(
		.INIT('h80)
	) name2313 (
		\wishbone_bd_ram_mem3_reg[139][30]/P0001 ,
		_w11936_,
		_w11955_,
		_w12826_
	);
	LUT3 #(
		.INIT('h80)
	) name2314 (
		\wishbone_bd_ram_mem3_reg[239][30]/P0001 ,
		_w11973_,
		_w11982_,
		_w12827_
	);
	LUT4 #(
		.INIT('h0001)
	) name2315 (
		_w12824_,
		_w12825_,
		_w12826_,
		_w12827_,
		_w12828_
	);
	LUT3 #(
		.INIT('h80)
	) name2316 (
		\wishbone_bd_ram_mem3_reg[59][30]/P0001 ,
		_w11936_,
		_w11979_,
		_w12829_
	);
	LUT3 #(
		.INIT('h80)
	) name2317 (
		\wishbone_bd_ram_mem3_reg[134][30]/P0001 ,
		_w11955_,
		_w11986_,
		_w12830_
	);
	LUT3 #(
		.INIT('h80)
	) name2318 (
		\wishbone_bd_ram_mem3_reg[23][30]/P0001 ,
		_w11935_,
		_w11975_,
		_w12831_
	);
	LUT3 #(
		.INIT('h80)
	) name2319 (
		\wishbone_bd_ram_mem3_reg[142][30]/P0001 ,
		_w11948_,
		_w11955_,
		_w12832_
	);
	LUT4 #(
		.INIT('h0001)
	) name2320 (
		_w12829_,
		_w12830_,
		_w12831_,
		_w12832_,
		_w12833_
	);
	LUT3 #(
		.INIT('h80)
	) name2321 (
		\wishbone_bd_ram_mem3_reg[179][30]/P0001 ,
		_w11938_,
		_w11942_,
		_w12834_
	);
	LUT3 #(
		.INIT('h80)
	) name2322 (
		\wishbone_bd_ram_mem3_reg[53][30]/P0001 ,
		_w11933_,
		_w11979_,
		_w12835_
	);
	LUT3 #(
		.INIT('h80)
	) name2323 (
		\wishbone_bd_ram_mem3_reg[6][30]/P0001 ,
		_w11932_,
		_w11986_,
		_w12836_
	);
	LUT3 #(
		.INIT('h80)
	) name2324 (
		\wishbone_bd_ram_mem3_reg[254][30]/P0001 ,
		_w11948_,
		_w11952_,
		_w12837_
	);
	LUT4 #(
		.INIT('h0001)
	) name2325 (
		_w12834_,
		_w12835_,
		_w12836_,
		_w12837_,
		_w12838_
	);
	LUT3 #(
		.INIT('h80)
	) name2326 (
		\wishbone_bd_ram_mem3_reg[243][30]/P0001 ,
		_w11938_,
		_w11952_,
		_w12839_
	);
	LUT3 #(
		.INIT('h80)
	) name2327 (
		\wishbone_bd_ram_mem3_reg[219][30]/P0001 ,
		_w11936_,
		_w11984_,
		_w12840_
	);
	LUT3 #(
		.INIT('h80)
	) name2328 (
		\wishbone_bd_ram_mem3_reg[189][30]/P0001 ,
		_w11942_,
		_w11966_,
		_w12841_
	);
	LUT3 #(
		.INIT('h80)
	) name2329 (
		\wishbone_bd_ram_mem3_reg[141][30]/P0001 ,
		_w11955_,
		_w11966_,
		_w12842_
	);
	LUT4 #(
		.INIT('h0001)
	) name2330 (
		_w12839_,
		_w12840_,
		_w12841_,
		_w12842_,
		_w12843_
	);
	LUT4 #(
		.INIT('h8000)
	) name2331 (
		_w12828_,
		_w12833_,
		_w12838_,
		_w12843_,
		_w12844_
	);
	LUT4 #(
		.INIT('h8000)
	) name2332 (
		_w12781_,
		_w12802_,
		_w12823_,
		_w12844_,
		_w12845_
	);
	LUT3 #(
		.INIT('h80)
	) name2333 (
		\wishbone_bd_ram_mem3_reg[42][30]/P0001 ,
		_w11944_,
		_w11957_,
		_w12846_
	);
	LUT3 #(
		.INIT('h80)
	) name2334 (
		\wishbone_bd_ram_mem3_reg[128][30]/P0001 ,
		_w11941_,
		_w11955_,
		_w12847_
	);
	LUT3 #(
		.INIT('h80)
	) name2335 (
		\wishbone_bd_ram_mem3_reg[137][30]/P0001 ,
		_w11955_,
		_w11968_,
		_w12848_
	);
	LUT3 #(
		.INIT('h80)
	) name2336 (
		\wishbone_bd_ram_mem3_reg[251][30]/P0001 ,
		_w11936_,
		_w11952_,
		_w12849_
	);
	LUT4 #(
		.INIT('h0001)
	) name2337 (
		_w12846_,
		_w12847_,
		_w12848_,
		_w12849_,
		_w12850_
	);
	LUT3 #(
		.INIT('h80)
	) name2338 (
		\wishbone_bd_ram_mem3_reg[85][30]/P0001 ,
		_w11933_,
		_w11972_,
		_w12851_
	);
	LUT3 #(
		.INIT('h80)
	) name2339 (
		\wishbone_bd_ram_mem3_reg[2][30]/P0001 ,
		_w11932_,
		_w11963_,
		_w12852_
	);
	LUT3 #(
		.INIT('h80)
	) name2340 (
		\wishbone_bd_ram_mem3_reg[238][30]/P0001 ,
		_w11948_,
		_w11982_,
		_w12853_
	);
	LUT3 #(
		.INIT('h80)
	) name2341 (
		\wishbone_bd_ram_mem3_reg[218][30]/P0001 ,
		_w11944_,
		_w11984_,
		_w12854_
	);
	LUT4 #(
		.INIT('h0001)
	) name2342 (
		_w12851_,
		_w12852_,
		_w12853_,
		_w12854_,
		_w12855_
	);
	LUT3 #(
		.INIT('h80)
	) name2343 (
		\wishbone_bd_ram_mem3_reg[108][30]/P0001 ,
		_w11954_,
		_w11965_,
		_w12856_
	);
	LUT3 #(
		.INIT('h80)
	) name2344 (
		\wishbone_bd_ram_mem3_reg[21][30]/P0001 ,
		_w11933_,
		_w11935_,
		_w12857_
	);
	LUT3 #(
		.INIT('h80)
	) name2345 (
		\wishbone_bd_ram_mem3_reg[114][30]/P0001 ,
		_w11963_,
		_w12012_,
		_w12858_
	);
	LUT3 #(
		.INIT('h80)
	) name2346 (
		\wishbone_bd_ram_mem3_reg[155][30]/P0001 ,
		_w11936_,
		_w11959_,
		_w12859_
	);
	LUT4 #(
		.INIT('h0001)
	) name2347 (
		_w12856_,
		_w12857_,
		_w12858_,
		_w12859_,
		_w12860_
	);
	LUT3 #(
		.INIT('h80)
	) name2348 (
		\wishbone_bd_ram_mem3_reg[80][30]/P0001 ,
		_w11941_,
		_w11972_,
		_w12861_
	);
	LUT3 #(
		.INIT('h80)
	) name2349 (
		\wishbone_bd_ram_mem3_reg[231][30]/P0001 ,
		_w11975_,
		_w11982_,
		_w12862_
	);
	LUT3 #(
		.INIT('h80)
	) name2350 (
		\wishbone_bd_ram_mem3_reg[198][30]/P0001 ,
		_w11945_,
		_w11986_,
		_w12863_
	);
	LUT3 #(
		.INIT('h80)
	) name2351 (
		\wishbone_bd_ram_mem3_reg[25][30]/P0001 ,
		_w11935_,
		_w11968_,
		_w12864_
	);
	LUT4 #(
		.INIT('h0001)
	) name2352 (
		_w12861_,
		_w12862_,
		_w12863_,
		_w12864_,
		_w12865_
	);
	LUT4 #(
		.INIT('h8000)
	) name2353 (
		_w12850_,
		_w12855_,
		_w12860_,
		_w12865_,
		_w12866_
	);
	LUT3 #(
		.INIT('h80)
	) name2354 (
		\wishbone_bd_ram_mem3_reg[245][30]/P0001 ,
		_w11933_,
		_w11952_,
		_w12867_
	);
	LUT3 #(
		.INIT('h80)
	) name2355 (
		\wishbone_bd_ram_mem3_reg[17][30]/P0001 ,
		_w11935_,
		_w11977_,
		_w12868_
	);
	LUT3 #(
		.INIT('h80)
	) name2356 (
		\wishbone_bd_ram_mem3_reg[69][30]/P0001 ,
		_w11933_,
		_w11949_,
		_w12869_
	);
	LUT3 #(
		.INIT('h80)
	) name2357 (
		\wishbone_bd_ram_mem3_reg[160][30]/P0001 ,
		_w11930_,
		_w11941_,
		_w12870_
	);
	LUT4 #(
		.INIT('h0001)
	) name2358 (
		_w12867_,
		_w12868_,
		_w12869_,
		_w12870_,
		_w12871_
	);
	LUT3 #(
		.INIT('h80)
	) name2359 (
		\wishbone_bd_ram_mem3_reg[201][30]/P0001 ,
		_w11945_,
		_w11968_,
		_w12872_
	);
	LUT3 #(
		.INIT('h80)
	) name2360 (
		\wishbone_bd_ram_mem3_reg[167][30]/P0001 ,
		_w11930_,
		_w11975_,
		_w12873_
	);
	LUT3 #(
		.INIT('h80)
	) name2361 (
		\wishbone_bd_ram_mem3_reg[105][30]/P0001 ,
		_w11965_,
		_w11968_,
		_w12874_
	);
	LUT3 #(
		.INIT('h80)
	) name2362 (
		\wishbone_bd_ram_mem3_reg[111][30]/P0001 ,
		_w11965_,
		_w11973_,
		_w12875_
	);
	LUT4 #(
		.INIT('h0001)
	) name2363 (
		_w12872_,
		_w12873_,
		_w12874_,
		_w12875_,
		_w12876_
	);
	LUT3 #(
		.INIT('h80)
	) name2364 (
		\wishbone_bd_ram_mem3_reg[223][30]/P0001 ,
		_w11973_,
		_w11984_,
		_w12877_
	);
	LUT3 #(
		.INIT('h80)
	) name2365 (
		\wishbone_bd_ram_mem3_reg[30][30]/P0001 ,
		_w11935_,
		_w11948_,
		_w12878_
	);
	LUT3 #(
		.INIT('h80)
	) name2366 (
		\wishbone_bd_ram_mem3_reg[165][30]/P0001 ,
		_w11930_,
		_w11933_,
		_w12879_
	);
	LUT3 #(
		.INIT('h80)
	) name2367 (
		\wishbone_bd_ram_mem3_reg[70][30]/P0001 ,
		_w11949_,
		_w11986_,
		_w12880_
	);
	LUT4 #(
		.INIT('h0001)
	) name2368 (
		_w12877_,
		_w12878_,
		_w12879_,
		_w12880_,
		_w12881_
	);
	LUT3 #(
		.INIT('h80)
	) name2369 (
		\wishbone_bd_ram_mem3_reg[51][30]/P0001 ,
		_w11938_,
		_w11979_,
		_w12882_
	);
	LUT3 #(
		.INIT('h80)
	) name2370 (
		\wishbone_bd_ram_mem3_reg[81][30]/P0001 ,
		_w11972_,
		_w11977_,
		_w12883_
	);
	LUT3 #(
		.INIT('h80)
	) name2371 (
		\wishbone_bd_ram_mem3_reg[76][30]/P0001 ,
		_w11949_,
		_w11954_,
		_w12884_
	);
	LUT3 #(
		.INIT('h80)
	) name2372 (
		\wishbone_bd_ram_mem3_reg[159][30]/P0001 ,
		_w11959_,
		_w11973_,
		_w12885_
	);
	LUT4 #(
		.INIT('h0001)
	) name2373 (
		_w12882_,
		_w12883_,
		_w12884_,
		_w12885_,
		_w12886_
	);
	LUT4 #(
		.INIT('h8000)
	) name2374 (
		_w12871_,
		_w12876_,
		_w12881_,
		_w12886_,
		_w12887_
	);
	LUT3 #(
		.INIT('h80)
	) name2375 (
		\wishbone_bd_ram_mem3_reg[214][30]/P0001 ,
		_w11984_,
		_w11986_,
		_w12888_
	);
	LUT3 #(
		.INIT('h80)
	) name2376 (
		\wishbone_bd_ram_mem3_reg[172][30]/P0001 ,
		_w11930_,
		_w11954_,
		_w12889_
	);
	LUT3 #(
		.INIT('h80)
	) name2377 (
		\wishbone_bd_ram_mem3_reg[24][30]/P0001 ,
		_w11935_,
		_w11990_,
		_w12890_
	);
	LUT3 #(
		.INIT('h80)
	) name2378 (
		\wishbone_bd_ram_mem3_reg[170][30]/P0001 ,
		_w11930_,
		_w11944_,
		_w12891_
	);
	LUT4 #(
		.INIT('h0001)
	) name2379 (
		_w12888_,
		_w12889_,
		_w12890_,
		_w12891_,
		_w12892_
	);
	LUT3 #(
		.INIT('h80)
	) name2380 (
		\wishbone_bd_ram_mem3_reg[240][30]/P0001 ,
		_w11941_,
		_w11952_,
		_w12893_
	);
	LUT3 #(
		.INIT('h80)
	) name2381 (
		\wishbone_bd_ram_mem3_reg[151][30]/P0001 ,
		_w11959_,
		_w11975_,
		_w12894_
	);
	LUT3 #(
		.INIT('h80)
	) name2382 (
		\wishbone_bd_ram_mem3_reg[195][30]/P0001 ,
		_w11938_,
		_w11945_,
		_w12895_
	);
	LUT3 #(
		.INIT('h80)
	) name2383 (
		\wishbone_bd_ram_mem3_reg[46][30]/P0001 ,
		_w11948_,
		_w11957_,
		_w12896_
	);
	LUT4 #(
		.INIT('h0001)
	) name2384 (
		_w12893_,
		_w12894_,
		_w12895_,
		_w12896_,
		_w12897_
	);
	LUT3 #(
		.INIT('h80)
	) name2385 (
		\wishbone_bd_ram_mem3_reg[44][30]/P0001 ,
		_w11954_,
		_w11957_,
		_w12898_
	);
	LUT3 #(
		.INIT('h80)
	) name2386 (
		\wishbone_bd_ram_mem3_reg[133][30]/P0001 ,
		_w11933_,
		_w11955_,
		_w12899_
	);
	LUT3 #(
		.INIT('h80)
	) name2387 (
		\wishbone_bd_ram_mem3_reg[57][30]/P0001 ,
		_w11968_,
		_w11979_,
		_w12900_
	);
	LUT3 #(
		.INIT('h80)
	) name2388 (
		\wishbone_bd_ram_mem3_reg[106][30]/P0001 ,
		_w11944_,
		_w11965_,
		_w12901_
	);
	LUT4 #(
		.INIT('h0001)
	) name2389 (
		_w12898_,
		_w12899_,
		_w12900_,
		_w12901_,
		_w12902_
	);
	LUT3 #(
		.INIT('h80)
	) name2390 (
		\wishbone_bd_ram_mem3_reg[161][30]/P0001 ,
		_w11930_,
		_w11977_,
		_w12903_
	);
	LUT3 #(
		.INIT('h80)
	) name2391 (
		\wishbone_bd_ram_mem3_reg[99][30]/P0001 ,
		_w11938_,
		_w11965_,
		_w12904_
	);
	LUT3 #(
		.INIT('h80)
	) name2392 (
		\wishbone_bd_ram_mem3_reg[101][30]/P0001 ,
		_w11933_,
		_w11965_,
		_w12905_
	);
	LUT3 #(
		.INIT('h80)
	) name2393 (
		\wishbone_bd_ram_mem3_reg[233][30]/P0001 ,
		_w11968_,
		_w11982_,
		_w12906_
	);
	LUT4 #(
		.INIT('h0001)
	) name2394 (
		_w12903_,
		_w12904_,
		_w12905_,
		_w12906_,
		_w12907_
	);
	LUT4 #(
		.INIT('h8000)
	) name2395 (
		_w12892_,
		_w12897_,
		_w12902_,
		_w12907_,
		_w12908_
	);
	LUT3 #(
		.INIT('h80)
	) name2396 (
		\wishbone_bd_ram_mem3_reg[113][30]/P0001 ,
		_w11977_,
		_w12012_,
		_w12909_
	);
	LUT3 #(
		.INIT('h80)
	) name2397 (
		\wishbone_bd_ram_mem3_reg[197][30]/P0001 ,
		_w11933_,
		_w11945_,
		_w12910_
	);
	LUT3 #(
		.INIT('h80)
	) name2398 (
		\wishbone_bd_ram_mem3_reg[152][30]/P0001 ,
		_w11959_,
		_w11990_,
		_w12911_
	);
	LUT3 #(
		.INIT('h80)
	) name2399 (
		\wishbone_bd_ram_mem3_reg[22][30]/P0001 ,
		_w11935_,
		_w11986_,
		_w12912_
	);
	LUT4 #(
		.INIT('h0001)
	) name2400 (
		_w12909_,
		_w12910_,
		_w12911_,
		_w12912_,
		_w12913_
	);
	LUT3 #(
		.INIT('h80)
	) name2401 (
		\wishbone_bd_ram_mem3_reg[84][30]/P0001 ,
		_w11929_,
		_w11972_,
		_w12914_
	);
	LUT3 #(
		.INIT('h80)
	) name2402 (
		\wishbone_bd_ram_mem3_reg[244][30]/P0001 ,
		_w11929_,
		_w11952_,
		_w12915_
	);
	LUT3 #(
		.INIT('h80)
	) name2403 (
		\wishbone_bd_ram_mem3_reg[221][30]/P0001 ,
		_w11966_,
		_w11984_,
		_w12916_
	);
	LUT3 #(
		.INIT('h80)
	) name2404 (
		\wishbone_bd_ram_mem3_reg[203][30]/P0001 ,
		_w11936_,
		_w11945_,
		_w12917_
	);
	LUT4 #(
		.INIT('h0001)
	) name2405 (
		_w12914_,
		_w12915_,
		_w12916_,
		_w12917_,
		_w12918_
	);
	LUT3 #(
		.INIT('h80)
	) name2406 (
		\wishbone_bd_ram_mem3_reg[253][30]/P0001 ,
		_w11952_,
		_w11966_,
		_w12919_
	);
	LUT3 #(
		.INIT('h80)
	) name2407 (
		\wishbone_bd_ram_mem3_reg[79][30]/P0001 ,
		_w11949_,
		_w11973_,
		_w12920_
	);
	LUT3 #(
		.INIT('h80)
	) name2408 (
		\wishbone_bd_ram_mem3_reg[55][30]/P0001 ,
		_w11975_,
		_w11979_,
		_w12921_
	);
	LUT3 #(
		.INIT('h80)
	) name2409 (
		\wishbone_bd_ram_mem3_reg[222][30]/P0001 ,
		_w11948_,
		_w11984_,
		_w12922_
	);
	LUT4 #(
		.INIT('h0001)
	) name2410 (
		_w12919_,
		_w12920_,
		_w12921_,
		_w12922_,
		_w12923_
	);
	LUT3 #(
		.INIT('h80)
	) name2411 (
		\wishbone_bd_ram_mem3_reg[48][30]/P0001 ,
		_w11941_,
		_w11979_,
		_w12924_
	);
	LUT3 #(
		.INIT('h80)
	) name2412 (
		\wishbone_bd_ram_mem3_reg[52][30]/P0001 ,
		_w11929_,
		_w11979_,
		_w12925_
	);
	LUT3 #(
		.INIT('h80)
	) name2413 (
		\wishbone_bd_ram_mem3_reg[5][30]/P0001 ,
		_w11932_,
		_w11933_,
		_w12926_
	);
	LUT3 #(
		.INIT('h80)
	) name2414 (
		\wishbone_bd_ram_mem3_reg[78][30]/P0001 ,
		_w11948_,
		_w11949_,
		_w12927_
	);
	LUT4 #(
		.INIT('h0001)
	) name2415 (
		_w12924_,
		_w12925_,
		_w12926_,
		_w12927_,
		_w12928_
	);
	LUT4 #(
		.INIT('h8000)
	) name2416 (
		_w12913_,
		_w12918_,
		_w12923_,
		_w12928_,
		_w12929_
	);
	LUT4 #(
		.INIT('h8000)
	) name2417 (
		_w12866_,
		_w12887_,
		_w12908_,
		_w12929_,
		_w12930_
	);
	LUT3 #(
		.INIT('h80)
	) name2418 (
		\wishbone_bd_ram_mem3_reg[29][30]/P0001 ,
		_w11935_,
		_w11966_,
		_w12931_
	);
	LUT3 #(
		.INIT('h80)
	) name2419 (
		\wishbone_bd_ram_mem3_reg[184][30]/P0001 ,
		_w11942_,
		_w11990_,
		_w12932_
	);
	LUT3 #(
		.INIT('h80)
	) name2420 (
		\wishbone_bd_ram_mem3_reg[82][30]/P0001 ,
		_w11963_,
		_w11972_,
		_w12933_
	);
	LUT3 #(
		.INIT('h80)
	) name2421 (
		\wishbone_bd_ram_mem3_reg[63][30]/P0001 ,
		_w11973_,
		_w11979_,
		_w12934_
	);
	LUT4 #(
		.INIT('h0001)
	) name2422 (
		_w12931_,
		_w12932_,
		_w12933_,
		_w12934_,
		_w12935_
	);
	LUT3 #(
		.INIT('h80)
	) name2423 (
		\wishbone_bd_ram_mem3_reg[143][30]/P0001 ,
		_w11955_,
		_w11973_,
		_w12936_
	);
	LUT3 #(
		.INIT('h80)
	) name2424 (
		\wishbone_bd_ram_mem3_reg[75][30]/P0001 ,
		_w11936_,
		_w11949_,
		_w12937_
	);
	LUT3 #(
		.INIT('h80)
	) name2425 (
		\wishbone_bd_ram_mem3_reg[118][30]/P0001 ,
		_w11986_,
		_w12012_,
		_w12938_
	);
	LUT3 #(
		.INIT('h80)
	) name2426 (
		\wishbone_bd_ram_mem3_reg[194][30]/P0001 ,
		_w11945_,
		_w11963_,
		_w12939_
	);
	LUT4 #(
		.INIT('h0001)
	) name2427 (
		_w12936_,
		_w12937_,
		_w12938_,
		_w12939_,
		_w12940_
	);
	LUT3 #(
		.INIT('h80)
	) name2428 (
		\wishbone_bd_ram_mem3_reg[45][30]/P0001 ,
		_w11957_,
		_w11966_,
		_w12941_
	);
	LUT3 #(
		.INIT('h80)
	) name2429 (
		\wishbone_bd_ram_mem3_reg[225][30]/P0001 ,
		_w11977_,
		_w11982_,
		_w12942_
	);
	LUT3 #(
		.INIT('h80)
	) name2430 (
		\wishbone_bd_ram_mem3_reg[35][30]/P0001 ,
		_w11938_,
		_w11957_,
		_w12943_
	);
	LUT3 #(
		.INIT('h80)
	) name2431 (
		\wishbone_bd_ram_mem3_reg[127][30]/P0001 ,
		_w11973_,
		_w12012_,
		_w12944_
	);
	LUT4 #(
		.INIT('h0001)
	) name2432 (
		_w12941_,
		_w12942_,
		_w12943_,
		_w12944_,
		_w12945_
	);
	LUT3 #(
		.INIT('h80)
	) name2433 (
		\wishbone_bd_ram_mem3_reg[115][30]/P0001 ,
		_w11938_,
		_w12012_,
		_w12946_
	);
	LUT3 #(
		.INIT('h80)
	) name2434 (
		\wishbone_bd_ram_mem3_reg[37][30]/P0001 ,
		_w11933_,
		_w11957_,
		_w12947_
	);
	LUT3 #(
		.INIT('h80)
	) name2435 (
		\wishbone_bd_ram_mem3_reg[7][30]/P0001 ,
		_w11932_,
		_w11975_,
		_w12948_
	);
	LUT3 #(
		.INIT('h80)
	) name2436 (
		\wishbone_bd_ram_mem3_reg[68][30]/P0001 ,
		_w11929_,
		_w11949_,
		_w12949_
	);
	LUT4 #(
		.INIT('h0001)
	) name2437 (
		_w12946_,
		_w12947_,
		_w12948_,
		_w12949_,
		_w12950_
	);
	LUT4 #(
		.INIT('h8000)
	) name2438 (
		_w12935_,
		_w12940_,
		_w12945_,
		_w12950_,
		_w12951_
	);
	LUT3 #(
		.INIT('h80)
	) name2439 (
		\wishbone_bd_ram_mem3_reg[121][30]/P0001 ,
		_w11968_,
		_w12012_,
		_w12952_
	);
	LUT3 #(
		.INIT('h80)
	) name2440 (
		\wishbone_bd_ram_mem3_reg[11][30]/P0001 ,
		_w11932_,
		_w11936_,
		_w12953_
	);
	LUT3 #(
		.INIT('h80)
	) name2441 (
		\wishbone_bd_ram_mem3_reg[49][30]/P0001 ,
		_w11977_,
		_w11979_,
		_w12954_
	);
	LUT3 #(
		.INIT('h80)
	) name2442 (
		\wishbone_bd_ram_mem3_reg[145][30]/P0001 ,
		_w11959_,
		_w11977_,
		_w12955_
	);
	LUT4 #(
		.INIT('h0001)
	) name2443 (
		_w12952_,
		_w12953_,
		_w12954_,
		_w12955_,
		_w12956_
	);
	LUT3 #(
		.INIT('h80)
	) name2444 (
		\wishbone_bd_ram_mem3_reg[125][30]/P0001 ,
		_w11966_,
		_w12012_,
		_w12957_
	);
	LUT3 #(
		.INIT('h80)
	) name2445 (
		\wishbone_bd_ram_mem3_reg[122][30]/P0001 ,
		_w11944_,
		_w12012_,
		_w12958_
	);
	LUT3 #(
		.INIT('h80)
	) name2446 (
		\wishbone_bd_ram_mem3_reg[147][30]/P0001 ,
		_w11938_,
		_w11959_,
		_w12959_
	);
	LUT3 #(
		.INIT('h80)
	) name2447 (
		\wishbone_bd_ram_mem3_reg[31][30]/P0001 ,
		_w11935_,
		_w11973_,
		_w12960_
	);
	LUT4 #(
		.INIT('h0001)
	) name2448 (
		_w12957_,
		_w12958_,
		_w12959_,
		_w12960_,
		_w12961_
	);
	LUT3 #(
		.INIT('h80)
	) name2449 (
		\wishbone_bd_ram_mem3_reg[220][30]/P0001 ,
		_w11954_,
		_w11984_,
		_w12962_
	);
	LUT3 #(
		.INIT('h80)
	) name2450 (
		\wishbone_bd_ram_mem3_reg[188][30]/P0001 ,
		_w11942_,
		_w11954_,
		_w12963_
	);
	LUT3 #(
		.INIT('h80)
	) name2451 (
		\wishbone_bd_ram_mem3_reg[12][30]/P0001 ,
		_w11932_,
		_w11954_,
		_w12964_
	);
	LUT3 #(
		.INIT('h80)
	) name2452 (
		\wishbone_bd_ram_mem3_reg[38][30]/P0001 ,
		_w11957_,
		_w11986_,
		_w12965_
	);
	LUT4 #(
		.INIT('h0001)
	) name2453 (
		_w12962_,
		_w12963_,
		_w12964_,
		_w12965_,
		_w12966_
	);
	LUT3 #(
		.INIT('h80)
	) name2454 (
		\wishbone_bd_ram_mem3_reg[8][30]/P0001 ,
		_w11932_,
		_w11990_,
		_w12967_
	);
	LUT3 #(
		.INIT('h80)
	) name2455 (
		\wishbone_bd_ram_mem3_reg[39][30]/P0001 ,
		_w11957_,
		_w11975_,
		_w12968_
	);
	LUT3 #(
		.INIT('h80)
	) name2456 (
		\wishbone_bd_ram_mem3_reg[246][30]/P0001 ,
		_w11952_,
		_w11986_,
		_w12969_
	);
	LUT3 #(
		.INIT('h80)
	) name2457 (
		\wishbone_bd_ram_mem3_reg[138][30]/P0001 ,
		_w11944_,
		_w11955_,
		_w12970_
	);
	LUT4 #(
		.INIT('h0001)
	) name2458 (
		_w12967_,
		_w12968_,
		_w12969_,
		_w12970_,
		_w12971_
	);
	LUT4 #(
		.INIT('h8000)
	) name2459 (
		_w12956_,
		_w12961_,
		_w12966_,
		_w12971_,
		_w12972_
	);
	LUT3 #(
		.INIT('h80)
	) name2460 (
		\wishbone_bd_ram_mem3_reg[209][30]/P0001 ,
		_w11977_,
		_w11984_,
		_w12973_
	);
	LUT3 #(
		.INIT('h80)
	) name2461 (
		\wishbone_bd_ram_mem3_reg[4][30]/P0001 ,
		_w11929_,
		_w11932_,
		_w12974_
	);
	LUT3 #(
		.INIT('h80)
	) name2462 (
		\wishbone_bd_ram_mem3_reg[191][30]/P0001 ,
		_w11942_,
		_w11973_,
		_w12975_
	);
	LUT3 #(
		.INIT('h80)
	) name2463 (
		\wishbone_bd_ram_mem3_reg[228][30]/P0001 ,
		_w11929_,
		_w11982_,
		_w12976_
	);
	LUT4 #(
		.INIT('h0001)
	) name2464 (
		_w12973_,
		_w12974_,
		_w12975_,
		_w12976_,
		_w12977_
	);
	LUT3 #(
		.INIT('h80)
	) name2465 (
		\wishbone_bd_ram_mem3_reg[120][30]/P0001 ,
		_w11990_,
		_w12012_,
		_w12978_
	);
	LUT3 #(
		.INIT('h80)
	) name2466 (
		\wishbone_bd_ram_mem3_reg[202][30]/P0001 ,
		_w11944_,
		_w11945_,
		_w12979_
	);
	LUT3 #(
		.INIT('h80)
	) name2467 (
		\wishbone_bd_ram_mem3_reg[168][30]/P0001 ,
		_w11930_,
		_w11990_,
		_w12980_
	);
	LUT3 #(
		.INIT('h80)
	) name2468 (
		\wishbone_bd_ram_mem3_reg[247][30]/P0001 ,
		_w11952_,
		_w11975_,
		_w12981_
	);
	LUT4 #(
		.INIT('h0001)
	) name2469 (
		_w12978_,
		_w12979_,
		_w12980_,
		_w12981_,
		_w12982_
	);
	LUT3 #(
		.INIT('h80)
	) name2470 (
		\wishbone_bd_ram_mem3_reg[88][30]/P0001 ,
		_w11972_,
		_w11990_,
		_w12983_
	);
	LUT3 #(
		.INIT('h80)
	) name2471 (
		\wishbone_bd_ram_mem3_reg[41][30]/P0001 ,
		_w11957_,
		_w11968_,
		_w12984_
	);
	LUT3 #(
		.INIT('h80)
	) name2472 (
		\wishbone_bd_ram_mem3_reg[40][30]/P0001 ,
		_w11957_,
		_w11990_,
		_w12985_
	);
	LUT3 #(
		.INIT('h80)
	) name2473 (
		\wishbone_bd_ram_mem3_reg[94][30]/P0001 ,
		_w11948_,
		_w11972_,
		_w12986_
	);
	LUT4 #(
		.INIT('h0001)
	) name2474 (
		_w12983_,
		_w12984_,
		_w12985_,
		_w12986_,
		_w12987_
	);
	LUT3 #(
		.INIT('h80)
	) name2475 (
		\wishbone_bd_ram_mem3_reg[217][30]/P0001 ,
		_w11968_,
		_w11984_,
		_w12988_
	);
	LUT3 #(
		.INIT('h80)
	) name2476 (
		\wishbone_bd_ram_mem3_reg[62][30]/P0001 ,
		_w11948_,
		_w11979_,
		_w12989_
	);
	LUT3 #(
		.INIT('h80)
	) name2477 (
		\wishbone_bd_ram_mem3_reg[207][30]/P0001 ,
		_w11945_,
		_w11973_,
		_w12990_
	);
	LUT3 #(
		.INIT('h80)
	) name2478 (
		\wishbone_bd_ram_mem3_reg[16][30]/P0001 ,
		_w11935_,
		_w11941_,
		_w12991_
	);
	LUT4 #(
		.INIT('h0001)
	) name2479 (
		_w12988_,
		_w12989_,
		_w12990_,
		_w12991_,
		_w12992_
	);
	LUT4 #(
		.INIT('h8000)
	) name2480 (
		_w12977_,
		_w12982_,
		_w12987_,
		_w12992_,
		_w12993_
	);
	LUT3 #(
		.INIT('h80)
	) name2481 (
		\wishbone_bd_ram_mem3_reg[171][30]/P0001 ,
		_w11930_,
		_w11936_,
		_w12994_
	);
	LUT3 #(
		.INIT('h80)
	) name2482 (
		\wishbone_bd_ram_mem3_reg[150][30]/P0001 ,
		_w11959_,
		_w11986_,
		_w12995_
	);
	LUT3 #(
		.INIT('h80)
	) name2483 (
		\wishbone_bd_ram_mem3_reg[95][30]/P0001 ,
		_w11972_,
		_w11973_,
		_w12996_
	);
	LUT3 #(
		.INIT('h80)
	) name2484 (
		\wishbone_bd_ram_mem3_reg[90][30]/P0001 ,
		_w11944_,
		_w11972_,
		_w12997_
	);
	LUT4 #(
		.INIT('h0001)
	) name2485 (
		_w12994_,
		_w12995_,
		_w12996_,
		_w12997_,
		_w12998_
	);
	LUT3 #(
		.INIT('h80)
	) name2486 (
		\wishbone_bd_ram_mem3_reg[248][30]/P0001 ,
		_w11952_,
		_w11990_,
		_w12999_
	);
	LUT3 #(
		.INIT('h80)
	) name2487 (
		\wishbone_bd_ram_mem3_reg[126][30]/P0001 ,
		_w11948_,
		_w12012_,
		_w13000_
	);
	LUT3 #(
		.INIT('h80)
	) name2488 (
		\wishbone_bd_ram_mem3_reg[93][30]/P0001 ,
		_w11966_,
		_w11972_,
		_w13001_
	);
	LUT3 #(
		.INIT('h80)
	) name2489 (
		\wishbone_bd_ram_mem3_reg[140][30]/P0001 ,
		_w11954_,
		_w11955_,
		_w13002_
	);
	LUT4 #(
		.INIT('h0001)
	) name2490 (
		_w12999_,
		_w13000_,
		_w13001_,
		_w13002_,
		_w13003_
	);
	LUT3 #(
		.INIT('h80)
	) name2491 (
		\wishbone_bd_ram_mem3_reg[14][30]/P0001 ,
		_w11932_,
		_w11948_,
		_w13004_
	);
	LUT3 #(
		.INIT('h80)
	) name2492 (
		\wishbone_bd_ram_mem3_reg[249][30]/P0001 ,
		_w11952_,
		_w11968_,
		_w13005_
	);
	LUT3 #(
		.INIT('h80)
	) name2493 (
		\wishbone_bd_ram_mem3_reg[162][30]/P0001 ,
		_w11930_,
		_w11963_,
		_w13006_
	);
	LUT3 #(
		.INIT('h80)
	) name2494 (
		\wishbone_bd_ram_mem3_reg[110][30]/P0001 ,
		_w11948_,
		_w11965_,
		_w13007_
	);
	LUT4 #(
		.INIT('h0001)
	) name2495 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13007_,
		_w13008_
	);
	LUT3 #(
		.INIT('h80)
	) name2496 (
		\wishbone_bd_ram_mem3_reg[71][30]/P0001 ,
		_w11949_,
		_w11975_,
		_w13009_
	);
	LUT3 #(
		.INIT('h80)
	) name2497 (
		\wishbone_bd_ram_mem3_reg[124][30]/P0001 ,
		_w11954_,
		_w12012_,
		_w13010_
	);
	LUT3 #(
		.INIT('h80)
	) name2498 (
		\wishbone_bd_ram_mem3_reg[65][30]/P0001 ,
		_w11949_,
		_w11977_,
		_w13011_
	);
	LUT3 #(
		.INIT('h80)
	) name2499 (
		\wishbone_bd_ram_mem3_reg[177][30]/P0001 ,
		_w11942_,
		_w11977_,
		_w13012_
	);
	LUT4 #(
		.INIT('h0001)
	) name2500 (
		_w13009_,
		_w13010_,
		_w13011_,
		_w13012_,
		_w13013_
	);
	LUT4 #(
		.INIT('h8000)
	) name2501 (
		_w12998_,
		_w13003_,
		_w13008_,
		_w13013_,
		_w13014_
	);
	LUT4 #(
		.INIT('h8000)
	) name2502 (
		_w12951_,
		_w12972_,
		_w12993_,
		_w13014_,
		_w13015_
	);
	LUT4 #(
		.INIT('h8000)
	) name2503 (
		_w12760_,
		_w12845_,
		_w12930_,
		_w13015_,
		_w13016_
	);
	LUT4 #(
		.INIT('he4a8)
	) name2504 (
		\wishbone_TxLength_reg[14]/NET0131 ,
		_w12319_,
		_w12669_,
		_w12672_,
		_w13017_
	);
	LUT3 #(
		.INIT('hf2)
	) name2505 (
		_w12303_,
		_w13016_,
		_w13017_,
		_w13018_
	);
	LUT3 #(
		.INIT('h7b)
	) name2506 (
		\rxethmac1_crcrx_Crc_reg[6]/NET0131 ,
		_w10582_,
		_w11574_,
		_w13019_
	);
	LUT3 #(
		.INIT('h7b)
	) name2507 (
		\rxethmac1_crcrx_Crc_reg[0]/NET0131 ,
		_w10582_,
		_w11574_,
		_w13020_
	);
	LUT4 #(
		.INIT('h1113)
	) name2508 (
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		\txethmac1_txstatem1_StatePAD_reg/NET0131 ,
		_w13021_
	);
	LUT3 #(
		.INIT('h70)
	) name2509 (
		_w10801_,
		_w10803_,
		_w13021_,
		_w13022_
	);
	LUT2 #(
		.INIT('h8)
	) name2510 (
		\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[7]/NET0131 ,
		_w13023_
	);
	LUT3 #(
		.INIT('h80)
	) name2511 (
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[8]/NET0131 ,
		_w13024_
	);
	LUT2 #(
		.INIT('h8)
	) name2512 (
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		_w13025_
	);
	LUT4 #(
		.INIT('h8000)
	) name2513 (
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		_w13026_
	);
	LUT2 #(
		.INIT('h8)
	) name2514 (
		\txethmac1_txcounters1_ByteCnt_reg[10]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[11]/NET0131 ,
		_w13027_
	);
	LUT3 #(
		.INIT('h80)
	) name2515 (
		\txethmac1_txcounters1_ByteCnt_reg[10]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[11]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 ,
		_w13028_
	);
	LUT4 #(
		.INIT('h8000)
	) name2516 (
		_w13023_,
		_w13024_,
		_w13026_,
		_w13028_,
		_w13029_
	);
	LUT4 #(
		.INIT('h8000)
	) name2517 (
		\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[13]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[14]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[15]/NET0131 ,
		_w13030_
	);
	LUT3 #(
		.INIT('h70)
	) name2518 (
		_w10801_,
		_w10803_,
		_w13030_,
		_w13031_
	);
	LUT3 #(
		.INIT('h15)
	) name2519 (
		_w13022_,
		_w13029_,
		_w13031_,
		_w13032_
	);
	LUT3 #(
		.INIT('h80)
	) name2520 (
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		_w13033_
	);
	LUT4 #(
		.INIT('h1500)
	) name2521 (
		_w13022_,
		_w13029_,
		_w13031_,
		_w13033_,
		_w13034_
	);
	LUT2 #(
		.INIT('h8)
	) name2522 (
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 ,
		_w13035_
	);
	LUT3 #(
		.INIT('h80)
	) name2523 (
		_w13023_,
		_w13024_,
		_w13035_,
		_w13036_
	);
	LUT3 #(
		.INIT('h80)
	) name2524 (
		\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[13]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[14]/NET0131 ,
		_w13037_
	);
	LUT2 #(
		.INIT('h8)
	) name2525 (
		_w13027_,
		_w13037_,
		_w13038_
	);
	LUT3 #(
		.INIT('h01)
	) name2526 (
		\txethmac1_PacketFinished_q_reg/NET0131 ,
		_w10936_,
		_w10937_,
		_w13039_
	);
	LUT3 #(
		.INIT('h70)
	) name2527 (
		_w10791_,
		_w10967_,
		_w13039_,
		_w13040_
	);
	LUT4 #(
		.INIT('h2a00)
	) name2528 (
		\txethmac1_txcounters1_ByteCnt_reg[15]/NET0131 ,
		_w10791_,
		_w10967_,
		_w13039_,
		_w13041_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2529 (
		_w13034_,
		_w13036_,
		_w13038_,
		_w13041_,
		_w13042_
	);
	LUT4 #(
		.INIT('h1500)
	) name2530 (
		\txethmac1_txcounters1_ByteCnt_reg[15]/NET0131 ,
		_w10791_,
		_w10967_,
		_w13039_,
		_w13043_
	);
	LUT4 #(
		.INIT('h8000)
	) name2531 (
		_w13034_,
		_w13036_,
		_w13038_,
		_w13043_,
		_w13044_
	);
	LUT2 #(
		.INIT('he)
	) name2532 (
		_w13042_,
		_w13044_,
		_w13045_
	);
	LUT3 #(
		.INIT('ha2)
	) name2533 (
		\wishbone_TxPointerMSB_reg[2]/NET0131 ,
		_w11900_,
		_w11909_,
		_w13046_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2534 (
		\m_wb_adr_o[2]_pad ,
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w13047_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2535 (
		\wishbone_RxPointerMSB_reg[2]/NET0131 ,
		_w11902_,
		_w11905_,
		_w13047_,
		_w13048_
	);
	LUT2 #(
		.INIT('h1)
	) name2536 (
		_w13046_,
		_w13048_,
		_w13049_
	);
	LUT3 #(
		.INIT('h07)
	) name2537 (
		_w11868_,
		_w11875_,
		_w11911_,
		_w13050_
	);
	LUT3 #(
		.INIT('h80)
	) name2538 (
		_w11870_,
		_w11873_,
		_w13050_,
		_w13051_
	);
	LUT4 #(
		.INIT('h80aa)
	) name2539 (
		\wishbone_TxPointerMSB_reg[2]/NET0131 ,
		_w11866_,
		_w11867_,
		_w11883_,
		_w13052_
	);
	LUT2 #(
		.INIT('h4)
	) name2540 (
		_w11882_,
		_w13052_,
		_w13053_
	);
	LUT4 #(
		.INIT('h5554)
	) name2541 (
		\m_wb_adr_o[2]_pad ,
		_w11887_,
		_w13051_,
		_w13053_,
		_w13054_
	);
	LUT3 #(
		.INIT('h07)
	) name2542 (
		\m_wb_adr_o[2]_pad ,
		_w11907_,
		_w13054_,
		_w13055_
	);
	LUT2 #(
		.INIT('h7)
	) name2543 (
		_w13049_,
		_w13055_,
		_w13056_
	);
	LUT3 #(
		.INIT('h80)
	) name2544 (
		\wishbone_bd_ram_mem3_reg[143][24]/P0001 ,
		_w11955_,
		_w11973_,
		_w13057_
	);
	LUT3 #(
		.INIT('h80)
	) name2545 (
		\wishbone_bd_ram_mem3_reg[8][24]/P0001 ,
		_w11932_,
		_w11990_,
		_w13058_
	);
	LUT3 #(
		.INIT('h80)
	) name2546 (
		\wishbone_bd_ram_mem3_reg[142][24]/P0001 ,
		_w11948_,
		_w11955_,
		_w13059_
	);
	LUT3 #(
		.INIT('h80)
	) name2547 (
		\wishbone_bd_ram_mem3_reg[115][24]/P0001 ,
		_w11938_,
		_w12012_,
		_w13060_
	);
	LUT4 #(
		.INIT('h0001)
	) name2548 (
		_w13057_,
		_w13058_,
		_w13059_,
		_w13060_,
		_w13061_
	);
	LUT3 #(
		.INIT('h80)
	) name2549 (
		\wishbone_bd_ram_mem3_reg[111][24]/P0001 ,
		_w11965_,
		_w11973_,
		_w13062_
	);
	LUT3 #(
		.INIT('h80)
	) name2550 (
		\wishbone_bd_ram_mem3_reg[228][24]/P0001 ,
		_w11929_,
		_w11982_,
		_w13063_
	);
	LUT3 #(
		.INIT('h80)
	) name2551 (
		\wishbone_bd_ram_mem3_reg[47][24]/P0001 ,
		_w11957_,
		_w11973_,
		_w13064_
	);
	LUT3 #(
		.INIT('h80)
	) name2552 (
		\wishbone_bd_ram_mem3_reg[185][24]/P0001 ,
		_w11942_,
		_w11968_,
		_w13065_
	);
	LUT4 #(
		.INIT('h0001)
	) name2553 (
		_w13062_,
		_w13063_,
		_w13064_,
		_w13065_,
		_w13066_
	);
	LUT3 #(
		.INIT('h80)
	) name2554 (
		\wishbone_bd_ram_mem3_reg[249][24]/P0001 ,
		_w11952_,
		_w11968_,
		_w13067_
	);
	LUT3 #(
		.INIT('h80)
	) name2555 (
		\wishbone_bd_ram_mem3_reg[106][24]/P0001 ,
		_w11944_,
		_w11965_,
		_w13068_
	);
	LUT3 #(
		.INIT('h80)
	) name2556 (
		\wishbone_bd_ram_mem3_reg[65][24]/P0001 ,
		_w11949_,
		_w11977_,
		_w13069_
	);
	LUT3 #(
		.INIT('h80)
	) name2557 (
		\wishbone_bd_ram_mem3_reg[150][24]/P0001 ,
		_w11959_,
		_w11986_,
		_w13070_
	);
	LUT4 #(
		.INIT('h0001)
	) name2558 (
		_w13067_,
		_w13068_,
		_w13069_,
		_w13070_,
		_w13071_
	);
	LUT3 #(
		.INIT('h80)
	) name2559 (
		\wishbone_bd_ram_mem3_reg[154][24]/P0001 ,
		_w11944_,
		_w11959_,
		_w13072_
	);
	LUT3 #(
		.INIT('h80)
	) name2560 (
		\wishbone_bd_ram_mem3_reg[129][24]/P0001 ,
		_w11955_,
		_w11977_,
		_w13073_
	);
	LUT3 #(
		.INIT('h80)
	) name2561 (
		\wishbone_bd_ram_mem3_reg[172][24]/P0001 ,
		_w11930_,
		_w11954_,
		_w13074_
	);
	LUT3 #(
		.INIT('h80)
	) name2562 (
		\wishbone_bd_ram_mem3_reg[28][24]/P0001 ,
		_w11935_,
		_w11954_,
		_w13075_
	);
	LUT4 #(
		.INIT('h0001)
	) name2563 (
		_w13072_,
		_w13073_,
		_w13074_,
		_w13075_,
		_w13076_
	);
	LUT4 #(
		.INIT('h8000)
	) name2564 (
		_w13061_,
		_w13066_,
		_w13071_,
		_w13076_,
		_w13077_
	);
	LUT3 #(
		.INIT('h80)
	) name2565 (
		\wishbone_bd_ram_mem3_reg[171][24]/P0001 ,
		_w11930_,
		_w11936_,
		_w13078_
	);
	LUT3 #(
		.INIT('h80)
	) name2566 (
		\wishbone_bd_ram_mem3_reg[40][24]/P0001 ,
		_w11957_,
		_w11990_,
		_w13079_
	);
	LUT3 #(
		.INIT('h80)
	) name2567 (
		\wishbone_bd_ram_mem3_reg[2][24]/P0001 ,
		_w11932_,
		_w11963_,
		_w13080_
	);
	LUT3 #(
		.INIT('h80)
	) name2568 (
		\wishbone_bd_ram_mem3_reg[75][24]/P0001 ,
		_w11936_,
		_w11949_,
		_w13081_
	);
	LUT4 #(
		.INIT('h0001)
	) name2569 (
		_w13078_,
		_w13079_,
		_w13080_,
		_w13081_,
		_w13082_
	);
	LUT3 #(
		.INIT('h80)
	) name2570 (
		\wishbone_bd_ram_mem3_reg[181][24]/P0001 ,
		_w11933_,
		_w11942_,
		_w13083_
	);
	LUT3 #(
		.INIT('h80)
	) name2571 (
		\wishbone_bd_ram_mem3_reg[244][24]/P0001 ,
		_w11929_,
		_w11952_,
		_w13084_
	);
	LUT3 #(
		.INIT('h80)
	) name2572 (
		\wishbone_bd_ram_mem3_reg[109][24]/P0001 ,
		_w11965_,
		_w11966_,
		_w13085_
	);
	LUT3 #(
		.INIT('h80)
	) name2573 (
		\wishbone_bd_ram_mem3_reg[88][24]/P0001 ,
		_w11972_,
		_w11990_,
		_w13086_
	);
	LUT4 #(
		.INIT('h0001)
	) name2574 (
		_w13083_,
		_w13084_,
		_w13085_,
		_w13086_,
		_w13087_
	);
	LUT3 #(
		.INIT('h80)
	) name2575 (
		\wishbone_bd_ram_mem3_reg[120][24]/P0001 ,
		_w11990_,
		_w12012_,
		_w13088_
	);
	LUT3 #(
		.INIT('h80)
	) name2576 (
		\wishbone_bd_ram_mem3_reg[250][24]/P0001 ,
		_w11944_,
		_w11952_,
		_w13089_
	);
	LUT3 #(
		.INIT('h80)
	) name2577 (
		\wishbone_bd_ram_mem3_reg[215][24]/P0001 ,
		_w11975_,
		_w11984_,
		_w13090_
	);
	LUT3 #(
		.INIT('h80)
	) name2578 (
		\wishbone_bd_ram_mem3_reg[67][24]/P0001 ,
		_w11938_,
		_w11949_,
		_w13091_
	);
	LUT4 #(
		.INIT('h0001)
	) name2579 (
		_w13088_,
		_w13089_,
		_w13090_,
		_w13091_,
		_w13092_
	);
	LUT3 #(
		.INIT('h80)
	) name2580 (
		\wishbone_bd_ram_mem3_reg[80][24]/P0001 ,
		_w11941_,
		_w11972_,
		_w13093_
	);
	LUT3 #(
		.INIT('h80)
	) name2581 (
		\wishbone_bd_ram_mem3_reg[140][24]/P0001 ,
		_w11954_,
		_w11955_,
		_w13094_
	);
	LUT3 #(
		.INIT('h80)
	) name2582 (
		\wishbone_bd_ram_mem3_reg[160][24]/P0001 ,
		_w11930_,
		_w11941_,
		_w13095_
	);
	LUT3 #(
		.INIT('h80)
	) name2583 (
		\wishbone_bd_ram_mem3_reg[219][24]/P0001 ,
		_w11936_,
		_w11984_,
		_w13096_
	);
	LUT4 #(
		.INIT('h0001)
	) name2584 (
		_w13093_,
		_w13094_,
		_w13095_,
		_w13096_,
		_w13097_
	);
	LUT4 #(
		.INIT('h8000)
	) name2585 (
		_w13082_,
		_w13087_,
		_w13092_,
		_w13097_,
		_w13098_
	);
	LUT3 #(
		.INIT('h80)
	) name2586 (
		\wishbone_bd_ram_mem3_reg[212][24]/P0001 ,
		_w11929_,
		_w11984_,
		_w13099_
	);
	LUT3 #(
		.INIT('h80)
	) name2587 (
		\wishbone_bd_ram_mem3_reg[10][24]/P0001 ,
		_w11932_,
		_w11944_,
		_w13100_
	);
	LUT3 #(
		.INIT('h80)
	) name2588 (
		\wishbone_bd_ram_mem3_reg[139][24]/P0001 ,
		_w11936_,
		_w11955_,
		_w13101_
	);
	LUT3 #(
		.INIT('h80)
	) name2589 (
		\wishbone_bd_ram_mem3_reg[30][24]/P0001 ,
		_w11935_,
		_w11948_,
		_w13102_
	);
	LUT4 #(
		.INIT('h0001)
	) name2590 (
		_w13099_,
		_w13100_,
		_w13101_,
		_w13102_,
		_w13103_
	);
	LUT3 #(
		.INIT('h80)
	) name2591 (
		\wishbone_bd_ram_mem3_reg[247][24]/P0001 ,
		_w11952_,
		_w11975_,
		_w13104_
	);
	LUT3 #(
		.INIT('h80)
	) name2592 (
		\wishbone_bd_ram_mem3_reg[29][24]/P0001 ,
		_w11935_,
		_w11966_,
		_w13105_
	);
	LUT3 #(
		.INIT('h80)
	) name2593 (
		\wishbone_bd_ram_mem3_reg[216][24]/P0001 ,
		_w11984_,
		_w11990_,
		_w13106_
	);
	LUT3 #(
		.INIT('h80)
	) name2594 (
		\wishbone_bd_ram_mem3_reg[145][24]/P0001 ,
		_w11959_,
		_w11977_,
		_w13107_
	);
	LUT4 #(
		.INIT('h0001)
	) name2595 (
		_w13104_,
		_w13105_,
		_w13106_,
		_w13107_,
		_w13108_
	);
	LUT3 #(
		.INIT('h80)
	) name2596 (
		\wishbone_bd_ram_mem3_reg[192][24]/P0001 ,
		_w11941_,
		_w11945_,
		_w13109_
	);
	LUT3 #(
		.INIT('h80)
	) name2597 (
		\wishbone_bd_ram_mem3_reg[162][24]/P0001 ,
		_w11930_,
		_w11963_,
		_w13110_
	);
	LUT3 #(
		.INIT('h80)
	) name2598 (
		\wishbone_bd_ram_mem3_reg[36][24]/P0001 ,
		_w11929_,
		_w11957_,
		_w13111_
	);
	LUT3 #(
		.INIT('h80)
	) name2599 (
		\wishbone_bd_ram_mem3_reg[9][24]/P0001 ,
		_w11932_,
		_w11968_,
		_w13112_
	);
	LUT4 #(
		.INIT('h0001)
	) name2600 (
		_w13109_,
		_w13110_,
		_w13111_,
		_w13112_,
		_w13113_
	);
	LUT3 #(
		.INIT('h80)
	) name2601 (
		\wishbone_bd_ram_mem3_reg[132][24]/P0001 ,
		_w11929_,
		_w11955_,
		_w13114_
	);
	LUT3 #(
		.INIT('h80)
	) name2602 (
		\wishbone_bd_ram_mem3_reg[187][24]/P0001 ,
		_w11936_,
		_w11942_,
		_w13115_
	);
	LUT3 #(
		.INIT('h80)
	) name2603 (
		\wishbone_bd_ram_mem3_reg[43][24]/P0001 ,
		_w11936_,
		_w11957_,
		_w13116_
	);
	LUT3 #(
		.INIT('h80)
	) name2604 (
		\wishbone_bd_ram_mem3_reg[239][24]/P0001 ,
		_w11973_,
		_w11982_,
		_w13117_
	);
	LUT4 #(
		.INIT('h0001)
	) name2605 (
		_w13114_,
		_w13115_,
		_w13116_,
		_w13117_,
		_w13118_
	);
	LUT4 #(
		.INIT('h8000)
	) name2606 (
		_w13103_,
		_w13108_,
		_w13113_,
		_w13118_,
		_w13119_
	);
	LUT3 #(
		.INIT('h80)
	) name2607 (
		\wishbone_bd_ram_mem3_reg[168][24]/P0001 ,
		_w11930_,
		_w11990_,
		_w13120_
	);
	LUT3 #(
		.INIT('h80)
	) name2608 (
		\wishbone_bd_ram_mem3_reg[182][24]/P0001 ,
		_w11942_,
		_w11986_,
		_w13121_
	);
	LUT3 #(
		.INIT('h80)
	) name2609 (
		\wishbone_bd_ram_mem3_reg[230][24]/P0001 ,
		_w11982_,
		_w11986_,
		_w13122_
	);
	LUT3 #(
		.INIT('h80)
	) name2610 (
		\wishbone_bd_ram_mem3_reg[21][24]/P0001 ,
		_w11933_,
		_w11935_,
		_w13123_
	);
	LUT4 #(
		.INIT('h0001)
	) name2611 (
		_w13120_,
		_w13121_,
		_w13122_,
		_w13123_,
		_w13124_
	);
	LUT3 #(
		.INIT('h80)
	) name2612 (
		\wishbone_bd_ram_mem3_reg[178][24]/P0001 ,
		_w11942_,
		_w11963_,
		_w13125_
	);
	LUT3 #(
		.INIT('h80)
	) name2613 (
		\wishbone_bd_ram_mem3_reg[127][24]/P0001 ,
		_w11973_,
		_w12012_,
		_w13126_
	);
	LUT3 #(
		.INIT('h80)
	) name2614 (
		\wishbone_bd_ram_mem3_reg[60][24]/P0001 ,
		_w11954_,
		_w11979_,
		_w13127_
	);
	LUT3 #(
		.INIT('h80)
	) name2615 (
		\wishbone_bd_ram_mem3_reg[18][24]/P0001 ,
		_w11935_,
		_w11963_,
		_w13128_
	);
	LUT4 #(
		.INIT('h0001)
	) name2616 (
		_w13125_,
		_w13126_,
		_w13127_,
		_w13128_,
		_w13129_
	);
	LUT3 #(
		.INIT('h80)
	) name2617 (
		\wishbone_bd_ram_mem3_reg[41][24]/P0001 ,
		_w11957_,
		_w11968_,
		_w13130_
	);
	LUT3 #(
		.INIT('h80)
	) name2618 (
		\wishbone_bd_ram_mem3_reg[52][24]/P0001 ,
		_w11929_,
		_w11979_,
		_w13131_
	);
	LUT3 #(
		.INIT('h80)
	) name2619 (
		\wishbone_bd_ram_mem3_reg[147][24]/P0001 ,
		_w11938_,
		_w11959_,
		_w13132_
	);
	LUT3 #(
		.INIT('h80)
	) name2620 (
		\wishbone_bd_ram_mem3_reg[20][24]/P0001 ,
		_w11929_,
		_w11935_,
		_w13133_
	);
	LUT4 #(
		.INIT('h0001)
	) name2621 (
		_w13130_,
		_w13131_,
		_w13132_,
		_w13133_,
		_w13134_
	);
	LUT3 #(
		.INIT('h80)
	) name2622 (
		\wishbone_bd_ram_mem3_reg[22][24]/P0001 ,
		_w11935_,
		_w11986_,
		_w13135_
	);
	LUT3 #(
		.INIT('h80)
	) name2623 (
		\wishbone_bd_ram_mem3_reg[97][24]/P0001 ,
		_w11965_,
		_w11977_,
		_w13136_
	);
	LUT3 #(
		.INIT('h80)
	) name2624 (
		\wishbone_bd_ram_mem3_reg[255][24]/P0001 ,
		_w11952_,
		_w11973_,
		_w13137_
	);
	LUT3 #(
		.INIT('h80)
	) name2625 (
		\wishbone_bd_ram_mem3_reg[164][24]/P0001 ,
		_w11929_,
		_w11930_,
		_w13138_
	);
	LUT4 #(
		.INIT('h0001)
	) name2626 (
		_w13135_,
		_w13136_,
		_w13137_,
		_w13138_,
		_w13139_
	);
	LUT4 #(
		.INIT('h8000)
	) name2627 (
		_w13124_,
		_w13129_,
		_w13134_,
		_w13139_,
		_w13140_
	);
	LUT4 #(
		.INIT('h8000)
	) name2628 (
		_w13077_,
		_w13098_,
		_w13119_,
		_w13140_,
		_w13141_
	);
	LUT3 #(
		.INIT('h80)
	) name2629 (
		\wishbone_bd_ram_mem3_reg[201][24]/P0001 ,
		_w11945_,
		_w11968_,
		_w13142_
	);
	LUT3 #(
		.INIT('h80)
	) name2630 (
		\wishbone_bd_ram_mem3_reg[91][24]/P0001 ,
		_w11936_,
		_w11972_,
		_w13143_
	);
	LUT3 #(
		.INIT('h80)
	) name2631 (
		\wishbone_bd_ram_mem3_reg[211][24]/P0001 ,
		_w11938_,
		_w11984_,
		_w13144_
	);
	LUT3 #(
		.INIT('h80)
	) name2632 (
		\wishbone_bd_ram_mem3_reg[149][24]/P0001 ,
		_w11933_,
		_w11959_,
		_w13145_
	);
	LUT4 #(
		.INIT('h0001)
	) name2633 (
		_w13142_,
		_w13143_,
		_w13144_,
		_w13145_,
		_w13146_
	);
	LUT3 #(
		.INIT('h80)
	) name2634 (
		\wishbone_bd_ram_mem3_reg[205][24]/P0001 ,
		_w11945_,
		_w11966_,
		_w13147_
	);
	LUT3 #(
		.INIT('h80)
	) name2635 (
		\wishbone_bd_ram_mem3_reg[176][24]/P0001 ,
		_w11941_,
		_w11942_,
		_w13148_
	);
	LUT3 #(
		.INIT('h80)
	) name2636 (
		\wishbone_bd_ram_mem3_reg[131][24]/P0001 ,
		_w11938_,
		_w11955_,
		_w13149_
	);
	LUT3 #(
		.INIT('h80)
	) name2637 (
		\wishbone_bd_ram_mem3_reg[39][24]/P0001 ,
		_w11957_,
		_w11975_,
		_w13150_
	);
	LUT4 #(
		.INIT('h0001)
	) name2638 (
		_w13147_,
		_w13148_,
		_w13149_,
		_w13150_,
		_w13151_
	);
	LUT3 #(
		.INIT('h80)
	) name2639 (
		\wishbone_bd_ram_mem3_reg[35][24]/P0001 ,
		_w11938_,
		_w11957_,
		_w13152_
	);
	LUT3 #(
		.INIT('h80)
	) name2640 (
		\wishbone_bd_ram_mem3_reg[218][24]/P0001 ,
		_w11944_,
		_w11984_,
		_w13153_
	);
	LUT3 #(
		.INIT('h80)
	) name2641 (
		\wishbone_bd_ram_mem3_reg[241][24]/P0001 ,
		_w11952_,
		_w11977_,
		_w13154_
	);
	LUT3 #(
		.INIT('h80)
	) name2642 (
		\wishbone_bd_ram_mem3_reg[170][24]/P0001 ,
		_w11930_,
		_w11944_,
		_w13155_
	);
	LUT4 #(
		.INIT('h0001)
	) name2643 (
		_w13152_,
		_w13153_,
		_w13154_,
		_w13155_,
		_w13156_
	);
	LUT3 #(
		.INIT('h80)
	) name2644 (
		\wishbone_bd_ram_mem3_reg[196][24]/P0001 ,
		_w11929_,
		_w11945_,
		_w13157_
	);
	LUT3 #(
		.INIT('h80)
	) name2645 (
		\wishbone_bd_ram_mem3_reg[84][24]/P0001 ,
		_w11929_,
		_w11972_,
		_w13158_
	);
	LUT3 #(
		.INIT('h80)
	) name2646 (
		\wishbone_bd_ram_mem3_reg[121][24]/P0001 ,
		_w11968_,
		_w12012_,
		_w13159_
	);
	LUT3 #(
		.INIT('h80)
	) name2647 (
		\wishbone_bd_ram_mem3_reg[83][24]/P0001 ,
		_w11938_,
		_w11972_,
		_w13160_
	);
	LUT4 #(
		.INIT('h0001)
	) name2648 (
		_w13157_,
		_w13158_,
		_w13159_,
		_w13160_,
		_w13161_
	);
	LUT4 #(
		.INIT('h8000)
	) name2649 (
		_w13146_,
		_w13151_,
		_w13156_,
		_w13161_,
		_w13162_
	);
	LUT3 #(
		.INIT('h80)
	) name2650 (
		\wishbone_bd_ram_mem3_reg[3][24]/P0001 ,
		_w11932_,
		_w11938_,
		_w13163_
	);
	LUT3 #(
		.INIT('h80)
	) name2651 (
		\wishbone_bd_ram_mem3_reg[126][24]/P0001 ,
		_w11948_,
		_w12012_,
		_w13164_
	);
	LUT3 #(
		.INIT('h80)
	) name2652 (
		\wishbone_bd_ram_mem3_reg[34][24]/P0001 ,
		_w11957_,
		_w11963_,
		_w13165_
	);
	LUT3 #(
		.INIT('h80)
	) name2653 (
		\wishbone_bd_ram_mem3_reg[55][24]/P0001 ,
		_w11975_,
		_w11979_,
		_w13166_
	);
	LUT4 #(
		.INIT('h0001)
	) name2654 (
		_w13163_,
		_w13164_,
		_w13165_,
		_w13166_,
		_w13167_
	);
	LUT3 #(
		.INIT('h80)
	) name2655 (
		\wishbone_bd_ram_mem3_reg[78][24]/P0001 ,
		_w11948_,
		_w11949_,
		_w13168_
	);
	LUT3 #(
		.INIT('h80)
	) name2656 (
		\wishbone_bd_ram_mem3_reg[157][24]/P0001 ,
		_w11959_,
		_w11966_,
		_w13169_
	);
	LUT3 #(
		.INIT('h80)
	) name2657 (
		\wishbone_bd_ram_mem3_reg[17][24]/P0001 ,
		_w11935_,
		_w11977_,
		_w13170_
	);
	LUT3 #(
		.INIT('h80)
	) name2658 (
		\wishbone_bd_ram_mem3_reg[0][24]/P0001 ,
		_w11932_,
		_w11941_,
		_w13171_
	);
	LUT4 #(
		.INIT('h0001)
	) name2659 (
		_w13168_,
		_w13169_,
		_w13170_,
		_w13171_,
		_w13172_
	);
	LUT3 #(
		.INIT('h80)
	) name2660 (
		\wishbone_bd_ram_mem3_reg[144][24]/P0001 ,
		_w11941_,
		_w11959_,
		_w13173_
	);
	LUT3 #(
		.INIT('h80)
	) name2661 (
		\wishbone_bd_ram_mem3_reg[227][24]/P0001 ,
		_w11938_,
		_w11982_,
		_w13174_
	);
	LUT3 #(
		.INIT('h80)
	) name2662 (
		\wishbone_bd_ram_mem3_reg[57][24]/P0001 ,
		_w11968_,
		_w11979_,
		_w13175_
	);
	LUT3 #(
		.INIT('h80)
	) name2663 (
		\wishbone_bd_ram_mem3_reg[188][24]/P0001 ,
		_w11942_,
		_w11954_,
		_w13176_
	);
	LUT4 #(
		.INIT('h0001)
	) name2664 (
		_w13173_,
		_w13174_,
		_w13175_,
		_w13176_,
		_w13177_
	);
	LUT3 #(
		.INIT('h80)
	) name2665 (
		\wishbone_bd_ram_mem3_reg[104][24]/P0001 ,
		_w11965_,
		_w11990_,
		_w13178_
	);
	LUT3 #(
		.INIT('h80)
	) name2666 (
		\wishbone_bd_ram_mem3_reg[252][24]/P0001 ,
		_w11952_,
		_w11954_,
		_w13179_
	);
	LUT3 #(
		.INIT('h80)
	) name2667 (
		\wishbone_bd_ram_mem3_reg[197][24]/P0001 ,
		_w11933_,
		_w11945_,
		_w13180_
	);
	LUT3 #(
		.INIT('h80)
	) name2668 (
		\wishbone_bd_ram_mem3_reg[137][24]/P0001 ,
		_w11955_,
		_w11968_,
		_w13181_
	);
	LUT4 #(
		.INIT('h0001)
	) name2669 (
		_w13178_,
		_w13179_,
		_w13180_,
		_w13181_,
		_w13182_
	);
	LUT4 #(
		.INIT('h8000)
	) name2670 (
		_w13167_,
		_w13172_,
		_w13177_,
		_w13182_,
		_w13183_
	);
	LUT3 #(
		.INIT('h80)
	) name2671 (
		\wishbone_bd_ram_mem3_reg[66][24]/P0001 ,
		_w11949_,
		_w11963_,
		_w13184_
	);
	LUT3 #(
		.INIT('h80)
	) name2672 (
		\wishbone_bd_ram_mem3_reg[105][24]/P0001 ,
		_w11965_,
		_w11968_,
		_w13185_
	);
	LUT3 #(
		.INIT('h80)
	) name2673 (
		\wishbone_bd_ram_mem3_reg[89][24]/P0001 ,
		_w11968_,
		_w11972_,
		_w13186_
	);
	LUT3 #(
		.INIT('h80)
	) name2674 (
		\wishbone_bd_ram_mem3_reg[224][24]/P0001 ,
		_w11941_,
		_w11982_,
		_w13187_
	);
	LUT4 #(
		.INIT('h0001)
	) name2675 (
		_w13184_,
		_w13185_,
		_w13186_,
		_w13187_,
		_w13188_
	);
	LUT3 #(
		.INIT('h80)
	) name2676 (
		\wishbone_bd_ram_mem3_reg[173][24]/P0001 ,
		_w11930_,
		_w11966_,
		_w13189_
	);
	LUT3 #(
		.INIT('h80)
	) name2677 (
		\wishbone_bd_ram_mem3_reg[226][24]/P0001 ,
		_w11963_,
		_w11982_,
		_w13190_
	);
	LUT3 #(
		.INIT('h80)
	) name2678 (
		\wishbone_bd_ram_mem3_reg[204][24]/P0001 ,
		_w11945_,
		_w11954_,
		_w13191_
	);
	LUT3 #(
		.INIT('h80)
	) name2679 (
		\wishbone_bd_ram_mem3_reg[24][24]/P0001 ,
		_w11935_,
		_w11990_,
		_w13192_
	);
	LUT4 #(
		.INIT('h0001)
	) name2680 (
		_w13189_,
		_w13190_,
		_w13191_,
		_w13192_,
		_w13193_
	);
	LUT3 #(
		.INIT('h80)
	) name2681 (
		\wishbone_bd_ram_mem3_reg[158][24]/P0001 ,
		_w11948_,
		_w11959_,
		_w13194_
	);
	LUT3 #(
		.INIT('h80)
	) name2682 (
		\wishbone_bd_ram_mem3_reg[26][24]/P0001 ,
		_w11935_,
		_w11944_,
		_w13195_
	);
	LUT3 #(
		.INIT('h80)
	) name2683 (
		\wishbone_bd_ram_mem3_reg[165][24]/P0001 ,
		_w11930_,
		_w11933_,
		_w13196_
	);
	LUT3 #(
		.INIT('h80)
	) name2684 (
		\wishbone_bd_ram_mem3_reg[209][24]/P0001 ,
		_w11977_,
		_w11984_,
		_w13197_
	);
	LUT4 #(
		.INIT('h0001)
	) name2685 (
		_w13194_,
		_w13195_,
		_w13196_,
		_w13197_,
		_w13198_
	);
	LUT3 #(
		.INIT('h80)
	) name2686 (
		\wishbone_bd_ram_mem3_reg[90][24]/P0001 ,
		_w11944_,
		_w11972_,
		_w13199_
	);
	LUT3 #(
		.INIT('h80)
	) name2687 (
		\wishbone_bd_ram_mem3_reg[184][24]/P0001 ,
		_w11942_,
		_w11990_,
		_w13200_
	);
	LUT3 #(
		.INIT('h80)
	) name2688 (
		\wishbone_bd_ram_mem3_reg[73][24]/P0001 ,
		_w11949_,
		_w11968_,
		_w13201_
	);
	LUT3 #(
		.INIT('h80)
	) name2689 (
		\wishbone_bd_ram_mem3_reg[31][24]/P0001 ,
		_w11935_,
		_w11973_,
		_w13202_
	);
	LUT4 #(
		.INIT('h0001)
	) name2690 (
		_w13199_,
		_w13200_,
		_w13201_,
		_w13202_,
		_w13203_
	);
	LUT4 #(
		.INIT('h8000)
	) name2691 (
		_w13188_,
		_w13193_,
		_w13198_,
		_w13203_,
		_w13204_
	);
	LUT3 #(
		.INIT('h80)
	) name2692 (
		\wishbone_bd_ram_mem3_reg[130][24]/P0001 ,
		_w11955_,
		_w11963_,
		_w13205_
	);
	LUT3 #(
		.INIT('h80)
	) name2693 (
		\wishbone_bd_ram_mem3_reg[133][24]/P0001 ,
		_w11933_,
		_w11955_,
		_w13206_
	);
	LUT3 #(
		.INIT('h80)
	) name2694 (
		\wishbone_bd_ram_mem3_reg[152][24]/P0001 ,
		_w11959_,
		_w11990_,
		_w13207_
	);
	LUT3 #(
		.INIT('h80)
	) name2695 (
		\wishbone_bd_ram_mem3_reg[25][24]/P0001 ,
		_w11935_,
		_w11968_,
		_w13208_
	);
	LUT4 #(
		.INIT('h0001)
	) name2696 (
		_w13205_,
		_w13206_,
		_w13207_,
		_w13208_,
		_w13209_
	);
	LUT3 #(
		.INIT('h80)
	) name2697 (
		\wishbone_bd_ram_mem3_reg[100][24]/P0001 ,
		_w11929_,
		_w11965_,
		_w13210_
	);
	LUT3 #(
		.INIT('h80)
	) name2698 (
		\wishbone_bd_ram_mem3_reg[229][24]/P0001 ,
		_w11933_,
		_w11982_,
		_w13211_
	);
	LUT3 #(
		.INIT('h80)
	) name2699 (
		\wishbone_bd_ram_mem3_reg[110][24]/P0001 ,
		_w11948_,
		_w11965_,
		_w13212_
	);
	LUT3 #(
		.INIT('h80)
	) name2700 (
		\wishbone_bd_ram_mem3_reg[99][24]/P0001 ,
		_w11938_,
		_w11965_,
		_w13213_
	);
	LUT4 #(
		.INIT('h0001)
	) name2701 (
		_w13210_,
		_w13211_,
		_w13212_,
		_w13213_,
		_w13214_
	);
	LUT3 #(
		.INIT('h80)
	) name2702 (
		\wishbone_bd_ram_mem3_reg[114][24]/P0001 ,
		_w11963_,
		_w12012_,
		_w13215_
	);
	LUT3 #(
		.INIT('h80)
	) name2703 (
		\wishbone_bd_ram_mem3_reg[93][24]/P0001 ,
		_w11966_,
		_w11972_,
		_w13216_
	);
	LUT3 #(
		.INIT('h80)
	) name2704 (
		\wishbone_bd_ram_mem3_reg[141][24]/P0001 ,
		_w11955_,
		_w11966_,
		_w13217_
	);
	LUT3 #(
		.INIT('h80)
	) name2705 (
		\wishbone_bd_ram_mem3_reg[146][24]/P0001 ,
		_w11959_,
		_w11963_,
		_w13218_
	);
	LUT4 #(
		.INIT('h0001)
	) name2706 (
		_w13215_,
		_w13216_,
		_w13217_,
		_w13218_,
		_w13219_
	);
	LUT3 #(
		.INIT('h80)
	) name2707 (
		\wishbone_bd_ram_mem3_reg[220][24]/P0001 ,
		_w11954_,
		_w11984_,
		_w13220_
	);
	LUT3 #(
		.INIT('h80)
	) name2708 (
		\wishbone_bd_ram_mem3_reg[245][24]/P0001 ,
		_w11933_,
		_w11952_,
		_w13221_
	);
	LUT3 #(
		.INIT('h80)
	) name2709 (
		\wishbone_bd_ram_mem3_reg[33][24]/P0001 ,
		_w11957_,
		_w11977_,
		_w13222_
	);
	LUT3 #(
		.INIT('h80)
	) name2710 (
		\wishbone_bd_ram_mem3_reg[61][24]/P0001 ,
		_w11966_,
		_w11979_,
		_w13223_
	);
	LUT4 #(
		.INIT('h0001)
	) name2711 (
		_w13220_,
		_w13221_,
		_w13222_,
		_w13223_,
		_w13224_
	);
	LUT4 #(
		.INIT('h8000)
	) name2712 (
		_w13209_,
		_w13214_,
		_w13219_,
		_w13224_,
		_w13225_
	);
	LUT4 #(
		.INIT('h8000)
	) name2713 (
		_w13162_,
		_w13183_,
		_w13204_,
		_w13225_,
		_w13226_
	);
	LUT3 #(
		.INIT('h80)
	) name2714 (
		\wishbone_bd_ram_mem3_reg[153][24]/P0001 ,
		_w11959_,
		_w11968_,
		_w13227_
	);
	LUT3 #(
		.INIT('h80)
	) name2715 (
		\wishbone_bd_ram_mem3_reg[44][24]/P0001 ,
		_w11954_,
		_w11957_,
		_w13228_
	);
	LUT3 #(
		.INIT('h80)
	) name2716 (
		\wishbone_bd_ram_mem3_reg[191][24]/P0001 ,
		_w11942_,
		_w11973_,
		_w13229_
	);
	LUT3 #(
		.INIT('h80)
	) name2717 (
		\wishbone_bd_ram_mem3_reg[217][24]/P0001 ,
		_w11968_,
		_w11984_,
		_w13230_
	);
	LUT4 #(
		.INIT('h0001)
	) name2718 (
		_w13227_,
		_w13228_,
		_w13229_,
		_w13230_,
		_w13231_
	);
	LUT3 #(
		.INIT('h80)
	) name2719 (
		\wishbone_bd_ram_mem3_reg[68][24]/P0001 ,
		_w11929_,
		_w11949_,
		_w13232_
	);
	LUT3 #(
		.INIT('h80)
	) name2720 (
		\wishbone_bd_ram_mem3_reg[38][24]/P0001 ,
		_w11957_,
		_w11986_,
		_w13233_
	);
	LUT3 #(
		.INIT('h80)
	) name2721 (
		\wishbone_bd_ram_mem3_reg[233][24]/P0001 ,
		_w11968_,
		_w11982_,
		_w13234_
	);
	LUT3 #(
		.INIT('h80)
	) name2722 (
		\wishbone_bd_ram_mem3_reg[117][24]/P0001 ,
		_w11933_,
		_w12012_,
		_w13235_
	);
	LUT4 #(
		.INIT('h0001)
	) name2723 (
		_w13232_,
		_w13233_,
		_w13234_,
		_w13235_,
		_w13236_
	);
	LUT3 #(
		.INIT('h80)
	) name2724 (
		\wishbone_bd_ram_mem3_reg[189][24]/P0001 ,
		_w11942_,
		_w11966_,
		_w13237_
	);
	LUT3 #(
		.INIT('h80)
	) name2725 (
		\wishbone_bd_ram_mem3_reg[180][24]/P0001 ,
		_w11929_,
		_w11942_,
		_w13238_
	);
	LUT3 #(
		.INIT('h80)
	) name2726 (
		\wishbone_bd_ram_mem3_reg[243][24]/P0001 ,
		_w11938_,
		_w11952_,
		_w13239_
	);
	LUT3 #(
		.INIT('h80)
	) name2727 (
		\wishbone_bd_ram_mem3_reg[116][24]/P0001 ,
		_w11929_,
		_w12012_,
		_w13240_
	);
	LUT4 #(
		.INIT('h0001)
	) name2728 (
		_w13237_,
		_w13238_,
		_w13239_,
		_w13240_,
		_w13241_
	);
	LUT3 #(
		.INIT('h80)
	) name2729 (
		\wishbone_bd_ram_mem3_reg[77][24]/P0001 ,
		_w11949_,
		_w11966_,
		_w13242_
	);
	LUT3 #(
		.INIT('h80)
	) name2730 (
		\wishbone_bd_ram_mem3_reg[125][24]/P0001 ,
		_w11966_,
		_w12012_,
		_w13243_
	);
	LUT3 #(
		.INIT('h80)
	) name2731 (
		\wishbone_bd_ram_mem3_reg[237][24]/P0001 ,
		_w11966_,
		_w11982_,
		_w13244_
	);
	LUT3 #(
		.INIT('h80)
	) name2732 (
		\wishbone_bd_ram_mem3_reg[195][24]/P0001 ,
		_w11938_,
		_w11945_,
		_w13245_
	);
	LUT4 #(
		.INIT('h0001)
	) name2733 (
		_w13242_,
		_w13243_,
		_w13244_,
		_w13245_,
		_w13246_
	);
	LUT4 #(
		.INIT('h8000)
	) name2734 (
		_w13231_,
		_w13236_,
		_w13241_,
		_w13246_,
		_w13247_
	);
	LUT3 #(
		.INIT('h80)
	) name2735 (
		\wishbone_bd_ram_mem3_reg[214][24]/P0001 ,
		_w11984_,
		_w11986_,
		_w13248_
	);
	LUT3 #(
		.INIT('h80)
	) name2736 (
		\wishbone_bd_ram_mem3_reg[177][24]/P0001 ,
		_w11942_,
		_w11977_,
		_w13249_
	);
	LUT3 #(
		.INIT('h80)
	) name2737 (
		\wishbone_bd_ram_mem3_reg[166][24]/P0001 ,
		_w11930_,
		_w11986_,
		_w13250_
	);
	LUT3 #(
		.INIT('h80)
	) name2738 (
		\wishbone_bd_ram_mem3_reg[102][24]/P0001 ,
		_w11965_,
		_w11986_,
		_w13251_
	);
	LUT4 #(
		.INIT('h0001)
	) name2739 (
		_w13248_,
		_w13249_,
		_w13250_,
		_w13251_,
		_w13252_
	);
	LUT3 #(
		.INIT('h80)
	) name2740 (
		\wishbone_bd_ram_mem3_reg[238][24]/P0001 ,
		_w11948_,
		_w11982_,
		_w13253_
	);
	LUT3 #(
		.INIT('h80)
	) name2741 (
		\wishbone_bd_ram_mem3_reg[124][24]/P0001 ,
		_w11954_,
		_w12012_,
		_w13254_
	);
	LUT3 #(
		.INIT('h80)
	) name2742 (
		\wishbone_bd_ram_mem3_reg[234][24]/P0001 ,
		_w11944_,
		_w11982_,
		_w13255_
	);
	LUT3 #(
		.INIT('h80)
	) name2743 (
		\wishbone_bd_ram_mem3_reg[232][24]/P0001 ,
		_w11982_,
		_w11990_,
		_w13256_
	);
	LUT4 #(
		.INIT('h0001)
	) name2744 (
		_w13253_,
		_w13254_,
		_w13255_,
		_w13256_,
		_w13257_
	);
	LUT3 #(
		.INIT('h80)
	) name2745 (
		\wishbone_bd_ram_mem3_reg[118][24]/P0001 ,
		_w11986_,
		_w12012_,
		_w13258_
	);
	LUT3 #(
		.INIT('h80)
	) name2746 (
		\wishbone_bd_ram_mem3_reg[50][24]/P0001 ,
		_w11963_,
		_w11979_,
		_w13259_
	);
	LUT3 #(
		.INIT('h80)
	) name2747 (
		\wishbone_bd_ram_mem3_reg[81][24]/P0001 ,
		_w11972_,
		_w11977_,
		_w13260_
	);
	LUT3 #(
		.INIT('h80)
	) name2748 (
		\wishbone_bd_ram_mem3_reg[82][24]/P0001 ,
		_w11963_,
		_w11972_,
		_w13261_
	);
	LUT4 #(
		.INIT('h0001)
	) name2749 (
		_w13258_,
		_w13259_,
		_w13260_,
		_w13261_,
		_w13262_
	);
	LUT3 #(
		.INIT('h80)
	) name2750 (
		\wishbone_bd_ram_mem3_reg[11][24]/P0001 ,
		_w11932_,
		_w11936_,
		_w13263_
	);
	LUT3 #(
		.INIT('h80)
	) name2751 (
		\wishbone_bd_ram_mem3_reg[53][24]/P0001 ,
		_w11933_,
		_w11979_,
		_w13264_
	);
	LUT3 #(
		.INIT('h80)
	) name2752 (
		\wishbone_bd_ram_mem3_reg[169][24]/P0001 ,
		_w11930_,
		_w11968_,
		_w13265_
	);
	LUT3 #(
		.INIT('h80)
	) name2753 (
		\wishbone_bd_ram_mem3_reg[59][24]/P0001 ,
		_w11936_,
		_w11979_,
		_w13266_
	);
	LUT4 #(
		.INIT('h0001)
	) name2754 (
		_w13263_,
		_w13264_,
		_w13265_,
		_w13266_,
		_w13267_
	);
	LUT4 #(
		.INIT('h8000)
	) name2755 (
		_w13252_,
		_w13257_,
		_w13262_,
		_w13267_,
		_w13268_
	);
	LUT3 #(
		.INIT('h80)
	) name2756 (
		\wishbone_bd_ram_mem3_reg[213][24]/P0001 ,
		_w11933_,
		_w11984_,
		_w13269_
	);
	LUT3 #(
		.INIT('h80)
	) name2757 (
		\wishbone_bd_ram_mem3_reg[76][24]/P0001 ,
		_w11949_,
		_w11954_,
		_w13270_
	);
	LUT3 #(
		.INIT('h80)
	) name2758 (
		\wishbone_bd_ram_mem3_reg[16][24]/P0001 ,
		_w11935_,
		_w11941_,
		_w13271_
	);
	LUT3 #(
		.INIT('h80)
	) name2759 (
		\wishbone_bd_ram_mem3_reg[175][24]/P0001 ,
		_w11930_,
		_w11973_,
		_w13272_
	);
	LUT4 #(
		.INIT('h0001)
	) name2760 (
		_w13269_,
		_w13270_,
		_w13271_,
		_w13272_,
		_w13273_
	);
	LUT3 #(
		.INIT('h80)
	) name2761 (
		\wishbone_bd_ram_mem3_reg[253][24]/P0001 ,
		_w11952_,
		_w11966_,
		_w13274_
	);
	LUT3 #(
		.INIT('h80)
	) name2762 (
		\wishbone_bd_ram_mem3_reg[62][24]/P0001 ,
		_w11948_,
		_w11979_,
		_w13275_
	);
	LUT3 #(
		.INIT('h80)
	) name2763 (
		\wishbone_bd_ram_mem3_reg[122][24]/P0001 ,
		_w11944_,
		_w12012_,
		_w13276_
	);
	LUT3 #(
		.INIT('h80)
	) name2764 (
		\wishbone_bd_ram_mem3_reg[6][24]/P0001 ,
		_w11932_,
		_w11986_,
		_w13277_
	);
	LUT4 #(
		.INIT('h0001)
	) name2765 (
		_w13274_,
		_w13275_,
		_w13276_,
		_w13277_,
		_w13278_
	);
	LUT3 #(
		.INIT('h80)
	) name2766 (
		\wishbone_bd_ram_mem3_reg[13][24]/P0001 ,
		_w11932_,
		_w11966_,
		_w13279_
	);
	LUT3 #(
		.INIT('h80)
	) name2767 (
		\wishbone_bd_ram_mem3_reg[193][24]/P0001 ,
		_w11945_,
		_w11977_,
		_w13280_
	);
	LUT3 #(
		.INIT('h80)
	) name2768 (
		\wishbone_bd_ram_mem3_reg[4][24]/P0001 ,
		_w11929_,
		_w11932_,
		_w13281_
	);
	LUT3 #(
		.INIT('h80)
	) name2769 (
		\wishbone_bd_ram_mem3_reg[236][24]/P0001 ,
		_w11954_,
		_w11982_,
		_w13282_
	);
	LUT4 #(
		.INIT('h0001)
	) name2770 (
		_w13279_,
		_w13280_,
		_w13281_,
		_w13282_,
		_w13283_
	);
	LUT3 #(
		.INIT('h80)
	) name2771 (
		\wishbone_bd_ram_mem3_reg[27][24]/P0001 ,
		_w11935_,
		_w11936_,
		_w13284_
	);
	LUT3 #(
		.INIT('h80)
	) name2772 (
		\wishbone_bd_ram_mem3_reg[159][24]/P0001 ,
		_w11959_,
		_w11973_,
		_w13285_
	);
	LUT3 #(
		.INIT('h80)
	) name2773 (
		\wishbone_bd_ram_mem3_reg[32][24]/P0001 ,
		_w11941_,
		_w11957_,
		_w13286_
	);
	LUT3 #(
		.INIT('h80)
	) name2774 (
		\wishbone_bd_ram_mem3_reg[14][24]/P0001 ,
		_w11932_,
		_w11948_,
		_w13287_
	);
	LUT4 #(
		.INIT('h0001)
	) name2775 (
		_w13284_,
		_w13285_,
		_w13286_,
		_w13287_,
		_w13288_
	);
	LUT4 #(
		.INIT('h8000)
	) name2776 (
		_w13273_,
		_w13278_,
		_w13283_,
		_w13288_,
		_w13289_
	);
	LUT3 #(
		.INIT('h80)
	) name2777 (
		\wishbone_bd_ram_mem3_reg[128][24]/P0001 ,
		_w11941_,
		_w11955_,
		_w13290_
	);
	LUT3 #(
		.INIT('h80)
	) name2778 (
		\wishbone_bd_ram_mem3_reg[113][24]/P0001 ,
		_w11977_,
		_w12012_,
		_w13291_
	);
	LUT3 #(
		.INIT('h80)
	) name2779 (
		\wishbone_bd_ram_mem3_reg[123][24]/P0001 ,
		_w11936_,
		_w12012_,
		_w13292_
	);
	LUT3 #(
		.INIT('h80)
	) name2780 (
		\wishbone_bd_ram_mem3_reg[206][24]/P0001 ,
		_w11945_,
		_w11948_,
		_w13293_
	);
	LUT4 #(
		.INIT('h0001)
	) name2781 (
		_w13290_,
		_w13291_,
		_w13292_,
		_w13293_,
		_w13294_
	);
	LUT3 #(
		.INIT('h80)
	) name2782 (
		\wishbone_bd_ram_mem3_reg[174][24]/P0001 ,
		_w11930_,
		_w11948_,
		_w13295_
	);
	LUT3 #(
		.INIT('h80)
	) name2783 (
		\wishbone_bd_ram_mem3_reg[242][24]/P0001 ,
		_w11952_,
		_w11963_,
		_w13296_
	);
	LUT3 #(
		.INIT('h80)
	) name2784 (
		\wishbone_bd_ram_mem3_reg[194][24]/P0001 ,
		_w11945_,
		_w11963_,
		_w13297_
	);
	LUT3 #(
		.INIT('h80)
	) name2785 (
		\wishbone_bd_ram_mem3_reg[223][24]/P0001 ,
		_w11973_,
		_w11984_,
		_w13298_
	);
	LUT4 #(
		.INIT('h0001)
	) name2786 (
		_w13295_,
		_w13296_,
		_w13297_,
		_w13298_,
		_w13299_
	);
	LUT3 #(
		.INIT('h80)
	) name2787 (
		\wishbone_bd_ram_mem3_reg[221][24]/P0001 ,
		_w11966_,
		_w11984_,
		_w13300_
	);
	LUT3 #(
		.INIT('h80)
	) name2788 (
		\wishbone_bd_ram_mem3_reg[85][24]/P0001 ,
		_w11933_,
		_w11972_,
		_w13301_
	);
	LUT3 #(
		.INIT('h80)
	) name2789 (
		\wishbone_bd_ram_mem3_reg[63][24]/P0001 ,
		_w11973_,
		_w11979_,
		_w13302_
	);
	LUT3 #(
		.INIT('h80)
	) name2790 (
		\wishbone_bd_ram_mem3_reg[71][24]/P0001 ,
		_w11949_,
		_w11975_,
		_w13303_
	);
	LUT4 #(
		.INIT('h0001)
	) name2791 (
		_w13300_,
		_w13301_,
		_w13302_,
		_w13303_,
		_w13304_
	);
	LUT3 #(
		.INIT('h80)
	) name2792 (
		\wishbone_bd_ram_mem3_reg[74][24]/P0001 ,
		_w11944_,
		_w11949_,
		_w13305_
	);
	LUT3 #(
		.INIT('h80)
	) name2793 (
		\wishbone_bd_ram_mem3_reg[56][24]/P0001 ,
		_w11979_,
		_w11990_,
		_w13306_
	);
	LUT3 #(
		.INIT('h80)
	) name2794 (
		\wishbone_bd_ram_mem3_reg[95][24]/P0001 ,
		_w11972_,
		_w11973_,
		_w13307_
	);
	LUT3 #(
		.INIT('h80)
	) name2795 (
		\wishbone_bd_ram_mem3_reg[49][24]/P0001 ,
		_w11977_,
		_w11979_,
		_w13308_
	);
	LUT4 #(
		.INIT('h0001)
	) name2796 (
		_w13305_,
		_w13306_,
		_w13307_,
		_w13308_,
		_w13309_
	);
	LUT4 #(
		.INIT('h8000)
	) name2797 (
		_w13294_,
		_w13299_,
		_w13304_,
		_w13309_,
		_w13310_
	);
	LUT4 #(
		.INIT('h8000)
	) name2798 (
		_w13247_,
		_w13268_,
		_w13289_,
		_w13310_,
		_w13311_
	);
	LUT3 #(
		.INIT('h80)
	) name2799 (
		\wishbone_bd_ram_mem3_reg[37][24]/P0001 ,
		_w11933_,
		_w11957_,
		_w13312_
	);
	LUT3 #(
		.INIT('h80)
	) name2800 (
		\wishbone_bd_ram_mem3_reg[222][24]/P0001 ,
		_w11948_,
		_w11984_,
		_w13313_
	);
	LUT3 #(
		.INIT('h80)
	) name2801 (
		\wishbone_bd_ram_mem3_reg[92][24]/P0001 ,
		_w11954_,
		_w11972_,
		_w13314_
	);
	LUT3 #(
		.INIT('h80)
	) name2802 (
		\wishbone_bd_ram_mem3_reg[208][24]/P0001 ,
		_w11941_,
		_w11984_,
		_w13315_
	);
	LUT4 #(
		.INIT('h0001)
	) name2803 (
		_w13312_,
		_w13313_,
		_w13314_,
		_w13315_,
		_w13316_
	);
	LUT3 #(
		.INIT('h80)
	) name2804 (
		\wishbone_bd_ram_mem3_reg[231][24]/P0001 ,
		_w11975_,
		_w11982_,
		_w13317_
	);
	LUT3 #(
		.INIT('h80)
	) name2805 (
		\wishbone_bd_ram_mem3_reg[48][24]/P0001 ,
		_w11941_,
		_w11979_,
		_w13318_
	);
	LUT3 #(
		.INIT('h80)
	) name2806 (
		\wishbone_bd_ram_mem3_reg[12][24]/P0001 ,
		_w11932_,
		_w11954_,
		_w13319_
	);
	LUT3 #(
		.INIT('h80)
	) name2807 (
		\wishbone_bd_ram_mem3_reg[240][24]/P0001 ,
		_w11941_,
		_w11952_,
		_w13320_
	);
	LUT4 #(
		.INIT('h0001)
	) name2808 (
		_w13317_,
		_w13318_,
		_w13319_,
		_w13320_,
		_w13321_
	);
	LUT3 #(
		.INIT('h80)
	) name2809 (
		\wishbone_bd_ram_mem3_reg[138][24]/P0001 ,
		_w11944_,
		_w11955_,
		_w13322_
	);
	LUT3 #(
		.INIT('h80)
	) name2810 (
		\wishbone_bd_ram_mem3_reg[246][24]/P0001 ,
		_w11952_,
		_w11986_,
		_w13323_
	);
	LUT3 #(
		.INIT('h80)
	) name2811 (
		\wishbone_bd_ram_mem3_reg[210][24]/P0001 ,
		_w11963_,
		_w11984_,
		_w13324_
	);
	LUT3 #(
		.INIT('h80)
	) name2812 (
		\wishbone_bd_ram_mem3_reg[107][24]/P0001 ,
		_w11936_,
		_w11965_,
		_w13325_
	);
	LUT4 #(
		.INIT('h0001)
	) name2813 (
		_w13322_,
		_w13323_,
		_w13324_,
		_w13325_,
		_w13326_
	);
	LUT3 #(
		.INIT('h80)
	) name2814 (
		\wishbone_bd_ram_mem3_reg[51][24]/P0001 ,
		_w11938_,
		_w11979_,
		_w13327_
	);
	LUT3 #(
		.INIT('h80)
	) name2815 (
		\wishbone_bd_ram_mem3_reg[5][24]/P0001 ,
		_w11932_,
		_w11933_,
		_w13328_
	);
	LUT3 #(
		.INIT('h80)
	) name2816 (
		\wishbone_bd_ram_mem3_reg[155][24]/P0001 ,
		_w11936_,
		_w11959_,
		_w13329_
	);
	LUT3 #(
		.INIT('h80)
	) name2817 (
		\wishbone_bd_ram_mem3_reg[72][24]/P0001 ,
		_w11949_,
		_w11990_,
		_w13330_
	);
	LUT4 #(
		.INIT('h0001)
	) name2818 (
		_w13327_,
		_w13328_,
		_w13329_,
		_w13330_,
		_w13331_
	);
	LUT4 #(
		.INIT('h8000)
	) name2819 (
		_w13316_,
		_w13321_,
		_w13326_,
		_w13331_,
		_w13332_
	);
	LUT3 #(
		.INIT('h80)
	) name2820 (
		\wishbone_bd_ram_mem3_reg[98][24]/P0001 ,
		_w11963_,
		_w11965_,
		_w13333_
	);
	LUT3 #(
		.INIT('h80)
	) name2821 (
		\wishbone_bd_ram_mem3_reg[45][24]/P0001 ,
		_w11957_,
		_w11966_,
		_w13334_
	);
	LUT3 #(
		.INIT('h80)
	) name2822 (
		\wishbone_bd_ram_mem3_reg[86][24]/P0001 ,
		_w11972_,
		_w11986_,
		_w13335_
	);
	LUT3 #(
		.INIT('h80)
	) name2823 (
		\wishbone_bd_ram_mem3_reg[64][24]/P0001 ,
		_w11941_,
		_w11949_,
		_w13336_
	);
	LUT4 #(
		.INIT('h0001)
	) name2824 (
		_w13333_,
		_w13334_,
		_w13335_,
		_w13336_,
		_w13337_
	);
	LUT3 #(
		.INIT('h80)
	) name2825 (
		\wishbone_bd_ram_mem3_reg[108][24]/P0001 ,
		_w11954_,
		_w11965_,
		_w13338_
	);
	LUT3 #(
		.INIT('h80)
	) name2826 (
		\wishbone_bd_ram_mem3_reg[19][24]/P0001 ,
		_w11935_,
		_w11938_,
		_w13339_
	);
	LUT3 #(
		.INIT('h80)
	) name2827 (
		\wishbone_bd_ram_mem3_reg[15][24]/P0001 ,
		_w11932_,
		_w11973_,
		_w13340_
	);
	LUT3 #(
		.INIT('h80)
	) name2828 (
		\wishbone_bd_ram_mem3_reg[23][24]/P0001 ,
		_w11935_,
		_w11975_,
		_w13341_
	);
	LUT4 #(
		.INIT('h0001)
	) name2829 (
		_w13338_,
		_w13339_,
		_w13340_,
		_w13341_,
		_w13342_
	);
	LUT3 #(
		.INIT('h80)
	) name2830 (
		\wishbone_bd_ram_mem3_reg[179][24]/P0001 ,
		_w11938_,
		_w11942_,
		_w13343_
	);
	LUT3 #(
		.INIT('h80)
	) name2831 (
		\wishbone_bd_ram_mem3_reg[167][24]/P0001 ,
		_w11930_,
		_w11975_,
		_w13344_
	);
	LUT3 #(
		.INIT('h80)
	) name2832 (
		\wishbone_bd_ram_mem3_reg[202][24]/P0001 ,
		_w11944_,
		_w11945_,
		_w13345_
	);
	LUT3 #(
		.INIT('h80)
	) name2833 (
		\wishbone_bd_ram_mem3_reg[119][24]/P0001 ,
		_w11975_,
		_w12012_,
		_w13346_
	);
	LUT4 #(
		.INIT('h0001)
	) name2834 (
		_w13343_,
		_w13344_,
		_w13345_,
		_w13346_,
		_w13347_
	);
	LUT3 #(
		.INIT('h80)
	) name2835 (
		\wishbone_bd_ram_mem3_reg[183][24]/P0001 ,
		_w11942_,
		_w11975_,
		_w13348_
	);
	LUT3 #(
		.INIT('h80)
	) name2836 (
		\wishbone_bd_ram_mem3_reg[161][24]/P0001 ,
		_w11930_,
		_w11977_,
		_w13349_
	);
	LUT3 #(
		.INIT('h80)
	) name2837 (
		\wishbone_bd_ram_mem3_reg[190][24]/P0001 ,
		_w11942_,
		_w11948_,
		_w13350_
	);
	LUT3 #(
		.INIT('h80)
	) name2838 (
		\wishbone_bd_ram_mem3_reg[54][24]/P0001 ,
		_w11979_,
		_w11986_,
		_w13351_
	);
	LUT4 #(
		.INIT('h0001)
	) name2839 (
		_w13348_,
		_w13349_,
		_w13350_,
		_w13351_,
		_w13352_
	);
	LUT4 #(
		.INIT('h8000)
	) name2840 (
		_w13337_,
		_w13342_,
		_w13347_,
		_w13352_,
		_w13353_
	);
	LUT3 #(
		.INIT('h80)
	) name2841 (
		\wishbone_bd_ram_mem3_reg[235][24]/P0001 ,
		_w11936_,
		_w11982_,
		_w13354_
	);
	LUT3 #(
		.INIT('h80)
	) name2842 (
		\wishbone_bd_ram_mem3_reg[42][24]/P0001 ,
		_w11944_,
		_w11957_,
		_w13355_
	);
	LUT3 #(
		.INIT('h80)
	) name2843 (
		\wishbone_bd_ram_mem3_reg[200][24]/P0001 ,
		_w11945_,
		_w11990_,
		_w13356_
	);
	LUT3 #(
		.INIT('h80)
	) name2844 (
		\wishbone_bd_ram_mem3_reg[112][24]/P0001 ,
		_w11941_,
		_w12012_,
		_w13357_
	);
	LUT4 #(
		.INIT('h0001)
	) name2845 (
		_w13354_,
		_w13355_,
		_w13356_,
		_w13357_,
		_w13358_
	);
	LUT3 #(
		.INIT('h80)
	) name2846 (
		\wishbone_bd_ram_mem3_reg[148][24]/P0001 ,
		_w11929_,
		_w11959_,
		_w13359_
	);
	LUT3 #(
		.INIT('h80)
	) name2847 (
		\wishbone_bd_ram_mem3_reg[134][24]/P0001 ,
		_w11955_,
		_w11986_,
		_w13360_
	);
	LUT3 #(
		.INIT('h80)
	) name2848 (
		\wishbone_bd_ram_mem3_reg[163][24]/P0001 ,
		_w11930_,
		_w11938_,
		_w13361_
	);
	LUT3 #(
		.INIT('h80)
	) name2849 (
		\wishbone_bd_ram_mem3_reg[186][24]/P0001 ,
		_w11942_,
		_w11944_,
		_w13362_
	);
	LUT4 #(
		.INIT('h0001)
	) name2850 (
		_w13359_,
		_w13360_,
		_w13361_,
		_w13362_,
		_w13363_
	);
	LUT3 #(
		.INIT('h80)
	) name2851 (
		\wishbone_bd_ram_mem3_reg[69][24]/P0001 ,
		_w11933_,
		_w11949_,
		_w13364_
	);
	LUT3 #(
		.INIT('h80)
	) name2852 (
		\wishbone_bd_ram_mem3_reg[225][24]/P0001 ,
		_w11977_,
		_w11982_,
		_w13365_
	);
	LUT3 #(
		.INIT('h80)
	) name2853 (
		\wishbone_bd_ram_mem3_reg[1][24]/P0001 ,
		_w11932_,
		_w11977_,
		_w13366_
	);
	LUT3 #(
		.INIT('h80)
	) name2854 (
		\wishbone_bd_ram_mem3_reg[70][24]/P0001 ,
		_w11949_,
		_w11986_,
		_w13367_
	);
	LUT4 #(
		.INIT('h0001)
	) name2855 (
		_w13364_,
		_w13365_,
		_w13366_,
		_w13367_,
		_w13368_
	);
	LUT3 #(
		.INIT('h80)
	) name2856 (
		\wishbone_bd_ram_mem3_reg[251][24]/P0001 ,
		_w11936_,
		_w11952_,
		_w13369_
	);
	LUT3 #(
		.INIT('h80)
	) name2857 (
		\wishbone_bd_ram_mem3_reg[151][24]/P0001 ,
		_w11959_,
		_w11975_,
		_w13370_
	);
	LUT3 #(
		.INIT('h80)
	) name2858 (
		\wishbone_bd_ram_mem3_reg[254][24]/P0001 ,
		_w11948_,
		_w11952_,
		_w13371_
	);
	LUT3 #(
		.INIT('h80)
	) name2859 (
		\wishbone_bd_ram_mem3_reg[103][24]/P0001 ,
		_w11965_,
		_w11975_,
		_w13372_
	);
	LUT4 #(
		.INIT('h0001)
	) name2860 (
		_w13369_,
		_w13370_,
		_w13371_,
		_w13372_,
		_w13373_
	);
	LUT4 #(
		.INIT('h8000)
	) name2861 (
		_w13358_,
		_w13363_,
		_w13368_,
		_w13373_,
		_w13374_
	);
	LUT3 #(
		.INIT('h80)
	) name2862 (
		\wishbone_bd_ram_mem3_reg[79][24]/P0001 ,
		_w11949_,
		_w11973_,
		_w13375_
	);
	LUT3 #(
		.INIT('h80)
	) name2863 (
		\wishbone_bd_ram_mem3_reg[101][24]/P0001 ,
		_w11933_,
		_w11965_,
		_w13376_
	);
	LUT3 #(
		.INIT('h80)
	) name2864 (
		\wishbone_bd_ram_mem3_reg[199][24]/P0001 ,
		_w11945_,
		_w11975_,
		_w13377_
	);
	LUT3 #(
		.INIT('h80)
	) name2865 (
		\wishbone_bd_ram_mem3_reg[58][24]/P0001 ,
		_w11944_,
		_w11979_,
		_w13378_
	);
	LUT4 #(
		.INIT('h0001)
	) name2866 (
		_w13375_,
		_w13376_,
		_w13377_,
		_w13378_,
		_w13379_
	);
	LUT3 #(
		.INIT('h80)
	) name2867 (
		\wishbone_bd_ram_mem3_reg[136][24]/P0001 ,
		_w11955_,
		_w11990_,
		_w13380_
	);
	LUT3 #(
		.INIT('h80)
	) name2868 (
		\wishbone_bd_ram_mem3_reg[135][24]/P0001 ,
		_w11955_,
		_w11975_,
		_w13381_
	);
	LUT3 #(
		.INIT('h80)
	) name2869 (
		\wishbone_bd_ram_mem3_reg[87][24]/P0001 ,
		_w11972_,
		_w11975_,
		_w13382_
	);
	LUT3 #(
		.INIT('h80)
	) name2870 (
		\wishbone_bd_ram_mem3_reg[156][24]/P0001 ,
		_w11954_,
		_w11959_,
		_w13383_
	);
	LUT4 #(
		.INIT('h0001)
	) name2871 (
		_w13380_,
		_w13381_,
		_w13382_,
		_w13383_,
		_w13384_
	);
	LUT3 #(
		.INIT('h80)
	) name2872 (
		\wishbone_bd_ram_mem3_reg[207][24]/P0001 ,
		_w11945_,
		_w11973_,
		_w13385_
	);
	LUT3 #(
		.INIT('h80)
	) name2873 (
		\wishbone_bd_ram_mem3_reg[248][24]/P0001 ,
		_w11952_,
		_w11990_,
		_w13386_
	);
	LUT3 #(
		.INIT('h80)
	) name2874 (
		\wishbone_bd_ram_mem3_reg[94][24]/P0001 ,
		_w11948_,
		_w11972_,
		_w13387_
	);
	LUT3 #(
		.INIT('h80)
	) name2875 (
		\wishbone_bd_ram_mem3_reg[7][24]/P0001 ,
		_w11932_,
		_w11975_,
		_w13388_
	);
	LUT4 #(
		.INIT('h0001)
	) name2876 (
		_w13385_,
		_w13386_,
		_w13387_,
		_w13388_,
		_w13389_
	);
	LUT3 #(
		.INIT('h80)
	) name2877 (
		\wishbone_bd_ram_mem3_reg[198][24]/P0001 ,
		_w11945_,
		_w11986_,
		_w13390_
	);
	LUT3 #(
		.INIT('h80)
	) name2878 (
		\wishbone_bd_ram_mem3_reg[46][24]/P0001 ,
		_w11948_,
		_w11957_,
		_w13391_
	);
	LUT3 #(
		.INIT('h80)
	) name2879 (
		\wishbone_bd_ram_mem3_reg[96][24]/P0001 ,
		_w11941_,
		_w11965_,
		_w13392_
	);
	LUT3 #(
		.INIT('h80)
	) name2880 (
		\wishbone_bd_ram_mem3_reg[203][24]/P0001 ,
		_w11936_,
		_w11945_,
		_w13393_
	);
	LUT4 #(
		.INIT('h0001)
	) name2881 (
		_w13390_,
		_w13391_,
		_w13392_,
		_w13393_,
		_w13394_
	);
	LUT4 #(
		.INIT('h8000)
	) name2882 (
		_w13379_,
		_w13384_,
		_w13389_,
		_w13394_,
		_w13395_
	);
	LUT4 #(
		.INIT('h8000)
	) name2883 (
		_w13332_,
		_w13353_,
		_w13374_,
		_w13395_,
		_w13396_
	);
	LUT4 #(
		.INIT('h8000)
	) name2884 (
		_w13141_,
		_w13226_,
		_w13311_,
		_w13396_,
		_w13397_
	);
	LUT3 #(
		.INIT('h01)
	) name2885 (
		\wishbone_TxLength_reg[5]/NET0131 ,
		\wishbone_TxLength_reg[6]/NET0131 ,
		\wishbone_TxLength_reg[7]/NET0131 ,
		_w13398_
	);
	LUT4 #(
		.INIT('h0800)
	) name2886 (
		_w12304_,
		_w12309_,
		_w12323_,
		_w13398_,
		_w13399_
	);
	LUT4 #(
		.INIT('h4055)
	) name2887 (
		\wishbone_TxLength_reg[8]/NET0131 ,
		_w12312_,
		_w12317_,
		_w13399_,
		_w13400_
	);
	LUT3 #(
		.INIT('h20)
	) name2888 (
		_w12309_,
		_w12323_,
		_w13398_,
		_w13401_
	);
	LUT3 #(
		.INIT('h80)
	) name2889 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_TxLength_reg[8]/NET0131 ,
		_w13402_
	);
	LUT4 #(
		.INIT('hf800)
	) name2890 (
		_w12312_,
		_w12317_,
		_w13401_,
		_w13402_,
		_w13403_
	);
	LUT3 #(
		.INIT('h01)
	) name2891 (
		_w12302_,
		_w13400_,
		_w13403_,
		_w13404_
	);
	LUT3 #(
		.INIT('hf2)
	) name2892 (
		_w12303_,
		_w13397_,
		_w13404_,
		_w13405_
	);
	LUT2 #(
		.INIT('h8)
	) name2893 (
		_w11854_,
		_w11855_,
		_w13406_
	);
	LUT3 #(
		.INIT('h80)
	) name2894 (
		_w11851_,
		_w11852_,
		_w13406_,
		_w13407_
	);
	LUT4 #(
		.INIT('h8000)
	) name2895 (
		\m_wb_adr_o[25]_pad ,
		_w11851_,
		_w11852_,
		_w13406_,
		_w13408_
	);
	LUT2 #(
		.INIT('h1)
	) name2896 (
		\m_wb_adr_o[26]_pad ,
		_w13408_,
		_w13409_
	);
	LUT4 #(
		.INIT('h80aa)
	) name2897 (
		\wishbone_TxPointerMSB_reg[26]/NET0131 ,
		_w11866_,
		_w11867_,
		_w11883_,
		_w13410_
	);
	LUT2 #(
		.INIT('h4)
	) name2898 (
		_w11882_,
		_w13410_,
		_w13411_
	);
	LUT4 #(
		.INIT('h5554)
	) name2899 (
		_w11858_,
		_w11887_,
		_w13051_,
		_w13411_,
		_w13412_
	);
	LUT2 #(
		.INIT('h4)
	) name2900 (
		_w13409_,
		_w13412_,
		_w13413_
	);
	LUT3 #(
		.INIT('ha2)
	) name2901 (
		\wishbone_TxPointerMSB_reg[26]/NET0131 ,
		_w11900_,
		_w11909_,
		_w13414_
	);
	LUT4 #(
		.INIT('h080a)
	) name2902 (
		\wishbone_RxPointerMSB_reg[26]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w13415_
	);
	LUT3 #(
		.INIT('he0)
	) name2903 (
		_w11902_,
		_w11905_,
		_w13415_,
		_w13416_
	);
	LUT4 #(
		.INIT('h0007)
	) name2904 (
		\m_wb_adr_o[26]_pad ,
		_w11907_,
		_w13414_,
		_w13416_,
		_w13417_
	);
	LUT2 #(
		.INIT('hb)
	) name2905 (
		_w13413_,
		_w13417_,
		_w13418_
	);
	LUT2 #(
		.INIT('h8)
	) name2906 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w13419_
	);
	LUT4 #(
		.INIT('h8000)
	) name2907 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w13420_
	);
	LUT3 #(
		.INIT('h40)
	) name2908 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_RxEnableWindow_reg/NET0131 ,
		_w13421_
	);
	LUT3 #(
		.INIT('h80)
	) name2909 (
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		\wishbone_RxByteCnt_reg[1]/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w13422_
	);
	LUT4 #(
		.INIT('h0777)
	) name2910 (
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w13420_,
		_w13421_,
		_w13422_,
		_w13423_
	);
	LUT4 #(
		.INIT('h8000)
	) name2911 (
		\wishbone_LastByteIn_reg/NET0131 ,
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		\wishbone_RxByteCnt_reg[1]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w13424_
	);
	LUT2 #(
		.INIT('h2)
	) name2912 (
		\wishbone_RxDataLatched2_reg[10]/NET0131 ,
		_w13424_,
		_w13425_
	);
	LUT2 #(
		.INIT('h8)
	) name2913 (
		_w13423_,
		_w13425_,
		_w13426_
	);
	LUT2 #(
		.INIT('h6)
	) name2914 (
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		_w13427_
	);
	LUT3 #(
		.INIT('he0)
	) name2915 (
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w13423_,
		_w13427_,
		_w13428_
	);
	LUT2 #(
		.INIT('hd)
	) name2916 (
		_w13423_,
		_w13424_,
		_w13429_
	);
	LUT3 #(
		.INIT('ha2)
	) name2917 (
		\wishbone_RxDataLatched1_reg[10]/NET0131 ,
		_w13423_,
		_w13424_,
		_w13430_
	);
	LUT3 #(
		.INIT('hba)
	) name2918 (
		_w13426_,
		_w13428_,
		_w13430_,
		_w13431_
	);
	LUT2 #(
		.INIT('h2)
	) name2919 (
		\wishbone_RxDataLatched2_reg[11]/NET0131 ,
		_w13424_,
		_w13432_
	);
	LUT2 #(
		.INIT('h8)
	) name2920 (
		_w13423_,
		_w13432_,
		_w13433_
	);
	LUT3 #(
		.INIT('ha2)
	) name2921 (
		\wishbone_RxDataLatched1_reg[11]/NET0131 ,
		_w13423_,
		_w13424_,
		_w13434_
	);
	LUT3 #(
		.INIT('hdc)
	) name2922 (
		_w13428_,
		_w13433_,
		_w13434_,
		_w13435_
	);
	LUT2 #(
		.INIT('h2)
	) name2923 (
		\wishbone_RxDataLatched2_reg[12]/NET0131 ,
		_w13424_,
		_w13436_
	);
	LUT2 #(
		.INIT('h8)
	) name2924 (
		_w13423_,
		_w13436_,
		_w13437_
	);
	LUT3 #(
		.INIT('ha2)
	) name2925 (
		\wishbone_RxDataLatched1_reg[12]/NET0131 ,
		_w13423_,
		_w13424_,
		_w13438_
	);
	LUT3 #(
		.INIT('hdc)
	) name2926 (
		_w13428_,
		_w13437_,
		_w13438_,
		_w13439_
	);
	LUT2 #(
		.INIT('h2)
	) name2927 (
		\wishbone_RxDataLatched2_reg[13]/NET0131 ,
		_w13424_,
		_w13440_
	);
	LUT2 #(
		.INIT('h8)
	) name2928 (
		_w13423_,
		_w13440_,
		_w13441_
	);
	LUT3 #(
		.INIT('ha2)
	) name2929 (
		\wishbone_RxDataLatched1_reg[13]/NET0131 ,
		_w13423_,
		_w13424_,
		_w13442_
	);
	LUT3 #(
		.INIT('hdc)
	) name2930 (
		_w13428_,
		_w13441_,
		_w13442_,
		_w13443_
	);
	LUT2 #(
		.INIT('h2)
	) name2931 (
		\wishbone_RxDataLatched2_reg[14]/NET0131 ,
		_w13424_,
		_w13444_
	);
	LUT2 #(
		.INIT('h8)
	) name2932 (
		_w13423_,
		_w13444_,
		_w13445_
	);
	LUT3 #(
		.INIT('ha2)
	) name2933 (
		\wishbone_RxDataLatched1_reg[14]/NET0131 ,
		_w13423_,
		_w13424_,
		_w13446_
	);
	LUT3 #(
		.INIT('hdc)
	) name2934 (
		_w13428_,
		_w13445_,
		_w13446_,
		_w13447_
	);
	LUT2 #(
		.INIT('h2)
	) name2935 (
		\wishbone_RxDataLatched2_reg[15]/NET0131 ,
		_w13424_,
		_w13448_
	);
	LUT2 #(
		.INIT('h8)
	) name2936 (
		_w13423_,
		_w13448_,
		_w13449_
	);
	LUT3 #(
		.INIT('ha2)
	) name2937 (
		\wishbone_RxDataLatched1_reg[15]/NET0131 ,
		_w13423_,
		_w13424_,
		_w13450_
	);
	LUT3 #(
		.INIT('hdc)
	) name2938 (
		_w13428_,
		_w13449_,
		_w13450_,
		_w13451_
	);
	LUT2 #(
		.INIT('h2)
	) name2939 (
		\wishbone_RxDataLatched2_reg[8]/NET0131 ,
		_w13424_,
		_w13452_
	);
	LUT2 #(
		.INIT('h8)
	) name2940 (
		_w13423_,
		_w13452_,
		_w13453_
	);
	LUT3 #(
		.INIT('ha2)
	) name2941 (
		\wishbone_RxDataLatched1_reg[8]/NET0131 ,
		_w13423_,
		_w13424_,
		_w13454_
	);
	LUT3 #(
		.INIT('hdc)
	) name2942 (
		_w13428_,
		_w13453_,
		_w13454_,
		_w13455_
	);
	LUT3 #(
		.INIT('h80)
	) name2943 (
		\wishbone_RxBDRead_reg/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		_w13456_
	);
	LUT2 #(
		.INIT('h2)
	) name2944 (
		\wishbone_RxBDReady_reg/NET0131 ,
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w13457_
	);
	LUT4 #(
		.INIT('h0080)
	) name2945 (
		\wishbone_RxBDRead_reg/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w13458_
	);
	LUT3 #(
		.INIT('h54)
	) name2946 (
		_w13456_,
		_w13457_,
		_w13458_,
		_w13459_
	);
	LUT3 #(
		.INIT('h80)
	) name2947 (
		\wishbone_bd_ram_mem1_reg[44][15]/P0001 ,
		_w11954_,
		_w11957_,
		_w13460_
	);
	LUT3 #(
		.INIT('h80)
	) name2948 (
		\wishbone_bd_ram_mem1_reg[243][15]/P0001 ,
		_w11938_,
		_w11952_,
		_w13461_
	);
	LUT3 #(
		.INIT('h80)
	) name2949 (
		\wishbone_bd_ram_mem1_reg[118][15]/P0001 ,
		_w11986_,
		_w12012_,
		_w13462_
	);
	LUT3 #(
		.INIT('h80)
	) name2950 (
		\wishbone_bd_ram_mem1_reg[193][15]/P0001 ,
		_w11945_,
		_w11977_,
		_w13463_
	);
	LUT4 #(
		.INIT('h0001)
	) name2951 (
		_w13460_,
		_w13461_,
		_w13462_,
		_w13463_,
		_w13464_
	);
	LUT3 #(
		.INIT('h80)
	) name2952 (
		\wishbone_bd_ram_mem1_reg[234][15]/P0001 ,
		_w11944_,
		_w11982_,
		_w13465_
	);
	LUT3 #(
		.INIT('h80)
	) name2953 (
		\wishbone_bd_ram_mem1_reg[162][15]/P0001 ,
		_w11930_,
		_w11963_,
		_w13466_
	);
	LUT3 #(
		.INIT('h80)
	) name2954 (
		\wishbone_bd_ram_mem1_reg[145][15]/P0001 ,
		_w11959_,
		_w11977_,
		_w13467_
	);
	LUT3 #(
		.INIT('h80)
	) name2955 (
		\wishbone_bd_ram_mem1_reg[72][15]/P0001 ,
		_w11949_,
		_w11990_,
		_w13468_
	);
	LUT4 #(
		.INIT('h0001)
	) name2956 (
		_w13465_,
		_w13466_,
		_w13467_,
		_w13468_,
		_w13469_
	);
	LUT3 #(
		.INIT('h80)
	) name2957 (
		\wishbone_bd_ram_mem1_reg[105][15]/P0001 ,
		_w11965_,
		_w11968_,
		_w13470_
	);
	LUT3 #(
		.INIT('h80)
	) name2958 (
		\wishbone_bd_ram_mem1_reg[141][15]/P0001 ,
		_w11955_,
		_w11966_,
		_w13471_
	);
	LUT3 #(
		.INIT('h80)
	) name2959 (
		\wishbone_bd_ram_mem1_reg[149][15]/P0001 ,
		_w11933_,
		_w11959_,
		_w13472_
	);
	LUT3 #(
		.INIT('h80)
	) name2960 (
		\wishbone_bd_ram_mem1_reg[194][15]/P0001 ,
		_w11945_,
		_w11963_,
		_w13473_
	);
	LUT4 #(
		.INIT('h0001)
	) name2961 (
		_w13470_,
		_w13471_,
		_w13472_,
		_w13473_,
		_w13474_
	);
	LUT3 #(
		.INIT('h80)
	) name2962 (
		\wishbone_bd_ram_mem1_reg[132][15]/P0001 ,
		_w11929_,
		_w11955_,
		_w13475_
	);
	LUT3 #(
		.INIT('h80)
	) name2963 (
		\wishbone_bd_ram_mem1_reg[83][15]/P0001 ,
		_w11938_,
		_w11972_,
		_w13476_
	);
	LUT3 #(
		.INIT('h80)
	) name2964 (
		\wishbone_bd_ram_mem1_reg[167][15]/P0001 ,
		_w11930_,
		_w11975_,
		_w13477_
	);
	LUT3 #(
		.INIT('h80)
	) name2965 (
		\wishbone_bd_ram_mem1_reg[151][15]/P0001 ,
		_w11959_,
		_w11975_,
		_w13478_
	);
	LUT4 #(
		.INIT('h0001)
	) name2966 (
		_w13475_,
		_w13476_,
		_w13477_,
		_w13478_,
		_w13479_
	);
	LUT4 #(
		.INIT('h8000)
	) name2967 (
		_w13464_,
		_w13469_,
		_w13474_,
		_w13479_,
		_w13480_
	);
	LUT3 #(
		.INIT('h80)
	) name2968 (
		\wishbone_bd_ram_mem1_reg[47][15]/P0001 ,
		_w11957_,
		_w11973_,
		_w13481_
	);
	LUT3 #(
		.INIT('h80)
	) name2969 (
		\wishbone_bd_ram_mem1_reg[21][15]/P0001 ,
		_w11933_,
		_w11935_,
		_w13482_
	);
	LUT3 #(
		.INIT('h80)
	) name2970 (
		\wishbone_bd_ram_mem1_reg[77][15]/P0001 ,
		_w11949_,
		_w11966_,
		_w13483_
	);
	LUT3 #(
		.INIT('h80)
	) name2971 (
		\wishbone_bd_ram_mem1_reg[206][15]/P0001 ,
		_w11945_,
		_w11948_,
		_w13484_
	);
	LUT4 #(
		.INIT('h0001)
	) name2972 (
		_w13481_,
		_w13482_,
		_w13483_,
		_w13484_,
		_w13485_
	);
	LUT3 #(
		.INIT('h80)
	) name2973 (
		\wishbone_bd_ram_mem1_reg[15][15]/P0001 ,
		_w11932_,
		_w11973_,
		_w13486_
	);
	LUT3 #(
		.INIT('h80)
	) name2974 (
		\wishbone_bd_ram_mem1_reg[26][15]/P0001 ,
		_w11935_,
		_w11944_,
		_w13487_
	);
	LUT3 #(
		.INIT('h80)
	) name2975 (
		\wishbone_bd_ram_mem1_reg[97][15]/P0001 ,
		_w11965_,
		_w11977_,
		_w13488_
	);
	LUT3 #(
		.INIT('h80)
	) name2976 (
		\wishbone_bd_ram_mem1_reg[160][15]/P0001 ,
		_w11930_,
		_w11941_,
		_w13489_
	);
	LUT4 #(
		.INIT('h0001)
	) name2977 (
		_w13486_,
		_w13487_,
		_w13488_,
		_w13489_,
		_w13490_
	);
	LUT3 #(
		.INIT('h80)
	) name2978 (
		\wishbone_bd_ram_mem1_reg[4][15]/P0001 ,
		_w11929_,
		_w11932_,
		_w13491_
	);
	LUT3 #(
		.INIT('h80)
	) name2979 (
		\wishbone_bd_ram_mem1_reg[117][15]/P0001 ,
		_w11933_,
		_w12012_,
		_w13492_
	);
	LUT3 #(
		.INIT('h80)
	) name2980 (
		\wishbone_bd_ram_mem1_reg[152][15]/P0001 ,
		_w11959_,
		_w11990_,
		_w13493_
	);
	LUT3 #(
		.INIT('h80)
	) name2981 (
		\wishbone_bd_ram_mem1_reg[103][15]/P0001 ,
		_w11965_,
		_w11975_,
		_w13494_
	);
	LUT4 #(
		.INIT('h0001)
	) name2982 (
		_w13491_,
		_w13492_,
		_w13493_,
		_w13494_,
		_w13495_
	);
	LUT3 #(
		.INIT('h80)
	) name2983 (
		\wishbone_bd_ram_mem1_reg[153][15]/P0001 ,
		_w11959_,
		_w11968_,
		_w13496_
	);
	LUT3 #(
		.INIT('h80)
	) name2984 (
		\wishbone_bd_ram_mem1_reg[98][15]/P0001 ,
		_w11963_,
		_w11965_,
		_w13497_
	);
	LUT3 #(
		.INIT('h80)
	) name2985 (
		\wishbone_bd_ram_mem1_reg[192][15]/P0001 ,
		_w11941_,
		_w11945_,
		_w13498_
	);
	LUT3 #(
		.INIT('h80)
	) name2986 (
		\wishbone_bd_ram_mem1_reg[142][15]/P0001 ,
		_w11948_,
		_w11955_,
		_w13499_
	);
	LUT4 #(
		.INIT('h0001)
	) name2987 (
		_w13496_,
		_w13497_,
		_w13498_,
		_w13499_,
		_w13500_
	);
	LUT4 #(
		.INIT('h8000)
	) name2988 (
		_w13485_,
		_w13490_,
		_w13495_,
		_w13500_,
		_w13501_
	);
	LUT3 #(
		.INIT('h80)
	) name2989 (
		\wishbone_bd_ram_mem1_reg[50][15]/P0001 ,
		_w11963_,
		_w11979_,
		_w13502_
	);
	LUT3 #(
		.INIT('h80)
	) name2990 (
		\wishbone_bd_ram_mem1_reg[213][15]/P0001 ,
		_w11933_,
		_w11984_,
		_w13503_
	);
	LUT3 #(
		.INIT('h80)
	) name2991 (
		\wishbone_bd_ram_mem1_reg[32][15]/P0001 ,
		_w11941_,
		_w11957_,
		_w13504_
	);
	LUT3 #(
		.INIT('h80)
	) name2992 (
		\wishbone_bd_ram_mem1_reg[182][15]/P0001 ,
		_w11942_,
		_w11986_,
		_w13505_
	);
	LUT4 #(
		.INIT('h0001)
	) name2993 (
		_w13502_,
		_w13503_,
		_w13504_,
		_w13505_,
		_w13506_
	);
	LUT3 #(
		.INIT('h80)
	) name2994 (
		\wishbone_bd_ram_mem1_reg[29][15]/P0001 ,
		_w11935_,
		_w11966_,
		_w13507_
	);
	LUT3 #(
		.INIT('h80)
	) name2995 (
		\wishbone_bd_ram_mem1_reg[39][15]/P0001 ,
		_w11957_,
		_w11975_,
		_w13508_
	);
	LUT3 #(
		.INIT('h80)
	) name2996 (
		\wishbone_bd_ram_mem1_reg[134][15]/P0001 ,
		_w11955_,
		_w11986_,
		_w13509_
	);
	LUT3 #(
		.INIT('h80)
	) name2997 (
		\wishbone_bd_ram_mem1_reg[43][15]/P0001 ,
		_w11936_,
		_w11957_,
		_w13510_
	);
	LUT4 #(
		.INIT('h0001)
	) name2998 (
		_w13507_,
		_w13508_,
		_w13509_,
		_w13510_,
		_w13511_
	);
	LUT3 #(
		.INIT('h80)
	) name2999 (
		\wishbone_bd_ram_mem1_reg[13][15]/P0001 ,
		_w11932_,
		_w11966_,
		_w13512_
	);
	LUT3 #(
		.INIT('h80)
	) name3000 (
		\wishbone_bd_ram_mem1_reg[46][15]/P0001 ,
		_w11948_,
		_w11957_,
		_w13513_
	);
	LUT3 #(
		.INIT('h80)
	) name3001 (
		\wishbone_bd_ram_mem1_reg[101][15]/P0001 ,
		_w11933_,
		_w11965_,
		_w13514_
	);
	LUT3 #(
		.INIT('h80)
	) name3002 (
		\wishbone_bd_ram_mem1_reg[202][15]/P0001 ,
		_w11944_,
		_w11945_,
		_w13515_
	);
	LUT4 #(
		.INIT('h0001)
	) name3003 (
		_w13512_,
		_w13513_,
		_w13514_,
		_w13515_,
		_w13516_
	);
	LUT3 #(
		.INIT('h80)
	) name3004 (
		\wishbone_bd_ram_mem1_reg[163][15]/P0001 ,
		_w11930_,
		_w11938_,
		_w13517_
	);
	LUT3 #(
		.INIT('h80)
	) name3005 (
		\wishbone_bd_ram_mem1_reg[75][15]/P0001 ,
		_w11936_,
		_w11949_,
		_w13518_
	);
	LUT3 #(
		.INIT('h80)
	) name3006 (
		\wishbone_bd_ram_mem1_reg[9][15]/P0001 ,
		_w11932_,
		_w11968_,
		_w13519_
	);
	LUT3 #(
		.INIT('h80)
	) name3007 (
		\wishbone_bd_ram_mem1_reg[14][15]/P0001 ,
		_w11932_,
		_w11948_,
		_w13520_
	);
	LUT4 #(
		.INIT('h0001)
	) name3008 (
		_w13517_,
		_w13518_,
		_w13519_,
		_w13520_,
		_w13521_
	);
	LUT4 #(
		.INIT('h8000)
	) name3009 (
		_w13506_,
		_w13511_,
		_w13516_,
		_w13521_,
		_w13522_
	);
	LUT3 #(
		.INIT('h80)
	) name3010 (
		\wishbone_bd_ram_mem1_reg[218][15]/P0001 ,
		_w11944_,
		_w11984_,
		_w13523_
	);
	LUT3 #(
		.INIT('h80)
	) name3011 (
		\wishbone_bd_ram_mem1_reg[90][15]/P0001 ,
		_w11944_,
		_w11972_,
		_w13524_
	);
	LUT3 #(
		.INIT('h80)
	) name3012 (
		\wishbone_bd_ram_mem1_reg[126][15]/P0001 ,
		_w11948_,
		_w12012_,
		_w13525_
	);
	LUT3 #(
		.INIT('h80)
	) name3013 (
		\wishbone_bd_ram_mem1_reg[119][15]/P0001 ,
		_w11975_,
		_w12012_,
		_w13526_
	);
	LUT4 #(
		.INIT('h0001)
	) name3014 (
		_w13523_,
		_w13524_,
		_w13525_,
		_w13526_,
		_w13527_
	);
	LUT3 #(
		.INIT('h80)
	) name3015 (
		\wishbone_bd_ram_mem1_reg[109][15]/P0001 ,
		_w11965_,
		_w11966_,
		_w13528_
	);
	LUT3 #(
		.INIT('h80)
	) name3016 (
		\wishbone_bd_ram_mem1_reg[42][15]/P0001 ,
		_w11944_,
		_w11957_,
		_w13529_
	);
	LUT3 #(
		.INIT('h80)
	) name3017 (
		\wishbone_bd_ram_mem1_reg[144][15]/P0001 ,
		_w11941_,
		_w11959_,
		_w13530_
	);
	LUT3 #(
		.INIT('h80)
	) name3018 (
		\wishbone_bd_ram_mem1_reg[166][15]/P0001 ,
		_w11930_,
		_w11986_,
		_w13531_
	);
	LUT4 #(
		.INIT('h0001)
	) name3019 (
		_w13528_,
		_w13529_,
		_w13530_,
		_w13531_,
		_w13532_
	);
	LUT3 #(
		.INIT('h80)
	) name3020 (
		\wishbone_bd_ram_mem1_reg[123][15]/P0001 ,
		_w11936_,
		_w12012_,
		_w13533_
	);
	LUT3 #(
		.INIT('h80)
	) name3021 (
		\wishbone_bd_ram_mem1_reg[247][15]/P0001 ,
		_w11952_,
		_w11975_,
		_w13534_
	);
	LUT3 #(
		.INIT('h80)
	) name3022 (
		\wishbone_bd_ram_mem1_reg[133][15]/P0001 ,
		_w11933_,
		_w11955_,
		_w13535_
	);
	LUT3 #(
		.INIT('h80)
	) name3023 (
		\wishbone_bd_ram_mem1_reg[49][15]/P0001 ,
		_w11977_,
		_w11979_,
		_w13536_
	);
	LUT4 #(
		.INIT('h0001)
	) name3024 (
		_w13533_,
		_w13534_,
		_w13535_,
		_w13536_,
		_w13537_
	);
	LUT3 #(
		.INIT('h80)
	) name3025 (
		\wishbone_bd_ram_mem1_reg[240][15]/P0001 ,
		_w11941_,
		_w11952_,
		_w13538_
	);
	LUT3 #(
		.INIT('h80)
	) name3026 (
		\wishbone_bd_ram_mem1_reg[76][15]/P0001 ,
		_w11949_,
		_w11954_,
		_w13539_
	);
	LUT3 #(
		.INIT('h80)
	) name3027 (
		\wishbone_bd_ram_mem1_reg[84][15]/P0001 ,
		_w11929_,
		_w11972_,
		_w13540_
	);
	LUT3 #(
		.INIT('h80)
	) name3028 (
		\wishbone_bd_ram_mem1_reg[177][15]/P0001 ,
		_w11942_,
		_w11977_,
		_w13541_
	);
	LUT4 #(
		.INIT('h0001)
	) name3029 (
		_w13538_,
		_w13539_,
		_w13540_,
		_w13541_,
		_w13542_
	);
	LUT4 #(
		.INIT('h8000)
	) name3030 (
		_w13527_,
		_w13532_,
		_w13537_,
		_w13542_,
		_w13543_
	);
	LUT4 #(
		.INIT('h8000)
	) name3031 (
		_w13480_,
		_w13501_,
		_w13522_,
		_w13543_,
		_w13544_
	);
	LUT3 #(
		.INIT('h80)
	) name3032 (
		\wishbone_bd_ram_mem1_reg[203][15]/P0001 ,
		_w11936_,
		_w11945_,
		_w13545_
	);
	LUT3 #(
		.INIT('h80)
	) name3033 (
		\wishbone_bd_ram_mem1_reg[147][15]/P0001 ,
		_w11938_,
		_w11959_,
		_w13546_
	);
	LUT3 #(
		.INIT('h80)
	) name3034 (
		\wishbone_bd_ram_mem1_reg[1][15]/P0001 ,
		_w11932_,
		_w11977_,
		_w13547_
	);
	LUT3 #(
		.INIT('h80)
	) name3035 (
		\wishbone_bd_ram_mem1_reg[179][15]/P0001 ,
		_w11938_,
		_w11942_,
		_w13548_
	);
	LUT4 #(
		.INIT('h0001)
	) name3036 (
		_w13545_,
		_w13546_,
		_w13547_,
		_w13548_,
		_w13549_
	);
	LUT3 #(
		.INIT('h80)
	) name3037 (
		\wishbone_bd_ram_mem1_reg[80][15]/P0001 ,
		_w11941_,
		_w11972_,
		_w13550_
	);
	LUT3 #(
		.INIT('h80)
	) name3038 (
		\wishbone_bd_ram_mem1_reg[237][15]/P0001 ,
		_w11966_,
		_w11982_,
		_w13551_
	);
	LUT3 #(
		.INIT('h80)
	) name3039 (
		\wishbone_bd_ram_mem1_reg[235][15]/P0001 ,
		_w11936_,
		_w11982_,
		_w13552_
	);
	LUT3 #(
		.INIT('h80)
	) name3040 (
		\wishbone_bd_ram_mem1_reg[86][15]/P0001 ,
		_w11972_,
		_w11986_,
		_w13553_
	);
	LUT4 #(
		.INIT('h0001)
	) name3041 (
		_w13550_,
		_w13551_,
		_w13552_,
		_w13553_,
		_w13554_
	);
	LUT3 #(
		.INIT('h80)
	) name3042 (
		\wishbone_bd_ram_mem1_reg[138][15]/P0001 ,
		_w11944_,
		_w11955_,
		_w13555_
	);
	LUT3 #(
		.INIT('h80)
	) name3043 (
		\wishbone_bd_ram_mem1_reg[252][15]/P0001 ,
		_w11952_,
		_w11954_,
		_w13556_
	);
	LUT3 #(
		.INIT('h80)
	) name3044 (
		\wishbone_bd_ram_mem1_reg[22][15]/P0001 ,
		_w11935_,
		_w11986_,
		_w13557_
	);
	LUT3 #(
		.INIT('h80)
	) name3045 (
		\wishbone_bd_ram_mem1_reg[62][15]/P0001 ,
		_w11948_,
		_w11979_,
		_w13558_
	);
	LUT4 #(
		.INIT('h0001)
	) name3046 (
		_w13555_,
		_w13556_,
		_w13557_,
		_w13558_,
		_w13559_
	);
	LUT3 #(
		.INIT('h80)
	) name3047 (
		\wishbone_bd_ram_mem1_reg[45][15]/P0001 ,
		_w11957_,
		_w11966_,
		_w13560_
	);
	LUT3 #(
		.INIT('h80)
	) name3048 (
		\wishbone_bd_ram_mem1_reg[180][15]/P0001 ,
		_w11929_,
		_w11942_,
		_w13561_
	);
	LUT3 #(
		.INIT('h80)
	) name3049 (
		\wishbone_bd_ram_mem1_reg[68][15]/P0001 ,
		_w11929_,
		_w11949_,
		_w13562_
	);
	LUT3 #(
		.INIT('h80)
	) name3050 (
		\wishbone_bd_ram_mem1_reg[233][15]/P0001 ,
		_w11968_,
		_w11982_,
		_w13563_
	);
	LUT4 #(
		.INIT('h0001)
	) name3051 (
		_w13560_,
		_w13561_,
		_w13562_,
		_w13563_,
		_w13564_
	);
	LUT4 #(
		.INIT('h8000)
	) name3052 (
		_w13549_,
		_w13554_,
		_w13559_,
		_w13564_,
		_w13565_
	);
	LUT3 #(
		.INIT('h80)
	) name3053 (
		\wishbone_bd_ram_mem1_reg[212][15]/P0001 ,
		_w11929_,
		_w11984_,
		_w13566_
	);
	LUT3 #(
		.INIT('h80)
	) name3054 (
		\wishbone_bd_ram_mem1_reg[85][15]/P0001 ,
		_w11933_,
		_w11972_,
		_w13567_
	);
	LUT3 #(
		.INIT('h80)
	) name3055 (
		\wishbone_bd_ram_mem1_reg[120][15]/P0001 ,
		_w11990_,
		_w12012_,
		_w13568_
	);
	LUT3 #(
		.INIT('h80)
	) name3056 (
		\wishbone_bd_ram_mem1_reg[169][15]/P0001 ,
		_w11930_,
		_w11968_,
		_w13569_
	);
	LUT4 #(
		.INIT('h0001)
	) name3057 (
		_w13566_,
		_w13567_,
		_w13568_,
		_w13569_,
		_w13570_
	);
	LUT3 #(
		.INIT('h80)
	) name3058 (
		\wishbone_bd_ram_mem1_reg[156][15]/P0001 ,
		_w11954_,
		_w11959_,
		_w13571_
	);
	LUT3 #(
		.INIT('h80)
	) name3059 (
		\wishbone_bd_ram_mem1_reg[242][15]/P0001 ,
		_w11952_,
		_w11963_,
		_w13572_
	);
	LUT3 #(
		.INIT('h80)
	) name3060 (
		\wishbone_bd_ram_mem1_reg[199][15]/P0001 ,
		_w11945_,
		_w11975_,
		_w13573_
	);
	LUT3 #(
		.INIT('h80)
	) name3061 (
		\wishbone_bd_ram_mem1_reg[173][15]/P0001 ,
		_w11930_,
		_w11966_,
		_w13574_
	);
	LUT4 #(
		.INIT('h0001)
	) name3062 (
		_w13571_,
		_w13572_,
		_w13573_,
		_w13574_,
		_w13575_
	);
	LUT3 #(
		.INIT('h80)
	) name3063 (
		\wishbone_bd_ram_mem1_reg[197][15]/P0001 ,
		_w11933_,
		_w11945_,
		_w13576_
	);
	LUT3 #(
		.INIT('h80)
	) name3064 (
		\wishbone_bd_ram_mem1_reg[155][15]/P0001 ,
		_w11936_,
		_w11959_,
		_w13577_
	);
	LUT3 #(
		.INIT('h80)
	) name3065 (
		\wishbone_bd_ram_mem1_reg[164][15]/P0001 ,
		_w11929_,
		_w11930_,
		_w13578_
	);
	LUT3 #(
		.INIT('h80)
	) name3066 (
		\wishbone_bd_ram_mem1_reg[226][15]/P0001 ,
		_w11963_,
		_w11982_,
		_w13579_
	);
	LUT4 #(
		.INIT('h0001)
	) name3067 (
		_w13576_,
		_w13577_,
		_w13578_,
		_w13579_,
		_w13580_
	);
	LUT3 #(
		.INIT('h80)
	) name3068 (
		\wishbone_bd_ram_mem1_reg[191][15]/P0001 ,
		_w11942_,
		_w11973_,
		_w13581_
	);
	LUT3 #(
		.INIT('h80)
	) name3069 (
		\wishbone_bd_ram_mem1_reg[217][15]/P0001 ,
		_w11968_,
		_w11984_,
		_w13582_
	);
	LUT3 #(
		.INIT('h80)
	) name3070 (
		\wishbone_bd_ram_mem1_reg[108][15]/P0001 ,
		_w11954_,
		_w11965_,
		_w13583_
	);
	LUT3 #(
		.INIT('h80)
	) name3071 (
		\wishbone_bd_ram_mem1_reg[139][15]/P0001 ,
		_w11936_,
		_w11955_,
		_w13584_
	);
	LUT4 #(
		.INIT('h0001)
	) name3072 (
		_w13581_,
		_w13582_,
		_w13583_,
		_w13584_,
		_w13585_
	);
	LUT4 #(
		.INIT('h8000)
	) name3073 (
		_w13570_,
		_w13575_,
		_w13580_,
		_w13585_,
		_w13586_
	);
	LUT3 #(
		.INIT('h80)
	) name3074 (
		\wishbone_bd_ram_mem1_reg[73][15]/P0001 ,
		_w11949_,
		_w11968_,
		_w13587_
	);
	LUT3 #(
		.INIT('h80)
	) name3075 (
		\wishbone_bd_ram_mem1_reg[201][15]/P0001 ,
		_w11945_,
		_w11968_,
		_w13588_
	);
	LUT3 #(
		.INIT('h80)
	) name3076 (
		\wishbone_bd_ram_mem1_reg[37][15]/P0001 ,
		_w11933_,
		_w11957_,
		_w13589_
	);
	LUT3 #(
		.INIT('h80)
	) name3077 (
		\wishbone_bd_ram_mem1_reg[104][15]/P0001 ,
		_w11965_,
		_w11990_,
		_w13590_
	);
	LUT4 #(
		.INIT('h0001)
	) name3078 (
		_w13587_,
		_w13588_,
		_w13589_,
		_w13590_,
		_w13591_
	);
	LUT3 #(
		.INIT('h80)
	) name3079 (
		\wishbone_bd_ram_mem1_reg[52][15]/P0001 ,
		_w11929_,
		_w11979_,
		_w13592_
	);
	LUT3 #(
		.INIT('h80)
	) name3080 (
		\wishbone_bd_ram_mem1_reg[112][15]/P0001 ,
		_w11941_,
		_w12012_,
		_w13593_
	);
	LUT3 #(
		.INIT('h80)
	) name3081 (
		\wishbone_bd_ram_mem1_reg[255][15]/P0001 ,
		_w11952_,
		_w11973_,
		_w13594_
	);
	LUT3 #(
		.INIT('h80)
	) name3082 (
		\wishbone_bd_ram_mem1_reg[175][15]/P0001 ,
		_w11930_,
		_w11973_,
		_w13595_
	);
	LUT4 #(
		.INIT('h0001)
	) name3083 (
		_w13592_,
		_w13593_,
		_w13594_,
		_w13595_,
		_w13596_
	);
	LUT3 #(
		.INIT('h80)
	) name3084 (
		\wishbone_bd_ram_mem1_reg[238][15]/P0001 ,
		_w11948_,
		_w11982_,
		_w13597_
	);
	LUT3 #(
		.INIT('h80)
	) name3085 (
		\wishbone_bd_ram_mem1_reg[58][15]/P0001 ,
		_w11944_,
		_w11979_,
		_w13598_
	);
	LUT3 #(
		.INIT('h80)
	) name3086 (
		\wishbone_bd_ram_mem1_reg[195][15]/P0001 ,
		_w11938_,
		_w11945_,
		_w13599_
	);
	LUT3 #(
		.INIT('h80)
	) name3087 (
		\wishbone_bd_ram_mem1_reg[60][15]/P0001 ,
		_w11954_,
		_w11979_,
		_w13600_
	);
	LUT4 #(
		.INIT('h0001)
	) name3088 (
		_w13597_,
		_w13598_,
		_w13599_,
		_w13600_,
		_w13601_
	);
	LUT3 #(
		.INIT('h80)
	) name3089 (
		\wishbone_bd_ram_mem1_reg[27][15]/P0001 ,
		_w11935_,
		_w11936_,
		_w13602_
	);
	LUT3 #(
		.INIT('h80)
	) name3090 (
		\wishbone_bd_ram_mem1_reg[7][15]/P0001 ,
		_w11932_,
		_w11975_,
		_w13603_
	);
	LUT3 #(
		.INIT('h80)
	) name3091 (
		\wishbone_bd_ram_mem1_reg[150][15]/P0001 ,
		_w11959_,
		_w11986_,
		_w13604_
	);
	LUT3 #(
		.INIT('h80)
	) name3092 (
		\wishbone_bd_ram_mem1_reg[215][15]/P0001 ,
		_w11975_,
		_w11984_,
		_w13605_
	);
	LUT4 #(
		.INIT('h0001)
	) name3093 (
		_w13602_,
		_w13603_,
		_w13604_,
		_w13605_,
		_w13606_
	);
	LUT4 #(
		.INIT('h8000)
	) name3094 (
		_w13591_,
		_w13596_,
		_w13601_,
		_w13606_,
		_w13607_
	);
	LUT3 #(
		.INIT('h80)
	) name3095 (
		\wishbone_bd_ram_mem1_reg[88][15]/P0001 ,
		_w11972_,
		_w11990_,
		_w13608_
	);
	LUT3 #(
		.INIT('h80)
	) name3096 (
		\wishbone_bd_ram_mem1_reg[172][15]/P0001 ,
		_w11930_,
		_w11954_,
		_w13609_
	);
	LUT3 #(
		.INIT('h80)
	) name3097 (
		\wishbone_bd_ram_mem1_reg[129][15]/P0001 ,
		_w11955_,
		_w11977_,
		_w13610_
	);
	LUT3 #(
		.INIT('h80)
	) name3098 (
		\wishbone_bd_ram_mem1_reg[227][15]/P0001 ,
		_w11938_,
		_w11982_,
		_w13611_
	);
	LUT4 #(
		.INIT('h0001)
	) name3099 (
		_w13608_,
		_w13609_,
		_w13610_,
		_w13611_,
		_w13612_
	);
	LUT3 #(
		.INIT('h80)
	) name3100 (
		\wishbone_bd_ram_mem1_reg[188][15]/P0001 ,
		_w11942_,
		_w11954_,
		_w13613_
	);
	LUT3 #(
		.INIT('h80)
	) name3101 (
		\wishbone_bd_ram_mem1_reg[198][15]/P0001 ,
		_w11945_,
		_w11986_,
		_w13614_
	);
	LUT3 #(
		.INIT('h80)
	) name3102 (
		\wishbone_bd_ram_mem1_reg[249][15]/P0001 ,
		_w11952_,
		_w11968_,
		_w13615_
	);
	LUT3 #(
		.INIT('h80)
	) name3103 (
		\wishbone_bd_ram_mem1_reg[196][15]/P0001 ,
		_w11929_,
		_w11945_,
		_w13616_
	);
	LUT4 #(
		.INIT('h0001)
	) name3104 (
		_w13613_,
		_w13614_,
		_w13615_,
		_w13616_,
		_w13617_
	);
	LUT3 #(
		.INIT('h80)
	) name3105 (
		\wishbone_bd_ram_mem1_reg[67][15]/P0001 ,
		_w11938_,
		_w11949_,
		_w13618_
	);
	LUT3 #(
		.INIT('h80)
	) name3106 (
		\wishbone_bd_ram_mem1_reg[41][15]/P0001 ,
		_w11957_,
		_w11968_,
		_w13619_
	);
	LUT3 #(
		.INIT('h80)
	) name3107 (
		\wishbone_bd_ram_mem1_reg[122][15]/P0001 ,
		_w11944_,
		_w12012_,
		_w13620_
	);
	LUT3 #(
		.INIT('h80)
	) name3108 (
		\wishbone_bd_ram_mem1_reg[25][15]/P0001 ,
		_w11935_,
		_w11968_,
		_w13621_
	);
	LUT4 #(
		.INIT('h0001)
	) name3109 (
		_w13618_,
		_w13619_,
		_w13620_,
		_w13621_,
		_w13622_
	);
	LUT3 #(
		.INIT('h80)
	) name3110 (
		\wishbone_bd_ram_mem1_reg[18][15]/P0001 ,
		_w11935_,
		_w11963_,
		_w13623_
	);
	LUT3 #(
		.INIT('h80)
	) name3111 (
		\wishbone_bd_ram_mem1_reg[181][15]/P0001 ,
		_w11933_,
		_w11942_,
		_w13624_
	);
	LUT3 #(
		.INIT('h80)
	) name3112 (
		\wishbone_bd_ram_mem1_reg[20][15]/P0001 ,
		_w11929_,
		_w11935_,
		_w13625_
	);
	LUT3 #(
		.INIT('h80)
	) name3113 (
		\wishbone_bd_ram_mem1_reg[189][15]/P0001 ,
		_w11942_,
		_w11966_,
		_w13626_
	);
	LUT4 #(
		.INIT('h0001)
	) name3114 (
		_w13623_,
		_w13624_,
		_w13625_,
		_w13626_,
		_w13627_
	);
	LUT4 #(
		.INIT('h8000)
	) name3115 (
		_w13612_,
		_w13617_,
		_w13622_,
		_w13627_,
		_w13628_
	);
	LUT4 #(
		.INIT('h8000)
	) name3116 (
		_w13565_,
		_w13586_,
		_w13607_,
		_w13628_,
		_w13629_
	);
	LUT3 #(
		.INIT('h80)
	) name3117 (
		\wishbone_bd_ram_mem1_reg[121][15]/P0001 ,
		_w11968_,
		_w12012_,
		_w13630_
	);
	LUT3 #(
		.INIT('h80)
	) name3118 (
		\wishbone_bd_ram_mem1_reg[65][15]/P0001 ,
		_w11949_,
		_w11977_,
		_w13631_
	);
	LUT3 #(
		.INIT('h80)
	) name3119 (
		\wishbone_bd_ram_mem1_reg[229][15]/P0001 ,
		_w11933_,
		_w11982_,
		_w13632_
	);
	LUT3 #(
		.INIT('h80)
	) name3120 (
		\wishbone_bd_ram_mem1_reg[100][15]/P0001 ,
		_w11929_,
		_w11965_,
		_w13633_
	);
	LUT4 #(
		.INIT('h0001)
	) name3121 (
		_w13630_,
		_w13631_,
		_w13632_,
		_w13633_,
		_w13634_
	);
	LUT3 #(
		.INIT('h80)
	) name3122 (
		\wishbone_bd_ram_mem1_reg[223][15]/P0001 ,
		_w11973_,
		_w11984_,
		_w13635_
	);
	LUT3 #(
		.INIT('h80)
	) name3123 (
		\wishbone_bd_ram_mem1_reg[89][15]/P0001 ,
		_w11968_,
		_w11972_,
		_w13636_
	);
	LUT3 #(
		.INIT('h80)
	) name3124 (
		\wishbone_bd_ram_mem1_reg[6][15]/P0001 ,
		_w11932_,
		_w11986_,
		_w13637_
	);
	LUT3 #(
		.INIT('h80)
	) name3125 (
		\wishbone_bd_ram_mem1_reg[70][15]/P0001 ,
		_w11949_,
		_w11986_,
		_w13638_
	);
	LUT4 #(
		.INIT('h0001)
	) name3126 (
		_w13635_,
		_w13636_,
		_w13637_,
		_w13638_,
		_w13639_
	);
	LUT3 #(
		.INIT('h80)
	) name3127 (
		\wishbone_bd_ram_mem1_reg[38][15]/P0001 ,
		_w11957_,
		_w11986_,
		_w13640_
	);
	LUT3 #(
		.INIT('h80)
	) name3128 (
		\wishbone_bd_ram_mem1_reg[34][15]/P0001 ,
		_w11957_,
		_w11963_,
		_w13641_
	);
	LUT3 #(
		.INIT('h80)
	) name3129 (
		\wishbone_bd_ram_mem1_reg[3][15]/P0001 ,
		_w11932_,
		_w11938_,
		_w13642_
	);
	LUT3 #(
		.INIT('h80)
	) name3130 (
		\wishbone_bd_ram_mem1_reg[63][15]/P0001 ,
		_w11973_,
		_w11979_,
		_w13643_
	);
	LUT4 #(
		.INIT('h0001)
	) name3131 (
		_w13640_,
		_w13641_,
		_w13642_,
		_w13643_,
		_w13644_
	);
	LUT3 #(
		.INIT('h80)
	) name3132 (
		\wishbone_bd_ram_mem1_reg[183][15]/P0001 ,
		_w11942_,
		_w11975_,
		_w13645_
	);
	LUT3 #(
		.INIT('h80)
	) name3133 (
		\wishbone_bd_ram_mem1_reg[96][15]/P0001 ,
		_w11941_,
		_w11965_,
		_w13646_
	);
	LUT3 #(
		.INIT('h80)
	) name3134 (
		\wishbone_bd_ram_mem1_reg[228][15]/P0001 ,
		_w11929_,
		_w11982_,
		_w13647_
	);
	LUT3 #(
		.INIT('h80)
	) name3135 (
		\wishbone_bd_ram_mem1_reg[59][15]/P0001 ,
		_w11936_,
		_w11979_,
		_w13648_
	);
	LUT4 #(
		.INIT('h0001)
	) name3136 (
		_w13645_,
		_w13646_,
		_w13647_,
		_w13648_,
		_w13649_
	);
	LUT4 #(
		.INIT('h8000)
	) name3137 (
		_w13634_,
		_w13639_,
		_w13644_,
		_w13649_,
		_w13650_
	);
	LUT3 #(
		.INIT('h80)
	) name3138 (
		\wishbone_bd_ram_mem1_reg[159][15]/P0001 ,
		_w11959_,
		_w11973_,
		_w13651_
	);
	LUT3 #(
		.INIT('h80)
	) name3139 (
		\wishbone_bd_ram_mem1_reg[56][15]/P0001 ,
		_w11979_,
		_w11990_,
		_w13652_
	);
	LUT3 #(
		.INIT('h80)
	) name3140 (
		\wishbone_bd_ram_mem1_reg[12][15]/P0001 ,
		_w11932_,
		_w11954_,
		_w13653_
	);
	LUT3 #(
		.INIT('h80)
	) name3141 (
		\wishbone_bd_ram_mem1_reg[161][15]/P0001 ,
		_w11930_,
		_w11977_,
		_w13654_
	);
	LUT4 #(
		.INIT('h0001)
	) name3142 (
		_w13651_,
		_w13652_,
		_w13653_,
		_w13654_,
		_w13655_
	);
	LUT3 #(
		.INIT('h80)
	) name3143 (
		\wishbone_bd_ram_mem1_reg[23][15]/P0001 ,
		_w11935_,
		_w11975_,
		_w13656_
	);
	LUT3 #(
		.INIT('h80)
	) name3144 (
		\wishbone_bd_ram_mem1_reg[208][15]/P0001 ,
		_w11941_,
		_w11984_,
		_w13657_
	);
	LUT3 #(
		.INIT('h80)
	) name3145 (
		\wishbone_bd_ram_mem1_reg[54][15]/P0001 ,
		_w11979_,
		_w11986_,
		_w13658_
	);
	LUT3 #(
		.INIT('h80)
	) name3146 (
		\wishbone_bd_ram_mem1_reg[248][15]/P0001 ,
		_w11952_,
		_w11990_,
		_w13659_
	);
	LUT4 #(
		.INIT('h0001)
	) name3147 (
		_w13656_,
		_w13657_,
		_w13658_,
		_w13659_,
		_w13660_
	);
	LUT3 #(
		.INIT('h80)
	) name3148 (
		\wishbone_bd_ram_mem1_reg[135][15]/P0001 ,
		_w11955_,
		_w11975_,
		_w13661_
	);
	LUT3 #(
		.INIT('h80)
	) name3149 (
		\wishbone_bd_ram_mem1_reg[2][15]/P0001 ,
		_w11932_,
		_w11963_,
		_w13662_
	);
	LUT3 #(
		.INIT('h80)
	) name3150 (
		\wishbone_bd_ram_mem1_reg[184][15]/P0001 ,
		_w11942_,
		_w11990_,
		_w13663_
	);
	LUT3 #(
		.INIT('h80)
	) name3151 (
		\wishbone_bd_ram_mem1_reg[154][15]/P0001 ,
		_w11944_,
		_w11959_,
		_w13664_
	);
	LUT4 #(
		.INIT('h0001)
	) name3152 (
		_w13661_,
		_w13662_,
		_w13663_,
		_w13664_,
		_w13665_
	);
	LUT3 #(
		.INIT('h80)
	) name3153 (
		\wishbone_bd_ram_mem1_reg[92][15]/P0001 ,
		_w11954_,
		_w11972_,
		_w13666_
	);
	LUT3 #(
		.INIT('h80)
	) name3154 (
		\wishbone_bd_ram_mem1_reg[186][15]/P0001 ,
		_w11942_,
		_w11944_,
		_w13667_
	);
	LUT3 #(
		.INIT('h80)
	) name3155 (
		\wishbone_bd_ram_mem1_reg[19][15]/P0001 ,
		_w11935_,
		_w11938_,
		_w13668_
	);
	LUT3 #(
		.INIT('h80)
	) name3156 (
		\wishbone_bd_ram_mem1_reg[232][15]/P0001 ,
		_w11982_,
		_w11990_,
		_w13669_
	);
	LUT4 #(
		.INIT('h0001)
	) name3157 (
		_w13666_,
		_w13667_,
		_w13668_,
		_w13669_,
		_w13670_
	);
	LUT4 #(
		.INIT('h8000)
	) name3158 (
		_w13655_,
		_w13660_,
		_w13665_,
		_w13670_,
		_w13671_
	);
	LUT3 #(
		.INIT('h80)
	) name3159 (
		\wishbone_bd_ram_mem1_reg[51][15]/P0001 ,
		_w11938_,
		_w11979_,
		_w13672_
	);
	LUT3 #(
		.INIT('h80)
	) name3160 (
		\wishbone_bd_ram_mem1_reg[250][15]/P0001 ,
		_w11944_,
		_w11952_,
		_w13673_
	);
	LUT3 #(
		.INIT('h80)
	) name3161 (
		\wishbone_bd_ram_mem1_reg[185][15]/P0001 ,
		_w11942_,
		_w11968_,
		_w13674_
	);
	LUT3 #(
		.INIT('h80)
	) name3162 (
		\wishbone_bd_ram_mem1_reg[148][15]/P0001 ,
		_w11929_,
		_w11959_,
		_w13675_
	);
	LUT4 #(
		.INIT('h0001)
	) name3163 (
		_w13672_,
		_w13673_,
		_w13674_,
		_w13675_,
		_w13676_
	);
	LUT3 #(
		.INIT('h80)
	) name3164 (
		\wishbone_bd_ram_mem1_reg[10][15]/P0001 ,
		_w11932_,
		_w11944_,
		_w13677_
	);
	LUT3 #(
		.INIT('h80)
	) name3165 (
		\wishbone_bd_ram_mem1_reg[102][15]/P0001 ,
		_w11965_,
		_w11986_,
		_w13678_
	);
	LUT3 #(
		.INIT('h80)
	) name3166 (
		\wishbone_bd_ram_mem1_reg[136][15]/P0001 ,
		_w11955_,
		_w11990_,
		_w13679_
	);
	LUT3 #(
		.INIT('h80)
	) name3167 (
		\wishbone_bd_ram_mem1_reg[190][15]/P0001 ,
		_w11942_,
		_w11948_,
		_w13680_
	);
	LUT4 #(
		.INIT('h0001)
	) name3168 (
		_w13677_,
		_w13678_,
		_w13679_,
		_w13680_,
		_w13681_
	);
	LUT3 #(
		.INIT('h80)
	) name3169 (
		\wishbone_bd_ram_mem1_reg[114][15]/P0001 ,
		_w11963_,
		_w12012_,
		_w13682_
	);
	LUT3 #(
		.INIT('h80)
	) name3170 (
		\wishbone_bd_ram_mem1_reg[94][15]/P0001 ,
		_w11948_,
		_w11972_,
		_w13683_
	);
	LUT3 #(
		.INIT('h80)
	) name3171 (
		\wishbone_bd_ram_mem1_reg[236][15]/P0001 ,
		_w11954_,
		_w11982_,
		_w13684_
	);
	LUT3 #(
		.INIT('h80)
	) name3172 (
		\wishbone_bd_ram_mem1_reg[113][15]/P0001 ,
		_w11977_,
		_w12012_,
		_w13685_
	);
	LUT4 #(
		.INIT('h0001)
	) name3173 (
		_w13682_,
		_w13683_,
		_w13684_,
		_w13685_,
		_w13686_
	);
	LUT3 #(
		.INIT('h80)
	) name3174 (
		\wishbone_bd_ram_mem1_reg[57][15]/P0001 ,
		_w11968_,
		_w11979_,
		_w13687_
	);
	LUT3 #(
		.INIT('h80)
	) name3175 (
		\wishbone_bd_ram_mem1_reg[254][15]/P0001 ,
		_w11948_,
		_w11952_,
		_w13688_
	);
	LUT3 #(
		.INIT('h80)
	) name3176 (
		\wishbone_bd_ram_mem1_reg[245][15]/P0001 ,
		_w11933_,
		_w11952_,
		_w13689_
	);
	LUT3 #(
		.INIT('h80)
	) name3177 (
		\wishbone_bd_ram_mem1_reg[253][15]/P0001 ,
		_w11952_,
		_w11966_,
		_w13690_
	);
	LUT4 #(
		.INIT('h0001)
	) name3178 (
		_w13687_,
		_w13688_,
		_w13689_,
		_w13690_,
		_w13691_
	);
	LUT4 #(
		.INIT('h8000)
	) name3179 (
		_w13676_,
		_w13681_,
		_w13686_,
		_w13691_,
		_w13692_
	);
	LUT3 #(
		.INIT('h80)
	) name3180 (
		\wishbone_bd_ram_mem1_reg[79][15]/P0001 ,
		_w11949_,
		_w11973_,
		_w13693_
	);
	LUT3 #(
		.INIT('h80)
	) name3181 (
		\wishbone_bd_ram_mem1_reg[5][15]/P0001 ,
		_w11932_,
		_w11933_,
		_w13694_
	);
	LUT3 #(
		.INIT('h80)
	) name3182 (
		\wishbone_bd_ram_mem1_reg[53][15]/P0001 ,
		_w11933_,
		_w11979_,
		_w13695_
	);
	LUT3 #(
		.INIT('h80)
	) name3183 (
		\wishbone_bd_ram_mem1_reg[225][15]/P0001 ,
		_w11977_,
		_w11982_,
		_w13696_
	);
	LUT4 #(
		.INIT('h0001)
	) name3184 (
		_w13693_,
		_w13694_,
		_w13695_,
		_w13696_,
		_w13697_
	);
	LUT3 #(
		.INIT('h80)
	) name3185 (
		\wishbone_bd_ram_mem1_reg[231][15]/P0001 ,
		_w11975_,
		_w11982_,
		_w13698_
	);
	LUT3 #(
		.INIT('h80)
	) name3186 (
		\wishbone_bd_ram_mem1_reg[209][15]/P0001 ,
		_w11977_,
		_w11984_,
		_w13699_
	);
	LUT3 #(
		.INIT('h80)
	) name3187 (
		\wishbone_bd_ram_mem1_reg[216][15]/P0001 ,
		_w11984_,
		_w11990_,
		_w13700_
	);
	LUT3 #(
		.INIT('h80)
	) name3188 (
		\wishbone_bd_ram_mem1_reg[8][15]/P0001 ,
		_w11932_,
		_w11990_,
		_w13701_
	);
	LUT4 #(
		.INIT('h0001)
	) name3189 (
		_w13698_,
		_w13699_,
		_w13700_,
		_w13701_,
		_w13702_
	);
	LUT3 #(
		.INIT('h80)
	) name3190 (
		\wishbone_bd_ram_mem1_reg[55][15]/P0001 ,
		_w11975_,
		_w11979_,
		_w13703_
	);
	LUT3 #(
		.INIT('h80)
	) name3191 (
		\wishbone_bd_ram_mem1_reg[157][15]/P0001 ,
		_w11959_,
		_w11966_,
		_w13704_
	);
	LUT3 #(
		.INIT('h80)
	) name3192 (
		\wishbone_bd_ram_mem1_reg[93][15]/P0001 ,
		_w11966_,
		_w11972_,
		_w13705_
	);
	LUT3 #(
		.INIT('h80)
	) name3193 (
		\wishbone_bd_ram_mem1_reg[176][15]/P0001 ,
		_w11941_,
		_w11942_,
		_w13706_
	);
	LUT4 #(
		.INIT('h0001)
	) name3194 (
		_w13703_,
		_w13704_,
		_w13705_,
		_w13706_,
		_w13707_
	);
	LUT3 #(
		.INIT('h80)
	) name3195 (
		\wishbone_bd_ram_mem1_reg[110][15]/P0001 ,
		_w11948_,
		_w11965_,
		_w13708_
	);
	LUT3 #(
		.INIT('h80)
	) name3196 (
		\wishbone_bd_ram_mem1_reg[230][15]/P0001 ,
		_w11982_,
		_w11986_,
		_w13709_
	);
	LUT3 #(
		.INIT('h80)
	) name3197 (
		\wishbone_bd_ram_mem1_reg[69][15]/P0001 ,
		_w11933_,
		_w11949_,
		_w13710_
	);
	LUT3 #(
		.INIT('h80)
	) name3198 (
		\wishbone_bd_ram_mem1_reg[146][15]/P0001 ,
		_w11959_,
		_w11963_,
		_w13711_
	);
	LUT4 #(
		.INIT('h0001)
	) name3199 (
		_w13708_,
		_w13709_,
		_w13710_,
		_w13711_,
		_w13712_
	);
	LUT4 #(
		.INIT('h8000)
	) name3200 (
		_w13697_,
		_w13702_,
		_w13707_,
		_w13712_,
		_w13713_
	);
	LUT4 #(
		.INIT('h8000)
	) name3201 (
		_w13650_,
		_w13671_,
		_w13692_,
		_w13713_,
		_w13714_
	);
	LUT3 #(
		.INIT('h80)
	) name3202 (
		\wishbone_bd_ram_mem1_reg[130][15]/P0001 ,
		_w11955_,
		_w11963_,
		_w13715_
	);
	LUT3 #(
		.INIT('h80)
	) name3203 (
		\wishbone_bd_ram_mem1_reg[48][15]/P0001 ,
		_w11941_,
		_w11979_,
		_w13716_
	);
	LUT3 #(
		.INIT('h80)
	) name3204 (
		\wishbone_bd_ram_mem1_reg[207][15]/P0001 ,
		_w11945_,
		_w11973_,
		_w13717_
	);
	LUT3 #(
		.INIT('h80)
	) name3205 (
		\wishbone_bd_ram_mem1_reg[71][15]/P0001 ,
		_w11949_,
		_w11975_,
		_w13718_
	);
	LUT4 #(
		.INIT('h0001)
	) name3206 (
		_w13715_,
		_w13716_,
		_w13717_,
		_w13718_,
		_w13719_
	);
	LUT3 #(
		.INIT('h80)
	) name3207 (
		\wishbone_bd_ram_mem1_reg[125][15]/P0001 ,
		_w11966_,
		_w12012_,
		_w13720_
	);
	LUT3 #(
		.INIT('h80)
	) name3208 (
		\wishbone_bd_ram_mem1_reg[28][15]/P0001 ,
		_w11935_,
		_w11954_,
		_w13721_
	);
	LUT3 #(
		.INIT('h80)
	) name3209 (
		\wishbone_bd_ram_mem1_reg[127][15]/P0001 ,
		_w11973_,
		_w12012_,
		_w13722_
	);
	LUT3 #(
		.INIT('h80)
	) name3210 (
		\wishbone_bd_ram_mem1_reg[74][15]/P0001 ,
		_w11944_,
		_w11949_,
		_w13723_
	);
	LUT4 #(
		.INIT('h0001)
	) name3211 (
		_w13720_,
		_w13721_,
		_w13722_,
		_w13723_,
		_w13724_
	);
	LUT3 #(
		.INIT('h80)
	) name3212 (
		\wishbone_bd_ram_mem1_reg[31][15]/P0001 ,
		_w11935_,
		_w11973_,
		_w13725_
	);
	LUT3 #(
		.INIT('h80)
	) name3213 (
		\wishbone_bd_ram_mem1_reg[82][15]/P0001 ,
		_w11963_,
		_w11972_,
		_w13726_
	);
	LUT3 #(
		.INIT('h80)
	) name3214 (
		\wishbone_bd_ram_mem1_reg[137][15]/P0001 ,
		_w11955_,
		_w11968_,
		_w13727_
	);
	LUT3 #(
		.INIT('h80)
	) name3215 (
		\wishbone_bd_ram_mem1_reg[200][15]/P0001 ,
		_w11945_,
		_w11990_,
		_w13728_
	);
	LUT4 #(
		.INIT('h0001)
	) name3216 (
		_w13725_,
		_w13726_,
		_w13727_,
		_w13728_,
		_w13729_
	);
	LUT3 #(
		.INIT('h80)
	) name3217 (
		\wishbone_bd_ram_mem1_reg[11][15]/P0001 ,
		_w11932_,
		_w11936_,
		_w13730_
	);
	LUT3 #(
		.INIT('h80)
	) name3218 (
		\wishbone_bd_ram_mem1_reg[106][15]/P0001 ,
		_w11944_,
		_w11965_,
		_w13731_
	);
	LUT3 #(
		.INIT('h80)
	) name3219 (
		\wishbone_bd_ram_mem1_reg[251][15]/P0001 ,
		_w11936_,
		_w11952_,
		_w13732_
	);
	LUT3 #(
		.INIT('h80)
	) name3220 (
		\wishbone_bd_ram_mem1_reg[204][15]/P0001 ,
		_w11945_,
		_w11954_,
		_w13733_
	);
	LUT4 #(
		.INIT('h0001)
	) name3221 (
		_w13730_,
		_w13731_,
		_w13732_,
		_w13733_,
		_w13734_
	);
	LUT4 #(
		.INIT('h8000)
	) name3222 (
		_w13719_,
		_w13724_,
		_w13729_,
		_w13734_,
		_w13735_
	);
	LUT3 #(
		.INIT('h80)
	) name3223 (
		\wishbone_bd_ram_mem1_reg[171][15]/P0001 ,
		_w11930_,
		_w11936_,
		_w13736_
	);
	LUT3 #(
		.INIT('h80)
	) name3224 (
		\wishbone_bd_ram_mem1_reg[91][15]/P0001 ,
		_w11936_,
		_w11972_,
		_w13737_
	);
	LUT3 #(
		.INIT('h80)
	) name3225 (
		\wishbone_bd_ram_mem1_reg[33][15]/P0001 ,
		_w11957_,
		_w11977_,
		_w13738_
	);
	LUT3 #(
		.INIT('h80)
	) name3226 (
		\wishbone_bd_ram_mem1_reg[174][15]/P0001 ,
		_w11930_,
		_w11948_,
		_w13739_
	);
	LUT4 #(
		.INIT('h0001)
	) name3227 (
		_w13736_,
		_w13737_,
		_w13738_,
		_w13739_,
		_w13740_
	);
	LUT3 #(
		.INIT('h80)
	) name3228 (
		\wishbone_bd_ram_mem1_reg[78][15]/P0001 ,
		_w11948_,
		_w11949_,
		_w13741_
	);
	LUT3 #(
		.INIT('h80)
	) name3229 (
		\wishbone_bd_ram_mem1_reg[178][15]/P0001 ,
		_w11942_,
		_w11963_,
		_w13742_
	);
	LUT3 #(
		.INIT('h80)
	) name3230 (
		\wishbone_bd_ram_mem1_reg[219][15]/P0001 ,
		_w11936_,
		_w11984_,
		_w13743_
	);
	LUT3 #(
		.INIT('h80)
	) name3231 (
		\wishbone_bd_ram_mem1_reg[187][15]/P0001 ,
		_w11936_,
		_w11942_,
		_w13744_
	);
	LUT4 #(
		.INIT('h0001)
	) name3232 (
		_w13741_,
		_w13742_,
		_w13743_,
		_w13744_,
		_w13745_
	);
	LUT3 #(
		.INIT('h80)
	) name3233 (
		\wishbone_bd_ram_mem1_reg[170][15]/P0001 ,
		_w11930_,
		_w11944_,
		_w13746_
	);
	LUT3 #(
		.INIT('h80)
	) name3234 (
		\wishbone_bd_ram_mem1_reg[241][15]/P0001 ,
		_w11952_,
		_w11977_,
		_w13747_
	);
	LUT3 #(
		.INIT('h80)
	) name3235 (
		\wishbone_bd_ram_mem1_reg[115][15]/P0001 ,
		_w11938_,
		_w12012_,
		_w13748_
	);
	LUT3 #(
		.INIT('h80)
	) name3236 (
		\wishbone_bd_ram_mem1_reg[24][15]/P0001 ,
		_w11935_,
		_w11990_,
		_w13749_
	);
	LUT4 #(
		.INIT('h0001)
	) name3237 (
		_w13746_,
		_w13747_,
		_w13748_,
		_w13749_,
		_w13750_
	);
	LUT3 #(
		.INIT('h80)
	) name3238 (
		\wishbone_bd_ram_mem1_reg[61][15]/P0001 ,
		_w11966_,
		_w11979_,
		_w13751_
	);
	LUT3 #(
		.INIT('h80)
	) name3239 (
		\wishbone_bd_ram_mem1_reg[64][15]/P0001 ,
		_w11941_,
		_w11949_,
		_w13752_
	);
	LUT3 #(
		.INIT('h80)
	) name3240 (
		\wishbone_bd_ram_mem1_reg[111][15]/P0001 ,
		_w11965_,
		_w11973_,
		_w13753_
	);
	LUT3 #(
		.INIT('h80)
	) name3241 (
		\wishbone_bd_ram_mem1_reg[222][15]/P0001 ,
		_w11948_,
		_w11984_,
		_w13754_
	);
	LUT4 #(
		.INIT('h0001)
	) name3242 (
		_w13751_,
		_w13752_,
		_w13753_,
		_w13754_,
		_w13755_
	);
	LUT4 #(
		.INIT('h8000)
	) name3243 (
		_w13740_,
		_w13745_,
		_w13750_,
		_w13755_,
		_w13756_
	);
	LUT3 #(
		.INIT('h80)
	) name3244 (
		\wishbone_bd_ram_mem1_reg[220][15]/P0001 ,
		_w11954_,
		_w11984_,
		_w13757_
	);
	LUT3 #(
		.INIT('h80)
	) name3245 (
		\wishbone_bd_ram_mem1_reg[95][15]/P0001 ,
		_w11972_,
		_w11973_,
		_w13758_
	);
	LUT3 #(
		.INIT('h80)
	) name3246 (
		\wishbone_bd_ram_mem1_reg[16][15]/P0001 ,
		_w11935_,
		_w11941_,
		_w13759_
	);
	LUT3 #(
		.INIT('h80)
	) name3247 (
		\wishbone_bd_ram_mem1_reg[81][15]/P0001 ,
		_w11972_,
		_w11977_,
		_w13760_
	);
	LUT4 #(
		.INIT('h0001)
	) name3248 (
		_w13757_,
		_w13758_,
		_w13759_,
		_w13760_,
		_w13761_
	);
	LUT3 #(
		.INIT('h80)
	) name3249 (
		\wishbone_bd_ram_mem1_reg[128][15]/P0001 ,
		_w11941_,
		_w11955_,
		_w13762_
	);
	LUT3 #(
		.INIT('h80)
	) name3250 (
		\wishbone_bd_ram_mem1_reg[124][15]/P0001 ,
		_w11954_,
		_w12012_,
		_w13763_
	);
	LUT3 #(
		.INIT('h80)
	) name3251 (
		\wishbone_bd_ram_mem1_reg[239][15]/P0001 ,
		_w11973_,
		_w11982_,
		_w13764_
	);
	LUT3 #(
		.INIT('h80)
	) name3252 (
		\wishbone_bd_ram_mem1_reg[17][15]/P0001 ,
		_w11935_,
		_w11977_,
		_w13765_
	);
	LUT4 #(
		.INIT('h0001)
	) name3253 (
		_w13762_,
		_w13763_,
		_w13764_,
		_w13765_,
		_w13766_
	);
	LUT3 #(
		.INIT('h80)
	) name3254 (
		\wishbone_bd_ram_mem1_reg[244][15]/P0001 ,
		_w11929_,
		_w11952_,
		_w13767_
	);
	LUT3 #(
		.INIT('h80)
	) name3255 (
		\wishbone_bd_ram_mem1_reg[87][15]/P0001 ,
		_w11972_,
		_w11975_,
		_w13768_
	);
	LUT3 #(
		.INIT('h80)
	) name3256 (
		\wishbone_bd_ram_mem1_reg[140][15]/P0001 ,
		_w11954_,
		_w11955_,
		_w13769_
	);
	LUT3 #(
		.INIT('h80)
	) name3257 (
		\wishbone_bd_ram_mem1_reg[158][15]/P0001 ,
		_w11948_,
		_w11959_,
		_w13770_
	);
	LUT4 #(
		.INIT('h0001)
	) name3258 (
		_w13767_,
		_w13768_,
		_w13769_,
		_w13770_,
		_w13771_
	);
	LUT3 #(
		.INIT('h80)
	) name3259 (
		\wishbone_bd_ram_mem1_reg[221][15]/P0001 ,
		_w11966_,
		_w11984_,
		_w13772_
	);
	LUT3 #(
		.INIT('h80)
	) name3260 (
		\wishbone_bd_ram_mem1_reg[30][15]/P0001 ,
		_w11935_,
		_w11948_,
		_w13773_
	);
	LUT3 #(
		.INIT('h80)
	) name3261 (
		\wishbone_bd_ram_mem1_reg[116][15]/P0001 ,
		_w11929_,
		_w12012_,
		_w13774_
	);
	LUT3 #(
		.INIT('h80)
	) name3262 (
		\wishbone_bd_ram_mem1_reg[224][15]/P0001 ,
		_w11941_,
		_w11982_,
		_w13775_
	);
	LUT4 #(
		.INIT('h0001)
	) name3263 (
		_w13772_,
		_w13773_,
		_w13774_,
		_w13775_,
		_w13776_
	);
	LUT4 #(
		.INIT('h8000)
	) name3264 (
		_w13761_,
		_w13766_,
		_w13771_,
		_w13776_,
		_w13777_
	);
	LUT3 #(
		.INIT('h80)
	) name3265 (
		\wishbone_bd_ram_mem1_reg[211][15]/P0001 ,
		_w11938_,
		_w11984_,
		_w13778_
	);
	LUT3 #(
		.INIT('h80)
	) name3266 (
		\wishbone_bd_ram_mem1_reg[165][15]/P0001 ,
		_w11930_,
		_w11933_,
		_w13779_
	);
	LUT3 #(
		.INIT('h80)
	) name3267 (
		\wishbone_bd_ram_mem1_reg[131][15]/P0001 ,
		_w11938_,
		_w11955_,
		_w13780_
	);
	LUT3 #(
		.INIT('h80)
	) name3268 (
		\wishbone_bd_ram_mem1_reg[107][15]/P0001 ,
		_w11936_,
		_w11965_,
		_w13781_
	);
	LUT4 #(
		.INIT('h0001)
	) name3269 (
		_w13778_,
		_w13779_,
		_w13780_,
		_w13781_,
		_w13782_
	);
	LUT3 #(
		.INIT('h80)
	) name3270 (
		\wishbone_bd_ram_mem1_reg[246][15]/P0001 ,
		_w11952_,
		_w11986_,
		_w13783_
	);
	LUT3 #(
		.INIT('h80)
	) name3271 (
		\wishbone_bd_ram_mem1_reg[205][15]/P0001 ,
		_w11945_,
		_w11966_,
		_w13784_
	);
	LUT3 #(
		.INIT('h80)
	) name3272 (
		\wishbone_bd_ram_mem1_reg[210][15]/P0001 ,
		_w11963_,
		_w11984_,
		_w13785_
	);
	LUT3 #(
		.INIT('h80)
	) name3273 (
		\wishbone_bd_ram_mem1_reg[0][15]/P0001 ,
		_w11932_,
		_w11941_,
		_w13786_
	);
	LUT4 #(
		.INIT('h0001)
	) name3274 (
		_w13783_,
		_w13784_,
		_w13785_,
		_w13786_,
		_w13787_
	);
	LUT3 #(
		.INIT('h80)
	) name3275 (
		\wishbone_bd_ram_mem1_reg[99][15]/P0001 ,
		_w11938_,
		_w11965_,
		_w13788_
	);
	LUT3 #(
		.INIT('h80)
	) name3276 (
		\wishbone_bd_ram_mem1_reg[168][15]/P0001 ,
		_w11930_,
		_w11990_,
		_w13789_
	);
	LUT3 #(
		.INIT('h80)
	) name3277 (
		\wishbone_bd_ram_mem1_reg[36][15]/P0001 ,
		_w11929_,
		_w11957_,
		_w13790_
	);
	LUT3 #(
		.INIT('h80)
	) name3278 (
		\wishbone_bd_ram_mem1_reg[214][15]/P0001 ,
		_w11984_,
		_w11986_,
		_w13791_
	);
	LUT4 #(
		.INIT('h0001)
	) name3279 (
		_w13788_,
		_w13789_,
		_w13790_,
		_w13791_,
		_w13792_
	);
	LUT3 #(
		.INIT('h80)
	) name3280 (
		\wishbone_bd_ram_mem1_reg[66][15]/P0001 ,
		_w11949_,
		_w11963_,
		_w13793_
	);
	LUT3 #(
		.INIT('h80)
	) name3281 (
		\wishbone_bd_ram_mem1_reg[35][15]/P0001 ,
		_w11938_,
		_w11957_,
		_w13794_
	);
	LUT3 #(
		.INIT('h80)
	) name3282 (
		\wishbone_bd_ram_mem1_reg[40][15]/P0001 ,
		_w11957_,
		_w11990_,
		_w13795_
	);
	LUT3 #(
		.INIT('h80)
	) name3283 (
		\wishbone_bd_ram_mem1_reg[143][15]/P0001 ,
		_w11955_,
		_w11973_,
		_w13796_
	);
	LUT4 #(
		.INIT('h0001)
	) name3284 (
		_w13793_,
		_w13794_,
		_w13795_,
		_w13796_,
		_w13797_
	);
	LUT4 #(
		.INIT('h8000)
	) name3285 (
		_w13782_,
		_w13787_,
		_w13792_,
		_w13797_,
		_w13798_
	);
	LUT4 #(
		.INIT('h8000)
	) name3286 (
		_w13735_,
		_w13756_,
		_w13777_,
		_w13798_,
		_w13799_
	);
	LUT4 #(
		.INIT('h8000)
	) name3287 (
		_w13544_,
		_w13629_,
		_w13714_,
		_w13799_,
		_w13800_
	);
	LUT3 #(
		.INIT('h54)
	) name3288 (
		wb_rst_i_pad,
		_w13457_,
		_w13458_,
		_w13801_
	);
	LUT3 #(
		.INIT('hba)
	) name3289 (
		_w13459_,
		_w13800_,
		_w13801_,
		_w13802_
	);
	LUT2 #(
		.INIT('h2)
	) name3290 (
		\wishbone_RxDataLatched2_reg[9]/NET0131 ,
		_w13424_,
		_w13803_
	);
	LUT2 #(
		.INIT('h8)
	) name3291 (
		_w13423_,
		_w13803_,
		_w13804_
	);
	LUT3 #(
		.INIT('ha2)
	) name3292 (
		\wishbone_RxDataLatched1_reg[9]/NET0131 ,
		_w13423_,
		_w13424_,
		_w13805_
	);
	LUT3 #(
		.INIT('hdc)
	) name3293 (
		_w13428_,
		_w13804_,
		_w13805_,
		_w13806_
	);
	LUT3 #(
		.INIT('h80)
	) name3294 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w13807_
	);
	LUT4 #(
		.INIT('h070f)
	) name3295 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w13808_
	);
	LUT2 #(
		.INIT('h8)
	) name3296 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		_w13809_
	);
	LUT3 #(
		.INIT('h02)
	) name3297 (
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w13807_,
		_w13809_,
		_w13810_
	);
	LUT3 #(
		.INIT('h80)
	) name3298 (
		\wishbone_bd_ram_mem0_reg[166][1]/P0001 ,
		_w11930_,
		_w11986_,
		_w13811_
	);
	LUT3 #(
		.INIT('h80)
	) name3299 (
		\wishbone_bd_ram_mem0_reg[57][1]/P0001 ,
		_w11968_,
		_w11979_,
		_w13812_
	);
	LUT3 #(
		.INIT('h80)
	) name3300 (
		\wishbone_bd_ram_mem0_reg[50][1]/P0001 ,
		_w11963_,
		_w11979_,
		_w13813_
	);
	LUT3 #(
		.INIT('h80)
	) name3301 (
		\wishbone_bd_ram_mem0_reg[216][1]/P0001 ,
		_w11984_,
		_w11990_,
		_w13814_
	);
	LUT4 #(
		.INIT('h0001)
	) name3302 (
		_w13811_,
		_w13812_,
		_w13813_,
		_w13814_,
		_w13815_
	);
	LUT3 #(
		.INIT('h80)
	) name3303 (
		\wishbone_bd_ram_mem0_reg[201][1]/P0001 ,
		_w11945_,
		_w11968_,
		_w13816_
	);
	LUT3 #(
		.INIT('h80)
	) name3304 (
		\wishbone_bd_ram_mem0_reg[122][1]/P0001 ,
		_w11944_,
		_w12012_,
		_w13817_
	);
	LUT3 #(
		.INIT('h80)
	) name3305 (
		\wishbone_bd_ram_mem0_reg[130][1]/P0001 ,
		_w11955_,
		_w11963_,
		_w13818_
	);
	LUT3 #(
		.INIT('h80)
	) name3306 (
		\wishbone_bd_ram_mem0_reg[13][1]/P0001 ,
		_w11932_,
		_w11966_,
		_w13819_
	);
	LUT4 #(
		.INIT('h0001)
	) name3307 (
		_w13816_,
		_w13817_,
		_w13818_,
		_w13819_,
		_w13820_
	);
	LUT3 #(
		.INIT('h80)
	) name3308 (
		\wishbone_bd_ram_mem0_reg[19][1]/P0001 ,
		_w11935_,
		_w11938_,
		_w13821_
	);
	LUT3 #(
		.INIT('h80)
	) name3309 (
		\wishbone_bd_ram_mem0_reg[40][1]/P0001 ,
		_w11957_,
		_w11990_,
		_w13822_
	);
	LUT3 #(
		.INIT('h80)
	) name3310 (
		\wishbone_bd_ram_mem0_reg[126][1]/P0001 ,
		_w11948_,
		_w12012_,
		_w13823_
	);
	LUT3 #(
		.INIT('h80)
	) name3311 (
		\wishbone_bd_ram_mem0_reg[222][1]/P0001 ,
		_w11948_,
		_w11984_,
		_w13824_
	);
	LUT4 #(
		.INIT('h0001)
	) name3312 (
		_w13821_,
		_w13822_,
		_w13823_,
		_w13824_,
		_w13825_
	);
	LUT3 #(
		.INIT('h80)
	) name3313 (
		\wishbone_bd_ram_mem0_reg[249][1]/P0001 ,
		_w11952_,
		_w11968_,
		_w13826_
	);
	LUT3 #(
		.INIT('h80)
	) name3314 (
		\wishbone_bd_ram_mem0_reg[241][1]/P0001 ,
		_w11952_,
		_w11977_,
		_w13827_
	);
	LUT3 #(
		.INIT('h80)
	) name3315 (
		\wishbone_bd_ram_mem0_reg[168][1]/P0001 ,
		_w11930_,
		_w11990_,
		_w13828_
	);
	LUT3 #(
		.INIT('h80)
	) name3316 (
		\wishbone_bd_ram_mem0_reg[244][1]/P0001 ,
		_w11929_,
		_w11952_,
		_w13829_
	);
	LUT4 #(
		.INIT('h0001)
	) name3317 (
		_w13826_,
		_w13827_,
		_w13828_,
		_w13829_,
		_w13830_
	);
	LUT4 #(
		.INIT('h8000)
	) name3318 (
		_w13815_,
		_w13820_,
		_w13825_,
		_w13830_,
		_w13831_
	);
	LUT3 #(
		.INIT('h80)
	) name3319 (
		\wishbone_bd_ram_mem0_reg[44][1]/P0001 ,
		_w11954_,
		_w11957_,
		_w13832_
	);
	LUT3 #(
		.INIT('h80)
	) name3320 (
		\wishbone_bd_ram_mem0_reg[33][1]/P0001 ,
		_w11957_,
		_w11977_,
		_w13833_
	);
	LUT3 #(
		.INIT('h80)
	) name3321 (
		\wishbone_bd_ram_mem0_reg[17][1]/P0001 ,
		_w11935_,
		_w11977_,
		_w13834_
	);
	LUT3 #(
		.INIT('h80)
	) name3322 (
		\wishbone_bd_ram_mem0_reg[31][1]/P0001 ,
		_w11935_,
		_w11973_,
		_w13835_
	);
	LUT4 #(
		.INIT('h0001)
	) name3323 (
		_w13832_,
		_w13833_,
		_w13834_,
		_w13835_,
		_w13836_
	);
	LUT3 #(
		.INIT('h80)
	) name3324 (
		\wishbone_bd_ram_mem0_reg[7][1]/P0001 ,
		_w11932_,
		_w11975_,
		_w13837_
	);
	LUT3 #(
		.INIT('h80)
	) name3325 (
		\wishbone_bd_ram_mem0_reg[21][1]/P0001 ,
		_w11933_,
		_w11935_,
		_w13838_
	);
	LUT3 #(
		.INIT('h80)
	) name3326 (
		\wishbone_bd_ram_mem0_reg[217][1]/P0001 ,
		_w11968_,
		_w11984_,
		_w13839_
	);
	LUT3 #(
		.INIT('h80)
	) name3327 (
		\wishbone_bd_ram_mem0_reg[85][1]/P0001 ,
		_w11933_,
		_w11972_,
		_w13840_
	);
	LUT4 #(
		.INIT('h0001)
	) name3328 (
		_w13837_,
		_w13838_,
		_w13839_,
		_w13840_,
		_w13841_
	);
	LUT3 #(
		.INIT('h80)
	) name3329 (
		\wishbone_bd_ram_mem0_reg[84][1]/P0001 ,
		_w11929_,
		_w11972_,
		_w13842_
	);
	LUT3 #(
		.INIT('h80)
	) name3330 (
		\wishbone_bd_ram_mem0_reg[35][1]/P0001 ,
		_w11938_,
		_w11957_,
		_w13843_
	);
	LUT3 #(
		.INIT('h80)
	) name3331 (
		\wishbone_bd_ram_mem0_reg[187][1]/P0001 ,
		_w11936_,
		_w11942_,
		_w13844_
	);
	LUT3 #(
		.INIT('h80)
	) name3332 (
		\wishbone_bd_ram_mem0_reg[205][1]/P0001 ,
		_w11945_,
		_w11966_,
		_w13845_
	);
	LUT4 #(
		.INIT('h0001)
	) name3333 (
		_w13842_,
		_w13843_,
		_w13844_,
		_w13845_,
		_w13846_
	);
	LUT3 #(
		.INIT('h80)
	) name3334 (
		\wishbone_bd_ram_mem0_reg[3][1]/P0001 ,
		_w11932_,
		_w11938_,
		_w13847_
	);
	LUT3 #(
		.INIT('h80)
	) name3335 (
		\wishbone_bd_ram_mem0_reg[79][1]/P0001 ,
		_w11949_,
		_w11973_,
		_w13848_
	);
	LUT3 #(
		.INIT('h80)
	) name3336 (
		\wishbone_bd_ram_mem0_reg[149][1]/P0001 ,
		_w11933_,
		_w11959_,
		_w13849_
	);
	LUT3 #(
		.INIT('h80)
	) name3337 (
		\wishbone_bd_ram_mem0_reg[46][1]/P0001 ,
		_w11948_,
		_w11957_,
		_w13850_
	);
	LUT4 #(
		.INIT('h0001)
	) name3338 (
		_w13847_,
		_w13848_,
		_w13849_,
		_w13850_,
		_w13851_
	);
	LUT4 #(
		.INIT('h8000)
	) name3339 (
		_w13836_,
		_w13841_,
		_w13846_,
		_w13851_,
		_w13852_
	);
	LUT3 #(
		.INIT('h80)
	) name3340 (
		\wishbone_bd_ram_mem0_reg[114][1]/P0001 ,
		_w11963_,
		_w12012_,
		_w13853_
	);
	LUT3 #(
		.INIT('h80)
	) name3341 (
		\wishbone_bd_ram_mem0_reg[226][1]/P0001 ,
		_w11963_,
		_w11982_,
		_w13854_
	);
	LUT3 #(
		.INIT('h80)
	) name3342 (
		\wishbone_bd_ram_mem0_reg[87][1]/P0001 ,
		_w11972_,
		_w11975_,
		_w13855_
	);
	LUT3 #(
		.INIT('h80)
	) name3343 (
		\wishbone_bd_ram_mem0_reg[170][1]/P0001 ,
		_w11930_,
		_w11944_,
		_w13856_
	);
	LUT4 #(
		.INIT('h0001)
	) name3344 (
		_w13853_,
		_w13854_,
		_w13855_,
		_w13856_,
		_w13857_
	);
	LUT3 #(
		.INIT('h80)
	) name3345 (
		\wishbone_bd_ram_mem0_reg[125][1]/P0001 ,
		_w11966_,
		_w12012_,
		_w13858_
	);
	LUT3 #(
		.INIT('h80)
	) name3346 (
		\wishbone_bd_ram_mem0_reg[88][1]/P0001 ,
		_w11972_,
		_w11990_,
		_w13859_
	);
	LUT3 #(
		.INIT('h80)
	) name3347 (
		\wishbone_bd_ram_mem0_reg[159][1]/P0001 ,
		_w11959_,
		_w11973_,
		_w13860_
	);
	LUT3 #(
		.INIT('h80)
	) name3348 (
		\wishbone_bd_ram_mem0_reg[62][1]/P0001 ,
		_w11948_,
		_w11979_,
		_w13861_
	);
	LUT4 #(
		.INIT('h0001)
	) name3349 (
		_w13858_,
		_w13859_,
		_w13860_,
		_w13861_,
		_w13862_
	);
	LUT3 #(
		.INIT('h80)
	) name3350 (
		\wishbone_bd_ram_mem0_reg[242][1]/P0001 ,
		_w11952_,
		_w11963_,
		_w13863_
	);
	LUT3 #(
		.INIT('h80)
	) name3351 (
		\wishbone_bd_ram_mem0_reg[245][1]/P0001 ,
		_w11933_,
		_w11952_,
		_w13864_
	);
	LUT3 #(
		.INIT('h80)
	) name3352 (
		\wishbone_bd_ram_mem0_reg[123][1]/P0001 ,
		_w11936_,
		_w12012_,
		_w13865_
	);
	LUT3 #(
		.INIT('h80)
	) name3353 (
		\wishbone_bd_ram_mem0_reg[250][1]/P0001 ,
		_w11944_,
		_w11952_,
		_w13866_
	);
	LUT4 #(
		.INIT('h0001)
	) name3354 (
		_w13863_,
		_w13864_,
		_w13865_,
		_w13866_,
		_w13867_
	);
	LUT3 #(
		.INIT('h80)
	) name3355 (
		\wishbone_bd_ram_mem0_reg[109][1]/P0001 ,
		_w11965_,
		_w11966_,
		_w13868_
	);
	LUT3 #(
		.INIT('h80)
	) name3356 (
		\wishbone_bd_ram_mem0_reg[22][1]/P0001 ,
		_w11935_,
		_w11986_,
		_w13869_
	);
	LUT3 #(
		.INIT('h80)
	) name3357 (
		\wishbone_bd_ram_mem0_reg[107][1]/P0001 ,
		_w11936_,
		_w11965_,
		_w13870_
	);
	LUT3 #(
		.INIT('h80)
	) name3358 (
		\wishbone_bd_ram_mem0_reg[184][1]/P0001 ,
		_w11942_,
		_w11990_,
		_w13871_
	);
	LUT4 #(
		.INIT('h0001)
	) name3359 (
		_w13868_,
		_w13869_,
		_w13870_,
		_w13871_,
		_w13872_
	);
	LUT4 #(
		.INIT('h8000)
	) name3360 (
		_w13857_,
		_w13862_,
		_w13867_,
		_w13872_,
		_w13873_
	);
	LUT3 #(
		.INIT('h80)
	) name3361 (
		\wishbone_bd_ram_mem0_reg[63][1]/P0001 ,
		_w11973_,
		_w11979_,
		_w13874_
	);
	LUT3 #(
		.INIT('h80)
	) name3362 (
		\wishbone_bd_ram_mem0_reg[135][1]/P0001 ,
		_w11955_,
		_w11975_,
		_w13875_
	);
	LUT3 #(
		.INIT('h80)
	) name3363 (
		\wishbone_bd_ram_mem0_reg[58][1]/P0001 ,
		_w11944_,
		_w11979_,
		_w13876_
	);
	LUT3 #(
		.INIT('h80)
	) name3364 (
		\wishbone_bd_ram_mem0_reg[175][1]/P0001 ,
		_w11930_,
		_w11973_,
		_w13877_
	);
	LUT4 #(
		.INIT('h0001)
	) name3365 (
		_w13874_,
		_w13875_,
		_w13876_,
		_w13877_,
		_w13878_
	);
	LUT3 #(
		.INIT('h80)
	) name3366 (
		\wishbone_bd_ram_mem0_reg[55][1]/P0001 ,
		_w11975_,
		_w11979_,
		_w13879_
	);
	LUT3 #(
		.INIT('h80)
	) name3367 (
		\wishbone_bd_ram_mem0_reg[18][1]/P0001 ,
		_w11935_,
		_w11963_,
		_w13880_
	);
	LUT3 #(
		.INIT('h80)
	) name3368 (
		\wishbone_bd_ram_mem0_reg[47][1]/P0001 ,
		_w11957_,
		_w11973_,
		_w13881_
	);
	LUT3 #(
		.INIT('h80)
	) name3369 (
		\wishbone_bd_ram_mem0_reg[143][1]/P0001 ,
		_w11955_,
		_w11973_,
		_w13882_
	);
	LUT4 #(
		.INIT('h0001)
	) name3370 (
		_w13879_,
		_w13880_,
		_w13881_,
		_w13882_,
		_w13883_
	);
	LUT3 #(
		.INIT('h80)
	) name3371 (
		\wishbone_bd_ram_mem0_reg[225][1]/P0001 ,
		_w11977_,
		_w11982_,
		_w13884_
	);
	LUT3 #(
		.INIT('h80)
	) name3372 (
		\wishbone_bd_ram_mem0_reg[27][1]/P0001 ,
		_w11935_,
		_w11936_,
		_w13885_
	);
	LUT3 #(
		.INIT('h80)
	) name3373 (
		\wishbone_bd_ram_mem0_reg[124][1]/P0001 ,
		_w11954_,
		_w12012_,
		_w13886_
	);
	LUT3 #(
		.INIT('h80)
	) name3374 (
		\wishbone_bd_ram_mem0_reg[177][1]/P0001 ,
		_w11942_,
		_w11977_,
		_w13887_
	);
	LUT4 #(
		.INIT('h0001)
	) name3375 (
		_w13884_,
		_w13885_,
		_w13886_,
		_w13887_,
		_w13888_
	);
	LUT3 #(
		.INIT('h80)
	) name3376 (
		\wishbone_bd_ram_mem0_reg[214][1]/P0001 ,
		_w11984_,
		_w11986_,
		_w13889_
	);
	LUT3 #(
		.INIT('h80)
	) name3377 (
		\wishbone_bd_ram_mem0_reg[196][1]/P0001 ,
		_w11929_,
		_w11945_,
		_w13890_
	);
	LUT3 #(
		.INIT('h80)
	) name3378 (
		\wishbone_bd_ram_mem0_reg[1][1]/P0001 ,
		_w11932_,
		_w11977_,
		_w13891_
	);
	LUT3 #(
		.INIT('h80)
	) name3379 (
		\wishbone_bd_ram_mem0_reg[160][1]/P0001 ,
		_w11930_,
		_w11941_,
		_w13892_
	);
	LUT4 #(
		.INIT('h0001)
	) name3380 (
		_w13889_,
		_w13890_,
		_w13891_,
		_w13892_,
		_w13893_
	);
	LUT4 #(
		.INIT('h8000)
	) name3381 (
		_w13878_,
		_w13883_,
		_w13888_,
		_w13893_,
		_w13894_
	);
	LUT4 #(
		.INIT('h8000)
	) name3382 (
		_w13831_,
		_w13852_,
		_w13873_,
		_w13894_,
		_w13895_
	);
	LUT3 #(
		.INIT('h80)
	) name3383 (
		\wishbone_bd_ram_mem0_reg[231][1]/P0001 ,
		_w11975_,
		_w11982_,
		_w13896_
	);
	LUT3 #(
		.INIT('h80)
	) name3384 (
		\wishbone_bd_ram_mem0_reg[45][1]/P0001 ,
		_w11957_,
		_w11966_,
		_w13897_
	);
	LUT3 #(
		.INIT('h80)
	) name3385 (
		\wishbone_bd_ram_mem0_reg[220][1]/P0001 ,
		_w11954_,
		_w11984_,
		_w13898_
	);
	LUT3 #(
		.INIT('h80)
	) name3386 (
		\wishbone_bd_ram_mem0_reg[145][1]/P0001 ,
		_w11959_,
		_w11977_,
		_w13899_
	);
	LUT4 #(
		.INIT('h0001)
	) name3387 (
		_w13896_,
		_w13897_,
		_w13898_,
		_w13899_,
		_w13900_
	);
	LUT3 #(
		.INIT('h80)
	) name3388 (
		\wishbone_bd_ram_mem0_reg[230][1]/P0001 ,
		_w11982_,
		_w11986_,
		_w13901_
	);
	LUT3 #(
		.INIT('h80)
	) name3389 (
		\wishbone_bd_ram_mem0_reg[111][1]/P0001 ,
		_w11965_,
		_w11973_,
		_w13902_
	);
	LUT3 #(
		.INIT('h80)
	) name3390 (
		\wishbone_bd_ram_mem0_reg[199][1]/P0001 ,
		_w11945_,
		_w11975_,
		_w13903_
	);
	LUT3 #(
		.INIT('h80)
	) name3391 (
		\wishbone_bd_ram_mem0_reg[146][1]/P0001 ,
		_w11959_,
		_w11963_,
		_w13904_
	);
	LUT4 #(
		.INIT('h0001)
	) name3392 (
		_w13901_,
		_w13902_,
		_w13903_,
		_w13904_,
		_w13905_
	);
	LUT3 #(
		.INIT('h80)
	) name3393 (
		\wishbone_bd_ram_mem0_reg[215][1]/P0001 ,
		_w11975_,
		_w11984_,
		_w13906_
	);
	LUT3 #(
		.INIT('h80)
	) name3394 (
		\wishbone_bd_ram_mem0_reg[238][1]/P0001 ,
		_w11948_,
		_w11982_,
		_w13907_
	);
	LUT3 #(
		.INIT('h80)
	) name3395 (
		\wishbone_bd_ram_mem0_reg[252][1]/P0001 ,
		_w11952_,
		_w11954_,
		_w13908_
	);
	LUT3 #(
		.INIT('h80)
	) name3396 (
		\wishbone_bd_ram_mem0_reg[52][1]/P0001 ,
		_w11929_,
		_w11979_,
		_w13909_
	);
	LUT4 #(
		.INIT('h0001)
	) name3397 (
		_w13906_,
		_w13907_,
		_w13908_,
		_w13909_,
		_w13910_
	);
	LUT3 #(
		.INIT('h80)
	) name3398 (
		\wishbone_bd_ram_mem0_reg[53][1]/P0001 ,
		_w11933_,
		_w11979_,
		_w13911_
	);
	LUT3 #(
		.INIT('h80)
	) name3399 (
		\wishbone_bd_ram_mem0_reg[69][1]/P0001 ,
		_w11933_,
		_w11949_,
		_w13912_
	);
	LUT3 #(
		.INIT('h80)
	) name3400 (
		\wishbone_bd_ram_mem0_reg[42][1]/P0001 ,
		_w11944_,
		_w11957_,
		_w13913_
	);
	LUT3 #(
		.INIT('h80)
	) name3401 (
		\wishbone_bd_ram_mem0_reg[213][1]/P0001 ,
		_w11933_,
		_w11984_,
		_w13914_
	);
	LUT4 #(
		.INIT('h0001)
	) name3402 (
		_w13911_,
		_w13912_,
		_w13913_,
		_w13914_,
		_w13915_
	);
	LUT4 #(
		.INIT('h8000)
	) name3403 (
		_w13900_,
		_w13905_,
		_w13910_,
		_w13915_,
		_w13916_
	);
	LUT3 #(
		.INIT('h80)
	) name3404 (
		\wishbone_bd_ram_mem0_reg[197][1]/P0001 ,
		_w11933_,
		_w11945_,
		_w13917_
	);
	LUT3 #(
		.INIT('h80)
	) name3405 (
		\wishbone_bd_ram_mem0_reg[16][1]/P0001 ,
		_w11935_,
		_w11941_,
		_w13918_
	);
	LUT3 #(
		.INIT('h80)
	) name3406 (
		\wishbone_bd_ram_mem0_reg[2][1]/P0001 ,
		_w11932_,
		_w11963_,
		_w13919_
	);
	LUT3 #(
		.INIT('h80)
	) name3407 (
		\wishbone_bd_ram_mem0_reg[198][1]/P0001 ,
		_w11945_,
		_w11986_,
		_w13920_
	);
	LUT4 #(
		.INIT('h0001)
	) name3408 (
		_w13917_,
		_w13918_,
		_w13919_,
		_w13920_,
		_w13921_
	);
	LUT3 #(
		.INIT('h80)
	) name3409 (
		\wishbone_bd_ram_mem0_reg[108][1]/P0001 ,
		_w11954_,
		_w11965_,
		_w13922_
	);
	LUT3 #(
		.INIT('h80)
	) name3410 (
		\wishbone_bd_ram_mem0_reg[200][1]/P0001 ,
		_w11945_,
		_w11990_,
		_w13923_
	);
	LUT3 #(
		.INIT('h80)
	) name3411 (
		\wishbone_bd_ram_mem0_reg[90][1]/P0001 ,
		_w11944_,
		_w11972_,
		_w13924_
	);
	LUT3 #(
		.INIT('h80)
	) name3412 (
		\wishbone_bd_ram_mem0_reg[247][1]/P0001 ,
		_w11952_,
		_w11975_,
		_w13925_
	);
	LUT4 #(
		.INIT('h0001)
	) name3413 (
		_w13922_,
		_w13923_,
		_w13924_,
		_w13925_,
		_w13926_
	);
	LUT3 #(
		.INIT('h80)
	) name3414 (
		\wishbone_bd_ram_mem0_reg[72][1]/P0001 ,
		_w11949_,
		_w11990_,
		_w13927_
	);
	LUT3 #(
		.INIT('h80)
	) name3415 (
		\wishbone_bd_ram_mem0_reg[163][1]/P0001 ,
		_w11930_,
		_w11938_,
		_w13928_
	);
	LUT3 #(
		.INIT('h80)
	) name3416 (
		\wishbone_bd_ram_mem0_reg[161][1]/P0001 ,
		_w11930_,
		_w11977_,
		_w13929_
	);
	LUT3 #(
		.INIT('h80)
	) name3417 (
		\wishbone_bd_ram_mem0_reg[75][1]/P0001 ,
		_w11936_,
		_w11949_,
		_w13930_
	);
	LUT4 #(
		.INIT('h0001)
	) name3418 (
		_w13927_,
		_w13928_,
		_w13929_,
		_w13930_,
		_w13931_
	);
	LUT3 #(
		.INIT('h80)
	) name3419 (
		\wishbone_bd_ram_mem0_reg[60][1]/P0001 ,
		_w11954_,
		_w11979_,
		_w13932_
	);
	LUT3 #(
		.INIT('h80)
	) name3420 (
		\wishbone_bd_ram_mem0_reg[229][1]/P0001 ,
		_w11933_,
		_w11982_,
		_w13933_
	);
	LUT3 #(
		.INIT('h80)
	) name3421 (
		\wishbone_bd_ram_mem0_reg[104][1]/P0001 ,
		_w11965_,
		_w11990_,
		_w13934_
	);
	LUT3 #(
		.INIT('h80)
	) name3422 (
		\wishbone_bd_ram_mem0_reg[11][1]/P0001 ,
		_w11932_,
		_w11936_,
		_w13935_
	);
	LUT4 #(
		.INIT('h0001)
	) name3423 (
		_w13932_,
		_w13933_,
		_w13934_,
		_w13935_,
		_w13936_
	);
	LUT4 #(
		.INIT('h8000)
	) name3424 (
		_w13921_,
		_w13926_,
		_w13931_,
		_w13936_,
		_w13937_
	);
	LUT3 #(
		.INIT('h80)
	) name3425 (
		\wishbone_bd_ram_mem0_reg[115][1]/P0001 ,
		_w11938_,
		_w12012_,
		_w13938_
	);
	LUT3 #(
		.INIT('h80)
	) name3426 (
		\wishbone_bd_ram_mem0_reg[100][1]/P0001 ,
		_w11929_,
		_w11965_,
		_w13939_
	);
	LUT3 #(
		.INIT('h80)
	) name3427 (
		\wishbone_bd_ram_mem0_reg[38][1]/P0001 ,
		_w11957_,
		_w11986_,
		_w13940_
	);
	LUT3 #(
		.INIT('h80)
	) name3428 (
		\wishbone_bd_ram_mem0_reg[12][1]/P0001 ,
		_w11932_,
		_w11954_,
		_w13941_
	);
	LUT4 #(
		.INIT('h0001)
	) name3429 (
		_w13938_,
		_w13939_,
		_w13940_,
		_w13941_,
		_w13942_
	);
	LUT3 #(
		.INIT('h80)
	) name3430 (
		\wishbone_bd_ram_mem0_reg[174][1]/P0001 ,
		_w11930_,
		_w11948_,
		_w13943_
	);
	LUT3 #(
		.INIT('h80)
	) name3431 (
		\wishbone_bd_ram_mem0_reg[105][1]/P0001 ,
		_w11965_,
		_w11968_,
		_w13944_
	);
	LUT3 #(
		.INIT('h80)
	) name3432 (
		\wishbone_bd_ram_mem0_reg[127][1]/P0001 ,
		_w11973_,
		_w12012_,
		_w13945_
	);
	LUT3 #(
		.INIT('h80)
	) name3433 (
		\wishbone_bd_ram_mem0_reg[140][1]/P0001 ,
		_w11954_,
		_w11955_,
		_w13946_
	);
	LUT4 #(
		.INIT('h0001)
	) name3434 (
		_w13943_,
		_w13944_,
		_w13945_,
		_w13946_,
		_w13947_
	);
	LUT3 #(
		.INIT('h80)
	) name3435 (
		\wishbone_bd_ram_mem0_reg[181][1]/P0001 ,
		_w11933_,
		_w11942_,
		_w13948_
	);
	LUT3 #(
		.INIT('h80)
	) name3436 (
		\wishbone_bd_ram_mem0_reg[151][1]/P0001 ,
		_w11959_,
		_w11975_,
		_w13949_
	);
	LUT3 #(
		.INIT('h80)
	) name3437 (
		\wishbone_bd_ram_mem0_reg[167][1]/P0001 ,
		_w11930_,
		_w11975_,
		_w13950_
	);
	LUT3 #(
		.INIT('h80)
	) name3438 (
		\wishbone_bd_ram_mem0_reg[171][1]/P0001 ,
		_w11930_,
		_w11936_,
		_w13951_
	);
	LUT4 #(
		.INIT('h0001)
	) name3439 (
		_w13948_,
		_w13949_,
		_w13950_,
		_w13951_,
		_w13952_
	);
	LUT3 #(
		.INIT('h80)
	) name3440 (
		\wishbone_bd_ram_mem0_reg[95][1]/P0001 ,
		_w11972_,
		_w11973_,
		_w13953_
	);
	LUT3 #(
		.INIT('h80)
	) name3441 (
		\wishbone_bd_ram_mem0_reg[14][1]/P0001 ,
		_w11932_,
		_w11948_,
		_w13954_
	);
	LUT3 #(
		.INIT('h80)
	) name3442 (
		\wishbone_bd_ram_mem0_reg[248][1]/P0001 ,
		_w11952_,
		_w11990_,
		_w13955_
	);
	LUT3 #(
		.INIT('h80)
	) name3443 (
		\wishbone_bd_ram_mem0_reg[190][1]/P0001 ,
		_w11942_,
		_w11948_,
		_w13956_
	);
	LUT4 #(
		.INIT('h0001)
	) name3444 (
		_w13953_,
		_w13954_,
		_w13955_,
		_w13956_,
		_w13957_
	);
	LUT4 #(
		.INIT('h8000)
	) name3445 (
		_w13942_,
		_w13947_,
		_w13952_,
		_w13957_,
		_w13958_
	);
	LUT3 #(
		.INIT('h80)
	) name3446 (
		\wishbone_bd_ram_mem0_reg[34][1]/P0001 ,
		_w11957_,
		_w11963_,
		_w13959_
	);
	LUT3 #(
		.INIT('h80)
	) name3447 (
		\wishbone_bd_ram_mem0_reg[137][1]/P0001 ,
		_w11955_,
		_w11968_,
		_w13960_
	);
	LUT3 #(
		.INIT('h80)
	) name3448 (
		\wishbone_bd_ram_mem0_reg[59][1]/P0001 ,
		_w11936_,
		_w11979_,
		_w13961_
	);
	LUT3 #(
		.INIT('h80)
	) name3449 (
		\wishbone_bd_ram_mem0_reg[94][1]/P0001 ,
		_w11948_,
		_w11972_,
		_w13962_
	);
	LUT4 #(
		.INIT('h0001)
	) name3450 (
		_w13959_,
		_w13960_,
		_w13961_,
		_w13962_,
		_w13963_
	);
	LUT3 #(
		.INIT('h80)
	) name3451 (
		\wishbone_bd_ram_mem0_reg[54][1]/P0001 ,
		_w11979_,
		_w11986_,
		_w13964_
	);
	LUT3 #(
		.INIT('h80)
	) name3452 (
		\wishbone_bd_ram_mem0_reg[73][1]/P0001 ,
		_w11949_,
		_w11968_,
		_w13965_
	);
	LUT3 #(
		.INIT('h80)
	) name3453 (
		\wishbone_bd_ram_mem0_reg[129][1]/P0001 ,
		_w11955_,
		_w11977_,
		_w13966_
	);
	LUT3 #(
		.INIT('h80)
	) name3454 (
		\wishbone_bd_ram_mem0_reg[91][1]/P0001 ,
		_w11936_,
		_w11972_,
		_w13967_
	);
	LUT4 #(
		.INIT('h0001)
	) name3455 (
		_w13964_,
		_w13965_,
		_w13966_,
		_w13967_,
		_w13968_
	);
	LUT3 #(
		.INIT('h80)
	) name3456 (
		\wishbone_bd_ram_mem0_reg[141][1]/P0001 ,
		_w11955_,
		_w11966_,
		_w13969_
	);
	LUT3 #(
		.INIT('h80)
	) name3457 (
		\wishbone_bd_ram_mem0_reg[193][1]/P0001 ,
		_w11945_,
		_w11977_,
		_w13970_
	);
	LUT3 #(
		.INIT('h80)
	) name3458 (
		\wishbone_bd_ram_mem0_reg[51][1]/P0001 ,
		_w11938_,
		_w11979_,
		_w13971_
	);
	LUT3 #(
		.INIT('h80)
	) name3459 (
		\wishbone_bd_ram_mem0_reg[218][1]/P0001 ,
		_w11944_,
		_w11984_,
		_w13972_
	);
	LUT4 #(
		.INIT('h0001)
	) name3460 (
		_w13969_,
		_w13970_,
		_w13971_,
		_w13972_,
		_w13973_
	);
	LUT3 #(
		.INIT('h80)
	) name3461 (
		\wishbone_bd_ram_mem0_reg[5][1]/P0001 ,
		_w11932_,
		_w11933_,
		_w13974_
	);
	LUT3 #(
		.INIT('h80)
	) name3462 (
		\wishbone_bd_ram_mem0_reg[155][1]/P0001 ,
		_w11936_,
		_w11959_,
		_w13975_
	);
	LUT3 #(
		.INIT('h80)
	) name3463 (
		\wishbone_bd_ram_mem0_reg[255][1]/P0001 ,
		_w11952_,
		_w11973_,
		_w13976_
	);
	LUT3 #(
		.INIT('h80)
	) name3464 (
		\wishbone_bd_ram_mem0_reg[89][1]/P0001 ,
		_w11968_,
		_w11972_,
		_w13977_
	);
	LUT4 #(
		.INIT('h0001)
	) name3465 (
		_w13974_,
		_w13975_,
		_w13976_,
		_w13977_,
		_w13978_
	);
	LUT4 #(
		.INIT('h8000)
	) name3466 (
		_w13963_,
		_w13968_,
		_w13973_,
		_w13978_,
		_w13979_
	);
	LUT4 #(
		.INIT('h8000)
	) name3467 (
		_w13916_,
		_w13937_,
		_w13958_,
		_w13979_,
		_w13980_
	);
	LUT3 #(
		.INIT('h80)
	) name3468 (
		\wishbone_bd_ram_mem0_reg[224][1]/P0001 ,
		_w11941_,
		_w11982_,
		_w13981_
	);
	LUT3 #(
		.INIT('h80)
	) name3469 (
		\wishbone_bd_ram_mem0_reg[30][1]/P0001 ,
		_w11935_,
		_w11948_,
		_w13982_
	);
	LUT3 #(
		.INIT('h80)
	) name3470 (
		\wishbone_bd_ram_mem0_reg[237][1]/P0001 ,
		_w11966_,
		_w11982_,
		_w13983_
	);
	LUT3 #(
		.INIT('h80)
	) name3471 (
		\wishbone_bd_ram_mem0_reg[234][1]/P0001 ,
		_w11944_,
		_w11982_,
		_w13984_
	);
	LUT4 #(
		.INIT('h0001)
	) name3472 (
		_w13981_,
		_w13982_,
		_w13983_,
		_w13984_,
		_w13985_
	);
	LUT3 #(
		.INIT('h80)
	) name3473 (
		\wishbone_bd_ram_mem0_reg[180][1]/P0001 ,
		_w11929_,
		_w11942_,
		_w13986_
	);
	LUT3 #(
		.INIT('h80)
	) name3474 (
		\wishbone_bd_ram_mem0_reg[120][1]/P0001 ,
		_w11990_,
		_w12012_,
		_w13987_
	);
	LUT3 #(
		.INIT('h80)
	) name3475 (
		\wishbone_bd_ram_mem0_reg[221][1]/P0001 ,
		_w11966_,
		_w11984_,
		_w13988_
	);
	LUT3 #(
		.INIT('h80)
	) name3476 (
		\wishbone_bd_ram_mem0_reg[202][1]/P0001 ,
		_w11944_,
		_w11945_,
		_w13989_
	);
	LUT4 #(
		.INIT('h0001)
	) name3477 (
		_w13986_,
		_w13987_,
		_w13988_,
		_w13989_,
		_w13990_
	);
	LUT3 #(
		.INIT('h80)
	) name3478 (
		\wishbone_bd_ram_mem0_reg[49][1]/P0001 ,
		_w11977_,
		_w11979_,
		_w13991_
	);
	LUT3 #(
		.INIT('h80)
	) name3479 (
		\wishbone_bd_ram_mem0_reg[153][1]/P0001 ,
		_w11959_,
		_w11968_,
		_w13992_
	);
	LUT3 #(
		.INIT('h80)
	) name3480 (
		\wishbone_bd_ram_mem0_reg[77][1]/P0001 ,
		_w11949_,
		_w11966_,
		_w13993_
	);
	LUT3 #(
		.INIT('h80)
	) name3481 (
		\wishbone_bd_ram_mem0_reg[172][1]/P0001 ,
		_w11930_,
		_w11954_,
		_w13994_
	);
	LUT4 #(
		.INIT('h0001)
	) name3482 (
		_w13991_,
		_w13992_,
		_w13993_,
		_w13994_,
		_w13995_
	);
	LUT3 #(
		.INIT('h80)
	) name3483 (
		\wishbone_bd_ram_mem0_reg[86][1]/P0001 ,
		_w11972_,
		_w11986_,
		_w13996_
	);
	LUT3 #(
		.INIT('h80)
	) name3484 (
		\wishbone_bd_ram_mem0_reg[118][1]/P0001 ,
		_w11986_,
		_w12012_,
		_w13997_
	);
	LUT3 #(
		.INIT('h80)
	) name3485 (
		\wishbone_bd_ram_mem0_reg[99][1]/P0001 ,
		_w11938_,
		_w11965_,
		_w13998_
	);
	LUT3 #(
		.INIT('h80)
	) name3486 (
		\wishbone_bd_ram_mem0_reg[206][1]/P0001 ,
		_w11945_,
		_w11948_,
		_w13999_
	);
	LUT4 #(
		.INIT('h0001)
	) name3487 (
		_w13996_,
		_w13997_,
		_w13998_,
		_w13999_,
		_w14000_
	);
	LUT4 #(
		.INIT('h8000)
	) name3488 (
		_w13985_,
		_w13990_,
		_w13995_,
		_w14000_,
		_w14001_
	);
	LUT3 #(
		.INIT('h80)
	) name3489 (
		\wishbone_bd_ram_mem0_reg[176][1]/P0001 ,
		_w11941_,
		_w11942_,
		_w14002_
	);
	LUT3 #(
		.INIT('h80)
	) name3490 (
		\wishbone_bd_ram_mem0_reg[204][1]/P0001 ,
		_w11945_,
		_w11954_,
		_w14003_
	);
	LUT3 #(
		.INIT('h80)
	) name3491 (
		\wishbone_bd_ram_mem0_reg[211][1]/P0001 ,
		_w11938_,
		_w11984_,
		_w14004_
	);
	LUT3 #(
		.INIT('h80)
	) name3492 (
		\wishbone_bd_ram_mem0_reg[121][1]/P0001 ,
		_w11968_,
		_w12012_,
		_w14005_
	);
	LUT4 #(
		.INIT('h0001)
	) name3493 (
		_w14002_,
		_w14003_,
		_w14004_,
		_w14005_,
		_w14006_
	);
	LUT3 #(
		.INIT('h80)
	) name3494 (
		\wishbone_bd_ram_mem0_reg[81][1]/P0001 ,
		_w11972_,
		_w11977_,
		_w14007_
	);
	LUT3 #(
		.INIT('h80)
	) name3495 (
		\wishbone_bd_ram_mem0_reg[132][1]/P0001 ,
		_w11929_,
		_w11955_,
		_w14008_
	);
	LUT3 #(
		.INIT('h80)
	) name3496 (
		\wishbone_bd_ram_mem0_reg[66][1]/P0001 ,
		_w11949_,
		_w11963_,
		_w14009_
	);
	LUT3 #(
		.INIT('h80)
	) name3497 (
		\wishbone_bd_ram_mem0_reg[70][1]/P0001 ,
		_w11949_,
		_w11986_,
		_w14010_
	);
	LUT4 #(
		.INIT('h0001)
	) name3498 (
		_w14007_,
		_w14008_,
		_w14009_,
		_w14010_,
		_w14011_
	);
	LUT3 #(
		.INIT('h80)
	) name3499 (
		\wishbone_bd_ram_mem0_reg[80][1]/P0001 ,
		_w11941_,
		_w11972_,
		_w14012_
	);
	LUT3 #(
		.INIT('h80)
	) name3500 (
		\wishbone_bd_ram_mem0_reg[144][1]/P0001 ,
		_w11941_,
		_w11959_,
		_w14013_
	);
	LUT3 #(
		.INIT('h80)
	) name3501 (
		\wishbone_bd_ram_mem0_reg[112][1]/P0001 ,
		_w11941_,
		_w12012_,
		_w14014_
	);
	LUT3 #(
		.INIT('h80)
	) name3502 (
		\wishbone_bd_ram_mem0_reg[10][1]/P0001 ,
		_w11932_,
		_w11944_,
		_w14015_
	);
	LUT4 #(
		.INIT('h0001)
	) name3503 (
		_w14012_,
		_w14013_,
		_w14014_,
		_w14015_,
		_w14016_
	);
	LUT3 #(
		.INIT('h80)
	) name3504 (
		\wishbone_bd_ram_mem0_reg[25][1]/P0001 ,
		_w11935_,
		_w11968_,
		_w14017_
	);
	LUT3 #(
		.INIT('h80)
	) name3505 (
		\wishbone_bd_ram_mem0_reg[207][1]/P0001 ,
		_w11945_,
		_w11973_,
		_w14018_
	);
	LUT3 #(
		.INIT('h80)
	) name3506 (
		\wishbone_bd_ram_mem0_reg[233][1]/P0001 ,
		_w11968_,
		_w11982_,
		_w14019_
	);
	LUT3 #(
		.INIT('h80)
	) name3507 (
		\wishbone_bd_ram_mem0_reg[194][1]/P0001 ,
		_w11945_,
		_w11963_,
		_w14020_
	);
	LUT4 #(
		.INIT('h0001)
	) name3508 (
		_w14017_,
		_w14018_,
		_w14019_,
		_w14020_,
		_w14021_
	);
	LUT4 #(
		.INIT('h8000)
	) name3509 (
		_w14006_,
		_w14011_,
		_w14016_,
		_w14021_,
		_w14022_
	);
	LUT3 #(
		.INIT('h80)
	) name3510 (
		\wishbone_bd_ram_mem0_reg[240][1]/P0001 ,
		_w11941_,
		_w11952_,
		_w14023_
	);
	LUT3 #(
		.INIT('h80)
	) name3511 (
		\wishbone_bd_ram_mem0_reg[32][1]/P0001 ,
		_w11941_,
		_w11957_,
		_w14024_
	);
	LUT3 #(
		.INIT('h80)
	) name3512 (
		\wishbone_bd_ram_mem0_reg[106][1]/P0001 ,
		_w11944_,
		_w11965_,
		_w14025_
	);
	LUT3 #(
		.INIT('h80)
	) name3513 (
		\wishbone_bd_ram_mem0_reg[185][1]/P0001 ,
		_w11942_,
		_w11968_,
		_w14026_
	);
	LUT4 #(
		.INIT('h0001)
	) name3514 (
		_w14023_,
		_w14024_,
		_w14025_,
		_w14026_,
		_w14027_
	);
	LUT3 #(
		.INIT('h80)
	) name3515 (
		\wishbone_bd_ram_mem0_reg[92][1]/P0001 ,
		_w11954_,
		_w11972_,
		_w14028_
	);
	LUT3 #(
		.INIT('h80)
	) name3516 (
		\wishbone_bd_ram_mem0_reg[37][1]/P0001 ,
		_w11933_,
		_w11957_,
		_w14029_
	);
	LUT3 #(
		.INIT('h80)
	) name3517 (
		\wishbone_bd_ram_mem0_reg[82][1]/P0001 ,
		_w11963_,
		_w11972_,
		_w14030_
	);
	LUT3 #(
		.INIT('h80)
	) name3518 (
		\wishbone_bd_ram_mem0_reg[117][1]/P0001 ,
		_w11933_,
		_w12012_,
		_w14031_
	);
	LUT4 #(
		.INIT('h0001)
	) name3519 (
		_w14028_,
		_w14029_,
		_w14030_,
		_w14031_,
		_w14032_
	);
	LUT3 #(
		.INIT('h80)
	) name3520 (
		\wishbone_bd_ram_mem0_reg[173][1]/P0001 ,
		_w11930_,
		_w11966_,
		_w14033_
	);
	LUT3 #(
		.INIT('h80)
	) name3521 (
		\wishbone_bd_ram_mem0_reg[136][1]/P0001 ,
		_w11955_,
		_w11990_,
		_w14034_
	);
	LUT3 #(
		.INIT('h80)
	) name3522 (
		\wishbone_bd_ram_mem0_reg[9][1]/P0001 ,
		_w11932_,
		_w11968_,
		_w14035_
	);
	LUT3 #(
		.INIT('h80)
	) name3523 (
		\wishbone_bd_ram_mem0_reg[131][1]/P0001 ,
		_w11938_,
		_w11955_,
		_w14036_
	);
	LUT4 #(
		.INIT('h0001)
	) name3524 (
		_w14033_,
		_w14034_,
		_w14035_,
		_w14036_,
		_w14037_
	);
	LUT3 #(
		.INIT('h80)
	) name3525 (
		\wishbone_bd_ram_mem0_reg[20][1]/P0001 ,
		_w11929_,
		_w11935_,
		_w14038_
	);
	LUT3 #(
		.INIT('h80)
	) name3526 (
		\wishbone_bd_ram_mem0_reg[36][1]/P0001 ,
		_w11929_,
		_w11957_,
		_w14039_
	);
	LUT3 #(
		.INIT('h80)
	) name3527 (
		\wishbone_bd_ram_mem0_reg[28][1]/P0001 ,
		_w11935_,
		_w11954_,
		_w14040_
	);
	LUT3 #(
		.INIT('h80)
	) name3528 (
		\wishbone_bd_ram_mem0_reg[101][1]/P0001 ,
		_w11933_,
		_w11965_,
		_w14041_
	);
	LUT4 #(
		.INIT('h0001)
	) name3529 (
		_w14038_,
		_w14039_,
		_w14040_,
		_w14041_,
		_w14042_
	);
	LUT4 #(
		.INIT('h8000)
	) name3530 (
		_w14027_,
		_w14032_,
		_w14037_,
		_w14042_,
		_w14043_
	);
	LUT3 #(
		.INIT('h80)
	) name3531 (
		\wishbone_bd_ram_mem0_reg[192][1]/P0001 ,
		_w11941_,
		_w11945_,
		_w14044_
	);
	LUT3 #(
		.INIT('h80)
	) name3532 (
		\wishbone_bd_ram_mem0_reg[0][1]/P0001 ,
		_w11932_,
		_w11941_,
		_w14045_
	);
	LUT3 #(
		.INIT('h80)
	) name3533 (
		\wishbone_bd_ram_mem0_reg[195][1]/P0001 ,
		_w11938_,
		_w11945_,
		_w14046_
	);
	LUT3 #(
		.INIT('h80)
	) name3534 (
		\wishbone_bd_ram_mem0_reg[178][1]/P0001 ,
		_w11942_,
		_w11963_,
		_w14047_
	);
	LUT4 #(
		.INIT('h0001)
	) name3535 (
		_w14044_,
		_w14045_,
		_w14046_,
		_w14047_,
		_w14048_
	);
	LUT3 #(
		.INIT('h80)
	) name3536 (
		\wishbone_bd_ram_mem0_reg[98][1]/P0001 ,
		_w11963_,
		_w11965_,
		_w14049_
	);
	LUT3 #(
		.INIT('h80)
	) name3537 (
		\wishbone_bd_ram_mem0_reg[203][1]/P0001 ,
		_w11936_,
		_w11945_,
		_w14050_
	);
	LUT3 #(
		.INIT('h80)
	) name3538 (
		\wishbone_bd_ram_mem0_reg[253][1]/P0001 ,
		_w11952_,
		_w11966_,
		_w14051_
	);
	LUT3 #(
		.INIT('h80)
	) name3539 (
		\wishbone_bd_ram_mem0_reg[156][1]/P0001 ,
		_w11954_,
		_w11959_,
		_w14052_
	);
	LUT4 #(
		.INIT('h0001)
	) name3540 (
		_w14049_,
		_w14050_,
		_w14051_,
		_w14052_,
		_w14053_
	);
	LUT3 #(
		.INIT('h80)
	) name3541 (
		\wishbone_bd_ram_mem0_reg[15][1]/P0001 ,
		_w11932_,
		_w11973_,
		_w14054_
	);
	LUT3 #(
		.INIT('h80)
	) name3542 (
		\wishbone_bd_ram_mem0_reg[39][1]/P0001 ,
		_w11957_,
		_w11975_,
		_w14055_
	);
	LUT3 #(
		.INIT('h80)
	) name3543 (
		\wishbone_bd_ram_mem0_reg[186][1]/P0001 ,
		_w11942_,
		_w11944_,
		_w14056_
	);
	LUT3 #(
		.INIT('h80)
	) name3544 (
		\wishbone_bd_ram_mem0_reg[138][1]/P0001 ,
		_w11944_,
		_w11955_,
		_w14057_
	);
	LUT4 #(
		.INIT('h0001)
	) name3545 (
		_w14054_,
		_w14055_,
		_w14056_,
		_w14057_,
		_w14058_
	);
	LUT3 #(
		.INIT('h80)
	) name3546 (
		\wishbone_bd_ram_mem0_reg[246][1]/P0001 ,
		_w11952_,
		_w11986_,
		_w14059_
	);
	LUT3 #(
		.INIT('h80)
	) name3547 (
		\wishbone_bd_ram_mem0_reg[179][1]/P0001 ,
		_w11938_,
		_w11942_,
		_w14060_
	);
	LUT3 #(
		.INIT('h80)
	) name3548 (
		\wishbone_bd_ram_mem0_reg[189][1]/P0001 ,
		_w11942_,
		_w11966_,
		_w14061_
	);
	LUT3 #(
		.INIT('h80)
	) name3549 (
		\wishbone_bd_ram_mem0_reg[183][1]/P0001 ,
		_w11942_,
		_w11975_,
		_w14062_
	);
	LUT4 #(
		.INIT('h0001)
	) name3550 (
		_w14059_,
		_w14060_,
		_w14061_,
		_w14062_,
		_w14063_
	);
	LUT4 #(
		.INIT('h8000)
	) name3551 (
		_w14048_,
		_w14053_,
		_w14058_,
		_w14063_,
		_w14064_
	);
	LUT4 #(
		.INIT('h8000)
	) name3552 (
		_w14001_,
		_w14022_,
		_w14043_,
		_w14064_,
		_w14065_
	);
	LUT3 #(
		.INIT('h80)
	) name3553 (
		\wishbone_bd_ram_mem0_reg[102][1]/P0001 ,
		_w11965_,
		_w11986_,
		_w14066_
	);
	LUT3 #(
		.INIT('h80)
	) name3554 (
		\wishbone_bd_ram_mem0_reg[134][1]/P0001 ,
		_w11955_,
		_w11986_,
		_w14067_
	);
	LUT3 #(
		.INIT('h80)
	) name3555 (
		\wishbone_bd_ram_mem0_reg[93][1]/P0001 ,
		_w11966_,
		_w11972_,
		_w14068_
	);
	LUT3 #(
		.INIT('h80)
	) name3556 (
		\wishbone_bd_ram_mem0_reg[162][1]/P0001 ,
		_w11930_,
		_w11963_,
		_w14069_
	);
	LUT4 #(
		.INIT('h0001)
	) name3557 (
		_w14066_,
		_w14067_,
		_w14068_,
		_w14069_,
		_w14070_
	);
	LUT3 #(
		.INIT('h80)
	) name3558 (
		\wishbone_bd_ram_mem0_reg[61][1]/P0001 ,
		_w11966_,
		_w11979_,
		_w14071_
	);
	LUT3 #(
		.INIT('h80)
	) name3559 (
		\wishbone_bd_ram_mem0_reg[158][1]/P0001 ,
		_w11948_,
		_w11959_,
		_w14072_
	);
	LUT3 #(
		.INIT('h80)
	) name3560 (
		\wishbone_bd_ram_mem0_reg[148][1]/P0001 ,
		_w11929_,
		_w11959_,
		_w14073_
	);
	LUT3 #(
		.INIT('h80)
	) name3561 (
		\wishbone_bd_ram_mem0_reg[142][1]/P0001 ,
		_w11948_,
		_w11955_,
		_w14074_
	);
	LUT4 #(
		.INIT('h0001)
	) name3562 (
		_w14071_,
		_w14072_,
		_w14073_,
		_w14074_,
		_w14075_
	);
	LUT3 #(
		.INIT('h80)
	) name3563 (
		\wishbone_bd_ram_mem0_reg[48][1]/P0001 ,
		_w11941_,
		_w11979_,
		_w14076_
	);
	LUT3 #(
		.INIT('h80)
	) name3564 (
		\wishbone_bd_ram_mem0_reg[232][1]/P0001 ,
		_w11982_,
		_w11990_,
		_w14077_
	);
	LUT3 #(
		.INIT('h80)
	) name3565 (
		\wishbone_bd_ram_mem0_reg[154][1]/P0001 ,
		_w11944_,
		_w11959_,
		_w14078_
	);
	LUT3 #(
		.INIT('h80)
	) name3566 (
		\wishbone_bd_ram_mem0_reg[113][1]/P0001 ,
		_w11977_,
		_w12012_,
		_w14079_
	);
	LUT4 #(
		.INIT('h0001)
	) name3567 (
		_w14076_,
		_w14077_,
		_w14078_,
		_w14079_,
		_w14080_
	);
	LUT3 #(
		.INIT('h80)
	) name3568 (
		\wishbone_bd_ram_mem0_reg[188][1]/P0001 ,
		_w11942_,
		_w11954_,
		_w14081_
	);
	LUT3 #(
		.INIT('h80)
	) name3569 (
		\wishbone_bd_ram_mem0_reg[223][1]/P0001 ,
		_w11973_,
		_w11984_,
		_w14082_
	);
	LUT3 #(
		.INIT('h80)
	) name3570 (
		\wishbone_bd_ram_mem0_reg[227][1]/P0001 ,
		_w11938_,
		_w11982_,
		_w14083_
	);
	LUT3 #(
		.INIT('h80)
	) name3571 (
		\wishbone_bd_ram_mem0_reg[24][1]/P0001 ,
		_w11935_,
		_w11990_,
		_w14084_
	);
	LUT4 #(
		.INIT('h0001)
	) name3572 (
		_w14081_,
		_w14082_,
		_w14083_,
		_w14084_,
		_w14085_
	);
	LUT4 #(
		.INIT('h8000)
	) name3573 (
		_w14070_,
		_w14075_,
		_w14080_,
		_w14085_,
		_w14086_
	);
	LUT3 #(
		.INIT('h80)
	) name3574 (
		\wishbone_bd_ram_mem0_reg[191][1]/P0001 ,
		_w11942_,
		_w11973_,
		_w14087_
	);
	LUT3 #(
		.INIT('h80)
	) name3575 (
		\wishbone_bd_ram_mem0_reg[139][1]/P0001 ,
		_w11936_,
		_w11955_,
		_w14088_
	);
	LUT3 #(
		.INIT('h80)
	) name3576 (
		\wishbone_bd_ram_mem0_reg[182][1]/P0001 ,
		_w11942_,
		_w11986_,
		_w14089_
	);
	LUT3 #(
		.INIT('h80)
	) name3577 (
		\wishbone_bd_ram_mem0_reg[119][1]/P0001 ,
		_w11975_,
		_w12012_,
		_w14090_
	);
	LUT4 #(
		.INIT('h0001)
	) name3578 (
		_w14087_,
		_w14088_,
		_w14089_,
		_w14090_,
		_w14091_
	);
	LUT3 #(
		.INIT('h80)
	) name3579 (
		\wishbone_bd_ram_mem0_reg[29][1]/P0001 ,
		_w11935_,
		_w11966_,
		_w14092_
	);
	LUT3 #(
		.INIT('h80)
	) name3580 (
		\wishbone_bd_ram_mem0_reg[152][1]/P0001 ,
		_w11959_,
		_w11990_,
		_w14093_
	);
	LUT3 #(
		.INIT('h80)
	) name3581 (
		\wishbone_bd_ram_mem0_reg[239][1]/P0001 ,
		_w11973_,
		_w11982_,
		_w14094_
	);
	LUT3 #(
		.INIT('h80)
	) name3582 (
		\wishbone_bd_ram_mem0_reg[219][1]/P0001 ,
		_w11936_,
		_w11984_,
		_w14095_
	);
	LUT4 #(
		.INIT('h0001)
	) name3583 (
		_w14092_,
		_w14093_,
		_w14094_,
		_w14095_,
		_w14096_
	);
	LUT3 #(
		.INIT('h80)
	) name3584 (
		\wishbone_bd_ram_mem0_reg[243][1]/P0001 ,
		_w11938_,
		_w11952_,
		_w14097_
	);
	LUT3 #(
		.INIT('h80)
	) name3585 (
		\wishbone_bd_ram_mem0_reg[150][1]/P0001 ,
		_w11959_,
		_w11986_,
		_w14098_
	);
	LUT3 #(
		.INIT('h80)
	) name3586 (
		\wishbone_bd_ram_mem0_reg[251][1]/P0001 ,
		_w11936_,
		_w11952_,
		_w14099_
	);
	LUT3 #(
		.INIT('h80)
	) name3587 (
		\wishbone_bd_ram_mem0_reg[43][1]/P0001 ,
		_w11936_,
		_w11957_,
		_w14100_
	);
	LUT4 #(
		.INIT('h0001)
	) name3588 (
		_w14097_,
		_w14098_,
		_w14099_,
		_w14100_,
		_w14101_
	);
	LUT3 #(
		.INIT('h80)
	) name3589 (
		\wishbone_bd_ram_mem0_reg[103][1]/P0001 ,
		_w11965_,
		_w11975_,
		_w14102_
	);
	LUT3 #(
		.INIT('h80)
	) name3590 (
		\wishbone_bd_ram_mem0_reg[96][1]/P0001 ,
		_w11941_,
		_w11965_,
		_w14103_
	);
	LUT3 #(
		.INIT('h80)
	) name3591 (
		\wishbone_bd_ram_mem0_reg[83][1]/P0001 ,
		_w11938_,
		_w11972_,
		_w14104_
	);
	LUT3 #(
		.INIT('h80)
	) name3592 (
		\wishbone_bd_ram_mem0_reg[133][1]/P0001 ,
		_w11933_,
		_w11955_,
		_w14105_
	);
	LUT4 #(
		.INIT('h0001)
	) name3593 (
		_w14102_,
		_w14103_,
		_w14104_,
		_w14105_,
		_w14106_
	);
	LUT4 #(
		.INIT('h8000)
	) name3594 (
		_w14091_,
		_w14096_,
		_w14101_,
		_w14106_,
		_w14107_
	);
	LUT3 #(
		.INIT('h80)
	) name3595 (
		\wishbone_bd_ram_mem0_reg[64][1]/P0001 ,
		_w11941_,
		_w11949_,
		_w14108_
	);
	LUT3 #(
		.INIT('h80)
	) name3596 (
		\wishbone_bd_ram_mem0_reg[209][1]/P0001 ,
		_w11977_,
		_w11984_,
		_w14109_
	);
	LUT3 #(
		.INIT('h80)
	) name3597 (
		\wishbone_bd_ram_mem0_reg[78][1]/P0001 ,
		_w11948_,
		_w11949_,
		_w14110_
	);
	LUT3 #(
		.INIT('h80)
	) name3598 (
		\wishbone_bd_ram_mem0_reg[116][1]/P0001 ,
		_w11929_,
		_w12012_,
		_w14111_
	);
	LUT4 #(
		.INIT('h0001)
	) name3599 (
		_w14108_,
		_w14109_,
		_w14110_,
		_w14111_,
		_w14112_
	);
	LUT3 #(
		.INIT('h80)
	) name3600 (
		\wishbone_bd_ram_mem0_reg[56][1]/P0001 ,
		_w11979_,
		_w11990_,
		_w14113_
	);
	LUT3 #(
		.INIT('h80)
	) name3601 (
		\wishbone_bd_ram_mem0_reg[147][1]/P0001 ,
		_w11938_,
		_w11959_,
		_w14114_
	);
	LUT3 #(
		.INIT('h80)
	) name3602 (
		\wishbone_bd_ram_mem0_reg[210][1]/P0001 ,
		_w11963_,
		_w11984_,
		_w14115_
	);
	LUT3 #(
		.INIT('h80)
	) name3603 (
		\wishbone_bd_ram_mem0_reg[157][1]/P0001 ,
		_w11959_,
		_w11966_,
		_w14116_
	);
	LUT4 #(
		.INIT('h0001)
	) name3604 (
		_w14113_,
		_w14114_,
		_w14115_,
		_w14116_,
		_w14117_
	);
	LUT3 #(
		.INIT('h80)
	) name3605 (
		\wishbone_bd_ram_mem0_reg[4][1]/P0001 ,
		_w11929_,
		_w11932_,
		_w14118_
	);
	LUT3 #(
		.INIT('h80)
	) name3606 (
		\wishbone_bd_ram_mem0_reg[6][1]/P0001 ,
		_w11932_,
		_w11986_,
		_w14119_
	);
	LUT3 #(
		.INIT('h80)
	) name3607 (
		\wishbone_bd_ram_mem0_reg[26][1]/P0001 ,
		_w11935_,
		_w11944_,
		_w14120_
	);
	LUT3 #(
		.INIT('h80)
	) name3608 (
		\wishbone_bd_ram_mem0_reg[74][1]/P0001 ,
		_w11944_,
		_w11949_,
		_w14121_
	);
	LUT4 #(
		.INIT('h0001)
	) name3609 (
		_w14118_,
		_w14119_,
		_w14120_,
		_w14121_,
		_w14122_
	);
	LUT3 #(
		.INIT('h80)
	) name3610 (
		\wishbone_bd_ram_mem0_reg[71][1]/P0001 ,
		_w11949_,
		_w11975_,
		_w14123_
	);
	LUT3 #(
		.INIT('h80)
	) name3611 (
		\wishbone_bd_ram_mem0_reg[235][1]/P0001 ,
		_w11936_,
		_w11982_,
		_w14124_
	);
	LUT3 #(
		.INIT('h80)
	) name3612 (
		\wishbone_bd_ram_mem0_reg[228][1]/P0001 ,
		_w11929_,
		_w11982_,
		_w14125_
	);
	LUT3 #(
		.INIT('h80)
	) name3613 (
		\wishbone_bd_ram_mem0_reg[128][1]/P0001 ,
		_w11941_,
		_w11955_,
		_w14126_
	);
	LUT4 #(
		.INIT('h0001)
	) name3614 (
		_w14123_,
		_w14124_,
		_w14125_,
		_w14126_,
		_w14127_
	);
	LUT4 #(
		.INIT('h8000)
	) name3615 (
		_w14112_,
		_w14117_,
		_w14122_,
		_w14127_,
		_w14128_
	);
	LUT3 #(
		.INIT('h80)
	) name3616 (
		\wishbone_bd_ram_mem0_reg[212][1]/P0001 ,
		_w11929_,
		_w11984_,
		_w14129_
	);
	LUT3 #(
		.INIT('h80)
	) name3617 (
		\wishbone_bd_ram_mem0_reg[208][1]/P0001 ,
		_w11941_,
		_w11984_,
		_w14130_
	);
	LUT3 #(
		.INIT('h80)
	) name3618 (
		\wishbone_bd_ram_mem0_reg[68][1]/P0001 ,
		_w11929_,
		_w11949_,
		_w14131_
	);
	LUT3 #(
		.INIT('h80)
	) name3619 (
		\wishbone_bd_ram_mem0_reg[67][1]/P0001 ,
		_w11938_,
		_w11949_,
		_w14132_
	);
	LUT4 #(
		.INIT('h0001)
	) name3620 (
		_w14129_,
		_w14130_,
		_w14131_,
		_w14132_,
		_w14133_
	);
	LUT3 #(
		.INIT('h80)
	) name3621 (
		\wishbone_bd_ram_mem0_reg[165][1]/P0001 ,
		_w11930_,
		_w11933_,
		_w14134_
	);
	LUT3 #(
		.INIT('h80)
	) name3622 (
		\wishbone_bd_ram_mem0_reg[164][1]/P0001 ,
		_w11929_,
		_w11930_,
		_w14135_
	);
	LUT3 #(
		.INIT('h80)
	) name3623 (
		\wishbone_bd_ram_mem0_reg[76][1]/P0001 ,
		_w11949_,
		_w11954_,
		_w14136_
	);
	LUT3 #(
		.INIT('h80)
	) name3624 (
		\wishbone_bd_ram_mem0_reg[8][1]/P0001 ,
		_w11932_,
		_w11990_,
		_w14137_
	);
	LUT4 #(
		.INIT('h0001)
	) name3625 (
		_w14134_,
		_w14135_,
		_w14136_,
		_w14137_,
		_w14138_
	);
	LUT3 #(
		.INIT('h80)
	) name3626 (
		\wishbone_bd_ram_mem0_reg[110][1]/P0001 ,
		_w11948_,
		_w11965_,
		_w14139_
	);
	LUT3 #(
		.INIT('h80)
	) name3627 (
		\wishbone_bd_ram_mem0_reg[23][1]/P0001 ,
		_w11935_,
		_w11975_,
		_w14140_
	);
	LUT3 #(
		.INIT('h80)
	) name3628 (
		\wishbone_bd_ram_mem0_reg[97][1]/P0001 ,
		_w11965_,
		_w11977_,
		_w14141_
	);
	LUT3 #(
		.INIT('h80)
	) name3629 (
		\wishbone_bd_ram_mem0_reg[254][1]/P0001 ,
		_w11948_,
		_w11952_,
		_w14142_
	);
	LUT4 #(
		.INIT('h0001)
	) name3630 (
		_w14139_,
		_w14140_,
		_w14141_,
		_w14142_,
		_w14143_
	);
	LUT3 #(
		.INIT('h80)
	) name3631 (
		\wishbone_bd_ram_mem0_reg[169][1]/P0001 ,
		_w11930_,
		_w11968_,
		_w14144_
	);
	LUT3 #(
		.INIT('h80)
	) name3632 (
		\wishbone_bd_ram_mem0_reg[41][1]/P0001 ,
		_w11957_,
		_w11968_,
		_w14145_
	);
	LUT3 #(
		.INIT('h80)
	) name3633 (
		\wishbone_bd_ram_mem0_reg[236][1]/P0001 ,
		_w11954_,
		_w11982_,
		_w14146_
	);
	LUT3 #(
		.INIT('h80)
	) name3634 (
		\wishbone_bd_ram_mem0_reg[65][1]/P0001 ,
		_w11949_,
		_w11977_,
		_w14147_
	);
	LUT4 #(
		.INIT('h0001)
	) name3635 (
		_w14144_,
		_w14145_,
		_w14146_,
		_w14147_,
		_w14148_
	);
	LUT4 #(
		.INIT('h8000)
	) name3636 (
		_w14133_,
		_w14138_,
		_w14143_,
		_w14148_,
		_w14149_
	);
	LUT4 #(
		.INIT('h8000)
	) name3637 (
		_w14086_,
		_w14107_,
		_w14128_,
		_w14149_,
		_w14150_
	);
	LUT4 #(
		.INIT('h8000)
	) name3638 (
		_w13895_,
		_w13980_,
		_w14065_,
		_w14150_,
		_w14151_
	);
	LUT3 #(
		.INIT('h01)
	) name3639 (
		wb_rst_i_pad,
		_w13808_,
		_w13809_,
		_w14152_
	);
	LUT3 #(
		.INIT('hba)
	) name3640 (
		_w13810_,
		_w14151_,
		_w14152_,
		_w14153_
	);
	LUT3 #(
		.INIT('h14)
	) name3641 (
		\rxethmac1_crcrx_Crc_reg[21]/NET0131 ,
		_w10590_,
		_w11047_,
		_w14154_
	);
	LUT4 #(
		.INIT('h7000)
	) name3642 (
		_w10554_,
		_w10573_,
		_w10577_,
		_w14154_,
		_w14155_
	);
	LUT2 #(
		.INIT('h4)
	) name3643 (
		\rxethmac1_crcrx_Crc_reg[21]/NET0131 ,
		_w10582_,
		_w14156_
	);
	LUT3 #(
		.INIT('hcd)
	) name3644 (
		_w11447_,
		_w14155_,
		_w14156_,
		_w14157_
	);
	LUT4 #(
		.INIT('h1000)
	) name3645 (
		\txethmac1_txcrc_Crc_reg[4]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11787_,
		_w11790_,
		_w14158_
	);
	LUT3 #(
		.INIT('h40)
	) name3646 (
		\txethmac1_txcrc_Crc_reg[4]/NET0131 ,
		_w10913_,
		_w10914_,
		_w14159_
	);
	LUT3 #(
		.INIT('hcd)
	) name3647 (
		_w11793_,
		_w14158_,
		_w14159_,
		_w14160_
	);
	LUT2 #(
		.INIT('h8)
	) name3648 (
		\m_wb_adr_o[16]_pad ,
		\m_wb_adr_o[17]_pad ,
		_w14161_
	);
	LUT2 #(
		.INIT('h8)
	) name3649 (
		_w11851_,
		_w14161_,
		_w14162_
	);
	LUT3 #(
		.INIT('h15)
	) name3650 (
		\m_wb_adr_o[18]_pad ,
		_w11851_,
		_w14161_,
		_w14163_
	);
	LUT3 #(
		.INIT('h80)
	) name3651 (
		\m_wb_adr_o[16]_pad ,
		\m_wb_adr_o[17]_pad ,
		\m_wb_adr_o[18]_pad ,
		_w14164_
	);
	LUT2 #(
		.INIT('h8)
	) name3652 (
		_w11851_,
		_w14164_,
		_w14165_
	);
	LUT4 #(
		.INIT('h000e)
	) name3653 (
		_w11887_,
		_w13051_,
		_w14163_,
		_w14165_,
		_w14166_
	);
	LUT4 #(
		.INIT('h080a)
	) name3654 (
		\wishbone_RxPointerMSB_reg[18]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w14167_
	);
	LUT3 #(
		.INIT('he0)
	) name3655 (
		_w11902_,
		_w11905_,
		_w14167_,
		_w14168_
	);
	LUT3 #(
		.INIT('ha2)
	) name3656 (
		\wishbone_TxPointerMSB_reg[18]/NET0131 ,
		_w11900_,
		_w11909_,
		_w14169_
	);
	LUT4 #(
		.INIT('h0007)
	) name3657 (
		\m_wb_adr_o[18]_pad ,
		_w11907_,
		_w14168_,
		_w14169_,
		_w14170_
	);
	LUT2 #(
		.INIT('hb)
	) name3658 (
		_w14166_,
		_w14170_,
		_w14171_
	);
	LUT3 #(
		.INIT('h80)
	) name3659 (
		\wishbone_bd_ram_mem2_reg[67][20]/P0001 ,
		_w11938_,
		_w11949_,
		_w14172_
	);
	LUT3 #(
		.INIT('h80)
	) name3660 (
		\wishbone_bd_ram_mem2_reg[113][20]/P0001 ,
		_w11977_,
		_w12012_,
		_w14173_
	);
	LUT3 #(
		.INIT('h80)
	) name3661 (
		\wishbone_bd_ram_mem2_reg[140][20]/P0001 ,
		_w11954_,
		_w11955_,
		_w14174_
	);
	LUT3 #(
		.INIT('h80)
	) name3662 (
		\wishbone_bd_ram_mem2_reg[245][20]/P0001 ,
		_w11933_,
		_w11952_,
		_w14175_
	);
	LUT4 #(
		.INIT('h0001)
	) name3663 (
		_w14172_,
		_w14173_,
		_w14174_,
		_w14175_,
		_w14176_
	);
	LUT3 #(
		.INIT('h80)
	) name3664 (
		\wishbone_bd_ram_mem2_reg[99][20]/P0001 ,
		_w11938_,
		_w11965_,
		_w14177_
	);
	LUT3 #(
		.INIT('h80)
	) name3665 (
		\wishbone_bd_ram_mem2_reg[133][20]/P0001 ,
		_w11933_,
		_w11955_,
		_w14178_
	);
	LUT3 #(
		.INIT('h80)
	) name3666 (
		\wishbone_bd_ram_mem2_reg[43][20]/P0001 ,
		_w11936_,
		_w11957_,
		_w14179_
	);
	LUT3 #(
		.INIT('h80)
	) name3667 (
		\wishbone_bd_ram_mem2_reg[34][20]/P0001 ,
		_w11957_,
		_w11963_,
		_w14180_
	);
	LUT4 #(
		.INIT('h0001)
	) name3668 (
		_w14177_,
		_w14178_,
		_w14179_,
		_w14180_,
		_w14181_
	);
	LUT3 #(
		.INIT('h80)
	) name3669 (
		\wishbone_bd_ram_mem2_reg[252][20]/P0001 ,
		_w11952_,
		_w11954_,
		_w14182_
	);
	LUT3 #(
		.INIT('h80)
	) name3670 (
		\wishbone_bd_ram_mem2_reg[3][20]/P0001 ,
		_w11932_,
		_w11938_,
		_w14183_
	);
	LUT3 #(
		.INIT('h80)
	) name3671 (
		\wishbone_bd_ram_mem2_reg[180][20]/P0001 ,
		_w11929_,
		_w11942_,
		_w14184_
	);
	LUT3 #(
		.INIT('h80)
	) name3672 (
		\wishbone_bd_ram_mem2_reg[83][20]/P0001 ,
		_w11938_,
		_w11972_,
		_w14185_
	);
	LUT4 #(
		.INIT('h0001)
	) name3673 (
		_w14182_,
		_w14183_,
		_w14184_,
		_w14185_,
		_w14186_
	);
	LUT3 #(
		.INIT('h80)
	) name3674 (
		\wishbone_bd_ram_mem2_reg[87][20]/P0001 ,
		_w11972_,
		_w11975_,
		_w14187_
	);
	LUT3 #(
		.INIT('h80)
	) name3675 (
		\wishbone_bd_ram_mem2_reg[194][20]/P0001 ,
		_w11945_,
		_w11963_,
		_w14188_
	);
	LUT3 #(
		.INIT('h80)
	) name3676 (
		\wishbone_bd_ram_mem2_reg[32][20]/P0001 ,
		_w11941_,
		_w11957_,
		_w14189_
	);
	LUT3 #(
		.INIT('h80)
	) name3677 (
		\wishbone_bd_ram_mem2_reg[29][20]/P0001 ,
		_w11935_,
		_w11966_,
		_w14190_
	);
	LUT4 #(
		.INIT('h0001)
	) name3678 (
		_w14187_,
		_w14188_,
		_w14189_,
		_w14190_,
		_w14191_
	);
	LUT4 #(
		.INIT('h8000)
	) name3679 (
		_w14176_,
		_w14181_,
		_w14186_,
		_w14191_,
		_w14192_
	);
	LUT3 #(
		.INIT('h80)
	) name3680 (
		\wishbone_bd_ram_mem2_reg[9][20]/P0001 ,
		_w11932_,
		_w11968_,
		_w14193_
	);
	LUT3 #(
		.INIT('h80)
	) name3681 (
		\wishbone_bd_ram_mem2_reg[135][20]/P0001 ,
		_w11955_,
		_w11975_,
		_w14194_
	);
	LUT3 #(
		.INIT('h80)
	) name3682 (
		\wishbone_bd_ram_mem2_reg[0][20]/P0001 ,
		_w11932_,
		_w11941_,
		_w14195_
	);
	LUT3 #(
		.INIT('h80)
	) name3683 (
		\wishbone_bd_ram_mem2_reg[19][20]/P0001 ,
		_w11935_,
		_w11938_,
		_w14196_
	);
	LUT4 #(
		.INIT('h0001)
	) name3684 (
		_w14193_,
		_w14194_,
		_w14195_,
		_w14196_,
		_w14197_
	);
	LUT3 #(
		.INIT('h80)
	) name3685 (
		\wishbone_bd_ram_mem2_reg[53][20]/P0001 ,
		_w11933_,
		_w11979_,
		_w14198_
	);
	LUT3 #(
		.INIT('h80)
	) name3686 (
		\wishbone_bd_ram_mem2_reg[164][20]/P0001 ,
		_w11929_,
		_w11930_,
		_w14199_
	);
	LUT3 #(
		.INIT('h80)
	) name3687 (
		\wishbone_bd_ram_mem2_reg[215][20]/P0001 ,
		_w11975_,
		_w11984_,
		_w14200_
	);
	LUT3 #(
		.INIT('h80)
	) name3688 (
		\wishbone_bd_ram_mem2_reg[4][20]/P0001 ,
		_w11929_,
		_w11932_,
		_w14201_
	);
	LUT4 #(
		.INIT('h0001)
	) name3689 (
		_w14198_,
		_w14199_,
		_w14200_,
		_w14201_,
		_w14202_
	);
	LUT3 #(
		.INIT('h80)
	) name3690 (
		\wishbone_bd_ram_mem2_reg[65][20]/P0001 ,
		_w11949_,
		_w11977_,
		_w14203_
	);
	LUT3 #(
		.INIT('h80)
	) name3691 (
		\wishbone_bd_ram_mem2_reg[165][20]/P0001 ,
		_w11930_,
		_w11933_,
		_w14204_
	);
	LUT3 #(
		.INIT('h80)
	) name3692 (
		\wishbone_bd_ram_mem2_reg[134][20]/P0001 ,
		_w11955_,
		_w11986_,
		_w14205_
	);
	LUT3 #(
		.INIT('h80)
	) name3693 (
		\wishbone_bd_ram_mem2_reg[146][20]/P0001 ,
		_w11959_,
		_w11963_,
		_w14206_
	);
	LUT4 #(
		.INIT('h0001)
	) name3694 (
		_w14203_,
		_w14204_,
		_w14205_,
		_w14206_,
		_w14207_
	);
	LUT3 #(
		.INIT('h80)
	) name3695 (
		\wishbone_bd_ram_mem2_reg[211][20]/P0001 ,
		_w11938_,
		_w11984_,
		_w14208_
	);
	LUT3 #(
		.INIT('h80)
	) name3696 (
		\wishbone_bd_ram_mem2_reg[235][20]/P0001 ,
		_w11936_,
		_w11982_,
		_w14209_
	);
	LUT3 #(
		.INIT('h80)
	) name3697 (
		\wishbone_bd_ram_mem2_reg[119][20]/P0001 ,
		_w11975_,
		_w12012_,
		_w14210_
	);
	LUT3 #(
		.INIT('h80)
	) name3698 (
		\wishbone_bd_ram_mem2_reg[10][20]/P0001 ,
		_w11932_,
		_w11944_,
		_w14211_
	);
	LUT4 #(
		.INIT('h0001)
	) name3699 (
		_w14208_,
		_w14209_,
		_w14210_,
		_w14211_,
		_w14212_
	);
	LUT4 #(
		.INIT('h8000)
	) name3700 (
		_w14197_,
		_w14202_,
		_w14207_,
		_w14212_,
		_w14213_
	);
	LUT3 #(
		.INIT('h80)
	) name3701 (
		\wishbone_bd_ram_mem2_reg[40][20]/P0001 ,
		_w11957_,
		_w11990_,
		_w14214_
	);
	LUT3 #(
		.INIT('h80)
	) name3702 (
		\wishbone_bd_ram_mem2_reg[229][20]/P0001 ,
		_w11933_,
		_w11982_,
		_w14215_
	);
	LUT3 #(
		.INIT('h80)
	) name3703 (
		\wishbone_bd_ram_mem2_reg[73][20]/P0001 ,
		_w11949_,
		_w11968_,
		_w14216_
	);
	LUT3 #(
		.INIT('h80)
	) name3704 (
		\wishbone_bd_ram_mem2_reg[236][20]/P0001 ,
		_w11954_,
		_w11982_,
		_w14217_
	);
	LUT4 #(
		.INIT('h0001)
	) name3705 (
		_w14214_,
		_w14215_,
		_w14216_,
		_w14217_,
		_w14218_
	);
	LUT3 #(
		.INIT('h80)
	) name3706 (
		\wishbone_bd_ram_mem2_reg[157][20]/P0001 ,
		_w11959_,
		_w11966_,
		_w14219_
	);
	LUT3 #(
		.INIT('h80)
	) name3707 (
		\wishbone_bd_ram_mem2_reg[90][20]/P0001 ,
		_w11944_,
		_w11972_,
		_w14220_
	);
	LUT3 #(
		.INIT('h80)
	) name3708 (
		\wishbone_bd_ram_mem2_reg[45][20]/P0001 ,
		_w11957_,
		_w11966_,
		_w14221_
	);
	LUT3 #(
		.INIT('h80)
	) name3709 (
		\wishbone_bd_ram_mem2_reg[125][20]/P0001 ,
		_w11966_,
		_w12012_,
		_w14222_
	);
	LUT4 #(
		.INIT('h0001)
	) name3710 (
		_w14219_,
		_w14220_,
		_w14221_,
		_w14222_,
		_w14223_
	);
	LUT3 #(
		.INIT('h80)
	) name3711 (
		\wishbone_bd_ram_mem2_reg[244][20]/P0001 ,
		_w11929_,
		_w11952_,
		_w14224_
	);
	LUT3 #(
		.INIT('h80)
	) name3712 (
		\wishbone_bd_ram_mem2_reg[193][20]/P0001 ,
		_w11945_,
		_w11977_,
		_w14225_
	);
	LUT3 #(
		.INIT('h80)
	) name3713 (
		\wishbone_bd_ram_mem2_reg[172][20]/P0001 ,
		_w11930_,
		_w11954_,
		_w14226_
	);
	LUT3 #(
		.INIT('h80)
	) name3714 (
		\wishbone_bd_ram_mem2_reg[116][20]/P0001 ,
		_w11929_,
		_w12012_,
		_w14227_
	);
	LUT4 #(
		.INIT('h0001)
	) name3715 (
		_w14224_,
		_w14225_,
		_w14226_,
		_w14227_,
		_w14228_
	);
	LUT3 #(
		.INIT('h80)
	) name3716 (
		\wishbone_bd_ram_mem2_reg[222][20]/P0001 ,
		_w11948_,
		_w11984_,
		_w14229_
	);
	LUT3 #(
		.INIT('h80)
	) name3717 (
		\wishbone_bd_ram_mem2_reg[137][20]/P0001 ,
		_w11955_,
		_w11968_,
		_w14230_
	);
	LUT3 #(
		.INIT('h80)
	) name3718 (
		\wishbone_bd_ram_mem2_reg[126][20]/P0001 ,
		_w11948_,
		_w12012_,
		_w14231_
	);
	LUT3 #(
		.INIT('h80)
	) name3719 (
		\wishbone_bd_ram_mem2_reg[109][20]/P0001 ,
		_w11965_,
		_w11966_,
		_w14232_
	);
	LUT4 #(
		.INIT('h0001)
	) name3720 (
		_w14229_,
		_w14230_,
		_w14231_,
		_w14232_,
		_w14233_
	);
	LUT4 #(
		.INIT('h8000)
	) name3721 (
		_w14218_,
		_w14223_,
		_w14228_,
		_w14233_,
		_w14234_
	);
	LUT3 #(
		.INIT('h80)
	) name3722 (
		\wishbone_bd_ram_mem2_reg[158][20]/P0001 ,
		_w11948_,
		_w11959_,
		_w14235_
	);
	LUT3 #(
		.INIT('h80)
	) name3723 (
		\wishbone_bd_ram_mem2_reg[8][20]/P0001 ,
		_w11932_,
		_w11990_,
		_w14236_
	);
	LUT3 #(
		.INIT('h80)
	) name3724 (
		\wishbone_bd_ram_mem2_reg[89][20]/P0001 ,
		_w11968_,
		_w11972_,
		_w14237_
	);
	LUT3 #(
		.INIT('h80)
	) name3725 (
		\wishbone_bd_ram_mem2_reg[204][20]/P0001 ,
		_w11945_,
		_w11954_,
		_w14238_
	);
	LUT4 #(
		.INIT('h0001)
	) name3726 (
		_w14235_,
		_w14236_,
		_w14237_,
		_w14238_,
		_w14239_
	);
	LUT3 #(
		.INIT('h80)
	) name3727 (
		\wishbone_bd_ram_mem2_reg[41][20]/P0001 ,
		_w11957_,
		_w11968_,
		_w14240_
	);
	LUT3 #(
		.INIT('h80)
	) name3728 (
		\wishbone_bd_ram_mem2_reg[33][20]/P0001 ,
		_w11957_,
		_w11977_,
		_w14241_
	);
	LUT3 #(
		.INIT('h80)
	) name3729 (
		\wishbone_bd_ram_mem2_reg[30][20]/P0001 ,
		_w11935_,
		_w11948_,
		_w14242_
	);
	LUT3 #(
		.INIT('h80)
	) name3730 (
		\wishbone_bd_ram_mem2_reg[5][20]/P0001 ,
		_w11932_,
		_w11933_,
		_w14243_
	);
	LUT4 #(
		.INIT('h0001)
	) name3731 (
		_w14240_,
		_w14241_,
		_w14242_,
		_w14243_,
		_w14244_
	);
	LUT3 #(
		.INIT('h80)
	) name3732 (
		\wishbone_bd_ram_mem2_reg[219][20]/P0001 ,
		_w11936_,
		_w11984_,
		_w14245_
	);
	LUT3 #(
		.INIT('h80)
	) name3733 (
		\wishbone_bd_ram_mem2_reg[189][20]/P0001 ,
		_w11942_,
		_w11966_,
		_w14246_
	);
	LUT3 #(
		.INIT('h80)
	) name3734 (
		\wishbone_bd_ram_mem2_reg[217][20]/P0001 ,
		_w11968_,
		_w11984_,
		_w14247_
	);
	LUT3 #(
		.INIT('h80)
	) name3735 (
		\wishbone_bd_ram_mem2_reg[26][20]/P0001 ,
		_w11935_,
		_w11944_,
		_w14248_
	);
	LUT4 #(
		.INIT('h0001)
	) name3736 (
		_w14245_,
		_w14246_,
		_w14247_,
		_w14248_,
		_w14249_
	);
	LUT3 #(
		.INIT('h80)
	) name3737 (
		\wishbone_bd_ram_mem2_reg[82][20]/P0001 ,
		_w11963_,
		_w11972_,
		_w14250_
	);
	LUT3 #(
		.INIT('h80)
	) name3738 (
		\wishbone_bd_ram_mem2_reg[202][20]/P0001 ,
		_w11944_,
		_w11945_,
		_w14251_
	);
	LUT3 #(
		.INIT('h80)
	) name3739 (
		\wishbone_bd_ram_mem2_reg[18][20]/P0001 ,
		_w11935_,
		_w11963_,
		_w14252_
	);
	LUT3 #(
		.INIT('h80)
	) name3740 (
		\wishbone_bd_ram_mem2_reg[108][20]/P0001 ,
		_w11954_,
		_w11965_,
		_w14253_
	);
	LUT4 #(
		.INIT('h0001)
	) name3741 (
		_w14250_,
		_w14251_,
		_w14252_,
		_w14253_,
		_w14254_
	);
	LUT4 #(
		.INIT('h8000)
	) name3742 (
		_w14239_,
		_w14244_,
		_w14249_,
		_w14254_,
		_w14255_
	);
	LUT4 #(
		.INIT('h8000)
	) name3743 (
		_w14192_,
		_w14213_,
		_w14234_,
		_w14255_,
		_w14256_
	);
	LUT3 #(
		.INIT('h80)
	) name3744 (
		\wishbone_bd_ram_mem2_reg[120][20]/P0001 ,
		_w11990_,
		_w12012_,
		_w14257_
	);
	LUT3 #(
		.INIT('h80)
	) name3745 (
		\wishbone_bd_ram_mem2_reg[239][20]/P0001 ,
		_w11973_,
		_w11982_,
		_w14258_
	);
	LUT3 #(
		.INIT('h80)
	) name3746 (
		\wishbone_bd_ram_mem2_reg[16][20]/P0001 ,
		_w11935_,
		_w11941_,
		_w14259_
	);
	LUT3 #(
		.INIT('h80)
	) name3747 (
		\wishbone_bd_ram_mem2_reg[79][20]/P0001 ,
		_w11949_,
		_w11973_,
		_w14260_
	);
	LUT4 #(
		.INIT('h0001)
	) name3748 (
		_w14257_,
		_w14258_,
		_w14259_,
		_w14260_,
		_w14261_
	);
	LUT3 #(
		.INIT('h80)
	) name3749 (
		\wishbone_bd_ram_mem2_reg[56][20]/P0001 ,
		_w11979_,
		_w11990_,
		_w14262_
	);
	LUT3 #(
		.INIT('h80)
	) name3750 (
		\wishbone_bd_ram_mem2_reg[100][20]/P0001 ,
		_w11929_,
		_w11965_,
		_w14263_
	);
	LUT3 #(
		.INIT('h80)
	) name3751 (
		\wishbone_bd_ram_mem2_reg[127][20]/P0001 ,
		_w11973_,
		_w12012_,
		_w14264_
	);
	LUT3 #(
		.INIT('h80)
	) name3752 (
		\wishbone_bd_ram_mem2_reg[144][20]/P0001 ,
		_w11941_,
		_w11959_,
		_w14265_
	);
	LUT4 #(
		.INIT('h0001)
	) name3753 (
		_w14262_,
		_w14263_,
		_w14264_,
		_w14265_,
		_w14266_
	);
	LUT3 #(
		.INIT('h80)
	) name3754 (
		\wishbone_bd_ram_mem2_reg[206][20]/P0001 ,
		_w11945_,
		_w11948_,
		_w14267_
	);
	LUT3 #(
		.INIT('h80)
	) name3755 (
		\wishbone_bd_ram_mem2_reg[169][20]/P0001 ,
		_w11930_,
		_w11968_,
		_w14268_
	);
	LUT3 #(
		.INIT('h80)
	) name3756 (
		\wishbone_bd_ram_mem2_reg[250][20]/P0001 ,
		_w11944_,
		_w11952_,
		_w14269_
	);
	LUT3 #(
		.INIT('h80)
	) name3757 (
		\wishbone_bd_ram_mem2_reg[38][20]/P0001 ,
		_w11957_,
		_w11986_,
		_w14270_
	);
	LUT4 #(
		.INIT('h0001)
	) name3758 (
		_w14267_,
		_w14268_,
		_w14269_,
		_w14270_,
		_w14271_
	);
	LUT3 #(
		.INIT('h80)
	) name3759 (
		\wishbone_bd_ram_mem2_reg[76][20]/P0001 ,
		_w11949_,
		_w11954_,
		_w14272_
	);
	LUT3 #(
		.INIT('h80)
	) name3760 (
		\wishbone_bd_ram_mem2_reg[39][20]/P0001 ,
		_w11957_,
		_w11975_,
		_w14273_
	);
	LUT3 #(
		.INIT('h80)
	) name3761 (
		\wishbone_bd_ram_mem2_reg[145][20]/P0001 ,
		_w11959_,
		_w11977_,
		_w14274_
	);
	LUT3 #(
		.INIT('h80)
	) name3762 (
		\wishbone_bd_ram_mem2_reg[111][20]/P0001 ,
		_w11965_,
		_w11973_,
		_w14275_
	);
	LUT4 #(
		.INIT('h0001)
	) name3763 (
		_w14272_,
		_w14273_,
		_w14274_,
		_w14275_,
		_w14276_
	);
	LUT4 #(
		.INIT('h8000)
	) name3764 (
		_w14261_,
		_w14266_,
		_w14271_,
		_w14276_,
		_w14277_
	);
	LUT3 #(
		.INIT('h80)
	) name3765 (
		\wishbone_bd_ram_mem2_reg[203][20]/P0001 ,
		_w11936_,
		_w11945_,
		_w14278_
	);
	LUT3 #(
		.INIT('h80)
	) name3766 (
		\wishbone_bd_ram_mem2_reg[118][20]/P0001 ,
		_w11986_,
		_w12012_,
		_w14279_
	);
	LUT3 #(
		.INIT('h80)
	) name3767 (
		\wishbone_bd_ram_mem2_reg[231][20]/P0001 ,
		_w11975_,
		_w11982_,
		_w14280_
	);
	LUT3 #(
		.INIT('h80)
	) name3768 (
		\wishbone_bd_ram_mem2_reg[15][20]/P0001 ,
		_w11932_,
		_w11973_,
		_w14281_
	);
	LUT4 #(
		.INIT('h0001)
	) name3769 (
		_w14278_,
		_w14279_,
		_w14280_,
		_w14281_,
		_w14282_
	);
	LUT3 #(
		.INIT('h80)
	) name3770 (
		\wishbone_bd_ram_mem2_reg[177][20]/P0001 ,
		_w11942_,
		_w11977_,
		_w14283_
	);
	LUT3 #(
		.INIT('h80)
	) name3771 (
		\wishbone_bd_ram_mem2_reg[166][20]/P0001 ,
		_w11930_,
		_w11986_,
		_w14284_
	);
	LUT3 #(
		.INIT('h80)
	) name3772 (
		\wishbone_bd_ram_mem2_reg[149][20]/P0001 ,
		_w11933_,
		_w11959_,
		_w14285_
	);
	LUT3 #(
		.INIT('h80)
	) name3773 (
		\wishbone_bd_ram_mem2_reg[121][20]/P0001 ,
		_w11968_,
		_w12012_,
		_w14286_
	);
	LUT4 #(
		.INIT('h0001)
	) name3774 (
		_w14283_,
		_w14284_,
		_w14285_,
		_w14286_,
		_w14287_
	);
	LUT3 #(
		.INIT('h80)
	) name3775 (
		\wishbone_bd_ram_mem2_reg[37][20]/P0001 ,
		_w11933_,
		_w11957_,
		_w14288_
	);
	LUT3 #(
		.INIT('h80)
	) name3776 (
		\wishbone_bd_ram_mem2_reg[234][20]/P0001 ,
		_w11944_,
		_w11982_,
		_w14289_
	);
	LUT3 #(
		.INIT('h80)
	) name3777 (
		\wishbone_bd_ram_mem2_reg[20][20]/P0001 ,
		_w11929_,
		_w11935_,
		_w14290_
	);
	LUT3 #(
		.INIT('h80)
	) name3778 (
		\wishbone_bd_ram_mem2_reg[147][20]/P0001 ,
		_w11938_,
		_w11959_,
		_w14291_
	);
	LUT4 #(
		.INIT('h0001)
	) name3779 (
		_w14288_,
		_w14289_,
		_w14290_,
		_w14291_,
		_w14292_
	);
	LUT3 #(
		.INIT('h80)
	) name3780 (
		\wishbone_bd_ram_mem2_reg[64][20]/P0001 ,
		_w11941_,
		_w11949_,
		_w14293_
	);
	LUT3 #(
		.INIT('h80)
	) name3781 (
		\wishbone_bd_ram_mem2_reg[225][20]/P0001 ,
		_w11977_,
		_w11982_,
		_w14294_
	);
	LUT3 #(
		.INIT('h80)
	) name3782 (
		\wishbone_bd_ram_mem2_reg[85][20]/P0001 ,
		_w11933_,
		_w11972_,
		_w14295_
	);
	LUT3 #(
		.INIT('h80)
	) name3783 (
		\wishbone_bd_ram_mem2_reg[237][20]/P0001 ,
		_w11966_,
		_w11982_,
		_w14296_
	);
	LUT4 #(
		.INIT('h0001)
	) name3784 (
		_w14293_,
		_w14294_,
		_w14295_,
		_w14296_,
		_w14297_
	);
	LUT4 #(
		.INIT('h8000)
	) name3785 (
		_w14282_,
		_w14287_,
		_w14292_,
		_w14297_,
		_w14298_
	);
	LUT3 #(
		.INIT('h80)
	) name3786 (
		\wishbone_bd_ram_mem2_reg[124][20]/P0001 ,
		_w11954_,
		_w12012_,
		_w14299_
	);
	LUT3 #(
		.INIT('h80)
	) name3787 (
		\wishbone_bd_ram_mem2_reg[71][20]/P0001 ,
		_w11949_,
		_w11975_,
		_w14300_
	);
	LUT3 #(
		.INIT('h80)
	) name3788 (
		\wishbone_bd_ram_mem2_reg[223][20]/P0001 ,
		_w11973_,
		_w11984_,
		_w14301_
	);
	LUT3 #(
		.INIT('h80)
	) name3789 (
		\wishbone_bd_ram_mem2_reg[242][20]/P0001 ,
		_w11952_,
		_w11963_,
		_w14302_
	);
	LUT4 #(
		.INIT('h0001)
	) name3790 (
		_w14299_,
		_w14300_,
		_w14301_,
		_w14302_,
		_w14303_
	);
	LUT3 #(
		.INIT('h80)
	) name3791 (
		\wishbone_bd_ram_mem2_reg[114][20]/P0001 ,
		_w11963_,
		_w12012_,
		_w14304_
	);
	LUT3 #(
		.INIT('h80)
	) name3792 (
		\wishbone_bd_ram_mem2_reg[168][20]/P0001 ,
		_w11930_,
		_w11990_,
		_w14305_
	);
	LUT3 #(
		.INIT('h80)
	) name3793 (
		\wishbone_bd_ram_mem2_reg[96][20]/P0001 ,
		_w11941_,
		_w11965_,
		_w14306_
	);
	LUT3 #(
		.INIT('h80)
	) name3794 (
		\wishbone_bd_ram_mem2_reg[247][20]/P0001 ,
		_w11952_,
		_w11975_,
		_w14307_
	);
	LUT4 #(
		.INIT('h0001)
	) name3795 (
		_w14304_,
		_w14305_,
		_w14306_,
		_w14307_,
		_w14308_
	);
	LUT3 #(
		.INIT('h80)
	) name3796 (
		\wishbone_bd_ram_mem2_reg[198][20]/P0001 ,
		_w11945_,
		_w11986_,
		_w14309_
	);
	LUT3 #(
		.INIT('h80)
	) name3797 (
		\wishbone_bd_ram_mem2_reg[128][20]/P0001 ,
		_w11941_,
		_w11955_,
		_w14310_
	);
	LUT3 #(
		.INIT('h80)
	) name3798 (
		\wishbone_bd_ram_mem2_reg[112][20]/P0001 ,
		_w11941_,
		_w12012_,
		_w14311_
	);
	LUT3 #(
		.INIT('h80)
	) name3799 (
		\wishbone_bd_ram_mem2_reg[44][20]/P0001 ,
		_w11954_,
		_w11957_,
		_w14312_
	);
	LUT4 #(
		.INIT('h0001)
	) name3800 (
		_w14309_,
		_w14310_,
		_w14311_,
		_w14312_,
		_w14313_
	);
	LUT3 #(
		.INIT('h80)
	) name3801 (
		\wishbone_bd_ram_mem2_reg[160][20]/P0001 ,
		_w11930_,
		_w11941_,
		_w14314_
	);
	LUT3 #(
		.INIT('h80)
	) name3802 (
		\wishbone_bd_ram_mem2_reg[92][20]/P0001 ,
		_w11954_,
		_w11972_,
		_w14315_
	);
	LUT3 #(
		.INIT('h80)
	) name3803 (
		\wishbone_bd_ram_mem2_reg[210][20]/P0001 ,
		_w11963_,
		_w11984_,
		_w14316_
	);
	LUT3 #(
		.INIT('h80)
	) name3804 (
		\wishbone_bd_ram_mem2_reg[254][20]/P0001 ,
		_w11948_,
		_w11952_,
		_w14317_
	);
	LUT4 #(
		.INIT('h0001)
	) name3805 (
		_w14314_,
		_w14315_,
		_w14316_,
		_w14317_,
		_w14318_
	);
	LUT4 #(
		.INIT('h8000)
	) name3806 (
		_w14303_,
		_w14308_,
		_w14313_,
		_w14318_,
		_w14319_
	);
	LUT3 #(
		.INIT('h80)
	) name3807 (
		\wishbone_bd_ram_mem2_reg[57][20]/P0001 ,
		_w11968_,
		_w11979_,
		_w14320_
	);
	LUT3 #(
		.INIT('h80)
	) name3808 (
		\wishbone_bd_ram_mem2_reg[101][20]/P0001 ,
		_w11933_,
		_w11965_,
		_w14321_
	);
	LUT3 #(
		.INIT('h80)
	) name3809 (
		\wishbone_bd_ram_mem2_reg[70][20]/P0001 ,
		_w11949_,
		_w11986_,
		_w14322_
	);
	LUT3 #(
		.INIT('h80)
	) name3810 (
		\wishbone_bd_ram_mem2_reg[150][20]/P0001 ,
		_w11959_,
		_w11986_,
		_w14323_
	);
	LUT4 #(
		.INIT('h0001)
	) name3811 (
		_w14320_,
		_w14321_,
		_w14322_,
		_w14323_,
		_w14324_
	);
	LUT3 #(
		.INIT('h80)
	) name3812 (
		\wishbone_bd_ram_mem2_reg[115][20]/P0001 ,
		_w11938_,
		_w12012_,
		_w14325_
	);
	LUT3 #(
		.INIT('h80)
	) name3813 (
		\wishbone_bd_ram_mem2_reg[154][20]/P0001 ,
		_w11944_,
		_w11959_,
		_w14326_
	);
	LUT3 #(
		.INIT('h80)
	) name3814 (
		\wishbone_bd_ram_mem2_reg[105][20]/P0001 ,
		_w11965_,
		_w11968_,
		_w14327_
	);
	LUT3 #(
		.INIT('h80)
	) name3815 (
		\wishbone_bd_ram_mem2_reg[152][20]/P0001 ,
		_w11959_,
		_w11990_,
		_w14328_
	);
	LUT4 #(
		.INIT('h0001)
	) name3816 (
		_w14325_,
		_w14326_,
		_w14327_,
		_w14328_,
		_w14329_
	);
	LUT3 #(
		.INIT('h80)
	) name3817 (
		\wishbone_bd_ram_mem2_reg[21][20]/P0001 ,
		_w11933_,
		_w11935_,
		_w14330_
	);
	LUT3 #(
		.INIT('h80)
	) name3818 (
		\wishbone_bd_ram_mem2_reg[201][20]/P0001 ,
		_w11945_,
		_w11968_,
		_w14331_
	);
	LUT3 #(
		.INIT('h80)
	) name3819 (
		\wishbone_bd_ram_mem2_reg[190][20]/P0001 ,
		_w11942_,
		_w11948_,
		_w14332_
	);
	LUT3 #(
		.INIT('h80)
	) name3820 (
		\wishbone_bd_ram_mem2_reg[22][20]/P0001 ,
		_w11935_,
		_w11986_,
		_w14333_
	);
	LUT4 #(
		.INIT('h0001)
	) name3821 (
		_w14330_,
		_w14331_,
		_w14332_,
		_w14333_,
		_w14334_
	);
	LUT3 #(
		.INIT('h80)
	) name3822 (
		\wishbone_bd_ram_mem2_reg[173][20]/P0001 ,
		_w11930_,
		_w11966_,
		_w14335_
	);
	LUT3 #(
		.INIT('h80)
	) name3823 (
		\wishbone_bd_ram_mem2_reg[142][20]/P0001 ,
		_w11948_,
		_w11955_,
		_w14336_
	);
	LUT3 #(
		.INIT('h80)
	) name3824 (
		\wishbone_bd_ram_mem2_reg[106][20]/P0001 ,
		_w11944_,
		_w11965_,
		_w14337_
	);
	LUT3 #(
		.INIT('h80)
	) name3825 (
		\wishbone_bd_ram_mem2_reg[148][20]/P0001 ,
		_w11929_,
		_w11959_,
		_w14338_
	);
	LUT4 #(
		.INIT('h0001)
	) name3826 (
		_w14335_,
		_w14336_,
		_w14337_,
		_w14338_,
		_w14339_
	);
	LUT4 #(
		.INIT('h8000)
	) name3827 (
		_w14324_,
		_w14329_,
		_w14334_,
		_w14339_,
		_w14340_
	);
	LUT4 #(
		.INIT('h8000)
	) name3828 (
		_w14277_,
		_w14298_,
		_w14319_,
		_w14340_,
		_w14341_
	);
	LUT3 #(
		.INIT('h80)
	) name3829 (
		\wishbone_bd_ram_mem2_reg[84][20]/P0001 ,
		_w11929_,
		_w11972_,
		_w14342_
	);
	LUT3 #(
		.INIT('h80)
	) name3830 (
		\wishbone_bd_ram_mem2_reg[102][20]/P0001 ,
		_w11965_,
		_w11986_,
		_w14343_
	);
	LUT3 #(
		.INIT('h80)
	) name3831 (
		\wishbone_bd_ram_mem2_reg[139][20]/P0001 ,
		_w11936_,
		_w11955_,
		_w14344_
	);
	LUT3 #(
		.INIT('h80)
	) name3832 (
		\wishbone_bd_ram_mem2_reg[66][20]/P0001 ,
		_w11949_,
		_w11963_,
		_w14345_
	);
	LUT4 #(
		.INIT('h0001)
	) name3833 (
		_w14342_,
		_w14343_,
		_w14344_,
		_w14345_,
		_w14346_
	);
	LUT3 #(
		.INIT('h80)
	) name3834 (
		\wishbone_bd_ram_mem2_reg[185][20]/P0001 ,
		_w11942_,
		_w11968_,
		_w14347_
	);
	LUT3 #(
		.INIT('h80)
	) name3835 (
		\wishbone_bd_ram_mem2_reg[1][20]/P0001 ,
		_w11932_,
		_w11977_,
		_w14348_
	);
	LUT3 #(
		.INIT('h80)
	) name3836 (
		\wishbone_bd_ram_mem2_reg[23][20]/P0001 ,
		_w11935_,
		_w11975_,
		_w14349_
	);
	LUT3 #(
		.INIT('h80)
	) name3837 (
		\wishbone_bd_ram_mem2_reg[129][20]/P0001 ,
		_w11955_,
		_w11977_,
		_w14350_
	);
	LUT4 #(
		.INIT('h0001)
	) name3838 (
		_w14347_,
		_w14348_,
		_w14349_,
		_w14350_,
		_w14351_
	);
	LUT3 #(
		.INIT('h80)
	) name3839 (
		\wishbone_bd_ram_mem2_reg[69][20]/P0001 ,
		_w11933_,
		_w11949_,
		_w14352_
	);
	LUT3 #(
		.INIT('h80)
	) name3840 (
		\wishbone_bd_ram_mem2_reg[197][20]/P0001 ,
		_w11933_,
		_w11945_,
		_w14353_
	);
	LUT3 #(
		.INIT('h80)
	) name3841 (
		\wishbone_bd_ram_mem2_reg[72][20]/P0001 ,
		_w11949_,
		_w11990_,
		_w14354_
	);
	LUT3 #(
		.INIT('h80)
	) name3842 (
		\wishbone_bd_ram_mem2_reg[94][20]/P0001 ,
		_w11948_,
		_w11972_,
		_w14355_
	);
	LUT4 #(
		.INIT('h0001)
	) name3843 (
		_w14352_,
		_w14353_,
		_w14354_,
		_w14355_,
		_w14356_
	);
	LUT3 #(
		.INIT('h80)
	) name3844 (
		\wishbone_bd_ram_mem2_reg[205][20]/P0001 ,
		_w11945_,
		_w11966_,
		_w14357_
	);
	LUT3 #(
		.INIT('h80)
	) name3845 (
		\wishbone_bd_ram_mem2_reg[130][20]/P0001 ,
		_w11955_,
		_w11963_,
		_w14358_
	);
	LUT3 #(
		.INIT('h80)
	) name3846 (
		\wishbone_bd_ram_mem2_reg[163][20]/P0001 ,
		_w11930_,
		_w11938_,
		_w14359_
	);
	LUT3 #(
		.INIT('h80)
	) name3847 (
		\wishbone_bd_ram_mem2_reg[253][20]/P0001 ,
		_w11952_,
		_w11966_,
		_w14360_
	);
	LUT4 #(
		.INIT('h0001)
	) name3848 (
		_w14357_,
		_w14358_,
		_w14359_,
		_w14360_,
		_w14361_
	);
	LUT4 #(
		.INIT('h8000)
	) name3849 (
		_w14346_,
		_w14351_,
		_w14356_,
		_w14361_,
		_w14362_
	);
	LUT3 #(
		.INIT('h80)
	) name3850 (
		\wishbone_bd_ram_mem2_reg[240][20]/P0001 ,
		_w11941_,
		_w11952_,
		_w14363_
	);
	LUT3 #(
		.INIT('h80)
	) name3851 (
		\wishbone_bd_ram_mem2_reg[243][20]/P0001 ,
		_w11938_,
		_w11952_,
		_w14364_
	);
	LUT3 #(
		.INIT('h80)
	) name3852 (
		\wishbone_bd_ram_mem2_reg[24][20]/P0001 ,
		_w11935_,
		_w11990_,
		_w14365_
	);
	LUT3 #(
		.INIT('h80)
	) name3853 (
		\wishbone_bd_ram_mem2_reg[103][20]/P0001 ,
		_w11965_,
		_w11975_,
		_w14366_
	);
	LUT4 #(
		.INIT('h0001)
	) name3854 (
		_w14363_,
		_w14364_,
		_w14365_,
		_w14366_,
		_w14367_
	);
	LUT3 #(
		.INIT('h80)
	) name3855 (
		\wishbone_bd_ram_mem2_reg[184][20]/P0001 ,
		_w11942_,
		_w11990_,
		_w14368_
	);
	LUT3 #(
		.INIT('h80)
	) name3856 (
		\wishbone_bd_ram_mem2_reg[110][20]/P0001 ,
		_w11948_,
		_w11965_,
		_w14369_
	);
	LUT3 #(
		.INIT('h80)
	) name3857 (
		\wishbone_bd_ram_mem2_reg[28][20]/P0001 ,
		_w11935_,
		_w11954_,
		_w14370_
	);
	LUT3 #(
		.INIT('h80)
	) name3858 (
		\wishbone_bd_ram_mem2_reg[91][20]/P0001 ,
		_w11936_,
		_w11972_,
		_w14371_
	);
	LUT4 #(
		.INIT('h0001)
	) name3859 (
		_w14368_,
		_w14369_,
		_w14370_,
		_w14371_,
		_w14372_
	);
	LUT3 #(
		.INIT('h80)
	) name3860 (
		\wishbone_bd_ram_mem2_reg[27][20]/P0001 ,
		_w11935_,
		_w11936_,
		_w14373_
	);
	LUT3 #(
		.INIT('h80)
	) name3861 (
		\wishbone_bd_ram_mem2_reg[170][20]/P0001 ,
		_w11930_,
		_w11944_,
		_w14374_
	);
	LUT3 #(
		.INIT('h80)
	) name3862 (
		\wishbone_bd_ram_mem2_reg[195][20]/P0001 ,
		_w11938_,
		_w11945_,
		_w14375_
	);
	LUT3 #(
		.INIT('h80)
	) name3863 (
		\wishbone_bd_ram_mem2_reg[233][20]/P0001 ,
		_w11968_,
		_w11982_,
		_w14376_
	);
	LUT4 #(
		.INIT('h0001)
	) name3864 (
		_w14373_,
		_w14374_,
		_w14375_,
		_w14376_,
		_w14377_
	);
	LUT3 #(
		.INIT('h80)
	) name3865 (
		\wishbone_bd_ram_mem2_reg[7][20]/P0001 ,
		_w11932_,
		_w11975_,
		_w14378_
	);
	LUT3 #(
		.INIT('h80)
	) name3866 (
		\wishbone_bd_ram_mem2_reg[97][20]/P0001 ,
		_w11965_,
		_w11977_,
		_w14379_
	);
	LUT3 #(
		.INIT('h80)
	) name3867 (
		\wishbone_bd_ram_mem2_reg[31][20]/P0001 ,
		_w11935_,
		_w11973_,
		_w14380_
	);
	LUT3 #(
		.INIT('h80)
	) name3868 (
		\wishbone_bd_ram_mem2_reg[54][20]/P0001 ,
		_w11979_,
		_w11986_,
		_w14381_
	);
	LUT4 #(
		.INIT('h0001)
	) name3869 (
		_w14378_,
		_w14379_,
		_w14380_,
		_w14381_,
		_w14382_
	);
	LUT4 #(
		.INIT('h8000)
	) name3870 (
		_w14367_,
		_w14372_,
		_w14377_,
		_w14382_,
		_w14383_
	);
	LUT3 #(
		.INIT('h80)
	) name3871 (
		\wishbone_bd_ram_mem2_reg[46][20]/P0001 ,
		_w11948_,
		_w11957_,
		_w14384_
	);
	LUT3 #(
		.INIT('h80)
	) name3872 (
		\wishbone_bd_ram_mem2_reg[207][20]/P0001 ,
		_w11945_,
		_w11973_,
		_w14385_
	);
	LUT3 #(
		.INIT('h80)
	) name3873 (
		\wishbone_bd_ram_mem2_reg[212][20]/P0001 ,
		_w11929_,
		_w11984_,
		_w14386_
	);
	LUT3 #(
		.INIT('h80)
	) name3874 (
		\wishbone_bd_ram_mem2_reg[62][20]/P0001 ,
		_w11948_,
		_w11979_,
		_w14387_
	);
	LUT4 #(
		.INIT('h0001)
	) name3875 (
		_w14384_,
		_w14385_,
		_w14386_,
		_w14387_,
		_w14388_
	);
	LUT3 #(
		.INIT('h80)
	) name3876 (
		\wishbone_bd_ram_mem2_reg[75][20]/P0001 ,
		_w11936_,
		_w11949_,
		_w14389_
	);
	LUT3 #(
		.INIT('h80)
	) name3877 (
		\wishbone_bd_ram_mem2_reg[161][20]/P0001 ,
		_w11930_,
		_w11977_,
		_w14390_
	);
	LUT3 #(
		.INIT('h80)
	) name3878 (
		\wishbone_bd_ram_mem2_reg[36][20]/P0001 ,
		_w11929_,
		_w11957_,
		_w14391_
	);
	LUT3 #(
		.INIT('h80)
	) name3879 (
		\wishbone_bd_ram_mem2_reg[51][20]/P0001 ,
		_w11938_,
		_w11979_,
		_w14392_
	);
	LUT4 #(
		.INIT('h0001)
	) name3880 (
		_w14389_,
		_w14390_,
		_w14391_,
		_w14392_,
		_w14393_
	);
	LUT3 #(
		.INIT('h80)
	) name3881 (
		\wishbone_bd_ram_mem2_reg[80][20]/P0001 ,
		_w11941_,
		_w11972_,
		_w14394_
	);
	LUT3 #(
		.INIT('h80)
	) name3882 (
		\wishbone_bd_ram_mem2_reg[14][20]/P0001 ,
		_w11932_,
		_w11948_,
		_w14395_
	);
	LUT3 #(
		.INIT('h80)
	) name3883 (
		\wishbone_bd_ram_mem2_reg[200][20]/P0001 ,
		_w11945_,
		_w11990_,
		_w14396_
	);
	LUT3 #(
		.INIT('h80)
	) name3884 (
		\wishbone_bd_ram_mem2_reg[141][20]/P0001 ,
		_w11955_,
		_w11966_,
		_w14397_
	);
	LUT4 #(
		.INIT('h0001)
	) name3885 (
		_w14394_,
		_w14395_,
		_w14396_,
		_w14397_,
		_w14398_
	);
	LUT3 #(
		.INIT('h80)
	) name3886 (
		\wishbone_bd_ram_mem2_reg[88][20]/P0001 ,
		_w11972_,
		_w11990_,
		_w14399_
	);
	LUT3 #(
		.INIT('h80)
	) name3887 (
		\wishbone_bd_ram_mem2_reg[196][20]/P0001 ,
		_w11929_,
		_w11945_,
		_w14400_
	);
	LUT3 #(
		.INIT('h80)
	) name3888 (
		\wishbone_bd_ram_mem2_reg[238][20]/P0001 ,
		_w11948_,
		_w11982_,
		_w14401_
	);
	LUT3 #(
		.INIT('h80)
	) name3889 (
		\wishbone_bd_ram_mem2_reg[181][20]/P0001 ,
		_w11933_,
		_w11942_,
		_w14402_
	);
	LUT4 #(
		.INIT('h0001)
	) name3890 (
		_w14399_,
		_w14400_,
		_w14401_,
		_w14402_,
		_w14403_
	);
	LUT4 #(
		.INIT('h8000)
	) name3891 (
		_w14388_,
		_w14393_,
		_w14398_,
		_w14403_,
		_w14404_
	);
	LUT3 #(
		.INIT('h80)
	) name3892 (
		\wishbone_bd_ram_mem2_reg[179][20]/P0001 ,
		_w11938_,
		_w11942_,
		_w14405_
	);
	LUT3 #(
		.INIT('h80)
	) name3893 (
		\wishbone_bd_ram_mem2_reg[49][20]/P0001 ,
		_w11977_,
		_w11979_,
		_w14406_
	);
	LUT3 #(
		.INIT('h80)
	) name3894 (
		\wishbone_bd_ram_mem2_reg[117][20]/P0001 ,
		_w11933_,
		_w12012_,
		_w14407_
	);
	LUT3 #(
		.INIT('h80)
	) name3895 (
		\wishbone_bd_ram_mem2_reg[162][20]/P0001 ,
		_w11930_,
		_w11963_,
		_w14408_
	);
	LUT4 #(
		.INIT('h0001)
	) name3896 (
		_w14405_,
		_w14406_,
		_w14407_,
		_w14408_,
		_w14409_
	);
	LUT3 #(
		.INIT('h80)
	) name3897 (
		\wishbone_bd_ram_mem2_reg[60][20]/P0001 ,
		_w11954_,
		_w11979_,
		_w14410_
	);
	LUT3 #(
		.INIT('h80)
	) name3898 (
		\wishbone_bd_ram_mem2_reg[255][20]/P0001 ,
		_w11952_,
		_w11973_,
		_w14411_
	);
	LUT3 #(
		.INIT('h80)
	) name3899 (
		\wishbone_bd_ram_mem2_reg[249][20]/P0001 ,
		_w11952_,
		_w11968_,
		_w14412_
	);
	LUT3 #(
		.INIT('h80)
	) name3900 (
		\wishbone_bd_ram_mem2_reg[42][20]/P0001 ,
		_w11944_,
		_w11957_,
		_w14413_
	);
	LUT4 #(
		.INIT('h0001)
	) name3901 (
		_w14410_,
		_w14411_,
		_w14412_,
		_w14413_,
		_w14414_
	);
	LUT3 #(
		.INIT('h80)
	) name3902 (
		\wishbone_bd_ram_mem2_reg[214][20]/P0001 ,
		_w11984_,
		_w11986_,
		_w14415_
	);
	LUT3 #(
		.INIT('h80)
	) name3903 (
		\wishbone_bd_ram_mem2_reg[107][20]/P0001 ,
		_w11936_,
		_w11965_,
		_w14416_
	);
	LUT3 #(
		.INIT('h80)
	) name3904 (
		\wishbone_bd_ram_mem2_reg[188][20]/P0001 ,
		_w11942_,
		_w11954_,
		_w14417_
	);
	LUT3 #(
		.INIT('h80)
	) name3905 (
		\wishbone_bd_ram_mem2_reg[25][20]/P0001 ,
		_w11935_,
		_w11968_,
		_w14418_
	);
	LUT4 #(
		.INIT('h0001)
	) name3906 (
		_w14415_,
		_w14416_,
		_w14417_,
		_w14418_,
		_w14419_
	);
	LUT3 #(
		.INIT('h80)
	) name3907 (
		\wishbone_bd_ram_mem2_reg[186][20]/P0001 ,
		_w11942_,
		_w11944_,
		_w14420_
	);
	LUT3 #(
		.INIT('h80)
	) name3908 (
		\wishbone_bd_ram_mem2_reg[47][20]/P0001 ,
		_w11957_,
		_w11973_,
		_w14421_
	);
	LUT3 #(
		.INIT('h80)
	) name3909 (
		\wishbone_bd_ram_mem2_reg[151][20]/P0001 ,
		_w11959_,
		_w11975_,
		_w14422_
	);
	LUT3 #(
		.INIT('h80)
	) name3910 (
		\wishbone_bd_ram_mem2_reg[95][20]/P0001 ,
		_w11972_,
		_w11973_,
		_w14423_
	);
	LUT4 #(
		.INIT('h0001)
	) name3911 (
		_w14420_,
		_w14421_,
		_w14422_,
		_w14423_,
		_w14424_
	);
	LUT4 #(
		.INIT('h8000)
	) name3912 (
		_w14409_,
		_w14414_,
		_w14419_,
		_w14424_,
		_w14425_
	);
	LUT4 #(
		.INIT('h8000)
	) name3913 (
		_w14362_,
		_w14383_,
		_w14404_,
		_w14425_,
		_w14426_
	);
	LUT3 #(
		.INIT('h80)
	) name3914 (
		\wishbone_bd_ram_mem2_reg[209][20]/P0001 ,
		_w11977_,
		_w11984_,
		_w14427_
	);
	LUT3 #(
		.INIT('h80)
	) name3915 (
		\wishbone_bd_ram_mem2_reg[228][20]/P0001 ,
		_w11929_,
		_w11982_,
		_w14428_
	);
	LUT3 #(
		.INIT('h80)
	) name3916 (
		\wishbone_bd_ram_mem2_reg[246][20]/P0001 ,
		_w11952_,
		_w11986_,
		_w14429_
	);
	LUT3 #(
		.INIT('h80)
	) name3917 (
		\wishbone_bd_ram_mem2_reg[81][20]/P0001 ,
		_w11972_,
		_w11977_,
		_w14430_
	);
	LUT4 #(
		.INIT('h0001)
	) name3918 (
		_w14427_,
		_w14428_,
		_w14429_,
		_w14430_,
		_w14431_
	);
	LUT3 #(
		.INIT('h80)
	) name3919 (
		\wishbone_bd_ram_mem2_reg[68][20]/P0001 ,
		_w11929_,
		_w11949_,
		_w14432_
	);
	LUT3 #(
		.INIT('h80)
	) name3920 (
		\wishbone_bd_ram_mem2_reg[248][20]/P0001 ,
		_w11952_,
		_w11990_,
		_w14433_
	);
	LUT3 #(
		.INIT('h80)
	) name3921 (
		\wishbone_bd_ram_mem2_reg[230][20]/P0001 ,
		_w11982_,
		_w11986_,
		_w14434_
	);
	LUT3 #(
		.INIT('h80)
	) name3922 (
		\wishbone_bd_ram_mem2_reg[35][20]/P0001 ,
		_w11938_,
		_w11957_,
		_w14435_
	);
	LUT4 #(
		.INIT('h0001)
	) name3923 (
		_w14432_,
		_w14433_,
		_w14434_,
		_w14435_,
		_w14436_
	);
	LUT3 #(
		.INIT('h80)
	) name3924 (
		\wishbone_bd_ram_mem2_reg[176][20]/P0001 ,
		_w11941_,
		_w11942_,
		_w14437_
	);
	LUT3 #(
		.INIT('h80)
	) name3925 (
		\wishbone_bd_ram_mem2_reg[59][20]/P0001 ,
		_w11936_,
		_w11979_,
		_w14438_
	);
	LUT3 #(
		.INIT('h80)
	) name3926 (
		\wishbone_bd_ram_mem2_reg[226][20]/P0001 ,
		_w11963_,
		_w11982_,
		_w14439_
	);
	LUT3 #(
		.INIT('h80)
	) name3927 (
		\wishbone_bd_ram_mem2_reg[143][20]/P0001 ,
		_w11955_,
		_w11973_,
		_w14440_
	);
	LUT4 #(
		.INIT('h0001)
	) name3928 (
		_w14437_,
		_w14438_,
		_w14439_,
		_w14440_,
		_w14441_
	);
	LUT3 #(
		.INIT('h80)
	) name3929 (
		\wishbone_bd_ram_mem2_reg[216][20]/P0001 ,
		_w11984_,
		_w11990_,
		_w14442_
	);
	LUT3 #(
		.INIT('h80)
	) name3930 (
		\wishbone_bd_ram_mem2_reg[2][20]/P0001 ,
		_w11932_,
		_w11963_,
		_w14443_
	);
	LUT3 #(
		.INIT('h80)
	) name3931 (
		\wishbone_bd_ram_mem2_reg[178][20]/P0001 ,
		_w11942_,
		_w11963_,
		_w14444_
	);
	LUT3 #(
		.INIT('h80)
	) name3932 (
		\wishbone_bd_ram_mem2_reg[12][20]/P0001 ,
		_w11932_,
		_w11954_,
		_w14445_
	);
	LUT4 #(
		.INIT('h0001)
	) name3933 (
		_w14442_,
		_w14443_,
		_w14444_,
		_w14445_,
		_w14446_
	);
	LUT4 #(
		.INIT('h8000)
	) name3934 (
		_w14431_,
		_w14436_,
		_w14441_,
		_w14446_,
		_w14447_
	);
	LUT3 #(
		.INIT('h80)
	) name3935 (
		\wishbone_bd_ram_mem2_reg[61][20]/P0001 ,
		_w11966_,
		_w11979_,
		_w14448_
	);
	LUT3 #(
		.INIT('h80)
	) name3936 (
		\wishbone_bd_ram_mem2_reg[6][20]/P0001 ,
		_w11932_,
		_w11986_,
		_w14449_
	);
	LUT3 #(
		.INIT('h80)
	) name3937 (
		\wishbone_bd_ram_mem2_reg[191][20]/P0001 ,
		_w11942_,
		_w11973_,
		_w14450_
	);
	LUT3 #(
		.INIT('h80)
	) name3938 (
		\wishbone_bd_ram_mem2_reg[17][20]/P0001 ,
		_w11935_,
		_w11977_,
		_w14451_
	);
	LUT4 #(
		.INIT('h0001)
	) name3939 (
		_w14448_,
		_w14449_,
		_w14450_,
		_w14451_,
		_w14452_
	);
	LUT3 #(
		.INIT('h80)
	) name3940 (
		\wishbone_bd_ram_mem2_reg[192][20]/P0001 ,
		_w11941_,
		_w11945_,
		_w14453_
	);
	LUT3 #(
		.INIT('h80)
	) name3941 (
		\wishbone_bd_ram_mem2_reg[232][20]/P0001 ,
		_w11982_,
		_w11990_,
		_w14454_
	);
	LUT3 #(
		.INIT('h80)
	) name3942 (
		\wishbone_bd_ram_mem2_reg[11][20]/P0001 ,
		_w11932_,
		_w11936_,
		_w14455_
	);
	LUT3 #(
		.INIT('h80)
	) name3943 (
		\wishbone_bd_ram_mem2_reg[213][20]/P0001 ,
		_w11933_,
		_w11984_,
		_w14456_
	);
	LUT4 #(
		.INIT('h0001)
	) name3944 (
		_w14453_,
		_w14454_,
		_w14455_,
		_w14456_,
		_w14457_
	);
	LUT3 #(
		.INIT('h80)
	) name3945 (
		\wishbone_bd_ram_mem2_reg[224][20]/P0001 ,
		_w11941_,
		_w11982_,
		_w14458_
	);
	LUT3 #(
		.INIT('h80)
	) name3946 (
		\wishbone_bd_ram_mem2_reg[138][20]/P0001 ,
		_w11944_,
		_w11955_,
		_w14459_
	);
	LUT3 #(
		.INIT('h80)
	) name3947 (
		\wishbone_bd_ram_mem2_reg[221][20]/P0001 ,
		_w11966_,
		_w11984_,
		_w14460_
	);
	LUT3 #(
		.INIT('h80)
	) name3948 (
		\wishbone_bd_ram_mem2_reg[174][20]/P0001 ,
		_w11930_,
		_w11948_,
		_w14461_
	);
	LUT4 #(
		.INIT('h0001)
	) name3949 (
		_w14458_,
		_w14459_,
		_w14460_,
		_w14461_,
		_w14462_
	);
	LUT3 #(
		.INIT('h80)
	) name3950 (
		\wishbone_bd_ram_mem2_reg[199][20]/P0001 ,
		_w11945_,
		_w11975_,
		_w14463_
	);
	LUT3 #(
		.INIT('h80)
	) name3951 (
		\wishbone_bd_ram_mem2_reg[78][20]/P0001 ,
		_w11948_,
		_w11949_,
		_w14464_
	);
	LUT3 #(
		.INIT('h80)
	) name3952 (
		\wishbone_bd_ram_mem2_reg[251][20]/P0001 ,
		_w11936_,
		_w11952_,
		_w14465_
	);
	LUT3 #(
		.INIT('h80)
	) name3953 (
		\wishbone_bd_ram_mem2_reg[48][20]/P0001 ,
		_w11941_,
		_w11979_,
		_w14466_
	);
	LUT4 #(
		.INIT('h0001)
	) name3954 (
		_w14463_,
		_w14464_,
		_w14465_,
		_w14466_,
		_w14467_
	);
	LUT4 #(
		.INIT('h8000)
	) name3955 (
		_w14452_,
		_w14457_,
		_w14462_,
		_w14467_,
		_w14468_
	);
	LUT3 #(
		.INIT('h80)
	) name3956 (
		\wishbone_bd_ram_mem2_reg[52][20]/P0001 ,
		_w11929_,
		_w11979_,
		_w14469_
	);
	LUT3 #(
		.INIT('h80)
	) name3957 (
		\wishbone_bd_ram_mem2_reg[175][20]/P0001 ,
		_w11930_,
		_w11973_,
		_w14470_
	);
	LUT3 #(
		.INIT('h80)
	) name3958 (
		\wishbone_bd_ram_mem2_reg[156][20]/P0001 ,
		_w11954_,
		_w11959_,
		_w14471_
	);
	LUT3 #(
		.INIT('h80)
	) name3959 (
		\wishbone_bd_ram_mem2_reg[241][20]/P0001 ,
		_w11952_,
		_w11977_,
		_w14472_
	);
	LUT4 #(
		.INIT('h0001)
	) name3960 (
		_w14469_,
		_w14470_,
		_w14471_,
		_w14472_,
		_w14473_
	);
	LUT3 #(
		.INIT('h80)
	) name3961 (
		\wishbone_bd_ram_mem2_reg[58][20]/P0001 ,
		_w11944_,
		_w11979_,
		_w14474_
	);
	LUT3 #(
		.INIT('h80)
	) name3962 (
		\wishbone_bd_ram_mem2_reg[208][20]/P0001 ,
		_w11941_,
		_w11984_,
		_w14475_
	);
	LUT3 #(
		.INIT('h80)
	) name3963 (
		\wishbone_bd_ram_mem2_reg[187][20]/P0001 ,
		_w11936_,
		_w11942_,
		_w14476_
	);
	LUT3 #(
		.INIT('h80)
	) name3964 (
		\wishbone_bd_ram_mem2_reg[13][20]/P0001 ,
		_w11932_,
		_w11966_,
		_w14477_
	);
	LUT4 #(
		.INIT('h0001)
	) name3965 (
		_w14474_,
		_w14475_,
		_w14476_,
		_w14477_,
		_w14478_
	);
	LUT3 #(
		.INIT('h80)
	) name3966 (
		\wishbone_bd_ram_mem2_reg[183][20]/P0001 ,
		_w11942_,
		_w11975_,
		_w14479_
	);
	LUT3 #(
		.INIT('h80)
	) name3967 (
		\wishbone_bd_ram_mem2_reg[55][20]/P0001 ,
		_w11975_,
		_w11979_,
		_w14480_
	);
	LUT3 #(
		.INIT('h80)
	) name3968 (
		\wishbone_bd_ram_mem2_reg[50][20]/P0001 ,
		_w11963_,
		_w11979_,
		_w14481_
	);
	LUT3 #(
		.INIT('h80)
	) name3969 (
		\wishbone_bd_ram_mem2_reg[155][20]/P0001 ,
		_w11936_,
		_w11959_,
		_w14482_
	);
	LUT4 #(
		.INIT('h0001)
	) name3970 (
		_w14479_,
		_w14480_,
		_w14481_,
		_w14482_,
		_w14483_
	);
	LUT3 #(
		.INIT('h80)
	) name3971 (
		\wishbone_bd_ram_mem2_reg[159][20]/P0001 ,
		_w11959_,
		_w11973_,
		_w14484_
	);
	LUT3 #(
		.INIT('h80)
	) name3972 (
		\wishbone_bd_ram_mem2_reg[220][20]/P0001 ,
		_w11954_,
		_w11984_,
		_w14485_
	);
	LUT3 #(
		.INIT('h80)
	) name3973 (
		\wishbone_bd_ram_mem2_reg[218][20]/P0001 ,
		_w11944_,
		_w11984_,
		_w14486_
	);
	LUT3 #(
		.INIT('h80)
	) name3974 (
		\wishbone_bd_ram_mem2_reg[104][20]/P0001 ,
		_w11965_,
		_w11990_,
		_w14487_
	);
	LUT4 #(
		.INIT('h0001)
	) name3975 (
		_w14484_,
		_w14485_,
		_w14486_,
		_w14487_,
		_w14488_
	);
	LUT4 #(
		.INIT('h8000)
	) name3976 (
		_w14473_,
		_w14478_,
		_w14483_,
		_w14488_,
		_w14489_
	);
	LUT3 #(
		.INIT('h80)
	) name3977 (
		\wishbone_bd_ram_mem2_reg[98][20]/P0001 ,
		_w11963_,
		_w11965_,
		_w14490_
	);
	LUT3 #(
		.INIT('h80)
	) name3978 (
		\wishbone_bd_ram_mem2_reg[123][20]/P0001 ,
		_w11936_,
		_w12012_,
		_w14491_
	);
	LUT3 #(
		.INIT('h80)
	) name3979 (
		\wishbone_bd_ram_mem2_reg[171][20]/P0001 ,
		_w11930_,
		_w11936_,
		_w14492_
	);
	LUT3 #(
		.INIT('h80)
	) name3980 (
		\wishbone_bd_ram_mem2_reg[131][20]/P0001 ,
		_w11938_,
		_w11955_,
		_w14493_
	);
	LUT4 #(
		.INIT('h0001)
	) name3981 (
		_w14490_,
		_w14491_,
		_w14492_,
		_w14493_,
		_w14494_
	);
	LUT3 #(
		.INIT('h80)
	) name3982 (
		\wishbone_bd_ram_mem2_reg[93][20]/P0001 ,
		_w11966_,
		_w11972_,
		_w14495_
	);
	LUT3 #(
		.INIT('h80)
	) name3983 (
		\wishbone_bd_ram_mem2_reg[86][20]/P0001 ,
		_w11972_,
		_w11986_,
		_w14496_
	);
	LUT3 #(
		.INIT('h80)
	) name3984 (
		\wishbone_bd_ram_mem2_reg[63][20]/P0001 ,
		_w11973_,
		_w11979_,
		_w14497_
	);
	LUT3 #(
		.INIT('h80)
	) name3985 (
		\wishbone_bd_ram_mem2_reg[77][20]/P0001 ,
		_w11949_,
		_w11966_,
		_w14498_
	);
	LUT4 #(
		.INIT('h0001)
	) name3986 (
		_w14495_,
		_w14496_,
		_w14497_,
		_w14498_,
		_w14499_
	);
	LUT3 #(
		.INIT('h80)
	) name3987 (
		\wishbone_bd_ram_mem2_reg[227][20]/P0001 ,
		_w11938_,
		_w11982_,
		_w14500_
	);
	LUT3 #(
		.INIT('h80)
	) name3988 (
		\wishbone_bd_ram_mem2_reg[122][20]/P0001 ,
		_w11944_,
		_w12012_,
		_w14501_
	);
	LUT3 #(
		.INIT('h80)
	) name3989 (
		\wishbone_bd_ram_mem2_reg[167][20]/P0001 ,
		_w11930_,
		_w11975_,
		_w14502_
	);
	LUT3 #(
		.INIT('h80)
	) name3990 (
		\wishbone_bd_ram_mem2_reg[132][20]/P0001 ,
		_w11929_,
		_w11955_,
		_w14503_
	);
	LUT4 #(
		.INIT('h0001)
	) name3991 (
		_w14500_,
		_w14501_,
		_w14502_,
		_w14503_,
		_w14504_
	);
	LUT3 #(
		.INIT('h80)
	) name3992 (
		\wishbone_bd_ram_mem2_reg[74][20]/P0001 ,
		_w11944_,
		_w11949_,
		_w14505_
	);
	LUT3 #(
		.INIT('h80)
	) name3993 (
		\wishbone_bd_ram_mem2_reg[136][20]/P0001 ,
		_w11955_,
		_w11990_,
		_w14506_
	);
	LUT3 #(
		.INIT('h80)
	) name3994 (
		\wishbone_bd_ram_mem2_reg[182][20]/P0001 ,
		_w11942_,
		_w11986_,
		_w14507_
	);
	LUT3 #(
		.INIT('h80)
	) name3995 (
		\wishbone_bd_ram_mem2_reg[153][20]/P0001 ,
		_w11959_,
		_w11968_,
		_w14508_
	);
	LUT4 #(
		.INIT('h0001)
	) name3996 (
		_w14505_,
		_w14506_,
		_w14507_,
		_w14508_,
		_w14509_
	);
	LUT4 #(
		.INIT('h8000)
	) name3997 (
		_w14494_,
		_w14499_,
		_w14504_,
		_w14509_,
		_w14510_
	);
	LUT4 #(
		.INIT('h8000)
	) name3998 (
		_w14447_,
		_w14468_,
		_w14489_,
		_w14510_,
		_w14511_
	);
	LUT4 #(
		.INIT('h8000)
	) name3999 (
		_w14256_,
		_w14341_,
		_w14426_,
		_w14511_,
		_w14512_
	);
	LUT3 #(
		.INIT('h70)
	) name4000 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w14513_
	);
	LUT4 #(
		.INIT('hd111)
	) name4001 (
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w12304_,
		_w12312_,
		_w12317_,
		_w14514_
	);
	LUT3 #(
		.INIT('h1e)
	) name4002 (
		\wishbone_TxLength_reg[2]/NET0131 ,
		\wishbone_TxLength_reg[3]/NET0131 ,
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w14515_
	);
	LUT2 #(
		.INIT('h8)
	) name4003 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		_w14516_
	);
	LUT2 #(
		.INIT('h2)
	) name4004 (
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w14517_
	);
	LUT4 #(
		.INIT('ha600)
	) name4005 (
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w12308_,
		_w14516_,
		_w14517_,
		_w14518_
	);
	LUT2 #(
		.INIT('h8)
	) name4006 (
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w14519_
	);
	LUT2 #(
		.INIT('h1)
	) name4007 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		_w14520_
	);
	LUT4 #(
		.INIT('h0001)
	) name4008 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		\wishbone_TxLength_reg[2]/NET0131 ,
		\wishbone_TxLength_reg[3]/NET0131 ,
		_w14521_
	);
	LUT4 #(
		.INIT('h60a0)
	) name4009 (
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w12308_,
		_w14519_,
		_w14520_,
		_w14522_
	);
	LUT2 #(
		.INIT('h1)
	) name4010 (
		_w14518_,
		_w14522_,
		_w14523_
	);
	LUT2 #(
		.INIT('h1)
	) name4011 (
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w14524_
	);
	LUT2 #(
		.INIT('h4)
	) name4012 (
		_w14515_,
		_w14524_,
		_w14525_
	);
	LUT2 #(
		.INIT('h4)
	) name4013 (
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w14526_
	);
	LUT4 #(
		.INIT('h0001)
	) name4014 (
		\wishbone_TxLength_reg[1]/NET0131 ,
		\wishbone_TxLength_reg[2]/NET0131 ,
		\wishbone_TxLength_reg[3]/NET0131 ,
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w14527_
	);
	LUT4 #(
		.INIT('h63ff)
	) name4015 (
		\wishbone_TxLength_reg[1]/NET0131 ,
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w12308_,
		_w14526_,
		_w14528_
	);
	LUT3 #(
		.INIT('h10)
	) name4016 (
		_w14513_,
		_w14525_,
		_w14528_,
		_w14529_
	);
	LUT4 #(
		.INIT('h0111)
	) name4017 (
		_w12302_,
		_w14514_,
		_w14523_,
		_w14529_,
		_w14530_
	);
	LUT3 #(
		.INIT('hf2)
	) name4018 (
		_w12303_,
		_w14512_,
		_w14530_,
		_w14531_
	);
	LUT3 #(
		.INIT('h80)
	) name4019 (
		\wishbone_bd_ram_mem3_reg[57][26]/P0001 ,
		_w11968_,
		_w11979_,
		_w14532_
	);
	LUT3 #(
		.INIT('h80)
	) name4020 (
		\wishbone_bd_ram_mem3_reg[185][26]/P0001 ,
		_w11942_,
		_w11968_,
		_w14533_
	);
	LUT3 #(
		.INIT('h80)
	) name4021 (
		\wishbone_bd_ram_mem3_reg[189][26]/P0001 ,
		_w11942_,
		_w11966_,
		_w14534_
	);
	LUT3 #(
		.INIT('h80)
	) name4022 (
		\wishbone_bd_ram_mem3_reg[55][26]/P0001 ,
		_w11975_,
		_w11979_,
		_w14535_
	);
	LUT4 #(
		.INIT('h0001)
	) name4023 (
		_w14532_,
		_w14533_,
		_w14534_,
		_w14535_,
		_w14536_
	);
	LUT3 #(
		.INIT('h80)
	) name4024 (
		\wishbone_bd_ram_mem3_reg[36][26]/P0001 ,
		_w11929_,
		_w11957_,
		_w14537_
	);
	LUT3 #(
		.INIT('h80)
	) name4025 (
		\wishbone_bd_ram_mem3_reg[159][26]/P0001 ,
		_w11959_,
		_w11973_,
		_w14538_
	);
	LUT3 #(
		.INIT('h80)
	) name4026 (
		\wishbone_bd_ram_mem3_reg[64][26]/P0001 ,
		_w11941_,
		_w11949_,
		_w14539_
	);
	LUT3 #(
		.INIT('h80)
	) name4027 (
		\wishbone_bd_ram_mem3_reg[204][26]/P0001 ,
		_w11945_,
		_w11954_,
		_w14540_
	);
	LUT4 #(
		.INIT('h0001)
	) name4028 (
		_w14537_,
		_w14538_,
		_w14539_,
		_w14540_,
		_w14541_
	);
	LUT3 #(
		.INIT('h80)
	) name4029 (
		\wishbone_bd_ram_mem3_reg[201][26]/P0001 ,
		_w11945_,
		_w11968_,
		_w14542_
	);
	LUT3 #(
		.INIT('h80)
	) name4030 (
		\wishbone_bd_ram_mem3_reg[127][26]/P0001 ,
		_w11973_,
		_w12012_,
		_w14543_
	);
	LUT3 #(
		.INIT('h80)
	) name4031 (
		\wishbone_bd_ram_mem3_reg[86][26]/P0001 ,
		_w11972_,
		_w11986_,
		_w14544_
	);
	LUT3 #(
		.INIT('h80)
	) name4032 (
		\wishbone_bd_ram_mem3_reg[111][26]/P0001 ,
		_w11965_,
		_w11973_,
		_w14545_
	);
	LUT4 #(
		.INIT('h0001)
	) name4033 (
		_w14542_,
		_w14543_,
		_w14544_,
		_w14545_,
		_w14546_
	);
	LUT3 #(
		.INIT('h80)
	) name4034 (
		\wishbone_bd_ram_mem3_reg[63][26]/P0001 ,
		_w11973_,
		_w11979_,
		_w14547_
	);
	LUT3 #(
		.INIT('h80)
	) name4035 (
		\wishbone_bd_ram_mem3_reg[207][26]/P0001 ,
		_w11945_,
		_w11973_,
		_w14548_
	);
	LUT3 #(
		.INIT('h80)
	) name4036 (
		\wishbone_bd_ram_mem3_reg[254][26]/P0001 ,
		_w11948_,
		_w11952_,
		_w14549_
	);
	LUT3 #(
		.INIT('h80)
	) name4037 (
		\wishbone_bd_ram_mem3_reg[119][26]/P0001 ,
		_w11975_,
		_w12012_,
		_w14550_
	);
	LUT4 #(
		.INIT('h0001)
	) name4038 (
		_w14547_,
		_w14548_,
		_w14549_,
		_w14550_,
		_w14551_
	);
	LUT4 #(
		.INIT('h8000)
	) name4039 (
		_w14536_,
		_w14541_,
		_w14546_,
		_w14551_,
		_w14552_
	);
	LUT3 #(
		.INIT('h80)
	) name4040 (
		\wishbone_bd_ram_mem3_reg[90][26]/P0001 ,
		_w11944_,
		_w11972_,
		_w14553_
	);
	LUT3 #(
		.INIT('h80)
	) name4041 (
		\wishbone_bd_ram_mem3_reg[143][26]/P0001 ,
		_w11955_,
		_w11973_,
		_w14554_
	);
	LUT3 #(
		.INIT('h80)
	) name4042 (
		\wishbone_bd_ram_mem3_reg[160][26]/P0001 ,
		_w11930_,
		_w11941_,
		_w14555_
	);
	LUT3 #(
		.INIT('h80)
	) name4043 (
		\wishbone_bd_ram_mem3_reg[75][26]/P0001 ,
		_w11936_,
		_w11949_,
		_w14556_
	);
	LUT4 #(
		.INIT('h0001)
	) name4044 (
		_w14553_,
		_w14554_,
		_w14555_,
		_w14556_,
		_w14557_
	);
	LUT3 #(
		.INIT('h80)
	) name4045 (
		\wishbone_bd_ram_mem3_reg[248][26]/P0001 ,
		_w11952_,
		_w11990_,
		_w14558_
	);
	LUT3 #(
		.INIT('h80)
	) name4046 (
		\wishbone_bd_ram_mem3_reg[209][26]/P0001 ,
		_w11977_,
		_w11984_,
		_w14559_
	);
	LUT3 #(
		.INIT('h80)
	) name4047 (
		\wishbone_bd_ram_mem3_reg[15][26]/P0001 ,
		_w11932_,
		_w11973_,
		_w14560_
	);
	LUT3 #(
		.INIT('h80)
	) name4048 (
		\wishbone_bd_ram_mem3_reg[247][26]/P0001 ,
		_w11952_,
		_w11975_,
		_w14561_
	);
	LUT4 #(
		.INIT('h0001)
	) name4049 (
		_w14558_,
		_w14559_,
		_w14560_,
		_w14561_,
		_w14562_
	);
	LUT3 #(
		.INIT('h80)
	) name4050 (
		\wishbone_bd_ram_mem3_reg[125][26]/P0001 ,
		_w11966_,
		_w12012_,
		_w14563_
	);
	LUT3 #(
		.INIT('h80)
	) name4051 (
		\wishbone_bd_ram_mem3_reg[217][26]/P0001 ,
		_w11968_,
		_w11984_,
		_w14564_
	);
	LUT3 #(
		.INIT('h80)
	) name4052 (
		\wishbone_bd_ram_mem3_reg[215][26]/P0001 ,
		_w11975_,
		_w11984_,
		_w14565_
	);
	LUT3 #(
		.INIT('h80)
	) name4053 (
		\wishbone_bd_ram_mem3_reg[65][26]/P0001 ,
		_w11949_,
		_w11977_,
		_w14566_
	);
	LUT4 #(
		.INIT('h0001)
	) name4054 (
		_w14563_,
		_w14564_,
		_w14565_,
		_w14566_,
		_w14567_
	);
	LUT3 #(
		.INIT('h80)
	) name4055 (
		\wishbone_bd_ram_mem3_reg[67][26]/P0001 ,
		_w11938_,
		_w11949_,
		_w14568_
	);
	LUT3 #(
		.INIT('h80)
	) name4056 (
		\wishbone_bd_ram_mem3_reg[242][26]/P0001 ,
		_w11952_,
		_w11963_,
		_w14569_
	);
	LUT3 #(
		.INIT('h80)
	) name4057 (
		\wishbone_bd_ram_mem3_reg[120][26]/P0001 ,
		_w11990_,
		_w12012_,
		_w14570_
	);
	LUT3 #(
		.INIT('h80)
	) name4058 (
		\wishbone_bd_ram_mem3_reg[178][26]/P0001 ,
		_w11942_,
		_w11963_,
		_w14571_
	);
	LUT4 #(
		.INIT('h0001)
	) name4059 (
		_w14568_,
		_w14569_,
		_w14570_,
		_w14571_,
		_w14572_
	);
	LUT4 #(
		.INIT('h8000)
	) name4060 (
		_w14557_,
		_w14562_,
		_w14567_,
		_w14572_,
		_w14573_
	);
	LUT3 #(
		.INIT('h80)
	) name4061 (
		\wishbone_bd_ram_mem3_reg[212][26]/P0001 ,
		_w11929_,
		_w11984_,
		_w14574_
	);
	LUT3 #(
		.INIT('h80)
	) name4062 (
		\wishbone_bd_ram_mem3_reg[54][26]/P0001 ,
		_w11979_,
		_w11986_,
		_w14575_
	);
	LUT3 #(
		.INIT('h80)
	) name4063 (
		\wishbone_bd_ram_mem3_reg[228][26]/P0001 ,
		_w11929_,
		_w11982_,
		_w14576_
	);
	LUT3 #(
		.INIT('h80)
	) name4064 (
		\wishbone_bd_ram_mem3_reg[18][26]/P0001 ,
		_w11935_,
		_w11963_,
		_w14577_
	);
	LUT4 #(
		.INIT('h0001)
	) name4065 (
		_w14574_,
		_w14575_,
		_w14576_,
		_w14577_,
		_w14578_
	);
	LUT3 #(
		.INIT('h80)
	) name4066 (
		\wishbone_bd_ram_mem3_reg[205][26]/P0001 ,
		_w11945_,
		_w11966_,
		_w14579_
	);
	LUT3 #(
		.INIT('h80)
	) name4067 (
		\wishbone_bd_ram_mem3_reg[26][26]/P0001 ,
		_w11935_,
		_w11944_,
		_w14580_
	);
	LUT3 #(
		.INIT('h80)
	) name4068 (
		\wishbone_bd_ram_mem3_reg[229][26]/P0001 ,
		_w11933_,
		_w11982_,
		_w14581_
	);
	LUT3 #(
		.INIT('h80)
	) name4069 (
		\wishbone_bd_ram_mem3_reg[146][26]/P0001 ,
		_w11959_,
		_w11963_,
		_w14582_
	);
	LUT4 #(
		.INIT('h0001)
	) name4070 (
		_w14579_,
		_w14580_,
		_w14581_,
		_w14582_,
		_w14583_
	);
	LUT3 #(
		.INIT('h80)
	) name4071 (
		\wishbone_bd_ram_mem3_reg[182][26]/P0001 ,
		_w11942_,
		_w11986_,
		_w14584_
	);
	LUT3 #(
		.INIT('h80)
	) name4072 (
		\wishbone_bd_ram_mem3_reg[188][26]/P0001 ,
		_w11942_,
		_w11954_,
		_w14585_
	);
	LUT3 #(
		.INIT('h80)
	) name4073 (
		\wishbone_bd_ram_mem3_reg[32][26]/P0001 ,
		_w11941_,
		_w11957_,
		_w14586_
	);
	LUT3 #(
		.INIT('h80)
	) name4074 (
		\wishbone_bd_ram_mem3_reg[138][26]/P0001 ,
		_w11944_,
		_w11955_,
		_w14587_
	);
	LUT4 #(
		.INIT('h0001)
	) name4075 (
		_w14584_,
		_w14585_,
		_w14586_,
		_w14587_,
		_w14588_
	);
	LUT3 #(
		.INIT('h80)
	) name4076 (
		\wishbone_bd_ram_mem3_reg[239][26]/P0001 ,
		_w11973_,
		_w11982_,
		_w14589_
	);
	LUT3 #(
		.INIT('h80)
	) name4077 (
		\wishbone_bd_ram_mem3_reg[206][26]/P0001 ,
		_w11945_,
		_w11948_,
		_w14590_
	);
	LUT3 #(
		.INIT('h80)
	) name4078 (
		\wishbone_bd_ram_mem3_reg[56][26]/P0001 ,
		_w11979_,
		_w11990_,
		_w14591_
	);
	LUT3 #(
		.INIT('h80)
	) name4079 (
		\wishbone_bd_ram_mem3_reg[253][26]/P0001 ,
		_w11952_,
		_w11966_,
		_w14592_
	);
	LUT4 #(
		.INIT('h0001)
	) name4080 (
		_w14589_,
		_w14590_,
		_w14591_,
		_w14592_,
		_w14593_
	);
	LUT4 #(
		.INIT('h8000)
	) name4081 (
		_w14578_,
		_w14583_,
		_w14588_,
		_w14593_,
		_w14594_
	);
	LUT3 #(
		.INIT('h80)
	) name4082 (
		\wishbone_bd_ram_mem3_reg[76][26]/P0001 ,
		_w11949_,
		_w11954_,
		_w14595_
	);
	LUT3 #(
		.INIT('h80)
	) name4083 (
		\wishbone_bd_ram_mem3_reg[157][26]/P0001 ,
		_w11959_,
		_w11966_,
		_w14596_
	);
	LUT3 #(
		.INIT('h80)
	) name4084 (
		\wishbone_bd_ram_mem3_reg[145][26]/P0001 ,
		_w11959_,
		_w11977_,
		_w14597_
	);
	LUT3 #(
		.INIT('h80)
	) name4085 (
		\wishbone_bd_ram_mem3_reg[104][26]/P0001 ,
		_w11965_,
		_w11990_,
		_w14598_
	);
	LUT4 #(
		.INIT('h0001)
	) name4086 (
		_w14595_,
		_w14596_,
		_w14597_,
		_w14598_,
		_w14599_
	);
	LUT3 #(
		.INIT('h80)
	) name4087 (
		\wishbone_bd_ram_mem3_reg[112][26]/P0001 ,
		_w11941_,
		_w12012_,
		_w14600_
	);
	LUT3 #(
		.INIT('h80)
	) name4088 (
		\wishbone_bd_ram_mem3_reg[108][26]/P0001 ,
		_w11954_,
		_w11965_,
		_w14601_
	);
	LUT3 #(
		.INIT('h80)
	) name4089 (
		\wishbone_bd_ram_mem3_reg[135][26]/P0001 ,
		_w11955_,
		_w11975_,
		_w14602_
	);
	LUT3 #(
		.INIT('h80)
	) name4090 (
		\wishbone_bd_ram_mem3_reg[12][26]/P0001 ,
		_w11932_,
		_w11954_,
		_w14603_
	);
	LUT4 #(
		.INIT('h0001)
	) name4091 (
		_w14600_,
		_w14601_,
		_w14602_,
		_w14603_,
		_w14604_
	);
	LUT3 #(
		.INIT('h80)
	) name4092 (
		\wishbone_bd_ram_mem3_reg[10][26]/P0001 ,
		_w11932_,
		_w11944_,
		_w14605_
	);
	LUT3 #(
		.INIT('h80)
	) name4093 (
		\wishbone_bd_ram_mem3_reg[29][26]/P0001 ,
		_w11935_,
		_w11966_,
		_w14606_
	);
	LUT3 #(
		.INIT('h80)
	) name4094 (
		\wishbone_bd_ram_mem3_reg[87][26]/P0001 ,
		_w11972_,
		_w11975_,
		_w14607_
	);
	LUT3 #(
		.INIT('h80)
	) name4095 (
		\wishbone_bd_ram_mem3_reg[141][26]/P0001 ,
		_w11955_,
		_w11966_,
		_w14608_
	);
	LUT4 #(
		.INIT('h0001)
	) name4096 (
		_w14605_,
		_w14606_,
		_w14607_,
		_w14608_,
		_w14609_
	);
	LUT3 #(
		.INIT('h80)
	) name4097 (
		\wishbone_bd_ram_mem3_reg[11][26]/P0001 ,
		_w11932_,
		_w11936_,
		_w14610_
	);
	LUT3 #(
		.INIT('h80)
	) name4098 (
		\wishbone_bd_ram_mem3_reg[41][26]/P0001 ,
		_w11957_,
		_w11968_,
		_w14611_
	);
	LUT3 #(
		.INIT('h80)
	) name4099 (
		\wishbone_bd_ram_mem3_reg[40][26]/P0001 ,
		_w11957_,
		_w11990_,
		_w14612_
	);
	LUT3 #(
		.INIT('h80)
	) name4100 (
		\wishbone_bd_ram_mem3_reg[151][26]/P0001 ,
		_w11959_,
		_w11975_,
		_w14613_
	);
	LUT4 #(
		.INIT('h0001)
	) name4101 (
		_w14610_,
		_w14611_,
		_w14612_,
		_w14613_,
		_w14614_
	);
	LUT4 #(
		.INIT('h8000)
	) name4102 (
		_w14599_,
		_w14604_,
		_w14609_,
		_w14614_,
		_w14615_
	);
	LUT4 #(
		.INIT('h8000)
	) name4103 (
		_w14552_,
		_w14573_,
		_w14594_,
		_w14615_,
		_w14616_
	);
	LUT3 #(
		.INIT('h80)
	) name4104 (
		\wishbone_bd_ram_mem3_reg[16][26]/P0001 ,
		_w11935_,
		_w11941_,
		_w14617_
	);
	LUT3 #(
		.INIT('h80)
	) name4105 (
		\wishbone_bd_ram_mem3_reg[81][26]/P0001 ,
		_w11972_,
		_w11977_,
		_w14618_
	);
	LUT3 #(
		.INIT('h80)
	) name4106 (
		\wishbone_bd_ram_mem3_reg[140][26]/P0001 ,
		_w11954_,
		_w11955_,
		_w14619_
	);
	LUT3 #(
		.INIT('h80)
	) name4107 (
		\wishbone_bd_ram_mem3_reg[98][26]/P0001 ,
		_w11963_,
		_w11965_,
		_w14620_
	);
	LUT4 #(
		.INIT('h0001)
	) name4108 (
		_w14617_,
		_w14618_,
		_w14619_,
		_w14620_,
		_w14621_
	);
	LUT3 #(
		.INIT('h80)
	) name4109 (
		\wishbone_bd_ram_mem3_reg[231][26]/P0001 ,
		_w11975_,
		_w11982_,
		_w14622_
	);
	LUT3 #(
		.INIT('h80)
	) name4110 (
		\wishbone_bd_ram_mem3_reg[176][26]/P0001 ,
		_w11941_,
		_w11942_,
		_w14623_
	);
	LUT3 #(
		.INIT('h80)
	) name4111 (
		\wishbone_bd_ram_mem3_reg[50][26]/P0001 ,
		_w11963_,
		_w11979_,
		_w14624_
	);
	LUT3 #(
		.INIT('h80)
	) name4112 (
		\wishbone_bd_ram_mem3_reg[153][26]/P0001 ,
		_w11959_,
		_w11968_,
		_w14625_
	);
	LUT4 #(
		.INIT('h0001)
	) name4113 (
		_w14622_,
		_w14623_,
		_w14624_,
		_w14625_,
		_w14626_
	);
	LUT3 #(
		.INIT('h80)
	) name4114 (
		\wishbone_bd_ram_mem3_reg[105][26]/P0001 ,
		_w11965_,
		_w11968_,
		_w14627_
	);
	LUT3 #(
		.INIT('h80)
	) name4115 (
		\wishbone_bd_ram_mem3_reg[92][26]/P0001 ,
		_w11954_,
		_w11972_,
		_w14628_
	);
	LUT3 #(
		.INIT('h80)
	) name4116 (
		\wishbone_bd_ram_mem3_reg[193][26]/P0001 ,
		_w11945_,
		_w11977_,
		_w14629_
	);
	LUT3 #(
		.INIT('h80)
	) name4117 (
		\wishbone_bd_ram_mem3_reg[203][26]/P0001 ,
		_w11936_,
		_w11945_,
		_w14630_
	);
	LUT4 #(
		.INIT('h0001)
	) name4118 (
		_w14627_,
		_w14628_,
		_w14629_,
		_w14630_,
		_w14631_
	);
	LUT3 #(
		.INIT('h80)
	) name4119 (
		\wishbone_bd_ram_mem3_reg[133][26]/P0001 ,
		_w11933_,
		_w11955_,
		_w14632_
	);
	LUT3 #(
		.INIT('h80)
	) name4120 (
		\wishbone_bd_ram_mem3_reg[1][26]/P0001 ,
		_w11932_,
		_w11977_,
		_w14633_
	);
	LUT3 #(
		.INIT('h80)
	) name4121 (
		\wishbone_bd_ram_mem3_reg[223][26]/P0001 ,
		_w11973_,
		_w11984_,
		_w14634_
	);
	LUT3 #(
		.INIT('h80)
	) name4122 (
		\wishbone_bd_ram_mem3_reg[137][26]/P0001 ,
		_w11955_,
		_w11968_,
		_w14635_
	);
	LUT4 #(
		.INIT('h0001)
	) name4123 (
		_w14632_,
		_w14633_,
		_w14634_,
		_w14635_,
		_w14636_
	);
	LUT4 #(
		.INIT('h8000)
	) name4124 (
		_w14621_,
		_w14626_,
		_w14631_,
		_w14636_,
		_w14637_
	);
	LUT3 #(
		.INIT('h80)
	) name4125 (
		\wishbone_bd_ram_mem3_reg[47][26]/P0001 ,
		_w11957_,
		_w11973_,
		_w14638_
	);
	LUT3 #(
		.INIT('h80)
	) name4126 (
		\wishbone_bd_ram_mem3_reg[113][26]/P0001 ,
		_w11977_,
		_w12012_,
		_w14639_
	);
	LUT3 #(
		.INIT('h80)
	) name4127 (
		\wishbone_bd_ram_mem3_reg[131][26]/P0001 ,
		_w11938_,
		_w11955_,
		_w14640_
	);
	LUT3 #(
		.INIT('h80)
	) name4128 (
		\wishbone_bd_ram_mem3_reg[19][26]/P0001 ,
		_w11935_,
		_w11938_,
		_w14641_
	);
	LUT4 #(
		.INIT('h0001)
	) name4129 (
		_w14638_,
		_w14639_,
		_w14640_,
		_w14641_,
		_w14642_
	);
	LUT3 #(
		.INIT('h80)
	) name4130 (
		\wishbone_bd_ram_mem3_reg[89][26]/P0001 ,
		_w11968_,
		_w11972_,
		_w14643_
	);
	LUT3 #(
		.INIT('h80)
	) name4131 (
		\wishbone_bd_ram_mem3_reg[77][26]/P0001 ,
		_w11949_,
		_w11966_,
		_w14644_
	);
	LUT3 #(
		.INIT('h80)
	) name4132 (
		\wishbone_bd_ram_mem3_reg[166][26]/P0001 ,
		_w11930_,
		_w11986_,
		_w14645_
	);
	LUT3 #(
		.INIT('h80)
	) name4133 (
		\wishbone_bd_ram_mem3_reg[107][26]/P0001 ,
		_w11936_,
		_w11965_,
		_w14646_
	);
	LUT4 #(
		.INIT('h0001)
	) name4134 (
		_w14643_,
		_w14644_,
		_w14645_,
		_w14646_,
		_w14647_
	);
	LUT3 #(
		.INIT('h80)
	) name4135 (
		\wishbone_bd_ram_mem3_reg[43][26]/P0001 ,
		_w11936_,
		_w11957_,
		_w14648_
	);
	LUT3 #(
		.INIT('h80)
	) name4136 (
		\wishbone_bd_ram_mem3_reg[132][26]/P0001 ,
		_w11929_,
		_w11955_,
		_w14649_
	);
	LUT3 #(
		.INIT('h80)
	) name4137 (
		\wishbone_bd_ram_mem3_reg[62][26]/P0001 ,
		_w11948_,
		_w11979_,
		_w14650_
	);
	LUT3 #(
		.INIT('h80)
	) name4138 (
		\wishbone_bd_ram_mem3_reg[48][26]/P0001 ,
		_w11941_,
		_w11979_,
		_w14651_
	);
	LUT4 #(
		.INIT('h0001)
	) name4139 (
		_w14648_,
		_w14649_,
		_w14650_,
		_w14651_,
		_w14652_
	);
	LUT3 #(
		.INIT('h80)
	) name4140 (
		\wishbone_bd_ram_mem3_reg[102][26]/P0001 ,
		_w11965_,
		_w11986_,
		_w14653_
	);
	LUT3 #(
		.INIT('h80)
	) name4141 (
		\wishbone_bd_ram_mem3_reg[233][26]/P0001 ,
		_w11968_,
		_w11982_,
		_w14654_
	);
	LUT3 #(
		.INIT('h80)
	) name4142 (
		\wishbone_bd_ram_mem3_reg[255][26]/P0001 ,
		_w11952_,
		_w11973_,
		_w14655_
	);
	LUT3 #(
		.INIT('h80)
	) name4143 (
		\wishbone_bd_ram_mem3_reg[155][26]/P0001 ,
		_w11936_,
		_w11959_,
		_w14656_
	);
	LUT4 #(
		.INIT('h0001)
	) name4144 (
		_w14653_,
		_w14654_,
		_w14655_,
		_w14656_,
		_w14657_
	);
	LUT4 #(
		.INIT('h8000)
	) name4145 (
		_w14642_,
		_w14647_,
		_w14652_,
		_w14657_,
		_w14658_
	);
	LUT3 #(
		.INIT('h80)
	) name4146 (
		\wishbone_bd_ram_mem3_reg[250][26]/P0001 ,
		_w11944_,
		_w11952_,
		_w14659_
	);
	LUT3 #(
		.INIT('h80)
	) name4147 (
		\wishbone_bd_ram_mem3_reg[124][26]/P0001 ,
		_w11954_,
		_w12012_,
		_w14660_
	);
	LUT3 #(
		.INIT('h80)
	) name4148 (
		\wishbone_bd_ram_mem3_reg[78][26]/P0001 ,
		_w11948_,
		_w11949_,
		_w14661_
	);
	LUT3 #(
		.INIT('h80)
	) name4149 (
		\wishbone_bd_ram_mem3_reg[191][26]/P0001 ,
		_w11942_,
		_w11973_,
		_w14662_
	);
	LUT4 #(
		.INIT('h0001)
	) name4150 (
		_w14659_,
		_w14660_,
		_w14661_,
		_w14662_,
		_w14663_
	);
	LUT3 #(
		.INIT('h80)
	) name4151 (
		\wishbone_bd_ram_mem3_reg[192][26]/P0001 ,
		_w11941_,
		_w11945_,
		_w14664_
	);
	LUT3 #(
		.INIT('h80)
	) name4152 (
		\wishbone_bd_ram_mem3_reg[225][26]/P0001 ,
		_w11977_,
		_w11982_,
		_w14665_
	);
	LUT3 #(
		.INIT('h80)
	) name4153 (
		\wishbone_bd_ram_mem3_reg[88][26]/P0001 ,
		_w11972_,
		_w11990_,
		_w14666_
	);
	LUT3 #(
		.INIT('h80)
	) name4154 (
		\wishbone_bd_ram_mem3_reg[148][26]/P0001 ,
		_w11929_,
		_w11959_,
		_w14667_
	);
	LUT4 #(
		.INIT('h0001)
	) name4155 (
		_w14664_,
		_w14665_,
		_w14666_,
		_w14667_,
		_w14668_
	);
	LUT3 #(
		.INIT('h80)
	) name4156 (
		\wishbone_bd_ram_mem3_reg[227][26]/P0001 ,
		_w11938_,
		_w11982_,
		_w14669_
	);
	LUT3 #(
		.INIT('h80)
	) name4157 (
		\wishbone_bd_ram_mem3_reg[180][26]/P0001 ,
		_w11929_,
		_w11942_,
		_w14670_
	);
	LUT3 #(
		.INIT('h80)
	) name4158 (
		\wishbone_bd_ram_mem3_reg[202][26]/P0001 ,
		_w11944_,
		_w11945_,
		_w14671_
	);
	LUT3 #(
		.INIT('h80)
	) name4159 (
		\wishbone_bd_ram_mem3_reg[200][26]/P0001 ,
		_w11945_,
		_w11990_,
		_w14672_
	);
	LUT4 #(
		.INIT('h0001)
	) name4160 (
		_w14669_,
		_w14670_,
		_w14671_,
		_w14672_,
		_w14673_
	);
	LUT3 #(
		.INIT('h80)
	) name4161 (
		\wishbone_bd_ram_mem3_reg[171][26]/P0001 ,
		_w11930_,
		_w11936_,
		_w14674_
	);
	LUT3 #(
		.INIT('h80)
	) name4162 (
		\wishbone_bd_ram_mem3_reg[214][26]/P0001 ,
		_w11984_,
		_w11986_,
		_w14675_
	);
	LUT3 #(
		.INIT('h80)
	) name4163 (
		\wishbone_bd_ram_mem3_reg[93][26]/P0001 ,
		_w11966_,
		_w11972_,
		_w14676_
	);
	LUT3 #(
		.INIT('h80)
	) name4164 (
		\wishbone_bd_ram_mem3_reg[152][26]/P0001 ,
		_w11959_,
		_w11990_,
		_w14677_
	);
	LUT4 #(
		.INIT('h0001)
	) name4165 (
		_w14674_,
		_w14675_,
		_w14676_,
		_w14677_,
		_w14678_
	);
	LUT4 #(
		.INIT('h8000)
	) name4166 (
		_w14663_,
		_w14668_,
		_w14673_,
		_w14678_,
		_w14679_
	);
	LUT3 #(
		.INIT('h80)
	) name4167 (
		\wishbone_bd_ram_mem3_reg[60][26]/P0001 ,
		_w11954_,
		_w11979_,
		_w14680_
	);
	LUT3 #(
		.INIT('h80)
	) name4168 (
		\wishbone_bd_ram_mem3_reg[100][26]/P0001 ,
		_w11929_,
		_w11965_,
		_w14681_
	);
	LUT3 #(
		.INIT('h80)
	) name4169 (
		\wishbone_bd_ram_mem3_reg[83][26]/P0001 ,
		_w11938_,
		_w11972_,
		_w14682_
	);
	LUT3 #(
		.INIT('h80)
	) name4170 (
		\wishbone_bd_ram_mem3_reg[169][26]/P0001 ,
		_w11930_,
		_w11968_,
		_w14683_
	);
	LUT4 #(
		.INIT('h0001)
	) name4171 (
		_w14680_,
		_w14681_,
		_w14682_,
		_w14683_,
		_w14684_
	);
	LUT3 #(
		.INIT('h80)
	) name4172 (
		\wishbone_bd_ram_mem3_reg[136][26]/P0001 ,
		_w11955_,
		_w11990_,
		_w14685_
	);
	LUT3 #(
		.INIT('h80)
	) name4173 (
		\wishbone_bd_ram_mem3_reg[216][26]/P0001 ,
		_w11984_,
		_w11990_,
		_w14686_
	);
	LUT3 #(
		.INIT('h80)
	) name4174 (
		\wishbone_bd_ram_mem3_reg[97][26]/P0001 ,
		_w11965_,
		_w11977_,
		_w14687_
	);
	LUT3 #(
		.INIT('h80)
	) name4175 (
		\wishbone_bd_ram_mem3_reg[53][26]/P0001 ,
		_w11933_,
		_w11979_,
		_w14688_
	);
	LUT4 #(
		.INIT('h0001)
	) name4176 (
		_w14685_,
		_w14686_,
		_w14687_,
		_w14688_,
		_w14689_
	);
	LUT3 #(
		.INIT('h80)
	) name4177 (
		\wishbone_bd_ram_mem3_reg[220][26]/P0001 ,
		_w11954_,
		_w11984_,
		_w14690_
	);
	LUT3 #(
		.INIT('h80)
	) name4178 (
		\wishbone_bd_ram_mem3_reg[82][26]/P0001 ,
		_w11963_,
		_w11972_,
		_w14691_
	);
	LUT3 #(
		.INIT('h80)
	) name4179 (
		\wishbone_bd_ram_mem3_reg[196][26]/P0001 ,
		_w11929_,
		_w11945_,
		_w14692_
	);
	LUT3 #(
		.INIT('h80)
	) name4180 (
		\wishbone_bd_ram_mem3_reg[226][26]/P0001 ,
		_w11963_,
		_w11982_,
		_w14693_
	);
	LUT4 #(
		.INIT('h0001)
	) name4181 (
		_w14690_,
		_w14691_,
		_w14692_,
		_w14693_,
		_w14694_
	);
	LUT3 #(
		.INIT('h80)
	) name4182 (
		\wishbone_bd_ram_mem3_reg[114][26]/P0001 ,
		_w11963_,
		_w12012_,
		_w14695_
	);
	LUT3 #(
		.INIT('h80)
	) name4183 (
		\wishbone_bd_ram_mem3_reg[251][26]/P0001 ,
		_w11936_,
		_w11952_,
		_w14696_
	);
	LUT3 #(
		.INIT('h80)
	) name4184 (
		\wishbone_bd_ram_mem3_reg[3][26]/P0001 ,
		_w11932_,
		_w11938_,
		_w14697_
	);
	LUT3 #(
		.INIT('h80)
	) name4185 (
		\wishbone_bd_ram_mem3_reg[49][26]/P0001 ,
		_w11977_,
		_w11979_,
		_w14698_
	);
	LUT4 #(
		.INIT('h0001)
	) name4186 (
		_w14695_,
		_w14696_,
		_w14697_,
		_w14698_,
		_w14699_
	);
	LUT4 #(
		.INIT('h8000)
	) name4187 (
		_w14684_,
		_w14689_,
		_w14694_,
		_w14699_,
		_w14700_
	);
	LUT4 #(
		.INIT('h8000)
	) name4188 (
		_w14637_,
		_w14658_,
		_w14679_,
		_w14700_,
		_w14701_
	);
	LUT3 #(
		.INIT('h80)
	) name4189 (
		\wishbone_bd_ram_mem3_reg[39][26]/P0001 ,
		_w11957_,
		_w11975_,
		_w14702_
	);
	LUT3 #(
		.INIT('h80)
	) name4190 (
		\wishbone_bd_ram_mem3_reg[244][26]/P0001 ,
		_w11929_,
		_w11952_,
		_w14703_
	);
	LUT3 #(
		.INIT('h80)
	) name4191 (
		\wishbone_bd_ram_mem3_reg[23][26]/P0001 ,
		_w11935_,
		_w11975_,
		_w14704_
	);
	LUT3 #(
		.INIT('h80)
	) name4192 (
		\wishbone_bd_ram_mem3_reg[238][26]/P0001 ,
		_w11948_,
		_w11982_,
		_w14705_
	);
	LUT4 #(
		.INIT('h0001)
	) name4193 (
		_w14702_,
		_w14703_,
		_w14704_,
		_w14705_,
		_w14706_
	);
	LUT3 #(
		.INIT('h80)
	) name4194 (
		\wishbone_bd_ram_mem3_reg[118][26]/P0001 ,
		_w11986_,
		_w12012_,
		_w14707_
	);
	LUT3 #(
		.INIT('h80)
	) name4195 (
		\wishbone_bd_ram_mem3_reg[37][26]/P0001 ,
		_w11933_,
		_w11957_,
		_w14708_
	);
	LUT3 #(
		.INIT('h80)
	) name4196 (
		\wishbone_bd_ram_mem3_reg[190][26]/P0001 ,
		_w11942_,
		_w11948_,
		_w14709_
	);
	LUT3 #(
		.INIT('h80)
	) name4197 (
		\wishbone_bd_ram_mem3_reg[210][26]/P0001 ,
		_w11963_,
		_w11984_,
		_w14710_
	);
	LUT4 #(
		.INIT('h0001)
	) name4198 (
		_w14707_,
		_w14708_,
		_w14709_,
		_w14710_,
		_w14711_
	);
	LUT3 #(
		.INIT('h80)
	) name4199 (
		\wishbone_bd_ram_mem3_reg[130][26]/P0001 ,
		_w11955_,
		_w11963_,
		_w14712_
	);
	LUT3 #(
		.INIT('h80)
	) name4200 (
		\wishbone_bd_ram_mem3_reg[13][26]/P0001 ,
		_w11932_,
		_w11966_,
		_w14713_
	);
	LUT3 #(
		.INIT('h80)
	) name4201 (
		\wishbone_bd_ram_mem3_reg[224][26]/P0001 ,
		_w11941_,
		_w11982_,
		_w14714_
	);
	LUT3 #(
		.INIT('h80)
	) name4202 (
		\wishbone_bd_ram_mem3_reg[117][26]/P0001 ,
		_w11933_,
		_w12012_,
		_w14715_
	);
	LUT4 #(
		.INIT('h0001)
	) name4203 (
		_w14712_,
		_w14713_,
		_w14714_,
		_w14715_,
		_w14716_
	);
	LUT3 #(
		.INIT('h80)
	) name4204 (
		\wishbone_bd_ram_mem3_reg[61][26]/P0001 ,
		_w11966_,
		_w11979_,
		_w14717_
	);
	LUT3 #(
		.INIT('h80)
	) name4205 (
		\wishbone_bd_ram_mem3_reg[52][26]/P0001 ,
		_w11929_,
		_w11979_,
		_w14718_
	);
	LUT3 #(
		.INIT('h80)
	) name4206 (
		\wishbone_bd_ram_mem3_reg[162][26]/P0001 ,
		_w11930_,
		_w11963_,
		_w14719_
	);
	LUT3 #(
		.INIT('h80)
	) name4207 (
		\wishbone_bd_ram_mem3_reg[109][26]/P0001 ,
		_w11965_,
		_w11966_,
		_w14720_
	);
	LUT4 #(
		.INIT('h0001)
	) name4208 (
		_w14717_,
		_w14718_,
		_w14719_,
		_w14720_,
		_w14721_
	);
	LUT4 #(
		.INIT('h8000)
	) name4209 (
		_w14706_,
		_w14711_,
		_w14716_,
		_w14721_,
		_w14722_
	);
	LUT3 #(
		.INIT('h80)
	) name4210 (
		\wishbone_bd_ram_mem3_reg[241][26]/P0001 ,
		_w11952_,
		_w11977_,
		_w14723_
	);
	LUT3 #(
		.INIT('h80)
	) name4211 (
		\wishbone_bd_ram_mem3_reg[42][26]/P0001 ,
		_w11944_,
		_w11957_,
		_w14724_
	);
	LUT3 #(
		.INIT('h80)
	) name4212 (
		\wishbone_bd_ram_mem3_reg[17][26]/P0001 ,
		_w11935_,
		_w11977_,
		_w14725_
	);
	LUT3 #(
		.INIT('h80)
	) name4213 (
		\wishbone_bd_ram_mem3_reg[38][26]/P0001 ,
		_w11957_,
		_w11986_,
		_w14726_
	);
	LUT4 #(
		.INIT('h0001)
	) name4214 (
		_w14723_,
		_w14724_,
		_w14725_,
		_w14726_,
		_w14727_
	);
	LUT3 #(
		.INIT('h80)
	) name4215 (
		\wishbone_bd_ram_mem3_reg[219][26]/P0001 ,
		_w11936_,
		_w11984_,
		_w14728_
	);
	LUT3 #(
		.INIT('h80)
	) name4216 (
		\wishbone_bd_ram_mem3_reg[45][26]/P0001 ,
		_w11957_,
		_w11966_,
		_w14729_
	);
	LUT3 #(
		.INIT('h80)
	) name4217 (
		\wishbone_bd_ram_mem3_reg[94][26]/P0001 ,
		_w11948_,
		_w11972_,
		_w14730_
	);
	LUT3 #(
		.INIT('h80)
	) name4218 (
		\wishbone_bd_ram_mem3_reg[222][26]/P0001 ,
		_w11948_,
		_w11984_,
		_w14731_
	);
	LUT4 #(
		.INIT('h0001)
	) name4219 (
		_w14728_,
		_w14729_,
		_w14730_,
		_w14731_,
		_w14732_
	);
	LUT3 #(
		.INIT('h80)
	) name4220 (
		\wishbone_bd_ram_mem3_reg[68][26]/P0001 ,
		_w11929_,
		_w11949_,
		_w14733_
	);
	LUT3 #(
		.INIT('h80)
	) name4221 (
		\wishbone_bd_ram_mem3_reg[58][26]/P0001 ,
		_w11944_,
		_w11979_,
		_w14734_
	);
	LUT3 #(
		.INIT('h80)
	) name4222 (
		\wishbone_bd_ram_mem3_reg[91][26]/P0001 ,
		_w11936_,
		_w11972_,
		_w14735_
	);
	LUT3 #(
		.INIT('h80)
	) name4223 (
		\wishbone_bd_ram_mem3_reg[74][26]/P0001 ,
		_w11944_,
		_w11949_,
		_w14736_
	);
	LUT4 #(
		.INIT('h0001)
	) name4224 (
		_w14733_,
		_w14734_,
		_w14735_,
		_w14736_,
		_w14737_
	);
	LUT3 #(
		.INIT('h80)
	) name4225 (
		\wishbone_bd_ram_mem3_reg[167][26]/P0001 ,
		_w11930_,
		_w11975_,
		_w14738_
	);
	LUT3 #(
		.INIT('h80)
	) name4226 (
		\wishbone_bd_ram_mem3_reg[14][26]/P0001 ,
		_w11932_,
		_w11948_,
		_w14739_
	);
	LUT3 #(
		.INIT('h80)
	) name4227 (
		\wishbone_bd_ram_mem3_reg[25][26]/P0001 ,
		_w11935_,
		_w11968_,
		_w14740_
	);
	LUT3 #(
		.INIT('h80)
	) name4228 (
		\wishbone_bd_ram_mem3_reg[31][26]/P0001 ,
		_w11935_,
		_w11973_,
		_w14741_
	);
	LUT4 #(
		.INIT('h0001)
	) name4229 (
		_w14738_,
		_w14739_,
		_w14740_,
		_w14741_,
		_w14742_
	);
	LUT4 #(
		.INIT('h8000)
	) name4230 (
		_w14727_,
		_w14732_,
		_w14737_,
		_w14742_,
		_w14743_
	);
	LUT3 #(
		.INIT('h80)
	) name4231 (
		\wishbone_bd_ram_mem3_reg[213][26]/P0001 ,
		_w11933_,
		_w11984_,
		_w14744_
	);
	LUT3 #(
		.INIT('h80)
	) name4232 (
		\wishbone_bd_ram_mem3_reg[168][26]/P0001 ,
		_w11930_,
		_w11990_,
		_w14745_
	);
	LUT3 #(
		.INIT('h80)
	) name4233 (
		\wishbone_bd_ram_mem3_reg[0][26]/P0001 ,
		_w11932_,
		_w11941_,
		_w14746_
	);
	LUT3 #(
		.INIT('h80)
	) name4234 (
		\wishbone_bd_ram_mem3_reg[175][26]/P0001 ,
		_w11930_,
		_w11973_,
		_w14747_
	);
	LUT4 #(
		.INIT('h0001)
	) name4235 (
		_w14744_,
		_w14745_,
		_w14746_,
		_w14747_,
		_w14748_
	);
	LUT3 #(
		.INIT('h80)
	) name4236 (
		\wishbone_bd_ram_mem3_reg[249][26]/P0001 ,
		_w11952_,
		_w11968_,
		_w14749_
	);
	LUT3 #(
		.INIT('h80)
	) name4237 (
		\wishbone_bd_ram_mem3_reg[230][26]/P0001 ,
		_w11982_,
		_w11986_,
		_w14750_
	);
	LUT3 #(
		.INIT('h80)
	) name4238 (
		\wishbone_bd_ram_mem3_reg[163][26]/P0001 ,
		_w11930_,
		_w11938_,
		_w14751_
	);
	LUT3 #(
		.INIT('h80)
	) name4239 (
		\wishbone_bd_ram_mem3_reg[66][26]/P0001 ,
		_w11949_,
		_w11963_,
		_w14752_
	);
	LUT4 #(
		.INIT('h0001)
	) name4240 (
		_w14749_,
		_w14750_,
		_w14751_,
		_w14752_,
		_w14753_
	);
	LUT3 #(
		.INIT('h80)
	) name4241 (
		\wishbone_bd_ram_mem3_reg[2][26]/P0001 ,
		_w11932_,
		_w11963_,
		_w14754_
	);
	LUT3 #(
		.INIT('h80)
	) name4242 (
		\wishbone_bd_ram_mem3_reg[218][26]/P0001 ,
		_w11944_,
		_w11984_,
		_w14755_
	);
	LUT3 #(
		.INIT('h80)
	) name4243 (
		\wishbone_bd_ram_mem3_reg[149][26]/P0001 ,
		_w11933_,
		_w11959_,
		_w14756_
	);
	LUT3 #(
		.INIT('h80)
	) name4244 (
		\wishbone_bd_ram_mem3_reg[235][26]/P0001 ,
		_w11936_,
		_w11982_,
		_w14757_
	);
	LUT4 #(
		.INIT('h0001)
	) name4245 (
		_w14754_,
		_w14755_,
		_w14756_,
		_w14757_,
		_w14758_
	);
	LUT3 #(
		.INIT('h80)
	) name4246 (
		\wishbone_bd_ram_mem3_reg[4][26]/P0001 ,
		_w11929_,
		_w11932_,
		_w14759_
	);
	LUT3 #(
		.INIT('h80)
	) name4247 (
		\wishbone_bd_ram_mem3_reg[116][26]/P0001 ,
		_w11929_,
		_w12012_,
		_w14760_
	);
	LUT3 #(
		.INIT('h80)
	) name4248 (
		\wishbone_bd_ram_mem3_reg[150][26]/P0001 ,
		_w11959_,
		_w11986_,
		_w14761_
	);
	LUT3 #(
		.INIT('h80)
	) name4249 (
		\wishbone_bd_ram_mem3_reg[187][26]/P0001 ,
		_w11936_,
		_w11942_,
		_w14762_
	);
	LUT4 #(
		.INIT('h0001)
	) name4250 (
		_w14759_,
		_w14760_,
		_w14761_,
		_w14762_,
		_w14763_
	);
	LUT4 #(
		.INIT('h8000)
	) name4251 (
		_w14748_,
		_w14753_,
		_w14758_,
		_w14763_,
		_w14764_
	);
	LUT3 #(
		.INIT('h80)
	) name4252 (
		\wishbone_bd_ram_mem3_reg[183][26]/P0001 ,
		_w11942_,
		_w11975_,
		_w14765_
	);
	LUT3 #(
		.INIT('h80)
	) name4253 (
		\wishbone_bd_ram_mem3_reg[126][26]/P0001 ,
		_w11948_,
		_w12012_,
		_w14766_
	);
	LUT3 #(
		.INIT('h80)
	) name4254 (
		\wishbone_bd_ram_mem3_reg[142][26]/P0001 ,
		_w11948_,
		_w11955_,
		_w14767_
	);
	LUT3 #(
		.INIT('h80)
	) name4255 (
		\wishbone_bd_ram_mem3_reg[172][26]/P0001 ,
		_w11930_,
		_w11954_,
		_w14768_
	);
	LUT4 #(
		.INIT('h0001)
	) name4256 (
		_w14765_,
		_w14766_,
		_w14767_,
		_w14768_,
		_w14769_
	);
	LUT3 #(
		.INIT('h80)
	) name4257 (
		\wishbone_bd_ram_mem3_reg[174][26]/P0001 ,
		_w11930_,
		_w11948_,
		_w14770_
	);
	LUT3 #(
		.INIT('h80)
	) name4258 (
		\wishbone_bd_ram_mem3_reg[211][26]/P0001 ,
		_w11938_,
		_w11984_,
		_w14771_
	);
	LUT3 #(
		.INIT('h80)
	) name4259 (
		\wishbone_bd_ram_mem3_reg[195][26]/P0001 ,
		_w11938_,
		_w11945_,
		_w14772_
	);
	LUT3 #(
		.INIT('h80)
	) name4260 (
		\wishbone_bd_ram_mem3_reg[243][26]/P0001 ,
		_w11938_,
		_w11952_,
		_w14773_
	);
	LUT4 #(
		.INIT('h0001)
	) name4261 (
		_w14770_,
		_w14771_,
		_w14772_,
		_w14773_,
		_w14774_
	);
	LUT3 #(
		.INIT('h80)
	) name4262 (
		\wishbone_bd_ram_mem3_reg[240][26]/P0001 ,
		_w11941_,
		_w11952_,
		_w14775_
	);
	LUT3 #(
		.INIT('h80)
	) name4263 (
		\wishbone_bd_ram_mem3_reg[69][26]/P0001 ,
		_w11933_,
		_w11949_,
		_w14776_
	);
	LUT3 #(
		.INIT('h80)
	) name4264 (
		\wishbone_bd_ram_mem3_reg[154][26]/P0001 ,
		_w11944_,
		_w11959_,
		_w14777_
	);
	LUT3 #(
		.INIT('h80)
	) name4265 (
		\wishbone_bd_ram_mem3_reg[110][26]/P0001 ,
		_w11948_,
		_w11965_,
		_w14778_
	);
	LUT4 #(
		.INIT('h0001)
	) name4266 (
		_w14775_,
		_w14776_,
		_w14777_,
		_w14778_,
		_w14779_
	);
	LUT3 #(
		.INIT('h80)
	) name4267 (
		\wishbone_bd_ram_mem3_reg[73][26]/P0001 ,
		_w11949_,
		_w11968_,
		_w14780_
	);
	LUT3 #(
		.INIT('h80)
	) name4268 (
		\wishbone_bd_ram_mem3_reg[24][26]/P0001 ,
		_w11935_,
		_w11990_,
		_w14781_
	);
	LUT3 #(
		.INIT('h80)
	) name4269 (
		\wishbone_bd_ram_mem3_reg[33][26]/P0001 ,
		_w11957_,
		_w11977_,
		_w14782_
	);
	LUT3 #(
		.INIT('h80)
	) name4270 (
		\wishbone_bd_ram_mem3_reg[8][26]/P0001 ,
		_w11932_,
		_w11990_,
		_w14783_
	);
	LUT4 #(
		.INIT('h0001)
	) name4271 (
		_w14780_,
		_w14781_,
		_w14782_,
		_w14783_,
		_w14784_
	);
	LUT4 #(
		.INIT('h8000)
	) name4272 (
		_w14769_,
		_w14774_,
		_w14779_,
		_w14784_,
		_w14785_
	);
	LUT4 #(
		.INIT('h8000)
	) name4273 (
		_w14722_,
		_w14743_,
		_w14764_,
		_w14785_,
		_w14786_
	);
	LUT3 #(
		.INIT('h80)
	) name4274 (
		\wishbone_bd_ram_mem3_reg[84][26]/P0001 ,
		_w11929_,
		_w11972_,
		_w14787_
	);
	LUT3 #(
		.INIT('h80)
	) name4275 (
		\wishbone_bd_ram_mem3_reg[186][26]/P0001 ,
		_w11942_,
		_w11944_,
		_w14788_
	);
	LUT3 #(
		.INIT('h80)
	) name4276 (
		\wishbone_bd_ram_mem3_reg[99][26]/P0001 ,
		_w11938_,
		_w11965_,
		_w14789_
	);
	LUT3 #(
		.INIT('h80)
	) name4277 (
		\wishbone_bd_ram_mem3_reg[123][26]/P0001 ,
		_w11936_,
		_w12012_,
		_w14790_
	);
	LUT4 #(
		.INIT('h0001)
	) name4278 (
		_w14787_,
		_w14788_,
		_w14789_,
		_w14790_,
		_w14791_
	);
	LUT3 #(
		.INIT('h80)
	) name4279 (
		\wishbone_bd_ram_mem3_reg[96][26]/P0001 ,
		_w11941_,
		_w11965_,
		_w14792_
	);
	LUT3 #(
		.INIT('h80)
	) name4280 (
		\wishbone_bd_ram_mem3_reg[59][26]/P0001 ,
		_w11936_,
		_w11979_,
		_w14793_
	);
	LUT3 #(
		.INIT('h80)
	) name4281 (
		\wishbone_bd_ram_mem3_reg[161][26]/P0001 ,
		_w11930_,
		_w11977_,
		_w14794_
	);
	LUT3 #(
		.INIT('h80)
	) name4282 (
		\wishbone_bd_ram_mem3_reg[221][26]/P0001 ,
		_w11966_,
		_w11984_,
		_w14795_
	);
	LUT4 #(
		.INIT('h0001)
	) name4283 (
		_w14792_,
		_w14793_,
		_w14794_,
		_w14795_,
		_w14796_
	);
	LUT3 #(
		.INIT('h80)
	) name4284 (
		\wishbone_bd_ram_mem3_reg[129][26]/P0001 ,
		_w11955_,
		_w11977_,
		_w14797_
	);
	LUT3 #(
		.INIT('h80)
	) name4285 (
		\wishbone_bd_ram_mem3_reg[237][26]/P0001 ,
		_w11966_,
		_w11982_,
		_w14798_
	);
	LUT3 #(
		.INIT('h80)
	) name4286 (
		\wishbone_bd_ram_mem3_reg[22][26]/P0001 ,
		_w11935_,
		_w11986_,
		_w14799_
	);
	LUT3 #(
		.INIT('h80)
	) name4287 (
		\wishbone_bd_ram_mem3_reg[199][26]/P0001 ,
		_w11945_,
		_w11975_,
		_w14800_
	);
	LUT4 #(
		.INIT('h0001)
	) name4288 (
		_w14797_,
		_w14798_,
		_w14799_,
		_w14800_,
		_w14801_
	);
	LUT3 #(
		.INIT('h80)
	) name4289 (
		\wishbone_bd_ram_mem3_reg[70][26]/P0001 ,
		_w11949_,
		_w11986_,
		_w14802_
	);
	LUT3 #(
		.INIT('h80)
	) name4290 (
		\wishbone_bd_ram_mem3_reg[9][26]/P0001 ,
		_w11932_,
		_w11968_,
		_w14803_
	);
	LUT3 #(
		.INIT('h80)
	) name4291 (
		\wishbone_bd_ram_mem3_reg[51][26]/P0001 ,
		_w11938_,
		_w11979_,
		_w14804_
	);
	LUT3 #(
		.INIT('h80)
	) name4292 (
		\wishbone_bd_ram_mem3_reg[72][26]/P0001 ,
		_w11949_,
		_w11990_,
		_w14805_
	);
	LUT4 #(
		.INIT('h0001)
	) name4293 (
		_w14802_,
		_w14803_,
		_w14804_,
		_w14805_,
		_w14806_
	);
	LUT4 #(
		.INIT('h8000)
	) name4294 (
		_w14791_,
		_w14796_,
		_w14801_,
		_w14806_,
		_w14807_
	);
	LUT3 #(
		.INIT('h80)
	) name4295 (
		\wishbone_bd_ram_mem3_reg[27][26]/P0001 ,
		_w11935_,
		_w11936_,
		_w14808_
	);
	LUT3 #(
		.INIT('h80)
	) name4296 (
		\wishbone_bd_ram_mem3_reg[147][26]/P0001 ,
		_w11938_,
		_w11959_,
		_w14809_
	);
	LUT3 #(
		.INIT('h80)
	) name4297 (
		\wishbone_bd_ram_mem3_reg[80][26]/P0001 ,
		_w11941_,
		_w11972_,
		_w14810_
	);
	LUT3 #(
		.INIT('h80)
	) name4298 (
		\wishbone_bd_ram_mem3_reg[103][26]/P0001 ,
		_w11965_,
		_w11975_,
		_w14811_
	);
	LUT4 #(
		.INIT('h0001)
	) name4299 (
		_w14808_,
		_w14809_,
		_w14810_,
		_w14811_,
		_w14812_
	);
	LUT3 #(
		.INIT('h80)
	) name4300 (
		\wishbone_bd_ram_mem3_reg[156][26]/P0001 ,
		_w11954_,
		_w11959_,
		_w14813_
	);
	LUT3 #(
		.INIT('h80)
	) name4301 (
		\wishbone_bd_ram_mem3_reg[208][26]/P0001 ,
		_w11941_,
		_w11984_,
		_w14814_
	);
	LUT3 #(
		.INIT('h80)
	) name4302 (
		\wishbone_bd_ram_mem3_reg[28][26]/P0001 ,
		_w11935_,
		_w11954_,
		_w14815_
	);
	LUT3 #(
		.INIT('h80)
	) name4303 (
		\wishbone_bd_ram_mem3_reg[7][26]/P0001 ,
		_w11932_,
		_w11975_,
		_w14816_
	);
	LUT4 #(
		.INIT('h0001)
	) name4304 (
		_w14813_,
		_w14814_,
		_w14815_,
		_w14816_,
		_w14817_
	);
	LUT3 #(
		.INIT('h80)
	) name4305 (
		\wishbone_bd_ram_mem3_reg[177][26]/P0001 ,
		_w11942_,
		_w11977_,
		_w14818_
	);
	LUT3 #(
		.INIT('h80)
	) name4306 (
		\wishbone_bd_ram_mem3_reg[139][26]/P0001 ,
		_w11936_,
		_w11955_,
		_w14819_
	);
	LUT3 #(
		.INIT('h80)
	) name4307 (
		\wishbone_bd_ram_mem3_reg[165][26]/P0001 ,
		_w11930_,
		_w11933_,
		_w14820_
	);
	LUT3 #(
		.INIT('h80)
	) name4308 (
		\wishbone_bd_ram_mem3_reg[128][26]/P0001 ,
		_w11941_,
		_w11955_,
		_w14821_
	);
	LUT4 #(
		.INIT('h0001)
	) name4309 (
		_w14818_,
		_w14819_,
		_w14820_,
		_w14821_,
		_w14822_
	);
	LUT3 #(
		.INIT('h80)
	) name4310 (
		\wishbone_bd_ram_mem3_reg[30][26]/P0001 ,
		_w11935_,
		_w11948_,
		_w14823_
	);
	LUT3 #(
		.INIT('h80)
	) name4311 (
		\wishbone_bd_ram_mem3_reg[20][26]/P0001 ,
		_w11929_,
		_w11935_,
		_w14824_
	);
	LUT3 #(
		.INIT('h80)
	) name4312 (
		\wishbone_bd_ram_mem3_reg[252][26]/P0001 ,
		_w11952_,
		_w11954_,
		_w14825_
	);
	LUT3 #(
		.INIT('h80)
	) name4313 (
		\wishbone_bd_ram_mem3_reg[71][26]/P0001 ,
		_w11949_,
		_w11975_,
		_w14826_
	);
	LUT4 #(
		.INIT('h0001)
	) name4314 (
		_w14823_,
		_w14824_,
		_w14825_,
		_w14826_,
		_w14827_
	);
	LUT4 #(
		.INIT('h8000)
	) name4315 (
		_w14812_,
		_w14817_,
		_w14822_,
		_w14827_,
		_w14828_
	);
	LUT3 #(
		.INIT('h80)
	) name4316 (
		\wishbone_bd_ram_mem3_reg[236][26]/P0001 ,
		_w11954_,
		_w11982_,
		_w14829_
	);
	LUT3 #(
		.INIT('h80)
	) name4317 (
		\wishbone_bd_ram_mem3_reg[5][26]/P0001 ,
		_w11932_,
		_w11933_,
		_w14830_
	);
	LUT3 #(
		.INIT('h80)
	) name4318 (
		\wishbone_bd_ram_mem3_reg[106][26]/P0001 ,
		_w11944_,
		_w11965_,
		_w14831_
	);
	LUT3 #(
		.INIT('h80)
	) name4319 (
		\wishbone_bd_ram_mem3_reg[184][26]/P0001 ,
		_w11942_,
		_w11990_,
		_w14832_
	);
	LUT4 #(
		.INIT('h0001)
	) name4320 (
		_w14829_,
		_w14830_,
		_w14831_,
		_w14832_,
		_w14833_
	);
	LUT3 #(
		.INIT('h80)
	) name4321 (
		\wishbone_bd_ram_mem3_reg[79][26]/P0001 ,
		_w11949_,
		_w11973_,
		_w14834_
	);
	LUT3 #(
		.INIT('h80)
	) name4322 (
		\wishbone_bd_ram_mem3_reg[232][26]/P0001 ,
		_w11982_,
		_w11990_,
		_w14835_
	);
	LUT3 #(
		.INIT('h80)
	) name4323 (
		\wishbone_bd_ram_mem3_reg[122][26]/P0001 ,
		_w11944_,
		_w12012_,
		_w14836_
	);
	LUT3 #(
		.INIT('h80)
	) name4324 (
		\wishbone_bd_ram_mem3_reg[197][26]/P0001 ,
		_w11933_,
		_w11945_,
		_w14837_
	);
	LUT4 #(
		.INIT('h0001)
	) name4325 (
		_w14834_,
		_w14835_,
		_w14836_,
		_w14837_,
		_w14838_
	);
	LUT3 #(
		.INIT('h80)
	) name4326 (
		\wishbone_bd_ram_mem3_reg[85][26]/P0001 ,
		_w11933_,
		_w11972_,
		_w14839_
	);
	LUT3 #(
		.INIT('h80)
	) name4327 (
		\wishbone_bd_ram_mem3_reg[46][26]/P0001 ,
		_w11948_,
		_w11957_,
		_w14840_
	);
	LUT3 #(
		.INIT('h80)
	) name4328 (
		\wishbone_bd_ram_mem3_reg[44][26]/P0001 ,
		_w11954_,
		_w11957_,
		_w14841_
	);
	LUT3 #(
		.INIT('h80)
	) name4329 (
		\wishbone_bd_ram_mem3_reg[35][26]/P0001 ,
		_w11938_,
		_w11957_,
		_w14842_
	);
	LUT4 #(
		.INIT('h0001)
	) name4330 (
		_w14839_,
		_w14840_,
		_w14841_,
		_w14842_,
		_w14843_
	);
	LUT3 #(
		.INIT('h80)
	) name4331 (
		\wishbone_bd_ram_mem3_reg[245][26]/P0001 ,
		_w11933_,
		_w11952_,
		_w14844_
	);
	LUT3 #(
		.INIT('h80)
	) name4332 (
		\wishbone_bd_ram_mem3_reg[164][26]/P0001 ,
		_w11929_,
		_w11930_,
		_w14845_
	);
	LUT3 #(
		.INIT('h80)
	) name4333 (
		\wishbone_bd_ram_mem3_reg[246][26]/P0001 ,
		_w11952_,
		_w11986_,
		_w14846_
	);
	LUT3 #(
		.INIT('h80)
	) name4334 (
		\wishbone_bd_ram_mem3_reg[95][26]/P0001 ,
		_w11972_,
		_w11973_,
		_w14847_
	);
	LUT4 #(
		.INIT('h0001)
	) name4335 (
		_w14844_,
		_w14845_,
		_w14846_,
		_w14847_,
		_w14848_
	);
	LUT4 #(
		.INIT('h8000)
	) name4336 (
		_w14833_,
		_w14838_,
		_w14843_,
		_w14848_,
		_w14849_
	);
	LUT3 #(
		.INIT('h80)
	) name4337 (
		\wishbone_bd_ram_mem3_reg[34][26]/P0001 ,
		_w11957_,
		_w11963_,
		_w14850_
	);
	LUT3 #(
		.INIT('h80)
	) name4338 (
		\wishbone_bd_ram_mem3_reg[134][26]/P0001 ,
		_w11955_,
		_w11986_,
		_w14851_
	);
	LUT3 #(
		.INIT('h80)
	) name4339 (
		\wishbone_bd_ram_mem3_reg[121][26]/P0001 ,
		_w11968_,
		_w12012_,
		_w14852_
	);
	LUT3 #(
		.INIT('h80)
	) name4340 (
		\wishbone_bd_ram_mem3_reg[21][26]/P0001 ,
		_w11933_,
		_w11935_,
		_w14853_
	);
	LUT4 #(
		.INIT('h0001)
	) name4341 (
		_w14850_,
		_w14851_,
		_w14852_,
		_w14853_,
		_w14854_
	);
	LUT3 #(
		.INIT('h80)
	) name4342 (
		\wishbone_bd_ram_mem3_reg[194][26]/P0001 ,
		_w11945_,
		_w11963_,
		_w14855_
	);
	LUT3 #(
		.INIT('h80)
	) name4343 (
		\wishbone_bd_ram_mem3_reg[179][26]/P0001 ,
		_w11938_,
		_w11942_,
		_w14856_
	);
	LUT3 #(
		.INIT('h80)
	) name4344 (
		\wishbone_bd_ram_mem3_reg[6][26]/P0001 ,
		_w11932_,
		_w11986_,
		_w14857_
	);
	LUT3 #(
		.INIT('h80)
	) name4345 (
		\wishbone_bd_ram_mem3_reg[173][26]/P0001 ,
		_w11930_,
		_w11966_,
		_w14858_
	);
	LUT4 #(
		.INIT('h0001)
	) name4346 (
		_w14855_,
		_w14856_,
		_w14857_,
		_w14858_,
		_w14859_
	);
	LUT3 #(
		.INIT('h80)
	) name4347 (
		\wishbone_bd_ram_mem3_reg[115][26]/P0001 ,
		_w11938_,
		_w12012_,
		_w14860_
	);
	LUT3 #(
		.INIT('h80)
	) name4348 (
		\wishbone_bd_ram_mem3_reg[181][26]/P0001 ,
		_w11933_,
		_w11942_,
		_w14861_
	);
	LUT3 #(
		.INIT('h80)
	) name4349 (
		\wishbone_bd_ram_mem3_reg[234][26]/P0001 ,
		_w11944_,
		_w11982_,
		_w14862_
	);
	LUT3 #(
		.INIT('h80)
	) name4350 (
		\wishbone_bd_ram_mem3_reg[158][26]/P0001 ,
		_w11948_,
		_w11959_,
		_w14863_
	);
	LUT4 #(
		.INIT('h0001)
	) name4351 (
		_w14860_,
		_w14861_,
		_w14862_,
		_w14863_,
		_w14864_
	);
	LUT3 #(
		.INIT('h80)
	) name4352 (
		\wishbone_bd_ram_mem3_reg[101][26]/P0001 ,
		_w11933_,
		_w11965_,
		_w14865_
	);
	LUT3 #(
		.INIT('h80)
	) name4353 (
		\wishbone_bd_ram_mem3_reg[198][26]/P0001 ,
		_w11945_,
		_w11986_,
		_w14866_
	);
	LUT3 #(
		.INIT('h80)
	) name4354 (
		\wishbone_bd_ram_mem3_reg[144][26]/P0001 ,
		_w11941_,
		_w11959_,
		_w14867_
	);
	LUT3 #(
		.INIT('h80)
	) name4355 (
		\wishbone_bd_ram_mem3_reg[170][26]/P0001 ,
		_w11930_,
		_w11944_,
		_w14868_
	);
	LUT4 #(
		.INIT('h0001)
	) name4356 (
		_w14865_,
		_w14866_,
		_w14867_,
		_w14868_,
		_w14869_
	);
	LUT4 #(
		.INIT('h8000)
	) name4357 (
		_w14854_,
		_w14859_,
		_w14864_,
		_w14869_,
		_w14870_
	);
	LUT4 #(
		.INIT('h8000)
	) name4358 (
		_w14807_,
		_w14828_,
		_w14849_,
		_w14870_,
		_w14871_
	);
	LUT4 #(
		.INIT('h8000)
	) name4359 (
		_w14616_,
		_w14701_,
		_w14786_,
		_w14871_,
		_w14872_
	);
	LUT4 #(
		.INIT('h040c)
	) name4360 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[10]/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		_w14873_
	);
	LUT2 #(
		.INIT('h2)
	) name4361 (
		\wishbone_TxLength_reg[10]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w14874_
	);
	LUT3 #(
		.INIT('h23)
	) name4362 (
		_w12322_,
		_w14873_,
		_w14874_,
		_w14875_
	);
	LUT4 #(
		.INIT('h8000)
	) name4363 (
		_w12304_,
		_w12307_,
		_w12309_,
		_w12310_,
		_w14876_
	);
	LUT3 #(
		.INIT('hb0)
	) name4364 (
		_w12317_,
		_w14875_,
		_w14876_,
		_w14877_
	);
	LUT4 #(
		.INIT('hef8f)
	) name4365 (
		\wishbone_TxLength_reg[1]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w12304_,
		_w12321_,
		_w14878_
	);
	LUT4 #(
		.INIT('h2232)
	) name4366 (
		\wishbone_TxLength_reg[10]/NET0131 ,
		_w12302_,
		_w12312_,
		_w14878_,
		_w14879_
	);
	LUT2 #(
		.INIT('h4)
	) name4367 (
		_w14877_,
		_w14879_,
		_w14880_
	);
	LUT3 #(
		.INIT('hf2)
	) name4368 (
		_w12303_,
		_w14872_,
		_w14880_,
		_w14881_
	);
	LUT3 #(
		.INIT('h80)
	) name4369 (
		\wishbone_bd_ram_mem3_reg[157][25]/P0001 ,
		_w11959_,
		_w11966_,
		_w14882_
	);
	LUT3 #(
		.INIT('h80)
	) name4370 (
		\wishbone_bd_ram_mem3_reg[183][25]/P0001 ,
		_w11942_,
		_w11975_,
		_w14883_
	);
	LUT3 #(
		.INIT('h80)
	) name4371 (
		\wishbone_bd_ram_mem3_reg[24][25]/P0001 ,
		_w11935_,
		_w11990_,
		_w14884_
	);
	LUT3 #(
		.INIT('h80)
	) name4372 (
		\wishbone_bd_ram_mem3_reg[51][25]/P0001 ,
		_w11938_,
		_w11979_,
		_w14885_
	);
	LUT4 #(
		.INIT('h0001)
	) name4373 (
		_w14882_,
		_w14883_,
		_w14884_,
		_w14885_,
		_w14886_
	);
	LUT3 #(
		.INIT('h80)
	) name4374 (
		\wishbone_bd_ram_mem3_reg[222][25]/P0001 ,
		_w11948_,
		_w11984_,
		_w14887_
	);
	LUT3 #(
		.INIT('h80)
	) name4375 (
		\wishbone_bd_ram_mem3_reg[172][25]/P0001 ,
		_w11930_,
		_w11954_,
		_w14888_
	);
	LUT3 #(
		.INIT('h80)
	) name4376 (
		\wishbone_bd_ram_mem3_reg[85][25]/P0001 ,
		_w11933_,
		_w11972_,
		_w14889_
	);
	LUT3 #(
		.INIT('h80)
	) name4377 (
		\wishbone_bd_ram_mem3_reg[242][25]/P0001 ,
		_w11952_,
		_w11963_,
		_w14890_
	);
	LUT4 #(
		.INIT('h0001)
	) name4378 (
		_w14887_,
		_w14888_,
		_w14889_,
		_w14890_,
		_w14891_
	);
	LUT3 #(
		.INIT('h80)
	) name4379 (
		\wishbone_bd_ram_mem3_reg[217][25]/P0001 ,
		_w11968_,
		_w11984_,
		_w14892_
	);
	LUT3 #(
		.INIT('h80)
	) name4380 (
		\wishbone_bd_ram_mem3_reg[140][25]/P0001 ,
		_w11954_,
		_w11955_,
		_w14893_
	);
	LUT3 #(
		.INIT('h80)
	) name4381 (
		\wishbone_bd_ram_mem3_reg[34][25]/P0001 ,
		_w11957_,
		_w11963_,
		_w14894_
	);
	LUT3 #(
		.INIT('h80)
	) name4382 (
		\wishbone_bd_ram_mem3_reg[93][25]/P0001 ,
		_w11966_,
		_w11972_,
		_w14895_
	);
	LUT4 #(
		.INIT('h0001)
	) name4383 (
		_w14892_,
		_w14893_,
		_w14894_,
		_w14895_,
		_w14896_
	);
	LUT3 #(
		.INIT('h80)
	) name4384 (
		\wishbone_bd_ram_mem3_reg[234][25]/P0001 ,
		_w11944_,
		_w11982_,
		_w14897_
	);
	LUT3 #(
		.INIT('h80)
	) name4385 (
		\wishbone_bd_ram_mem3_reg[105][25]/P0001 ,
		_w11965_,
		_w11968_,
		_w14898_
	);
	LUT3 #(
		.INIT('h80)
	) name4386 (
		\wishbone_bd_ram_mem3_reg[253][25]/P0001 ,
		_w11952_,
		_w11966_,
		_w14899_
	);
	LUT3 #(
		.INIT('h80)
	) name4387 (
		\wishbone_bd_ram_mem3_reg[108][25]/P0001 ,
		_w11954_,
		_w11965_,
		_w14900_
	);
	LUT4 #(
		.INIT('h0001)
	) name4388 (
		_w14897_,
		_w14898_,
		_w14899_,
		_w14900_,
		_w14901_
	);
	LUT4 #(
		.INIT('h8000)
	) name4389 (
		_w14886_,
		_w14891_,
		_w14896_,
		_w14901_,
		_w14902_
	);
	LUT3 #(
		.INIT('h80)
	) name4390 (
		\wishbone_bd_ram_mem3_reg[61][25]/P0001 ,
		_w11966_,
		_w11979_,
		_w14903_
	);
	LUT3 #(
		.INIT('h80)
	) name4391 (
		\wishbone_bd_ram_mem3_reg[98][25]/P0001 ,
		_w11963_,
		_w11965_,
		_w14904_
	);
	LUT3 #(
		.INIT('h80)
	) name4392 (
		\wishbone_bd_ram_mem3_reg[79][25]/P0001 ,
		_w11949_,
		_w11973_,
		_w14905_
	);
	LUT3 #(
		.INIT('h80)
	) name4393 (
		\wishbone_bd_ram_mem3_reg[202][25]/P0001 ,
		_w11944_,
		_w11945_,
		_w14906_
	);
	LUT4 #(
		.INIT('h0001)
	) name4394 (
		_w14903_,
		_w14904_,
		_w14905_,
		_w14906_,
		_w14907_
	);
	LUT3 #(
		.INIT('h80)
	) name4395 (
		\wishbone_bd_ram_mem3_reg[213][25]/P0001 ,
		_w11933_,
		_w11984_,
		_w14908_
	);
	LUT3 #(
		.INIT('h80)
	) name4396 (
		\wishbone_bd_ram_mem3_reg[90][25]/P0001 ,
		_w11944_,
		_w11972_,
		_w14909_
	);
	LUT3 #(
		.INIT('h80)
	) name4397 (
		\wishbone_bd_ram_mem3_reg[110][25]/P0001 ,
		_w11948_,
		_w11965_,
		_w14910_
	);
	LUT3 #(
		.INIT('h80)
	) name4398 (
		\wishbone_bd_ram_mem3_reg[243][25]/P0001 ,
		_w11938_,
		_w11952_,
		_w14911_
	);
	LUT4 #(
		.INIT('h0001)
	) name4399 (
		_w14908_,
		_w14909_,
		_w14910_,
		_w14911_,
		_w14912_
	);
	LUT3 #(
		.INIT('h80)
	) name4400 (
		\wishbone_bd_ram_mem3_reg[153][25]/P0001 ,
		_w11959_,
		_w11968_,
		_w14913_
	);
	LUT3 #(
		.INIT('h80)
	) name4401 (
		\wishbone_bd_ram_mem3_reg[94][25]/P0001 ,
		_w11948_,
		_w11972_,
		_w14914_
	);
	LUT3 #(
		.INIT('h80)
	) name4402 (
		\wishbone_bd_ram_mem3_reg[122][25]/P0001 ,
		_w11944_,
		_w12012_,
		_w14915_
	);
	LUT3 #(
		.INIT('h80)
	) name4403 (
		\wishbone_bd_ram_mem3_reg[144][25]/P0001 ,
		_w11941_,
		_w11959_,
		_w14916_
	);
	LUT4 #(
		.INIT('h0001)
	) name4404 (
		_w14913_,
		_w14914_,
		_w14915_,
		_w14916_,
		_w14917_
	);
	LUT3 #(
		.INIT('h80)
	) name4405 (
		\wishbone_bd_ram_mem3_reg[1][25]/P0001 ,
		_w11932_,
		_w11977_,
		_w14918_
	);
	LUT3 #(
		.INIT('h80)
	) name4406 (
		\wishbone_bd_ram_mem3_reg[220][25]/P0001 ,
		_w11954_,
		_w11984_,
		_w14919_
	);
	LUT3 #(
		.INIT('h80)
	) name4407 (
		\wishbone_bd_ram_mem3_reg[64][25]/P0001 ,
		_w11941_,
		_w11949_,
		_w14920_
	);
	LUT3 #(
		.INIT('h80)
	) name4408 (
		\wishbone_bd_ram_mem3_reg[190][25]/P0001 ,
		_w11942_,
		_w11948_,
		_w14921_
	);
	LUT4 #(
		.INIT('h0001)
	) name4409 (
		_w14918_,
		_w14919_,
		_w14920_,
		_w14921_,
		_w14922_
	);
	LUT4 #(
		.INIT('h8000)
	) name4410 (
		_w14907_,
		_w14912_,
		_w14917_,
		_w14922_,
		_w14923_
	);
	LUT3 #(
		.INIT('h80)
	) name4411 (
		\wishbone_bd_ram_mem3_reg[127][25]/P0001 ,
		_w11973_,
		_w12012_,
		_w14924_
	);
	LUT3 #(
		.INIT('h80)
	) name4412 (
		\wishbone_bd_ram_mem3_reg[101][25]/P0001 ,
		_w11933_,
		_w11965_,
		_w14925_
	);
	LUT3 #(
		.INIT('h80)
	) name4413 (
		\wishbone_bd_ram_mem3_reg[154][25]/P0001 ,
		_w11944_,
		_w11959_,
		_w14926_
	);
	LUT3 #(
		.INIT('h80)
	) name4414 (
		\wishbone_bd_ram_mem3_reg[50][25]/P0001 ,
		_w11963_,
		_w11979_,
		_w14927_
	);
	LUT4 #(
		.INIT('h0001)
	) name4415 (
		_w14924_,
		_w14925_,
		_w14926_,
		_w14927_,
		_w14928_
	);
	LUT3 #(
		.INIT('h80)
	) name4416 (
		\wishbone_bd_ram_mem3_reg[211][25]/P0001 ,
		_w11938_,
		_w11984_,
		_w14929_
	);
	LUT3 #(
		.INIT('h80)
	) name4417 (
		\wishbone_bd_ram_mem3_reg[149][25]/P0001 ,
		_w11933_,
		_w11959_,
		_w14930_
	);
	LUT3 #(
		.INIT('h80)
	) name4418 (
		\wishbone_bd_ram_mem3_reg[227][25]/P0001 ,
		_w11938_,
		_w11982_,
		_w14931_
	);
	LUT3 #(
		.INIT('h80)
	) name4419 (
		\wishbone_bd_ram_mem3_reg[96][25]/P0001 ,
		_w11941_,
		_w11965_,
		_w14932_
	);
	LUT4 #(
		.INIT('h0001)
	) name4420 (
		_w14929_,
		_w14930_,
		_w14931_,
		_w14932_,
		_w14933_
	);
	LUT3 #(
		.INIT('h80)
	) name4421 (
		\wishbone_bd_ram_mem3_reg[52][25]/P0001 ,
		_w11929_,
		_w11979_,
		_w14934_
	);
	LUT3 #(
		.INIT('h80)
	) name4422 (
		\wishbone_bd_ram_mem3_reg[196][25]/P0001 ,
		_w11929_,
		_w11945_,
		_w14935_
	);
	LUT3 #(
		.INIT('h80)
	) name4423 (
		\wishbone_bd_ram_mem3_reg[74][25]/P0001 ,
		_w11944_,
		_w11949_,
		_w14936_
	);
	LUT3 #(
		.INIT('h80)
	) name4424 (
		\wishbone_bd_ram_mem3_reg[112][25]/P0001 ,
		_w11941_,
		_w12012_,
		_w14937_
	);
	LUT4 #(
		.INIT('h0001)
	) name4425 (
		_w14934_,
		_w14935_,
		_w14936_,
		_w14937_,
		_w14938_
	);
	LUT3 #(
		.INIT('h80)
	) name4426 (
		\wishbone_bd_ram_mem3_reg[165][25]/P0001 ,
		_w11930_,
		_w11933_,
		_w14939_
	);
	LUT3 #(
		.INIT('h80)
	) name4427 (
		\wishbone_bd_ram_mem3_reg[252][25]/P0001 ,
		_w11952_,
		_w11954_,
		_w14940_
	);
	LUT3 #(
		.INIT('h80)
	) name4428 (
		\wishbone_bd_ram_mem3_reg[29][25]/P0001 ,
		_w11935_,
		_w11966_,
		_w14941_
	);
	LUT3 #(
		.INIT('h80)
	) name4429 (
		\wishbone_bd_ram_mem3_reg[205][25]/P0001 ,
		_w11945_,
		_w11966_,
		_w14942_
	);
	LUT4 #(
		.INIT('h0001)
	) name4430 (
		_w14939_,
		_w14940_,
		_w14941_,
		_w14942_,
		_w14943_
	);
	LUT4 #(
		.INIT('h8000)
	) name4431 (
		_w14928_,
		_w14933_,
		_w14938_,
		_w14943_,
		_w14944_
	);
	LUT3 #(
		.INIT('h80)
	) name4432 (
		\wishbone_bd_ram_mem3_reg[59][25]/P0001 ,
		_w11936_,
		_w11979_,
		_w14945_
	);
	LUT3 #(
		.INIT('h80)
	) name4433 (
		\wishbone_bd_ram_mem3_reg[128][25]/P0001 ,
		_w11941_,
		_w11955_,
		_w14946_
	);
	LUT3 #(
		.INIT('h80)
	) name4434 (
		\wishbone_bd_ram_mem3_reg[47][25]/P0001 ,
		_w11957_,
		_w11973_,
		_w14947_
	);
	LUT3 #(
		.INIT('h80)
	) name4435 (
		\wishbone_bd_ram_mem3_reg[177][25]/P0001 ,
		_w11942_,
		_w11977_,
		_w14948_
	);
	LUT4 #(
		.INIT('h0001)
	) name4436 (
		_w14945_,
		_w14946_,
		_w14947_,
		_w14948_,
		_w14949_
	);
	LUT3 #(
		.INIT('h80)
	) name4437 (
		\wishbone_bd_ram_mem3_reg[100][25]/P0001 ,
		_w11929_,
		_w11965_,
		_w14950_
	);
	LUT3 #(
		.INIT('h80)
	) name4438 (
		\wishbone_bd_ram_mem3_reg[60][25]/P0001 ,
		_w11954_,
		_w11979_,
		_w14951_
	);
	LUT3 #(
		.INIT('h80)
	) name4439 (
		\wishbone_bd_ram_mem3_reg[39][25]/P0001 ,
		_w11957_,
		_w11975_,
		_w14952_
	);
	LUT3 #(
		.INIT('h80)
	) name4440 (
		\wishbone_bd_ram_mem3_reg[166][25]/P0001 ,
		_w11930_,
		_w11986_,
		_w14953_
	);
	LUT4 #(
		.INIT('h0001)
	) name4441 (
		_w14950_,
		_w14951_,
		_w14952_,
		_w14953_,
		_w14954_
	);
	LUT3 #(
		.INIT('h80)
	) name4442 (
		\wishbone_bd_ram_mem3_reg[176][25]/P0001 ,
		_w11941_,
		_w11942_,
		_w14955_
	);
	LUT3 #(
		.INIT('h80)
	) name4443 (
		\wishbone_bd_ram_mem3_reg[3][25]/P0001 ,
		_w11932_,
		_w11938_,
		_w14956_
	);
	LUT3 #(
		.INIT('h80)
	) name4444 (
		\wishbone_bd_ram_mem3_reg[81][25]/P0001 ,
		_w11972_,
		_w11977_,
		_w14957_
	);
	LUT3 #(
		.INIT('h80)
	) name4445 (
		\wishbone_bd_ram_mem3_reg[77][25]/P0001 ,
		_w11949_,
		_w11966_,
		_w14958_
	);
	LUT4 #(
		.INIT('h0001)
	) name4446 (
		_w14955_,
		_w14956_,
		_w14957_,
		_w14958_,
		_w14959_
	);
	LUT3 #(
		.INIT('h80)
	) name4447 (
		\wishbone_bd_ram_mem3_reg[36][25]/P0001 ,
		_w11929_,
		_w11957_,
		_w14960_
	);
	LUT3 #(
		.INIT('h80)
	) name4448 (
		\wishbone_bd_ram_mem3_reg[55][25]/P0001 ,
		_w11975_,
		_w11979_,
		_w14961_
	);
	LUT3 #(
		.INIT('h80)
	) name4449 (
		\wishbone_bd_ram_mem3_reg[106][25]/P0001 ,
		_w11944_,
		_w11965_,
		_w14962_
	);
	LUT3 #(
		.INIT('h80)
	) name4450 (
		\wishbone_bd_ram_mem3_reg[143][25]/P0001 ,
		_w11955_,
		_w11973_,
		_w14963_
	);
	LUT4 #(
		.INIT('h0001)
	) name4451 (
		_w14960_,
		_w14961_,
		_w14962_,
		_w14963_,
		_w14964_
	);
	LUT4 #(
		.INIT('h8000)
	) name4452 (
		_w14949_,
		_w14954_,
		_w14959_,
		_w14964_,
		_w14965_
	);
	LUT4 #(
		.INIT('h8000)
	) name4453 (
		_w14902_,
		_w14923_,
		_w14944_,
		_w14965_,
		_w14966_
	);
	LUT3 #(
		.INIT('h80)
	) name4454 (
		\wishbone_bd_ram_mem3_reg[38][25]/P0001 ,
		_w11957_,
		_w11986_,
		_w14967_
	);
	LUT3 #(
		.INIT('h80)
	) name4455 (
		\wishbone_bd_ram_mem3_reg[229][25]/P0001 ,
		_w11933_,
		_w11982_,
		_w14968_
	);
	LUT3 #(
		.INIT('h80)
	) name4456 (
		\wishbone_bd_ram_mem3_reg[126][25]/P0001 ,
		_w11948_,
		_w12012_,
		_w14969_
	);
	LUT3 #(
		.INIT('h80)
	) name4457 (
		\wishbone_bd_ram_mem3_reg[86][25]/P0001 ,
		_w11972_,
		_w11986_,
		_w14970_
	);
	LUT4 #(
		.INIT('h0001)
	) name4458 (
		_w14967_,
		_w14968_,
		_w14969_,
		_w14970_,
		_w14971_
	);
	LUT3 #(
		.INIT('h80)
	) name4459 (
		\wishbone_bd_ram_mem3_reg[130][25]/P0001 ,
		_w11955_,
		_w11963_,
		_w14972_
	);
	LUT3 #(
		.INIT('h80)
	) name4460 (
		\wishbone_bd_ram_mem3_reg[124][25]/P0001 ,
		_w11954_,
		_w12012_,
		_w14973_
	);
	LUT3 #(
		.INIT('h80)
	) name4461 (
		\wishbone_bd_ram_mem3_reg[0][25]/P0001 ,
		_w11932_,
		_w11941_,
		_w14974_
	);
	LUT3 #(
		.INIT('h80)
	) name4462 (
		\wishbone_bd_ram_mem3_reg[5][25]/P0001 ,
		_w11932_,
		_w11933_,
		_w14975_
	);
	LUT4 #(
		.INIT('h0001)
	) name4463 (
		_w14972_,
		_w14973_,
		_w14974_,
		_w14975_,
		_w14976_
	);
	LUT3 #(
		.INIT('h80)
	) name4464 (
		\wishbone_bd_ram_mem3_reg[195][25]/P0001 ,
		_w11938_,
		_w11945_,
		_w14977_
	);
	LUT3 #(
		.INIT('h80)
	) name4465 (
		\wishbone_bd_ram_mem3_reg[251][25]/P0001 ,
		_w11936_,
		_w11952_,
		_w14978_
	);
	LUT3 #(
		.INIT('h80)
	) name4466 (
		\wishbone_bd_ram_mem3_reg[159][25]/P0001 ,
		_w11959_,
		_w11973_,
		_w14979_
	);
	LUT3 #(
		.INIT('h80)
	) name4467 (
		\wishbone_bd_ram_mem3_reg[199][25]/P0001 ,
		_w11945_,
		_w11975_,
		_w14980_
	);
	LUT4 #(
		.INIT('h0001)
	) name4468 (
		_w14977_,
		_w14978_,
		_w14979_,
		_w14980_,
		_w14981_
	);
	LUT3 #(
		.INIT('h80)
	) name4469 (
		\wishbone_bd_ram_mem3_reg[152][25]/P0001 ,
		_w11959_,
		_w11990_,
		_w14982_
	);
	LUT3 #(
		.INIT('h80)
	) name4470 (
		\wishbone_bd_ram_mem3_reg[230][25]/P0001 ,
		_w11982_,
		_w11986_,
		_w14983_
	);
	LUT3 #(
		.INIT('h80)
	) name4471 (
		\wishbone_bd_ram_mem3_reg[164][25]/P0001 ,
		_w11929_,
		_w11930_,
		_w14984_
	);
	LUT3 #(
		.INIT('h80)
	) name4472 (
		\wishbone_bd_ram_mem3_reg[109][25]/P0001 ,
		_w11965_,
		_w11966_,
		_w14985_
	);
	LUT4 #(
		.INIT('h0001)
	) name4473 (
		_w14982_,
		_w14983_,
		_w14984_,
		_w14985_,
		_w14986_
	);
	LUT4 #(
		.INIT('h8000)
	) name4474 (
		_w14971_,
		_w14976_,
		_w14981_,
		_w14986_,
		_w14987_
	);
	LUT3 #(
		.INIT('h80)
	) name4475 (
		\wishbone_bd_ram_mem3_reg[57][25]/P0001 ,
		_w11968_,
		_w11979_,
		_w14988_
	);
	LUT3 #(
		.INIT('h80)
	) name4476 (
		\wishbone_bd_ram_mem3_reg[179][25]/P0001 ,
		_w11938_,
		_w11942_,
		_w14989_
	);
	LUT3 #(
		.INIT('h80)
	) name4477 (
		\wishbone_bd_ram_mem3_reg[160][25]/P0001 ,
		_w11930_,
		_w11941_,
		_w14990_
	);
	LUT3 #(
		.INIT('h80)
	) name4478 (
		\wishbone_bd_ram_mem3_reg[169][25]/P0001 ,
		_w11930_,
		_w11968_,
		_w14991_
	);
	LUT4 #(
		.INIT('h0001)
	) name4479 (
		_w14988_,
		_w14989_,
		_w14990_,
		_w14991_,
		_w14992_
	);
	LUT3 #(
		.INIT('h80)
	) name4480 (
		\wishbone_bd_ram_mem3_reg[17][25]/P0001 ,
		_w11935_,
		_w11977_,
		_w14993_
	);
	LUT3 #(
		.INIT('h80)
	) name4481 (
		\wishbone_bd_ram_mem3_reg[235][25]/P0001 ,
		_w11936_,
		_w11982_,
		_w14994_
	);
	LUT3 #(
		.INIT('h80)
	) name4482 (
		\wishbone_bd_ram_mem3_reg[141][25]/P0001 ,
		_w11955_,
		_w11966_,
		_w14995_
	);
	LUT3 #(
		.INIT('h80)
	) name4483 (
		\wishbone_bd_ram_mem3_reg[49][25]/P0001 ,
		_w11977_,
		_w11979_,
		_w14996_
	);
	LUT4 #(
		.INIT('h0001)
	) name4484 (
		_w14993_,
		_w14994_,
		_w14995_,
		_w14996_,
		_w14997_
	);
	LUT3 #(
		.INIT('h80)
	) name4485 (
		\wishbone_bd_ram_mem3_reg[12][25]/P0001 ,
		_w11932_,
		_w11954_,
		_w14998_
	);
	LUT3 #(
		.INIT('h80)
	) name4486 (
		\wishbone_bd_ram_mem3_reg[237][25]/P0001 ,
		_w11966_,
		_w11982_,
		_w14999_
	);
	LUT3 #(
		.INIT('h80)
	) name4487 (
		\wishbone_bd_ram_mem3_reg[68][25]/P0001 ,
		_w11929_,
		_w11949_,
		_w15000_
	);
	LUT3 #(
		.INIT('h80)
	) name4488 (
		\wishbone_bd_ram_mem3_reg[19][25]/P0001 ,
		_w11935_,
		_w11938_,
		_w15001_
	);
	LUT4 #(
		.INIT('h0001)
	) name4489 (
		_w14998_,
		_w14999_,
		_w15000_,
		_w15001_,
		_w15002_
	);
	LUT3 #(
		.INIT('h80)
	) name4490 (
		\wishbone_bd_ram_mem3_reg[13][25]/P0001 ,
		_w11932_,
		_w11966_,
		_w15003_
	);
	LUT3 #(
		.INIT('h80)
	) name4491 (
		\wishbone_bd_ram_mem3_reg[214][25]/P0001 ,
		_w11984_,
		_w11986_,
		_w15004_
	);
	LUT3 #(
		.INIT('h80)
	) name4492 (
		\wishbone_bd_ram_mem3_reg[156][25]/P0001 ,
		_w11954_,
		_w11959_,
		_w15005_
	);
	LUT3 #(
		.INIT('h80)
	) name4493 (
		\wishbone_bd_ram_mem3_reg[167][25]/P0001 ,
		_w11930_,
		_w11975_,
		_w15006_
	);
	LUT4 #(
		.INIT('h0001)
	) name4494 (
		_w15003_,
		_w15004_,
		_w15005_,
		_w15006_,
		_w15007_
	);
	LUT4 #(
		.INIT('h8000)
	) name4495 (
		_w14992_,
		_w14997_,
		_w15002_,
		_w15007_,
		_w15008_
	);
	LUT3 #(
		.INIT('h80)
	) name4496 (
		\wishbone_bd_ram_mem3_reg[225][25]/P0001 ,
		_w11977_,
		_w11982_,
		_w15009_
	);
	LUT3 #(
		.INIT('h80)
	) name4497 (
		\wishbone_bd_ram_mem3_reg[22][25]/P0001 ,
		_w11935_,
		_w11986_,
		_w15010_
	);
	LUT3 #(
		.INIT('h80)
	) name4498 (
		\wishbone_bd_ram_mem3_reg[203][25]/P0001 ,
		_w11936_,
		_w11945_,
		_w15011_
	);
	LUT3 #(
		.INIT('h80)
	) name4499 (
		\wishbone_bd_ram_mem3_reg[209][25]/P0001 ,
		_w11977_,
		_w11984_,
		_w15012_
	);
	LUT4 #(
		.INIT('h0001)
	) name4500 (
		_w15009_,
		_w15010_,
		_w15011_,
		_w15012_,
		_w15013_
	);
	LUT3 #(
		.INIT('h80)
	) name4501 (
		\wishbone_bd_ram_mem3_reg[161][25]/P0001 ,
		_w11930_,
		_w11977_,
		_w15014_
	);
	LUT3 #(
		.INIT('h80)
	) name4502 (
		\wishbone_bd_ram_mem3_reg[184][25]/P0001 ,
		_w11942_,
		_w11990_,
		_w15015_
	);
	LUT3 #(
		.INIT('h80)
	) name4503 (
		\wishbone_bd_ram_mem3_reg[89][25]/P0001 ,
		_w11968_,
		_w11972_,
		_w15016_
	);
	LUT3 #(
		.INIT('h80)
	) name4504 (
		\wishbone_bd_ram_mem3_reg[26][25]/P0001 ,
		_w11935_,
		_w11944_,
		_w15017_
	);
	LUT4 #(
		.INIT('h0001)
	) name4505 (
		_w15014_,
		_w15015_,
		_w15016_,
		_w15017_,
		_w15018_
	);
	LUT3 #(
		.INIT('h80)
	) name4506 (
		\wishbone_bd_ram_mem3_reg[240][25]/P0001 ,
		_w11941_,
		_w11952_,
		_w15019_
	);
	LUT3 #(
		.INIT('h80)
	) name4507 (
		\wishbone_bd_ram_mem3_reg[84][25]/P0001 ,
		_w11929_,
		_w11972_,
		_w15020_
	);
	LUT3 #(
		.INIT('h80)
	) name4508 (
		\wishbone_bd_ram_mem3_reg[198][25]/P0001 ,
		_w11945_,
		_w11986_,
		_w15021_
	);
	LUT3 #(
		.INIT('h80)
	) name4509 (
		\wishbone_bd_ram_mem3_reg[197][25]/P0001 ,
		_w11933_,
		_w11945_,
		_w15022_
	);
	LUT4 #(
		.INIT('h0001)
	) name4510 (
		_w15019_,
		_w15020_,
		_w15021_,
		_w15022_,
		_w15023_
	);
	LUT3 #(
		.INIT('h80)
	) name4511 (
		\wishbone_bd_ram_mem3_reg[192][25]/P0001 ,
		_w11941_,
		_w11945_,
		_w15024_
	);
	LUT3 #(
		.INIT('h80)
	) name4512 (
		\wishbone_bd_ram_mem3_reg[215][25]/P0001 ,
		_w11975_,
		_w11984_,
		_w15025_
	);
	LUT3 #(
		.INIT('h80)
	) name4513 (
		\wishbone_bd_ram_mem3_reg[137][25]/P0001 ,
		_w11955_,
		_w11968_,
		_w15026_
	);
	LUT3 #(
		.INIT('h80)
	) name4514 (
		\wishbone_bd_ram_mem3_reg[117][25]/P0001 ,
		_w11933_,
		_w12012_,
		_w15027_
	);
	LUT4 #(
		.INIT('h0001)
	) name4515 (
		_w15024_,
		_w15025_,
		_w15026_,
		_w15027_,
		_w15028_
	);
	LUT4 #(
		.INIT('h8000)
	) name4516 (
		_w15013_,
		_w15018_,
		_w15023_,
		_w15028_,
		_w15029_
	);
	LUT3 #(
		.INIT('h80)
	) name4517 (
		\wishbone_bd_ram_mem3_reg[43][25]/P0001 ,
		_w11936_,
		_w11957_,
		_w15030_
	);
	LUT3 #(
		.INIT('h80)
	) name4518 (
		\wishbone_bd_ram_mem3_reg[48][25]/P0001 ,
		_w11941_,
		_w11979_,
		_w15031_
	);
	LUT3 #(
		.INIT('h80)
	) name4519 (
		\wishbone_bd_ram_mem3_reg[75][25]/P0001 ,
		_w11936_,
		_w11949_,
		_w15032_
	);
	LUT3 #(
		.INIT('h80)
	) name4520 (
		\wishbone_bd_ram_mem3_reg[142][25]/P0001 ,
		_w11948_,
		_w11955_,
		_w15033_
	);
	LUT4 #(
		.INIT('h0001)
	) name4521 (
		_w15030_,
		_w15031_,
		_w15032_,
		_w15033_,
		_w15034_
	);
	LUT3 #(
		.INIT('h80)
	) name4522 (
		\wishbone_bd_ram_mem3_reg[63][25]/P0001 ,
		_w11973_,
		_w11979_,
		_w15035_
	);
	LUT3 #(
		.INIT('h80)
	) name4523 (
		\wishbone_bd_ram_mem3_reg[201][25]/P0001 ,
		_w11945_,
		_w11968_,
		_w15036_
	);
	LUT3 #(
		.INIT('h80)
	) name4524 (
		\wishbone_bd_ram_mem3_reg[76][25]/P0001 ,
		_w11949_,
		_w11954_,
		_w15037_
	);
	LUT3 #(
		.INIT('h80)
	) name4525 (
		\wishbone_bd_ram_mem3_reg[134][25]/P0001 ,
		_w11955_,
		_w11986_,
		_w15038_
	);
	LUT4 #(
		.INIT('h0001)
	) name4526 (
		_w15035_,
		_w15036_,
		_w15037_,
		_w15038_,
		_w15039_
	);
	LUT3 #(
		.INIT('h80)
	) name4527 (
		\wishbone_bd_ram_mem3_reg[224][25]/P0001 ,
		_w11941_,
		_w11982_,
		_w15040_
	);
	LUT3 #(
		.INIT('h80)
	) name4528 (
		\wishbone_bd_ram_mem3_reg[35][25]/P0001 ,
		_w11938_,
		_w11957_,
		_w15041_
	);
	LUT3 #(
		.INIT('h80)
	) name4529 (
		\wishbone_bd_ram_mem3_reg[31][25]/P0001 ,
		_w11935_,
		_w11973_,
		_w15042_
	);
	LUT3 #(
		.INIT('h80)
	) name4530 (
		\wishbone_bd_ram_mem3_reg[187][25]/P0001 ,
		_w11936_,
		_w11942_,
		_w15043_
	);
	LUT4 #(
		.INIT('h0001)
	) name4531 (
		_w15040_,
		_w15041_,
		_w15042_,
		_w15043_,
		_w15044_
	);
	LUT3 #(
		.INIT('h80)
	) name4532 (
		\wishbone_bd_ram_mem3_reg[236][25]/P0001 ,
		_w11954_,
		_w11982_,
		_w15045_
	);
	LUT3 #(
		.INIT('h80)
	) name4533 (
		\wishbone_bd_ram_mem3_reg[238][25]/P0001 ,
		_w11948_,
		_w11982_,
		_w15046_
	);
	LUT3 #(
		.INIT('h80)
	) name4534 (
		\wishbone_bd_ram_mem3_reg[174][25]/P0001 ,
		_w11930_,
		_w11948_,
		_w15047_
	);
	LUT3 #(
		.INIT('h80)
	) name4535 (
		\wishbone_bd_ram_mem3_reg[62][25]/P0001 ,
		_w11948_,
		_w11979_,
		_w15048_
	);
	LUT4 #(
		.INIT('h0001)
	) name4536 (
		_w15045_,
		_w15046_,
		_w15047_,
		_w15048_,
		_w15049_
	);
	LUT4 #(
		.INIT('h8000)
	) name4537 (
		_w15034_,
		_w15039_,
		_w15044_,
		_w15049_,
		_w15050_
	);
	LUT4 #(
		.INIT('h8000)
	) name4538 (
		_w14987_,
		_w15008_,
		_w15029_,
		_w15050_,
		_w15051_
	);
	LUT3 #(
		.INIT('h80)
	) name4539 (
		\wishbone_bd_ram_mem3_reg[171][25]/P0001 ,
		_w11930_,
		_w11936_,
		_w15052_
	);
	LUT3 #(
		.INIT('h80)
	) name4540 (
		\wishbone_bd_ram_mem3_reg[255][25]/P0001 ,
		_w11952_,
		_w11973_,
		_w15053_
	);
	LUT3 #(
		.INIT('h80)
	) name4541 (
		\wishbone_bd_ram_mem3_reg[45][25]/P0001 ,
		_w11957_,
		_w11966_,
		_w15054_
	);
	LUT3 #(
		.INIT('h80)
	) name4542 (
		\wishbone_bd_ram_mem3_reg[226][25]/P0001 ,
		_w11963_,
		_w11982_,
		_w15055_
	);
	LUT4 #(
		.INIT('h0001)
	) name4543 (
		_w15052_,
		_w15053_,
		_w15054_,
		_w15055_,
		_w15056_
	);
	LUT3 #(
		.INIT('h80)
	) name4544 (
		\wishbone_bd_ram_mem3_reg[135][25]/P0001 ,
		_w11955_,
		_w11975_,
		_w15057_
	);
	LUT3 #(
		.INIT('h80)
	) name4545 (
		\wishbone_bd_ram_mem3_reg[2][25]/P0001 ,
		_w11932_,
		_w11963_,
		_w15058_
	);
	LUT3 #(
		.INIT('h80)
	) name4546 (
		\wishbone_bd_ram_mem3_reg[248][25]/P0001 ,
		_w11952_,
		_w11990_,
		_w15059_
	);
	LUT3 #(
		.INIT('h80)
	) name4547 (
		\wishbone_bd_ram_mem3_reg[87][25]/P0001 ,
		_w11972_,
		_w11975_,
		_w15060_
	);
	LUT4 #(
		.INIT('h0001)
	) name4548 (
		_w15057_,
		_w15058_,
		_w15059_,
		_w15060_,
		_w15061_
	);
	LUT3 #(
		.INIT('h80)
	) name4549 (
		\wishbone_bd_ram_mem3_reg[148][25]/P0001 ,
		_w11929_,
		_w11959_,
		_w15062_
	);
	LUT3 #(
		.INIT('h80)
	) name4550 (
		\wishbone_bd_ram_mem3_reg[95][25]/P0001 ,
		_w11972_,
		_w11973_,
		_w15063_
	);
	LUT3 #(
		.INIT('h80)
	) name4551 (
		\wishbone_bd_ram_mem3_reg[113][25]/P0001 ,
		_w11977_,
		_w12012_,
		_w15064_
	);
	LUT3 #(
		.INIT('h80)
	) name4552 (
		\wishbone_bd_ram_mem3_reg[150][25]/P0001 ,
		_w11959_,
		_w11986_,
		_w15065_
	);
	LUT4 #(
		.INIT('h0001)
	) name4553 (
		_w15062_,
		_w15063_,
		_w15064_,
		_w15065_,
		_w15066_
	);
	LUT3 #(
		.INIT('h80)
	) name4554 (
		\wishbone_bd_ram_mem3_reg[119][25]/P0001 ,
		_w11975_,
		_w12012_,
		_w15067_
	);
	LUT3 #(
		.INIT('h80)
	) name4555 (
		\wishbone_bd_ram_mem3_reg[88][25]/P0001 ,
		_w11972_,
		_w11990_,
		_w15068_
	);
	LUT3 #(
		.INIT('h80)
	) name4556 (
		\wishbone_bd_ram_mem3_reg[82][25]/P0001 ,
		_w11963_,
		_w11972_,
		_w15069_
	);
	LUT3 #(
		.INIT('h80)
	) name4557 (
		\wishbone_bd_ram_mem3_reg[155][25]/P0001 ,
		_w11936_,
		_w11959_,
		_w15070_
	);
	LUT4 #(
		.INIT('h0001)
	) name4558 (
		_w15067_,
		_w15068_,
		_w15069_,
		_w15070_,
		_w15071_
	);
	LUT4 #(
		.INIT('h8000)
	) name4559 (
		_w15056_,
		_w15061_,
		_w15066_,
		_w15071_,
		_w15072_
	);
	LUT3 #(
		.INIT('h80)
	) name4560 (
		\wishbone_bd_ram_mem3_reg[208][25]/P0001 ,
		_w11941_,
		_w11984_,
		_w15073_
	);
	LUT3 #(
		.INIT('h80)
	) name4561 (
		\wishbone_bd_ram_mem3_reg[66][25]/P0001 ,
		_w11949_,
		_w11963_,
		_w15074_
	);
	LUT3 #(
		.INIT('h80)
	) name4562 (
		\wishbone_bd_ram_mem3_reg[30][25]/P0001 ,
		_w11935_,
		_w11948_,
		_w15075_
	);
	LUT3 #(
		.INIT('h80)
	) name4563 (
		\wishbone_bd_ram_mem3_reg[40][25]/P0001 ,
		_w11957_,
		_w11990_,
		_w15076_
	);
	LUT4 #(
		.INIT('h0001)
	) name4564 (
		_w15073_,
		_w15074_,
		_w15075_,
		_w15076_,
		_w15077_
	);
	LUT3 #(
		.INIT('h80)
	) name4565 (
		\wishbone_bd_ram_mem3_reg[239][25]/P0001 ,
		_w11973_,
		_w11982_,
		_w15078_
	);
	LUT3 #(
		.INIT('h80)
	) name4566 (
		\wishbone_bd_ram_mem3_reg[46][25]/P0001 ,
		_w11948_,
		_w11957_,
		_w15079_
	);
	LUT3 #(
		.INIT('h80)
	) name4567 (
		\wishbone_bd_ram_mem3_reg[99][25]/P0001 ,
		_w11938_,
		_w11965_,
		_w15080_
	);
	LUT3 #(
		.INIT('h80)
	) name4568 (
		\wishbone_bd_ram_mem3_reg[54][25]/P0001 ,
		_w11979_,
		_w11986_,
		_w15081_
	);
	LUT4 #(
		.INIT('h0001)
	) name4569 (
		_w15078_,
		_w15079_,
		_w15080_,
		_w15081_,
		_w15082_
	);
	LUT3 #(
		.INIT('h80)
	) name4570 (
		\wishbone_bd_ram_mem3_reg[9][25]/P0001 ,
		_w11932_,
		_w11968_,
		_w15083_
	);
	LUT3 #(
		.INIT('h80)
	) name4571 (
		\wishbone_bd_ram_mem3_reg[65][25]/P0001 ,
		_w11949_,
		_w11977_,
		_w15084_
	);
	LUT3 #(
		.INIT('h80)
	) name4572 (
		\wishbone_bd_ram_mem3_reg[25][25]/P0001 ,
		_w11935_,
		_w11968_,
		_w15085_
	);
	LUT3 #(
		.INIT('h80)
	) name4573 (
		\wishbone_bd_ram_mem3_reg[6][25]/P0001 ,
		_w11932_,
		_w11986_,
		_w15086_
	);
	LUT4 #(
		.INIT('h0001)
	) name4574 (
		_w15083_,
		_w15084_,
		_w15085_,
		_w15086_,
		_w15087_
	);
	LUT3 #(
		.INIT('h80)
	) name4575 (
		\wishbone_bd_ram_mem3_reg[83][25]/P0001 ,
		_w11938_,
		_w11972_,
		_w15088_
	);
	LUT3 #(
		.INIT('h80)
	) name4576 (
		\wishbone_bd_ram_mem3_reg[139][25]/P0001 ,
		_w11936_,
		_w11955_,
		_w15089_
	);
	LUT3 #(
		.INIT('h80)
	) name4577 (
		\wishbone_bd_ram_mem3_reg[115][25]/P0001 ,
		_w11938_,
		_w12012_,
		_w15090_
	);
	LUT3 #(
		.INIT('h80)
	) name4578 (
		\wishbone_bd_ram_mem3_reg[158][25]/P0001 ,
		_w11948_,
		_w11959_,
		_w15091_
	);
	LUT4 #(
		.INIT('h0001)
	) name4579 (
		_w15088_,
		_w15089_,
		_w15090_,
		_w15091_,
		_w15092_
	);
	LUT4 #(
		.INIT('h8000)
	) name4580 (
		_w15077_,
		_w15082_,
		_w15087_,
		_w15092_,
		_w15093_
	);
	LUT3 #(
		.INIT('h80)
	) name4581 (
		\wishbone_bd_ram_mem3_reg[178][25]/P0001 ,
		_w11942_,
		_w11963_,
		_w15094_
	);
	LUT3 #(
		.INIT('h80)
	) name4582 (
		\wishbone_bd_ram_mem3_reg[14][25]/P0001 ,
		_w11932_,
		_w11948_,
		_w15095_
	);
	LUT3 #(
		.INIT('h80)
	) name4583 (
		\wishbone_bd_ram_mem3_reg[204][25]/P0001 ,
		_w11945_,
		_w11954_,
		_w15096_
	);
	LUT3 #(
		.INIT('h80)
	) name4584 (
		\wishbone_bd_ram_mem3_reg[118][25]/P0001 ,
		_w11986_,
		_w12012_,
		_w15097_
	);
	LUT4 #(
		.INIT('h0001)
	) name4585 (
		_w15094_,
		_w15095_,
		_w15096_,
		_w15097_,
		_w15098_
	);
	LUT3 #(
		.INIT('h80)
	) name4586 (
		\wishbone_bd_ram_mem3_reg[181][25]/P0001 ,
		_w11933_,
		_w11942_,
		_w15099_
	);
	LUT3 #(
		.INIT('h80)
	) name4587 (
		\wishbone_bd_ram_mem3_reg[193][25]/P0001 ,
		_w11945_,
		_w11977_,
		_w15100_
	);
	LUT3 #(
		.INIT('h80)
	) name4588 (
		\wishbone_bd_ram_mem3_reg[28][25]/P0001 ,
		_w11935_,
		_w11954_,
		_w15101_
	);
	LUT3 #(
		.INIT('h80)
	) name4589 (
		\wishbone_bd_ram_mem3_reg[210][25]/P0001 ,
		_w11963_,
		_w11984_,
		_w15102_
	);
	LUT4 #(
		.INIT('h0001)
	) name4590 (
		_w15099_,
		_w15100_,
		_w15101_,
		_w15102_,
		_w15103_
	);
	LUT3 #(
		.INIT('h80)
	) name4591 (
		\wishbone_bd_ram_mem3_reg[27][25]/P0001 ,
		_w11935_,
		_w11936_,
		_w15104_
	);
	LUT3 #(
		.INIT('h80)
	) name4592 (
		\wishbone_bd_ram_mem3_reg[129][25]/P0001 ,
		_w11955_,
		_w11977_,
		_w15105_
	);
	LUT3 #(
		.INIT('h80)
	) name4593 (
		\wishbone_bd_ram_mem3_reg[20][25]/P0001 ,
		_w11929_,
		_w11935_,
		_w15106_
	);
	LUT3 #(
		.INIT('h80)
	) name4594 (
		\wishbone_bd_ram_mem3_reg[200][25]/P0001 ,
		_w11945_,
		_w11990_,
		_w15107_
	);
	LUT4 #(
		.INIT('h0001)
	) name4595 (
		_w15104_,
		_w15105_,
		_w15106_,
		_w15107_,
		_w15108_
	);
	LUT3 #(
		.INIT('h80)
	) name4596 (
		\wishbone_bd_ram_mem3_reg[67][25]/P0001 ,
		_w11938_,
		_w11949_,
		_w15109_
	);
	LUT3 #(
		.INIT('h80)
	) name4597 (
		\wishbone_bd_ram_mem3_reg[10][25]/P0001 ,
		_w11932_,
		_w11944_,
		_w15110_
	);
	LUT3 #(
		.INIT('h80)
	) name4598 (
		\wishbone_bd_ram_mem3_reg[123][25]/P0001 ,
		_w11936_,
		_w12012_,
		_w15111_
	);
	LUT3 #(
		.INIT('h80)
	) name4599 (
		\wishbone_bd_ram_mem3_reg[207][25]/P0001 ,
		_w11945_,
		_w11973_,
		_w15112_
	);
	LUT4 #(
		.INIT('h0001)
	) name4600 (
		_w15109_,
		_w15110_,
		_w15111_,
		_w15112_,
		_w15113_
	);
	LUT4 #(
		.INIT('h8000)
	) name4601 (
		_w15098_,
		_w15103_,
		_w15108_,
		_w15113_,
		_w15114_
	);
	LUT3 #(
		.INIT('h80)
	) name4602 (
		\wishbone_bd_ram_mem3_reg[104][25]/P0001 ,
		_w11965_,
		_w11990_,
		_w15115_
	);
	LUT3 #(
		.INIT('h80)
	) name4603 (
		\wishbone_bd_ram_mem3_reg[212][25]/P0001 ,
		_w11929_,
		_w11984_,
		_w15116_
	);
	LUT3 #(
		.INIT('h80)
	) name4604 (
		\wishbone_bd_ram_mem3_reg[92][25]/P0001 ,
		_w11954_,
		_w11972_,
		_w15117_
	);
	LUT3 #(
		.INIT('h80)
	) name4605 (
		\wishbone_bd_ram_mem3_reg[91][25]/P0001 ,
		_w11936_,
		_w11972_,
		_w15118_
	);
	LUT4 #(
		.INIT('h0001)
	) name4606 (
		_w15115_,
		_w15116_,
		_w15117_,
		_w15118_,
		_w15119_
	);
	LUT3 #(
		.INIT('h80)
	) name4607 (
		\wishbone_bd_ram_mem3_reg[102][25]/P0001 ,
		_w11965_,
		_w11986_,
		_w15120_
	);
	LUT3 #(
		.INIT('h80)
	) name4608 (
		\wishbone_bd_ram_mem3_reg[173][25]/P0001 ,
		_w11930_,
		_w11966_,
		_w15121_
	);
	LUT3 #(
		.INIT('h80)
	) name4609 (
		\wishbone_bd_ram_mem3_reg[216][25]/P0001 ,
		_w11984_,
		_w11990_,
		_w15122_
	);
	LUT3 #(
		.INIT('h80)
	) name4610 (
		\wishbone_bd_ram_mem3_reg[246][25]/P0001 ,
		_w11952_,
		_w11986_,
		_w15123_
	);
	LUT4 #(
		.INIT('h0001)
	) name4611 (
		_w15120_,
		_w15121_,
		_w15122_,
		_w15123_,
		_w15124_
	);
	LUT3 #(
		.INIT('h80)
	) name4612 (
		\wishbone_bd_ram_mem3_reg[245][25]/P0001 ,
		_w11933_,
		_w11952_,
		_w15125_
	);
	LUT3 #(
		.INIT('h80)
	) name4613 (
		\wishbone_bd_ram_mem3_reg[56][25]/P0001 ,
		_w11979_,
		_w11990_,
		_w15126_
	);
	LUT3 #(
		.INIT('h80)
	) name4614 (
		\wishbone_bd_ram_mem3_reg[15][25]/P0001 ,
		_w11932_,
		_w11973_,
		_w15127_
	);
	LUT3 #(
		.INIT('h80)
	) name4615 (
		\wishbone_bd_ram_mem3_reg[132][25]/P0001 ,
		_w11929_,
		_w11955_,
		_w15128_
	);
	LUT4 #(
		.INIT('h0001)
	) name4616 (
		_w15125_,
		_w15126_,
		_w15127_,
		_w15128_,
		_w15129_
	);
	LUT3 #(
		.INIT('h80)
	) name4617 (
		\wishbone_bd_ram_mem3_reg[188][25]/P0001 ,
		_w11942_,
		_w11954_,
		_w15130_
	);
	LUT3 #(
		.INIT('h80)
	) name4618 (
		\wishbone_bd_ram_mem3_reg[107][25]/P0001 ,
		_w11936_,
		_w11965_,
		_w15131_
	);
	LUT3 #(
		.INIT('h80)
	) name4619 (
		\wishbone_bd_ram_mem3_reg[18][25]/P0001 ,
		_w11935_,
		_w11963_,
		_w15132_
	);
	LUT3 #(
		.INIT('h80)
	) name4620 (
		\wishbone_bd_ram_mem3_reg[120][25]/P0001 ,
		_w11990_,
		_w12012_,
		_w15133_
	);
	LUT4 #(
		.INIT('h0001)
	) name4621 (
		_w15130_,
		_w15131_,
		_w15132_,
		_w15133_,
		_w15134_
	);
	LUT4 #(
		.INIT('h8000)
	) name4622 (
		_w15119_,
		_w15124_,
		_w15129_,
		_w15134_,
		_w15135_
	);
	LUT4 #(
		.INIT('h8000)
	) name4623 (
		_w15072_,
		_w15093_,
		_w15114_,
		_w15135_,
		_w15136_
	);
	LUT3 #(
		.INIT('h80)
	) name4624 (
		\wishbone_bd_ram_mem3_reg[78][25]/P0001 ,
		_w11948_,
		_w11949_,
		_w15137_
	);
	LUT3 #(
		.INIT('h80)
	) name4625 (
		\wishbone_bd_ram_mem3_reg[162][25]/P0001 ,
		_w11930_,
		_w11963_,
		_w15138_
	);
	LUT3 #(
		.INIT('h80)
	) name4626 (
		\wishbone_bd_ram_mem3_reg[138][25]/P0001 ,
		_w11944_,
		_w11955_,
		_w15139_
	);
	LUT3 #(
		.INIT('h80)
	) name4627 (
		\wishbone_bd_ram_mem3_reg[41][25]/P0001 ,
		_w11957_,
		_w11968_,
		_w15140_
	);
	LUT4 #(
		.INIT('h0001)
	) name4628 (
		_w15137_,
		_w15138_,
		_w15139_,
		_w15140_,
		_w15141_
	);
	LUT3 #(
		.INIT('h80)
	) name4629 (
		\wishbone_bd_ram_mem3_reg[80][25]/P0001 ,
		_w11941_,
		_w11972_,
		_w15142_
	);
	LUT3 #(
		.INIT('h80)
	) name4630 (
		\wishbone_bd_ram_mem3_reg[116][25]/P0001 ,
		_w11929_,
		_w12012_,
		_w15143_
	);
	LUT3 #(
		.INIT('h80)
	) name4631 (
		\wishbone_bd_ram_mem3_reg[131][25]/P0001 ,
		_w11938_,
		_w11955_,
		_w15144_
	);
	LUT3 #(
		.INIT('h80)
	) name4632 (
		\wishbone_bd_ram_mem3_reg[249][25]/P0001 ,
		_w11952_,
		_w11968_,
		_w15145_
	);
	LUT4 #(
		.INIT('h0001)
	) name4633 (
		_w15142_,
		_w15143_,
		_w15144_,
		_w15145_,
		_w15146_
	);
	LUT3 #(
		.INIT('h80)
	) name4634 (
		\wishbone_bd_ram_mem3_reg[147][25]/P0001 ,
		_w11938_,
		_w11959_,
		_w15147_
	);
	LUT3 #(
		.INIT('h80)
	) name4635 (
		\wishbone_bd_ram_mem3_reg[133][25]/P0001 ,
		_w11933_,
		_w11955_,
		_w15148_
	);
	LUT3 #(
		.INIT('h80)
	) name4636 (
		\wishbone_bd_ram_mem3_reg[97][25]/P0001 ,
		_w11965_,
		_w11977_,
		_w15149_
	);
	LUT3 #(
		.INIT('h80)
	) name4637 (
		\wishbone_bd_ram_mem3_reg[114][25]/P0001 ,
		_w11963_,
		_w12012_,
		_w15150_
	);
	LUT4 #(
		.INIT('h0001)
	) name4638 (
		_w15147_,
		_w15148_,
		_w15149_,
		_w15150_,
		_w15151_
	);
	LUT3 #(
		.INIT('h80)
	) name4639 (
		\wishbone_bd_ram_mem3_reg[73][25]/P0001 ,
		_w11949_,
		_w11968_,
		_w15152_
	);
	LUT3 #(
		.INIT('h80)
	) name4640 (
		\wishbone_bd_ram_mem3_reg[58][25]/P0001 ,
		_w11944_,
		_w11979_,
		_w15153_
	);
	LUT3 #(
		.INIT('h80)
	) name4641 (
		\wishbone_bd_ram_mem3_reg[7][25]/P0001 ,
		_w11932_,
		_w11975_,
		_w15154_
	);
	LUT3 #(
		.INIT('h80)
	) name4642 (
		\wishbone_bd_ram_mem3_reg[151][25]/P0001 ,
		_w11959_,
		_w11975_,
		_w15155_
	);
	LUT4 #(
		.INIT('h0001)
	) name4643 (
		_w15152_,
		_w15153_,
		_w15154_,
		_w15155_,
		_w15156_
	);
	LUT4 #(
		.INIT('h8000)
	) name4644 (
		_w15141_,
		_w15146_,
		_w15151_,
		_w15156_,
		_w15157_
	);
	LUT3 #(
		.INIT('h80)
	) name4645 (
		\wishbone_bd_ram_mem3_reg[145][25]/P0001 ,
		_w11959_,
		_w11977_,
		_w15158_
	);
	LUT3 #(
		.INIT('h80)
	) name4646 (
		\wishbone_bd_ram_mem3_reg[11][25]/P0001 ,
		_w11932_,
		_w11936_,
		_w15159_
	);
	LUT3 #(
		.INIT('h80)
	) name4647 (
		\wishbone_bd_ram_mem3_reg[21][25]/P0001 ,
		_w11933_,
		_w11935_,
		_w15160_
	);
	LUT3 #(
		.INIT('h80)
	) name4648 (
		\wishbone_bd_ram_mem3_reg[121][25]/P0001 ,
		_w11968_,
		_w12012_,
		_w15161_
	);
	LUT4 #(
		.INIT('h0001)
	) name4649 (
		_w15158_,
		_w15159_,
		_w15160_,
		_w15161_,
		_w15162_
	);
	LUT3 #(
		.INIT('h80)
	) name4650 (
		\wishbone_bd_ram_mem3_reg[125][25]/P0001 ,
		_w11966_,
		_w12012_,
		_w15163_
	);
	LUT3 #(
		.INIT('h80)
	) name4651 (
		\wishbone_bd_ram_mem3_reg[44][25]/P0001 ,
		_w11954_,
		_w11957_,
		_w15164_
	);
	LUT3 #(
		.INIT('h80)
	) name4652 (
		\wishbone_bd_ram_mem3_reg[70][25]/P0001 ,
		_w11949_,
		_w11986_,
		_w15165_
	);
	LUT3 #(
		.INIT('h80)
	) name4653 (
		\wishbone_bd_ram_mem3_reg[206][25]/P0001 ,
		_w11945_,
		_w11948_,
		_w15166_
	);
	LUT4 #(
		.INIT('h0001)
	) name4654 (
		_w15163_,
		_w15164_,
		_w15165_,
		_w15166_,
		_w15167_
	);
	LUT3 #(
		.INIT('h80)
	) name4655 (
		\wishbone_bd_ram_mem3_reg[170][25]/P0001 ,
		_w11930_,
		_w11944_,
		_w15168_
	);
	LUT3 #(
		.INIT('h80)
	) name4656 (
		\wishbone_bd_ram_mem3_reg[71][25]/P0001 ,
		_w11949_,
		_w11975_,
		_w15169_
	);
	LUT3 #(
		.INIT('h80)
	) name4657 (
		\wishbone_bd_ram_mem3_reg[186][25]/P0001 ,
		_w11942_,
		_w11944_,
		_w15170_
	);
	LUT3 #(
		.INIT('h80)
	) name4658 (
		\wishbone_bd_ram_mem3_reg[37][25]/P0001 ,
		_w11933_,
		_w11957_,
		_w15171_
	);
	LUT4 #(
		.INIT('h0001)
	) name4659 (
		_w15168_,
		_w15169_,
		_w15170_,
		_w15171_,
		_w15172_
	);
	LUT3 #(
		.INIT('h80)
	) name4660 (
		\wishbone_bd_ram_mem3_reg[4][25]/P0001 ,
		_w11929_,
		_w11932_,
		_w15173_
	);
	LUT3 #(
		.INIT('h80)
	) name4661 (
		\wishbone_bd_ram_mem3_reg[33][25]/P0001 ,
		_w11957_,
		_w11977_,
		_w15174_
	);
	LUT3 #(
		.INIT('h80)
	) name4662 (
		\wishbone_bd_ram_mem3_reg[221][25]/P0001 ,
		_w11966_,
		_w11984_,
		_w15175_
	);
	LUT3 #(
		.INIT('h80)
	) name4663 (
		\wishbone_bd_ram_mem3_reg[168][25]/P0001 ,
		_w11930_,
		_w11990_,
		_w15176_
	);
	LUT4 #(
		.INIT('h0001)
	) name4664 (
		_w15173_,
		_w15174_,
		_w15175_,
		_w15176_,
		_w15177_
	);
	LUT4 #(
		.INIT('h8000)
	) name4665 (
		_w15162_,
		_w15167_,
		_w15172_,
		_w15177_,
		_w15178_
	);
	LUT3 #(
		.INIT('h80)
	) name4666 (
		\wishbone_bd_ram_mem3_reg[247][25]/P0001 ,
		_w11952_,
		_w11975_,
		_w15179_
	);
	LUT3 #(
		.INIT('h80)
	) name4667 (
		\wishbone_bd_ram_mem3_reg[103][25]/P0001 ,
		_w11965_,
		_w11975_,
		_w15180_
	);
	LUT3 #(
		.INIT('h80)
	) name4668 (
		\wishbone_bd_ram_mem3_reg[223][25]/P0001 ,
		_w11973_,
		_w11984_,
		_w15181_
	);
	LUT3 #(
		.INIT('h80)
	) name4669 (
		\wishbone_bd_ram_mem3_reg[228][25]/P0001 ,
		_w11929_,
		_w11982_,
		_w15182_
	);
	LUT4 #(
		.INIT('h0001)
	) name4670 (
		_w15179_,
		_w15180_,
		_w15181_,
		_w15182_,
		_w15183_
	);
	LUT3 #(
		.INIT('h80)
	) name4671 (
		\wishbone_bd_ram_mem3_reg[72][25]/P0001 ,
		_w11949_,
		_w11990_,
		_w15184_
	);
	LUT3 #(
		.INIT('h80)
	) name4672 (
		\wishbone_bd_ram_mem3_reg[182][25]/P0001 ,
		_w11942_,
		_w11986_,
		_w15185_
	);
	LUT3 #(
		.INIT('h80)
	) name4673 (
		\wishbone_bd_ram_mem3_reg[136][25]/P0001 ,
		_w11955_,
		_w11990_,
		_w15186_
	);
	LUT3 #(
		.INIT('h80)
	) name4674 (
		\wishbone_bd_ram_mem3_reg[185][25]/P0001 ,
		_w11942_,
		_w11968_,
		_w15187_
	);
	LUT4 #(
		.INIT('h0001)
	) name4675 (
		_w15184_,
		_w15185_,
		_w15186_,
		_w15187_,
		_w15188_
	);
	LUT3 #(
		.INIT('h80)
	) name4676 (
		\wishbone_bd_ram_mem3_reg[8][25]/P0001 ,
		_w11932_,
		_w11990_,
		_w15189_
	);
	LUT3 #(
		.INIT('h80)
	) name4677 (
		\wishbone_bd_ram_mem3_reg[219][25]/P0001 ,
		_w11936_,
		_w11984_,
		_w15190_
	);
	LUT3 #(
		.INIT('h80)
	) name4678 (
		\wishbone_bd_ram_mem3_reg[180][25]/P0001 ,
		_w11929_,
		_w11942_,
		_w15191_
	);
	LUT3 #(
		.INIT('h80)
	) name4679 (
		\wishbone_bd_ram_mem3_reg[23][25]/P0001 ,
		_w11935_,
		_w11975_,
		_w15192_
	);
	LUT4 #(
		.INIT('h0001)
	) name4680 (
		_w15189_,
		_w15190_,
		_w15191_,
		_w15192_,
		_w15193_
	);
	LUT3 #(
		.INIT('h80)
	) name4681 (
		\wishbone_bd_ram_mem3_reg[254][25]/P0001 ,
		_w11948_,
		_w11952_,
		_w15194_
	);
	LUT3 #(
		.INIT('h80)
	) name4682 (
		\wishbone_bd_ram_mem3_reg[146][25]/P0001 ,
		_w11959_,
		_w11963_,
		_w15195_
	);
	LUT3 #(
		.INIT('h80)
	) name4683 (
		\wishbone_bd_ram_mem3_reg[233][25]/P0001 ,
		_w11968_,
		_w11982_,
		_w15196_
	);
	LUT3 #(
		.INIT('h80)
	) name4684 (
		\wishbone_bd_ram_mem3_reg[69][25]/P0001 ,
		_w11933_,
		_w11949_,
		_w15197_
	);
	LUT4 #(
		.INIT('h0001)
	) name4685 (
		_w15194_,
		_w15195_,
		_w15196_,
		_w15197_,
		_w15198_
	);
	LUT4 #(
		.INIT('h8000)
	) name4686 (
		_w15183_,
		_w15188_,
		_w15193_,
		_w15198_,
		_w15199_
	);
	LUT3 #(
		.INIT('h80)
	) name4687 (
		\wishbone_bd_ram_mem3_reg[42][25]/P0001 ,
		_w11944_,
		_w11957_,
		_w15200_
	);
	LUT3 #(
		.INIT('h80)
	) name4688 (
		\wishbone_bd_ram_mem3_reg[163][25]/P0001 ,
		_w11930_,
		_w11938_,
		_w15201_
	);
	LUT3 #(
		.INIT('h80)
	) name4689 (
		\wishbone_bd_ram_mem3_reg[231][25]/P0001 ,
		_w11975_,
		_w11982_,
		_w15202_
	);
	LUT3 #(
		.INIT('h80)
	) name4690 (
		\wishbone_bd_ram_mem3_reg[16][25]/P0001 ,
		_w11935_,
		_w11941_,
		_w15203_
	);
	LUT4 #(
		.INIT('h0001)
	) name4691 (
		_w15200_,
		_w15201_,
		_w15202_,
		_w15203_,
		_w15204_
	);
	LUT3 #(
		.INIT('h80)
	) name4692 (
		\wishbone_bd_ram_mem3_reg[250][25]/P0001 ,
		_w11944_,
		_w11952_,
		_w15205_
	);
	LUT3 #(
		.INIT('h80)
	) name4693 (
		\wishbone_bd_ram_mem3_reg[244][25]/P0001 ,
		_w11929_,
		_w11952_,
		_w15206_
	);
	LUT3 #(
		.INIT('h80)
	) name4694 (
		\wishbone_bd_ram_mem3_reg[232][25]/P0001 ,
		_w11982_,
		_w11990_,
		_w15207_
	);
	LUT3 #(
		.INIT('h80)
	) name4695 (
		\wishbone_bd_ram_mem3_reg[175][25]/P0001 ,
		_w11930_,
		_w11973_,
		_w15208_
	);
	LUT4 #(
		.INIT('h0001)
	) name4696 (
		_w15205_,
		_w15206_,
		_w15207_,
		_w15208_,
		_w15209_
	);
	LUT3 #(
		.INIT('h80)
	) name4697 (
		\wishbone_bd_ram_mem3_reg[32][25]/P0001 ,
		_w11941_,
		_w11957_,
		_w15210_
	);
	LUT3 #(
		.INIT('h80)
	) name4698 (
		\wishbone_bd_ram_mem3_reg[194][25]/P0001 ,
		_w11945_,
		_w11963_,
		_w15211_
	);
	LUT3 #(
		.INIT('h80)
	) name4699 (
		\wishbone_bd_ram_mem3_reg[241][25]/P0001 ,
		_w11952_,
		_w11977_,
		_w15212_
	);
	LUT3 #(
		.INIT('h80)
	) name4700 (
		\wishbone_bd_ram_mem3_reg[53][25]/P0001 ,
		_w11933_,
		_w11979_,
		_w15213_
	);
	LUT4 #(
		.INIT('h0001)
	) name4701 (
		_w15210_,
		_w15211_,
		_w15212_,
		_w15213_,
		_w15214_
	);
	LUT3 #(
		.INIT('h80)
	) name4702 (
		\wishbone_bd_ram_mem3_reg[218][25]/P0001 ,
		_w11944_,
		_w11984_,
		_w15215_
	);
	LUT3 #(
		.INIT('h80)
	) name4703 (
		\wishbone_bd_ram_mem3_reg[111][25]/P0001 ,
		_w11965_,
		_w11973_,
		_w15216_
	);
	LUT3 #(
		.INIT('h80)
	) name4704 (
		\wishbone_bd_ram_mem3_reg[189][25]/P0001 ,
		_w11942_,
		_w11966_,
		_w15217_
	);
	LUT3 #(
		.INIT('h80)
	) name4705 (
		\wishbone_bd_ram_mem3_reg[191][25]/P0001 ,
		_w11942_,
		_w11973_,
		_w15218_
	);
	LUT4 #(
		.INIT('h0001)
	) name4706 (
		_w15215_,
		_w15216_,
		_w15217_,
		_w15218_,
		_w15219_
	);
	LUT4 #(
		.INIT('h8000)
	) name4707 (
		_w15204_,
		_w15209_,
		_w15214_,
		_w15219_,
		_w15220_
	);
	LUT4 #(
		.INIT('h8000)
	) name4708 (
		_w15157_,
		_w15178_,
		_w15199_,
		_w15220_,
		_w15221_
	);
	LUT4 #(
		.INIT('h8000)
	) name4709 (
		_w14966_,
		_w15051_,
		_w15136_,
		_w15221_,
		_w15222_
	);
	LUT3 #(
		.INIT('h10)
	) name4710 (
		\wishbone_TxLength_reg[7]/NET0131 ,
		\wishbone_TxLength_reg[8]/NET0131 ,
		\wishbone_TxLength_reg[9]/NET0131 ,
		_w15223_
	);
	LUT3 #(
		.INIT('h80)
	) name4711 (
		_w12309_,
		_w12310_,
		_w15223_,
		_w15224_
	);
	LUT3 #(
		.INIT('h0e)
	) name4712 (
		\wishbone_TxLength_reg[7]/NET0131 ,
		\wishbone_TxLength_reg[8]/NET0131 ,
		\wishbone_TxLength_reg[9]/NET0131 ,
		_w15225_
	);
	LUT4 #(
		.INIT('h00ea)
	) name4713 (
		\wishbone_TxLength_reg[9]/NET0131 ,
		_w12309_,
		_w12310_,
		_w15225_,
		_w15226_
	);
	LUT3 #(
		.INIT('hb0)
	) name4714 (
		_w14878_,
		_w15224_,
		_w15226_,
		_w15227_
	);
	LUT2 #(
		.INIT('h4)
	) name4715 (
		\wishbone_TxLength_reg[9]/NET0131 ,
		_w14878_,
		_w15228_
	);
	LUT2 #(
		.INIT('ha)
	) name4716 (
		_w12302_,
		_w12304_,
		_w15229_
	);
	LUT4 #(
		.INIT('he000)
	) name4717 (
		_w12302_,
		_w12304_,
		_w12314_,
		_w12316_,
		_w15230_
	);
	LUT3 #(
		.INIT('h13)
	) name4718 (
		_w12312_,
		_w15229_,
		_w15230_,
		_w15231_
	);
	LUT3 #(
		.INIT('h20)
	) name4719 (
		_w15227_,
		_w15228_,
		_w15231_,
		_w15232_
	);
	LUT3 #(
		.INIT('hf2)
	) name4720 (
		_w12303_,
		_w15222_,
		_w15232_,
		_w15233_
	);
	LUT2 #(
		.INIT('h2)
	) name4721 (
		\wishbone_RxDataLatched2_reg[0]/NET0131 ,
		_w13424_,
		_w15234_
	);
	LUT2 #(
		.INIT('h8)
	) name4722 (
		_w13423_,
		_w15234_,
		_w15235_
	);
	LUT3 #(
		.INIT('h02)
	) name4723 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w13423_,
		_w15236_
	);
	LUT3 #(
		.INIT('h02)
	) name4724 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		_w15237_
	);
	LUT3 #(
		.INIT('hd0)
	) name4725 (
		_w13423_,
		_w13424_,
		_w15237_,
		_w15238_
	);
	LUT3 #(
		.INIT('hfe)
	) name4726 (
		_w15235_,
		_w15236_,
		_w15238_,
		_w15239_
	);
	LUT2 #(
		.INIT('h2)
	) name4727 (
		\wishbone_RxDataLatched2_reg[1]/NET0131 ,
		_w13424_,
		_w15240_
	);
	LUT2 #(
		.INIT('h8)
	) name4728 (
		_w13423_,
		_w15240_,
		_w15241_
	);
	LUT3 #(
		.INIT('h02)
	) name4729 (
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w13423_,
		_w15242_
	);
	LUT3 #(
		.INIT('h02)
	) name4730 (
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		_w15243_
	);
	LUT3 #(
		.INIT('hd0)
	) name4731 (
		_w13423_,
		_w13424_,
		_w15243_,
		_w15244_
	);
	LUT3 #(
		.INIT('hfe)
	) name4732 (
		_w15241_,
		_w15242_,
		_w15244_,
		_w15245_
	);
	LUT2 #(
		.INIT('h2)
	) name4733 (
		\wishbone_RxDataLatched2_reg[2]/NET0131 ,
		_w13424_,
		_w15246_
	);
	LUT2 #(
		.INIT('h8)
	) name4734 (
		_w13423_,
		_w15246_,
		_w15247_
	);
	LUT3 #(
		.INIT('h02)
	) name4735 (
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w13423_,
		_w15248_
	);
	LUT3 #(
		.INIT('h02)
	) name4736 (
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		_w15249_
	);
	LUT3 #(
		.INIT('hd0)
	) name4737 (
		_w13423_,
		_w13424_,
		_w15249_,
		_w15250_
	);
	LUT3 #(
		.INIT('hfe)
	) name4738 (
		_w15247_,
		_w15248_,
		_w15250_,
		_w15251_
	);
	LUT2 #(
		.INIT('h2)
	) name4739 (
		\wishbone_RxDataLatched2_reg[3]/NET0131 ,
		_w13424_,
		_w15252_
	);
	LUT2 #(
		.INIT('h8)
	) name4740 (
		_w13423_,
		_w15252_,
		_w15253_
	);
	LUT3 #(
		.INIT('h02)
	) name4741 (
		\rxethmac1_RxData_reg[3]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w13423_,
		_w15254_
	);
	LUT3 #(
		.INIT('h02)
	) name4742 (
		\rxethmac1_RxData_reg[3]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		_w15255_
	);
	LUT3 #(
		.INIT('hd0)
	) name4743 (
		_w13423_,
		_w13424_,
		_w15255_,
		_w15256_
	);
	LUT3 #(
		.INIT('hfe)
	) name4744 (
		_w15253_,
		_w15254_,
		_w15256_,
		_w15257_
	);
	LUT2 #(
		.INIT('h2)
	) name4745 (
		\wishbone_RxDataLatched2_reg[5]/NET0131 ,
		_w13424_,
		_w15258_
	);
	LUT2 #(
		.INIT('h8)
	) name4746 (
		_w13423_,
		_w15258_,
		_w15259_
	);
	LUT3 #(
		.INIT('h02)
	) name4747 (
		\rxethmac1_RxData_reg[5]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w13423_,
		_w15260_
	);
	LUT3 #(
		.INIT('h02)
	) name4748 (
		\rxethmac1_RxData_reg[5]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		_w15261_
	);
	LUT3 #(
		.INIT('hd0)
	) name4749 (
		_w13423_,
		_w13424_,
		_w15261_,
		_w15262_
	);
	LUT3 #(
		.INIT('hfe)
	) name4750 (
		_w15259_,
		_w15260_,
		_w15262_,
		_w15263_
	);
	LUT2 #(
		.INIT('h2)
	) name4751 (
		\wishbone_RxDataLatched2_reg[4]/NET0131 ,
		_w13424_,
		_w15264_
	);
	LUT2 #(
		.INIT('h8)
	) name4752 (
		_w13423_,
		_w15264_,
		_w15265_
	);
	LUT3 #(
		.INIT('h02)
	) name4753 (
		\rxethmac1_RxData_reg[4]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w13423_,
		_w15266_
	);
	LUT3 #(
		.INIT('h02)
	) name4754 (
		\rxethmac1_RxData_reg[4]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		_w15267_
	);
	LUT3 #(
		.INIT('hd0)
	) name4755 (
		_w13423_,
		_w13424_,
		_w15267_,
		_w15268_
	);
	LUT3 #(
		.INIT('hfe)
	) name4756 (
		_w15265_,
		_w15266_,
		_w15268_,
		_w15269_
	);
	LUT2 #(
		.INIT('h2)
	) name4757 (
		\wishbone_RxDataLatched2_reg[6]/NET0131 ,
		_w13424_,
		_w15270_
	);
	LUT2 #(
		.INIT('h8)
	) name4758 (
		_w13423_,
		_w15270_,
		_w15271_
	);
	LUT3 #(
		.INIT('h02)
	) name4759 (
		\rxethmac1_RxData_reg[6]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w13423_,
		_w15272_
	);
	LUT3 #(
		.INIT('h02)
	) name4760 (
		\rxethmac1_RxData_reg[6]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		_w15273_
	);
	LUT3 #(
		.INIT('hd0)
	) name4761 (
		_w13423_,
		_w13424_,
		_w15273_,
		_w15274_
	);
	LUT3 #(
		.INIT('hfe)
	) name4762 (
		_w15271_,
		_w15272_,
		_w15274_,
		_w15275_
	);
	LUT2 #(
		.INIT('h2)
	) name4763 (
		\wishbone_RxDataLatched2_reg[7]/NET0131 ,
		_w13424_,
		_w15276_
	);
	LUT2 #(
		.INIT('h8)
	) name4764 (
		_w13423_,
		_w15276_,
		_w15277_
	);
	LUT3 #(
		.INIT('h02)
	) name4765 (
		\rxethmac1_RxData_reg[7]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w13423_,
		_w15278_
	);
	LUT3 #(
		.INIT('h02)
	) name4766 (
		\rxethmac1_RxData_reg[7]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		_w15279_
	);
	LUT3 #(
		.INIT('hd0)
	) name4767 (
		_w13423_,
		_w13424_,
		_w15279_,
		_w15280_
	);
	LUT3 #(
		.INIT('hfe)
	) name4768 (
		_w15277_,
		_w15278_,
		_w15280_,
		_w15281_
	);
	LUT4 #(
		.INIT('h4000)
	) name4769 (
		wb_rst_i_pad,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w15282_
	);
	LUT4 #(
		.INIT('h8000)
	) name4770 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_RxPointerMSB_reg[2]/NET0131 ,
		\wishbone_RxPointerMSB_reg[3]/NET0131 ,
		_w15283_
	);
	LUT3 #(
		.INIT('h80)
	) name4771 (
		\wishbone_RxPointerMSB_reg[4]/NET0131 ,
		\wishbone_RxPointerMSB_reg[5]/NET0131 ,
		\wishbone_RxPointerMSB_reg[6]/NET0131 ,
		_w15284_
	);
	LUT4 #(
		.INIT('h8000)
	) name4772 (
		\wishbone_RxPointerMSB_reg[10]/NET0131 ,
		\wishbone_RxPointerMSB_reg[7]/NET0131 ,
		\wishbone_RxPointerMSB_reg[8]/NET0131 ,
		\wishbone_RxPointerMSB_reg[9]/NET0131 ,
		_w15285_
	);
	LUT3 #(
		.INIT('h80)
	) name4773 (
		_w15283_,
		_w15284_,
		_w15285_,
		_w15286_
	);
	LUT4 #(
		.INIT('h8000)
	) name4774 (
		\wishbone_RxPointerMSB_reg[11]/NET0131 ,
		\wishbone_RxPointerMSB_reg[12]/NET0131 ,
		\wishbone_RxPointerMSB_reg[13]/NET0131 ,
		\wishbone_RxPointerMSB_reg[14]/NET0131 ,
		_w15287_
	);
	LUT4 #(
		.INIT('h8000)
	) name4775 (
		_w15283_,
		_w15284_,
		_w15285_,
		_w15287_,
		_w15288_
	);
	LUT4 #(
		.INIT('h8000)
	) name4776 (
		\wishbone_RxPointerMSB_reg[16]/NET0131 ,
		\wishbone_RxPointerMSB_reg[17]/NET0131 ,
		\wishbone_RxPointerMSB_reg[18]/NET0131 ,
		\wishbone_RxPointerMSB_reg[19]/NET0131 ,
		_w15289_
	);
	LUT2 #(
		.INIT('h8)
	) name4777 (
		\wishbone_RxPointerMSB_reg[15]/NET0131 ,
		\wishbone_RxPointerMSB_reg[20]/NET0131 ,
		_w15290_
	);
	LUT2 #(
		.INIT('h8)
	) name4778 (
		_w15289_,
		_w15290_,
		_w15291_
	);
	LUT2 #(
		.INIT('h8)
	) name4779 (
		\wishbone_RxPointerMSB_reg[21]/NET0131 ,
		\wishbone_RxPointerMSB_reg[22]/NET0131 ,
		_w15292_
	);
	LUT4 #(
		.INIT('h8000)
	) name4780 (
		\wishbone_RxPointerMSB_reg[21]/NET0131 ,
		\wishbone_RxPointerMSB_reg[22]/NET0131 ,
		\wishbone_RxPointerMSB_reg[23]/NET0131 ,
		\wishbone_RxPointerMSB_reg[24]/NET0131 ,
		_w15293_
	);
	LUT3 #(
		.INIT('h80)
	) name4781 (
		\wishbone_RxPointerMSB_reg[26]/NET0131 ,
		\wishbone_RxPointerMSB_reg[27]/NET0131 ,
		\wishbone_RxPointerMSB_reg[28]/NET0131 ,
		_w15294_
	);
	LUT2 #(
		.INIT('h8)
	) name4782 (
		\wishbone_RxPointerMSB_reg[25]/NET0131 ,
		\wishbone_RxPointerMSB_reg[29]/NET0131 ,
		_w15295_
	);
	LUT2 #(
		.INIT('h8)
	) name4783 (
		_w15294_,
		_w15295_,
		_w15296_
	);
	LUT4 #(
		.INIT('h8000)
	) name4784 (
		_w15288_,
		_w15291_,
		_w15293_,
		_w15296_,
		_w15297_
	);
	LUT3 #(
		.INIT('h80)
	) name4785 (
		\wishbone_RxPointerMSB_reg[25]/NET0131 ,
		\wishbone_RxPointerMSB_reg[29]/NET0131 ,
		\wishbone_RxPointerMSB_reg[30]/NET0131 ,
		_w15298_
	);
	LUT2 #(
		.INIT('h8)
	) name4786 (
		_w15294_,
		_w15298_,
		_w15299_
	);
	LUT4 #(
		.INIT('h8000)
	) name4787 (
		_w15288_,
		_w15291_,
		_w15293_,
		_w15299_,
		_w15300_
	);
	LUT4 #(
		.INIT('h0032)
	) name4788 (
		\wishbone_RxPointerMSB_reg[30]/NET0131 ,
		_w13807_,
		_w15297_,
		_w15300_,
		_w15301_
	);
	LUT3 #(
		.INIT('hf4)
	) name4789 (
		_w13016_,
		_w15282_,
		_w15301_,
		_w15302_
	);
	LUT3 #(
		.INIT('h80)
	) name4790 (
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w15303_
	);
	LUT2 #(
		.INIT('h4)
	) name4791 (
		\wishbone_BlockingIncrementTxPointer_reg/NET0131 ,
		\wishbone_IncrTxPointer_reg/NET0131 ,
		_w15304_
	);
	LUT4 #(
		.INIT('h4000)
	) name4792 (
		\wishbone_BlockingIncrementTxPointer_reg/NET0131 ,
		\wishbone_IncrTxPointer_reg/NET0131 ,
		\wishbone_TxPointerMSB_reg[2]/NET0131 ,
		\wishbone_TxPointerMSB_reg[3]/NET0131 ,
		_w15305_
	);
	LUT3 #(
		.INIT('h80)
	) name4793 (
		\wishbone_TxPointerMSB_reg[4]/NET0131 ,
		\wishbone_TxPointerMSB_reg[5]/NET0131 ,
		\wishbone_TxPointerMSB_reg[6]/NET0131 ,
		_w15306_
	);
	LUT3 #(
		.INIT('h80)
	) name4794 (
		\wishbone_TxPointerMSB_reg[7]/NET0131 ,
		\wishbone_TxPointerMSB_reg[8]/NET0131 ,
		\wishbone_TxPointerMSB_reg[9]/NET0131 ,
		_w15307_
	);
	LUT3 #(
		.INIT('h80)
	) name4795 (
		_w15305_,
		_w15306_,
		_w15307_,
		_w15308_
	);
	LUT3 #(
		.INIT('h80)
	) name4796 (
		\wishbone_TxPointerMSB_reg[10]/NET0131 ,
		\wishbone_TxPointerMSB_reg[11]/NET0131 ,
		\wishbone_TxPointerMSB_reg[12]/NET0131 ,
		_w15309_
	);
	LUT4 #(
		.INIT('h8000)
	) name4797 (
		_w15305_,
		_w15306_,
		_w15307_,
		_w15309_,
		_w15310_
	);
	LUT2 #(
		.INIT('h8)
	) name4798 (
		\wishbone_TxPointerMSB_reg[15]/NET0131 ,
		\wishbone_TxPointerMSB_reg[16]/NET0131 ,
		_w15311_
	);
	LUT2 #(
		.INIT('h8)
	) name4799 (
		\wishbone_TxPointerMSB_reg[13]/NET0131 ,
		\wishbone_TxPointerMSB_reg[14]/NET0131 ,
		_w15312_
	);
	LUT3 #(
		.INIT('h80)
	) name4800 (
		\wishbone_TxPointerMSB_reg[13]/NET0131 ,
		\wishbone_TxPointerMSB_reg[14]/NET0131 ,
		\wishbone_TxPointerMSB_reg[17]/NET0131 ,
		_w15313_
	);
	LUT2 #(
		.INIT('h8)
	) name4801 (
		_w15311_,
		_w15313_,
		_w15314_
	);
	LUT3 #(
		.INIT('h80)
	) name4802 (
		\wishbone_TxPointerMSB_reg[18]/NET0131 ,
		\wishbone_TxPointerMSB_reg[19]/NET0131 ,
		\wishbone_TxPointerMSB_reg[20]/NET0131 ,
		_w15315_
	);
	LUT2 #(
		.INIT('h8)
	) name4803 (
		\wishbone_TxPointerMSB_reg[21]/NET0131 ,
		\wishbone_TxPointerMSB_reg[22]/NET0131 ,
		_w15316_
	);
	LUT2 #(
		.INIT('h8)
	) name4804 (
		_w15315_,
		_w15316_,
		_w15317_
	);
	LUT3 #(
		.INIT('h80)
	) name4805 (
		_w15310_,
		_w15314_,
		_w15317_,
		_w15318_
	);
	LUT2 #(
		.INIT('h8)
	) name4806 (
		\wishbone_TxPointerMSB_reg[25]/NET0131 ,
		\wishbone_TxPointerMSB_reg[26]/NET0131 ,
		_w15319_
	);
	LUT2 #(
		.INIT('h8)
	) name4807 (
		\wishbone_TxPointerMSB_reg[23]/NET0131 ,
		\wishbone_TxPointerMSB_reg[24]/NET0131 ,
		_w15320_
	);
	LUT4 #(
		.INIT('h8000)
	) name4808 (
		\wishbone_TxPointerMSB_reg[23]/NET0131 ,
		\wishbone_TxPointerMSB_reg[24]/NET0131 ,
		\wishbone_TxPointerMSB_reg[27]/NET0131 ,
		\wishbone_TxPointerMSB_reg[28]/NET0131 ,
		_w15321_
	);
	LUT2 #(
		.INIT('h8)
	) name4809 (
		_w15319_,
		_w15321_,
		_w15322_
	);
	LUT4 #(
		.INIT('h8000)
	) name4810 (
		_w15310_,
		_w15314_,
		_w15317_,
		_w15322_,
		_w15323_
	);
	LUT2 #(
		.INIT('h6)
	) name4811 (
		\wishbone_TxPointerMSB_reg[29]/NET0131 ,
		\wishbone_TxPointerMSB_reg[30]/NET0131 ,
		_w15324_
	);
	LUT2 #(
		.INIT('h1)
	) name4812 (
		_w15303_,
		_w15324_,
		_w15325_
	);
	LUT4 #(
		.INIT('h070f)
	) name4813 (
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		\wishbone_TxPointerMSB_reg[30]/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w15326_
	);
	LUT4 #(
		.INIT('h060c)
	) name4814 (
		\wishbone_TxPointerMSB_reg[29]/NET0131 ,
		\wishbone_TxPointerMSB_reg[30]/NET0131 ,
		_w15303_,
		_w15323_,
		_w15327_
	);
	LUT4 #(
		.INIT('h0415)
	) name4815 (
		wb_rst_i_pad,
		_w15323_,
		_w15325_,
		_w15326_,
		_w15328_
	);
	LUT3 #(
		.INIT('hdc)
	) name4816 (
		_w13016_,
		_w15327_,
		_w15328_,
		_w15329_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4817 (
		\wishbone_RxDataLatched1_reg[16]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w15330_
	);
	LUT4 #(
		.INIT('hfb08)
	) name4818 (
		\wishbone_RxDataLatched2_reg[16]/NET0131 ,
		_w13423_,
		_w13424_,
		_w15330_,
		_w15331_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4819 (
		\wishbone_RxDataLatched1_reg[17]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w15332_
	);
	LUT4 #(
		.INIT('hfb08)
	) name4820 (
		\wishbone_RxDataLatched2_reg[17]/NET0131 ,
		_w13423_,
		_w13424_,
		_w15332_,
		_w15333_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4821 (
		\wishbone_RxDataLatched1_reg[18]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w15334_
	);
	LUT4 #(
		.INIT('hfb08)
	) name4822 (
		\wishbone_RxDataLatched2_reg[18]/NET0131 ,
		_w13423_,
		_w13424_,
		_w15334_,
		_w15335_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4823 (
		\wishbone_RxDataLatched1_reg[19]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w15336_
	);
	LUT4 #(
		.INIT('hfb08)
	) name4824 (
		\wishbone_RxDataLatched2_reg[19]/NET0131 ,
		_w13423_,
		_w13424_,
		_w15336_,
		_w15337_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4825 (
		\wishbone_RxDataLatched1_reg[20]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w15338_
	);
	LUT4 #(
		.INIT('hfb08)
	) name4826 (
		\wishbone_RxDataLatched2_reg[20]/NET0131 ,
		_w13423_,
		_w13424_,
		_w15338_,
		_w15339_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4827 (
		\wishbone_RxDataLatched1_reg[21]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w15340_
	);
	LUT4 #(
		.INIT('hfb08)
	) name4828 (
		\wishbone_RxDataLatched2_reg[21]/NET0131 ,
		_w13423_,
		_w13424_,
		_w15340_,
		_w15341_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4829 (
		\wishbone_RxDataLatched1_reg[22]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w15342_
	);
	LUT4 #(
		.INIT('hfb08)
	) name4830 (
		\wishbone_RxDataLatched2_reg[22]/NET0131 ,
		_w13423_,
		_w13424_,
		_w15342_,
		_w15343_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4831 (
		\wishbone_RxDataLatched1_reg[23]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w15344_
	);
	LUT4 #(
		.INIT('hfb08)
	) name4832 (
		\wishbone_RxDataLatched2_reg[23]/NET0131 ,
		_w13423_,
		_w13424_,
		_w15344_,
		_w15345_
	);
	LUT4 #(
		.INIT('h0001)
	) name4833 (
		\wishbone_RxPointerMSB_reg[13]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w15346_
	);
	LUT3 #(
		.INIT('h07)
	) name4834 (
		_w11868_,
		_w11875_,
		_w15346_,
		_w15347_
	);
	LUT3 #(
		.INIT('h80)
	) name4835 (
		_w11870_,
		_w11873_,
		_w15347_,
		_w15348_
	);
	LUT2 #(
		.INIT('h8)
	) name4836 (
		\m_wb_adr_o[12]_pad ,
		\m_wb_adr_o[13]_pad ,
		_w15349_
	);
	LUT4 #(
		.INIT('h8000)
	) name4837 (
		_w11845_,
		_w11846_,
		_w11848_,
		_w15349_,
		_w15350_
	);
	LUT3 #(
		.INIT('h6c)
	) name4838 (
		\m_wb_adr_o[12]_pad ,
		\m_wb_adr_o[13]_pad ,
		_w11849_,
		_w15351_
	);
	LUT3 #(
		.INIT('he0)
	) name4839 (
		_w11887_,
		_w15348_,
		_w15351_,
		_w15352_
	);
	LUT3 #(
		.INIT('ha2)
	) name4840 (
		\wishbone_TxPointerMSB_reg[13]/NET0131 ,
		_w11900_,
		_w11909_,
		_w15353_
	);
	LUT4 #(
		.INIT('h080a)
	) name4841 (
		\wishbone_RxPointerMSB_reg[13]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w15354_
	);
	LUT3 #(
		.INIT('he0)
	) name4842 (
		_w11902_,
		_w11905_,
		_w15354_,
		_w15355_
	);
	LUT4 #(
		.INIT('h0007)
	) name4843 (
		\m_wb_adr_o[13]_pad ,
		_w11907_,
		_w15353_,
		_w15355_,
		_w15356_
	);
	LUT2 #(
		.INIT('hb)
	) name4844 (
		_w15352_,
		_w15356_,
		_w15357_
	);
	LUT3 #(
		.INIT('h80)
	) name4845 (
		\m_wb_adr_o[12]_pad ,
		\m_wb_adr_o[13]_pad ,
		\m_wb_adr_o[14]_pad ,
		_w15358_
	);
	LUT4 #(
		.INIT('h8000)
	) name4846 (
		_w11845_,
		_w11846_,
		_w11848_,
		_w15358_,
		_w15359_
	);
	LUT3 #(
		.INIT('h0e)
	) name4847 (
		\m_wb_adr_o[14]_pad ,
		_w15350_,
		_w15359_,
		_w15360_
	);
	LUT3 #(
		.INIT('he0)
	) name4848 (
		_w11887_,
		_w13051_,
		_w15360_,
		_w15361_
	);
	LUT3 #(
		.INIT('h07)
	) name4849 (
		\m_wb_adr_o[14]_pad ,
		_w11907_,
		_w15361_,
		_w15362_
	);
	LUT3 #(
		.INIT('h04)
	) name4850 (
		_w11885_,
		_w11900_,
		_w15360_,
		_w15363_
	);
	LUT3 #(
		.INIT('h8a)
	) name4851 (
		\wishbone_TxPointerMSB_reg[14]/NET0131 ,
		_w11890_,
		_w11900_,
		_w15364_
	);
	LUT2 #(
		.INIT('h1)
	) name4852 (
		_w11914_,
		_w15360_,
		_w15365_
	);
	LUT3 #(
		.INIT('ha8)
	) name4853 (
		\wishbone_RxPointerMSB_reg[14]/NET0131 ,
		_w11902_,
		_w11905_,
		_w15366_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4854 (
		_w15363_,
		_w15364_,
		_w15365_,
		_w15366_,
		_w15367_
	);
	LUT2 #(
		.INIT('h7)
	) name4855 (
		_w15362_,
		_w15367_,
		_w15368_
	);
	LUT4 #(
		.INIT('h080a)
	) name4856 (
		\wishbone_RxPointerMSB_reg[8]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w15369_
	);
	LUT3 #(
		.INIT('he0)
	) name4857 (
		_w11902_,
		_w11905_,
		_w15369_,
		_w15370_
	);
	LUT3 #(
		.INIT('h07)
	) name4858 (
		\m_wb_adr_o[8]_pad ,
		_w11907_,
		_w15370_,
		_w15371_
	);
	LUT3 #(
		.INIT('ha2)
	) name4859 (
		\wishbone_TxPointerMSB_reg[8]/NET0131 ,
		_w11900_,
		_w11909_,
		_w15372_
	);
	LUT4 #(
		.INIT('h78f0)
	) name4860 (
		\m_wb_adr_o[6]_pad ,
		\m_wb_adr_o[7]_pad ,
		\m_wb_adr_o[8]_pad ,
		_w11845_,
		_w15373_
	);
	LUT3 #(
		.INIT('he0)
	) name4861 (
		_w11887_,
		_w13051_,
		_w15373_,
		_w15374_
	);
	LUT2 #(
		.INIT('h1)
	) name4862 (
		_w15372_,
		_w15374_,
		_w15375_
	);
	LUT2 #(
		.INIT('h7)
	) name4863 (
		_w15371_,
		_w15375_,
		_w15376_
	);
	LUT4 #(
		.INIT('h0001)
	) name4864 (
		\wishbone_RxPointerMSB_reg[11]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w15377_
	);
	LUT3 #(
		.INIT('h07)
	) name4865 (
		_w11868_,
		_w11875_,
		_w15377_,
		_w15378_
	);
	LUT3 #(
		.INIT('h80)
	) name4866 (
		_w11870_,
		_w11873_,
		_w15378_,
		_w15379_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name4867 (
		\m_wb_adr_o[11]_pad ,
		_w11845_,
		_w11846_,
		_w11847_,
		_w15380_
	);
	LUT3 #(
		.INIT('he0)
	) name4868 (
		_w11887_,
		_w15379_,
		_w15380_,
		_w15381_
	);
	LUT3 #(
		.INIT('ha2)
	) name4869 (
		\wishbone_TxPointerMSB_reg[11]/NET0131 ,
		_w11900_,
		_w11909_,
		_w15382_
	);
	LUT4 #(
		.INIT('h080a)
	) name4870 (
		\wishbone_RxPointerMSB_reg[11]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w15383_
	);
	LUT3 #(
		.INIT('he0)
	) name4871 (
		_w11902_,
		_w11905_,
		_w15383_,
		_w15384_
	);
	LUT4 #(
		.INIT('h0007)
	) name4872 (
		\m_wb_adr_o[11]_pad ,
		_w11907_,
		_w15382_,
		_w15384_,
		_w15385_
	);
	LUT2 #(
		.INIT('hb)
	) name4873 (
		_w15381_,
		_w15385_,
		_w15386_
	);
	LUT4 #(
		.INIT('h80aa)
	) name4874 (
		\wishbone_TxPointerMSB_reg[15]/NET0131 ,
		_w11866_,
		_w11867_,
		_w11883_,
		_w15387_
	);
	LUT2 #(
		.INIT('h4)
	) name4875 (
		_w11882_,
		_w15387_,
		_w15388_
	);
	LUT3 #(
		.INIT('h32)
	) name4876 (
		\m_wb_adr_o[15]_pad ,
		_w11851_,
		_w15359_,
		_w15389_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4877 (
		_w11887_,
		_w13051_,
		_w15388_,
		_w15389_,
		_w15390_
	);
	LUT3 #(
		.INIT('ha2)
	) name4878 (
		\wishbone_TxPointerMSB_reg[15]/NET0131 ,
		_w11900_,
		_w11909_,
		_w15391_
	);
	LUT4 #(
		.INIT('h080a)
	) name4879 (
		\wishbone_RxPointerMSB_reg[15]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w15392_
	);
	LUT3 #(
		.INIT('he0)
	) name4880 (
		_w11902_,
		_w11905_,
		_w15392_,
		_w15393_
	);
	LUT4 #(
		.INIT('h0007)
	) name4881 (
		\m_wb_adr_o[15]_pad ,
		_w11907_,
		_w15391_,
		_w15393_,
		_w15394_
	);
	LUT2 #(
		.INIT('hb)
	) name4882 (
		_w15390_,
		_w15394_,
		_w15395_
	);
	LUT4 #(
		.INIT('h080a)
	) name4883 (
		\wishbone_RxPointerMSB_reg[4]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w15396_
	);
	LUT3 #(
		.INIT('he0)
	) name4884 (
		_w11902_,
		_w11905_,
		_w15396_,
		_w15397_
	);
	LUT3 #(
		.INIT('h07)
	) name4885 (
		\m_wb_adr_o[4]_pad ,
		_w11907_,
		_w15397_,
		_w15398_
	);
	LUT3 #(
		.INIT('ha2)
	) name4886 (
		\wishbone_TxPointerMSB_reg[4]/NET0131 ,
		_w11900_,
		_w11909_,
		_w15399_
	);
	LUT3 #(
		.INIT('h78)
	) name4887 (
		\m_wb_adr_o[2]_pad ,
		\m_wb_adr_o[3]_pad ,
		\m_wb_adr_o[4]_pad ,
		_w15400_
	);
	LUT3 #(
		.INIT('he0)
	) name4888 (
		_w11887_,
		_w13051_,
		_w15400_,
		_w15401_
	);
	LUT2 #(
		.INIT('h1)
	) name4889 (
		_w15399_,
		_w15401_,
		_w15402_
	);
	LUT2 #(
		.INIT('h7)
	) name4890 (
		_w15398_,
		_w15402_,
		_w15403_
	);
	LUT4 #(
		.INIT('h8000)
	) name4891 (
		\m_wb_adr_o[27]_pad ,
		_w11851_,
		_w11852_,
		_w11857_,
		_w15404_
	);
	LUT4 #(
		.INIT('h1555)
	) name4892 (
		\m_wb_adr_o[27]_pad ,
		_w11851_,
		_w11852_,
		_w11857_,
		_w15405_
	);
	LUT4 #(
		.INIT('h80aa)
	) name4893 (
		\wishbone_TxPointerMSB_reg[27]/NET0131 ,
		_w11866_,
		_w11867_,
		_w11883_,
		_w15406_
	);
	LUT2 #(
		.INIT('h4)
	) name4894 (
		_w11882_,
		_w15406_,
		_w15407_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name4895 (
		_w11887_,
		_w13051_,
		_w15405_,
		_w15407_,
		_w15408_
	);
	LUT2 #(
		.INIT('h4)
	) name4896 (
		_w15404_,
		_w15408_,
		_w15409_
	);
	LUT3 #(
		.INIT('ha2)
	) name4897 (
		\wishbone_TxPointerMSB_reg[27]/NET0131 ,
		_w11900_,
		_w11909_,
		_w15410_
	);
	LUT4 #(
		.INIT('h080a)
	) name4898 (
		\wishbone_RxPointerMSB_reg[27]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w15411_
	);
	LUT3 #(
		.INIT('he0)
	) name4899 (
		_w11902_,
		_w11905_,
		_w15411_,
		_w15412_
	);
	LUT4 #(
		.INIT('h0007)
	) name4900 (
		\m_wb_adr_o[27]_pad ,
		_w11907_,
		_w15410_,
		_w15412_,
		_w15413_
	);
	LUT2 #(
		.INIT('hb)
	) name4901 (
		_w15409_,
		_w15413_,
		_w15414_
	);
	LUT4 #(
		.INIT('h0001)
	) name4902 (
		\wishbone_RxPointerMSB_reg[31]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w15415_
	);
	LUT3 #(
		.INIT('h07)
	) name4903 (
		_w11868_,
		_w11875_,
		_w15415_,
		_w15416_
	);
	LUT3 #(
		.INIT('h80)
	) name4904 (
		_w11870_,
		_w11873_,
		_w15416_,
		_w15417_
	);
	LUT4 #(
		.INIT('h999f)
	) name4905 (
		\m_wb_adr_o[31]_pad ,
		_w11864_,
		_w11887_,
		_w15417_,
		_w15418_
	);
	LUT4 #(
		.INIT('h080a)
	) name4906 (
		\wishbone_RxPointerMSB_reg[31]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w15419_
	);
	LUT3 #(
		.INIT('he0)
	) name4907 (
		_w11902_,
		_w11905_,
		_w15419_,
		_w15420_
	);
	LUT3 #(
		.INIT('ha2)
	) name4908 (
		\wishbone_TxPointerMSB_reg[31]/NET0131 ,
		_w11900_,
		_w11909_,
		_w15421_
	);
	LUT4 #(
		.INIT('h0007)
	) name4909 (
		\m_wb_adr_o[31]_pad ,
		_w11907_,
		_w15420_,
		_w15421_,
		_w15422_
	);
	LUT2 #(
		.INIT('h7)
	) name4910 (
		_w15418_,
		_w15422_,
		_w15423_
	);
	LUT2 #(
		.INIT('h4)
	) name4911 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		_w15424_
	);
	LUT4 #(
		.INIT('h0222)
	) name4912 (
		\maccontrol1_receivecontrol1_TypeLengthOK_reg/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w11486_,
		_w15424_,
		_w15425_
	);
	LUT2 #(
		.INIT('h4)
	) name4913 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w15426_
	);
	LUT4 #(
		.INIT('h0200)
	) name4914 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w15427_
	);
	LUT3 #(
		.INIT('h80)
	) name4915 (
		_w11455_,
		_w11456_,
		_w15427_,
		_w15428_
	);
	LUT3 #(
		.INIT('h80)
	) name4916 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_receivecontrol1_TypeLengthOK_reg/NET0131 ,
		_w11486_,
		_w15429_
	);
	LUT3 #(
		.INIT('h15)
	) name4917 (
		_w15425_,
		_w15428_,
		_w15429_,
		_w15430_
	);
	LUT4 #(
		.INIT('h0001)
	) name4918 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w15431_
	);
	LUT3 #(
		.INIT('h80)
	) name4919 (
		_w11469_,
		_w15426_,
		_w15431_,
		_w15432_
	);
	LUT2 #(
		.INIT('h8)
	) name4920 (
		_w11924_,
		_w15432_,
		_w15433_
	);
	LUT2 #(
		.INIT('hd)
	) name4921 (
		_w15430_,
		_w15433_,
		_w15434_
	);
	LUT3 #(
		.INIT('h80)
	) name4922 (
		\wishbone_bd_ram_mem2_reg[85][18]/P0001 ,
		_w11933_,
		_w11972_,
		_w15435_
	);
	LUT3 #(
		.INIT('h80)
	) name4923 (
		\wishbone_bd_ram_mem2_reg[106][18]/P0001 ,
		_w11944_,
		_w11965_,
		_w15436_
	);
	LUT3 #(
		.INIT('h80)
	) name4924 (
		\wishbone_bd_ram_mem2_reg[197][18]/P0001 ,
		_w11933_,
		_w11945_,
		_w15437_
	);
	LUT3 #(
		.INIT('h80)
	) name4925 (
		\wishbone_bd_ram_mem2_reg[176][18]/P0001 ,
		_w11941_,
		_w11942_,
		_w15438_
	);
	LUT4 #(
		.INIT('h0001)
	) name4926 (
		_w15435_,
		_w15436_,
		_w15437_,
		_w15438_,
		_w15439_
	);
	LUT3 #(
		.INIT('h80)
	) name4927 (
		\wishbone_bd_ram_mem2_reg[221][18]/P0001 ,
		_w11966_,
		_w11984_,
		_w15440_
	);
	LUT3 #(
		.INIT('h80)
	) name4928 (
		\wishbone_bd_ram_mem2_reg[55][18]/P0001 ,
		_w11975_,
		_w11979_,
		_w15441_
	);
	LUT3 #(
		.INIT('h80)
	) name4929 (
		\wishbone_bd_ram_mem2_reg[102][18]/P0001 ,
		_w11965_,
		_w11986_,
		_w15442_
	);
	LUT3 #(
		.INIT('h80)
	) name4930 (
		\wishbone_bd_ram_mem2_reg[157][18]/P0001 ,
		_w11959_,
		_w11966_,
		_w15443_
	);
	LUT4 #(
		.INIT('h0001)
	) name4931 (
		_w15440_,
		_w15441_,
		_w15442_,
		_w15443_,
		_w15444_
	);
	LUT3 #(
		.INIT('h80)
	) name4932 (
		\wishbone_bd_ram_mem2_reg[7][18]/P0001 ,
		_w11932_,
		_w11975_,
		_w15445_
	);
	LUT3 #(
		.INIT('h80)
	) name4933 (
		\wishbone_bd_ram_mem2_reg[3][18]/P0001 ,
		_w11932_,
		_w11938_,
		_w15446_
	);
	LUT3 #(
		.INIT('h80)
	) name4934 (
		\wishbone_bd_ram_mem2_reg[191][18]/P0001 ,
		_w11942_,
		_w11973_,
		_w15447_
	);
	LUT3 #(
		.INIT('h80)
	) name4935 (
		\wishbone_bd_ram_mem2_reg[254][18]/P0001 ,
		_w11948_,
		_w11952_,
		_w15448_
	);
	LUT4 #(
		.INIT('h0001)
	) name4936 (
		_w15445_,
		_w15446_,
		_w15447_,
		_w15448_,
		_w15449_
	);
	LUT3 #(
		.INIT('h80)
	) name4937 (
		\wishbone_bd_ram_mem2_reg[6][18]/P0001 ,
		_w11932_,
		_w11986_,
		_w15450_
	);
	LUT3 #(
		.INIT('h80)
	) name4938 (
		\wishbone_bd_ram_mem2_reg[222][18]/P0001 ,
		_w11948_,
		_w11984_,
		_w15451_
	);
	LUT3 #(
		.INIT('h80)
	) name4939 (
		\wishbone_bd_ram_mem2_reg[32][18]/P0001 ,
		_w11941_,
		_w11957_,
		_w15452_
	);
	LUT3 #(
		.INIT('h80)
	) name4940 (
		\wishbone_bd_ram_mem2_reg[119][18]/P0001 ,
		_w11975_,
		_w12012_,
		_w15453_
	);
	LUT4 #(
		.INIT('h0001)
	) name4941 (
		_w15450_,
		_w15451_,
		_w15452_,
		_w15453_,
		_w15454_
	);
	LUT4 #(
		.INIT('h8000)
	) name4942 (
		_w15439_,
		_w15444_,
		_w15449_,
		_w15454_,
		_w15455_
	);
	LUT3 #(
		.INIT('h80)
	) name4943 (
		\wishbone_bd_ram_mem2_reg[40][18]/P0001 ,
		_w11957_,
		_w11990_,
		_w15456_
	);
	LUT3 #(
		.INIT('h80)
	) name4944 (
		\wishbone_bd_ram_mem2_reg[42][18]/P0001 ,
		_w11944_,
		_w11957_,
		_w15457_
	);
	LUT3 #(
		.INIT('h80)
	) name4945 (
		\wishbone_bd_ram_mem2_reg[179][18]/P0001 ,
		_w11938_,
		_w11942_,
		_w15458_
	);
	LUT3 #(
		.INIT('h80)
	) name4946 (
		\wishbone_bd_ram_mem2_reg[210][18]/P0001 ,
		_w11963_,
		_w11984_,
		_w15459_
	);
	LUT4 #(
		.INIT('h0001)
	) name4947 (
		_w15456_,
		_w15457_,
		_w15458_,
		_w15459_,
		_w15460_
	);
	LUT3 #(
		.INIT('h80)
	) name4948 (
		\wishbone_bd_ram_mem2_reg[14][18]/P0001 ,
		_w11932_,
		_w11948_,
		_w15461_
	);
	LUT3 #(
		.INIT('h80)
	) name4949 (
		\wishbone_bd_ram_mem2_reg[61][18]/P0001 ,
		_w11966_,
		_w11979_,
		_w15462_
	);
	LUT3 #(
		.INIT('h80)
	) name4950 (
		\wishbone_bd_ram_mem2_reg[234][18]/P0001 ,
		_w11944_,
		_w11982_,
		_w15463_
	);
	LUT3 #(
		.INIT('h80)
	) name4951 (
		\wishbone_bd_ram_mem2_reg[4][18]/P0001 ,
		_w11929_,
		_w11932_,
		_w15464_
	);
	LUT4 #(
		.INIT('h0001)
	) name4952 (
		_w15461_,
		_w15462_,
		_w15463_,
		_w15464_,
		_w15465_
	);
	LUT3 #(
		.INIT('h80)
	) name4953 (
		\wishbone_bd_ram_mem2_reg[80][18]/P0001 ,
		_w11941_,
		_w11972_,
		_w15466_
	);
	LUT3 #(
		.INIT('h80)
	) name4954 (
		\wishbone_bd_ram_mem2_reg[99][18]/P0001 ,
		_w11938_,
		_w11965_,
		_w15467_
	);
	LUT3 #(
		.INIT('h80)
	) name4955 (
		\wishbone_bd_ram_mem2_reg[159][18]/P0001 ,
		_w11959_,
		_w11973_,
		_w15468_
	);
	LUT3 #(
		.INIT('h80)
	) name4956 (
		\wishbone_bd_ram_mem2_reg[107][18]/P0001 ,
		_w11936_,
		_w11965_,
		_w15469_
	);
	LUT4 #(
		.INIT('h0001)
	) name4957 (
		_w15466_,
		_w15467_,
		_w15468_,
		_w15469_,
		_w15470_
	);
	LUT3 #(
		.INIT('h80)
	) name4958 (
		\wishbone_bd_ram_mem2_reg[146][18]/P0001 ,
		_w11959_,
		_w11963_,
		_w15471_
	);
	LUT3 #(
		.INIT('h80)
	) name4959 (
		\wishbone_bd_ram_mem2_reg[65][18]/P0001 ,
		_w11949_,
		_w11977_,
		_w15472_
	);
	LUT3 #(
		.INIT('h80)
	) name4960 (
		\wishbone_bd_ram_mem2_reg[13][18]/P0001 ,
		_w11932_,
		_w11966_,
		_w15473_
	);
	LUT3 #(
		.INIT('h80)
	) name4961 (
		\wishbone_bd_ram_mem2_reg[10][18]/P0001 ,
		_w11932_,
		_w11944_,
		_w15474_
	);
	LUT4 #(
		.INIT('h0001)
	) name4962 (
		_w15471_,
		_w15472_,
		_w15473_,
		_w15474_,
		_w15475_
	);
	LUT4 #(
		.INIT('h8000)
	) name4963 (
		_w15460_,
		_w15465_,
		_w15470_,
		_w15475_,
		_w15476_
	);
	LUT3 #(
		.INIT('h80)
	) name4964 (
		\wishbone_bd_ram_mem2_reg[12][18]/P0001 ,
		_w11932_,
		_w11954_,
		_w15477_
	);
	LUT3 #(
		.INIT('h80)
	) name4965 (
		\wishbone_bd_ram_mem2_reg[184][18]/P0001 ,
		_w11942_,
		_w11990_,
		_w15478_
	);
	LUT3 #(
		.INIT('h80)
	) name4966 (
		\wishbone_bd_ram_mem2_reg[82][18]/P0001 ,
		_w11963_,
		_w11972_,
		_w15479_
	);
	LUT3 #(
		.INIT('h80)
	) name4967 (
		\wishbone_bd_ram_mem2_reg[174][18]/P0001 ,
		_w11930_,
		_w11948_,
		_w15480_
	);
	LUT4 #(
		.INIT('h0001)
	) name4968 (
		_w15477_,
		_w15478_,
		_w15479_,
		_w15480_,
		_w15481_
	);
	LUT3 #(
		.INIT('h80)
	) name4969 (
		\wishbone_bd_ram_mem2_reg[79][18]/P0001 ,
		_w11949_,
		_w11973_,
		_w15482_
	);
	LUT3 #(
		.INIT('h80)
	) name4970 (
		\wishbone_bd_ram_mem2_reg[90][18]/P0001 ,
		_w11944_,
		_w11972_,
		_w15483_
	);
	LUT3 #(
		.INIT('h80)
	) name4971 (
		\wishbone_bd_ram_mem2_reg[45][18]/P0001 ,
		_w11957_,
		_w11966_,
		_w15484_
	);
	LUT3 #(
		.INIT('h80)
	) name4972 (
		\wishbone_bd_ram_mem2_reg[128][18]/P0001 ,
		_w11941_,
		_w11955_,
		_w15485_
	);
	LUT4 #(
		.INIT('h0001)
	) name4973 (
		_w15482_,
		_w15483_,
		_w15484_,
		_w15485_,
		_w15486_
	);
	LUT3 #(
		.INIT('h80)
	) name4974 (
		\wishbone_bd_ram_mem2_reg[84][18]/P0001 ,
		_w11929_,
		_w11972_,
		_w15487_
	);
	LUT3 #(
		.INIT('h80)
	) name4975 (
		\wishbone_bd_ram_mem2_reg[193][18]/P0001 ,
		_w11945_,
		_w11977_,
		_w15488_
	);
	LUT3 #(
		.INIT('h80)
	) name4976 (
		\wishbone_bd_ram_mem2_reg[241][18]/P0001 ,
		_w11952_,
		_w11977_,
		_w15489_
	);
	LUT3 #(
		.INIT('h80)
	) name4977 (
		\wishbone_bd_ram_mem2_reg[138][18]/P0001 ,
		_w11944_,
		_w11955_,
		_w15490_
	);
	LUT4 #(
		.INIT('h0001)
	) name4978 (
		_w15487_,
		_w15488_,
		_w15489_,
		_w15490_,
		_w15491_
	);
	LUT3 #(
		.INIT('h80)
	) name4979 (
		\wishbone_bd_ram_mem2_reg[11][18]/P0001 ,
		_w11932_,
		_w11936_,
		_w15492_
	);
	LUT3 #(
		.INIT('h80)
	) name4980 (
		\wishbone_bd_ram_mem2_reg[218][18]/P0001 ,
		_w11944_,
		_w11984_,
		_w15493_
	);
	LUT3 #(
		.INIT('h80)
	) name4981 (
		\wishbone_bd_ram_mem2_reg[126][18]/P0001 ,
		_w11948_,
		_w12012_,
		_w15494_
	);
	LUT3 #(
		.INIT('h80)
	) name4982 (
		\wishbone_bd_ram_mem2_reg[115][18]/P0001 ,
		_w11938_,
		_w12012_,
		_w15495_
	);
	LUT4 #(
		.INIT('h0001)
	) name4983 (
		_w15492_,
		_w15493_,
		_w15494_,
		_w15495_,
		_w15496_
	);
	LUT4 #(
		.INIT('h8000)
	) name4984 (
		_w15481_,
		_w15486_,
		_w15491_,
		_w15496_,
		_w15497_
	);
	LUT3 #(
		.INIT('h80)
	) name4985 (
		\wishbone_bd_ram_mem2_reg[195][18]/P0001 ,
		_w11938_,
		_w11945_,
		_w15498_
	);
	LUT3 #(
		.INIT('h80)
	) name4986 (
		\wishbone_bd_ram_mem2_reg[103][18]/P0001 ,
		_w11965_,
		_w11975_,
		_w15499_
	);
	LUT3 #(
		.INIT('h80)
	) name4987 (
		\wishbone_bd_ram_mem2_reg[86][18]/P0001 ,
		_w11972_,
		_w11986_,
		_w15500_
	);
	LUT3 #(
		.INIT('h80)
	) name4988 (
		\wishbone_bd_ram_mem2_reg[170][18]/P0001 ,
		_w11930_,
		_w11944_,
		_w15501_
	);
	LUT4 #(
		.INIT('h0001)
	) name4989 (
		_w15498_,
		_w15499_,
		_w15500_,
		_w15501_,
		_w15502_
	);
	LUT3 #(
		.INIT('h80)
	) name4990 (
		\wishbone_bd_ram_mem2_reg[48][18]/P0001 ,
		_w11941_,
		_w11979_,
		_w15503_
	);
	LUT3 #(
		.INIT('h80)
	) name4991 (
		\wishbone_bd_ram_mem2_reg[43][18]/P0001 ,
		_w11936_,
		_w11957_,
		_w15504_
	);
	LUT3 #(
		.INIT('h80)
	) name4992 (
		\wishbone_bd_ram_mem2_reg[230][18]/P0001 ,
		_w11982_,
		_w11986_,
		_w15505_
	);
	LUT3 #(
		.INIT('h80)
	) name4993 (
		\wishbone_bd_ram_mem2_reg[242][18]/P0001 ,
		_w11952_,
		_w11963_,
		_w15506_
	);
	LUT4 #(
		.INIT('h0001)
	) name4994 (
		_w15503_,
		_w15504_,
		_w15505_,
		_w15506_,
		_w15507_
	);
	LUT3 #(
		.INIT('h80)
	) name4995 (
		\wishbone_bd_ram_mem2_reg[178][18]/P0001 ,
		_w11942_,
		_w11963_,
		_w15508_
	);
	LUT3 #(
		.INIT('h80)
	) name4996 (
		\wishbone_bd_ram_mem2_reg[29][18]/P0001 ,
		_w11935_,
		_w11966_,
		_w15509_
	);
	LUT3 #(
		.INIT('h80)
	) name4997 (
		\wishbone_bd_ram_mem2_reg[229][18]/P0001 ,
		_w11933_,
		_w11982_,
		_w15510_
	);
	LUT3 #(
		.INIT('h80)
	) name4998 (
		\wishbone_bd_ram_mem2_reg[130][18]/P0001 ,
		_w11955_,
		_w11963_,
		_w15511_
	);
	LUT4 #(
		.INIT('h0001)
	) name4999 (
		_w15508_,
		_w15509_,
		_w15510_,
		_w15511_,
		_w15512_
	);
	LUT3 #(
		.INIT('h80)
	) name5000 (
		\wishbone_bd_ram_mem2_reg[251][18]/P0001 ,
		_w11936_,
		_w11952_,
		_w15513_
	);
	LUT3 #(
		.INIT('h80)
	) name5001 (
		\wishbone_bd_ram_mem2_reg[206][18]/P0001 ,
		_w11945_,
		_w11948_,
		_w15514_
	);
	LUT3 #(
		.INIT('h80)
	) name5002 (
		\wishbone_bd_ram_mem2_reg[224][18]/P0001 ,
		_w11941_,
		_w11982_,
		_w15515_
	);
	LUT3 #(
		.INIT('h80)
	) name5003 (
		\wishbone_bd_ram_mem2_reg[185][18]/P0001 ,
		_w11942_,
		_w11968_,
		_w15516_
	);
	LUT4 #(
		.INIT('h0001)
	) name5004 (
		_w15513_,
		_w15514_,
		_w15515_,
		_w15516_,
		_w15517_
	);
	LUT4 #(
		.INIT('h8000)
	) name5005 (
		_w15502_,
		_w15507_,
		_w15512_,
		_w15517_,
		_w15518_
	);
	LUT4 #(
		.INIT('h8000)
	) name5006 (
		_w15455_,
		_w15476_,
		_w15497_,
		_w15518_,
		_w15519_
	);
	LUT3 #(
		.INIT('h80)
	) name5007 (
		\wishbone_bd_ram_mem2_reg[16][18]/P0001 ,
		_w11935_,
		_w11941_,
		_w15520_
	);
	LUT3 #(
		.INIT('h80)
	) name5008 (
		\wishbone_bd_ram_mem2_reg[167][18]/P0001 ,
		_w11930_,
		_w11975_,
		_w15521_
	);
	LUT3 #(
		.INIT('h80)
	) name5009 (
		\wishbone_bd_ram_mem2_reg[120][18]/P0001 ,
		_w11990_,
		_w12012_,
		_w15522_
	);
	LUT3 #(
		.INIT('h80)
	) name5010 (
		\wishbone_bd_ram_mem2_reg[247][18]/P0001 ,
		_w11952_,
		_w11975_,
		_w15523_
	);
	LUT4 #(
		.INIT('h0001)
	) name5011 (
		_w15520_,
		_w15521_,
		_w15522_,
		_w15523_,
		_w15524_
	);
	LUT3 #(
		.INIT('h80)
	) name5012 (
		\wishbone_bd_ram_mem2_reg[113][18]/P0001 ,
		_w11977_,
		_w12012_,
		_w15525_
	);
	LUT3 #(
		.INIT('h80)
	) name5013 (
		\wishbone_bd_ram_mem2_reg[134][18]/P0001 ,
		_w11955_,
		_w11986_,
		_w15526_
	);
	LUT3 #(
		.INIT('h80)
	) name5014 (
		\wishbone_bd_ram_mem2_reg[47][18]/P0001 ,
		_w11957_,
		_w11973_,
		_w15527_
	);
	LUT3 #(
		.INIT('h80)
	) name5015 (
		\wishbone_bd_ram_mem2_reg[153][18]/P0001 ,
		_w11959_,
		_w11968_,
		_w15528_
	);
	LUT4 #(
		.INIT('h0001)
	) name5016 (
		_w15525_,
		_w15526_,
		_w15527_,
		_w15528_,
		_w15529_
	);
	LUT3 #(
		.INIT('h80)
	) name5017 (
		\wishbone_bd_ram_mem2_reg[216][18]/P0001 ,
		_w11984_,
		_w11990_,
		_w15530_
	);
	LUT3 #(
		.INIT('h80)
	) name5018 (
		\wishbone_bd_ram_mem2_reg[238][18]/P0001 ,
		_w11948_,
		_w11982_,
		_w15531_
	);
	LUT3 #(
		.INIT('h80)
	) name5019 (
		\wishbone_bd_ram_mem2_reg[87][18]/P0001 ,
		_w11972_,
		_w11975_,
		_w15532_
	);
	LUT3 #(
		.INIT('h80)
	) name5020 (
		\wishbone_bd_ram_mem2_reg[38][18]/P0001 ,
		_w11957_,
		_w11986_,
		_w15533_
	);
	LUT4 #(
		.INIT('h0001)
	) name5021 (
		_w15530_,
		_w15531_,
		_w15532_,
		_w15533_,
		_w15534_
	);
	LUT3 #(
		.INIT('h80)
	) name5022 (
		\wishbone_bd_ram_mem2_reg[75][18]/P0001 ,
		_w11936_,
		_w11949_,
		_w15535_
	);
	LUT3 #(
		.INIT('h80)
	) name5023 (
		\wishbone_bd_ram_mem2_reg[39][18]/P0001 ,
		_w11957_,
		_w11975_,
		_w15536_
	);
	LUT3 #(
		.INIT('h80)
	) name5024 (
		\wishbone_bd_ram_mem2_reg[2][18]/P0001 ,
		_w11932_,
		_w11963_,
		_w15537_
	);
	LUT3 #(
		.INIT('h80)
	) name5025 (
		\wishbone_bd_ram_mem2_reg[111][18]/P0001 ,
		_w11965_,
		_w11973_,
		_w15538_
	);
	LUT4 #(
		.INIT('h0001)
	) name5026 (
		_w15535_,
		_w15536_,
		_w15537_,
		_w15538_,
		_w15539_
	);
	LUT4 #(
		.INIT('h8000)
	) name5027 (
		_w15524_,
		_w15529_,
		_w15534_,
		_w15539_,
		_w15540_
	);
	LUT3 #(
		.INIT('h80)
	) name5028 (
		\wishbone_bd_ram_mem2_reg[156][18]/P0001 ,
		_w11954_,
		_w11959_,
		_w15541_
	);
	LUT3 #(
		.INIT('h80)
	) name5029 (
		\wishbone_bd_ram_mem2_reg[37][18]/P0001 ,
		_w11933_,
		_w11957_,
		_w15542_
	);
	LUT3 #(
		.INIT('h80)
	) name5030 (
		\wishbone_bd_ram_mem2_reg[88][18]/P0001 ,
		_w11972_,
		_w11990_,
		_w15543_
	);
	LUT3 #(
		.INIT('h80)
	) name5031 (
		\wishbone_bd_ram_mem2_reg[252][18]/P0001 ,
		_w11952_,
		_w11954_,
		_w15544_
	);
	LUT4 #(
		.INIT('h0001)
	) name5032 (
		_w15541_,
		_w15542_,
		_w15543_,
		_w15544_,
		_w15545_
	);
	LUT3 #(
		.INIT('h80)
	) name5033 (
		\wishbone_bd_ram_mem2_reg[211][18]/P0001 ,
		_w11938_,
		_w11984_,
		_w15546_
	);
	LUT3 #(
		.INIT('h80)
	) name5034 (
		\wishbone_bd_ram_mem2_reg[200][18]/P0001 ,
		_w11945_,
		_w11990_,
		_w15547_
	);
	LUT3 #(
		.INIT('h80)
	) name5035 (
		\wishbone_bd_ram_mem2_reg[96][18]/P0001 ,
		_w11941_,
		_w11965_,
		_w15548_
	);
	LUT3 #(
		.INIT('h80)
	) name5036 (
		\wishbone_bd_ram_mem2_reg[5][18]/P0001 ,
		_w11932_,
		_w11933_,
		_w15549_
	);
	LUT4 #(
		.INIT('h0001)
	) name5037 (
		_w15546_,
		_w15547_,
		_w15548_,
		_w15549_,
		_w15550_
	);
	LUT3 #(
		.INIT('h80)
	) name5038 (
		\wishbone_bd_ram_mem2_reg[68][18]/P0001 ,
		_w11929_,
		_w11949_,
		_w15551_
	);
	LUT3 #(
		.INIT('h80)
	) name5039 (
		\wishbone_bd_ram_mem2_reg[76][18]/P0001 ,
		_w11949_,
		_w11954_,
		_w15552_
	);
	LUT3 #(
		.INIT('h80)
	) name5040 (
		\wishbone_bd_ram_mem2_reg[125][18]/P0001 ,
		_w11966_,
		_w12012_,
		_w15553_
	);
	LUT3 #(
		.INIT('h80)
	) name5041 (
		\wishbone_bd_ram_mem2_reg[163][18]/P0001 ,
		_w11930_,
		_w11938_,
		_w15554_
	);
	LUT4 #(
		.INIT('h0001)
	) name5042 (
		_w15551_,
		_w15552_,
		_w15553_,
		_w15554_,
		_w15555_
	);
	LUT3 #(
		.INIT('h80)
	) name5043 (
		\wishbone_bd_ram_mem2_reg[95][18]/P0001 ,
		_w11972_,
		_w11973_,
		_w15556_
	);
	LUT3 #(
		.INIT('h80)
	) name5044 (
		\wishbone_bd_ram_mem2_reg[101][18]/P0001 ,
		_w11933_,
		_w11965_,
		_w15557_
	);
	LUT3 #(
		.INIT('h80)
	) name5045 (
		\wishbone_bd_ram_mem2_reg[89][18]/P0001 ,
		_w11968_,
		_w11972_,
		_w15558_
	);
	LUT3 #(
		.INIT('h80)
	) name5046 (
		\wishbone_bd_ram_mem2_reg[172][18]/P0001 ,
		_w11930_,
		_w11954_,
		_w15559_
	);
	LUT4 #(
		.INIT('h0001)
	) name5047 (
		_w15556_,
		_w15557_,
		_w15558_,
		_w15559_,
		_w15560_
	);
	LUT4 #(
		.INIT('h8000)
	) name5048 (
		_w15545_,
		_w15550_,
		_w15555_,
		_w15560_,
		_w15561_
	);
	LUT3 #(
		.INIT('h80)
	) name5049 (
		\wishbone_bd_ram_mem2_reg[41][18]/P0001 ,
		_w11957_,
		_w11968_,
		_w15562_
	);
	LUT3 #(
		.INIT('h80)
	) name5050 (
		\wishbone_bd_ram_mem2_reg[97][18]/P0001 ,
		_w11965_,
		_w11977_,
		_w15563_
	);
	LUT3 #(
		.INIT('h80)
	) name5051 (
		\wishbone_bd_ram_mem2_reg[160][18]/P0001 ,
		_w11930_,
		_w11941_,
		_w15564_
	);
	LUT3 #(
		.INIT('h80)
	) name5052 (
		\wishbone_bd_ram_mem2_reg[0][18]/P0001 ,
		_w11932_,
		_w11941_,
		_w15565_
	);
	LUT4 #(
		.INIT('h0001)
	) name5053 (
		_w15562_,
		_w15563_,
		_w15564_,
		_w15565_,
		_w15566_
	);
	LUT3 #(
		.INIT('h80)
	) name5054 (
		\wishbone_bd_ram_mem2_reg[114][18]/P0001 ,
		_w11963_,
		_w12012_,
		_w15567_
	);
	LUT3 #(
		.INIT('h80)
	) name5055 (
		\wishbone_bd_ram_mem2_reg[91][18]/P0001 ,
		_w11936_,
		_w11972_,
		_w15568_
	);
	LUT3 #(
		.INIT('h80)
	) name5056 (
		\wishbone_bd_ram_mem2_reg[151][18]/P0001 ,
		_w11959_,
		_w11975_,
		_w15569_
	);
	LUT3 #(
		.INIT('h80)
	) name5057 (
		\wishbone_bd_ram_mem2_reg[244][18]/P0001 ,
		_w11929_,
		_w11952_,
		_w15570_
	);
	LUT4 #(
		.INIT('h0001)
	) name5058 (
		_w15567_,
		_w15568_,
		_w15569_,
		_w15570_,
		_w15571_
	);
	LUT3 #(
		.INIT('h80)
	) name5059 (
		\wishbone_bd_ram_mem2_reg[208][18]/P0001 ,
		_w11941_,
		_w11984_,
		_w15572_
	);
	LUT3 #(
		.INIT('h80)
	) name5060 (
		\wishbone_bd_ram_mem2_reg[121][18]/P0001 ,
		_w11968_,
		_w12012_,
		_w15573_
	);
	LUT3 #(
		.INIT('h80)
	) name5061 (
		\wishbone_bd_ram_mem2_reg[187][18]/P0001 ,
		_w11936_,
		_w11942_,
		_w15574_
	);
	LUT3 #(
		.INIT('h80)
	) name5062 (
		\wishbone_bd_ram_mem2_reg[131][18]/P0001 ,
		_w11938_,
		_w11955_,
		_w15575_
	);
	LUT4 #(
		.INIT('h0001)
	) name5063 (
		_w15572_,
		_w15573_,
		_w15574_,
		_w15575_,
		_w15576_
	);
	LUT3 #(
		.INIT('h80)
	) name5064 (
		\wishbone_bd_ram_mem2_reg[9][18]/P0001 ,
		_w11932_,
		_w11968_,
		_w15577_
	);
	LUT3 #(
		.INIT('h80)
	) name5065 (
		\wishbone_bd_ram_mem2_reg[25][18]/P0001 ,
		_w11935_,
		_w11968_,
		_w15578_
	);
	LUT3 #(
		.INIT('h80)
	) name5066 (
		\wishbone_bd_ram_mem2_reg[201][18]/P0001 ,
		_w11945_,
		_w11968_,
		_w15579_
	);
	LUT3 #(
		.INIT('h80)
	) name5067 (
		\wishbone_bd_ram_mem2_reg[250][18]/P0001 ,
		_w11944_,
		_w11952_,
		_w15580_
	);
	LUT4 #(
		.INIT('h0001)
	) name5068 (
		_w15577_,
		_w15578_,
		_w15579_,
		_w15580_,
		_w15581_
	);
	LUT4 #(
		.INIT('h8000)
	) name5069 (
		_w15566_,
		_w15571_,
		_w15576_,
		_w15581_,
		_w15582_
	);
	LUT3 #(
		.INIT('h80)
	) name5070 (
		\wishbone_bd_ram_mem2_reg[20][18]/P0001 ,
		_w11929_,
		_w11935_,
		_w15583_
	);
	LUT3 #(
		.INIT('h80)
	) name5071 (
		\wishbone_bd_ram_mem2_reg[123][18]/P0001 ,
		_w11936_,
		_w12012_,
		_w15584_
	);
	LUT3 #(
		.INIT('h80)
	) name5072 (
		\wishbone_bd_ram_mem2_reg[122][18]/P0001 ,
		_w11944_,
		_w12012_,
		_w15585_
	);
	LUT3 #(
		.INIT('h80)
	) name5073 (
		\wishbone_bd_ram_mem2_reg[162][18]/P0001 ,
		_w11930_,
		_w11963_,
		_w15586_
	);
	LUT4 #(
		.INIT('h0001)
	) name5074 (
		_w15583_,
		_w15584_,
		_w15585_,
		_w15586_,
		_w15587_
	);
	LUT3 #(
		.INIT('h80)
	) name5075 (
		\wishbone_bd_ram_mem2_reg[232][18]/P0001 ,
		_w11982_,
		_w11990_,
		_w15588_
	);
	LUT3 #(
		.INIT('h80)
	) name5076 (
		\wishbone_bd_ram_mem2_reg[70][18]/P0001 ,
		_w11949_,
		_w11986_,
		_w15589_
	);
	LUT3 #(
		.INIT('h80)
	) name5077 (
		\wishbone_bd_ram_mem2_reg[59][18]/P0001 ,
		_w11936_,
		_w11979_,
		_w15590_
	);
	LUT3 #(
		.INIT('h80)
	) name5078 (
		\wishbone_bd_ram_mem2_reg[169][18]/P0001 ,
		_w11930_,
		_w11968_,
		_w15591_
	);
	LUT4 #(
		.INIT('h0001)
	) name5079 (
		_w15588_,
		_w15589_,
		_w15590_,
		_w15591_,
		_w15592_
	);
	LUT3 #(
		.INIT('h80)
	) name5080 (
		\wishbone_bd_ram_mem2_reg[149][18]/P0001 ,
		_w11933_,
		_w11959_,
		_w15593_
	);
	LUT3 #(
		.INIT('h80)
	) name5081 (
		\wishbone_bd_ram_mem2_reg[100][18]/P0001 ,
		_w11929_,
		_w11965_,
		_w15594_
	);
	LUT3 #(
		.INIT('h80)
	) name5082 (
		\wishbone_bd_ram_mem2_reg[226][18]/P0001 ,
		_w11963_,
		_w11982_,
		_w15595_
	);
	LUT3 #(
		.INIT('h80)
	) name5083 (
		\wishbone_bd_ram_mem2_reg[196][18]/P0001 ,
		_w11929_,
		_w11945_,
		_w15596_
	);
	LUT4 #(
		.INIT('h0001)
	) name5084 (
		_w15593_,
		_w15594_,
		_w15595_,
		_w15596_,
		_w15597_
	);
	LUT3 #(
		.INIT('h80)
	) name5085 (
		\wishbone_bd_ram_mem2_reg[34][18]/P0001 ,
		_w11957_,
		_w11963_,
		_w15598_
	);
	LUT3 #(
		.INIT('h80)
	) name5086 (
		\wishbone_bd_ram_mem2_reg[207][18]/P0001 ,
		_w11945_,
		_w11973_,
		_w15599_
	);
	LUT3 #(
		.INIT('h80)
	) name5087 (
		\wishbone_bd_ram_mem2_reg[127][18]/P0001 ,
		_w11973_,
		_w12012_,
		_w15600_
	);
	LUT3 #(
		.INIT('h80)
	) name5088 (
		\wishbone_bd_ram_mem2_reg[166][18]/P0001 ,
		_w11930_,
		_w11986_,
		_w15601_
	);
	LUT4 #(
		.INIT('h0001)
	) name5089 (
		_w15598_,
		_w15599_,
		_w15600_,
		_w15601_,
		_w15602_
	);
	LUT4 #(
		.INIT('h8000)
	) name5090 (
		_w15587_,
		_w15592_,
		_w15597_,
		_w15602_,
		_w15603_
	);
	LUT4 #(
		.INIT('h8000)
	) name5091 (
		_w15540_,
		_w15561_,
		_w15582_,
		_w15603_,
		_w15604_
	);
	LUT3 #(
		.INIT('h80)
	) name5092 (
		\wishbone_bd_ram_mem2_reg[1][18]/P0001 ,
		_w11932_,
		_w11977_,
		_w15605_
	);
	LUT3 #(
		.INIT('h80)
	) name5093 (
		\wishbone_bd_ram_mem2_reg[33][18]/P0001 ,
		_w11957_,
		_w11977_,
		_w15606_
	);
	LUT3 #(
		.INIT('h80)
	) name5094 (
		\wishbone_bd_ram_mem2_reg[23][18]/P0001 ,
		_w11935_,
		_w11975_,
		_w15607_
	);
	LUT3 #(
		.INIT('h80)
	) name5095 (
		\wishbone_bd_ram_mem2_reg[155][18]/P0001 ,
		_w11936_,
		_w11959_,
		_w15608_
	);
	LUT4 #(
		.INIT('h0001)
	) name5096 (
		_w15605_,
		_w15606_,
		_w15607_,
		_w15608_,
		_w15609_
	);
	LUT3 #(
		.INIT('h80)
	) name5097 (
		\wishbone_bd_ram_mem2_reg[108][18]/P0001 ,
		_w11954_,
		_w11965_,
		_w15610_
	);
	LUT3 #(
		.INIT('h80)
	) name5098 (
		\wishbone_bd_ram_mem2_reg[50][18]/P0001 ,
		_w11963_,
		_w11979_,
		_w15611_
	);
	LUT3 #(
		.INIT('h80)
	) name5099 (
		\wishbone_bd_ram_mem2_reg[139][18]/P0001 ,
		_w11936_,
		_w11955_,
		_w15612_
	);
	LUT3 #(
		.INIT('h80)
	) name5100 (
		\wishbone_bd_ram_mem2_reg[132][18]/P0001 ,
		_w11929_,
		_w11955_,
		_w15613_
	);
	LUT4 #(
		.INIT('h0001)
	) name5101 (
		_w15610_,
		_w15611_,
		_w15612_,
		_w15613_,
		_w15614_
	);
	LUT3 #(
		.INIT('h80)
	) name5102 (
		\wishbone_bd_ram_mem2_reg[72][18]/P0001 ,
		_w11949_,
		_w11990_,
		_w15615_
	);
	LUT3 #(
		.INIT('h80)
	) name5103 (
		\wishbone_bd_ram_mem2_reg[140][18]/P0001 ,
		_w11954_,
		_w11955_,
		_w15616_
	);
	LUT3 #(
		.INIT('h80)
	) name5104 (
		\wishbone_bd_ram_mem2_reg[67][18]/P0001 ,
		_w11938_,
		_w11949_,
		_w15617_
	);
	LUT3 #(
		.INIT('h80)
	) name5105 (
		\wishbone_bd_ram_mem2_reg[94][18]/P0001 ,
		_w11948_,
		_w11972_,
		_w15618_
	);
	LUT4 #(
		.INIT('h0001)
	) name5106 (
		_w15615_,
		_w15616_,
		_w15617_,
		_w15618_,
		_w15619_
	);
	LUT3 #(
		.INIT('h80)
	) name5107 (
		\wishbone_bd_ram_mem2_reg[205][18]/P0001 ,
		_w11945_,
		_w11966_,
		_w15620_
	);
	LUT3 #(
		.INIT('h80)
	) name5108 (
		\wishbone_bd_ram_mem2_reg[18][18]/P0001 ,
		_w11935_,
		_w11963_,
		_w15621_
	);
	LUT3 #(
		.INIT('h80)
	) name5109 (
		\wishbone_bd_ram_mem2_reg[188][18]/P0001 ,
		_w11942_,
		_w11954_,
		_w15622_
	);
	LUT3 #(
		.INIT('h80)
	) name5110 (
		\wishbone_bd_ram_mem2_reg[198][18]/P0001 ,
		_w11945_,
		_w11986_,
		_w15623_
	);
	LUT4 #(
		.INIT('h0001)
	) name5111 (
		_w15620_,
		_w15621_,
		_w15622_,
		_w15623_,
		_w15624_
	);
	LUT4 #(
		.INIT('h8000)
	) name5112 (
		_w15609_,
		_w15614_,
		_w15619_,
		_w15624_,
		_w15625_
	);
	LUT3 #(
		.INIT('h80)
	) name5113 (
		\wishbone_bd_ram_mem2_reg[240][18]/P0001 ,
		_w11941_,
		_w11952_,
		_w15626_
	);
	LUT3 #(
		.INIT('h80)
	) name5114 (
		\wishbone_bd_ram_mem2_reg[143][18]/P0001 ,
		_w11955_,
		_w11973_,
		_w15627_
	);
	LUT3 #(
		.INIT('h80)
	) name5115 (
		\wishbone_bd_ram_mem2_reg[24][18]/P0001 ,
		_w11935_,
		_w11990_,
		_w15628_
	);
	LUT3 #(
		.INIT('h80)
	) name5116 (
		\wishbone_bd_ram_mem2_reg[104][18]/P0001 ,
		_w11965_,
		_w11990_,
		_w15629_
	);
	LUT4 #(
		.INIT('h0001)
	) name5117 (
		_w15626_,
		_w15627_,
		_w15628_,
		_w15629_,
		_w15630_
	);
	LUT3 #(
		.INIT('h80)
	) name5118 (
		\wishbone_bd_ram_mem2_reg[165][18]/P0001 ,
		_w11930_,
		_w11933_,
		_w15631_
	);
	LUT3 #(
		.INIT('h80)
	) name5119 (
		\wishbone_bd_ram_mem2_reg[105][18]/P0001 ,
		_w11965_,
		_w11968_,
		_w15632_
	);
	LUT3 #(
		.INIT('h80)
	) name5120 (
		\wishbone_bd_ram_mem2_reg[46][18]/P0001 ,
		_w11948_,
		_w11957_,
		_w15633_
	);
	LUT3 #(
		.INIT('h80)
	) name5121 (
		\wishbone_bd_ram_mem2_reg[93][18]/P0001 ,
		_w11966_,
		_w11972_,
		_w15634_
	);
	LUT4 #(
		.INIT('h0001)
	) name5122 (
		_w15631_,
		_w15632_,
		_w15633_,
		_w15634_,
		_w15635_
	);
	LUT3 #(
		.INIT('h80)
	) name5123 (
		\wishbone_bd_ram_mem2_reg[209][18]/P0001 ,
		_w11977_,
		_w11984_,
		_w15636_
	);
	LUT3 #(
		.INIT('h80)
	) name5124 (
		\wishbone_bd_ram_mem2_reg[21][18]/P0001 ,
		_w11933_,
		_w11935_,
		_w15637_
	);
	LUT3 #(
		.INIT('h80)
	) name5125 (
		\wishbone_bd_ram_mem2_reg[233][18]/P0001 ,
		_w11968_,
		_w11982_,
		_w15638_
	);
	LUT3 #(
		.INIT('h80)
	) name5126 (
		\wishbone_bd_ram_mem2_reg[186][18]/P0001 ,
		_w11942_,
		_w11944_,
		_w15639_
	);
	LUT4 #(
		.INIT('h0001)
	) name5127 (
		_w15636_,
		_w15637_,
		_w15638_,
		_w15639_,
		_w15640_
	);
	LUT3 #(
		.INIT('h80)
	) name5128 (
		\wishbone_bd_ram_mem2_reg[194][18]/P0001 ,
		_w11945_,
		_w11963_,
		_w15641_
	);
	LUT3 #(
		.INIT('h80)
	) name5129 (
		\wishbone_bd_ram_mem2_reg[71][18]/P0001 ,
		_w11949_,
		_w11975_,
		_w15642_
	);
	LUT3 #(
		.INIT('h80)
	) name5130 (
		\wishbone_bd_ram_mem2_reg[31][18]/P0001 ,
		_w11935_,
		_w11973_,
		_w15643_
	);
	LUT3 #(
		.INIT('h80)
	) name5131 (
		\wishbone_bd_ram_mem2_reg[53][18]/P0001 ,
		_w11933_,
		_w11979_,
		_w15644_
	);
	LUT4 #(
		.INIT('h0001)
	) name5132 (
		_w15641_,
		_w15642_,
		_w15643_,
		_w15644_,
		_w15645_
	);
	LUT4 #(
		.INIT('h8000)
	) name5133 (
		_w15630_,
		_w15635_,
		_w15640_,
		_w15645_,
		_w15646_
	);
	LUT3 #(
		.INIT('h80)
	) name5134 (
		\wishbone_bd_ram_mem2_reg[19][18]/P0001 ,
		_w11935_,
		_w11938_,
		_w15647_
	);
	LUT3 #(
		.INIT('h80)
	) name5135 (
		\wishbone_bd_ram_mem2_reg[239][18]/P0001 ,
		_w11973_,
		_w11982_,
		_w15648_
	);
	LUT3 #(
		.INIT('h80)
	) name5136 (
		\wishbone_bd_ram_mem2_reg[78][18]/P0001 ,
		_w11948_,
		_w11949_,
		_w15649_
	);
	LUT3 #(
		.INIT('h80)
	) name5137 (
		\wishbone_bd_ram_mem2_reg[52][18]/P0001 ,
		_w11929_,
		_w11979_,
		_w15650_
	);
	LUT4 #(
		.INIT('h0001)
	) name5138 (
		_w15647_,
		_w15648_,
		_w15649_,
		_w15650_,
		_w15651_
	);
	LUT3 #(
		.INIT('h80)
	) name5139 (
		\wishbone_bd_ram_mem2_reg[74][18]/P0001 ,
		_w11944_,
		_w11949_,
		_w15652_
	);
	LUT3 #(
		.INIT('h80)
	) name5140 (
		\wishbone_bd_ram_mem2_reg[199][18]/P0001 ,
		_w11945_,
		_w11975_,
		_w15653_
	);
	LUT3 #(
		.INIT('h80)
	) name5141 (
		\wishbone_bd_ram_mem2_reg[217][18]/P0001 ,
		_w11968_,
		_w11984_,
		_w15654_
	);
	LUT3 #(
		.INIT('h80)
	) name5142 (
		\wishbone_bd_ram_mem2_reg[214][18]/P0001 ,
		_w11984_,
		_w11986_,
		_w15655_
	);
	LUT4 #(
		.INIT('h0001)
	) name5143 (
		_w15652_,
		_w15653_,
		_w15654_,
		_w15655_,
		_w15656_
	);
	LUT3 #(
		.INIT('h80)
	) name5144 (
		\wishbone_bd_ram_mem2_reg[235][18]/P0001 ,
		_w11936_,
		_w11982_,
		_w15657_
	);
	LUT3 #(
		.INIT('h80)
	) name5145 (
		\wishbone_bd_ram_mem2_reg[110][18]/P0001 ,
		_w11948_,
		_w11965_,
		_w15658_
	);
	LUT3 #(
		.INIT('h80)
	) name5146 (
		\wishbone_bd_ram_mem2_reg[27][18]/P0001 ,
		_w11935_,
		_w11936_,
		_w15659_
	);
	LUT3 #(
		.INIT('h80)
	) name5147 (
		\wishbone_bd_ram_mem2_reg[183][18]/P0001 ,
		_w11942_,
		_w11975_,
		_w15660_
	);
	LUT4 #(
		.INIT('h0001)
	) name5148 (
		_w15657_,
		_w15658_,
		_w15659_,
		_w15660_,
		_w15661_
	);
	LUT3 #(
		.INIT('h80)
	) name5149 (
		\wishbone_bd_ram_mem2_reg[192][18]/P0001 ,
		_w11941_,
		_w11945_,
		_w15662_
	);
	LUT3 #(
		.INIT('h80)
	) name5150 (
		\wishbone_bd_ram_mem2_reg[116][18]/P0001 ,
		_w11929_,
		_w12012_,
		_w15663_
	);
	LUT3 #(
		.INIT('h80)
	) name5151 (
		\wishbone_bd_ram_mem2_reg[36][18]/P0001 ,
		_w11929_,
		_w11957_,
		_w15664_
	);
	LUT3 #(
		.INIT('h80)
	) name5152 (
		\wishbone_bd_ram_mem2_reg[219][18]/P0001 ,
		_w11936_,
		_w11984_,
		_w15665_
	);
	LUT4 #(
		.INIT('h0001)
	) name5153 (
		_w15662_,
		_w15663_,
		_w15664_,
		_w15665_,
		_w15666_
	);
	LUT4 #(
		.INIT('h8000)
	) name5154 (
		_w15651_,
		_w15656_,
		_w15661_,
		_w15666_,
		_w15667_
	);
	LUT3 #(
		.INIT('h80)
	) name5155 (
		\wishbone_bd_ram_mem2_reg[145][18]/P0001 ,
		_w11959_,
		_w11977_,
		_w15668_
	);
	LUT3 #(
		.INIT('h80)
	) name5156 (
		\wishbone_bd_ram_mem2_reg[8][18]/P0001 ,
		_w11932_,
		_w11990_,
		_w15669_
	);
	LUT3 #(
		.INIT('h80)
	) name5157 (
		\wishbone_bd_ram_mem2_reg[133][18]/P0001 ,
		_w11933_,
		_w11955_,
		_w15670_
	);
	LUT3 #(
		.INIT('h80)
	) name5158 (
		\wishbone_bd_ram_mem2_reg[202][18]/P0001 ,
		_w11944_,
		_w11945_,
		_w15671_
	);
	LUT4 #(
		.INIT('h0001)
	) name5159 (
		_w15668_,
		_w15669_,
		_w15670_,
		_w15671_,
		_w15672_
	);
	LUT3 #(
		.INIT('h80)
	) name5160 (
		\wishbone_bd_ram_mem2_reg[62][18]/P0001 ,
		_w11948_,
		_w11979_,
		_w15673_
	);
	LUT3 #(
		.INIT('h80)
	) name5161 (
		\wishbone_bd_ram_mem2_reg[57][18]/P0001 ,
		_w11968_,
		_w11979_,
		_w15674_
	);
	LUT3 #(
		.INIT('h80)
	) name5162 (
		\wishbone_bd_ram_mem2_reg[117][18]/P0001 ,
		_w11933_,
		_w12012_,
		_w15675_
	);
	LUT3 #(
		.INIT('h80)
	) name5163 (
		\wishbone_bd_ram_mem2_reg[30][18]/P0001 ,
		_w11935_,
		_w11948_,
		_w15676_
	);
	LUT4 #(
		.INIT('h0001)
	) name5164 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15677_
	);
	LUT3 #(
		.INIT('h80)
	) name5165 (
		\wishbone_bd_ram_mem2_reg[137][18]/P0001 ,
		_w11955_,
		_w11968_,
		_w15678_
	);
	LUT3 #(
		.INIT('h80)
	) name5166 (
		\wishbone_bd_ram_mem2_reg[177][18]/P0001 ,
		_w11942_,
		_w11977_,
		_w15679_
	);
	LUT3 #(
		.INIT('h80)
	) name5167 (
		\wishbone_bd_ram_mem2_reg[154][18]/P0001 ,
		_w11944_,
		_w11959_,
		_w15680_
	);
	LUT3 #(
		.INIT('h80)
	) name5168 (
		\wishbone_bd_ram_mem2_reg[152][18]/P0001 ,
		_w11959_,
		_w11990_,
		_w15681_
	);
	LUT4 #(
		.INIT('h0001)
	) name5169 (
		_w15678_,
		_w15679_,
		_w15680_,
		_w15681_,
		_w15682_
	);
	LUT3 #(
		.INIT('h80)
	) name5170 (
		\wishbone_bd_ram_mem2_reg[158][18]/P0001 ,
		_w11948_,
		_w11959_,
		_w15683_
	);
	LUT3 #(
		.INIT('h80)
	) name5171 (
		\wishbone_bd_ram_mem2_reg[49][18]/P0001 ,
		_w11977_,
		_w11979_,
		_w15684_
	);
	LUT3 #(
		.INIT('h80)
	) name5172 (
		\wishbone_bd_ram_mem2_reg[204][18]/P0001 ,
		_w11945_,
		_w11954_,
		_w15685_
	);
	LUT3 #(
		.INIT('h80)
	) name5173 (
		\wishbone_bd_ram_mem2_reg[64][18]/P0001 ,
		_w11941_,
		_w11949_,
		_w15686_
	);
	LUT4 #(
		.INIT('h0001)
	) name5174 (
		_w15683_,
		_w15684_,
		_w15685_,
		_w15686_,
		_w15687_
	);
	LUT4 #(
		.INIT('h8000)
	) name5175 (
		_w15672_,
		_w15677_,
		_w15682_,
		_w15687_,
		_w15688_
	);
	LUT4 #(
		.INIT('h8000)
	) name5176 (
		_w15625_,
		_w15646_,
		_w15667_,
		_w15688_,
		_w15689_
	);
	LUT3 #(
		.INIT('h80)
	) name5177 (
		\wishbone_bd_ram_mem2_reg[203][18]/P0001 ,
		_w11936_,
		_w11945_,
		_w15690_
	);
	LUT3 #(
		.INIT('h80)
	) name5178 (
		\wishbone_bd_ram_mem2_reg[129][18]/P0001 ,
		_w11955_,
		_w11977_,
		_w15691_
	);
	LUT3 #(
		.INIT('h80)
	) name5179 (
		\wishbone_bd_ram_mem2_reg[246][18]/P0001 ,
		_w11952_,
		_w11986_,
		_w15692_
	);
	LUT3 #(
		.INIT('h80)
	) name5180 (
		\wishbone_bd_ram_mem2_reg[245][18]/P0001 ,
		_w11933_,
		_w11952_,
		_w15693_
	);
	LUT4 #(
		.INIT('h0001)
	) name5181 (
		_w15690_,
		_w15691_,
		_w15692_,
		_w15693_,
		_w15694_
	);
	LUT3 #(
		.INIT('h80)
	) name5182 (
		\wishbone_bd_ram_mem2_reg[144][18]/P0001 ,
		_w11941_,
		_w11959_,
		_w15695_
	);
	LUT3 #(
		.INIT('h80)
	) name5183 (
		\wishbone_bd_ram_mem2_reg[248][18]/P0001 ,
		_w11952_,
		_w11990_,
		_w15696_
	);
	LUT3 #(
		.INIT('h80)
	) name5184 (
		\wishbone_bd_ram_mem2_reg[135][18]/P0001 ,
		_w11955_,
		_w11975_,
		_w15697_
	);
	LUT3 #(
		.INIT('h80)
	) name5185 (
		\wishbone_bd_ram_mem2_reg[150][18]/P0001 ,
		_w11959_,
		_w11986_,
		_w15698_
	);
	LUT4 #(
		.INIT('h0001)
	) name5186 (
		_w15695_,
		_w15696_,
		_w15697_,
		_w15698_,
		_w15699_
	);
	LUT3 #(
		.INIT('h80)
	) name5187 (
		\wishbone_bd_ram_mem2_reg[215][18]/P0001 ,
		_w11975_,
		_w11984_,
		_w15700_
	);
	LUT3 #(
		.INIT('h80)
	) name5188 (
		\wishbone_bd_ram_mem2_reg[181][18]/P0001 ,
		_w11933_,
		_w11942_,
		_w15701_
	);
	LUT3 #(
		.INIT('h80)
	) name5189 (
		\wishbone_bd_ram_mem2_reg[190][18]/P0001 ,
		_w11942_,
		_w11948_,
		_w15702_
	);
	LUT3 #(
		.INIT('h80)
	) name5190 (
		\wishbone_bd_ram_mem2_reg[161][18]/P0001 ,
		_w11930_,
		_w11977_,
		_w15703_
	);
	LUT4 #(
		.INIT('h0001)
	) name5191 (
		_w15700_,
		_w15701_,
		_w15702_,
		_w15703_,
		_w15704_
	);
	LUT3 #(
		.INIT('h80)
	) name5192 (
		\wishbone_bd_ram_mem2_reg[35][18]/P0001 ,
		_w11938_,
		_w11957_,
		_w15705_
	);
	LUT3 #(
		.INIT('h80)
	) name5193 (
		\wishbone_bd_ram_mem2_reg[255][18]/P0001 ,
		_w11952_,
		_w11973_,
		_w15706_
	);
	LUT3 #(
		.INIT('h80)
	) name5194 (
		\wishbone_bd_ram_mem2_reg[54][18]/P0001 ,
		_w11979_,
		_w11986_,
		_w15707_
	);
	LUT3 #(
		.INIT('h80)
	) name5195 (
		\wishbone_bd_ram_mem2_reg[180][18]/P0001 ,
		_w11929_,
		_w11942_,
		_w15708_
	);
	LUT4 #(
		.INIT('h0001)
	) name5196 (
		_w15705_,
		_w15706_,
		_w15707_,
		_w15708_,
		_w15709_
	);
	LUT4 #(
		.INIT('h8000)
	) name5197 (
		_w15694_,
		_w15699_,
		_w15704_,
		_w15709_,
		_w15710_
	);
	LUT3 #(
		.INIT('h80)
	) name5198 (
		\wishbone_bd_ram_mem2_reg[220][18]/P0001 ,
		_w11954_,
		_w11984_,
		_w15711_
	);
	LUT3 #(
		.INIT('h80)
	) name5199 (
		\wishbone_bd_ram_mem2_reg[51][18]/P0001 ,
		_w11938_,
		_w11979_,
		_w15712_
	);
	LUT3 #(
		.INIT('h80)
	) name5200 (
		\wishbone_bd_ram_mem2_reg[60][18]/P0001 ,
		_w11954_,
		_w11979_,
		_w15713_
	);
	LUT3 #(
		.INIT('h80)
	) name5201 (
		\wishbone_bd_ram_mem2_reg[148][18]/P0001 ,
		_w11929_,
		_w11959_,
		_w15714_
	);
	LUT4 #(
		.INIT('h0001)
	) name5202 (
		_w15711_,
		_w15712_,
		_w15713_,
		_w15714_,
		_w15715_
	);
	LUT3 #(
		.INIT('h80)
	) name5203 (
		\wishbone_bd_ram_mem2_reg[231][18]/P0001 ,
		_w11975_,
		_w11982_,
		_w15716_
	);
	LUT3 #(
		.INIT('h80)
	) name5204 (
		\wishbone_bd_ram_mem2_reg[136][18]/P0001 ,
		_w11955_,
		_w11990_,
		_w15717_
	);
	LUT3 #(
		.INIT('h80)
	) name5205 (
		\wishbone_bd_ram_mem2_reg[225][18]/P0001 ,
		_w11977_,
		_w11982_,
		_w15718_
	);
	LUT3 #(
		.INIT('h80)
	) name5206 (
		\wishbone_bd_ram_mem2_reg[81][18]/P0001 ,
		_w11972_,
		_w11977_,
		_w15719_
	);
	LUT4 #(
		.INIT('h0001)
	) name5207 (
		_w15716_,
		_w15717_,
		_w15718_,
		_w15719_,
		_w15720_
	);
	LUT3 #(
		.INIT('h80)
	) name5208 (
		\wishbone_bd_ram_mem2_reg[26][18]/P0001 ,
		_w11935_,
		_w11944_,
		_w15721_
	);
	LUT3 #(
		.INIT('h80)
	) name5209 (
		\wishbone_bd_ram_mem2_reg[22][18]/P0001 ,
		_w11935_,
		_w11986_,
		_w15722_
	);
	LUT3 #(
		.INIT('h80)
	) name5210 (
		\wishbone_bd_ram_mem2_reg[92][18]/P0001 ,
		_w11954_,
		_w11972_,
		_w15723_
	);
	LUT3 #(
		.INIT('h80)
	) name5211 (
		\wishbone_bd_ram_mem2_reg[175][18]/P0001 ,
		_w11930_,
		_w11973_,
		_w15724_
	);
	LUT4 #(
		.INIT('h0001)
	) name5212 (
		_w15721_,
		_w15722_,
		_w15723_,
		_w15724_,
		_w15725_
	);
	LUT3 #(
		.INIT('h80)
	) name5213 (
		\wishbone_bd_ram_mem2_reg[243][18]/P0001 ,
		_w11938_,
		_w11952_,
		_w15726_
	);
	LUT3 #(
		.INIT('h80)
	) name5214 (
		\wishbone_bd_ram_mem2_reg[236][18]/P0001 ,
		_w11954_,
		_w11982_,
		_w15727_
	);
	LUT3 #(
		.INIT('h80)
	) name5215 (
		\wishbone_bd_ram_mem2_reg[73][18]/P0001 ,
		_w11949_,
		_w11968_,
		_w15728_
	);
	LUT3 #(
		.INIT('h80)
	) name5216 (
		\wishbone_bd_ram_mem2_reg[124][18]/P0001 ,
		_w11954_,
		_w12012_,
		_w15729_
	);
	LUT4 #(
		.INIT('h0001)
	) name5217 (
		_w15726_,
		_w15727_,
		_w15728_,
		_w15729_,
		_w15730_
	);
	LUT4 #(
		.INIT('h8000)
	) name5218 (
		_w15715_,
		_w15720_,
		_w15725_,
		_w15730_,
		_w15731_
	);
	LUT3 #(
		.INIT('h80)
	) name5219 (
		\wishbone_bd_ram_mem2_reg[141][18]/P0001 ,
		_w11955_,
		_w11966_,
		_w15732_
	);
	LUT3 #(
		.INIT('h80)
	) name5220 (
		\wishbone_bd_ram_mem2_reg[171][18]/P0001 ,
		_w11930_,
		_w11936_,
		_w15733_
	);
	LUT3 #(
		.INIT('h80)
	) name5221 (
		\wishbone_bd_ram_mem2_reg[164][18]/P0001 ,
		_w11929_,
		_w11930_,
		_w15734_
	);
	LUT3 #(
		.INIT('h80)
	) name5222 (
		\wishbone_bd_ram_mem2_reg[237][18]/P0001 ,
		_w11966_,
		_w11982_,
		_w15735_
	);
	LUT4 #(
		.INIT('h0001)
	) name5223 (
		_w15732_,
		_w15733_,
		_w15734_,
		_w15735_,
		_w15736_
	);
	LUT3 #(
		.INIT('h80)
	) name5224 (
		\wishbone_bd_ram_mem2_reg[118][18]/P0001 ,
		_w11986_,
		_w12012_,
		_w15737_
	);
	LUT3 #(
		.INIT('h80)
	) name5225 (
		\wishbone_bd_ram_mem2_reg[227][18]/P0001 ,
		_w11938_,
		_w11982_,
		_w15738_
	);
	LUT3 #(
		.INIT('h80)
	) name5226 (
		\wishbone_bd_ram_mem2_reg[112][18]/P0001 ,
		_w11941_,
		_w12012_,
		_w15739_
	);
	LUT3 #(
		.INIT('h80)
	) name5227 (
		\wishbone_bd_ram_mem2_reg[189][18]/P0001 ,
		_w11942_,
		_w11966_,
		_w15740_
	);
	LUT4 #(
		.INIT('h0001)
	) name5228 (
		_w15737_,
		_w15738_,
		_w15739_,
		_w15740_,
		_w15741_
	);
	LUT3 #(
		.INIT('h80)
	) name5229 (
		\wishbone_bd_ram_mem2_reg[223][18]/P0001 ,
		_w11973_,
		_w11984_,
		_w15742_
	);
	LUT3 #(
		.INIT('h80)
	) name5230 (
		\wishbone_bd_ram_mem2_reg[249][18]/P0001 ,
		_w11952_,
		_w11968_,
		_w15743_
	);
	LUT3 #(
		.INIT('h80)
	) name5231 (
		\wishbone_bd_ram_mem2_reg[173][18]/P0001 ,
		_w11930_,
		_w11966_,
		_w15744_
	);
	LUT3 #(
		.INIT('h80)
	) name5232 (
		\wishbone_bd_ram_mem2_reg[66][18]/P0001 ,
		_w11949_,
		_w11963_,
		_w15745_
	);
	LUT4 #(
		.INIT('h0001)
	) name5233 (
		_w15742_,
		_w15743_,
		_w15744_,
		_w15745_,
		_w15746_
	);
	LUT3 #(
		.INIT('h80)
	) name5234 (
		\wishbone_bd_ram_mem2_reg[142][18]/P0001 ,
		_w11948_,
		_w11955_,
		_w15747_
	);
	LUT3 #(
		.INIT('h80)
	) name5235 (
		\wishbone_bd_ram_mem2_reg[77][18]/P0001 ,
		_w11949_,
		_w11966_,
		_w15748_
	);
	LUT3 #(
		.INIT('h80)
	) name5236 (
		\wishbone_bd_ram_mem2_reg[83][18]/P0001 ,
		_w11938_,
		_w11972_,
		_w15749_
	);
	LUT3 #(
		.INIT('h80)
	) name5237 (
		\wishbone_bd_ram_mem2_reg[56][18]/P0001 ,
		_w11979_,
		_w11990_,
		_w15750_
	);
	LUT4 #(
		.INIT('h0001)
	) name5238 (
		_w15747_,
		_w15748_,
		_w15749_,
		_w15750_,
		_w15751_
	);
	LUT4 #(
		.INIT('h8000)
	) name5239 (
		_w15736_,
		_w15741_,
		_w15746_,
		_w15751_,
		_w15752_
	);
	LUT3 #(
		.INIT('h80)
	) name5240 (
		\wishbone_bd_ram_mem2_reg[98][18]/P0001 ,
		_w11963_,
		_w11965_,
		_w15753_
	);
	LUT3 #(
		.INIT('h80)
	) name5241 (
		\wishbone_bd_ram_mem2_reg[228][18]/P0001 ,
		_w11929_,
		_w11982_,
		_w15754_
	);
	LUT3 #(
		.INIT('h80)
	) name5242 (
		\wishbone_bd_ram_mem2_reg[69][18]/P0001 ,
		_w11933_,
		_w11949_,
		_w15755_
	);
	LUT3 #(
		.INIT('h80)
	) name5243 (
		\wishbone_bd_ram_mem2_reg[44][18]/P0001 ,
		_w11954_,
		_w11957_,
		_w15756_
	);
	LUT4 #(
		.INIT('h0001)
	) name5244 (
		_w15753_,
		_w15754_,
		_w15755_,
		_w15756_,
		_w15757_
	);
	LUT3 #(
		.INIT('h80)
	) name5245 (
		\wishbone_bd_ram_mem2_reg[213][18]/P0001 ,
		_w11933_,
		_w11984_,
		_w15758_
	);
	LUT3 #(
		.INIT('h80)
	) name5246 (
		\wishbone_bd_ram_mem2_reg[212][18]/P0001 ,
		_w11929_,
		_w11984_,
		_w15759_
	);
	LUT3 #(
		.INIT('h80)
	) name5247 (
		\wishbone_bd_ram_mem2_reg[63][18]/P0001 ,
		_w11973_,
		_w11979_,
		_w15760_
	);
	LUT3 #(
		.INIT('h80)
	) name5248 (
		\wishbone_bd_ram_mem2_reg[17][18]/P0001 ,
		_w11935_,
		_w11977_,
		_w15761_
	);
	LUT4 #(
		.INIT('h0001)
	) name5249 (
		_w15758_,
		_w15759_,
		_w15760_,
		_w15761_,
		_w15762_
	);
	LUT3 #(
		.INIT('h80)
	) name5250 (
		\wishbone_bd_ram_mem2_reg[253][18]/P0001 ,
		_w11952_,
		_w11966_,
		_w15763_
	);
	LUT3 #(
		.INIT('h80)
	) name5251 (
		\wishbone_bd_ram_mem2_reg[147][18]/P0001 ,
		_w11938_,
		_w11959_,
		_w15764_
	);
	LUT3 #(
		.INIT('h80)
	) name5252 (
		\wishbone_bd_ram_mem2_reg[28][18]/P0001 ,
		_w11935_,
		_w11954_,
		_w15765_
	);
	LUT3 #(
		.INIT('h80)
	) name5253 (
		\wishbone_bd_ram_mem2_reg[15][18]/P0001 ,
		_w11932_,
		_w11973_,
		_w15766_
	);
	LUT4 #(
		.INIT('h0001)
	) name5254 (
		_w15763_,
		_w15764_,
		_w15765_,
		_w15766_,
		_w15767_
	);
	LUT3 #(
		.INIT('h80)
	) name5255 (
		\wishbone_bd_ram_mem2_reg[168][18]/P0001 ,
		_w11930_,
		_w11990_,
		_w15768_
	);
	LUT3 #(
		.INIT('h80)
	) name5256 (
		\wishbone_bd_ram_mem2_reg[109][18]/P0001 ,
		_w11965_,
		_w11966_,
		_w15769_
	);
	LUT3 #(
		.INIT('h80)
	) name5257 (
		\wishbone_bd_ram_mem2_reg[182][18]/P0001 ,
		_w11942_,
		_w11986_,
		_w15770_
	);
	LUT3 #(
		.INIT('h80)
	) name5258 (
		\wishbone_bd_ram_mem2_reg[58][18]/P0001 ,
		_w11944_,
		_w11979_,
		_w15771_
	);
	LUT4 #(
		.INIT('h0001)
	) name5259 (
		_w15768_,
		_w15769_,
		_w15770_,
		_w15771_,
		_w15772_
	);
	LUT4 #(
		.INIT('h8000)
	) name5260 (
		_w15757_,
		_w15762_,
		_w15767_,
		_w15772_,
		_w15773_
	);
	LUT4 #(
		.INIT('h8000)
	) name5261 (
		_w15710_,
		_w15731_,
		_w15752_,
		_w15773_,
		_w15774_
	);
	LUT4 #(
		.INIT('h8000)
	) name5262 (
		_w15519_,
		_w15604_,
		_w15689_,
		_w15774_,
		_w15775_
	);
	LUT3 #(
		.INIT('h80)
	) name5263 (
		_w12304_,
		_w12314_,
		_w12316_,
		_w15776_
	);
	LUT3 #(
		.INIT('h15)
	) name5264 (
		_w12302_,
		_w12312_,
		_w15776_,
		_w15777_
	);
	LUT2 #(
		.INIT('h9)
	) name5265 (
		\wishbone_TxLength_reg[2]/NET0131 ,
		_w14878_,
		_w15778_
	);
	LUT2 #(
		.INIT('h8)
	) name5266 (
		_w15777_,
		_w15778_,
		_w15779_
	);
	LUT3 #(
		.INIT('hf2)
	) name5267 (
		_w12303_,
		_w15775_,
		_w15779_,
		_w15780_
	);
	LUT2 #(
		.INIT('hd)
	) name5268 (
		_w10582_,
		_w11368_,
		_w15781_
	);
	LUT3 #(
		.INIT('h80)
	) name5269 (
		\wishbone_bd_ram_mem2_reg[128][16]/P0001 ,
		_w11941_,
		_w11955_,
		_w15782_
	);
	LUT3 #(
		.INIT('h80)
	) name5270 (
		\wishbone_bd_ram_mem2_reg[55][16]/P0001 ,
		_w11975_,
		_w11979_,
		_w15783_
	);
	LUT3 #(
		.INIT('h80)
	) name5271 (
		\wishbone_bd_ram_mem2_reg[34][16]/P0001 ,
		_w11957_,
		_w11963_,
		_w15784_
	);
	LUT3 #(
		.INIT('h80)
	) name5272 (
		\wishbone_bd_ram_mem2_reg[125][16]/P0001 ,
		_w11966_,
		_w12012_,
		_w15785_
	);
	LUT4 #(
		.INIT('h0001)
	) name5273 (
		_w15782_,
		_w15783_,
		_w15784_,
		_w15785_,
		_w15786_
	);
	LUT3 #(
		.INIT('h80)
	) name5274 (
		\wishbone_bd_ram_mem2_reg[220][16]/P0001 ,
		_w11954_,
		_w11984_,
		_w15787_
	);
	LUT3 #(
		.INIT('h80)
	) name5275 (
		\wishbone_bd_ram_mem2_reg[118][16]/P0001 ,
		_w11986_,
		_w12012_,
		_w15788_
	);
	LUT3 #(
		.INIT('h80)
	) name5276 (
		\wishbone_bd_ram_mem2_reg[138][16]/P0001 ,
		_w11944_,
		_w11955_,
		_w15789_
	);
	LUT3 #(
		.INIT('h80)
	) name5277 (
		\wishbone_bd_ram_mem2_reg[127][16]/P0001 ,
		_w11973_,
		_w12012_,
		_w15790_
	);
	LUT4 #(
		.INIT('h0001)
	) name5278 (
		_w15787_,
		_w15788_,
		_w15789_,
		_w15790_,
		_w15791_
	);
	LUT3 #(
		.INIT('h80)
	) name5279 (
		\wishbone_bd_ram_mem2_reg[103][16]/P0001 ,
		_w11965_,
		_w11975_,
		_w15792_
	);
	LUT3 #(
		.INIT('h80)
	) name5280 (
		\wishbone_bd_ram_mem2_reg[69][16]/P0001 ,
		_w11933_,
		_w11949_,
		_w15793_
	);
	LUT3 #(
		.INIT('h80)
	) name5281 (
		\wishbone_bd_ram_mem2_reg[254][16]/P0001 ,
		_w11948_,
		_w11952_,
		_w15794_
	);
	LUT3 #(
		.INIT('h80)
	) name5282 (
		\wishbone_bd_ram_mem2_reg[39][16]/P0001 ,
		_w11957_,
		_w11975_,
		_w15795_
	);
	LUT4 #(
		.INIT('h0001)
	) name5283 (
		_w15792_,
		_w15793_,
		_w15794_,
		_w15795_,
		_w15796_
	);
	LUT3 #(
		.INIT('h80)
	) name5284 (
		\wishbone_bd_ram_mem2_reg[137][16]/P0001 ,
		_w11955_,
		_w11968_,
		_w15797_
	);
	LUT3 #(
		.INIT('h80)
	) name5285 (
		\wishbone_bd_ram_mem2_reg[20][16]/P0001 ,
		_w11929_,
		_w11935_,
		_w15798_
	);
	LUT3 #(
		.INIT('h80)
	) name5286 (
		\wishbone_bd_ram_mem2_reg[31][16]/P0001 ,
		_w11935_,
		_w11973_,
		_w15799_
	);
	LUT3 #(
		.INIT('h80)
	) name5287 (
		\wishbone_bd_ram_mem2_reg[237][16]/P0001 ,
		_w11966_,
		_w11982_,
		_w15800_
	);
	LUT4 #(
		.INIT('h0001)
	) name5288 (
		_w15797_,
		_w15798_,
		_w15799_,
		_w15800_,
		_w15801_
	);
	LUT4 #(
		.INIT('h8000)
	) name5289 (
		_w15786_,
		_w15791_,
		_w15796_,
		_w15801_,
		_w15802_
	);
	LUT3 #(
		.INIT('h80)
	) name5290 (
		\wishbone_bd_ram_mem2_reg[204][16]/P0001 ,
		_w11945_,
		_w11954_,
		_w15803_
	);
	LUT3 #(
		.INIT('h80)
	) name5291 (
		\wishbone_bd_ram_mem2_reg[120][16]/P0001 ,
		_w11990_,
		_w12012_,
		_w15804_
	);
	LUT3 #(
		.INIT('h80)
	) name5292 (
		\wishbone_bd_ram_mem2_reg[79][16]/P0001 ,
		_w11949_,
		_w11973_,
		_w15805_
	);
	LUT3 #(
		.INIT('h80)
	) name5293 (
		\wishbone_bd_ram_mem2_reg[6][16]/P0001 ,
		_w11932_,
		_w11986_,
		_w15806_
	);
	LUT4 #(
		.INIT('h0001)
	) name5294 (
		_w15803_,
		_w15804_,
		_w15805_,
		_w15806_,
		_w15807_
	);
	LUT3 #(
		.INIT('h80)
	) name5295 (
		\wishbone_bd_ram_mem2_reg[221][16]/P0001 ,
		_w11966_,
		_w11984_,
		_w15808_
	);
	LUT3 #(
		.INIT('h80)
	) name5296 (
		\wishbone_bd_ram_mem2_reg[0][16]/P0001 ,
		_w11932_,
		_w11941_,
		_w15809_
	);
	LUT3 #(
		.INIT('h80)
	) name5297 (
		\wishbone_bd_ram_mem2_reg[8][16]/P0001 ,
		_w11932_,
		_w11990_,
		_w15810_
	);
	LUT3 #(
		.INIT('h80)
	) name5298 (
		\wishbone_bd_ram_mem2_reg[100][16]/P0001 ,
		_w11929_,
		_w11965_,
		_w15811_
	);
	LUT4 #(
		.INIT('h0001)
	) name5299 (
		_w15808_,
		_w15809_,
		_w15810_,
		_w15811_,
		_w15812_
	);
	LUT3 #(
		.INIT('h80)
	) name5300 (
		\wishbone_bd_ram_mem2_reg[164][16]/P0001 ,
		_w11929_,
		_w11930_,
		_w15813_
	);
	LUT3 #(
		.INIT('h80)
	) name5301 (
		\wishbone_bd_ram_mem2_reg[188][16]/P0001 ,
		_w11942_,
		_w11954_,
		_w15814_
	);
	LUT3 #(
		.INIT('h80)
	) name5302 (
		\wishbone_bd_ram_mem2_reg[241][16]/P0001 ,
		_w11952_,
		_w11977_,
		_w15815_
	);
	LUT3 #(
		.INIT('h80)
	) name5303 (
		\wishbone_bd_ram_mem2_reg[197][16]/P0001 ,
		_w11933_,
		_w11945_,
		_w15816_
	);
	LUT4 #(
		.INIT('h0001)
	) name5304 (
		_w15813_,
		_w15814_,
		_w15815_,
		_w15816_,
		_w15817_
	);
	LUT3 #(
		.INIT('h80)
	) name5305 (
		\wishbone_bd_ram_mem2_reg[122][16]/P0001 ,
		_w11944_,
		_w12012_,
		_w15818_
	);
	LUT3 #(
		.INIT('h80)
	) name5306 (
		\wishbone_bd_ram_mem2_reg[33][16]/P0001 ,
		_w11957_,
		_w11977_,
		_w15819_
	);
	LUT3 #(
		.INIT('h80)
	) name5307 (
		\wishbone_bd_ram_mem2_reg[91][16]/P0001 ,
		_w11936_,
		_w11972_,
		_w15820_
	);
	LUT3 #(
		.INIT('h80)
	) name5308 (
		\wishbone_bd_ram_mem2_reg[161][16]/P0001 ,
		_w11930_,
		_w11977_,
		_w15821_
	);
	LUT4 #(
		.INIT('h0001)
	) name5309 (
		_w15818_,
		_w15819_,
		_w15820_,
		_w15821_,
		_w15822_
	);
	LUT4 #(
		.INIT('h8000)
	) name5310 (
		_w15807_,
		_w15812_,
		_w15817_,
		_w15822_,
		_w15823_
	);
	LUT3 #(
		.INIT('h80)
	) name5311 (
		\wishbone_bd_ram_mem2_reg[170][16]/P0001 ,
		_w11930_,
		_w11944_,
		_w15824_
	);
	LUT3 #(
		.INIT('h80)
	) name5312 (
		\wishbone_bd_ram_mem2_reg[71][16]/P0001 ,
		_w11949_,
		_w11975_,
		_w15825_
	);
	LUT3 #(
		.INIT('h80)
	) name5313 (
		\wishbone_bd_ram_mem2_reg[52][16]/P0001 ,
		_w11929_,
		_w11979_,
		_w15826_
	);
	LUT3 #(
		.INIT('h80)
	) name5314 (
		\wishbone_bd_ram_mem2_reg[40][16]/P0001 ,
		_w11957_,
		_w11990_,
		_w15827_
	);
	LUT4 #(
		.INIT('h0001)
	) name5315 (
		_w15824_,
		_w15825_,
		_w15826_,
		_w15827_,
		_w15828_
	);
	LUT3 #(
		.INIT('h80)
	) name5316 (
		\wishbone_bd_ram_mem2_reg[244][16]/P0001 ,
		_w11929_,
		_w11952_,
		_w15829_
	);
	LUT3 #(
		.INIT('h80)
	) name5317 (
		\wishbone_bd_ram_mem2_reg[129][16]/P0001 ,
		_w11955_,
		_w11977_,
		_w15830_
	);
	LUT3 #(
		.INIT('h80)
	) name5318 (
		\wishbone_bd_ram_mem2_reg[242][16]/P0001 ,
		_w11952_,
		_w11963_,
		_w15831_
	);
	LUT3 #(
		.INIT('h80)
	) name5319 (
		\wishbone_bd_ram_mem2_reg[11][16]/P0001 ,
		_w11932_,
		_w11936_,
		_w15832_
	);
	LUT4 #(
		.INIT('h0001)
	) name5320 (
		_w15829_,
		_w15830_,
		_w15831_,
		_w15832_,
		_w15833_
	);
	LUT3 #(
		.INIT('h80)
	) name5321 (
		\wishbone_bd_ram_mem2_reg[41][16]/P0001 ,
		_w11957_,
		_w11968_,
		_w15834_
	);
	LUT3 #(
		.INIT('h80)
	) name5322 (
		\wishbone_bd_ram_mem2_reg[240][16]/P0001 ,
		_w11941_,
		_w11952_,
		_w15835_
	);
	LUT3 #(
		.INIT('h80)
	) name5323 (
		\wishbone_bd_ram_mem2_reg[143][16]/P0001 ,
		_w11955_,
		_w11973_,
		_w15836_
	);
	LUT3 #(
		.INIT('h80)
	) name5324 (
		\wishbone_bd_ram_mem2_reg[139][16]/P0001 ,
		_w11936_,
		_w11955_,
		_w15837_
	);
	LUT4 #(
		.INIT('h0001)
	) name5325 (
		_w15834_,
		_w15835_,
		_w15836_,
		_w15837_,
		_w15838_
	);
	LUT3 #(
		.INIT('h80)
	) name5326 (
		\wishbone_bd_ram_mem2_reg[19][16]/P0001 ,
		_w11935_,
		_w11938_,
		_w15839_
	);
	LUT3 #(
		.INIT('h80)
	) name5327 (
		\wishbone_bd_ram_mem2_reg[247][16]/P0001 ,
		_w11952_,
		_w11975_,
		_w15840_
	);
	LUT3 #(
		.INIT('h80)
	) name5328 (
		\wishbone_bd_ram_mem2_reg[192][16]/P0001 ,
		_w11941_,
		_w11945_,
		_w15841_
	);
	LUT3 #(
		.INIT('h80)
	) name5329 (
		\wishbone_bd_ram_mem2_reg[81][16]/P0001 ,
		_w11972_,
		_w11977_,
		_w15842_
	);
	LUT4 #(
		.INIT('h0001)
	) name5330 (
		_w15839_,
		_w15840_,
		_w15841_,
		_w15842_,
		_w15843_
	);
	LUT4 #(
		.INIT('h8000)
	) name5331 (
		_w15828_,
		_w15833_,
		_w15838_,
		_w15843_,
		_w15844_
	);
	LUT3 #(
		.INIT('h80)
	) name5332 (
		\wishbone_bd_ram_mem2_reg[121][16]/P0001 ,
		_w11968_,
		_w12012_,
		_w15845_
	);
	LUT3 #(
		.INIT('h80)
	) name5333 (
		\wishbone_bd_ram_mem2_reg[102][16]/P0001 ,
		_w11965_,
		_w11986_,
		_w15846_
	);
	LUT3 #(
		.INIT('h80)
	) name5334 (
		\wishbone_bd_ram_mem2_reg[93][16]/P0001 ,
		_w11966_,
		_w11972_,
		_w15847_
	);
	LUT3 #(
		.INIT('h80)
	) name5335 (
		\wishbone_bd_ram_mem2_reg[158][16]/P0001 ,
		_w11948_,
		_w11959_,
		_w15848_
	);
	LUT4 #(
		.INIT('h0001)
	) name5336 (
		_w15845_,
		_w15846_,
		_w15847_,
		_w15848_,
		_w15849_
	);
	LUT3 #(
		.INIT('h80)
	) name5337 (
		\wishbone_bd_ram_mem2_reg[202][16]/P0001 ,
		_w11944_,
		_w11945_,
		_w15850_
	);
	LUT3 #(
		.INIT('h80)
	) name5338 (
		\wishbone_bd_ram_mem2_reg[99][16]/P0001 ,
		_w11938_,
		_w11965_,
		_w15851_
	);
	LUT3 #(
		.INIT('h80)
	) name5339 (
		\wishbone_bd_ram_mem2_reg[13][16]/P0001 ,
		_w11932_,
		_w11966_,
		_w15852_
	);
	LUT3 #(
		.INIT('h80)
	) name5340 (
		\wishbone_bd_ram_mem2_reg[193][16]/P0001 ,
		_w11945_,
		_w11977_,
		_w15853_
	);
	LUT4 #(
		.INIT('h0001)
	) name5341 (
		_w15850_,
		_w15851_,
		_w15852_,
		_w15853_,
		_w15854_
	);
	LUT3 #(
		.INIT('h80)
	) name5342 (
		\wishbone_bd_ram_mem2_reg[229][16]/P0001 ,
		_w11933_,
		_w11982_,
		_w15855_
	);
	LUT3 #(
		.INIT('h80)
	) name5343 (
		\wishbone_bd_ram_mem2_reg[206][16]/P0001 ,
		_w11945_,
		_w11948_,
		_w15856_
	);
	LUT3 #(
		.INIT('h80)
	) name5344 (
		\wishbone_bd_ram_mem2_reg[239][16]/P0001 ,
		_w11973_,
		_w11982_,
		_w15857_
	);
	LUT3 #(
		.INIT('h80)
	) name5345 (
		\wishbone_bd_ram_mem2_reg[48][16]/P0001 ,
		_w11941_,
		_w11979_,
		_w15858_
	);
	LUT4 #(
		.INIT('h0001)
	) name5346 (
		_w15855_,
		_w15856_,
		_w15857_,
		_w15858_,
		_w15859_
	);
	LUT3 #(
		.INIT('h80)
	) name5347 (
		\wishbone_bd_ram_mem2_reg[28][16]/P0001 ,
		_w11935_,
		_w11954_,
		_w15860_
	);
	LUT3 #(
		.INIT('h80)
	) name5348 (
		\wishbone_bd_ram_mem2_reg[105][16]/P0001 ,
		_w11965_,
		_w11968_,
		_w15861_
	);
	LUT3 #(
		.INIT('h80)
	) name5349 (
		\wishbone_bd_ram_mem2_reg[252][16]/P0001 ,
		_w11952_,
		_w11954_,
		_w15862_
	);
	LUT3 #(
		.INIT('h80)
	) name5350 (
		\wishbone_bd_ram_mem2_reg[149][16]/P0001 ,
		_w11933_,
		_w11959_,
		_w15863_
	);
	LUT4 #(
		.INIT('h0001)
	) name5351 (
		_w15860_,
		_w15861_,
		_w15862_,
		_w15863_,
		_w15864_
	);
	LUT4 #(
		.INIT('h8000)
	) name5352 (
		_w15849_,
		_w15854_,
		_w15859_,
		_w15864_,
		_w15865_
	);
	LUT4 #(
		.INIT('h8000)
	) name5353 (
		_w15802_,
		_w15823_,
		_w15844_,
		_w15865_,
		_w15866_
	);
	LUT3 #(
		.INIT('h80)
	) name5354 (
		\wishbone_bd_ram_mem2_reg[182][16]/P0001 ,
		_w11942_,
		_w11986_,
		_w15867_
	);
	LUT3 #(
		.INIT('h80)
	) name5355 (
		\wishbone_bd_ram_mem2_reg[42][16]/P0001 ,
		_w11944_,
		_w11957_,
		_w15868_
	);
	LUT3 #(
		.INIT('h80)
	) name5356 (
		\wishbone_bd_ram_mem2_reg[23][16]/P0001 ,
		_w11935_,
		_w11975_,
		_w15869_
	);
	LUT3 #(
		.INIT('h80)
	) name5357 (
		\wishbone_bd_ram_mem2_reg[213][16]/P0001 ,
		_w11933_,
		_w11984_,
		_w15870_
	);
	LUT4 #(
		.INIT('h0001)
	) name5358 (
		_w15867_,
		_w15868_,
		_w15869_,
		_w15870_,
		_w15871_
	);
	LUT3 #(
		.INIT('h80)
	) name5359 (
		\wishbone_bd_ram_mem2_reg[74][16]/P0001 ,
		_w11944_,
		_w11949_,
		_w15872_
	);
	LUT3 #(
		.INIT('h80)
	) name5360 (
		\wishbone_bd_ram_mem2_reg[116][16]/P0001 ,
		_w11929_,
		_w12012_,
		_w15873_
	);
	LUT3 #(
		.INIT('h80)
	) name5361 (
		\wishbone_bd_ram_mem2_reg[101][16]/P0001 ,
		_w11933_,
		_w11965_,
		_w15874_
	);
	LUT3 #(
		.INIT('h80)
	) name5362 (
		\wishbone_bd_ram_mem2_reg[58][16]/P0001 ,
		_w11944_,
		_w11979_,
		_w15875_
	);
	LUT4 #(
		.INIT('h0001)
	) name5363 (
		_w15872_,
		_w15873_,
		_w15874_,
		_w15875_,
		_w15876_
	);
	LUT3 #(
		.INIT('h80)
	) name5364 (
		\wishbone_bd_ram_mem2_reg[196][16]/P0001 ,
		_w11929_,
		_w11945_,
		_w15877_
	);
	LUT3 #(
		.INIT('h80)
	) name5365 (
		\wishbone_bd_ram_mem2_reg[1][16]/P0001 ,
		_w11932_,
		_w11977_,
		_w15878_
	);
	LUT3 #(
		.INIT('h80)
	) name5366 (
		\wishbone_bd_ram_mem2_reg[17][16]/P0001 ,
		_w11935_,
		_w11977_,
		_w15879_
	);
	LUT3 #(
		.INIT('h80)
	) name5367 (
		\wishbone_bd_ram_mem2_reg[2][16]/P0001 ,
		_w11932_,
		_w11963_,
		_w15880_
	);
	LUT4 #(
		.INIT('h0001)
	) name5368 (
		_w15877_,
		_w15878_,
		_w15879_,
		_w15880_,
		_w15881_
	);
	LUT3 #(
		.INIT('h80)
	) name5369 (
		\wishbone_bd_ram_mem2_reg[218][16]/P0001 ,
		_w11944_,
		_w11984_,
		_w15882_
	);
	LUT3 #(
		.INIT('h80)
	) name5370 (
		\wishbone_bd_ram_mem2_reg[10][16]/P0001 ,
		_w11932_,
		_w11944_,
		_w15883_
	);
	LUT3 #(
		.INIT('h80)
	) name5371 (
		\wishbone_bd_ram_mem2_reg[75][16]/P0001 ,
		_w11936_,
		_w11949_,
		_w15884_
	);
	LUT3 #(
		.INIT('h80)
	) name5372 (
		\wishbone_bd_ram_mem2_reg[184][16]/P0001 ,
		_w11942_,
		_w11990_,
		_w15885_
	);
	LUT4 #(
		.INIT('h0001)
	) name5373 (
		_w15882_,
		_w15883_,
		_w15884_,
		_w15885_,
		_w15886_
	);
	LUT4 #(
		.INIT('h8000)
	) name5374 (
		_w15871_,
		_w15876_,
		_w15881_,
		_w15886_,
		_w15887_
	);
	LUT3 #(
		.INIT('h80)
	) name5375 (
		\wishbone_bd_ram_mem2_reg[126][16]/P0001 ,
		_w11948_,
		_w12012_,
		_w15888_
	);
	LUT3 #(
		.INIT('h80)
	) name5376 (
		\wishbone_bd_ram_mem2_reg[235][16]/P0001 ,
		_w11936_,
		_w11982_,
		_w15889_
	);
	LUT3 #(
		.INIT('h80)
	) name5377 (
		\wishbone_bd_ram_mem2_reg[32][16]/P0001 ,
		_w11941_,
		_w11957_,
		_w15890_
	);
	LUT3 #(
		.INIT('h80)
	) name5378 (
		\wishbone_bd_ram_mem2_reg[185][16]/P0001 ,
		_w11942_,
		_w11968_,
		_w15891_
	);
	LUT4 #(
		.INIT('h0001)
	) name5379 (
		_w15888_,
		_w15889_,
		_w15890_,
		_w15891_,
		_w15892_
	);
	LUT3 #(
		.INIT('h80)
	) name5380 (
		\wishbone_bd_ram_mem2_reg[24][16]/P0001 ,
		_w11935_,
		_w11990_,
		_w15893_
	);
	LUT3 #(
		.INIT('h80)
	) name5381 (
		\wishbone_bd_ram_mem2_reg[108][16]/P0001 ,
		_w11954_,
		_w11965_,
		_w15894_
	);
	LUT3 #(
		.INIT('h80)
	) name5382 (
		\wishbone_bd_ram_mem2_reg[77][16]/P0001 ,
		_w11949_,
		_w11966_,
		_w15895_
	);
	LUT3 #(
		.INIT('h80)
	) name5383 (
		\wishbone_bd_ram_mem2_reg[147][16]/P0001 ,
		_w11938_,
		_w11959_,
		_w15896_
	);
	LUT4 #(
		.INIT('h0001)
	) name5384 (
		_w15893_,
		_w15894_,
		_w15895_,
		_w15896_,
		_w15897_
	);
	LUT3 #(
		.INIT('h80)
	) name5385 (
		\wishbone_bd_ram_mem2_reg[219][16]/P0001 ,
		_w11936_,
		_w11984_,
		_w15898_
	);
	LUT3 #(
		.INIT('h80)
	) name5386 (
		\wishbone_bd_ram_mem2_reg[47][16]/P0001 ,
		_w11957_,
		_w11973_,
		_w15899_
	);
	LUT3 #(
		.INIT('h80)
	) name5387 (
		\wishbone_bd_ram_mem2_reg[30][16]/P0001 ,
		_w11935_,
		_w11948_,
		_w15900_
	);
	LUT3 #(
		.INIT('h80)
	) name5388 (
		\wishbone_bd_ram_mem2_reg[7][16]/P0001 ,
		_w11932_,
		_w11975_,
		_w15901_
	);
	LUT4 #(
		.INIT('h0001)
	) name5389 (
		_w15898_,
		_w15899_,
		_w15900_,
		_w15901_,
		_w15902_
	);
	LUT3 #(
		.INIT('h80)
	) name5390 (
		\wishbone_bd_ram_mem2_reg[148][16]/P0001 ,
		_w11929_,
		_w11959_,
		_w15903_
	);
	LUT3 #(
		.INIT('h80)
	) name5391 (
		\wishbone_bd_ram_mem2_reg[117][16]/P0001 ,
		_w11933_,
		_w12012_,
		_w15904_
	);
	LUT3 #(
		.INIT('h80)
	) name5392 (
		\wishbone_bd_ram_mem2_reg[59][16]/P0001 ,
		_w11936_,
		_w11979_,
		_w15905_
	);
	LUT3 #(
		.INIT('h80)
	) name5393 (
		\wishbone_bd_ram_mem2_reg[160][16]/P0001 ,
		_w11930_,
		_w11941_,
		_w15906_
	);
	LUT4 #(
		.INIT('h0001)
	) name5394 (
		_w15903_,
		_w15904_,
		_w15905_,
		_w15906_,
		_w15907_
	);
	LUT4 #(
		.INIT('h8000)
	) name5395 (
		_w15892_,
		_w15897_,
		_w15902_,
		_w15907_,
		_w15908_
	);
	LUT3 #(
		.INIT('h80)
	) name5396 (
		\wishbone_bd_ram_mem2_reg[124][16]/P0001 ,
		_w11954_,
		_w12012_,
		_w15909_
	);
	LUT3 #(
		.INIT('h80)
	) name5397 (
		\wishbone_bd_ram_mem2_reg[57][16]/P0001 ,
		_w11968_,
		_w11979_,
		_w15910_
	);
	LUT3 #(
		.INIT('h80)
	) name5398 (
		\wishbone_bd_ram_mem2_reg[45][16]/P0001 ,
		_w11957_,
		_w11966_,
		_w15911_
	);
	LUT3 #(
		.INIT('h80)
	) name5399 (
		\wishbone_bd_ram_mem2_reg[190][16]/P0001 ,
		_w11942_,
		_w11948_,
		_w15912_
	);
	LUT4 #(
		.INIT('h0001)
	) name5400 (
		_w15909_,
		_w15910_,
		_w15911_,
		_w15912_,
		_w15913_
	);
	LUT3 #(
		.INIT('h80)
	) name5401 (
		\wishbone_bd_ram_mem2_reg[134][16]/P0001 ,
		_w11955_,
		_w11986_,
		_w15914_
	);
	LUT3 #(
		.INIT('h80)
	) name5402 (
		\wishbone_bd_ram_mem2_reg[234][16]/P0001 ,
		_w11944_,
		_w11982_,
		_w15915_
	);
	LUT3 #(
		.INIT('h80)
	) name5403 (
		\wishbone_bd_ram_mem2_reg[203][16]/P0001 ,
		_w11936_,
		_w11945_,
		_w15916_
	);
	LUT3 #(
		.INIT('h80)
	) name5404 (
		\wishbone_bd_ram_mem2_reg[49][16]/P0001 ,
		_w11977_,
		_w11979_,
		_w15917_
	);
	LUT4 #(
		.INIT('h0001)
	) name5405 (
		_w15914_,
		_w15915_,
		_w15916_,
		_w15917_,
		_w15918_
	);
	LUT3 #(
		.INIT('h80)
	) name5406 (
		\wishbone_bd_ram_mem2_reg[36][16]/P0001 ,
		_w11929_,
		_w11957_,
		_w15919_
	);
	LUT3 #(
		.INIT('h80)
	) name5407 (
		\wishbone_bd_ram_mem2_reg[150][16]/P0001 ,
		_w11959_,
		_w11986_,
		_w15920_
	);
	LUT3 #(
		.INIT('h80)
	) name5408 (
		\wishbone_bd_ram_mem2_reg[115][16]/P0001 ,
		_w11938_,
		_w12012_,
		_w15921_
	);
	LUT3 #(
		.INIT('h80)
	) name5409 (
		\wishbone_bd_ram_mem2_reg[163][16]/P0001 ,
		_w11930_,
		_w11938_,
		_w15922_
	);
	LUT4 #(
		.INIT('h0001)
	) name5410 (
		_w15919_,
		_w15920_,
		_w15921_,
		_w15922_,
		_w15923_
	);
	LUT3 #(
		.INIT('h80)
	) name5411 (
		\wishbone_bd_ram_mem2_reg[200][16]/P0001 ,
		_w11945_,
		_w11990_,
		_w15924_
	);
	LUT3 #(
		.INIT('h80)
	) name5412 (
		\wishbone_bd_ram_mem2_reg[44][16]/P0001 ,
		_w11954_,
		_w11957_,
		_w15925_
	);
	LUT3 #(
		.INIT('h80)
	) name5413 (
		\wishbone_bd_ram_mem2_reg[96][16]/P0001 ,
		_w11941_,
		_w11965_,
		_w15926_
	);
	LUT3 #(
		.INIT('h80)
	) name5414 (
		\wishbone_bd_ram_mem2_reg[38][16]/P0001 ,
		_w11957_,
		_w11986_,
		_w15927_
	);
	LUT4 #(
		.INIT('h0001)
	) name5415 (
		_w15924_,
		_w15925_,
		_w15926_,
		_w15927_,
		_w15928_
	);
	LUT4 #(
		.INIT('h8000)
	) name5416 (
		_w15913_,
		_w15918_,
		_w15923_,
		_w15928_,
		_w15929_
	);
	LUT3 #(
		.INIT('h80)
	) name5417 (
		\wishbone_bd_ram_mem2_reg[62][16]/P0001 ,
		_w11948_,
		_w11979_,
		_w15930_
	);
	LUT3 #(
		.INIT('h80)
	) name5418 (
		\wishbone_bd_ram_mem2_reg[21][16]/P0001 ,
		_w11933_,
		_w11935_,
		_w15931_
	);
	LUT3 #(
		.INIT('h80)
	) name5419 (
		\wishbone_bd_ram_mem2_reg[67][16]/P0001 ,
		_w11938_,
		_w11949_,
		_w15932_
	);
	LUT3 #(
		.INIT('h80)
	) name5420 (
		\wishbone_bd_ram_mem2_reg[159][16]/P0001 ,
		_w11959_,
		_w11973_,
		_w15933_
	);
	LUT4 #(
		.INIT('h0001)
	) name5421 (
		_w15930_,
		_w15931_,
		_w15932_,
		_w15933_,
		_w15934_
	);
	LUT3 #(
		.INIT('h80)
	) name5422 (
		\wishbone_bd_ram_mem2_reg[191][16]/P0001 ,
		_w11942_,
		_w11973_,
		_w15935_
	);
	LUT3 #(
		.INIT('h80)
	) name5423 (
		\wishbone_bd_ram_mem2_reg[80][16]/P0001 ,
		_w11941_,
		_w11972_,
		_w15936_
	);
	LUT3 #(
		.INIT('h80)
	) name5424 (
		\wishbone_bd_ram_mem2_reg[214][16]/P0001 ,
		_w11984_,
		_w11986_,
		_w15937_
	);
	LUT3 #(
		.INIT('h80)
	) name5425 (
		\wishbone_bd_ram_mem2_reg[194][16]/P0001 ,
		_w11945_,
		_w11963_,
		_w15938_
	);
	LUT4 #(
		.INIT('h0001)
	) name5426 (
		_w15935_,
		_w15936_,
		_w15937_,
		_w15938_,
		_w15939_
	);
	LUT3 #(
		.INIT('h80)
	) name5427 (
		\wishbone_bd_ram_mem2_reg[246][16]/P0001 ,
		_w11952_,
		_w11986_,
		_w15940_
	);
	LUT3 #(
		.INIT('h80)
	) name5428 (
		\wishbone_bd_ram_mem2_reg[151][16]/P0001 ,
		_w11959_,
		_w11975_,
		_w15941_
	);
	LUT3 #(
		.INIT('h80)
	) name5429 (
		\wishbone_bd_ram_mem2_reg[172][16]/P0001 ,
		_w11930_,
		_w11954_,
		_w15942_
	);
	LUT3 #(
		.INIT('h80)
	) name5430 (
		\wishbone_bd_ram_mem2_reg[86][16]/P0001 ,
		_w11972_,
		_w11986_,
		_w15943_
	);
	LUT4 #(
		.INIT('h0001)
	) name5431 (
		_w15940_,
		_w15941_,
		_w15942_,
		_w15943_,
		_w15944_
	);
	LUT3 #(
		.INIT('h80)
	) name5432 (
		\wishbone_bd_ram_mem2_reg[231][16]/P0001 ,
		_w11975_,
		_w11982_,
		_w15945_
	);
	LUT3 #(
		.INIT('h80)
	) name5433 (
		\wishbone_bd_ram_mem2_reg[183][16]/P0001 ,
		_w11942_,
		_w11975_,
		_w15946_
	);
	LUT3 #(
		.INIT('h80)
	) name5434 (
		\wishbone_bd_ram_mem2_reg[112][16]/P0001 ,
		_w11941_,
		_w12012_,
		_w15947_
	);
	LUT3 #(
		.INIT('h80)
	) name5435 (
		\wishbone_bd_ram_mem2_reg[88][16]/P0001 ,
		_w11972_,
		_w11990_,
		_w15948_
	);
	LUT4 #(
		.INIT('h0001)
	) name5436 (
		_w15945_,
		_w15946_,
		_w15947_,
		_w15948_,
		_w15949_
	);
	LUT4 #(
		.INIT('h8000)
	) name5437 (
		_w15934_,
		_w15939_,
		_w15944_,
		_w15949_,
		_w15950_
	);
	LUT4 #(
		.INIT('h8000)
	) name5438 (
		_w15887_,
		_w15908_,
		_w15929_,
		_w15950_,
		_w15951_
	);
	LUT3 #(
		.INIT('h80)
	) name5439 (
		\wishbone_bd_ram_mem2_reg[3][16]/P0001 ,
		_w11932_,
		_w11938_,
		_w15952_
	);
	LUT3 #(
		.INIT('h80)
	) name5440 (
		\wishbone_bd_ram_mem2_reg[98][16]/P0001 ,
		_w11963_,
		_w11965_,
		_w15953_
	);
	LUT3 #(
		.INIT('h80)
	) name5441 (
		\wishbone_bd_ram_mem2_reg[168][16]/P0001 ,
		_w11930_,
		_w11990_,
		_w15954_
	);
	LUT3 #(
		.INIT('h80)
	) name5442 (
		\wishbone_bd_ram_mem2_reg[64][16]/P0001 ,
		_w11941_,
		_w11949_,
		_w15955_
	);
	LUT4 #(
		.INIT('h0001)
	) name5443 (
		_w15952_,
		_w15953_,
		_w15954_,
		_w15955_,
		_w15956_
	);
	LUT3 #(
		.INIT('h80)
	) name5444 (
		\wishbone_bd_ram_mem2_reg[18][16]/P0001 ,
		_w11935_,
		_w11963_,
		_w15957_
	);
	LUT3 #(
		.INIT('h80)
	) name5445 (
		\wishbone_bd_ram_mem2_reg[136][16]/P0001 ,
		_w11955_,
		_w11990_,
		_w15958_
	);
	LUT3 #(
		.INIT('h80)
	) name5446 (
		\wishbone_bd_ram_mem2_reg[152][16]/P0001 ,
		_w11959_,
		_w11990_,
		_w15959_
	);
	LUT3 #(
		.INIT('h80)
	) name5447 (
		\wishbone_bd_ram_mem2_reg[146][16]/P0001 ,
		_w11959_,
		_w11963_,
		_w15960_
	);
	LUT4 #(
		.INIT('h0001)
	) name5448 (
		_w15957_,
		_w15958_,
		_w15959_,
		_w15960_,
		_w15961_
	);
	LUT3 #(
		.INIT('h80)
	) name5449 (
		\wishbone_bd_ram_mem2_reg[51][16]/P0001 ,
		_w11938_,
		_w11979_,
		_w15962_
	);
	LUT3 #(
		.INIT('h80)
	) name5450 (
		\wishbone_bd_ram_mem2_reg[223][16]/P0001 ,
		_w11973_,
		_w11984_,
		_w15963_
	);
	LUT3 #(
		.INIT('h80)
	) name5451 (
		\wishbone_bd_ram_mem2_reg[9][16]/P0001 ,
		_w11932_,
		_w11968_,
		_w15964_
	);
	LUT3 #(
		.INIT('h80)
	) name5452 (
		\wishbone_bd_ram_mem2_reg[70][16]/P0001 ,
		_w11949_,
		_w11986_,
		_w15965_
	);
	LUT4 #(
		.INIT('h0001)
	) name5453 (
		_w15962_,
		_w15963_,
		_w15964_,
		_w15965_,
		_w15966_
	);
	LUT3 #(
		.INIT('h80)
	) name5454 (
		\wishbone_bd_ram_mem2_reg[215][16]/P0001 ,
		_w11975_,
		_w11984_,
		_w15967_
	);
	LUT3 #(
		.INIT('h80)
	) name5455 (
		\wishbone_bd_ram_mem2_reg[176][16]/P0001 ,
		_w11941_,
		_w11942_,
		_w15968_
	);
	LUT3 #(
		.INIT('h80)
	) name5456 (
		\wishbone_bd_ram_mem2_reg[37][16]/P0001 ,
		_w11933_,
		_w11957_,
		_w15969_
	);
	LUT3 #(
		.INIT('h80)
	) name5457 (
		\wishbone_bd_ram_mem2_reg[54][16]/P0001 ,
		_w11979_,
		_w11986_,
		_w15970_
	);
	LUT4 #(
		.INIT('h0001)
	) name5458 (
		_w15967_,
		_w15968_,
		_w15969_,
		_w15970_,
		_w15971_
	);
	LUT4 #(
		.INIT('h8000)
	) name5459 (
		_w15956_,
		_w15961_,
		_w15966_,
		_w15971_,
		_w15972_
	);
	LUT3 #(
		.INIT('h80)
	) name5460 (
		\wishbone_bd_ram_mem2_reg[50][16]/P0001 ,
		_w11963_,
		_w11979_,
		_w15973_
	);
	LUT3 #(
		.INIT('h80)
	) name5461 (
		\wishbone_bd_ram_mem2_reg[162][16]/P0001 ,
		_w11930_,
		_w11963_,
		_w15974_
	);
	LUT3 #(
		.INIT('h80)
	) name5462 (
		\wishbone_bd_ram_mem2_reg[157][16]/P0001 ,
		_w11959_,
		_w11966_,
		_w15975_
	);
	LUT3 #(
		.INIT('h80)
	) name5463 (
		\wishbone_bd_ram_mem2_reg[253][16]/P0001 ,
		_w11952_,
		_w11966_,
		_w15976_
	);
	LUT4 #(
		.INIT('h0001)
	) name5464 (
		_w15973_,
		_w15974_,
		_w15975_,
		_w15976_,
		_w15977_
	);
	LUT3 #(
		.INIT('h80)
	) name5465 (
		\wishbone_bd_ram_mem2_reg[22][16]/P0001 ,
		_w11935_,
		_w11986_,
		_w15978_
	);
	LUT3 #(
		.INIT('h80)
	) name5466 (
		\wishbone_bd_ram_mem2_reg[236][16]/P0001 ,
		_w11954_,
		_w11982_,
		_w15979_
	);
	LUT3 #(
		.INIT('h80)
	) name5467 (
		\wishbone_bd_ram_mem2_reg[255][16]/P0001 ,
		_w11952_,
		_w11973_,
		_w15980_
	);
	LUT3 #(
		.INIT('h80)
	) name5468 (
		\wishbone_bd_ram_mem2_reg[211][16]/P0001 ,
		_w11938_,
		_w11984_,
		_w15981_
	);
	LUT4 #(
		.INIT('h0001)
	) name5469 (
		_w15978_,
		_w15979_,
		_w15980_,
		_w15981_,
		_w15982_
	);
	LUT3 #(
		.INIT('h80)
	) name5470 (
		\wishbone_bd_ram_mem2_reg[72][16]/P0001 ,
		_w11949_,
		_w11990_,
		_w15983_
	);
	LUT3 #(
		.INIT('h80)
	) name5471 (
		\wishbone_bd_ram_mem2_reg[174][16]/P0001 ,
		_w11930_,
		_w11948_,
		_w15984_
	);
	LUT3 #(
		.INIT('h80)
	) name5472 (
		\wishbone_bd_ram_mem2_reg[27][16]/P0001 ,
		_w11935_,
		_w11936_,
		_w15985_
	);
	LUT3 #(
		.INIT('h80)
	) name5473 (
		\wishbone_bd_ram_mem2_reg[154][16]/P0001 ,
		_w11944_,
		_w11959_,
		_w15986_
	);
	LUT4 #(
		.INIT('h0001)
	) name5474 (
		_w15983_,
		_w15984_,
		_w15985_,
		_w15986_,
		_w15987_
	);
	LUT3 #(
		.INIT('h80)
	) name5475 (
		\wishbone_bd_ram_mem2_reg[156][16]/P0001 ,
		_w11954_,
		_w11959_,
		_w15988_
	);
	LUT3 #(
		.INIT('h80)
	) name5476 (
		\wishbone_bd_ram_mem2_reg[166][16]/P0001 ,
		_w11930_,
		_w11986_,
		_w15989_
	);
	LUT3 #(
		.INIT('h80)
	) name5477 (
		\wishbone_bd_ram_mem2_reg[53][16]/P0001 ,
		_w11933_,
		_w11979_,
		_w15990_
	);
	LUT3 #(
		.INIT('h80)
	) name5478 (
		\wishbone_bd_ram_mem2_reg[123][16]/P0001 ,
		_w11936_,
		_w12012_,
		_w15991_
	);
	LUT4 #(
		.INIT('h0001)
	) name5479 (
		_w15988_,
		_w15989_,
		_w15990_,
		_w15991_,
		_w15992_
	);
	LUT4 #(
		.INIT('h8000)
	) name5480 (
		_w15977_,
		_w15982_,
		_w15987_,
		_w15992_,
		_w15993_
	);
	LUT3 #(
		.INIT('h80)
	) name5481 (
		\wishbone_bd_ram_mem2_reg[4][16]/P0001 ,
		_w11929_,
		_w11932_,
		_w15994_
	);
	LUT3 #(
		.INIT('h80)
	) name5482 (
		\wishbone_bd_ram_mem2_reg[224][16]/P0001 ,
		_w11941_,
		_w11982_,
		_w15995_
	);
	LUT3 #(
		.INIT('h80)
	) name5483 (
		\wishbone_bd_ram_mem2_reg[107][16]/P0001 ,
		_w11936_,
		_w11965_,
		_w15996_
	);
	LUT3 #(
		.INIT('h80)
	) name5484 (
		\wishbone_bd_ram_mem2_reg[145][16]/P0001 ,
		_w11959_,
		_w11977_,
		_w15997_
	);
	LUT4 #(
		.INIT('h0001)
	) name5485 (
		_w15994_,
		_w15995_,
		_w15996_,
		_w15997_,
		_w15998_
	);
	LUT3 #(
		.INIT('h80)
	) name5486 (
		\wishbone_bd_ram_mem2_reg[84][16]/P0001 ,
		_w11929_,
		_w11972_,
		_w15999_
	);
	LUT3 #(
		.INIT('h80)
	) name5487 (
		\wishbone_bd_ram_mem2_reg[83][16]/P0001 ,
		_w11938_,
		_w11972_,
		_w16000_
	);
	LUT3 #(
		.INIT('h80)
	) name5488 (
		\wishbone_bd_ram_mem2_reg[179][16]/P0001 ,
		_w11938_,
		_w11942_,
		_w16001_
	);
	LUT3 #(
		.INIT('h80)
	) name5489 (
		\wishbone_bd_ram_mem2_reg[130][16]/P0001 ,
		_w11955_,
		_w11963_,
		_w16002_
	);
	LUT4 #(
		.INIT('h0001)
	) name5490 (
		_w15999_,
		_w16000_,
		_w16001_,
		_w16002_,
		_w16003_
	);
	LUT3 #(
		.INIT('h80)
	) name5491 (
		\wishbone_bd_ram_mem2_reg[94][16]/P0001 ,
		_w11948_,
		_w11972_,
		_w16004_
	);
	LUT3 #(
		.INIT('h80)
	) name5492 (
		\wishbone_bd_ram_mem2_reg[217][16]/P0001 ,
		_w11968_,
		_w11984_,
		_w16005_
	);
	LUT3 #(
		.INIT('h80)
	) name5493 (
		\wishbone_bd_ram_mem2_reg[144][16]/P0001 ,
		_w11941_,
		_w11959_,
		_w16006_
	);
	LUT3 #(
		.INIT('h80)
	) name5494 (
		\wishbone_bd_ram_mem2_reg[73][16]/P0001 ,
		_w11949_,
		_w11968_,
		_w16007_
	);
	LUT4 #(
		.INIT('h0001)
	) name5495 (
		_w16004_,
		_w16005_,
		_w16006_,
		_w16007_,
		_w16008_
	);
	LUT3 #(
		.INIT('h80)
	) name5496 (
		\wishbone_bd_ram_mem2_reg[210][16]/P0001 ,
		_w11963_,
		_w11984_,
		_w16009_
	);
	LUT3 #(
		.INIT('h80)
	) name5497 (
		\wishbone_bd_ram_mem2_reg[198][16]/P0001 ,
		_w11945_,
		_w11986_,
		_w16010_
	);
	LUT3 #(
		.INIT('h80)
	) name5498 (
		\wishbone_bd_ram_mem2_reg[153][16]/P0001 ,
		_w11959_,
		_w11968_,
		_w16011_
	);
	LUT3 #(
		.INIT('h80)
	) name5499 (
		\wishbone_bd_ram_mem2_reg[131][16]/P0001 ,
		_w11938_,
		_w11955_,
		_w16012_
	);
	LUT4 #(
		.INIT('h0001)
	) name5500 (
		_w16009_,
		_w16010_,
		_w16011_,
		_w16012_,
		_w16013_
	);
	LUT4 #(
		.INIT('h8000)
	) name5501 (
		_w15998_,
		_w16003_,
		_w16008_,
		_w16013_,
		_w16014_
	);
	LUT3 #(
		.INIT('h80)
	) name5502 (
		\wishbone_bd_ram_mem2_reg[187][16]/P0001 ,
		_w11936_,
		_w11942_,
		_w16015_
	);
	LUT3 #(
		.INIT('h80)
	) name5503 (
		\wishbone_bd_ram_mem2_reg[68][16]/P0001 ,
		_w11929_,
		_w11949_,
		_w16016_
	);
	LUT3 #(
		.INIT('h80)
	) name5504 (
		\wishbone_bd_ram_mem2_reg[66][16]/P0001 ,
		_w11949_,
		_w11963_,
		_w16017_
	);
	LUT3 #(
		.INIT('h80)
	) name5505 (
		\wishbone_bd_ram_mem2_reg[14][16]/P0001 ,
		_w11932_,
		_w11948_,
		_w16018_
	);
	LUT4 #(
		.INIT('h0001)
	) name5506 (
		_w16015_,
		_w16016_,
		_w16017_,
		_w16018_,
		_w16019_
	);
	LUT3 #(
		.INIT('h80)
	) name5507 (
		\wishbone_bd_ram_mem2_reg[222][16]/P0001 ,
		_w11948_,
		_w11984_,
		_w16020_
	);
	LUT3 #(
		.INIT('h80)
	) name5508 (
		\wishbone_bd_ram_mem2_reg[155][16]/P0001 ,
		_w11936_,
		_w11959_,
		_w16021_
	);
	LUT3 #(
		.INIT('h80)
	) name5509 (
		\wishbone_bd_ram_mem2_reg[78][16]/P0001 ,
		_w11948_,
		_w11949_,
		_w16022_
	);
	LUT3 #(
		.INIT('h80)
	) name5510 (
		\wishbone_bd_ram_mem2_reg[177][16]/P0001 ,
		_w11942_,
		_w11977_,
		_w16023_
	);
	LUT4 #(
		.INIT('h0001)
	) name5511 (
		_w16020_,
		_w16021_,
		_w16022_,
		_w16023_,
		_w16024_
	);
	LUT3 #(
		.INIT('h80)
	) name5512 (
		\wishbone_bd_ram_mem2_reg[238][16]/P0001 ,
		_w11948_,
		_w11982_,
		_w16025_
	);
	LUT3 #(
		.INIT('h80)
	) name5513 (
		\wishbone_bd_ram_mem2_reg[5][16]/P0001 ,
		_w11932_,
		_w11933_,
		_w16026_
	);
	LUT3 #(
		.INIT('h80)
	) name5514 (
		\wishbone_bd_ram_mem2_reg[133][16]/P0001 ,
		_w11933_,
		_w11955_,
		_w16027_
	);
	LUT3 #(
		.INIT('h80)
	) name5515 (
		\wishbone_bd_ram_mem2_reg[114][16]/P0001 ,
		_w11963_,
		_w12012_,
		_w16028_
	);
	LUT4 #(
		.INIT('h0001)
	) name5516 (
		_w16025_,
		_w16026_,
		_w16027_,
		_w16028_,
		_w16029_
	);
	LUT3 #(
		.INIT('h80)
	) name5517 (
		\wishbone_bd_ram_mem2_reg[232][16]/P0001 ,
		_w11982_,
		_w11990_,
		_w16030_
	);
	LUT3 #(
		.INIT('h80)
	) name5518 (
		\wishbone_bd_ram_mem2_reg[16][16]/P0001 ,
		_w11935_,
		_w11941_,
		_w16031_
	);
	LUT3 #(
		.INIT('h80)
	) name5519 (
		\wishbone_bd_ram_mem2_reg[109][16]/P0001 ,
		_w11965_,
		_w11966_,
		_w16032_
	);
	LUT3 #(
		.INIT('h80)
	) name5520 (
		\wishbone_bd_ram_mem2_reg[216][16]/P0001 ,
		_w11984_,
		_w11990_,
		_w16033_
	);
	LUT4 #(
		.INIT('h0001)
	) name5521 (
		_w16030_,
		_w16031_,
		_w16032_,
		_w16033_,
		_w16034_
	);
	LUT4 #(
		.INIT('h8000)
	) name5522 (
		_w16019_,
		_w16024_,
		_w16029_,
		_w16034_,
		_w16035_
	);
	LUT4 #(
		.INIT('h8000)
	) name5523 (
		_w15972_,
		_w15993_,
		_w16014_,
		_w16035_,
		_w16036_
	);
	LUT3 #(
		.INIT('h80)
	) name5524 (
		\wishbone_bd_ram_mem2_reg[65][16]/P0001 ,
		_w11949_,
		_w11977_,
		_w16037_
	);
	LUT3 #(
		.INIT('h80)
	) name5525 (
		\wishbone_bd_ram_mem2_reg[207][16]/P0001 ,
		_w11945_,
		_w11973_,
		_w16038_
	);
	LUT3 #(
		.INIT('h80)
	) name5526 (
		\wishbone_bd_ram_mem2_reg[142][16]/P0001 ,
		_w11948_,
		_w11955_,
		_w16039_
	);
	LUT3 #(
		.INIT('h80)
	) name5527 (
		\wishbone_bd_ram_mem2_reg[181][16]/P0001 ,
		_w11933_,
		_w11942_,
		_w16040_
	);
	LUT4 #(
		.INIT('h0001)
	) name5528 (
		_w16037_,
		_w16038_,
		_w16039_,
		_w16040_,
		_w16041_
	);
	LUT3 #(
		.INIT('h80)
	) name5529 (
		\wishbone_bd_ram_mem2_reg[15][16]/P0001 ,
		_w11932_,
		_w11973_,
		_w16042_
	);
	LUT3 #(
		.INIT('h80)
	) name5530 (
		\wishbone_bd_ram_mem2_reg[230][16]/P0001 ,
		_w11982_,
		_w11986_,
		_w16043_
	);
	LUT3 #(
		.INIT('h80)
	) name5531 (
		\wishbone_bd_ram_mem2_reg[189][16]/P0001 ,
		_w11942_,
		_w11966_,
		_w16044_
	);
	LUT3 #(
		.INIT('h80)
	) name5532 (
		\wishbone_bd_ram_mem2_reg[243][16]/P0001 ,
		_w11938_,
		_w11952_,
		_w16045_
	);
	LUT4 #(
		.INIT('h0001)
	) name5533 (
		_w16042_,
		_w16043_,
		_w16044_,
		_w16045_,
		_w16046_
	);
	LUT3 #(
		.INIT('h80)
	) name5534 (
		\wishbone_bd_ram_mem2_reg[25][16]/P0001 ,
		_w11935_,
		_w11968_,
		_w16047_
	);
	LUT3 #(
		.INIT('h80)
	) name5535 (
		\wishbone_bd_ram_mem2_reg[97][16]/P0001 ,
		_w11965_,
		_w11977_,
		_w16048_
	);
	LUT3 #(
		.INIT('h80)
	) name5536 (
		\wishbone_bd_ram_mem2_reg[251][16]/P0001 ,
		_w11936_,
		_w11952_,
		_w16049_
	);
	LUT3 #(
		.INIT('h80)
	) name5537 (
		\wishbone_bd_ram_mem2_reg[61][16]/P0001 ,
		_w11966_,
		_w11979_,
		_w16050_
	);
	LUT4 #(
		.INIT('h0001)
	) name5538 (
		_w16047_,
		_w16048_,
		_w16049_,
		_w16050_,
		_w16051_
	);
	LUT3 #(
		.INIT('h80)
	) name5539 (
		\wishbone_bd_ram_mem2_reg[249][16]/P0001 ,
		_w11952_,
		_w11968_,
		_w16052_
	);
	LUT3 #(
		.INIT('h80)
	) name5540 (
		\wishbone_bd_ram_mem2_reg[110][16]/P0001 ,
		_w11948_,
		_w11965_,
		_w16053_
	);
	LUT3 #(
		.INIT('h80)
	) name5541 (
		\wishbone_bd_ram_mem2_reg[63][16]/P0001 ,
		_w11973_,
		_w11979_,
		_w16054_
	);
	LUT3 #(
		.INIT('h80)
	) name5542 (
		\wishbone_bd_ram_mem2_reg[104][16]/P0001 ,
		_w11965_,
		_w11990_,
		_w16055_
	);
	LUT4 #(
		.INIT('h0001)
	) name5543 (
		_w16052_,
		_w16053_,
		_w16054_,
		_w16055_,
		_w16056_
	);
	LUT4 #(
		.INIT('h8000)
	) name5544 (
		_w16041_,
		_w16046_,
		_w16051_,
		_w16056_,
		_w16057_
	);
	LUT3 #(
		.INIT('h80)
	) name5545 (
		\wishbone_bd_ram_mem2_reg[225][16]/P0001 ,
		_w11977_,
		_w11982_,
		_w16058_
	);
	LUT3 #(
		.INIT('h80)
	) name5546 (
		\wishbone_bd_ram_mem2_reg[135][16]/P0001 ,
		_w11955_,
		_w11975_,
		_w16059_
	);
	LUT3 #(
		.INIT('h80)
	) name5547 (
		\wishbone_bd_ram_mem2_reg[199][16]/P0001 ,
		_w11945_,
		_w11975_,
		_w16060_
	);
	LUT3 #(
		.INIT('h80)
	) name5548 (
		\wishbone_bd_ram_mem2_reg[186][16]/P0001 ,
		_w11942_,
		_w11944_,
		_w16061_
	);
	LUT4 #(
		.INIT('h0001)
	) name5549 (
		_w16058_,
		_w16059_,
		_w16060_,
		_w16061_,
		_w16062_
	);
	LUT3 #(
		.INIT('h80)
	) name5550 (
		\wishbone_bd_ram_mem2_reg[180][16]/P0001 ,
		_w11929_,
		_w11942_,
		_w16063_
	);
	LUT3 #(
		.INIT('h80)
	) name5551 (
		\wishbone_bd_ram_mem2_reg[167][16]/P0001 ,
		_w11930_,
		_w11975_,
		_w16064_
	);
	LUT3 #(
		.INIT('h80)
	) name5552 (
		\wishbone_bd_ram_mem2_reg[113][16]/P0001 ,
		_w11977_,
		_w12012_,
		_w16065_
	);
	LUT3 #(
		.INIT('h80)
	) name5553 (
		\wishbone_bd_ram_mem2_reg[95][16]/P0001 ,
		_w11972_,
		_w11973_,
		_w16066_
	);
	LUT4 #(
		.INIT('h0001)
	) name5554 (
		_w16063_,
		_w16064_,
		_w16065_,
		_w16066_,
		_w16067_
	);
	LUT3 #(
		.INIT('h80)
	) name5555 (
		\wishbone_bd_ram_mem2_reg[26][16]/P0001 ,
		_w11935_,
		_w11944_,
		_w16068_
	);
	LUT3 #(
		.INIT('h80)
	) name5556 (
		\wishbone_bd_ram_mem2_reg[250][16]/P0001 ,
		_w11944_,
		_w11952_,
		_w16069_
	);
	LUT3 #(
		.INIT('h80)
	) name5557 (
		\wishbone_bd_ram_mem2_reg[82][16]/P0001 ,
		_w11963_,
		_w11972_,
		_w16070_
	);
	LUT3 #(
		.INIT('h80)
	) name5558 (
		\wishbone_bd_ram_mem2_reg[248][16]/P0001 ,
		_w11952_,
		_w11990_,
		_w16071_
	);
	LUT4 #(
		.INIT('h0001)
	) name5559 (
		_w16068_,
		_w16069_,
		_w16070_,
		_w16071_,
		_w16072_
	);
	LUT3 #(
		.INIT('h80)
	) name5560 (
		\wishbone_bd_ram_mem2_reg[60][16]/P0001 ,
		_w11954_,
		_w11979_,
		_w16073_
	);
	LUT3 #(
		.INIT('h80)
	) name5561 (
		\wishbone_bd_ram_mem2_reg[35][16]/P0001 ,
		_w11938_,
		_w11957_,
		_w16074_
	);
	LUT3 #(
		.INIT('h80)
	) name5562 (
		\wishbone_bd_ram_mem2_reg[89][16]/P0001 ,
		_w11968_,
		_w11972_,
		_w16075_
	);
	LUT3 #(
		.INIT('h80)
	) name5563 (
		\wishbone_bd_ram_mem2_reg[165][16]/P0001 ,
		_w11930_,
		_w11933_,
		_w16076_
	);
	LUT4 #(
		.INIT('h0001)
	) name5564 (
		_w16073_,
		_w16074_,
		_w16075_,
		_w16076_,
		_w16077_
	);
	LUT4 #(
		.INIT('h8000)
	) name5565 (
		_w16062_,
		_w16067_,
		_w16072_,
		_w16077_,
		_w16078_
	);
	LUT3 #(
		.INIT('h80)
	) name5566 (
		\wishbone_bd_ram_mem2_reg[201][16]/P0001 ,
		_w11945_,
		_w11968_,
		_w16079_
	);
	LUT3 #(
		.INIT('h80)
	) name5567 (
		\wishbone_bd_ram_mem2_reg[208][16]/P0001 ,
		_w11941_,
		_w11984_,
		_w16080_
	);
	LUT3 #(
		.INIT('h80)
	) name5568 (
		\wishbone_bd_ram_mem2_reg[29][16]/P0001 ,
		_w11935_,
		_w11966_,
		_w16081_
	);
	LUT3 #(
		.INIT('h80)
	) name5569 (
		\wishbone_bd_ram_mem2_reg[132][16]/P0001 ,
		_w11929_,
		_w11955_,
		_w16082_
	);
	LUT4 #(
		.INIT('h0001)
	) name5570 (
		_w16079_,
		_w16080_,
		_w16081_,
		_w16082_,
		_w16083_
	);
	LUT3 #(
		.INIT('h80)
	) name5571 (
		\wishbone_bd_ram_mem2_reg[92][16]/P0001 ,
		_w11954_,
		_w11972_,
		_w16084_
	);
	LUT3 #(
		.INIT('h80)
	) name5572 (
		\wishbone_bd_ram_mem2_reg[227][16]/P0001 ,
		_w11938_,
		_w11982_,
		_w16085_
	);
	LUT3 #(
		.INIT('h80)
	) name5573 (
		\wishbone_bd_ram_mem2_reg[245][16]/P0001 ,
		_w11933_,
		_w11952_,
		_w16086_
	);
	LUT3 #(
		.INIT('h80)
	) name5574 (
		\wishbone_bd_ram_mem2_reg[111][16]/P0001 ,
		_w11965_,
		_w11973_,
		_w16087_
	);
	LUT4 #(
		.INIT('h0001)
	) name5575 (
		_w16084_,
		_w16085_,
		_w16086_,
		_w16087_,
		_w16088_
	);
	LUT3 #(
		.INIT('h80)
	) name5576 (
		\wishbone_bd_ram_mem2_reg[12][16]/P0001 ,
		_w11932_,
		_w11954_,
		_w16089_
	);
	LUT3 #(
		.INIT('h80)
	) name5577 (
		\wishbone_bd_ram_mem2_reg[90][16]/P0001 ,
		_w11944_,
		_w11972_,
		_w16090_
	);
	LUT3 #(
		.INIT('h80)
	) name5578 (
		\wishbone_bd_ram_mem2_reg[85][16]/P0001 ,
		_w11933_,
		_w11972_,
		_w16091_
	);
	LUT3 #(
		.INIT('h80)
	) name5579 (
		\wishbone_bd_ram_mem2_reg[87][16]/P0001 ,
		_w11972_,
		_w11975_,
		_w16092_
	);
	LUT4 #(
		.INIT('h0001)
	) name5580 (
		_w16089_,
		_w16090_,
		_w16091_,
		_w16092_,
		_w16093_
	);
	LUT3 #(
		.INIT('h80)
	) name5581 (
		\wishbone_bd_ram_mem2_reg[212][16]/P0001 ,
		_w11929_,
		_w11984_,
		_w16094_
	);
	LUT3 #(
		.INIT('h80)
	) name5582 (
		\wishbone_bd_ram_mem2_reg[173][16]/P0001 ,
		_w11930_,
		_w11966_,
		_w16095_
	);
	LUT3 #(
		.INIT('h80)
	) name5583 (
		\wishbone_bd_ram_mem2_reg[43][16]/P0001 ,
		_w11936_,
		_w11957_,
		_w16096_
	);
	LUT3 #(
		.INIT('h80)
	) name5584 (
		\wishbone_bd_ram_mem2_reg[233][16]/P0001 ,
		_w11968_,
		_w11982_,
		_w16097_
	);
	LUT4 #(
		.INIT('h0001)
	) name5585 (
		_w16094_,
		_w16095_,
		_w16096_,
		_w16097_,
		_w16098_
	);
	LUT4 #(
		.INIT('h8000)
	) name5586 (
		_w16083_,
		_w16088_,
		_w16093_,
		_w16098_,
		_w16099_
	);
	LUT3 #(
		.INIT('h80)
	) name5587 (
		\wishbone_bd_ram_mem2_reg[76][16]/P0001 ,
		_w11949_,
		_w11954_,
		_w16100_
	);
	LUT3 #(
		.INIT('h80)
	) name5588 (
		\wishbone_bd_ram_mem2_reg[106][16]/P0001 ,
		_w11944_,
		_w11965_,
		_w16101_
	);
	LUT3 #(
		.INIT('h80)
	) name5589 (
		\wishbone_bd_ram_mem2_reg[228][16]/P0001 ,
		_w11929_,
		_w11982_,
		_w16102_
	);
	LUT3 #(
		.INIT('h80)
	) name5590 (
		\wishbone_bd_ram_mem2_reg[169][16]/P0001 ,
		_w11930_,
		_w11968_,
		_w16103_
	);
	LUT4 #(
		.INIT('h0001)
	) name5591 (
		_w16100_,
		_w16101_,
		_w16102_,
		_w16103_,
		_w16104_
	);
	LUT3 #(
		.INIT('h80)
	) name5592 (
		\wishbone_bd_ram_mem2_reg[209][16]/P0001 ,
		_w11977_,
		_w11984_,
		_w16105_
	);
	LUT3 #(
		.INIT('h80)
	) name5593 (
		\wishbone_bd_ram_mem2_reg[178][16]/P0001 ,
		_w11942_,
		_w11963_,
		_w16106_
	);
	LUT3 #(
		.INIT('h80)
	) name5594 (
		\wishbone_bd_ram_mem2_reg[205][16]/P0001 ,
		_w11945_,
		_w11966_,
		_w16107_
	);
	LUT3 #(
		.INIT('h80)
	) name5595 (
		\wishbone_bd_ram_mem2_reg[141][16]/P0001 ,
		_w11955_,
		_w11966_,
		_w16108_
	);
	LUT4 #(
		.INIT('h0001)
	) name5596 (
		_w16105_,
		_w16106_,
		_w16107_,
		_w16108_,
		_w16109_
	);
	LUT3 #(
		.INIT('h80)
	) name5597 (
		\wishbone_bd_ram_mem2_reg[140][16]/P0001 ,
		_w11954_,
		_w11955_,
		_w16110_
	);
	LUT3 #(
		.INIT('h80)
	) name5598 (
		\wishbone_bd_ram_mem2_reg[56][16]/P0001 ,
		_w11979_,
		_w11990_,
		_w16111_
	);
	LUT3 #(
		.INIT('h80)
	) name5599 (
		\wishbone_bd_ram_mem2_reg[175][16]/P0001 ,
		_w11930_,
		_w11973_,
		_w16112_
	);
	LUT3 #(
		.INIT('h80)
	) name5600 (
		\wishbone_bd_ram_mem2_reg[46][16]/P0001 ,
		_w11948_,
		_w11957_,
		_w16113_
	);
	LUT4 #(
		.INIT('h0001)
	) name5601 (
		_w16110_,
		_w16111_,
		_w16112_,
		_w16113_,
		_w16114_
	);
	LUT3 #(
		.INIT('h80)
	) name5602 (
		\wishbone_bd_ram_mem2_reg[195][16]/P0001 ,
		_w11938_,
		_w11945_,
		_w16115_
	);
	LUT3 #(
		.INIT('h80)
	) name5603 (
		\wishbone_bd_ram_mem2_reg[119][16]/P0001 ,
		_w11975_,
		_w12012_,
		_w16116_
	);
	LUT3 #(
		.INIT('h80)
	) name5604 (
		\wishbone_bd_ram_mem2_reg[171][16]/P0001 ,
		_w11930_,
		_w11936_,
		_w16117_
	);
	LUT3 #(
		.INIT('h80)
	) name5605 (
		\wishbone_bd_ram_mem2_reg[226][16]/P0001 ,
		_w11963_,
		_w11982_,
		_w16118_
	);
	LUT4 #(
		.INIT('h0001)
	) name5606 (
		_w16115_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16119_
	);
	LUT4 #(
		.INIT('h8000)
	) name5607 (
		_w16104_,
		_w16109_,
		_w16114_,
		_w16119_,
		_w16120_
	);
	LUT4 #(
		.INIT('h8000)
	) name5608 (
		_w16057_,
		_w16078_,
		_w16099_,
		_w16120_,
		_w16121_
	);
	LUT4 #(
		.INIT('h8000)
	) name5609 (
		_w15866_,
		_w15951_,
		_w16036_,
		_w16121_,
		_w16122_
	);
	LUT2 #(
		.INIT('h6)
	) name5610 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		_w16123_
	);
	LUT3 #(
		.INIT('h40)
	) name5611 (
		_w12302_,
		_w12304_,
		_w16123_,
		_w16124_
	);
	LUT3 #(
		.INIT('h70)
	) name5612 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_TxLength_reg[0]/NET0131 ,
		_w16125_
	);
	LUT2 #(
		.INIT('h4)
	) name5613 (
		_w12302_,
		_w16125_,
		_w16126_
	);
	LUT4 #(
		.INIT('h008f)
	) name5614 (
		_w12312_,
		_w12317_,
		_w16124_,
		_w16126_,
		_w16127_
	);
	LUT3 #(
		.INIT('h2f)
	) name5615 (
		_w12303_,
		_w16122_,
		_w16127_,
		_w16128_
	);
	LUT3 #(
		.INIT('h80)
	) name5616 (
		\wishbone_bd_ram_mem3_reg[128][31]/P0001 ,
		_w11941_,
		_w11955_,
		_w16129_
	);
	LUT3 #(
		.INIT('h80)
	) name5617 (
		\wishbone_bd_ram_mem3_reg[68][31]/P0001 ,
		_w11929_,
		_w11949_,
		_w16130_
	);
	LUT3 #(
		.INIT('h80)
	) name5618 (
		\wishbone_bd_ram_mem3_reg[52][31]/P0001 ,
		_w11929_,
		_w11979_,
		_w16131_
	);
	LUT3 #(
		.INIT('h80)
	) name5619 (
		\wishbone_bd_ram_mem3_reg[7][31]/P0001 ,
		_w11932_,
		_w11975_,
		_w16132_
	);
	LUT4 #(
		.INIT('h0001)
	) name5620 (
		_w16129_,
		_w16130_,
		_w16131_,
		_w16132_,
		_w16133_
	);
	LUT3 #(
		.INIT('h80)
	) name5621 (
		\wishbone_bd_ram_mem3_reg[184][31]/P0001 ,
		_w11942_,
		_w11990_,
		_w16134_
	);
	LUT3 #(
		.INIT('h80)
	) name5622 (
		\wishbone_bd_ram_mem3_reg[139][31]/P0001 ,
		_w11936_,
		_w11955_,
		_w16135_
	);
	LUT3 #(
		.INIT('h80)
	) name5623 (
		\wishbone_bd_ram_mem3_reg[39][31]/P0001 ,
		_w11957_,
		_w11975_,
		_w16136_
	);
	LUT3 #(
		.INIT('h80)
	) name5624 (
		\wishbone_bd_ram_mem3_reg[220][31]/P0001 ,
		_w11954_,
		_w11984_,
		_w16137_
	);
	LUT4 #(
		.INIT('h0001)
	) name5625 (
		_w16134_,
		_w16135_,
		_w16136_,
		_w16137_,
		_w16138_
	);
	LUT3 #(
		.INIT('h80)
	) name5626 (
		\wishbone_bd_ram_mem3_reg[226][31]/P0001 ,
		_w11963_,
		_w11982_,
		_w16139_
	);
	LUT3 #(
		.INIT('h80)
	) name5627 (
		\wishbone_bd_ram_mem3_reg[247][31]/P0001 ,
		_w11952_,
		_w11975_,
		_w16140_
	);
	LUT3 #(
		.INIT('h80)
	) name5628 (
		\wishbone_bd_ram_mem3_reg[85][31]/P0001 ,
		_w11933_,
		_w11972_,
		_w16141_
	);
	LUT3 #(
		.INIT('h80)
	) name5629 (
		\wishbone_bd_ram_mem3_reg[193][31]/P0001 ,
		_w11945_,
		_w11977_,
		_w16142_
	);
	LUT4 #(
		.INIT('h0001)
	) name5630 (
		_w16139_,
		_w16140_,
		_w16141_,
		_w16142_,
		_w16143_
	);
	LUT3 #(
		.INIT('h80)
	) name5631 (
		\wishbone_bd_ram_mem3_reg[66][31]/P0001 ,
		_w11949_,
		_w11963_,
		_w16144_
	);
	LUT3 #(
		.INIT('h80)
	) name5632 (
		\wishbone_bd_ram_mem3_reg[227][31]/P0001 ,
		_w11938_,
		_w11982_,
		_w16145_
	);
	LUT3 #(
		.INIT('h80)
	) name5633 (
		\wishbone_bd_ram_mem3_reg[25][31]/P0001 ,
		_w11935_,
		_w11968_,
		_w16146_
	);
	LUT3 #(
		.INIT('h80)
	) name5634 (
		\wishbone_bd_ram_mem3_reg[180][31]/P0001 ,
		_w11929_,
		_w11942_,
		_w16147_
	);
	LUT4 #(
		.INIT('h0001)
	) name5635 (
		_w16144_,
		_w16145_,
		_w16146_,
		_w16147_,
		_w16148_
	);
	LUT4 #(
		.INIT('h8000)
	) name5636 (
		_w16133_,
		_w16138_,
		_w16143_,
		_w16148_,
		_w16149_
	);
	LUT3 #(
		.INIT('h80)
	) name5637 (
		\wishbone_bd_ram_mem3_reg[89][31]/P0001 ,
		_w11968_,
		_w11972_,
		_w16150_
	);
	LUT3 #(
		.INIT('h80)
	) name5638 (
		\wishbone_bd_ram_mem3_reg[186][31]/P0001 ,
		_w11942_,
		_w11944_,
		_w16151_
	);
	LUT3 #(
		.INIT('h80)
	) name5639 (
		\wishbone_bd_ram_mem3_reg[13][31]/P0001 ,
		_w11932_,
		_w11966_,
		_w16152_
	);
	LUT3 #(
		.INIT('h80)
	) name5640 (
		\wishbone_bd_ram_mem3_reg[93][31]/P0001 ,
		_w11966_,
		_w11972_,
		_w16153_
	);
	LUT4 #(
		.INIT('h0001)
	) name5641 (
		_w16150_,
		_w16151_,
		_w16152_,
		_w16153_,
		_w16154_
	);
	LUT3 #(
		.INIT('h80)
	) name5642 (
		\wishbone_bd_ram_mem3_reg[240][31]/P0001 ,
		_w11941_,
		_w11952_,
		_w16155_
	);
	LUT3 #(
		.INIT('h80)
	) name5643 (
		\wishbone_bd_ram_mem3_reg[185][31]/P0001 ,
		_w11942_,
		_w11968_,
		_w16156_
	);
	LUT3 #(
		.INIT('h80)
	) name5644 (
		\wishbone_bd_ram_mem3_reg[15][31]/P0001 ,
		_w11932_,
		_w11973_,
		_w16157_
	);
	LUT3 #(
		.INIT('h80)
	) name5645 (
		\wishbone_bd_ram_mem3_reg[17][31]/P0001 ,
		_w11935_,
		_w11977_,
		_w16158_
	);
	LUT4 #(
		.INIT('h0001)
	) name5646 (
		_w16155_,
		_w16156_,
		_w16157_,
		_w16158_,
		_w16159_
	);
	LUT3 #(
		.INIT('h80)
	) name5647 (
		\wishbone_bd_ram_mem3_reg[121][31]/P0001 ,
		_w11968_,
		_w12012_,
		_w16160_
	);
	LUT3 #(
		.INIT('h80)
	) name5648 (
		\wishbone_bd_ram_mem3_reg[187][31]/P0001 ,
		_w11936_,
		_w11942_,
		_w16161_
	);
	LUT3 #(
		.INIT('h80)
	) name5649 (
		\wishbone_bd_ram_mem3_reg[245][31]/P0001 ,
		_w11933_,
		_w11952_,
		_w16162_
	);
	LUT3 #(
		.INIT('h80)
	) name5650 (
		\wishbone_bd_ram_mem3_reg[72][31]/P0001 ,
		_w11949_,
		_w11990_,
		_w16163_
	);
	LUT4 #(
		.INIT('h0001)
	) name5651 (
		_w16160_,
		_w16161_,
		_w16162_,
		_w16163_,
		_w16164_
	);
	LUT3 #(
		.INIT('h80)
	) name5652 (
		\wishbone_bd_ram_mem3_reg[69][31]/P0001 ,
		_w11933_,
		_w11949_,
		_w16165_
	);
	LUT3 #(
		.INIT('h80)
	) name5653 (
		\wishbone_bd_ram_mem3_reg[179][31]/P0001 ,
		_w11938_,
		_w11942_,
		_w16166_
	);
	LUT3 #(
		.INIT('h80)
	) name5654 (
		\wishbone_bd_ram_mem3_reg[107][31]/P0001 ,
		_w11936_,
		_w11965_,
		_w16167_
	);
	LUT3 #(
		.INIT('h80)
	) name5655 (
		\wishbone_bd_ram_mem3_reg[254][31]/P0001 ,
		_w11948_,
		_w11952_,
		_w16168_
	);
	LUT4 #(
		.INIT('h0001)
	) name5656 (
		_w16165_,
		_w16166_,
		_w16167_,
		_w16168_,
		_w16169_
	);
	LUT4 #(
		.INIT('h8000)
	) name5657 (
		_w16154_,
		_w16159_,
		_w16164_,
		_w16169_,
		_w16170_
	);
	LUT3 #(
		.INIT('h80)
	) name5658 (
		\wishbone_bd_ram_mem3_reg[235][31]/P0001 ,
		_w11936_,
		_w11982_,
		_w16171_
	);
	LUT3 #(
		.INIT('h80)
	) name5659 (
		\wishbone_bd_ram_mem3_reg[218][31]/P0001 ,
		_w11944_,
		_w11984_,
		_w16172_
	);
	LUT3 #(
		.INIT('h80)
	) name5660 (
		\wishbone_bd_ram_mem3_reg[132][31]/P0001 ,
		_w11929_,
		_w11955_,
		_w16173_
	);
	LUT3 #(
		.INIT('h80)
	) name5661 (
		\wishbone_bd_ram_mem3_reg[0][31]/P0001 ,
		_w11932_,
		_w11941_,
		_w16174_
	);
	LUT4 #(
		.INIT('h0001)
	) name5662 (
		_w16171_,
		_w16172_,
		_w16173_,
		_w16174_,
		_w16175_
	);
	LUT3 #(
		.INIT('h80)
	) name5663 (
		\wishbone_bd_ram_mem3_reg[173][31]/P0001 ,
		_w11930_,
		_w11966_,
		_w16176_
	);
	LUT3 #(
		.INIT('h80)
	) name5664 (
		\wishbone_bd_ram_mem3_reg[57][31]/P0001 ,
		_w11968_,
		_w11979_,
		_w16177_
	);
	LUT3 #(
		.INIT('h80)
	) name5665 (
		\wishbone_bd_ram_mem3_reg[238][31]/P0001 ,
		_w11948_,
		_w11982_,
		_w16178_
	);
	LUT3 #(
		.INIT('h80)
	) name5666 (
		\wishbone_bd_ram_mem3_reg[189][31]/P0001 ,
		_w11942_,
		_w11966_,
		_w16179_
	);
	LUT4 #(
		.INIT('h0001)
	) name5667 (
		_w16176_,
		_w16177_,
		_w16178_,
		_w16179_,
		_w16180_
	);
	LUT3 #(
		.INIT('h80)
	) name5668 (
		\wishbone_bd_ram_mem3_reg[88][31]/P0001 ,
		_w11972_,
		_w11990_,
		_w16181_
	);
	LUT3 #(
		.INIT('h80)
	) name5669 (
		\wishbone_bd_ram_mem3_reg[14][31]/P0001 ,
		_w11932_,
		_w11948_,
		_w16182_
	);
	LUT3 #(
		.INIT('h80)
	) name5670 (
		\wishbone_bd_ram_mem3_reg[155][31]/P0001 ,
		_w11936_,
		_w11959_,
		_w16183_
	);
	LUT3 #(
		.INIT('h80)
	) name5671 (
		\wishbone_bd_ram_mem3_reg[210][31]/P0001 ,
		_w11963_,
		_w11984_,
		_w16184_
	);
	LUT4 #(
		.INIT('h0001)
	) name5672 (
		_w16181_,
		_w16182_,
		_w16183_,
		_w16184_,
		_w16185_
	);
	LUT3 #(
		.INIT('h80)
	) name5673 (
		\wishbone_bd_ram_mem3_reg[232][31]/P0001 ,
		_w11982_,
		_w11990_,
		_w16186_
	);
	LUT3 #(
		.INIT('h80)
	) name5674 (
		\wishbone_bd_ram_mem3_reg[221][31]/P0001 ,
		_w11966_,
		_w11984_,
		_w16187_
	);
	LUT3 #(
		.INIT('h80)
	) name5675 (
		\wishbone_bd_ram_mem3_reg[34][31]/P0001 ,
		_w11957_,
		_w11963_,
		_w16188_
	);
	LUT3 #(
		.INIT('h80)
	) name5676 (
		\wishbone_bd_ram_mem3_reg[239][31]/P0001 ,
		_w11973_,
		_w11982_,
		_w16189_
	);
	LUT4 #(
		.INIT('h0001)
	) name5677 (
		_w16186_,
		_w16187_,
		_w16188_,
		_w16189_,
		_w16190_
	);
	LUT4 #(
		.INIT('h8000)
	) name5678 (
		_w16175_,
		_w16180_,
		_w16185_,
		_w16190_,
		_w16191_
	);
	LUT3 #(
		.INIT('h80)
	) name5679 (
		\wishbone_bd_ram_mem3_reg[82][31]/P0001 ,
		_w11963_,
		_w11972_,
		_w16192_
	);
	LUT3 #(
		.INIT('h80)
	) name5680 (
		\wishbone_bd_ram_mem3_reg[103][31]/P0001 ,
		_w11965_,
		_w11975_,
		_w16193_
	);
	LUT3 #(
		.INIT('h80)
	) name5681 (
		\wishbone_bd_ram_mem3_reg[145][31]/P0001 ,
		_w11959_,
		_w11977_,
		_w16194_
	);
	LUT3 #(
		.INIT('h80)
	) name5682 (
		\wishbone_bd_ram_mem3_reg[104][31]/P0001 ,
		_w11965_,
		_w11990_,
		_w16195_
	);
	LUT4 #(
		.INIT('h0001)
	) name5683 (
		_w16192_,
		_w16193_,
		_w16194_,
		_w16195_,
		_w16196_
	);
	LUT3 #(
		.INIT('h80)
	) name5684 (
		\wishbone_bd_ram_mem3_reg[216][31]/P0001 ,
		_w11984_,
		_w11990_,
		_w16197_
	);
	LUT3 #(
		.INIT('h80)
	) name5685 (
		\wishbone_bd_ram_mem3_reg[170][31]/P0001 ,
		_w11930_,
		_w11944_,
		_w16198_
	);
	LUT3 #(
		.INIT('h80)
	) name5686 (
		\wishbone_bd_ram_mem3_reg[28][31]/P0001 ,
		_w11935_,
		_w11954_,
		_w16199_
	);
	LUT3 #(
		.INIT('h80)
	) name5687 (
		\wishbone_bd_ram_mem3_reg[42][31]/P0001 ,
		_w11944_,
		_w11957_,
		_w16200_
	);
	LUT4 #(
		.INIT('h0001)
	) name5688 (
		_w16197_,
		_w16198_,
		_w16199_,
		_w16200_,
		_w16201_
	);
	LUT3 #(
		.INIT('h80)
	) name5689 (
		\wishbone_bd_ram_mem3_reg[111][31]/P0001 ,
		_w11965_,
		_w11973_,
		_w16202_
	);
	LUT3 #(
		.INIT('h80)
	) name5690 (
		\wishbone_bd_ram_mem3_reg[60][31]/P0001 ,
		_w11954_,
		_w11979_,
		_w16203_
	);
	LUT3 #(
		.INIT('h80)
	) name5691 (
		\wishbone_bd_ram_mem3_reg[71][31]/P0001 ,
		_w11949_,
		_w11975_,
		_w16204_
	);
	LUT3 #(
		.INIT('h80)
	) name5692 (
		\wishbone_bd_ram_mem3_reg[119][31]/P0001 ,
		_w11975_,
		_w12012_,
		_w16205_
	);
	LUT4 #(
		.INIT('h0001)
	) name5693 (
		_w16202_,
		_w16203_,
		_w16204_,
		_w16205_,
		_w16206_
	);
	LUT3 #(
		.INIT('h80)
	) name5694 (
		\wishbone_bd_ram_mem3_reg[55][31]/P0001 ,
		_w11975_,
		_w11979_,
		_w16207_
	);
	LUT3 #(
		.INIT('h80)
	) name5695 (
		\wishbone_bd_ram_mem3_reg[51][31]/P0001 ,
		_w11938_,
		_w11979_,
		_w16208_
	);
	LUT3 #(
		.INIT('h80)
	) name5696 (
		\wishbone_bd_ram_mem3_reg[30][31]/P0001 ,
		_w11935_,
		_w11948_,
		_w16209_
	);
	LUT3 #(
		.INIT('h80)
	) name5697 (
		\wishbone_bd_ram_mem3_reg[144][31]/P0001 ,
		_w11941_,
		_w11959_,
		_w16210_
	);
	LUT4 #(
		.INIT('h0001)
	) name5698 (
		_w16207_,
		_w16208_,
		_w16209_,
		_w16210_,
		_w16211_
	);
	LUT4 #(
		.INIT('h8000)
	) name5699 (
		_w16196_,
		_w16201_,
		_w16206_,
		_w16211_,
		_w16212_
	);
	LUT4 #(
		.INIT('h8000)
	) name5700 (
		_w16149_,
		_w16170_,
		_w16191_,
		_w16212_,
		_w16213_
	);
	LUT3 #(
		.INIT('h80)
	) name5701 (
		\wishbone_bd_ram_mem3_reg[160][31]/P0001 ,
		_w11930_,
		_w11941_,
		_w16214_
	);
	LUT3 #(
		.INIT('h80)
	) name5702 (
		\wishbone_bd_ram_mem3_reg[234][31]/P0001 ,
		_w11944_,
		_w11982_,
		_w16215_
	);
	LUT3 #(
		.INIT('h80)
	) name5703 (
		\wishbone_bd_ram_mem3_reg[183][31]/P0001 ,
		_w11942_,
		_w11975_,
		_w16216_
	);
	LUT3 #(
		.INIT('h80)
	) name5704 (
		\wishbone_bd_ram_mem3_reg[182][31]/P0001 ,
		_w11942_,
		_w11986_,
		_w16217_
	);
	LUT4 #(
		.INIT('h0001)
	) name5705 (
		_w16214_,
		_w16215_,
		_w16216_,
		_w16217_,
		_w16218_
	);
	LUT3 #(
		.INIT('h80)
	) name5706 (
		\wishbone_bd_ram_mem3_reg[113][31]/P0001 ,
		_w11977_,
		_w12012_,
		_w16219_
	);
	LUT3 #(
		.INIT('h80)
	) name5707 (
		\wishbone_bd_ram_mem3_reg[94][31]/P0001 ,
		_w11948_,
		_w11972_,
		_w16220_
	);
	LUT3 #(
		.INIT('h80)
	) name5708 (
		\wishbone_bd_ram_mem3_reg[47][31]/P0001 ,
		_w11957_,
		_w11973_,
		_w16221_
	);
	LUT3 #(
		.INIT('h80)
	) name5709 (
		\wishbone_bd_ram_mem3_reg[37][31]/P0001 ,
		_w11933_,
		_w11957_,
		_w16222_
	);
	LUT4 #(
		.INIT('h0001)
	) name5710 (
		_w16219_,
		_w16220_,
		_w16221_,
		_w16222_,
		_w16223_
	);
	LUT3 #(
		.INIT('h80)
	) name5711 (
		\wishbone_bd_ram_mem3_reg[105][31]/P0001 ,
		_w11965_,
		_w11968_,
		_w16224_
	);
	LUT3 #(
		.INIT('h80)
	) name5712 (
		\wishbone_bd_ram_mem3_reg[45][31]/P0001 ,
		_w11957_,
		_w11966_,
		_w16225_
	);
	LUT3 #(
		.INIT('h80)
	) name5713 (
		\wishbone_bd_ram_mem3_reg[172][31]/P0001 ,
		_w11930_,
		_w11954_,
		_w16226_
	);
	LUT3 #(
		.INIT('h80)
	) name5714 (
		\wishbone_bd_ram_mem3_reg[200][31]/P0001 ,
		_w11945_,
		_w11990_,
		_w16227_
	);
	LUT4 #(
		.INIT('h0001)
	) name5715 (
		_w16224_,
		_w16225_,
		_w16226_,
		_w16227_,
		_w16228_
	);
	LUT3 #(
		.INIT('h80)
	) name5716 (
		\wishbone_bd_ram_mem3_reg[228][31]/P0001 ,
		_w11929_,
		_w11982_,
		_w16229_
	);
	LUT3 #(
		.INIT('h80)
	) name5717 (
		\wishbone_bd_ram_mem3_reg[118][31]/P0001 ,
		_w11986_,
		_w12012_,
		_w16230_
	);
	LUT3 #(
		.INIT('h80)
	) name5718 (
		\wishbone_bd_ram_mem3_reg[230][31]/P0001 ,
		_w11982_,
		_w11986_,
		_w16231_
	);
	LUT3 #(
		.INIT('h80)
	) name5719 (
		\wishbone_bd_ram_mem3_reg[202][31]/P0001 ,
		_w11944_,
		_w11945_,
		_w16232_
	);
	LUT4 #(
		.INIT('h0001)
	) name5720 (
		_w16229_,
		_w16230_,
		_w16231_,
		_w16232_,
		_w16233_
	);
	LUT4 #(
		.INIT('h8000)
	) name5721 (
		_w16218_,
		_w16223_,
		_w16228_,
		_w16233_,
		_w16234_
	);
	LUT3 #(
		.INIT('h80)
	) name5722 (
		\wishbone_bd_ram_mem3_reg[157][31]/P0001 ,
		_w11959_,
		_w11966_,
		_w16235_
	);
	LUT3 #(
		.INIT('h80)
	) name5723 (
		\wishbone_bd_ram_mem3_reg[244][31]/P0001 ,
		_w11929_,
		_w11952_,
		_w16236_
	);
	LUT3 #(
		.INIT('h80)
	) name5724 (
		\wishbone_bd_ram_mem3_reg[84][31]/P0001 ,
		_w11929_,
		_w11972_,
		_w16237_
	);
	LUT3 #(
		.INIT('h80)
	) name5725 (
		\wishbone_bd_ram_mem3_reg[109][31]/P0001 ,
		_w11965_,
		_w11966_,
		_w16238_
	);
	LUT4 #(
		.INIT('h0001)
	) name5726 (
		_w16235_,
		_w16236_,
		_w16237_,
		_w16238_,
		_w16239_
	);
	LUT3 #(
		.INIT('h80)
	) name5727 (
		\wishbone_bd_ram_mem3_reg[67][31]/P0001 ,
		_w11938_,
		_w11949_,
		_w16240_
	);
	LUT3 #(
		.INIT('h80)
	) name5728 (
		\wishbone_bd_ram_mem3_reg[38][31]/P0001 ,
		_w11957_,
		_w11986_,
		_w16241_
	);
	LUT3 #(
		.INIT('h80)
	) name5729 (
		\wishbone_bd_ram_mem3_reg[58][31]/P0001 ,
		_w11944_,
		_w11979_,
		_w16242_
	);
	LUT3 #(
		.INIT('h80)
	) name5730 (
		\wishbone_bd_ram_mem3_reg[143][31]/P0001 ,
		_w11955_,
		_w11973_,
		_w16243_
	);
	LUT4 #(
		.INIT('h0001)
	) name5731 (
		_w16240_,
		_w16241_,
		_w16242_,
		_w16243_,
		_w16244_
	);
	LUT3 #(
		.INIT('h80)
	) name5732 (
		\wishbone_bd_ram_mem3_reg[43][31]/P0001 ,
		_w11936_,
		_w11957_,
		_w16245_
	);
	LUT3 #(
		.INIT('h80)
	) name5733 (
		\wishbone_bd_ram_mem3_reg[133][31]/P0001 ,
		_w11933_,
		_w11955_,
		_w16246_
	);
	LUT3 #(
		.INIT('h80)
	) name5734 (
		\wishbone_bd_ram_mem3_reg[161][31]/P0001 ,
		_w11930_,
		_w11977_,
		_w16247_
	);
	LUT3 #(
		.INIT('h80)
	) name5735 (
		\wishbone_bd_ram_mem3_reg[48][31]/P0001 ,
		_w11941_,
		_w11979_,
		_w16248_
	);
	LUT4 #(
		.INIT('h0001)
	) name5736 (
		_w16245_,
		_w16246_,
		_w16247_,
		_w16248_,
		_w16249_
	);
	LUT3 #(
		.INIT('h80)
	) name5737 (
		\wishbone_bd_ram_mem3_reg[192][31]/P0001 ,
		_w11941_,
		_w11945_,
		_w16250_
	);
	LUT3 #(
		.INIT('h80)
	) name5738 (
		\wishbone_bd_ram_mem3_reg[190][31]/P0001 ,
		_w11942_,
		_w11948_,
		_w16251_
	);
	LUT3 #(
		.INIT('h80)
	) name5739 (
		\wishbone_bd_ram_mem3_reg[242][31]/P0001 ,
		_w11952_,
		_w11963_,
		_w16252_
	);
	LUT3 #(
		.INIT('h80)
	) name5740 (
		\wishbone_bd_ram_mem3_reg[87][31]/P0001 ,
		_w11972_,
		_w11975_,
		_w16253_
	);
	LUT4 #(
		.INIT('h0001)
	) name5741 (
		_w16250_,
		_w16251_,
		_w16252_,
		_w16253_,
		_w16254_
	);
	LUT4 #(
		.INIT('h8000)
	) name5742 (
		_w16239_,
		_w16244_,
		_w16249_,
		_w16254_,
		_w16255_
	);
	LUT3 #(
		.INIT('h80)
	) name5743 (
		\wishbone_bd_ram_mem3_reg[41][31]/P0001 ,
		_w11957_,
		_w11968_,
		_w16256_
	);
	LUT3 #(
		.INIT('h80)
	) name5744 (
		\wishbone_bd_ram_mem3_reg[241][31]/P0001 ,
		_w11952_,
		_w11977_,
		_w16257_
	);
	LUT3 #(
		.INIT('h80)
	) name5745 (
		\wishbone_bd_ram_mem3_reg[171][31]/P0001 ,
		_w11930_,
		_w11936_,
		_w16258_
	);
	LUT3 #(
		.INIT('h80)
	) name5746 (
		\wishbone_bd_ram_mem3_reg[197][31]/P0001 ,
		_w11933_,
		_w11945_,
		_w16259_
	);
	LUT4 #(
		.INIT('h0001)
	) name5747 (
		_w16256_,
		_w16257_,
		_w16258_,
		_w16259_,
		_w16260_
	);
	LUT3 #(
		.INIT('h80)
	) name5748 (
		\wishbone_bd_ram_mem3_reg[203][31]/P0001 ,
		_w11936_,
		_w11945_,
		_w16261_
	);
	LUT3 #(
		.INIT('h80)
	) name5749 (
		\wishbone_bd_ram_mem3_reg[252][31]/P0001 ,
		_w11952_,
		_w11954_,
		_w16262_
	);
	LUT3 #(
		.INIT('h80)
	) name5750 (
		\wishbone_bd_ram_mem3_reg[3][31]/P0001 ,
		_w11932_,
		_w11938_,
		_w16263_
	);
	LUT3 #(
		.INIT('h80)
	) name5751 (
		\wishbone_bd_ram_mem3_reg[149][31]/P0001 ,
		_w11933_,
		_w11959_,
		_w16264_
	);
	LUT4 #(
		.INIT('h0001)
	) name5752 (
		_w16261_,
		_w16262_,
		_w16263_,
		_w16264_,
		_w16265_
	);
	LUT3 #(
		.INIT('h80)
	) name5753 (
		\wishbone_bd_ram_mem3_reg[191][31]/P0001 ,
		_w11942_,
		_w11973_,
		_w16266_
	);
	LUT3 #(
		.INIT('h80)
	) name5754 (
		\wishbone_bd_ram_mem3_reg[29][31]/P0001 ,
		_w11935_,
		_w11966_,
		_w16267_
	);
	LUT3 #(
		.INIT('h80)
	) name5755 (
		\wishbone_bd_ram_mem3_reg[188][31]/P0001 ,
		_w11942_,
		_w11954_,
		_w16268_
	);
	LUT3 #(
		.INIT('h80)
	) name5756 (
		\wishbone_bd_ram_mem3_reg[127][31]/P0001 ,
		_w11973_,
		_w12012_,
		_w16269_
	);
	LUT4 #(
		.INIT('h0001)
	) name5757 (
		_w16266_,
		_w16267_,
		_w16268_,
		_w16269_,
		_w16270_
	);
	LUT3 #(
		.INIT('h80)
	) name5758 (
		\wishbone_bd_ram_mem3_reg[174][31]/P0001 ,
		_w11930_,
		_w11948_,
		_w16271_
	);
	LUT3 #(
		.INIT('h80)
	) name5759 (
		\wishbone_bd_ram_mem3_reg[248][31]/P0001 ,
		_w11952_,
		_w11990_,
		_w16272_
	);
	LUT3 #(
		.INIT('h80)
	) name5760 (
		\wishbone_bd_ram_mem3_reg[168][31]/P0001 ,
		_w11930_,
		_w11990_,
		_w16273_
	);
	LUT3 #(
		.INIT('h80)
	) name5761 (
		\wishbone_bd_ram_mem3_reg[150][31]/P0001 ,
		_w11959_,
		_w11986_,
		_w16274_
	);
	LUT4 #(
		.INIT('h0001)
	) name5762 (
		_w16271_,
		_w16272_,
		_w16273_,
		_w16274_,
		_w16275_
	);
	LUT4 #(
		.INIT('h8000)
	) name5763 (
		_w16260_,
		_w16265_,
		_w16270_,
		_w16275_,
		_w16276_
	);
	LUT3 #(
		.INIT('h80)
	) name5764 (
		\wishbone_bd_ram_mem3_reg[135][31]/P0001 ,
		_w11955_,
		_w11975_,
		_w16277_
	);
	LUT3 #(
		.INIT('h80)
	) name5765 (
		\wishbone_bd_ram_mem3_reg[136][31]/P0001 ,
		_w11955_,
		_w11990_,
		_w16278_
	);
	LUT3 #(
		.INIT('h80)
	) name5766 (
		\wishbone_bd_ram_mem3_reg[97][31]/P0001 ,
		_w11965_,
		_w11977_,
		_w16279_
	);
	LUT3 #(
		.INIT('h80)
	) name5767 (
		\wishbone_bd_ram_mem3_reg[70][31]/P0001 ,
		_w11949_,
		_w11986_,
		_w16280_
	);
	LUT4 #(
		.INIT('h0001)
	) name5768 (
		_w16277_,
		_w16278_,
		_w16279_,
		_w16280_,
		_w16281_
	);
	LUT3 #(
		.INIT('h80)
	) name5769 (
		\wishbone_bd_ram_mem3_reg[9][31]/P0001 ,
		_w11932_,
		_w11968_,
		_w16282_
	);
	LUT3 #(
		.INIT('h80)
	) name5770 (
		\wishbone_bd_ram_mem3_reg[217][31]/P0001 ,
		_w11968_,
		_w11984_,
		_w16283_
	);
	LUT3 #(
		.INIT('h80)
	) name5771 (
		\wishbone_bd_ram_mem3_reg[32][31]/P0001 ,
		_w11941_,
		_w11957_,
		_w16284_
	);
	LUT3 #(
		.INIT('h80)
	) name5772 (
		\wishbone_bd_ram_mem3_reg[53][31]/P0001 ,
		_w11933_,
		_w11979_,
		_w16285_
	);
	LUT4 #(
		.INIT('h0001)
	) name5773 (
		_w16282_,
		_w16283_,
		_w16284_,
		_w16285_,
		_w16286_
	);
	LUT3 #(
		.INIT('h80)
	) name5774 (
		\wishbone_bd_ram_mem3_reg[204][31]/P0001 ,
		_w11945_,
		_w11954_,
		_w16287_
	);
	LUT3 #(
		.INIT('h80)
	) name5775 (
		\wishbone_bd_ram_mem3_reg[81][31]/P0001 ,
		_w11972_,
		_w11977_,
		_w16288_
	);
	LUT3 #(
		.INIT('h80)
	) name5776 (
		\wishbone_bd_ram_mem3_reg[159][31]/P0001 ,
		_w11959_,
		_w11973_,
		_w16289_
	);
	LUT3 #(
		.INIT('h80)
	) name5777 (
		\wishbone_bd_ram_mem3_reg[233][31]/P0001 ,
		_w11968_,
		_w11982_,
		_w16290_
	);
	LUT4 #(
		.INIT('h0001)
	) name5778 (
		_w16287_,
		_w16288_,
		_w16289_,
		_w16290_,
		_w16291_
	);
	LUT3 #(
		.INIT('h80)
	) name5779 (
		\wishbone_bd_ram_mem3_reg[205][31]/P0001 ,
		_w11945_,
		_w11966_,
		_w16292_
	);
	LUT3 #(
		.INIT('h80)
	) name5780 (
		\wishbone_bd_ram_mem3_reg[215][31]/P0001 ,
		_w11975_,
		_w11984_,
		_w16293_
	);
	LUT3 #(
		.INIT('h80)
	) name5781 (
		\wishbone_bd_ram_mem3_reg[98][31]/P0001 ,
		_w11963_,
		_w11965_,
		_w16294_
	);
	LUT3 #(
		.INIT('h80)
	) name5782 (
		\wishbone_bd_ram_mem3_reg[49][31]/P0001 ,
		_w11977_,
		_w11979_,
		_w16295_
	);
	LUT4 #(
		.INIT('h0001)
	) name5783 (
		_w16292_,
		_w16293_,
		_w16294_,
		_w16295_,
		_w16296_
	);
	LUT4 #(
		.INIT('h8000)
	) name5784 (
		_w16281_,
		_w16286_,
		_w16291_,
		_w16296_,
		_w16297_
	);
	LUT4 #(
		.INIT('h8000)
	) name5785 (
		_w16234_,
		_w16255_,
		_w16276_,
		_w16297_,
		_w16298_
	);
	LUT3 #(
		.INIT('h80)
	) name5786 (
		\wishbone_bd_ram_mem3_reg[44][31]/P0001 ,
		_w11954_,
		_w11957_,
		_w16299_
	);
	LUT3 #(
		.INIT('h80)
	) name5787 (
		\wishbone_bd_ram_mem3_reg[33][31]/P0001 ,
		_w11957_,
		_w11977_,
		_w16300_
	);
	LUT3 #(
		.INIT('h80)
	) name5788 (
		\wishbone_bd_ram_mem3_reg[167][31]/P0001 ,
		_w11930_,
		_w11975_,
		_w16301_
	);
	LUT3 #(
		.INIT('h80)
	) name5789 (
		\wishbone_bd_ram_mem3_reg[178][31]/P0001 ,
		_w11942_,
		_w11963_,
		_w16302_
	);
	LUT4 #(
		.INIT('h0001)
	) name5790 (
		_w16299_,
		_w16300_,
		_w16301_,
		_w16302_,
		_w16303_
	);
	LUT3 #(
		.INIT('h80)
	) name5791 (
		\wishbone_bd_ram_mem3_reg[61][31]/P0001 ,
		_w11966_,
		_w11979_,
		_w16304_
	);
	LUT3 #(
		.INIT('h80)
	) name5792 (
		\wishbone_bd_ram_mem3_reg[27][31]/P0001 ,
		_w11935_,
		_w11936_,
		_w16305_
	);
	LUT3 #(
		.INIT('h80)
	) name5793 (
		\wishbone_bd_ram_mem3_reg[207][31]/P0001 ,
		_w11945_,
		_w11973_,
		_w16306_
	);
	LUT3 #(
		.INIT('h80)
	) name5794 (
		\wishbone_bd_ram_mem3_reg[116][31]/P0001 ,
		_w11929_,
		_w12012_,
		_w16307_
	);
	LUT4 #(
		.INIT('h0001)
	) name5795 (
		_w16304_,
		_w16305_,
		_w16306_,
		_w16307_,
		_w16308_
	);
	LUT3 #(
		.INIT('h80)
	) name5796 (
		\wishbone_bd_ram_mem3_reg[125][31]/P0001 ,
		_w11966_,
		_w12012_,
		_w16309_
	);
	LUT3 #(
		.INIT('h80)
	) name5797 (
		\wishbone_bd_ram_mem3_reg[40][31]/P0001 ,
		_w11957_,
		_w11990_,
		_w16310_
	);
	LUT3 #(
		.INIT('h80)
	) name5798 (
		\wishbone_bd_ram_mem3_reg[224][31]/P0001 ,
		_w11941_,
		_w11982_,
		_w16311_
	);
	LUT3 #(
		.INIT('h80)
	) name5799 (
		\wishbone_bd_ram_mem3_reg[101][31]/P0001 ,
		_w11933_,
		_w11965_,
		_w16312_
	);
	LUT4 #(
		.INIT('h0001)
	) name5800 (
		_w16309_,
		_w16310_,
		_w16311_,
		_w16312_,
		_w16313_
	);
	LUT3 #(
		.INIT('h80)
	) name5801 (
		\wishbone_bd_ram_mem3_reg[56][31]/P0001 ,
		_w11979_,
		_w11990_,
		_w16314_
	);
	LUT3 #(
		.INIT('h80)
	) name5802 (
		\wishbone_bd_ram_mem3_reg[120][31]/P0001 ,
		_w11990_,
		_w12012_,
		_w16315_
	);
	LUT3 #(
		.INIT('h80)
	) name5803 (
		\wishbone_bd_ram_mem3_reg[112][31]/P0001 ,
		_w11941_,
		_w12012_,
		_w16316_
	);
	LUT3 #(
		.INIT('h80)
	) name5804 (
		\wishbone_bd_ram_mem3_reg[19][31]/P0001 ,
		_w11935_,
		_w11938_,
		_w16317_
	);
	LUT4 #(
		.INIT('h0001)
	) name5805 (
		_w16314_,
		_w16315_,
		_w16316_,
		_w16317_,
		_w16318_
	);
	LUT4 #(
		.INIT('h8000)
	) name5806 (
		_w16303_,
		_w16308_,
		_w16313_,
		_w16318_,
		_w16319_
	);
	LUT3 #(
		.INIT('h80)
	) name5807 (
		\wishbone_bd_ram_mem3_reg[229][31]/P0001 ,
		_w11933_,
		_w11982_,
		_w16320_
	);
	LUT3 #(
		.INIT('h80)
	) name5808 (
		\wishbone_bd_ram_mem3_reg[12][31]/P0001 ,
		_w11932_,
		_w11954_,
		_w16321_
	);
	LUT3 #(
		.INIT('h80)
	) name5809 (
		\wishbone_bd_ram_mem3_reg[21][31]/P0001 ,
		_w11933_,
		_w11935_,
		_w16322_
	);
	LUT3 #(
		.INIT('h80)
	) name5810 (
		\wishbone_bd_ram_mem3_reg[166][31]/P0001 ,
		_w11930_,
		_w11986_,
		_w16323_
	);
	LUT4 #(
		.INIT('h0001)
	) name5811 (
		_w16320_,
		_w16321_,
		_w16322_,
		_w16323_,
		_w16324_
	);
	LUT3 #(
		.INIT('h80)
	) name5812 (
		\wishbone_bd_ram_mem3_reg[219][31]/P0001 ,
		_w11936_,
		_w11984_,
		_w16325_
	);
	LUT3 #(
		.INIT('h80)
	) name5813 (
		\wishbone_bd_ram_mem3_reg[169][31]/P0001 ,
		_w11930_,
		_w11968_,
		_w16326_
	);
	LUT3 #(
		.INIT('h80)
	) name5814 (
		\wishbone_bd_ram_mem3_reg[91][31]/P0001 ,
		_w11936_,
		_w11972_,
		_w16327_
	);
	LUT3 #(
		.INIT('h80)
	) name5815 (
		\wishbone_bd_ram_mem3_reg[222][31]/P0001 ,
		_w11948_,
		_w11984_,
		_w16328_
	);
	LUT4 #(
		.INIT('h0001)
	) name5816 (
		_w16325_,
		_w16326_,
		_w16327_,
		_w16328_,
		_w16329_
	);
	LUT3 #(
		.INIT('h80)
	) name5817 (
		\wishbone_bd_ram_mem3_reg[77][31]/P0001 ,
		_w11949_,
		_w11966_,
		_w16330_
	);
	LUT3 #(
		.INIT('h80)
	) name5818 (
		\wishbone_bd_ram_mem3_reg[24][31]/P0001 ,
		_w11935_,
		_w11990_,
		_w16331_
	);
	LUT3 #(
		.INIT('h80)
	) name5819 (
		\wishbone_bd_ram_mem3_reg[74][31]/P0001 ,
		_w11944_,
		_w11949_,
		_w16332_
	);
	LUT3 #(
		.INIT('h80)
	) name5820 (
		\wishbone_bd_ram_mem3_reg[76][31]/P0001 ,
		_w11949_,
		_w11954_,
		_w16333_
	);
	LUT4 #(
		.INIT('h0001)
	) name5821 (
		_w16330_,
		_w16331_,
		_w16332_,
		_w16333_,
		_w16334_
	);
	LUT3 #(
		.INIT('h80)
	) name5822 (
		\wishbone_bd_ram_mem3_reg[22][31]/P0001 ,
		_w11935_,
		_w11986_,
		_w16335_
	);
	LUT3 #(
		.INIT('h80)
	) name5823 (
		\wishbone_bd_ram_mem3_reg[6][31]/P0001 ,
		_w11932_,
		_w11986_,
		_w16336_
	);
	LUT3 #(
		.INIT('h80)
	) name5824 (
		\wishbone_bd_ram_mem3_reg[35][31]/P0001 ,
		_w11938_,
		_w11957_,
		_w16337_
	);
	LUT3 #(
		.INIT('h80)
	) name5825 (
		\wishbone_bd_ram_mem3_reg[165][31]/P0001 ,
		_w11930_,
		_w11933_,
		_w16338_
	);
	LUT4 #(
		.INIT('h0001)
	) name5826 (
		_w16335_,
		_w16336_,
		_w16337_,
		_w16338_,
		_w16339_
	);
	LUT4 #(
		.INIT('h8000)
	) name5827 (
		_w16324_,
		_w16329_,
		_w16334_,
		_w16339_,
		_w16340_
	);
	LUT3 #(
		.INIT('h80)
	) name5828 (
		\wishbone_bd_ram_mem3_reg[251][31]/P0001 ,
		_w11936_,
		_w11952_,
		_w16341_
	);
	LUT3 #(
		.INIT('h80)
	) name5829 (
		\wishbone_bd_ram_mem3_reg[73][31]/P0001 ,
		_w11949_,
		_w11968_,
		_w16342_
	);
	LUT3 #(
		.INIT('h80)
	) name5830 (
		\wishbone_bd_ram_mem3_reg[2][31]/P0001 ,
		_w11932_,
		_w11963_,
		_w16343_
	);
	LUT3 #(
		.INIT('h80)
	) name5831 (
		\wishbone_bd_ram_mem3_reg[236][31]/P0001 ,
		_w11954_,
		_w11982_,
		_w16344_
	);
	LUT4 #(
		.INIT('h0001)
	) name5832 (
		_w16341_,
		_w16342_,
		_w16343_,
		_w16344_,
		_w16345_
	);
	LUT3 #(
		.INIT('h80)
	) name5833 (
		\wishbone_bd_ram_mem3_reg[249][31]/P0001 ,
		_w11952_,
		_w11968_,
		_w16346_
	);
	LUT3 #(
		.INIT('h80)
	) name5834 (
		\wishbone_bd_ram_mem3_reg[177][31]/P0001 ,
		_w11942_,
		_w11977_,
		_w16347_
	);
	LUT3 #(
		.INIT('h80)
	) name5835 (
		\wishbone_bd_ram_mem3_reg[92][31]/P0001 ,
		_w11954_,
		_w11972_,
		_w16348_
	);
	LUT3 #(
		.INIT('h80)
	) name5836 (
		\wishbone_bd_ram_mem3_reg[83][31]/P0001 ,
		_w11938_,
		_w11972_,
		_w16349_
	);
	LUT4 #(
		.INIT('h0001)
	) name5837 (
		_w16346_,
		_w16347_,
		_w16348_,
		_w16349_,
		_w16350_
	);
	LUT3 #(
		.INIT('h80)
	) name5838 (
		\wishbone_bd_ram_mem3_reg[18][31]/P0001 ,
		_w11935_,
		_w11963_,
		_w16351_
	);
	LUT3 #(
		.INIT('h80)
	) name5839 (
		\wishbone_bd_ram_mem3_reg[110][31]/P0001 ,
		_w11948_,
		_w11965_,
		_w16352_
	);
	LUT3 #(
		.INIT('h80)
	) name5840 (
		\wishbone_bd_ram_mem3_reg[148][31]/P0001 ,
		_w11929_,
		_w11959_,
		_w16353_
	);
	LUT3 #(
		.INIT('h80)
	) name5841 (
		\wishbone_bd_ram_mem3_reg[175][31]/P0001 ,
		_w11930_,
		_w11973_,
		_w16354_
	);
	LUT4 #(
		.INIT('h0001)
	) name5842 (
		_w16351_,
		_w16352_,
		_w16353_,
		_w16354_,
		_w16355_
	);
	LUT3 #(
		.INIT('h80)
	) name5843 (
		\wishbone_bd_ram_mem3_reg[131][31]/P0001 ,
		_w11938_,
		_w11955_,
		_w16356_
	);
	LUT3 #(
		.INIT('h80)
	) name5844 (
		\wishbone_bd_ram_mem3_reg[100][31]/P0001 ,
		_w11929_,
		_w11965_,
		_w16357_
	);
	LUT3 #(
		.INIT('h80)
	) name5845 (
		\wishbone_bd_ram_mem3_reg[152][31]/P0001 ,
		_w11959_,
		_w11990_,
		_w16358_
	);
	LUT3 #(
		.INIT('h80)
	) name5846 (
		\wishbone_bd_ram_mem3_reg[163][31]/P0001 ,
		_w11930_,
		_w11938_,
		_w16359_
	);
	LUT4 #(
		.INIT('h0001)
	) name5847 (
		_w16356_,
		_w16357_,
		_w16358_,
		_w16359_,
		_w16360_
	);
	LUT4 #(
		.INIT('h8000)
	) name5848 (
		_w16345_,
		_w16350_,
		_w16355_,
		_w16360_,
		_w16361_
	);
	LUT3 #(
		.INIT('h80)
	) name5849 (
		\wishbone_bd_ram_mem3_reg[199][31]/P0001 ,
		_w11945_,
		_w11975_,
		_w16362_
	);
	LUT3 #(
		.INIT('h80)
	) name5850 (
		\wishbone_bd_ram_mem3_reg[114][31]/P0001 ,
		_w11963_,
		_w12012_,
		_w16363_
	);
	LUT3 #(
		.INIT('h80)
	) name5851 (
		\wishbone_bd_ram_mem3_reg[138][31]/P0001 ,
		_w11944_,
		_w11955_,
		_w16364_
	);
	LUT3 #(
		.INIT('h80)
	) name5852 (
		\wishbone_bd_ram_mem3_reg[10][31]/P0001 ,
		_w11932_,
		_w11944_,
		_w16365_
	);
	LUT4 #(
		.INIT('h0001)
	) name5853 (
		_w16362_,
		_w16363_,
		_w16364_,
		_w16365_,
		_w16366_
	);
	LUT3 #(
		.INIT('h80)
	) name5854 (
		\wishbone_bd_ram_mem3_reg[90][31]/P0001 ,
		_w11944_,
		_w11972_,
		_w16367_
	);
	LUT3 #(
		.INIT('h80)
	) name5855 (
		\wishbone_bd_ram_mem3_reg[140][31]/P0001 ,
		_w11954_,
		_w11955_,
		_w16368_
	);
	LUT3 #(
		.INIT('h80)
	) name5856 (
		\wishbone_bd_ram_mem3_reg[253][31]/P0001 ,
		_w11952_,
		_w11966_,
		_w16369_
	);
	LUT3 #(
		.INIT('h80)
	) name5857 (
		\wishbone_bd_ram_mem3_reg[223][31]/P0001 ,
		_w11973_,
		_w11984_,
		_w16370_
	);
	LUT4 #(
		.INIT('h0001)
	) name5858 (
		_w16367_,
		_w16368_,
		_w16369_,
		_w16370_,
		_w16371_
	);
	LUT3 #(
		.INIT('h80)
	) name5859 (
		\wishbone_bd_ram_mem3_reg[246][31]/P0001 ,
		_w11952_,
		_w11986_,
		_w16372_
	);
	LUT3 #(
		.INIT('h80)
	) name5860 (
		\wishbone_bd_ram_mem3_reg[80][31]/P0001 ,
		_w11941_,
		_w11972_,
		_w16373_
	);
	LUT3 #(
		.INIT('h80)
	) name5861 (
		\wishbone_bd_ram_mem3_reg[147][31]/P0001 ,
		_w11938_,
		_w11959_,
		_w16374_
	);
	LUT3 #(
		.INIT('h80)
	) name5862 (
		\wishbone_bd_ram_mem3_reg[237][31]/P0001 ,
		_w11966_,
		_w11982_,
		_w16375_
	);
	LUT4 #(
		.INIT('h0001)
	) name5863 (
		_w16372_,
		_w16373_,
		_w16374_,
		_w16375_,
		_w16376_
	);
	LUT3 #(
		.INIT('h80)
	) name5864 (
		\wishbone_bd_ram_mem3_reg[75][31]/P0001 ,
		_w11936_,
		_w11949_,
		_w16377_
	);
	LUT3 #(
		.INIT('h80)
	) name5865 (
		\wishbone_bd_ram_mem3_reg[164][31]/P0001 ,
		_w11929_,
		_w11930_,
		_w16378_
	);
	LUT3 #(
		.INIT('h80)
	) name5866 (
		\wishbone_bd_ram_mem3_reg[50][31]/P0001 ,
		_w11963_,
		_w11979_,
		_w16379_
	);
	LUT3 #(
		.INIT('h80)
	) name5867 (
		\wishbone_bd_ram_mem3_reg[1][31]/P0001 ,
		_w11932_,
		_w11977_,
		_w16380_
	);
	LUT4 #(
		.INIT('h0001)
	) name5868 (
		_w16377_,
		_w16378_,
		_w16379_,
		_w16380_,
		_w16381_
	);
	LUT4 #(
		.INIT('h8000)
	) name5869 (
		_w16366_,
		_w16371_,
		_w16376_,
		_w16381_,
		_w16382_
	);
	LUT4 #(
		.INIT('h8000)
	) name5870 (
		_w16319_,
		_w16340_,
		_w16361_,
		_w16382_,
		_w16383_
	);
	LUT3 #(
		.INIT('h80)
	) name5871 (
		\wishbone_bd_ram_mem3_reg[64][31]/P0001 ,
		_w11941_,
		_w11949_,
		_w16384_
	);
	LUT3 #(
		.INIT('h80)
	) name5872 (
		\wishbone_bd_ram_mem3_reg[196][31]/P0001 ,
		_w11929_,
		_w11945_,
		_w16385_
	);
	LUT3 #(
		.INIT('h80)
	) name5873 (
		\wishbone_bd_ram_mem3_reg[59][31]/P0001 ,
		_w11936_,
		_w11979_,
		_w16386_
	);
	LUT3 #(
		.INIT('h80)
	) name5874 (
		\wishbone_bd_ram_mem3_reg[123][31]/P0001 ,
		_w11936_,
		_w12012_,
		_w16387_
	);
	LUT4 #(
		.INIT('h0001)
	) name5875 (
		_w16384_,
		_w16385_,
		_w16386_,
		_w16387_,
		_w16388_
	);
	LUT3 #(
		.INIT('h80)
	) name5876 (
		\wishbone_bd_ram_mem3_reg[108][31]/P0001 ,
		_w11954_,
		_w11965_,
		_w16389_
	);
	LUT3 #(
		.INIT('h80)
	) name5877 (
		\wishbone_bd_ram_mem3_reg[137][31]/P0001 ,
		_w11955_,
		_w11968_,
		_w16390_
	);
	LUT3 #(
		.INIT('h80)
	) name5878 (
		\wishbone_bd_ram_mem3_reg[62][31]/P0001 ,
		_w11948_,
		_w11979_,
		_w16391_
	);
	LUT3 #(
		.INIT('h80)
	) name5879 (
		\wishbone_bd_ram_mem3_reg[206][31]/P0001 ,
		_w11945_,
		_w11948_,
		_w16392_
	);
	LUT4 #(
		.INIT('h0001)
	) name5880 (
		_w16389_,
		_w16390_,
		_w16391_,
		_w16392_,
		_w16393_
	);
	LUT3 #(
		.INIT('h80)
	) name5881 (
		\wishbone_bd_ram_mem3_reg[117][31]/P0001 ,
		_w11933_,
		_w12012_,
		_w16394_
	);
	LUT3 #(
		.INIT('h80)
	) name5882 (
		\wishbone_bd_ram_mem3_reg[181][31]/P0001 ,
		_w11933_,
		_w11942_,
		_w16395_
	);
	LUT3 #(
		.INIT('h80)
	) name5883 (
		\wishbone_bd_ram_mem3_reg[46][31]/P0001 ,
		_w11948_,
		_w11957_,
		_w16396_
	);
	LUT3 #(
		.INIT('h80)
	) name5884 (
		\wishbone_bd_ram_mem3_reg[201][31]/P0001 ,
		_w11945_,
		_w11968_,
		_w16397_
	);
	LUT4 #(
		.INIT('h0001)
	) name5885 (
		_w16394_,
		_w16395_,
		_w16396_,
		_w16397_,
		_w16398_
	);
	LUT3 #(
		.INIT('h80)
	) name5886 (
		\wishbone_bd_ram_mem3_reg[31][31]/P0001 ,
		_w11935_,
		_w11973_,
		_w16399_
	);
	LUT3 #(
		.INIT('h80)
	) name5887 (
		\wishbone_bd_ram_mem3_reg[16][31]/P0001 ,
		_w11935_,
		_w11941_,
		_w16400_
	);
	LUT3 #(
		.INIT('h80)
	) name5888 (
		\wishbone_bd_ram_mem3_reg[54][31]/P0001 ,
		_w11979_,
		_w11986_,
		_w16401_
	);
	LUT3 #(
		.INIT('h80)
	) name5889 (
		\wishbone_bd_ram_mem3_reg[86][31]/P0001 ,
		_w11972_,
		_w11986_,
		_w16402_
	);
	LUT4 #(
		.INIT('h0001)
	) name5890 (
		_w16399_,
		_w16400_,
		_w16401_,
		_w16402_,
		_w16403_
	);
	LUT4 #(
		.INIT('h8000)
	) name5891 (
		_w16388_,
		_w16393_,
		_w16398_,
		_w16403_,
		_w16404_
	);
	LUT3 #(
		.INIT('h80)
	) name5892 (
		\wishbone_bd_ram_mem3_reg[156][31]/P0001 ,
		_w11954_,
		_w11959_,
		_w16405_
	);
	LUT3 #(
		.INIT('h80)
	) name5893 (
		\wishbone_bd_ram_mem3_reg[36][31]/P0001 ,
		_w11929_,
		_w11957_,
		_w16406_
	);
	LUT3 #(
		.INIT('h80)
	) name5894 (
		\wishbone_bd_ram_mem3_reg[78][31]/P0001 ,
		_w11948_,
		_w11949_,
		_w16407_
	);
	LUT3 #(
		.INIT('h80)
	) name5895 (
		\wishbone_bd_ram_mem3_reg[231][31]/P0001 ,
		_w11975_,
		_w11982_,
		_w16408_
	);
	LUT4 #(
		.INIT('h0001)
	) name5896 (
		_w16405_,
		_w16406_,
		_w16407_,
		_w16408_,
		_w16409_
	);
	LUT3 #(
		.INIT('h80)
	) name5897 (
		\wishbone_bd_ram_mem3_reg[153][31]/P0001 ,
		_w11959_,
		_w11968_,
		_w16410_
	);
	LUT3 #(
		.INIT('h80)
	) name5898 (
		\wishbone_bd_ram_mem3_reg[134][31]/P0001 ,
		_w11955_,
		_w11986_,
		_w16411_
	);
	LUT3 #(
		.INIT('h80)
	) name5899 (
		\wishbone_bd_ram_mem3_reg[23][31]/P0001 ,
		_w11935_,
		_w11975_,
		_w16412_
	);
	LUT3 #(
		.INIT('h80)
	) name5900 (
		\wishbone_bd_ram_mem3_reg[11][31]/P0001 ,
		_w11932_,
		_w11936_,
		_w16413_
	);
	LUT4 #(
		.INIT('h0001)
	) name5901 (
		_w16410_,
		_w16411_,
		_w16412_,
		_w16413_,
		_w16414_
	);
	LUT3 #(
		.INIT('h80)
	) name5902 (
		\wishbone_bd_ram_mem3_reg[243][31]/P0001 ,
		_w11938_,
		_w11952_,
		_w16415_
	);
	LUT3 #(
		.INIT('h80)
	) name5903 (
		\wishbone_bd_ram_mem3_reg[158][31]/P0001 ,
		_w11948_,
		_w11959_,
		_w16416_
	);
	LUT3 #(
		.INIT('h80)
	) name5904 (
		\wishbone_bd_ram_mem3_reg[162][31]/P0001 ,
		_w11930_,
		_w11963_,
		_w16417_
	);
	LUT3 #(
		.INIT('h80)
	) name5905 (
		\wishbone_bd_ram_mem3_reg[26][31]/P0001 ,
		_w11935_,
		_w11944_,
		_w16418_
	);
	LUT4 #(
		.INIT('h0001)
	) name5906 (
		_w16415_,
		_w16416_,
		_w16417_,
		_w16418_,
		_w16419_
	);
	LUT3 #(
		.INIT('h80)
	) name5907 (
		\wishbone_bd_ram_mem3_reg[142][31]/P0001 ,
		_w11948_,
		_w11955_,
		_w16420_
	);
	LUT3 #(
		.INIT('h80)
	) name5908 (
		\wishbone_bd_ram_mem3_reg[20][31]/P0001 ,
		_w11929_,
		_w11935_,
		_w16421_
	);
	LUT3 #(
		.INIT('h80)
	) name5909 (
		\wishbone_bd_ram_mem3_reg[194][31]/P0001 ,
		_w11945_,
		_w11963_,
		_w16422_
	);
	LUT3 #(
		.INIT('h80)
	) name5910 (
		\wishbone_bd_ram_mem3_reg[63][31]/P0001 ,
		_w11973_,
		_w11979_,
		_w16423_
	);
	LUT4 #(
		.INIT('h0001)
	) name5911 (
		_w16420_,
		_w16421_,
		_w16422_,
		_w16423_,
		_w16424_
	);
	LUT4 #(
		.INIT('h8000)
	) name5912 (
		_w16409_,
		_w16414_,
		_w16419_,
		_w16424_,
		_w16425_
	);
	LUT3 #(
		.INIT('h80)
	) name5913 (
		\wishbone_bd_ram_mem3_reg[212][31]/P0001 ,
		_w11929_,
		_w11984_,
		_w16426_
	);
	LUT3 #(
		.INIT('h80)
	) name5914 (
		\wishbone_bd_ram_mem3_reg[5][31]/P0001 ,
		_w11932_,
		_w11933_,
		_w16427_
	);
	LUT3 #(
		.INIT('h80)
	) name5915 (
		\wishbone_bd_ram_mem3_reg[106][31]/P0001 ,
		_w11944_,
		_w11965_,
		_w16428_
	);
	LUT3 #(
		.INIT('h80)
	) name5916 (
		\wishbone_bd_ram_mem3_reg[154][31]/P0001 ,
		_w11944_,
		_w11959_,
		_w16429_
	);
	LUT4 #(
		.INIT('h0001)
	) name5917 (
		_w16426_,
		_w16427_,
		_w16428_,
		_w16429_,
		_w16430_
	);
	LUT3 #(
		.INIT('h80)
	) name5918 (
		\wishbone_bd_ram_mem3_reg[95][31]/P0001 ,
		_w11972_,
		_w11973_,
		_w16431_
	);
	LUT3 #(
		.INIT('h80)
	) name5919 (
		\wishbone_bd_ram_mem3_reg[195][31]/P0001 ,
		_w11938_,
		_w11945_,
		_w16432_
	);
	LUT3 #(
		.INIT('h80)
	) name5920 (
		\wishbone_bd_ram_mem3_reg[99][31]/P0001 ,
		_w11938_,
		_w11965_,
		_w16433_
	);
	LUT3 #(
		.INIT('h80)
	) name5921 (
		\wishbone_bd_ram_mem3_reg[211][31]/P0001 ,
		_w11938_,
		_w11984_,
		_w16434_
	);
	LUT4 #(
		.INIT('h0001)
	) name5922 (
		_w16431_,
		_w16432_,
		_w16433_,
		_w16434_,
		_w16435_
	);
	LUT3 #(
		.INIT('h80)
	) name5923 (
		\wishbone_bd_ram_mem3_reg[65][31]/P0001 ,
		_w11949_,
		_w11977_,
		_w16436_
	);
	LUT3 #(
		.INIT('h80)
	) name5924 (
		\wishbone_bd_ram_mem3_reg[115][31]/P0001 ,
		_w11938_,
		_w12012_,
		_w16437_
	);
	LUT3 #(
		.INIT('h80)
	) name5925 (
		\wishbone_bd_ram_mem3_reg[79][31]/P0001 ,
		_w11949_,
		_w11973_,
		_w16438_
	);
	LUT3 #(
		.INIT('h80)
	) name5926 (
		\wishbone_bd_ram_mem3_reg[124][31]/P0001 ,
		_w11954_,
		_w12012_,
		_w16439_
	);
	LUT4 #(
		.INIT('h0001)
	) name5927 (
		_w16436_,
		_w16437_,
		_w16438_,
		_w16439_,
		_w16440_
	);
	LUT3 #(
		.INIT('h80)
	) name5928 (
		\wishbone_bd_ram_mem3_reg[213][31]/P0001 ,
		_w11933_,
		_w11984_,
		_w16441_
	);
	LUT3 #(
		.INIT('h80)
	) name5929 (
		\wishbone_bd_ram_mem3_reg[96][31]/P0001 ,
		_w11941_,
		_w11965_,
		_w16442_
	);
	LUT3 #(
		.INIT('h80)
	) name5930 (
		\wishbone_bd_ram_mem3_reg[214][31]/P0001 ,
		_w11984_,
		_w11986_,
		_w16443_
	);
	LUT3 #(
		.INIT('h80)
	) name5931 (
		\wishbone_bd_ram_mem3_reg[4][31]/P0001 ,
		_w11929_,
		_w11932_,
		_w16444_
	);
	LUT4 #(
		.INIT('h0001)
	) name5932 (
		_w16441_,
		_w16442_,
		_w16443_,
		_w16444_,
		_w16445_
	);
	LUT4 #(
		.INIT('h8000)
	) name5933 (
		_w16430_,
		_w16435_,
		_w16440_,
		_w16445_,
		_w16446_
	);
	LUT3 #(
		.INIT('h80)
	) name5934 (
		\wishbone_bd_ram_mem3_reg[151][31]/P0001 ,
		_w11959_,
		_w11975_,
		_w16447_
	);
	LUT3 #(
		.INIT('h80)
	) name5935 (
		\wishbone_bd_ram_mem3_reg[208][31]/P0001 ,
		_w11941_,
		_w11984_,
		_w16448_
	);
	LUT3 #(
		.INIT('h80)
	) name5936 (
		\wishbone_bd_ram_mem3_reg[130][31]/P0001 ,
		_w11955_,
		_w11963_,
		_w16449_
	);
	LUT3 #(
		.INIT('h80)
	) name5937 (
		\wishbone_bd_ram_mem3_reg[102][31]/P0001 ,
		_w11965_,
		_w11986_,
		_w16450_
	);
	LUT4 #(
		.INIT('h0001)
	) name5938 (
		_w16447_,
		_w16448_,
		_w16449_,
		_w16450_,
		_w16451_
	);
	LUT3 #(
		.INIT('h80)
	) name5939 (
		\wishbone_bd_ram_mem3_reg[225][31]/P0001 ,
		_w11977_,
		_w11982_,
		_w16452_
	);
	LUT3 #(
		.INIT('h80)
	) name5940 (
		\wishbone_bd_ram_mem3_reg[255][31]/P0001 ,
		_w11952_,
		_w11973_,
		_w16453_
	);
	LUT3 #(
		.INIT('h80)
	) name5941 (
		\wishbone_bd_ram_mem3_reg[122][31]/P0001 ,
		_w11944_,
		_w12012_,
		_w16454_
	);
	LUT3 #(
		.INIT('h80)
	) name5942 (
		\wishbone_bd_ram_mem3_reg[126][31]/P0001 ,
		_w11948_,
		_w12012_,
		_w16455_
	);
	LUT4 #(
		.INIT('h0001)
	) name5943 (
		_w16452_,
		_w16453_,
		_w16454_,
		_w16455_,
		_w16456_
	);
	LUT3 #(
		.INIT('h80)
	) name5944 (
		\wishbone_bd_ram_mem3_reg[141][31]/P0001 ,
		_w11955_,
		_w11966_,
		_w16457_
	);
	LUT3 #(
		.INIT('h80)
	) name5945 (
		\wishbone_bd_ram_mem3_reg[250][31]/P0001 ,
		_w11944_,
		_w11952_,
		_w16458_
	);
	LUT3 #(
		.INIT('h80)
	) name5946 (
		\wishbone_bd_ram_mem3_reg[176][31]/P0001 ,
		_w11941_,
		_w11942_,
		_w16459_
	);
	LUT3 #(
		.INIT('h80)
	) name5947 (
		\wishbone_bd_ram_mem3_reg[198][31]/P0001 ,
		_w11945_,
		_w11986_,
		_w16460_
	);
	LUT4 #(
		.INIT('h0001)
	) name5948 (
		_w16457_,
		_w16458_,
		_w16459_,
		_w16460_,
		_w16461_
	);
	LUT3 #(
		.INIT('h80)
	) name5949 (
		\wishbone_bd_ram_mem3_reg[129][31]/P0001 ,
		_w11955_,
		_w11977_,
		_w16462_
	);
	LUT3 #(
		.INIT('h80)
	) name5950 (
		\wishbone_bd_ram_mem3_reg[146][31]/P0001 ,
		_w11959_,
		_w11963_,
		_w16463_
	);
	LUT3 #(
		.INIT('h80)
	) name5951 (
		\wishbone_bd_ram_mem3_reg[8][31]/P0001 ,
		_w11932_,
		_w11990_,
		_w16464_
	);
	LUT3 #(
		.INIT('h80)
	) name5952 (
		\wishbone_bd_ram_mem3_reg[209][31]/P0001 ,
		_w11977_,
		_w11984_,
		_w16465_
	);
	LUT4 #(
		.INIT('h0001)
	) name5953 (
		_w16462_,
		_w16463_,
		_w16464_,
		_w16465_,
		_w16466_
	);
	LUT4 #(
		.INIT('h8000)
	) name5954 (
		_w16451_,
		_w16456_,
		_w16461_,
		_w16466_,
		_w16467_
	);
	LUT4 #(
		.INIT('h8000)
	) name5955 (
		_w16404_,
		_w16425_,
		_w16446_,
		_w16467_,
		_w16468_
	);
	LUT4 #(
		.INIT('h8000)
	) name5956 (
		_w16213_,
		_w16298_,
		_w16383_,
		_w16468_,
		_w16469_
	);
	LUT4 #(
		.INIT('h007f)
	) name5957 (
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		\wishbone_TxLength_reg[15]/NET0131 ,
		_w16470_
	);
	LUT3 #(
		.INIT('h40)
	) name5958 (
		_w12302_,
		_w12314_,
		_w12315_,
		_w16471_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name5959 (
		_w12312_,
		_w14878_,
		_w16470_,
		_w16471_,
		_w16472_
	);
	LUT4 #(
		.INIT('h3700)
	) name5960 (
		wb_rst_i_pad,
		_w12302_,
		_w16469_,
		_w16472_,
		_w16473_
	);
	LUT3 #(
		.INIT('h80)
	) name5961 (
		\wishbone_bd_ram_mem2_reg[173][17]/P0001 ,
		_w11930_,
		_w11966_,
		_w16474_
	);
	LUT3 #(
		.INIT('h80)
	) name5962 (
		\wishbone_bd_ram_mem2_reg[105][17]/P0001 ,
		_w11965_,
		_w11968_,
		_w16475_
	);
	LUT3 #(
		.INIT('h80)
	) name5963 (
		\wishbone_bd_ram_mem2_reg[212][17]/P0001 ,
		_w11929_,
		_w11984_,
		_w16476_
	);
	LUT3 #(
		.INIT('h80)
	) name5964 (
		\wishbone_bd_ram_mem2_reg[209][17]/P0001 ,
		_w11977_,
		_w11984_,
		_w16477_
	);
	LUT4 #(
		.INIT('h0001)
	) name5965 (
		_w16474_,
		_w16475_,
		_w16476_,
		_w16477_,
		_w16478_
	);
	LUT3 #(
		.INIT('h80)
	) name5966 (
		\wishbone_bd_ram_mem2_reg[13][17]/P0001 ,
		_w11932_,
		_w11966_,
		_w16479_
	);
	LUT3 #(
		.INIT('h80)
	) name5967 (
		\wishbone_bd_ram_mem2_reg[12][17]/P0001 ,
		_w11932_,
		_w11954_,
		_w16480_
	);
	LUT3 #(
		.INIT('h80)
	) name5968 (
		\wishbone_bd_ram_mem2_reg[51][17]/P0001 ,
		_w11938_,
		_w11979_,
		_w16481_
	);
	LUT3 #(
		.INIT('h80)
	) name5969 (
		\wishbone_bd_ram_mem2_reg[183][17]/P0001 ,
		_w11942_,
		_w11975_,
		_w16482_
	);
	LUT4 #(
		.INIT('h0001)
	) name5970 (
		_w16479_,
		_w16480_,
		_w16481_,
		_w16482_,
		_w16483_
	);
	LUT3 #(
		.INIT('h80)
	) name5971 (
		\wishbone_bd_ram_mem2_reg[161][17]/P0001 ,
		_w11930_,
		_w11977_,
		_w16484_
	);
	LUT3 #(
		.INIT('h80)
	) name5972 (
		\wishbone_bd_ram_mem2_reg[33][17]/P0001 ,
		_w11957_,
		_w11977_,
		_w16485_
	);
	LUT3 #(
		.INIT('h80)
	) name5973 (
		\wishbone_bd_ram_mem2_reg[76][17]/P0001 ,
		_w11949_,
		_w11954_,
		_w16486_
	);
	LUT3 #(
		.INIT('h80)
	) name5974 (
		\wishbone_bd_ram_mem2_reg[57][17]/P0001 ,
		_w11968_,
		_w11979_,
		_w16487_
	);
	LUT4 #(
		.INIT('h0001)
	) name5975 (
		_w16484_,
		_w16485_,
		_w16486_,
		_w16487_,
		_w16488_
	);
	LUT3 #(
		.INIT('h80)
	) name5976 (
		\wishbone_bd_ram_mem2_reg[213][17]/P0001 ,
		_w11933_,
		_w11984_,
		_w16489_
	);
	LUT3 #(
		.INIT('h80)
	) name5977 (
		\wishbone_bd_ram_mem2_reg[166][17]/P0001 ,
		_w11930_,
		_w11986_,
		_w16490_
	);
	LUT3 #(
		.INIT('h80)
	) name5978 (
		\wishbone_bd_ram_mem2_reg[117][17]/P0001 ,
		_w11933_,
		_w12012_,
		_w16491_
	);
	LUT3 #(
		.INIT('h80)
	) name5979 (
		\wishbone_bd_ram_mem2_reg[23][17]/P0001 ,
		_w11935_,
		_w11975_,
		_w16492_
	);
	LUT4 #(
		.INIT('h0001)
	) name5980 (
		_w16489_,
		_w16490_,
		_w16491_,
		_w16492_,
		_w16493_
	);
	LUT4 #(
		.INIT('h8000)
	) name5981 (
		_w16478_,
		_w16483_,
		_w16488_,
		_w16493_,
		_w16494_
	);
	LUT3 #(
		.INIT('h80)
	) name5982 (
		\wishbone_bd_ram_mem2_reg[143][17]/P0001 ,
		_w11955_,
		_w11973_,
		_w16495_
	);
	LUT3 #(
		.INIT('h80)
	) name5983 (
		\wishbone_bd_ram_mem2_reg[102][17]/P0001 ,
		_w11965_,
		_w11986_,
		_w16496_
	);
	LUT3 #(
		.INIT('h80)
	) name5984 (
		\wishbone_bd_ram_mem2_reg[90][17]/P0001 ,
		_w11944_,
		_w11972_,
		_w16497_
	);
	LUT3 #(
		.INIT('h80)
	) name5985 (
		\wishbone_bd_ram_mem2_reg[176][17]/P0001 ,
		_w11941_,
		_w11942_,
		_w16498_
	);
	LUT4 #(
		.INIT('h0001)
	) name5986 (
		_w16495_,
		_w16496_,
		_w16497_,
		_w16498_,
		_w16499_
	);
	LUT3 #(
		.INIT('h80)
	) name5987 (
		\wishbone_bd_ram_mem2_reg[22][17]/P0001 ,
		_w11935_,
		_w11986_,
		_w16500_
	);
	LUT3 #(
		.INIT('h80)
	) name5988 (
		\wishbone_bd_ram_mem2_reg[84][17]/P0001 ,
		_w11929_,
		_w11972_,
		_w16501_
	);
	LUT3 #(
		.INIT('h80)
	) name5989 (
		\wishbone_bd_ram_mem2_reg[60][17]/P0001 ,
		_w11954_,
		_w11979_,
		_w16502_
	);
	LUT3 #(
		.INIT('h80)
	) name5990 (
		\wishbone_bd_ram_mem2_reg[10][17]/P0001 ,
		_w11932_,
		_w11944_,
		_w16503_
	);
	LUT4 #(
		.INIT('h0001)
	) name5991 (
		_w16500_,
		_w16501_,
		_w16502_,
		_w16503_,
		_w16504_
	);
	LUT3 #(
		.INIT('h80)
	) name5992 (
		\wishbone_bd_ram_mem2_reg[9][17]/P0001 ,
		_w11932_,
		_w11968_,
		_w16505_
	);
	LUT3 #(
		.INIT('h80)
	) name5993 (
		\wishbone_bd_ram_mem2_reg[234][17]/P0001 ,
		_w11944_,
		_w11982_,
		_w16506_
	);
	LUT3 #(
		.INIT('h80)
	) name5994 (
		\wishbone_bd_ram_mem2_reg[168][17]/P0001 ,
		_w11930_,
		_w11990_,
		_w16507_
	);
	LUT3 #(
		.INIT('h80)
	) name5995 (
		\wishbone_bd_ram_mem2_reg[231][17]/P0001 ,
		_w11975_,
		_w11982_,
		_w16508_
	);
	LUT4 #(
		.INIT('h0001)
	) name5996 (
		_w16505_,
		_w16506_,
		_w16507_,
		_w16508_,
		_w16509_
	);
	LUT3 #(
		.INIT('h80)
	) name5997 (
		\wishbone_bd_ram_mem2_reg[19][17]/P0001 ,
		_w11935_,
		_w11938_,
		_w16510_
	);
	LUT3 #(
		.INIT('h80)
	) name5998 (
		\wishbone_bd_ram_mem2_reg[243][17]/P0001 ,
		_w11938_,
		_w11952_,
		_w16511_
	);
	LUT3 #(
		.INIT('h80)
	) name5999 (
		\wishbone_bd_ram_mem2_reg[122][17]/P0001 ,
		_w11944_,
		_w12012_,
		_w16512_
	);
	LUT3 #(
		.INIT('h80)
	) name6000 (
		\wishbone_bd_ram_mem2_reg[34][17]/P0001 ,
		_w11957_,
		_w11963_,
		_w16513_
	);
	LUT4 #(
		.INIT('h0001)
	) name6001 (
		_w16510_,
		_w16511_,
		_w16512_,
		_w16513_,
		_w16514_
	);
	LUT4 #(
		.INIT('h8000)
	) name6002 (
		_w16499_,
		_w16504_,
		_w16509_,
		_w16514_,
		_w16515_
	);
	LUT3 #(
		.INIT('h80)
	) name6003 (
		\wishbone_bd_ram_mem2_reg[146][17]/P0001 ,
		_w11959_,
		_w11963_,
		_w16516_
	);
	LUT3 #(
		.INIT('h80)
	) name6004 (
		\wishbone_bd_ram_mem2_reg[15][17]/P0001 ,
		_w11932_,
		_w11973_,
		_w16517_
	);
	LUT3 #(
		.INIT('h80)
	) name6005 (
		\wishbone_bd_ram_mem2_reg[44][17]/P0001 ,
		_w11954_,
		_w11957_,
		_w16518_
	);
	LUT3 #(
		.INIT('h80)
	) name6006 (
		\wishbone_bd_ram_mem2_reg[64][17]/P0001 ,
		_w11941_,
		_w11949_,
		_w16519_
	);
	LUT4 #(
		.INIT('h0001)
	) name6007 (
		_w16516_,
		_w16517_,
		_w16518_,
		_w16519_,
		_w16520_
	);
	LUT3 #(
		.INIT('h80)
	) name6008 (
		\wishbone_bd_ram_mem2_reg[119][17]/P0001 ,
		_w11975_,
		_w12012_,
		_w16521_
	);
	LUT3 #(
		.INIT('h80)
	) name6009 (
		\wishbone_bd_ram_mem2_reg[214][17]/P0001 ,
		_w11984_,
		_w11986_,
		_w16522_
	);
	LUT3 #(
		.INIT('h80)
	) name6010 (
		\wishbone_bd_ram_mem2_reg[96][17]/P0001 ,
		_w11941_,
		_w11965_,
		_w16523_
	);
	LUT3 #(
		.INIT('h80)
	) name6011 (
		\wishbone_bd_ram_mem2_reg[92][17]/P0001 ,
		_w11954_,
		_w11972_,
		_w16524_
	);
	LUT4 #(
		.INIT('h0001)
	) name6012 (
		_w16521_,
		_w16522_,
		_w16523_,
		_w16524_,
		_w16525_
	);
	LUT3 #(
		.INIT('h80)
	) name6013 (
		\wishbone_bd_ram_mem2_reg[253][17]/P0001 ,
		_w11952_,
		_w11966_,
		_w16526_
	);
	LUT3 #(
		.INIT('h80)
	) name6014 (
		\wishbone_bd_ram_mem2_reg[132][17]/P0001 ,
		_w11929_,
		_w11955_,
		_w16527_
	);
	LUT3 #(
		.INIT('h80)
	) name6015 (
		\wishbone_bd_ram_mem2_reg[149][17]/P0001 ,
		_w11933_,
		_w11959_,
		_w16528_
	);
	LUT3 #(
		.INIT('h80)
	) name6016 (
		\wishbone_bd_ram_mem2_reg[124][17]/P0001 ,
		_w11954_,
		_w12012_,
		_w16529_
	);
	LUT4 #(
		.INIT('h0001)
	) name6017 (
		_w16526_,
		_w16527_,
		_w16528_,
		_w16529_,
		_w16530_
	);
	LUT3 #(
		.INIT('h80)
	) name6018 (
		\wishbone_bd_ram_mem2_reg[63][17]/P0001 ,
		_w11973_,
		_w11979_,
		_w16531_
	);
	LUT3 #(
		.INIT('h80)
	) name6019 (
		\wishbone_bd_ram_mem2_reg[69][17]/P0001 ,
		_w11933_,
		_w11949_,
		_w16532_
	);
	LUT3 #(
		.INIT('h80)
	) name6020 (
		\wishbone_bd_ram_mem2_reg[85][17]/P0001 ,
		_w11933_,
		_w11972_,
		_w16533_
	);
	LUT3 #(
		.INIT('h80)
	) name6021 (
		\wishbone_bd_ram_mem2_reg[229][17]/P0001 ,
		_w11933_,
		_w11982_,
		_w16534_
	);
	LUT4 #(
		.INIT('h0001)
	) name6022 (
		_w16531_,
		_w16532_,
		_w16533_,
		_w16534_,
		_w16535_
	);
	LUT4 #(
		.INIT('h8000)
	) name6023 (
		_w16520_,
		_w16525_,
		_w16530_,
		_w16535_,
		_w16536_
	);
	LUT3 #(
		.INIT('h80)
	) name6024 (
		\wishbone_bd_ram_mem2_reg[49][17]/P0001 ,
		_w11977_,
		_w11979_,
		_w16537_
	);
	LUT3 #(
		.INIT('h80)
	) name6025 (
		\wishbone_bd_ram_mem2_reg[107][17]/P0001 ,
		_w11936_,
		_w11965_,
		_w16538_
	);
	LUT3 #(
		.INIT('h80)
	) name6026 (
		\wishbone_bd_ram_mem2_reg[184][17]/P0001 ,
		_w11942_,
		_w11990_,
		_w16539_
	);
	LUT3 #(
		.INIT('h80)
	) name6027 (
		\wishbone_bd_ram_mem2_reg[97][17]/P0001 ,
		_w11965_,
		_w11977_,
		_w16540_
	);
	LUT4 #(
		.INIT('h0001)
	) name6028 (
		_w16537_,
		_w16538_,
		_w16539_,
		_w16540_,
		_w16541_
	);
	LUT3 #(
		.INIT('h80)
	) name6029 (
		\wishbone_bd_ram_mem2_reg[134][17]/P0001 ,
		_w11955_,
		_w11986_,
		_w16542_
	);
	LUT3 #(
		.INIT('h80)
	) name6030 (
		\wishbone_bd_ram_mem2_reg[93][17]/P0001 ,
		_w11966_,
		_w11972_,
		_w16543_
	);
	LUT3 #(
		.INIT('h80)
	) name6031 (
		\wishbone_bd_ram_mem2_reg[56][17]/P0001 ,
		_w11979_,
		_w11990_,
		_w16544_
	);
	LUT3 #(
		.INIT('h80)
	) name6032 (
		\wishbone_bd_ram_mem2_reg[133][17]/P0001 ,
		_w11933_,
		_w11955_,
		_w16545_
	);
	LUT4 #(
		.INIT('h0001)
	) name6033 (
		_w16542_,
		_w16543_,
		_w16544_,
		_w16545_,
		_w16546_
	);
	LUT3 #(
		.INIT('h80)
	) name6034 (
		\wishbone_bd_ram_mem2_reg[195][17]/P0001 ,
		_w11938_,
		_w11945_,
		_w16547_
	);
	LUT3 #(
		.INIT('h80)
	) name6035 (
		\wishbone_bd_ram_mem2_reg[198][17]/P0001 ,
		_w11945_,
		_w11986_,
		_w16548_
	);
	LUT3 #(
		.INIT('h80)
	) name6036 (
		\wishbone_bd_ram_mem2_reg[240][17]/P0001 ,
		_w11941_,
		_w11952_,
		_w16549_
	);
	LUT3 #(
		.INIT('h80)
	) name6037 (
		\wishbone_bd_ram_mem2_reg[210][17]/P0001 ,
		_w11963_,
		_w11984_,
		_w16550_
	);
	LUT4 #(
		.INIT('h0001)
	) name6038 (
		_w16547_,
		_w16548_,
		_w16549_,
		_w16550_,
		_w16551_
	);
	LUT3 #(
		.INIT('h80)
	) name6039 (
		\wishbone_bd_ram_mem2_reg[45][17]/P0001 ,
		_w11957_,
		_w11966_,
		_w16552_
	);
	LUT3 #(
		.INIT('h80)
	) name6040 (
		\wishbone_bd_ram_mem2_reg[233][17]/P0001 ,
		_w11968_,
		_w11982_,
		_w16553_
	);
	LUT3 #(
		.INIT('h80)
	) name6041 (
		\wishbone_bd_ram_mem2_reg[162][17]/P0001 ,
		_w11930_,
		_w11963_,
		_w16554_
	);
	LUT3 #(
		.INIT('h80)
	) name6042 (
		\wishbone_bd_ram_mem2_reg[29][17]/P0001 ,
		_w11935_,
		_w11966_,
		_w16555_
	);
	LUT4 #(
		.INIT('h0001)
	) name6043 (
		_w16552_,
		_w16553_,
		_w16554_,
		_w16555_,
		_w16556_
	);
	LUT4 #(
		.INIT('h8000)
	) name6044 (
		_w16541_,
		_w16546_,
		_w16551_,
		_w16556_,
		_w16557_
	);
	LUT4 #(
		.INIT('h8000)
	) name6045 (
		_w16494_,
		_w16515_,
		_w16536_,
		_w16557_,
		_w16558_
	);
	LUT3 #(
		.INIT('h80)
	) name6046 (
		\wishbone_bd_ram_mem2_reg[130][17]/P0001 ,
		_w11955_,
		_w11963_,
		_w16559_
	);
	LUT3 #(
		.INIT('h80)
	) name6047 (
		\wishbone_bd_ram_mem2_reg[192][17]/P0001 ,
		_w11941_,
		_w11945_,
		_w16560_
	);
	LUT3 #(
		.INIT('h80)
	) name6048 (
		\wishbone_bd_ram_mem2_reg[218][17]/P0001 ,
		_w11944_,
		_w11984_,
		_w16561_
	);
	LUT3 #(
		.INIT('h80)
	) name6049 (
		\wishbone_bd_ram_mem2_reg[181][17]/P0001 ,
		_w11933_,
		_w11942_,
		_w16562_
	);
	LUT4 #(
		.INIT('h0001)
	) name6050 (
		_w16559_,
		_w16560_,
		_w16561_,
		_w16562_,
		_w16563_
	);
	LUT3 #(
		.INIT('h80)
	) name6051 (
		\wishbone_bd_ram_mem2_reg[147][17]/P0001 ,
		_w11938_,
		_w11959_,
		_w16564_
	);
	LUT3 #(
		.INIT('h80)
	) name6052 (
		\wishbone_bd_ram_mem2_reg[14][17]/P0001 ,
		_w11932_,
		_w11948_,
		_w16565_
	);
	LUT3 #(
		.INIT('h80)
	) name6053 (
		\wishbone_bd_ram_mem2_reg[48][17]/P0001 ,
		_w11941_,
		_w11979_,
		_w16566_
	);
	LUT3 #(
		.INIT('h80)
	) name6054 (
		\wishbone_bd_ram_mem2_reg[175][17]/P0001 ,
		_w11930_,
		_w11973_,
		_w16567_
	);
	LUT4 #(
		.INIT('h0001)
	) name6055 (
		_w16564_,
		_w16565_,
		_w16566_,
		_w16567_,
		_w16568_
	);
	LUT3 #(
		.INIT('h80)
	) name6056 (
		\wishbone_bd_ram_mem2_reg[250][17]/P0001 ,
		_w11944_,
		_w11952_,
		_w16569_
	);
	LUT3 #(
		.INIT('h80)
	) name6057 (
		\wishbone_bd_ram_mem2_reg[174][17]/P0001 ,
		_w11930_,
		_w11948_,
		_w16570_
	);
	LUT3 #(
		.INIT('h80)
	) name6058 (
		\wishbone_bd_ram_mem2_reg[223][17]/P0001 ,
		_w11973_,
		_w11984_,
		_w16571_
	);
	LUT3 #(
		.INIT('h80)
	) name6059 (
		\wishbone_bd_ram_mem2_reg[77][17]/P0001 ,
		_w11949_,
		_w11966_,
		_w16572_
	);
	LUT4 #(
		.INIT('h0001)
	) name6060 (
		_w16569_,
		_w16570_,
		_w16571_,
		_w16572_,
		_w16573_
	);
	LUT3 #(
		.INIT('h80)
	) name6061 (
		\wishbone_bd_ram_mem2_reg[226][17]/P0001 ,
		_w11963_,
		_w11982_,
		_w16574_
	);
	LUT3 #(
		.INIT('h80)
	) name6062 (
		\wishbone_bd_ram_mem2_reg[249][17]/P0001 ,
		_w11952_,
		_w11968_,
		_w16575_
	);
	LUT3 #(
		.INIT('h80)
	) name6063 (
		\wishbone_bd_ram_mem2_reg[25][17]/P0001 ,
		_w11935_,
		_w11968_,
		_w16576_
	);
	LUT3 #(
		.INIT('h80)
	) name6064 (
		\wishbone_bd_ram_mem2_reg[227][17]/P0001 ,
		_w11938_,
		_w11982_,
		_w16577_
	);
	LUT4 #(
		.INIT('h0001)
	) name6065 (
		_w16574_,
		_w16575_,
		_w16576_,
		_w16577_,
		_w16578_
	);
	LUT4 #(
		.INIT('h8000)
	) name6066 (
		_w16563_,
		_w16568_,
		_w16573_,
		_w16578_,
		_w16579_
	);
	LUT3 #(
		.INIT('h80)
	) name6067 (
		\wishbone_bd_ram_mem2_reg[145][17]/P0001 ,
		_w11959_,
		_w11977_,
		_w16580_
	);
	LUT3 #(
		.INIT('h80)
	) name6068 (
		\wishbone_bd_ram_mem2_reg[61][17]/P0001 ,
		_w11966_,
		_w11979_,
		_w16581_
	);
	LUT3 #(
		.INIT('h80)
	) name6069 (
		\wishbone_bd_ram_mem2_reg[55][17]/P0001 ,
		_w11975_,
		_w11979_,
		_w16582_
	);
	LUT3 #(
		.INIT('h80)
	) name6070 (
		\wishbone_bd_ram_mem2_reg[242][17]/P0001 ,
		_w11952_,
		_w11963_,
		_w16583_
	);
	LUT4 #(
		.INIT('h0001)
	) name6071 (
		_w16580_,
		_w16581_,
		_w16582_,
		_w16583_,
		_w16584_
	);
	LUT3 #(
		.INIT('h80)
	) name6072 (
		\wishbone_bd_ram_mem2_reg[26][17]/P0001 ,
		_w11935_,
		_w11944_,
		_w16585_
	);
	LUT3 #(
		.INIT('h80)
	) name6073 (
		\wishbone_bd_ram_mem2_reg[125][17]/P0001 ,
		_w11966_,
		_w12012_,
		_w16586_
	);
	LUT3 #(
		.INIT('h80)
	) name6074 (
		\wishbone_bd_ram_mem2_reg[89][17]/P0001 ,
		_w11968_,
		_w11972_,
		_w16587_
	);
	LUT3 #(
		.INIT('h80)
	) name6075 (
		\wishbone_bd_ram_mem2_reg[136][17]/P0001 ,
		_w11955_,
		_w11990_,
		_w16588_
	);
	LUT4 #(
		.INIT('h0001)
	) name6076 (
		_w16585_,
		_w16586_,
		_w16587_,
		_w16588_,
		_w16589_
	);
	LUT3 #(
		.INIT('h80)
	) name6077 (
		\wishbone_bd_ram_mem2_reg[167][17]/P0001 ,
		_w11930_,
		_w11975_,
		_w16590_
	);
	LUT3 #(
		.INIT('h80)
	) name6078 (
		\wishbone_bd_ram_mem2_reg[42][17]/P0001 ,
		_w11944_,
		_w11957_,
		_w16591_
	);
	LUT3 #(
		.INIT('h80)
	) name6079 (
		\wishbone_bd_ram_mem2_reg[27][17]/P0001 ,
		_w11935_,
		_w11936_,
		_w16592_
	);
	LUT3 #(
		.INIT('h80)
	) name6080 (
		\wishbone_bd_ram_mem2_reg[87][17]/P0001 ,
		_w11972_,
		_w11975_,
		_w16593_
	);
	LUT4 #(
		.INIT('h0001)
	) name6081 (
		_w16590_,
		_w16591_,
		_w16592_,
		_w16593_,
		_w16594_
	);
	LUT3 #(
		.INIT('h80)
	) name6082 (
		\wishbone_bd_ram_mem2_reg[30][17]/P0001 ,
		_w11935_,
		_w11948_,
		_w16595_
	);
	LUT3 #(
		.INIT('h80)
	) name6083 (
		\wishbone_bd_ram_mem2_reg[70][17]/P0001 ,
		_w11949_,
		_w11986_,
		_w16596_
	);
	LUT3 #(
		.INIT('h80)
	) name6084 (
		\wishbone_bd_ram_mem2_reg[46][17]/P0001 ,
		_w11948_,
		_w11957_,
		_w16597_
	);
	LUT3 #(
		.INIT('h80)
	) name6085 (
		\wishbone_bd_ram_mem2_reg[131][17]/P0001 ,
		_w11938_,
		_w11955_,
		_w16598_
	);
	LUT4 #(
		.INIT('h0001)
	) name6086 (
		_w16595_,
		_w16596_,
		_w16597_,
		_w16598_,
		_w16599_
	);
	LUT4 #(
		.INIT('h8000)
	) name6087 (
		_w16584_,
		_w16589_,
		_w16594_,
		_w16599_,
		_w16600_
	);
	LUT3 #(
		.INIT('h80)
	) name6088 (
		\wishbone_bd_ram_mem2_reg[158][17]/P0001 ,
		_w11948_,
		_w11959_,
		_w16601_
	);
	LUT3 #(
		.INIT('h80)
	) name6089 (
		\wishbone_bd_ram_mem2_reg[43][17]/P0001 ,
		_w11936_,
		_w11957_,
		_w16602_
	);
	LUT3 #(
		.INIT('h80)
	) name6090 (
		\wishbone_bd_ram_mem2_reg[11][17]/P0001 ,
		_w11932_,
		_w11936_,
		_w16603_
	);
	LUT3 #(
		.INIT('h80)
	) name6091 (
		\wishbone_bd_ram_mem2_reg[178][17]/P0001 ,
		_w11942_,
		_w11963_,
		_w16604_
	);
	LUT4 #(
		.INIT('h0001)
	) name6092 (
		_w16601_,
		_w16602_,
		_w16603_,
		_w16604_,
		_w16605_
	);
	LUT3 #(
		.INIT('h80)
	) name6093 (
		\wishbone_bd_ram_mem2_reg[111][17]/P0001 ,
		_w11965_,
		_w11973_,
		_w16606_
	);
	LUT3 #(
		.INIT('h80)
	) name6094 (
		\wishbone_bd_ram_mem2_reg[152][17]/P0001 ,
		_w11959_,
		_w11990_,
		_w16607_
	);
	LUT3 #(
		.INIT('h80)
	) name6095 (
		\wishbone_bd_ram_mem2_reg[177][17]/P0001 ,
		_w11942_,
		_w11977_,
		_w16608_
	);
	LUT3 #(
		.INIT('h80)
	) name6096 (
		\wishbone_bd_ram_mem2_reg[52][17]/P0001 ,
		_w11929_,
		_w11979_,
		_w16609_
	);
	LUT4 #(
		.INIT('h0001)
	) name6097 (
		_w16606_,
		_w16607_,
		_w16608_,
		_w16609_,
		_w16610_
	);
	LUT3 #(
		.INIT('h80)
	) name6098 (
		\wishbone_bd_ram_mem2_reg[139][17]/P0001 ,
		_w11936_,
		_w11955_,
		_w16611_
	);
	LUT3 #(
		.INIT('h80)
	) name6099 (
		\wishbone_bd_ram_mem2_reg[116][17]/P0001 ,
		_w11929_,
		_w12012_,
		_w16612_
	);
	LUT3 #(
		.INIT('h80)
	) name6100 (
		\wishbone_bd_ram_mem2_reg[36][17]/P0001 ,
		_w11929_,
		_w11957_,
		_w16613_
	);
	LUT3 #(
		.INIT('h80)
	) name6101 (
		\wishbone_bd_ram_mem2_reg[201][17]/P0001 ,
		_w11945_,
		_w11968_,
		_w16614_
	);
	LUT4 #(
		.INIT('h0001)
	) name6102 (
		_w16611_,
		_w16612_,
		_w16613_,
		_w16614_,
		_w16615_
	);
	LUT3 #(
		.INIT('h80)
	) name6103 (
		\wishbone_bd_ram_mem2_reg[67][17]/P0001 ,
		_w11938_,
		_w11949_,
		_w16616_
	);
	LUT3 #(
		.INIT('h80)
	) name6104 (
		\wishbone_bd_ram_mem2_reg[0][17]/P0001 ,
		_w11932_,
		_w11941_,
		_w16617_
	);
	LUT3 #(
		.INIT('h80)
	) name6105 (
		\wishbone_bd_ram_mem2_reg[72][17]/P0001 ,
		_w11949_,
		_w11990_,
		_w16618_
	);
	LUT3 #(
		.INIT('h80)
	) name6106 (
		\wishbone_bd_ram_mem2_reg[2][17]/P0001 ,
		_w11932_,
		_w11963_,
		_w16619_
	);
	LUT4 #(
		.INIT('h0001)
	) name6107 (
		_w16616_,
		_w16617_,
		_w16618_,
		_w16619_,
		_w16620_
	);
	LUT4 #(
		.INIT('h8000)
	) name6108 (
		_w16605_,
		_w16610_,
		_w16615_,
		_w16620_,
		_w16621_
	);
	LUT3 #(
		.INIT('h80)
	) name6109 (
		\wishbone_bd_ram_mem2_reg[98][17]/P0001 ,
		_w11963_,
		_w11965_,
		_w16622_
	);
	LUT3 #(
		.INIT('h80)
	) name6110 (
		\wishbone_bd_ram_mem2_reg[236][17]/P0001 ,
		_w11954_,
		_w11982_,
		_w16623_
	);
	LUT3 #(
		.INIT('h80)
	) name6111 (
		\wishbone_bd_ram_mem2_reg[37][17]/P0001 ,
		_w11933_,
		_w11957_,
		_w16624_
	);
	LUT3 #(
		.INIT('h80)
	) name6112 (
		\wishbone_bd_ram_mem2_reg[66][17]/P0001 ,
		_w11949_,
		_w11963_,
		_w16625_
	);
	LUT4 #(
		.INIT('h0001)
	) name6113 (
		_w16622_,
		_w16623_,
		_w16624_,
		_w16625_,
		_w16626_
	);
	LUT3 #(
		.INIT('h80)
	) name6114 (
		\wishbone_bd_ram_mem2_reg[185][17]/P0001 ,
		_w11942_,
		_w11968_,
		_w16627_
	);
	LUT3 #(
		.INIT('h80)
	) name6115 (
		\wishbone_bd_ram_mem2_reg[21][17]/P0001 ,
		_w11933_,
		_w11935_,
		_w16628_
	);
	LUT3 #(
		.INIT('h80)
	) name6116 (
		\wishbone_bd_ram_mem2_reg[73][17]/P0001 ,
		_w11949_,
		_w11968_,
		_w16629_
	);
	LUT3 #(
		.INIT('h80)
	) name6117 (
		\wishbone_bd_ram_mem2_reg[219][17]/P0001 ,
		_w11936_,
		_w11984_,
		_w16630_
	);
	LUT4 #(
		.INIT('h0001)
	) name6118 (
		_w16627_,
		_w16628_,
		_w16629_,
		_w16630_,
		_w16631_
	);
	LUT3 #(
		.INIT('h80)
	) name6119 (
		\wishbone_bd_ram_mem2_reg[129][17]/P0001 ,
		_w11955_,
		_w11977_,
		_w16632_
	);
	LUT3 #(
		.INIT('h80)
	) name6120 (
		\wishbone_bd_ram_mem2_reg[62][17]/P0001 ,
		_w11948_,
		_w11979_,
		_w16633_
	);
	LUT3 #(
		.INIT('h80)
	) name6121 (
		\wishbone_bd_ram_mem2_reg[82][17]/P0001 ,
		_w11963_,
		_w11972_,
		_w16634_
	);
	LUT3 #(
		.INIT('h80)
	) name6122 (
		\wishbone_bd_ram_mem2_reg[156][17]/P0001 ,
		_w11954_,
		_w11959_,
		_w16635_
	);
	LUT4 #(
		.INIT('h0001)
	) name6123 (
		_w16632_,
		_w16633_,
		_w16634_,
		_w16635_,
		_w16636_
	);
	LUT3 #(
		.INIT('h80)
	) name6124 (
		\wishbone_bd_ram_mem2_reg[16][17]/P0001 ,
		_w11935_,
		_w11941_,
		_w16637_
	);
	LUT3 #(
		.INIT('h80)
	) name6125 (
		\wishbone_bd_ram_mem2_reg[126][17]/P0001 ,
		_w11948_,
		_w12012_,
		_w16638_
	);
	LUT3 #(
		.INIT('h80)
	) name6126 (
		\wishbone_bd_ram_mem2_reg[228][17]/P0001 ,
		_w11929_,
		_w11982_,
		_w16639_
	);
	LUT3 #(
		.INIT('h80)
	) name6127 (
		\wishbone_bd_ram_mem2_reg[80][17]/P0001 ,
		_w11941_,
		_w11972_,
		_w16640_
	);
	LUT4 #(
		.INIT('h0001)
	) name6128 (
		_w16637_,
		_w16638_,
		_w16639_,
		_w16640_,
		_w16641_
	);
	LUT4 #(
		.INIT('h8000)
	) name6129 (
		_w16626_,
		_w16631_,
		_w16636_,
		_w16641_,
		_w16642_
	);
	LUT4 #(
		.INIT('h8000)
	) name6130 (
		_w16579_,
		_w16600_,
		_w16621_,
		_w16642_,
		_w16643_
	);
	LUT3 #(
		.INIT('h80)
	) name6131 (
		\wishbone_bd_ram_mem2_reg[224][17]/P0001 ,
		_w11941_,
		_w11982_,
		_w16644_
	);
	LUT3 #(
		.INIT('h80)
	) name6132 (
		\wishbone_bd_ram_mem2_reg[179][17]/P0001 ,
		_w11938_,
		_w11942_,
		_w16645_
	);
	LUT3 #(
		.INIT('h80)
	) name6133 (
		\wishbone_bd_ram_mem2_reg[54][17]/P0001 ,
		_w11979_,
		_w11986_,
		_w16646_
	);
	LUT3 #(
		.INIT('h80)
	) name6134 (
		\wishbone_bd_ram_mem2_reg[5][17]/P0001 ,
		_w11932_,
		_w11933_,
		_w16647_
	);
	LUT4 #(
		.INIT('h0001)
	) name6135 (
		_w16644_,
		_w16645_,
		_w16646_,
		_w16647_,
		_w16648_
	);
	LUT3 #(
		.INIT('h80)
	) name6136 (
		\wishbone_bd_ram_mem2_reg[104][17]/P0001 ,
		_w11965_,
		_w11990_,
		_w16649_
	);
	LUT3 #(
		.INIT('h80)
	) name6137 (
		\wishbone_bd_ram_mem2_reg[154][17]/P0001 ,
		_w11944_,
		_w11959_,
		_w16650_
	);
	LUT3 #(
		.INIT('h80)
	) name6138 (
		\wishbone_bd_ram_mem2_reg[115][17]/P0001 ,
		_w11938_,
		_w12012_,
		_w16651_
	);
	LUT3 #(
		.INIT('h80)
	) name6139 (
		\wishbone_bd_ram_mem2_reg[108][17]/P0001 ,
		_w11954_,
		_w11965_,
		_w16652_
	);
	LUT4 #(
		.INIT('h0001)
	) name6140 (
		_w16649_,
		_w16650_,
		_w16651_,
		_w16652_,
		_w16653_
	);
	LUT3 #(
		.INIT('h80)
	) name6141 (
		\wishbone_bd_ram_mem2_reg[196][17]/P0001 ,
		_w11929_,
		_w11945_,
		_w16654_
	);
	LUT3 #(
		.INIT('h80)
	) name6142 (
		\wishbone_bd_ram_mem2_reg[114][17]/P0001 ,
		_w11963_,
		_w12012_,
		_w16655_
	);
	LUT3 #(
		.INIT('h80)
	) name6143 (
		\wishbone_bd_ram_mem2_reg[38][17]/P0001 ,
		_w11957_,
		_w11986_,
		_w16656_
	);
	LUT3 #(
		.INIT('h80)
	) name6144 (
		\wishbone_bd_ram_mem2_reg[215][17]/P0001 ,
		_w11975_,
		_w11984_,
		_w16657_
	);
	LUT4 #(
		.INIT('h0001)
	) name6145 (
		_w16654_,
		_w16655_,
		_w16656_,
		_w16657_,
		_w16658_
	);
	LUT3 #(
		.INIT('h80)
	) name6146 (
		\wishbone_bd_ram_mem2_reg[202][17]/P0001 ,
		_w11944_,
		_w11945_,
		_w16659_
	);
	LUT3 #(
		.INIT('h80)
	) name6147 (
		\wishbone_bd_ram_mem2_reg[110][17]/P0001 ,
		_w11948_,
		_w11965_,
		_w16660_
	);
	LUT3 #(
		.INIT('h80)
	) name6148 (
		\wishbone_bd_ram_mem2_reg[135][17]/P0001 ,
		_w11955_,
		_w11975_,
		_w16661_
	);
	LUT3 #(
		.INIT('h80)
	) name6149 (
		\wishbone_bd_ram_mem2_reg[109][17]/P0001 ,
		_w11965_,
		_w11966_,
		_w16662_
	);
	LUT4 #(
		.INIT('h0001)
	) name6150 (
		_w16659_,
		_w16660_,
		_w16661_,
		_w16662_,
		_w16663_
	);
	LUT4 #(
		.INIT('h8000)
	) name6151 (
		_w16648_,
		_w16653_,
		_w16658_,
		_w16663_,
		_w16664_
	);
	LUT3 #(
		.INIT('h80)
	) name6152 (
		\wishbone_bd_ram_mem2_reg[189][17]/P0001 ,
		_w11942_,
		_w11966_,
		_w16665_
	);
	LUT3 #(
		.INIT('h80)
	) name6153 (
		\wishbone_bd_ram_mem2_reg[75][17]/P0001 ,
		_w11936_,
		_w11949_,
		_w16666_
	);
	LUT3 #(
		.INIT('h80)
	) name6154 (
		\wishbone_bd_ram_mem2_reg[197][17]/P0001 ,
		_w11933_,
		_w11945_,
		_w16667_
	);
	LUT3 #(
		.INIT('h80)
	) name6155 (
		\wishbone_bd_ram_mem2_reg[254][17]/P0001 ,
		_w11948_,
		_w11952_,
		_w16668_
	);
	LUT4 #(
		.INIT('h0001)
	) name6156 (
		_w16665_,
		_w16666_,
		_w16667_,
		_w16668_,
		_w16669_
	);
	LUT3 #(
		.INIT('h80)
	) name6157 (
		\wishbone_bd_ram_mem2_reg[59][17]/P0001 ,
		_w11936_,
		_w11979_,
		_w16670_
	);
	LUT3 #(
		.INIT('h80)
	) name6158 (
		\wishbone_bd_ram_mem2_reg[204][17]/P0001 ,
		_w11945_,
		_w11954_,
		_w16671_
	);
	LUT3 #(
		.INIT('h80)
	) name6159 (
		\wishbone_bd_ram_mem2_reg[88][17]/P0001 ,
		_w11972_,
		_w11990_,
		_w16672_
	);
	LUT3 #(
		.INIT('h80)
	) name6160 (
		\wishbone_bd_ram_mem2_reg[182][17]/P0001 ,
		_w11942_,
		_w11986_,
		_w16673_
	);
	LUT4 #(
		.INIT('h0001)
	) name6161 (
		_w16670_,
		_w16671_,
		_w16672_,
		_w16673_,
		_w16674_
	);
	LUT3 #(
		.INIT('h80)
	) name6162 (
		\wishbone_bd_ram_mem2_reg[17][17]/P0001 ,
		_w11935_,
		_w11977_,
		_w16675_
	);
	LUT3 #(
		.INIT('h80)
	) name6163 (
		\wishbone_bd_ram_mem2_reg[103][17]/P0001 ,
		_w11965_,
		_w11975_,
		_w16676_
	);
	LUT3 #(
		.INIT('h80)
	) name6164 (
		\wishbone_bd_ram_mem2_reg[120][17]/P0001 ,
		_w11990_,
		_w12012_,
		_w16677_
	);
	LUT3 #(
		.INIT('h80)
	) name6165 (
		\wishbone_bd_ram_mem2_reg[190][17]/P0001 ,
		_w11942_,
		_w11948_,
		_w16678_
	);
	LUT4 #(
		.INIT('h0001)
	) name6166 (
		_w16675_,
		_w16676_,
		_w16677_,
		_w16678_,
		_w16679_
	);
	LUT3 #(
		.INIT('h80)
	) name6167 (
		\wishbone_bd_ram_mem2_reg[199][17]/P0001 ,
		_w11945_,
		_w11975_,
		_w16680_
	);
	LUT3 #(
		.INIT('h80)
	) name6168 (
		\wishbone_bd_ram_mem2_reg[141][17]/P0001 ,
		_w11955_,
		_w11966_,
		_w16681_
	);
	LUT3 #(
		.INIT('h80)
	) name6169 (
		\wishbone_bd_ram_mem2_reg[159][17]/P0001 ,
		_w11959_,
		_w11973_,
		_w16682_
	);
	LUT3 #(
		.INIT('h80)
	) name6170 (
		\wishbone_bd_ram_mem2_reg[169][17]/P0001 ,
		_w11930_,
		_w11968_,
		_w16683_
	);
	LUT4 #(
		.INIT('h0001)
	) name6171 (
		_w16680_,
		_w16681_,
		_w16682_,
		_w16683_,
		_w16684_
	);
	LUT4 #(
		.INIT('h8000)
	) name6172 (
		_w16669_,
		_w16674_,
		_w16679_,
		_w16684_,
		_w16685_
	);
	LUT3 #(
		.INIT('h80)
	) name6173 (
		\wishbone_bd_ram_mem2_reg[18][17]/P0001 ,
		_w11935_,
		_w11963_,
		_w16686_
	);
	LUT3 #(
		.INIT('h80)
	) name6174 (
		\wishbone_bd_ram_mem2_reg[68][17]/P0001 ,
		_w11929_,
		_w11949_,
		_w16687_
	);
	LUT3 #(
		.INIT('h80)
	) name6175 (
		\wishbone_bd_ram_mem2_reg[95][17]/P0001 ,
		_w11972_,
		_w11973_,
		_w16688_
	);
	LUT3 #(
		.INIT('h80)
	) name6176 (
		\wishbone_bd_ram_mem2_reg[170][17]/P0001 ,
		_w11930_,
		_w11944_,
		_w16689_
	);
	LUT4 #(
		.INIT('h0001)
	) name6177 (
		_w16686_,
		_w16687_,
		_w16688_,
		_w16689_,
		_w16690_
	);
	LUT3 #(
		.INIT('h80)
	) name6178 (
		\wishbone_bd_ram_mem2_reg[235][17]/P0001 ,
		_w11936_,
		_w11982_,
		_w16691_
	);
	LUT3 #(
		.INIT('h80)
	) name6179 (
		\wishbone_bd_ram_mem2_reg[94][17]/P0001 ,
		_w11948_,
		_w11972_,
		_w16692_
	);
	LUT3 #(
		.INIT('h80)
	) name6180 (
		\wishbone_bd_ram_mem2_reg[106][17]/P0001 ,
		_w11944_,
		_w11965_,
		_w16693_
	);
	LUT3 #(
		.INIT('h80)
	) name6181 (
		\wishbone_bd_ram_mem2_reg[79][17]/P0001 ,
		_w11949_,
		_w11973_,
		_w16694_
	);
	LUT4 #(
		.INIT('h0001)
	) name6182 (
		_w16691_,
		_w16692_,
		_w16693_,
		_w16694_,
		_w16695_
	);
	LUT3 #(
		.INIT('h80)
	) name6183 (
		\wishbone_bd_ram_mem2_reg[188][17]/P0001 ,
		_w11942_,
		_w11954_,
		_w16696_
	);
	LUT3 #(
		.INIT('h80)
	) name6184 (
		\wishbone_bd_ram_mem2_reg[81][17]/P0001 ,
		_w11972_,
		_w11977_,
		_w16697_
	);
	LUT3 #(
		.INIT('h80)
	) name6185 (
		\wishbone_bd_ram_mem2_reg[171][17]/P0001 ,
		_w11930_,
		_w11936_,
		_w16698_
	);
	LUT3 #(
		.INIT('h80)
	) name6186 (
		\wishbone_bd_ram_mem2_reg[238][17]/P0001 ,
		_w11948_,
		_w11982_,
		_w16699_
	);
	LUT4 #(
		.INIT('h0001)
	) name6187 (
		_w16696_,
		_w16697_,
		_w16698_,
		_w16699_,
		_w16700_
	);
	LUT3 #(
		.INIT('h80)
	) name6188 (
		\wishbone_bd_ram_mem2_reg[246][17]/P0001 ,
		_w11952_,
		_w11986_,
		_w16701_
	);
	LUT3 #(
		.INIT('h80)
	) name6189 (
		\wishbone_bd_ram_mem2_reg[150][17]/P0001 ,
		_w11959_,
		_w11986_,
		_w16702_
	);
	LUT3 #(
		.INIT('h80)
	) name6190 (
		\wishbone_bd_ram_mem2_reg[140][17]/P0001 ,
		_w11954_,
		_w11955_,
		_w16703_
	);
	LUT3 #(
		.INIT('h80)
	) name6191 (
		\wishbone_bd_ram_mem2_reg[255][17]/P0001 ,
		_w11952_,
		_w11973_,
		_w16704_
	);
	LUT4 #(
		.INIT('h0001)
	) name6192 (
		_w16701_,
		_w16702_,
		_w16703_,
		_w16704_,
		_w16705_
	);
	LUT4 #(
		.INIT('h8000)
	) name6193 (
		_w16690_,
		_w16695_,
		_w16700_,
		_w16705_,
		_w16706_
	);
	LUT3 #(
		.INIT('h80)
	) name6194 (
		\wishbone_bd_ram_mem2_reg[252][17]/P0001 ,
		_w11952_,
		_w11954_,
		_w16707_
	);
	LUT3 #(
		.INIT('h80)
	) name6195 (
		\wishbone_bd_ram_mem2_reg[191][17]/P0001 ,
		_w11942_,
		_w11973_,
		_w16708_
	);
	LUT3 #(
		.INIT('h80)
	) name6196 (
		\wishbone_bd_ram_mem2_reg[7][17]/P0001 ,
		_w11932_,
		_w11975_,
		_w16709_
	);
	LUT3 #(
		.INIT('h80)
	) name6197 (
		\wishbone_bd_ram_mem2_reg[100][17]/P0001 ,
		_w11929_,
		_w11965_,
		_w16710_
	);
	LUT4 #(
		.INIT('h0001)
	) name6198 (
		_w16707_,
		_w16708_,
		_w16709_,
		_w16710_,
		_w16711_
	);
	LUT3 #(
		.INIT('h80)
	) name6199 (
		\wishbone_bd_ram_mem2_reg[216][17]/P0001 ,
		_w11984_,
		_w11990_,
		_w16712_
	);
	LUT3 #(
		.INIT('h80)
	) name6200 (
		\wishbone_bd_ram_mem2_reg[225][17]/P0001 ,
		_w11977_,
		_w11982_,
		_w16713_
	);
	LUT3 #(
		.INIT('h80)
	) name6201 (
		\wishbone_bd_ram_mem2_reg[203][17]/P0001 ,
		_w11936_,
		_w11945_,
		_w16714_
	);
	LUT3 #(
		.INIT('h80)
	) name6202 (
		\wishbone_bd_ram_mem2_reg[4][17]/P0001 ,
		_w11929_,
		_w11932_,
		_w16715_
	);
	LUT4 #(
		.INIT('h0001)
	) name6203 (
		_w16712_,
		_w16713_,
		_w16714_,
		_w16715_,
		_w16716_
	);
	LUT3 #(
		.INIT('h80)
	) name6204 (
		\wishbone_bd_ram_mem2_reg[74][17]/P0001 ,
		_w11944_,
		_w11949_,
		_w16717_
	);
	LUT3 #(
		.INIT('h80)
	) name6205 (
		\wishbone_bd_ram_mem2_reg[164][17]/P0001 ,
		_w11929_,
		_w11930_,
		_w16718_
	);
	LUT3 #(
		.INIT('h80)
	) name6206 (
		\wishbone_bd_ram_mem2_reg[83][17]/P0001 ,
		_w11938_,
		_w11972_,
		_w16719_
	);
	LUT3 #(
		.INIT('h80)
	) name6207 (
		\wishbone_bd_ram_mem2_reg[121][17]/P0001 ,
		_w11968_,
		_w12012_,
		_w16720_
	);
	LUT4 #(
		.INIT('h0001)
	) name6208 (
		_w16717_,
		_w16718_,
		_w16719_,
		_w16720_,
		_w16721_
	);
	LUT3 #(
		.INIT('h80)
	) name6209 (
		\wishbone_bd_ram_mem2_reg[6][17]/P0001 ,
		_w11932_,
		_w11986_,
		_w16722_
	);
	LUT3 #(
		.INIT('h80)
	) name6210 (
		\wishbone_bd_ram_mem2_reg[157][17]/P0001 ,
		_w11959_,
		_w11966_,
		_w16723_
	);
	LUT3 #(
		.INIT('h80)
	) name6211 (
		\wishbone_bd_ram_mem2_reg[241][17]/P0001 ,
		_w11952_,
		_w11977_,
		_w16724_
	);
	LUT3 #(
		.INIT('h80)
	) name6212 (
		\wishbone_bd_ram_mem2_reg[186][17]/P0001 ,
		_w11942_,
		_w11944_,
		_w16725_
	);
	LUT4 #(
		.INIT('h0001)
	) name6213 (
		_w16722_,
		_w16723_,
		_w16724_,
		_w16725_,
		_w16726_
	);
	LUT4 #(
		.INIT('h8000)
	) name6214 (
		_w16711_,
		_w16716_,
		_w16721_,
		_w16726_,
		_w16727_
	);
	LUT4 #(
		.INIT('h8000)
	) name6215 (
		_w16664_,
		_w16685_,
		_w16706_,
		_w16727_,
		_w16728_
	);
	LUT3 #(
		.INIT('h80)
	) name6216 (
		\wishbone_bd_ram_mem2_reg[200][17]/P0001 ,
		_w11945_,
		_w11990_,
		_w16729_
	);
	LUT3 #(
		.INIT('h80)
	) name6217 (
		\wishbone_bd_ram_mem2_reg[248][17]/P0001 ,
		_w11952_,
		_w11990_,
		_w16730_
	);
	LUT3 #(
		.INIT('h80)
	) name6218 (
		\wishbone_bd_ram_mem2_reg[31][17]/P0001 ,
		_w11935_,
		_w11973_,
		_w16731_
	);
	LUT3 #(
		.INIT('h80)
	) name6219 (
		\wishbone_bd_ram_mem2_reg[232][17]/P0001 ,
		_w11982_,
		_w11990_,
		_w16732_
	);
	LUT4 #(
		.INIT('h0001)
	) name6220 (
		_w16729_,
		_w16730_,
		_w16731_,
		_w16732_,
		_w16733_
	);
	LUT3 #(
		.INIT('h80)
	) name6221 (
		\wishbone_bd_ram_mem2_reg[165][17]/P0001 ,
		_w11930_,
		_w11933_,
		_w16734_
	);
	LUT3 #(
		.INIT('h80)
	) name6222 (
		\wishbone_bd_ram_mem2_reg[1][17]/P0001 ,
		_w11932_,
		_w11977_,
		_w16735_
	);
	LUT3 #(
		.INIT('h80)
	) name6223 (
		\wishbone_bd_ram_mem2_reg[244][17]/P0001 ,
		_w11929_,
		_w11952_,
		_w16736_
	);
	LUT3 #(
		.INIT('h80)
	) name6224 (
		\wishbone_bd_ram_mem2_reg[247][17]/P0001 ,
		_w11952_,
		_w11975_,
		_w16737_
	);
	LUT4 #(
		.INIT('h0001)
	) name6225 (
		_w16734_,
		_w16735_,
		_w16736_,
		_w16737_,
		_w16738_
	);
	LUT3 #(
		.INIT('h80)
	) name6226 (
		\wishbone_bd_ram_mem2_reg[239][17]/P0001 ,
		_w11973_,
		_w11982_,
		_w16739_
	);
	LUT3 #(
		.INIT('h80)
	) name6227 (
		\wishbone_bd_ram_mem2_reg[123][17]/P0001 ,
		_w11936_,
		_w12012_,
		_w16740_
	);
	LUT3 #(
		.INIT('h80)
	) name6228 (
		\wishbone_bd_ram_mem2_reg[99][17]/P0001 ,
		_w11938_,
		_w11965_,
		_w16741_
	);
	LUT3 #(
		.INIT('h80)
	) name6229 (
		\wishbone_bd_ram_mem2_reg[86][17]/P0001 ,
		_w11972_,
		_w11986_,
		_w16742_
	);
	LUT4 #(
		.INIT('h0001)
	) name6230 (
		_w16739_,
		_w16740_,
		_w16741_,
		_w16742_,
		_w16743_
	);
	LUT3 #(
		.INIT('h80)
	) name6231 (
		\wishbone_bd_ram_mem2_reg[163][17]/P0001 ,
		_w11930_,
		_w11938_,
		_w16744_
	);
	LUT3 #(
		.INIT('h80)
	) name6232 (
		\wishbone_bd_ram_mem2_reg[208][17]/P0001 ,
		_w11941_,
		_w11984_,
		_w16745_
	);
	LUT3 #(
		.INIT('h80)
	) name6233 (
		\wishbone_bd_ram_mem2_reg[101][17]/P0001 ,
		_w11933_,
		_w11965_,
		_w16746_
	);
	LUT3 #(
		.INIT('h80)
	) name6234 (
		\wishbone_bd_ram_mem2_reg[211][17]/P0001 ,
		_w11938_,
		_w11984_,
		_w16747_
	);
	LUT4 #(
		.INIT('h0001)
	) name6235 (
		_w16744_,
		_w16745_,
		_w16746_,
		_w16747_,
		_w16748_
	);
	LUT4 #(
		.INIT('h8000)
	) name6236 (
		_w16733_,
		_w16738_,
		_w16743_,
		_w16748_,
		_w16749_
	);
	LUT3 #(
		.INIT('h80)
	) name6237 (
		\wishbone_bd_ram_mem2_reg[172][17]/P0001 ,
		_w11930_,
		_w11954_,
		_w16750_
	);
	LUT3 #(
		.INIT('h80)
	) name6238 (
		\wishbone_bd_ram_mem2_reg[153][17]/P0001 ,
		_w11959_,
		_w11968_,
		_w16751_
	);
	LUT3 #(
		.INIT('h80)
	) name6239 (
		\wishbone_bd_ram_mem2_reg[220][17]/P0001 ,
		_w11954_,
		_w11984_,
		_w16752_
	);
	LUT3 #(
		.INIT('h80)
	) name6240 (
		\wishbone_bd_ram_mem2_reg[112][17]/P0001 ,
		_w11941_,
		_w12012_,
		_w16753_
	);
	LUT4 #(
		.INIT('h0001)
	) name6241 (
		_w16750_,
		_w16751_,
		_w16752_,
		_w16753_,
		_w16754_
	);
	LUT3 #(
		.INIT('h80)
	) name6242 (
		\wishbone_bd_ram_mem2_reg[205][17]/P0001 ,
		_w11945_,
		_w11966_,
		_w16755_
	);
	LUT3 #(
		.INIT('h80)
	) name6243 (
		\wishbone_bd_ram_mem2_reg[155][17]/P0001 ,
		_w11936_,
		_w11959_,
		_w16756_
	);
	LUT3 #(
		.INIT('h80)
	) name6244 (
		\wishbone_bd_ram_mem2_reg[230][17]/P0001 ,
		_w11982_,
		_w11986_,
		_w16757_
	);
	LUT3 #(
		.INIT('h80)
	) name6245 (
		\wishbone_bd_ram_mem2_reg[20][17]/P0001 ,
		_w11929_,
		_w11935_,
		_w16758_
	);
	LUT4 #(
		.INIT('h0001)
	) name6246 (
		_w16755_,
		_w16756_,
		_w16757_,
		_w16758_,
		_w16759_
	);
	LUT3 #(
		.INIT('h80)
	) name6247 (
		\wishbone_bd_ram_mem2_reg[58][17]/P0001 ,
		_w11944_,
		_w11979_,
		_w16760_
	);
	LUT3 #(
		.INIT('h80)
	) name6248 (
		\wishbone_bd_ram_mem2_reg[138][17]/P0001 ,
		_w11944_,
		_w11955_,
		_w16761_
	);
	LUT3 #(
		.INIT('h80)
	) name6249 (
		\wishbone_bd_ram_mem2_reg[35][17]/P0001 ,
		_w11938_,
		_w11957_,
		_w16762_
	);
	LUT3 #(
		.INIT('h80)
	) name6250 (
		\wishbone_bd_ram_mem2_reg[222][17]/P0001 ,
		_w11948_,
		_w11984_,
		_w16763_
	);
	LUT4 #(
		.INIT('h0001)
	) name6251 (
		_w16760_,
		_w16761_,
		_w16762_,
		_w16763_,
		_w16764_
	);
	LUT3 #(
		.INIT('h80)
	) name6252 (
		\wishbone_bd_ram_mem2_reg[3][17]/P0001 ,
		_w11932_,
		_w11938_,
		_w16765_
	);
	LUT3 #(
		.INIT('h80)
	) name6253 (
		\wishbone_bd_ram_mem2_reg[245][17]/P0001 ,
		_w11933_,
		_w11952_,
		_w16766_
	);
	LUT3 #(
		.INIT('h80)
	) name6254 (
		\wishbone_bd_ram_mem2_reg[118][17]/P0001 ,
		_w11986_,
		_w12012_,
		_w16767_
	);
	LUT3 #(
		.INIT('h80)
	) name6255 (
		\wishbone_bd_ram_mem2_reg[28][17]/P0001 ,
		_w11935_,
		_w11954_,
		_w16768_
	);
	LUT4 #(
		.INIT('h0001)
	) name6256 (
		_w16765_,
		_w16766_,
		_w16767_,
		_w16768_,
		_w16769_
	);
	LUT4 #(
		.INIT('h8000)
	) name6257 (
		_w16754_,
		_w16759_,
		_w16764_,
		_w16769_,
		_w16770_
	);
	LUT3 #(
		.INIT('h80)
	) name6258 (
		\wishbone_bd_ram_mem2_reg[187][17]/P0001 ,
		_w11936_,
		_w11942_,
		_w16771_
	);
	LUT3 #(
		.INIT('h80)
	) name6259 (
		\wishbone_bd_ram_mem2_reg[137][17]/P0001 ,
		_w11955_,
		_w11968_,
		_w16772_
	);
	LUT3 #(
		.INIT('h80)
	) name6260 (
		\wishbone_bd_ram_mem2_reg[8][17]/P0001 ,
		_w11932_,
		_w11990_,
		_w16773_
	);
	LUT3 #(
		.INIT('h80)
	) name6261 (
		\wishbone_bd_ram_mem2_reg[53][17]/P0001 ,
		_w11933_,
		_w11979_,
		_w16774_
	);
	LUT4 #(
		.INIT('h0001)
	) name6262 (
		_w16771_,
		_w16772_,
		_w16773_,
		_w16774_,
		_w16775_
	);
	LUT3 #(
		.INIT('h80)
	) name6263 (
		\wishbone_bd_ram_mem2_reg[91][17]/P0001 ,
		_w11936_,
		_w11972_,
		_w16776_
	);
	LUT3 #(
		.INIT('h80)
	) name6264 (
		\wishbone_bd_ram_mem2_reg[221][17]/P0001 ,
		_w11966_,
		_w11984_,
		_w16777_
	);
	LUT3 #(
		.INIT('h80)
	) name6265 (
		\wishbone_bd_ram_mem2_reg[206][17]/P0001 ,
		_w11945_,
		_w11948_,
		_w16778_
	);
	LUT3 #(
		.INIT('h80)
	) name6266 (
		\wishbone_bd_ram_mem2_reg[194][17]/P0001 ,
		_w11945_,
		_w11963_,
		_w16779_
	);
	LUT4 #(
		.INIT('h0001)
	) name6267 (
		_w16776_,
		_w16777_,
		_w16778_,
		_w16779_,
		_w16780_
	);
	LUT3 #(
		.INIT('h80)
	) name6268 (
		\wishbone_bd_ram_mem2_reg[39][17]/P0001 ,
		_w11957_,
		_w11975_,
		_w16781_
	);
	LUT3 #(
		.INIT('h80)
	) name6269 (
		\wishbone_bd_ram_mem2_reg[144][17]/P0001 ,
		_w11941_,
		_w11959_,
		_w16782_
	);
	LUT3 #(
		.INIT('h80)
	) name6270 (
		\wishbone_bd_ram_mem2_reg[47][17]/P0001 ,
		_w11957_,
		_w11973_,
		_w16783_
	);
	LUT3 #(
		.INIT('h80)
	) name6271 (
		\wishbone_bd_ram_mem2_reg[251][17]/P0001 ,
		_w11936_,
		_w11952_,
		_w16784_
	);
	LUT4 #(
		.INIT('h0001)
	) name6272 (
		_w16781_,
		_w16782_,
		_w16783_,
		_w16784_,
		_w16785_
	);
	LUT3 #(
		.INIT('h80)
	) name6273 (
		\wishbone_bd_ram_mem2_reg[113][17]/P0001 ,
		_w11977_,
		_w12012_,
		_w16786_
	);
	LUT3 #(
		.INIT('h80)
	) name6274 (
		\wishbone_bd_ram_mem2_reg[65][17]/P0001 ,
		_w11949_,
		_w11977_,
		_w16787_
	);
	LUT3 #(
		.INIT('h80)
	) name6275 (
		\wishbone_bd_ram_mem2_reg[180][17]/P0001 ,
		_w11929_,
		_w11942_,
		_w16788_
	);
	LUT3 #(
		.INIT('h80)
	) name6276 (
		\wishbone_bd_ram_mem2_reg[193][17]/P0001 ,
		_w11945_,
		_w11977_,
		_w16789_
	);
	LUT4 #(
		.INIT('h0001)
	) name6277 (
		_w16786_,
		_w16787_,
		_w16788_,
		_w16789_,
		_w16790_
	);
	LUT4 #(
		.INIT('h8000)
	) name6278 (
		_w16775_,
		_w16780_,
		_w16785_,
		_w16790_,
		_w16791_
	);
	LUT3 #(
		.INIT('h80)
	) name6279 (
		\wishbone_bd_ram_mem2_reg[41][17]/P0001 ,
		_w11957_,
		_w11968_,
		_w16792_
	);
	LUT3 #(
		.INIT('h80)
	) name6280 (
		\wishbone_bd_ram_mem2_reg[160][17]/P0001 ,
		_w11930_,
		_w11941_,
		_w16793_
	);
	LUT3 #(
		.INIT('h80)
	) name6281 (
		\wishbone_bd_ram_mem2_reg[217][17]/P0001 ,
		_w11968_,
		_w11984_,
		_w16794_
	);
	LUT3 #(
		.INIT('h80)
	) name6282 (
		\wishbone_bd_ram_mem2_reg[142][17]/P0001 ,
		_w11948_,
		_w11955_,
		_w16795_
	);
	LUT4 #(
		.INIT('h0001)
	) name6283 (
		_w16792_,
		_w16793_,
		_w16794_,
		_w16795_,
		_w16796_
	);
	LUT3 #(
		.INIT('h80)
	) name6284 (
		\wishbone_bd_ram_mem2_reg[78][17]/P0001 ,
		_w11948_,
		_w11949_,
		_w16797_
	);
	LUT3 #(
		.INIT('h80)
	) name6285 (
		\wishbone_bd_ram_mem2_reg[207][17]/P0001 ,
		_w11945_,
		_w11973_,
		_w16798_
	);
	LUT3 #(
		.INIT('h80)
	) name6286 (
		\wishbone_bd_ram_mem2_reg[128][17]/P0001 ,
		_w11941_,
		_w11955_,
		_w16799_
	);
	LUT3 #(
		.INIT('h80)
	) name6287 (
		\wishbone_bd_ram_mem2_reg[24][17]/P0001 ,
		_w11935_,
		_w11990_,
		_w16800_
	);
	LUT4 #(
		.INIT('h0001)
	) name6288 (
		_w16797_,
		_w16798_,
		_w16799_,
		_w16800_,
		_w16801_
	);
	LUT3 #(
		.INIT('h80)
	) name6289 (
		\wishbone_bd_ram_mem2_reg[127][17]/P0001 ,
		_w11973_,
		_w12012_,
		_w16802_
	);
	LUT3 #(
		.INIT('h80)
	) name6290 (
		\wishbone_bd_ram_mem2_reg[40][17]/P0001 ,
		_w11957_,
		_w11990_,
		_w16803_
	);
	LUT3 #(
		.INIT('h80)
	) name6291 (
		\wishbone_bd_ram_mem2_reg[151][17]/P0001 ,
		_w11959_,
		_w11975_,
		_w16804_
	);
	LUT3 #(
		.INIT('h80)
	) name6292 (
		\wishbone_bd_ram_mem2_reg[71][17]/P0001 ,
		_w11949_,
		_w11975_,
		_w16805_
	);
	LUT4 #(
		.INIT('h0001)
	) name6293 (
		_w16802_,
		_w16803_,
		_w16804_,
		_w16805_,
		_w16806_
	);
	LUT3 #(
		.INIT('h80)
	) name6294 (
		\wishbone_bd_ram_mem2_reg[32][17]/P0001 ,
		_w11941_,
		_w11957_,
		_w16807_
	);
	LUT3 #(
		.INIT('h80)
	) name6295 (
		\wishbone_bd_ram_mem2_reg[50][17]/P0001 ,
		_w11963_,
		_w11979_,
		_w16808_
	);
	LUT3 #(
		.INIT('h80)
	) name6296 (
		\wishbone_bd_ram_mem2_reg[148][17]/P0001 ,
		_w11929_,
		_w11959_,
		_w16809_
	);
	LUT3 #(
		.INIT('h80)
	) name6297 (
		\wishbone_bd_ram_mem2_reg[237][17]/P0001 ,
		_w11966_,
		_w11982_,
		_w16810_
	);
	LUT4 #(
		.INIT('h0001)
	) name6298 (
		_w16807_,
		_w16808_,
		_w16809_,
		_w16810_,
		_w16811_
	);
	LUT4 #(
		.INIT('h8000)
	) name6299 (
		_w16796_,
		_w16801_,
		_w16806_,
		_w16811_,
		_w16812_
	);
	LUT4 #(
		.INIT('h8000)
	) name6300 (
		_w16749_,
		_w16770_,
		_w16791_,
		_w16812_,
		_w16813_
	);
	LUT4 #(
		.INIT('h8000)
	) name6301 (
		_w16558_,
		_w16643_,
		_w16728_,
		_w16813_,
		_w16814_
	);
	LUT4 #(
		.INIT('h936c)
	) name6302 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w16815_
	);
	LUT3 #(
		.INIT('h40)
	) name6303 (
		_w12302_,
		_w12304_,
		_w16815_,
		_w16816_
	);
	LUT3 #(
		.INIT('h70)
	) name6304 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		_w16817_
	);
	LUT2 #(
		.INIT('h4)
	) name6305 (
		_w12302_,
		_w16817_,
		_w16818_
	);
	LUT4 #(
		.INIT('h008f)
	) name6306 (
		_w12312_,
		_w12317_,
		_w16816_,
		_w16818_,
		_w16819_
	);
	LUT3 #(
		.INIT('h2f)
	) name6307 (
		_w12303_,
		_w16814_,
		_w16819_,
		_w16820_
	);
	LUT4 #(
		.INIT('h1333)
	) name6308 (
		\txethmac1_txcounters1_ByteCnt_reg[10]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[11]/NET0131 ,
		_w13034_,
		_w13036_,
		_w16821_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6309 (
		_w13027_,
		_w13034_,
		_w13036_,
		_w13040_,
		_w16822_
	);
	LUT2 #(
		.INIT('h4)
	) name6310 (
		_w16821_,
		_w16822_,
		_w16823_
	);
	LUT2 #(
		.INIT('h1)
	) name6311 (
		\txethmac1_txcrc_Crc_reg[5]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w16824_
	);
	LUT3 #(
		.INIT('h60)
	) name6312 (
		_w11105_,
		_w11106_,
		_w16824_,
		_w16825_
	);
	LUT3 #(
		.INIT('h40)
	) name6313 (
		\txethmac1_txcrc_Crc_reg[5]/NET0131 ,
		_w10913_,
		_w10914_,
		_w16826_
	);
	LUT4 #(
		.INIT('h090f)
	) name6314 (
		_w11105_,
		_w11106_,
		_w16826_,
		_w11110_,
		_w16827_
	);
	LUT2 #(
		.INIT('he)
	) name6315 (
		_w16825_,
		_w16827_,
		_w16828_
	);
	LUT4 #(
		.INIT('h0001)
	) name6316 (
		\wishbone_RxPointerMSB_reg[12]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w16829_
	);
	LUT3 #(
		.INIT('h07)
	) name6317 (
		_w11868_,
		_w11875_,
		_w16829_,
		_w16830_
	);
	LUT3 #(
		.INIT('h80)
	) name6318 (
		_w11870_,
		_w11873_,
		_w16830_,
		_w16831_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name6319 (
		\m_wb_adr_o[12]_pad ,
		_w11845_,
		_w11846_,
		_w11848_,
		_w16832_
	);
	LUT3 #(
		.INIT('he0)
	) name6320 (
		_w11887_,
		_w16831_,
		_w16832_,
		_w16833_
	);
	LUT4 #(
		.INIT('h080a)
	) name6321 (
		\wishbone_RxPointerMSB_reg[12]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16834_
	);
	LUT3 #(
		.INIT('he0)
	) name6322 (
		_w11902_,
		_w11905_,
		_w16834_,
		_w16835_
	);
	LUT3 #(
		.INIT('ha2)
	) name6323 (
		\wishbone_TxPointerMSB_reg[12]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16836_
	);
	LUT4 #(
		.INIT('h0007)
	) name6324 (
		\m_wb_adr_o[12]_pad ,
		_w11907_,
		_w16835_,
		_w16836_,
		_w16837_
	);
	LUT2 #(
		.INIT('hb)
	) name6325 (
		_w16833_,
		_w16837_,
		_w16838_
	);
	LUT4 #(
		.INIT('h0001)
	) name6326 (
		\wishbone_TxPointerMSB_reg[16]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w16839_
	);
	LUT4 #(
		.INIT('h008f)
	) name6327 (
		_w11866_,
		_w11867_,
		_w11883_,
		_w16839_,
		_w16840_
	);
	LUT2 #(
		.INIT('h4)
	) name6328 (
		_w11882_,
		_w16840_,
		_w16841_
	);
	LUT2 #(
		.INIT('h6)
	) name6329 (
		\m_wb_adr_o[16]_pad ,
		_w11851_,
		_w16842_
	);
	LUT3 #(
		.INIT('he0)
	) name6330 (
		_w13051_,
		_w16841_,
		_w16842_,
		_w16843_
	);
	LUT3 #(
		.INIT('ha2)
	) name6331 (
		\wishbone_TxPointerMSB_reg[16]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16844_
	);
	LUT4 #(
		.INIT('h080a)
	) name6332 (
		\wishbone_RxPointerMSB_reg[16]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16845_
	);
	LUT3 #(
		.INIT('he0)
	) name6333 (
		_w11902_,
		_w11905_,
		_w16845_,
		_w16846_
	);
	LUT4 #(
		.INIT('h0007)
	) name6334 (
		\m_wb_adr_o[16]_pad ,
		_w11907_,
		_w16844_,
		_w16846_,
		_w16847_
	);
	LUT2 #(
		.INIT('hb)
	) name6335 (
		_w16843_,
		_w16847_,
		_w16848_
	);
	LUT3 #(
		.INIT('h13)
	) name6336 (
		\m_wb_adr_o[16]_pad ,
		\m_wb_adr_o[17]_pad ,
		_w11851_,
		_w16849_
	);
	LUT4 #(
		.INIT('h0001)
	) name6337 (
		\wishbone_TxPointerMSB_reg[17]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w16850_
	);
	LUT4 #(
		.INIT('h008f)
	) name6338 (
		_w11866_,
		_w11867_,
		_w11883_,
		_w16850_,
		_w16851_
	);
	LUT2 #(
		.INIT('h4)
	) name6339 (
		_w11882_,
		_w16851_,
		_w16852_
	);
	LUT4 #(
		.INIT('h0302)
	) name6340 (
		_w13051_,
		_w14162_,
		_w16849_,
		_w16852_,
		_w16853_
	);
	LUT3 #(
		.INIT('ha2)
	) name6341 (
		\wishbone_TxPointerMSB_reg[17]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16854_
	);
	LUT4 #(
		.INIT('h080a)
	) name6342 (
		\wishbone_RxPointerMSB_reg[17]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16855_
	);
	LUT3 #(
		.INIT('he0)
	) name6343 (
		_w11902_,
		_w11905_,
		_w16855_,
		_w16856_
	);
	LUT4 #(
		.INIT('h0007)
	) name6344 (
		\m_wb_adr_o[17]_pad ,
		_w11907_,
		_w16854_,
		_w16856_,
		_w16857_
	);
	LUT2 #(
		.INIT('hb)
	) name6345 (
		_w16853_,
		_w16857_,
		_w16858_
	);
	LUT3 #(
		.INIT('h15)
	) name6346 (
		\m_wb_adr_o[19]_pad ,
		_w11851_,
		_w14164_,
		_w16859_
	);
	LUT4 #(
		.INIT('h0001)
	) name6347 (
		\wishbone_TxPointerMSB_reg[19]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w16860_
	);
	LUT4 #(
		.INIT('h008f)
	) name6348 (
		_w11866_,
		_w11867_,
		_w11883_,
		_w16860_,
		_w16861_
	);
	LUT2 #(
		.INIT('h4)
	) name6349 (
		_w11882_,
		_w16861_,
		_w16862_
	);
	LUT4 #(
		.INIT('h0504)
	) name6350 (
		_w11853_,
		_w13051_,
		_w16859_,
		_w16862_,
		_w16863_
	);
	LUT3 #(
		.INIT('ha2)
	) name6351 (
		\wishbone_TxPointerMSB_reg[19]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16864_
	);
	LUT4 #(
		.INIT('h080a)
	) name6352 (
		\wishbone_RxPointerMSB_reg[19]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16865_
	);
	LUT3 #(
		.INIT('he0)
	) name6353 (
		_w11902_,
		_w11905_,
		_w16865_,
		_w16866_
	);
	LUT4 #(
		.INIT('h0007)
	) name6354 (
		\m_wb_adr_o[19]_pad ,
		_w11907_,
		_w16864_,
		_w16866_,
		_w16867_
	);
	LUT2 #(
		.INIT('hb)
	) name6355 (
		_w16863_,
		_w16867_,
		_w16868_
	);
	LUT4 #(
		.INIT('h0001)
	) name6356 (
		\wishbone_RxPointerMSB_reg[20]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w16869_
	);
	LUT3 #(
		.INIT('h07)
	) name6357 (
		_w11868_,
		_w11875_,
		_w16869_,
		_w16870_
	);
	LUT3 #(
		.INIT('h80)
	) name6358 (
		_w11870_,
		_w11873_,
		_w16870_,
		_w16871_
	);
	LUT4 #(
		.INIT('h6660)
	) name6359 (
		\m_wb_adr_o[20]_pad ,
		_w11853_,
		_w11887_,
		_w16871_,
		_w16872_
	);
	LUT3 #(
		.INIT('ha2)
	) name6360 (
		\wishbone_TxPointerMSB_reg[20]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16873_
	);
	LUT4 #(
		.INIT('h080a)
	) name6361 (
		\wishbone_RxPointerMSB_reg[20]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16874_
	);
	LUT3 #(
		.INIT('he0)
	) name6362 (
		_w11902_,
		_w11905_,
		_w16874_,
		_w16875_
	);
	LUT4 #(
		.INIT('h0007)
	) name6363 (
		\m_wb_adr_o[20]_pad ,
		_w11907_,
		_w16873_,
		_w16875_,
		_w16876_
	);
	LUT2 #(
		.INIT('hb)
	) name6364 (
		_w16872_,
		_w16876_,
		_w16877_
	);
	LUT4 #(
		.INIT('h1333)
	) name6365 (
		\m_wb_adr_o[20]_pad ,
		\m_wb_adr_o[21]_pad ,
		_w11851_,
		_w11852_,
		_w16878_
	);
	LUT3 #(
		.INIT('h80)
	) name6366 (
		_w11851_,
		_w11852_,
		_w11854_,
		_w16879_
	);
	LUT4 #(
		.INIT('h0001)
	) name6367 (
		\wishbone_TxPointerMSB_reg[21]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w16880_
	);
	LUT4 #(
		.INIT('h008f)
	) name6368 (
		_w11866_,
		_w11867_,
		_w11883_,
		_w16880_,
		_w16881_
	);
	LUT2 #(
		.INIT('h4)
	) name6369 (
		_w11882_,
		_w16881_,
		_w16882_
	);
	LUT4 #(
		.INIT('h0302)
	) name6370 (
		_w13051_,
		_w16878_,
		_w16879_,
		_w16882_,
		_w16883_
	);
	LUT3 #(
		.INIT('ha2)
	) name6371 (
		\wishbone_TxPointerMSB_reg[21]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16884_
	);
	LUT4 #(
		.INIT('h080a)
	) name6372 (
		\wishbone_RxPointerMSB_reg[21]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16885_
	);
	LUT3 #(
		.INIT('he0)
	) name6373 (
		_w11902_,
		_w11905_,
		_w16885_,
		_w16886_
	);
	LUT4 #(
		.INIT('h0007)
	) name6374 (
		\m_wb_adr_o[21]_pad ,
		_w11907_,
		_w16884_,
		_w16886_,
		_w16887_
	);
	LUT2 #(
		.INIT('hb)
	) name6375 (
		_w16883_,
		_w16887_,
		_w16888_
	);
	LUT4 #(
		.INIT('h080a)
	) name6376 (
		\wishbone_RxPointerMSB_reg[3]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16889_
	);
	LUT3 #(
		.INIT('he0)
	) name6377 (
		_w11902_,
		_w11905_,
		_w16889_,
		_w16890_
	);
	LUT3 #(
		.INIT('h07)
	) name6378 (
		\m_wb_adr_o[3]_pad ,
		_w11907_,
		_w16890_,
		_w16891_
	);
	LUT3 #(
		.INIT('ha2)
	) name6379 (
		\wishbone_TxPointerMSB_reg[3]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16892_
	);
	LUT2 #(
		.INIT('h6)
	) name6380 (
		\m_wb_adr_o[2]_pad ,
		\m_wb_adr_o[3]_pad ,
		_w16893_
	);
	LUT3 #(
		.INIT('he0)
	) name6381 (
		_w11887_,
		_w13051_,
		_w16893_,
		_w16894_
	);
	LUT2 #(
		.INIT('h1)
	) name6382 (
		_w16892_,
		_w16894_,
		_w16895_
	);
	LUT2 #(
		.INIT('h7)
	) name6383 (
		_w16891_,
		_w16895_,
		_w16896_
	);
	LUT4 #(
		.INIT('h1555)
	) name6384 (
		\m_wb_adr_o[22]_pad ,
		_w11851_,
		_w11852_,
		_w11854_,
		_w16897_
	);
	LUT4 #(
		.INIT('h0001)
	) name6385 (
		\wishbone_TxPointerMSB_reg[22]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w16898_
	);
	LUT4 #(
		.INIT('h008f)
	) name6386 (
		_w11866_,
		_w11867_,
		_w11883_,
		_w16898_,
		_w16899_
	);
	LUT2 #(
		.INIT('h4)
	) name6387 (
		_w11882_,
		_w16899_,
		_w16900_
	);
	LUT3 #(
		.INIT('h80)
	) name6388 (
		\m_wb_adr_o[20]_pad ,
		\m_wb_adr_o[21]_pad ,
		\m_wb_adr_o[22]_pad ,
		_w16901_
	);
	LUT3 #(
		.INIT('h80)
	) name6389 (
		_w11851_,
		_w11852_,
		_w16901_,
		_w16902_
	);
	LUT4 #(
		.INIT('h0032)
	) name6390 (
		_w13051_,
		_w16897_,
		_w16900_,
		_w16902_,
		_w16903_
	);
	LUT3 #(
		.INIT('ha2)
	) name6391 (
		\wishbone_TxPointerMSB_reg[22]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16904_
	);
	LUT4 #(
		.INIT('h080a)
	) name6392 (
		\wishbone_RxPointerMSB_reg[22]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16905_
	);
	LUT3 #(
		.INIT('he0)
	) name6393 (
		_w11902_,
		_w11905_,
		_w16905_,
		_w16906_
	);
	LUT4 #(
		.INIT('h0007)
	) name6394 (
		\m_wb_adr_o[22]_pad ,
		_w11907_,
		_w16904_,
		_w16906_,
		_w16907_
	);
	LUT2 #(
		.INIT('hb)
	) name6395 (
		_w16903_,
		_w16907_,
		_w16908_
	);
	LUT4 #(
		.INIT('h8000)
	) name6396 (
		\m_wb_adr_o[23]_pad ,
		_w11851_,
		_w11852_,
		_w16901_,
		_w16909_
	);
	LUT4 #(
		.INIT('h54a8)
	) name6397 (
		\m_wb_adr_o[23]_pad ,
		_w11887_,
		_w13051_,
		_w16902_,
		_w16910_
	);
	LUT4 #(
		.INIT('h080a)
	) name6398 (
		\wishbone_RxPointerMSB_reg[23]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16911_
	);
	LUT3 #(
		.INIT('he0)
	) name6399 (
		_w11902_,
		_w11905_,
		_w16911_,
		_w16912_
	);
	LUT3 #(
		.INIT('ha2)
	) name6400 (
		\wishbone_TxPointerMSB_reg[23]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16913_
	);
	LUT4 #(
		.INIT('h0007)
	) name6401 (
		\m_wb_adr_o[23]_pad ,
		_w11907_,
		_w16912_,
		_w16913_,
		_w16914_
	);
	LUT2 #(
		.INIT('hb)
	) name6402 (
		_w16910_,
		_w16914_,
		_w16915_
	);
	LUT2 #(
		.INIT('h1)
	) name6403 (
		\m_wb_adr_o[24]_pad ,
		_w16909_,
		_w16916_
	);
	LUT4 #(
		.INIT('h0001)
	) name6404 (
		\wishbone_RxPointerMSB_reg[24]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w16917_
	);
	LUT3 #(
		.INIT('h07)
	) name6405 (
		_w11868_,
		_w11875_,
		_w16917_,
		_w16918_
	);
	LUT3 #(
		.INIT('h80)
	) name6406 (
		_w11870_,
		_w11873_,
		_w16918_,
		_w16919_
	);
	LUT3 #(
		.INIT('h32)
	) name6407 (
		_w11887_,
		_w13407_,
		_w16919_,
		_w16920_
	);
	LUT2 #(
		.INIT('h4)
	) name6408 (
		_w16916_,
		_w16920_,
		_w16921_
	);
	LUT3 #(
		.INIT('ha2)
	) name6409 (
		\wishbone_TxPointerMSB_reg[24]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16922_
	);
	LUT4 #(
		.INIT('h080a)
	) name6410 (
		\wishbone_RxPointerMSB_reg[24]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16923_
	);
	LUT3 #(
		.INIT('he0)
	) name6411 (
		_w11902_,
		_w11905_,
		_w16923_,
		_w16924_
	);
	LUT4 #(
		.INIT('h0007)
	) name6412 (
		\m_wb_adr_o[24]_pad ,
		_w11907_,
		_w16922_,
		_w16924_,
		_w16925_
	);
	LUT2 #(
		.INIT('hb)
	) name6413 (
		_w16921_,
		_w16925_,
		_w16926_
	);
	LUT4 #(
		.INIT('h5554)
	) name6414 (
		\m_wb_adr_o[25]_pad ,
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w16927_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6415 (
		_w11851_,
		_w11852_,
		_w13406_,
		_w16927_,
		_w16928_
	);
	LUT4 #(
		.INIT('haaa8)
	) name6416 (
		\m_wb_adr_o[25]_pad ,
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w16929_
	);
	LUT4 #(
		.INIT('h8000)
	) name6417 (
		_w11851_,
		_w11852_,
		_w13406_,
		_w16929_,
		_w16930_
	);
	LUT4 #(
		.INIT('h0001)
	) name6418 (
		\wishbone_RxPointerMSB_reg[25]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w16931_
	);
	LUT3 #(
		.INIT('h07)
	) name6419 (
		_w11868_,
		_w11875_,
		_w16931_,
		_w16932_
	);
	LUT3 #(
		.INIT('h80)
	) name6420 (
		_w11870_,
		_w11873_,
		_w16932_,
		_w16933_
	);
	LUT3 #(
		.INIT('h10)
	) name6421 (
		_w16928_,
		_w16930_,
		_w16933_,
		_w16934_
	);
	LUT4 #(
		.INIT('h5554)
	) name6422 (
		\m_wb_adr_o[25]_pad ,
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w16935_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6423 (
		_w11851_,
		_w11852_,
		_w13406_,
		_w16935_,
		_w16936_
	);
	LUT4 #(
		.INIT('haaa8)
	) name6424 (
		\m_wb_adr_o[25]_pad ,
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w16937_
	);
	LUT4 #(
		.INIT('h8000)
	) name6425 (
		_w11851_,
		_w11852_,
		_w13406_,
		_w16937_,
		_w16938_
	);
	LUT4 #(
		.INIT('h0001)
	) name6426 (
		\wishbone_TxPointerMSB_reg[25]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w16939_
	);
	LUT4 #(
		.INIT('h008f)
	) name6427 (
		_w11866_,
		_w11867_,
		_w11883_,
		_w16939_,
		_w16940_
	);
	LUT2 #(
		.INIT('h4)
	) name6428 (
		_w11882_,
		_w16940_,
		_w16941_
	);
	LUT3 #(
		.INIT('h10)
	) name6429 (
		_w16936_,
		_w16938_,
		_w16941_,
		_w16942_
	);
	LUT4 #(
		.INIT('h0222)
	) name6430 (
		\wishbone_RxPointerMSB_reg[25]/NET0131 ,
		\wishbone_rx_burst_en_reg/NET0131 ,
		_w11866_,
		_w11867_,
		_w16943_
	);
	LUT3 #(
		.INIT('he0)
	) name6431 (
		_w11894_,
		_w11904_,
		_w16943_,
		_w16944_
	);
	LUT3 #(
		.INIT('h0d)
	) name6432 (
		\wishbone_TxPointerMSB_reg[25]/NET0131 ,
		_w11900_,
		_w16944_,
		_w16945_
	);
	LUT4 #(
		.INIT('h0700)
	) name6433 (
		\m_wb_adr_o[25]_pad ,
		_w11907_,
		_w16942_,
		_w16945_,
		_w16946_
	);
	LUT2 #(
		.INIT('hb)
	) name6434 (
		_w16934_,
		_w16946_,
		_w16947_
	);
	LUT2 #(
		.INIT('h1)
	) name6435 (
		\m_wb_adr_o[28]_pad ,
		_w15404_,
		_w16948_
	);
	LUT4 #(
		.INIT('h8000)
	) name6436 (
		_w11851_,
		_w11852_,
		_w11857_,
		_w11859_,
		_w16949_
	);
	LUT4 #(
		.INIT('h0001)
	) name6437 (
		\wishbone_RxPointerMSB_reg[28]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w16950_
	);
	LUT3 #(
		.INIT('h07)
	) name6438 (
		_w11868_,
		_w11875_,
		_w16950_,
		_w16951_
	);
	LUT3 #(
		.INIT('h80)
	) name6439 (
		_w11870_,
		_w11873_,
		_w16951_,
		_w16952_
	);
	LUT3 #(
		.INIT('h32)
	) name6440 (
		_w11887_,
		_w16949_,
		_w16952_,
		_w16953_
	);
	LUT2 #(
		.INIT('h4)
	) name6441 (
		_w16948_,
		_w16953_,
		_w16954_
	);
	LUT3 #(
		.INIT('ha2)
	) name6442 (
		\wishbone_TxPointerMSB_reg[28]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16955_
	);
	LUT4 #(
		.INIT('h080a)
	) name6443 (
		\wishbone_RxPointerMSB_reg[28]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16956_
	);
	LUT3 #(
		.INIT('he0)
	) name6444 (
		_w11902_,
		_w11905_,
		_w16956_,
		_w16957_
	);
	LUT4 #(
		.INIT('h0007)
	) name6445 (
		\m_wb_adr_o[28]_pad ,
		_w11907_,
		_w16955_,
		_w16957_,
		_w16958_
	);
	LUT2 #(
		.INIT('hb)
	) name6446 (
		_w16954_,
		_w16958_,
		_w16959_
	);
	LUT2 #(
		.INIT('h1)
	) name6447 (
		\m_wb_adr_o[29]_pad ,
		_w16949_,
		_w16960_
	);
	LUT4 #(
		.INIT('h0001)
	) name6448 (
		\wishbone_RxPointerMSB_reg[29]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w16961_
	);
	LUT3 #(
		.INIT('h07)
	) name6449 (
		_w11868_,
		_w11875_,
		_w16961_,
		_w16962_
	);
	LUT3 #(
		.INIT('h80)
	) name6450 (
		_w11870_,
		_w11873_,
		_w16962_,
		_w16963_
	);
	LUT3 #(
		.INIT('h54)
	) name6451 (
		_w11861_,
		_w11887_,
		_w16963_,
		_w16964_
	);
	LUT2 #(
		.INIT('h4)
	) name6452 (
		_w16960_,
		_w16964_,
		_w16965_
	);
	LUT4 #(
		.INIT('h080a)
	) name6453 (
		\wishbone_RxPointerMSB_reg[29]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16966_
	);
	LUT3 #(
		.INIT('he0)
	) name6454 (
		_w11902_,
		_w11905_,
		_w16966_,
		_w16967_
	);
	LUT3 #(
		.INIT('ha2)
	) name6455 (
		\wishbone_TxPointerMSB_reg[29]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16968_
	);
	LUT4 #(
		.INIT('h0007)
	) name6456 (
		\m_wb_adr_o[29]_pad ,
		_w11907_,
		_w16967_,
		_w16968_,
		_w16969_
	);
	LUT2 #(
		.INIT('hb)
	) name6457 (
		_w16965_,
		_w16969_,
		_w16970_
	);
	LUT4 #(
		.INIT('h080a)
	) name6458 (
		\wishbone_RxPointerMSB_reg[5]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16971_
	);
	LUT3 #(
		.INIT('he0)
	) name6459 (
		_w11902_,
		_w11905_,
		_w16971_,
		_w16972_
	);
	LUT3 #(
		.INIT('h07)
	) name6460 (
		\m_wb_adr_o[5]_pad ,
		_w11907_,
		_w16972_,
		_w16973_
	);
	LUT3 #(
		.INIT('ha2)
	) name6461 (
		\wishbone_TxPointerMSB_reg[5]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16974_
	);
	LUT4 #(
		.INIT('h7f80)
	) name6462 (
		\m_wb_adr_o[2]_pad ,
		\m_wb_adr_o[3]_pad ,
		\m_wb_adr_o[4]_pad ,
		\m_wb_adr_o[5]_pad ,
		_w16975_
	);
	LUT3 #(
		.INIT('he0)
	) name6463 (
		_w11887_,
		_w13051_,
		_w16975_,
		_w16976_
	);
	LUT2 #(
		.INIT('h1)
	) name6464 (
		_w16974_,
		_w16976_,
		_w16977_
	);
	LUT2 #(
		.INIT('h7)
	) name6465 (
		_w16973_,
		_w16977_,
		_w16978_
	);
	LUT4 #(
		.INIT('h080a)
	) name6466 (
		\wishbone_RxPointerMSB_reg[6]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16979_
	);
	LUT3 #(
		.INIT('he0)
	) name6467 (
		_w11902_,
		_w11905_,
		_w16979_,
		_w16980_
	);
	LUT3 #(
		.INIT('h07)
	) name6468 (
		\m_wb_adr_o[6]_pad ,
		_w11907_,
		_w16980_,
		_w16981_
	);
	LUT3 #(
		.INIT('ha2)
	) name6469 (
		\wishbone_TxPointerMSB_reg[6]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16982_
	);
	LUT2 #(
		.INIT('h6)
	) name6470 (
		\m_wb_adr_o[6]_pad ,
		_w11845_,
		_w16983_
	);
	LUT3 #(
		.INIT('he0)
	) name6471 (
		_w11887_,
		_w13051_,
		_w16983_,
		_w16984_
	);
	LUT2 #(
		.INIT('h1)
	) name6472 (
		_w16982_,
		_w16984_,
		_w16985_
	);
	LUT2 #(
		.INIT('h7)
	) name6473 (
		_w16981_,
		_w16985_,
		_w16986_
	);
	LUT4 #(
		.INIT('h080a)
	) name6474 (
		\wishbone_RxPointerMSB_reg[7]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16987_
	);
	LUT3 #(
		.INIT('he0)
	) name6475 (
		_w11902_,
		_w11905_,
		_w16987_,
		_w16988_
	);
	LUT3 #(
		.INIT('h07)
	) name6476 (
		\m_wb_adr_o[7]_pad ,
		_w11907_,
		_w16988_,
		_w16989_
	);
	LUT3 #(
		.INIT('ha2)
	) name6477 (
		\wishbone_TxPointerMSB_reg[7]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16990_
	);
	LUT3 #(
		.INIT('h6c)
	) name6478 (
		\m_wb_adr_o[6]_pad ,
		\m_wb_adr_o[7]_pad ,
		_w11845_,
		_w16991_
	);
	LUT3 #(
		.INIT('he0)
	) name6479 (
		_w11887_,
		_w13051_,
		_w16991_,
		_w16992_
	);
	LUT2 #(
		.INIT('h1)
	) name6480 (
		_w16990_,
		_w16992_,
		_w16993_
	);
	LUT2 #(
		.INIT('h7)
	) name6481 (
		_w16989_,
		_w16993_,
		_w16994_
	);
	LUT3 #(
		.INIT('ha2)
	) name6482 (
		\wishbone_TxPointerMSB_reg[9]/NET0131 ,
		_w11900_,
		_w11909_,
		_w16995_
	);
	LUT4 #(
		.INIT('h080a)
	) name6483 (
		\wishbone_RxPointerMSB_reg[9]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w16996_
	);
	LUT3 #(
		.INIT('he0)
	) name6484 (
		_w11902_,
		_w11905_,
		_w16996_,
		_w16997_
	);
	LUT2 #(
		.INIT('h1)
	) name6485 (
		_w16995_,
		_w16997_,
		_w16998_
	);
	LUT3 #(
		.INIT('h6a)
	) name6486 (
		\m_wb_adr_o[9]_pad ,
		_w11845_,
		_w11846_,
		_w16999_
	);
	LUT3 #(
		.INIT('he0)
	) name6487 (
		_w11887_,
		_w13051_,
		_w16999_,
		_w17000_
	);
	LUT3 #(
		.INIT('h07)
	) name6488 (
		\m_wb_adr_o[9]_pad ,
		_w11907_,
		_w17000_,
		_w17001_
	);
	LUT2 #(
		.INIT('h7)
	) name6489 (
		_w16998_,
		_w17001_,
		_w17002_
	);
	LUT3 #(
		.INIT('ha2)
	) name6490 (
		\wishbone_TxPointerMSB_reg[10]/NET0131 ,
		_w11900_,
		_w11909_,
		_w17003_
	);
	LUT4 #(
		.INIT('h080a)
	) name6491 (
		\wishbone_RxPointerMSB_reg[10]/NET0131 ,
		_w11904_,
		_w11912_,
		_w11913_,
		_w17004_
	);
	LUT3 #(
		.INIT('he0)
	) name6492 (
		_w11902_,
		_w11905_,
		_w17004_,
		_w17005_
	);
	LUT2 #(
		.INIT('h1)
	) name6493 (
		_w17003_,
		_w17005_,
		_w17006_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name6494 (
		\m_wb_adr_o[10]_pad ,
		\m_wb_adr_o[9]_pad ,
		_w11845_,
		_w11846_,
		_w17007_
	);
	LUT3 #(
		.INIT('he0)
	) name6495 (
		_w11887_,
		_w13051_,
		_w17007_,
		_w17008_
	);
	LUT3 #(
		.INIT('h07)
	) name6496 (
		\m_wb_adr_o[10]_pad ,
		_w11907_,
		_w17008_,
		_w17009_
	);
	LUT2 #(
		.INIT('h7)
	) name6497 (
		_w17006_,
		_w17009_,
		_w17010_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6498 (
		\wishbone_LatchedTxLength_reg[0]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w17011_
	);
	LUT3 #(
		.INIT('hf2)
	) name6499 (
		_w12303_,
		_w16122_,
		_w17011_,
		_w17012_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6500 (
		\wishbone_LatchedTxLength_reg[10]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w17013_
	);
	LUT3 #(
		.INIT('hf2)
	) name6501 (
		_w12303_,
		_w14872_,
		_w17013_,
		_w17014_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6502 (
		\wishbone_LatchedTxLength_reg[11]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w17015_
	);
	LUT3 #(
		.INIT('h80)
	) name6503 (
		\wishbone_bd_ram_mem3_reg[80][27]/P0001 ,
		_w11941_,
		_w11972_,
		_w17016_
	);
	LUT3 #(
		.INIT('h80)
	) name6504 (
		\wishbone_bd_ram_mem3_reg[3][27]/P0001 ,
		_w11932_,
		_w11938_,
		_w17017_
	);
	LUT3 #(
		.INIT('h80)
	) name6505 (
		\wishbone_bd_ram_mem3_reg[52][27]/P0001 ,
		_w11929_,
		_w11979_,
		_w17018_
	);
	LUT3 #(
		.INIT('h80)
	) name6506 (
		\wishbone_bd_ram_mem3_reg[73][27]/P0001 ,
		_w11949_,
		_w11968_,
		_w17019_
	);
	LUT4 #(
		.INIT('h0001)
	) name6507 (
		_w17016_,
		_w17017_,
		_w17018_,
		_w17019_,
		_w17020_
	);
	LUT3 #(
		.INIT('h80)
	) name6508 (
		\wishbone_bd_ram_mem3_reg[124][27]/P0001 ,
		_w11954_,
		_w12012_,
		_w17021_
	);
	LUT3 #(
		.INIT('h80)
	) name6509 (
		\wishbone_bd_ram_mem3_reg[169][27]/P0001 ,
		_w11930_,
		_w11968_,
		_w17022_
	);
	LUT3 #(
		.INIT('h80)
	) name6510 (
		\wishbone_bd_ram_mem3_reg[128][27]/P0001 ,
		_w11941_,
		_w11955_,
		_w17023_
	);
	LUT3 #(
		.INIT('h80)
	) name6511 (
		\wishbone_bd_ram_mem3_reg[200][27]/P0001 ,
		_w11945_,
		_w11990_,
		_w17024_
	);
	LUT4 #(
		.INIT('h0001)
	) name6512 (
		_w17021_,
		_w17022_,
		_w17023_,
		_w17024_,
		_w17025_
	);
	LUT3 #(
		.INIT('h80)
	) name6513 (
		\wishbone_bd_ram_mem3_reg[214][27]/P0001 ,
		_w11984_,
		_w11986_,
		_w17026_
	);
	LUT3 #(
		.INIT('h80)
	) name6514 (
		\wishbone_bd_ram_mem3_reg[113][27]/P0001 ,
		_w11977_,
		_w12012_,
		_w17027_
	);
	LUT3 #(
		.INIT('h80)
	) name6515 (
		\wishbone_bd_ram_mem3_reg[119][27]/P0001 ,
		_w11975_,
		_w12012_,
		_w17028_
	);
	LUT3 #(
		.INIT('h80)
	) name6516 (
		\wishbone_bd_ram_mem3_reg[132][27]/P0001 ,
		_w11929_,
		_w11955_,
		_w17029_
	);
	LUT4 #(
		.INIT('h0001)
	) name6517 (
		_w17026_,
		_w17027_,
		_w17028_,
		_w17029_,
		_w17030_
	);
	LUT3 #(
		.INIT('h80)
	) name6518 (
		\wishbone_bd_ram_mem3_reg[55][27]/P0001 ,
		_w11975_,
		_w11979_,
		_w17031_
	);
	LUT3 #(
		.INIT('h80)
	) name6519 (
		\wishbone_bd_ram_mem3_reg[219][27]/P0001 ,
		_w11936_,
		_w11984_,
		_w17032_
	);
	LUT3 #(
		.INIT('h80)
	) name6520 (
		\wishbone_bd_ram_mem3_reg[147][27]/P0001 ,
		_w11938_,
		_w11959_,
		_w17033_
	);
	LUT3 #(
		.INIT('h80)
	) name6521 (
		\wishbone_bd_ram_mem3_reg[180][27]/P0001 ,
		_w11929_,
		_w11942_,
		_w17034_
	);
	LUT4 #(
		.INIT('h0001)
	) name6522 (
		_w17031_,
		_w17032_,
		_w17033_,
		_w17034_,
		_w17035_
	);
	LUT4 #(
		.INIT('h8000)
	) name6523 (
		_w17020_,
		_w17025_,
		_w17030_,
		_w17035_,
		_w17036_
	);
	LUT3 #(
		.INIT('h80)
	) name6524 (
		\wishbone_bd_ram_mem3_reg[120][27]/P0001 ,
		_w11990_,
		_w12012_,
		_w17037_
	);
	LUT3 #(
		.INIT('h80)
	) name6525 (
		\wishbone_bd_ram_mem3_reg[177][27]/P0001 ,
		_w11942_,
		_w11977_,
		_w17038_
	);
	LUT3 #(
		.INIT('h80)
	) name6526 (
		\wishbone_bd_ram_mem3_reg[68][27]/P0001 ,
		_w11929_,
		_w11949_,
		_w17039_
	);
	LUT3 #(
		.INIT('h80)
	) name6527 (
		\wishbone_bd_ram_mem3_reg[136][27]/P0001 ,
		_w11955_,
		_w11990_,
		_w17040_
	);
	LUT4 #(
		.INIT('h0001)
	) name6528 (
		_w17037_,
		_w17038_,
		_w17039_,
		_w17040_,
		_w17041_
	);
	LUT3 #(
		.INIT('h80)
	) name6529 (
		\wishbone_bd_ram_mem3_reg[225][27]/P0001 ,
		_w11977_,
		_w11982_,
		_w17042_
	);
	LUT3 #(
		.INIT('h80)
	) name6530 (
		\wishbone_bd_ram_mem3_reg[242][27]/P0001 ,
		_w11952_,
		_w11963_,
		_w17043_
	);
	LUT3 #(
		.INIT('h80)
	) name6531 (
		\wishbone_bd_ram_mem3_reg[74][27]/P0001 ,
		_w11944_,
		_w11949_,
		_w17044_
	);
	LUT3 #(
		.INIT('h80)
	) name6532 (
		\wishbone_bd_ram_mem3_reg[37][27]/P0001 ,
		_w11933_,
		_w11957_,
		_w17045_
	);
	LUT4 #(
		.INIT('h0001)
	) name6533 (
		_w17042_,
		_w17043_,
		_w17044_,
		_w17045_,
		_w17046_
	);
	LUT3 #(
		.INIT('h80)
	) name6534 (
		\wishbone_bd_ram_mem3_reg[89][27]/P0001 ,
		_w11968_,
		_w11972_,
		_w17047_
	);
	LUT3 #(
		.INIT('h80)
	) name6535 (
		\wishbone_bd_ram_mem3_reg[252][27]/P0001 ,
		_w11952_,
		_w11954_,
		_w17048_
	);
	LUT3 #(
		.INIT('h80)
	) name6536 (
		\wishbone_bd_ram_mem3_reg[227][27]/P0001 ,
		_w11938_,
		_w11982_,
		_w17049_
	);
	LUT3 #(
		.INIT('h80)
	) name6537 (
		\wishbone_bd_ram_mem3_reg[13][27]/P0001 ,
		_w11932_,
		_w11966_,
		_w17050_
	);
	LUT4 #(
		.INIT('h0001)
	) name6538 (
		_w17047_,
		_w17048_,
		_w17049_,
		_w17050_,
		_w17051_
	);
	LUT3 #(
		.INIT('h80)
	) name6539 (
		\wishbone_bd_ram_mem3_reg[16][27]/P0001 ,
		_w11935_,
		_w11941_,
		_w17052_
	);
	LUT3 #(
		.INIT('h80)
	) name6540 (
		\wishbone_bd_ram_mem3_reg[175][27]/P0001 ,
		_w11930_,
		_w11973_,
		_w17053_
	);
	LUT3 #(
		.INIT('h80)
	) name6541 (
		\wishbone_bd_ram_mem3_reg[107][27]/P0001 ,
		_w11936_,
		_w11965_,
		_w17054_
	);
	LUT3 #(
		.INIT('h80)
	) name6542 (
		\wishbone_bd_ram_mem3_reg[181][27]/P0001 ,
		_w11933_,
		_w11942_,
		_w17055_
	);
	LUT4 #(
		.INIT('h0001)
	) name6543 (
		_w17052_,
		_w17053_,
		_w17054_,
		_w17055_,
		_w17056_
	);
	LUT4 #(
		.INIT('h8000)
	) name6544 (
		_w17041_,
		_w17046_,
		_w17051_,
		_w17056_,
		_w17057_
	);
	LUT3 #(
		.INIT('h80)
	) name6545 (
		\wishbone_bd_ram_mem3_reg[243][27]/P0001 ,
		_w11938_,
		_w11952_,
		_w17058_
	);
	LUT3 #(
		.INIT('h80)
	) name6546 (
		\wishbone_bd_ram_mem3_reg[122][27]/P0001 ,
		_w11944_,
		_w12012_,
		_w17059_
	);
	LUT3 #(
		.INIT('h80)
	) name6547 (
		\wishbone_bd_ram_mem3_reg[91][27]/P0001 ,
		_w11936_,
		_w11972_,
		_w17060_
	);
	LUT3 #(
		.INIT('h80)
	) name6548 (
		\wishbone_bd_ram_mem3_reg[65][27]/P0001 ,
		_w11949_,
		_w11977_,
		_w17061_
	);
	LUT4 #(
		.INIT('h0001)
	) name6549 (
		_w17058_,
		_w17059_,
		_w17060_,
		_w17061_,
		_w17062_
	);
	LUT3 #(
		.INIT('h80)
	) name6550 (
		\wishbone_bd_ram_mem3_reg[205][27]/P0001 ,
		_w11945_,
		_w11966_,
		_w17063_
	);
	LUT3 #(
		.INIT('h80)
	) name6551 (
		\wishbone_bd_ram_mem3_reg[78][27]/P0001 ,
		_w11948_,
		_w11949_,
		_w17064_
	);
	LUT3 #(
		.INIT('h80)
	) name6552 (
		\wishbone_bd_ram_mem3_reg[221][27]/P0001 ,
		_w11966_,
		_w11984_,
		_w17065_
	);
	LUT3 #(
		.INIT('h80)
	) name6553 (
		\wishbone_bd_ram_mem3_reg[88][27]/P0001 ,
		_w11972_,
		_w11990_,
		_w17066_
	);
	LUT4 #(
		.INIT('h0001)
	) name6554 (
		_w17063_,
		_w17064_,
		_w17065_,
		_w17066_,
		_w17067_
	);
	LUT3 #(
		.INIT('h80)
	) name6555 (
		\wishbone_bd_ram_mem3_reg[182][27]/P0001 ,
		_w11942_,
		_w11986_,
		_w17068_
	);
	LUT3 #(
		.INIT('h80)
	) name6556 (
		\wishbone_bd_ram_mem3_reg[51][27]/P0001 ,
		_w11938_,
		_w11979_,
		_w17069_
	);
	LUT3 #(
		.INIT('h80)
	) name6557 (
		\wishbone_bd_ram_mem3_reg[101][27]/P0001 ,
		_w11933_,
		_w11965_,
		_w17070_
	);
	LUT3 #(
		.INIT('h80)
	) name6558 (
		\wishbone_bd_ram_mem3_reg[210][27]/P0001 ,
		_w11963_,
		_w11984_,
		_w17071_
	);
	LUT4 #(
		.INIT('h0001)
	) name6559 (
		_w17068_,
		_w17069_,
		_w17070_,
		_w17071_,
		_w17072_
	);
	LUT3 #(
		.INIT('h80)
	) name6560 (
		\wishbone_bd_ram_mem3_reg[162][27]/P0001 ,
		_w11930_,
		_w11963_,
		_w17073_
	);
	LUT3 #(
		.INIT('h80)
	) name6561 (
		\wishbone_bd_ram_mem3_reg[238][27]/P0001 ,
		_w11948_,
		_w11982_,
		_w17074_
	);
	LUT3 #(
		.INIT('h80)
	) name6562 (
		\wishbone_bd_ram_mem3_reg[47][27]/P0001 ,
		_w11957_,
		_w11973_,
		_w17075_
	);
	LUT3 #(
		.INIT('h80)
	) name6563 (
		\wishbone_bd_ram_mem3_reg[201][27]/P0001 ,
		_w11945_,
		_w11968_,
		_w17076_
	);
	LUT4 #(
		.INIT('h0001)
	) name6564 (
		_w17073_,
		_w17074_,
		_w17075_,
		_w17076_,
		_w17077_
	);
	LUT4 #(
		.INIT('h8000)
	) name6565 (
		_w17062_,
		_w17067_,
		_w17072_,
		_w17077_,
		_w17078_
	);
	LUT3 #(
		.INIT('h80)
	) name6566 (
		\wishbone_bd_ram_mem3_reg[208][27]/P0001 ,
		_w11941_,
		_w11984_,
		_w17079_
	);
	LUT3 #(
		.INIT('h80)
	) name6567 (
		\wishbone_bd_ram_mem3_reg[192][27]/P0001 ,
		_w11941_,
		_w11945_,
		_w17080_
	);
	LUT3 #(
		.INIT('h80)
	) name6568 (
		\wishbone_bd_ram_mem3_reg[171][27]/P0001 ,
		_w11930_,
		_w11936_,
		_w17081_
	);
	LUT3 #(
		.INIT('h80)
	) name6569 (
		\wishbone_bd_ram_mem3_reg[98][27]/P0001 ,
		_w11963_,
		_w11965_,
		_w17082_
	);
	LUT4 #(
		.INIT('h0001)
	) name6570 (
		_w17079_,
		_w17080_,
		_w17081_,
		_w17082_,
		_w17083_
	);
	LUT3 #(
		.INIT('h80)
	) name6571 (
		\wishbone_bd_ram_mem3_reg[248][27]/P0001 ,
		_w11952_,
		_w11990_,
		_w17084_
	);
	LUT3 #(
		.INIT('h80)
	) name6572 (
		\wishbone_bd_ram_mem3_reg[126][27]/P0001 ,
		_w11948_,
		_w12012_,
		_w17085_
	);
	LUT3 #(
		.INIT('h80)
	) name6573 (
		\wishbone_bd_ram_mem3_reg[62][27]/P0001 ,
		_w11948_,
		_w11979_,
		_w17086_
	);
	LUT3 #(
		.INIT('h80)
	) name6574 (
		\wishbone_bd_ram_mem3_reg[58][27]/P0001 ,
		_w11944_,
		_w11979_,
		_w17087_
	);
	LUT4 #(
		.INIT('h0001)
	) name6575 (
		_w17084_,
		_w17085_,
		_w17086_,
		_w17087_,
		_w17088_
	);
	LUT3 #(
		.INIT('h80)
	) name6576 (
		\wishbone_bd_ram_mem3_reg[133][27]/P0001 ,
		_w11933_,
		_w11955_,
		_w17089_
	);
	LUT3 #(
		.INIT('h80)
	) name6577 (
		\wishbone_bd_ram_mem3_reg[60][27]/P0001 ,
		_w11954_,
		_w11979_,
		_w17090_
	);
	LUT3 #(
		.INIT('h80)
	) name6578 (
		\wishbone_bd_ram_mem3_reg[123][27]/P0001 ,
		_w11936_,
		_w12012_,
		_w17091_
	);
	LUT3 #(
		.INIT('h80)
	) name6579 (
		\wishbone_bd_ram_mem3_reg[84][27]/P0001 ,
		_w11929_,
		_w11972_,
		_w17092_
	);
	LUT4 #(
		.INIT('h0001)
	) name6580 (
		_w17089_,
		_w17090_,
		_w17091_,
		_w17092_,
		_w17093_
	);
	LUT3 #(
		.INIT('h80)
	) name6581 (
		\wishbone_bd_ram_mem3_reg[75][27]/P0001 ,
		_w11936_,
		_w11949_,
		_w17094_
	);
	LUT3 #(
		.INIT('h80)
	) name6582 (
		\wishbone_bd_ram_mem3_reg[25][27]/P0001 ,
		_w11935_,
		_w11968_,
		_w17095_
	);
	LUT3 #(
		.INIT('h80)
	) name6583 (
		\wishbone_bd_ram_mem3_reg[43][27]/P0001 ,
		_w11936_,
		_w11957_,
		_w17096_
	);
	LUT3 #(
		.INIT('h80)
	) name6584 (
		\wishbone_bd_ram_mem3_reg[153][27]/P0001 ,
		_w11959_,
		_w11968_,
		_w17097_
	);
	LUT4 #(
		.INIT('h0001)
	) name6585 (
		_w17094_,
		_w17095_,
		_w17096_,
		_w17097_,
		_w17098_
	);
	LUT4 #(
		.INIT('h8000)
	) name6586 (
		_w17083_,
		_w17088_,
		_w17093_,
		_w17098_,
		_w17099_
	);
	LUT4 #(
		.INIT('h8000)
	) name6587 (
		_w17036_,
		_w17057_,
		_w17078_,
		_w17099_,
		_w17100_
	);
	LUT3 #(
		.INIT('h80)
	) name6588 (
		\wishbone_bd_ram_mem3_reg[160][27]/P0001 ,
		_w11930_,
		_w11941_,
		_w17101_
	);
	LUT3 #(
		.INIT('h80)
	) name6589 (
		\wishbone_bd_ram_mem3_reg[198][27]/P0001 ,
		_w11945_,
		_w11986_,
		_w17102_
	);
	LUT3 #(
		.INIT('h80)
	) name6590 (
		\wishbone_bd_ram_mem3_reg[183][27]/P0001 ,
		_w11942_,
		_w11975_,
		_w17103_
	);
	LUT3 #(
		.INIT('h80)
	) name6591 (
		\wishbone_bd_ram_mem3_reg[121][27]/P0001 ,
		_w11968_,
		_w12012_,
		_w17104_
	);
	LUT4 #(
		.INIT('h0001)
	) name6592 (
		_w17101_,
		_w17102_,
		_w17103_,
		_w17104_,
		_w17105_
	);
	LUT3 #(
		.INIT('h80)
	) name6593 (
		\wishbone_bd_ram_mem3_reg[247][27]/P0001 ,
		_w11952_,
		_w11975_,
		_w17106_
	);
	LUT3 #(
		.INIT('h80)
	) name6594 (
		\wishbone_bd_ram_mem3_reg[232][27]/P0001 ,
		_w11982_,
		_w11990_,
		_w17107_
	);
	LUT3 #(
		.INIT('h80)
	) name6595 (
		\wishbone_bd_ram_mem3_reg[34][27]/P0001 ,
		_w11957_,
		_w11963_,
		_w17108_
	);
	LUT3 #(
		.INIT('h80)
	) name6596 (
		\wishbone_bd_ram_mem3_reg[8][27]/P0001 ,
		_w11932_,
		_w11990_,
		_w17109_
	);
	LUT4 #(
		.INIT('h0001)
	) name6597 (
		_w17106_,
		_w17107_,
		_w17108_,
		_w17109_,
		_w17110_
	);
	LUT3 #(
		.INIT('h80)
	) name6598 (
		\wishbone_bd_ram_mem3_reg[111][27]/P0001 ,
		_w11965_,
		_w11973_,
		_w17111_
	);
	LUT3 #(
		.INIT('h80)
	) name6599 (
		\wishbone_bd_ram_mem3_reg[117][27]/P0001 ,
		_w11933_,
		_w12012_,
		_w17112_
	);
	LUT3 #(
		.INIT('h80)
	) name6600 (
		\wishbone_bd_ram_mem3_reg[193][27]/P0001 ,
		_w11945_,
		_w11977_,
		_w17113_
	);
	LUT3 #(
		.INIT('h80)
	) name6601 (
		\wishbone_bd_ram_mem3_reg[220][27]/P0001 ,
		_w11954_,
		_w11984_,
		_w17114_
	);
	LUT4 #(
		.INIT('h0001)
	) name6602 (
		_w17111_,
		_w17112_,
		_w17113_,
		_w17114_,
		_w17115_
	);
	LUT3 #(
		.INIT('h80)
	) name6603 (
		\wishbone_bd_ram_mem3_reg[176][27]/P0001 ,
		_w11941_,
		_w11942_,
		_w17116_
	);
	LUT3 #(
		.INIT('h80)
	) name6604 (
		\wishbone_bd_ram_mem3_reg[148][27]/P0001 ,
		_w11929_,
		_w11959_,
		_w17117_
	);
	LUT3 #(
		.INIT('h80)
	) name6605 (
		\wishbone_bd_ram_mem3_reg[96][27]/P0001 ,
		_w11941_,
		_w11965_,
		_w17118_
	);
	LUT3 #(
		.INIT('h80)
	) name6606 (
		\wishbone_bd_ram_mem3_reg[184][27]/P0001 ,
		_w11942_,
		_w11990_,
		_w17119_
	);
	LUT4 #(
		.INIT('h0001)
	) name6607 (
		_w17116_,
		_w17117_,
		_w17118_,
		_w17119_,
		_w17120_
	);
	LUT4 #(
		.INIT('h8000)
	) name6608 (
		_w17105_,
		_w17110_,
		_w17115_,
		_w17120_,
		_w17121_
	);
	LUT3 #(
		.INIT('h80)
	) name6609 (
		\wishbone_bd_ram_mem3_reg[118][27]/P0001 ,
		_w11986_,
		_w12012_,
		_w17122_
	);
	LUT3 #(
		.INIT('h80)
	) name6610 (
		\wishbone_bd_ram_mem3_reg[203][27]/P0001 ,
		_w11936_,
		_w11945_,
		_w17123_
	);
	LUT3 #(
		.INIT('h80)
	) name6611 (
		\wishbone_bd_ram_mem3_reg[131][27]/P0001 ,
		_w11938_,
		_w11955_,
		_w17124_
	);
	LUT3 #(
		.INIT('h80)
	) name6612 (
		\wishbone_bd_ram_mem3_reg[70][27]/P0001 ,
		_w11949_,
		_w11986_,
		_w17125_
	);
	LUT4 #(
		.INIT('h0001)
	) name6613 (
		_w17122_,
		_w17123_,
		_w17124_,
		_w17125_,
		_w17126_
	);
	LUT3 #(
		.INIT('h80)
	) name6614 (
		\wishbone_bd_ram_mem3_reg[30][27]/P0001 ,
		_w11935_,
		_w11948_,
		_w17127_
	);
	LUT3 #(
		.INIT('h80)
	) name6615 (
		\wishbone_bd_ram_mem3_reg[26][27]/P0001 ,
		_w11935_,
		_w11944_,
		_w17128_
	);
	LUT3 #(
		.INIT('h80)
	) name6616 (
		\wishbone_bd_ram_mem3_reg[24][27]/P0001 ,
		_w11935_,
		_w11990_,
		_w17129_
	);
	LUT3 #(
		.INIT('h80)
	) name6617 (
		\wishbone_bd_ram_mem3_reg[104][27]/P0001 ,
		_w11965_,
		_w11990_,
		_w17130_
	);
	LUT4 #(
		.INIT('h0001)
	) name6618 (
		_w17127_,
		_w17128_,
		_w17129_,
		_w17130_,
		_w17131_
	);
	LUT3 #(
		.INIT('h80)
	) name6619 (
		\wishbone_bd_ram_mem3_reg[4][27]/P0001 ,
		_w11929_,
		_w11932_,
		_w17132_
	);
	LUT3 #(
		.INIT('h80)
	) name6620 (
		\wishbone_bd_ram_mem3_reg[94][27]/P0001 ,
		_w11948_,
		_w11972_,
		_w17133_
	);
	LUT3 #(
		.INIT('h80)
	) name6621 (
		\wishbone_bd_ram_mem3_reg[77][27]/P0001 ,
		_w11949_,
		_w11966_,
		_w17134_
	);
	LUT3 #(
		.INIT('h80)
	) name6622 (
		\wishbone_bd_ram_mem3_reg[32][27]/P0001 ,
		_w11941_,
		_w11957_,
		_w17135_
	);
	LUT4 #(
		.INIT('h0001)
	) name6623 (
		_w17132_,
		_w17133_,
		_w17134_,
		_w17135_,
		_w17136_
	);
	LUT3 #(
		.INIT('h80)
	) name6624 (
		\wishbone_bd_ram_mem3_reg[103][27]/P0001 ,
		_w11965_,
		_w11975_,
		_w17137_
	);
	LUT3 #(
		.INIT('h80)
	) name6625 (
		\wishbone_bd_ram_mem3_reg[216][27]/P0001 ,
		_w11984_,
		_w11990_,
		_w17138_
	);
	LUT3 #(
		.INIT('h80)
	) name6626 (
		\wishbone_bd_ram_mem3_reg[212][27]/P0001 ,
		_w11929_,
		_w11984_,
		_w17139_
	);
	LUT3 #(
		.INIT('h80)
	) name6627 (
		\wishbone_bd_ram_mem3_reg[155][27]/P0001 ,
		_w11936_,
		_w11959_,
		_w17140_
	);
	LUT4 #(
		.INIT('h0001)
	) name6628 (
		_w17137_,
		_w17138_,
		_w17139_,
		_w17140_,
		_w17141_
	);
	LUT4 #(
		.INIT('h8000)
	) name6629 (
		_w17126_,
		_w17131_,
		_w17136_,
		_w17141_,
		_w17142_
	);
	LUT3 #(
		.INIT('h80)
	) name6630 (
		\wishbone_bd_ram_mem3_reg[6][27]/P0001 ,
		_w11932_,
		_w11986_,
		_w17143_
	);
	LUT3 #(
		.INIT('h80)
	) name6631 (
		\wishbone_bd_ram_mem3_reg[110][27]/P0001 ,
		_w11948_,
		_w11965_,
		_w17144_
	);
	LUT3 #(
		.INIT('h80)
	) name6632 (
		\wishbone_bd_ram_mem3_reg[143][27]/P0001 ,
		_w11955_,
		_w11973_,
		_w17145_
	);
	LUT3 #(
		.INIT('h80)
	) name6633 (
		\wishbone_bd_ram_mem3_reg[173][27]/P0001 ,
		_w11930_,
		_w11966_,
		_w17146_
	);
	LUT4 #(
		.INIT('h0001)
	) name6634 (
		_w17143_,
		_w17144_,
		_w17145_,
		_w17146_,
		_w17147_
	);
	LUT3 #(
		.INIT('h80)
	) name6635 (
		\wishbone_bd_ram_mem3_reg[204][27]/P0001 ,
		_w11945_,
		_w11954_,
		_w17148_
	);
	LUT3 #(
		.INIT('h80)
	) name6636 (
		\wishbone_bd_ram_mem3_reg[213][27]/P0001 ,
		_w11933_,
		_w11984_,
		_w17149_
	);
	LUT3 #(
		.INIT('h80)
	) name6637 (
		\wishbone_bd_ram_mem3_reg[5][27]/P0001 ,
		_w11932_,
		_w11933_,
		_w17150_
	);
	LUT3 #(
		.INIT('h80)
	) name6638 (
		\wishbone_bd_ram_mem3_reg[61][27]/P0001 ,
		_w11966_,
		_w11979_,
		_w17151_
	);
	LUT4 #(
		.INIT('h0001)
	) name6639 (
		_w17148_,
		_w17149_,
		_w17150_,
		_w17151_,
		_w17152_
	);
	LUT3 #(
		.INIT('h80)
	) name6640 (
		\wishbone_bd_ram_mem3_reg[239][27]/P0001 ,
		_w11973_,
		_w11982_,
		_w17153_
	);
	LUT3 #(
		.INIT('h80)
	) name6641 (
		\wishbone_bd_ram_mem3_reg[164][27]/P0001 ,
		_w11929_,
		_w11930_,
		_w17154_
	);
	LUT3 #(
		.INIT('h80)
	) name6642 (
		\wishbone_bd_ram_mem3_reg[154][27]/P0001 ,
		_w11944_,
		_w11959_,
		_w17155_
	);
	LUT3 #(
		.INIT('h80)
	) name6643 (
		\wishbone_bd_ram_mem3_reg[244][27]/P0001 ,
		_w11929_,
		_w11952_,
		_w17156_
	);
	LUT4 #(
		.INIT('h0001)
	) name6644 (
		_w17153_,
		_w17154_,
		_w17155_,
		_w17156_,
		_w17157_
	);
	LUT3 #(
		.INIT('h80)
	) name6645 (
		\wishbone_bd_ram_mem3_reg[189][27]/P0001 ,
		_w11942_,
		_w11966_,
		_w17158_
	);
	LUT3 #(
		.INIT('h80)
	) name6646 (
		\wishbone_bd_ram_mem3_reg[249][27]/P0001 ,
		_w11952_,
		_w11968_,
		_w17159_
	);
	LUT3 #(
		.INIT('h80)
	) name6647 (
		\wishbone_bd_ram_mem3_reg[138][27]/P0001 ,
		_w11944_,
		_w11955_,
		_w17160_
	);
	LUT3 #(
		.INIT('h80)
	) name6648 (
		\wishbone_bd_ram_mem3_reg[99][27]/P0001 ,
		_w11938_,
		_w11965_,
		_w17161_
	);
	LUT4 #(
		.INIT('h0001)
	) name6649 (
		_w17158_,
		_w17159_,
		_w17160_,
		_w17161_,
		_w17162_
	);
	LUT4 #(
		.INIT('h8000)
	) name6650 (
		_w17147_,
		_w17152_,
		_w17157_,
		_w17162_,
		_w17163_
	);
	LUT3 #(
		.INIT('h80)
	) name6651 (
		\wishbone_bd_ram_mem3_reg[49][27]/P0001 ,
		_w11977_,
		_w11979_,
		_w17164_
	);
	LUT3 #(
		.INIT('h80)
	) name6652 (
		\wishbone_bd_ram_mem3_reg[53][27]/P0001 ,
		_w11933_,
		_w11979_,
		_w17165_
	);
	LUT3 #(
		.INIT('h80)
	) name6653 (
		\wishbone_bd_ram_mem3_reg[222][27]/P0001 ,
		_w11948_,
		_w11984_,
		_w17166_
	);
	LUT3 #(
		.INIT('h80)
	) name6654 (
		\wishbone_bd_ram_mem3_reg[31][27]/P0001 ,
		_w11935_,
		_w11973_,
		_w17167_
	);
	LUT4 #(
		.INIT('h0001)
	) name6655 (
		_w17164_,
		_w17165_,
		_w17166_,
		_w17167_,
		_w17168_
	);
	LUT3 #(
		.INIT('h80)
	) name6656 (
		\wishbone_bd_ram_mem3_reg[134][27]/P0001 ,
		_w11955_,
		_w11986_,
		_w17169_
	);
	LUT3 #(
		.INIT('h80)
	) name6657 (
		\wishbone_bd_ram_mem3_reg[187][27]/P0001 ,
		_w11936_,
		_w11942_,
		_w17170_
	);
	LUT3 #(
		.INIT('h80)
	) name6658 (
		\wishbone_bd_ram_mem3_reg[7][27]/P0001 ,
		_w11932_,
		_w11975_,
		_w17171_
	);
	LUT3 #(
		.INIT('h80)
	) name6659 (
		\wishbone_bd_ram_mem3_reg[63][27]/P0001 ,
		_w11973_,
		_w11979_,
		_w17172_
	);
	LUT4 #(
		.INIT('h0001)
	) name6660 (
		_w17169_,
		_w17170_,
		_w17171_,
		_w17172_,
		_w17173_
	);
	LUT3 #(
		.INIT('h80)
	) name6661 (
		\wishbone_bd_ram_mem3_reg[127][27]/P0001 ,
		_w11973_,
		_w12012_,
		_w17174_
	);
	LUT3 #(
		.INIT('h80)
	) name6662 (
		\wishbone_bd_ram_mem3_reg[116][27]/P0001 ,
		_w11929_,
		_w12012_,
		_w17175_
	);
	LUT3 #(
		.INIT('h80)
	) name6663 (
		\wishbone_bd_ram_mem3_reg[159][27]/P0001 ,
		_w11959_,
		_w11973_,
		_w17176_
	);
	LUT3 #(
		.INIT('h80)
	) name6664 (
		\wishbone_bd_ram_mem3_reg[233][27]/P0001 ,
		_w11968_,
		_w11982_,
		_w17177_
	);
	LUT4 #(
		.INIT('h0001)
	) name6665 (
		_w17174_,
		_w17175_,
		_w17176_,
		_w17177_,
		_w17178_
	);
	LUT3 #(
		.INIT('h80)
	) name6666 (
		\wishbone_bd_ram_mem3_reg[179][27]/P0001 ,
		_w11938_,
		_w11942_,
		_w17179_
	);
	LUT3 #(
		.INIT('h80)
	) name6667 (
		\wishbone_bd_ram_mem3_reg[190][27]/P0001 ,
		_w11942_,
		_w11948_,
		_w17180_
	);
	LUT3 #(
		.INIT('h80)
	) name6668 (
		\wishbone_bd_ram_mem3_reg[130][27]/P0001 ,
		_w11955_,
		_w11963_,
		_w17181_
	);
	LUT3 #(
		.INIT('h80)
	) name6669 (
		\wishbone_bd_ram_mem3_reg[39][27]/P0001 ,
		_w11957_,
		_w11975_,
		_w17182_
	);
	LUT4 #(
		.INIT('h0001)
	) name6670 (
		_w17179_,
		_w17180_,
		_w17181_,
		_w17182_,
		_w17183_
	);
	LUT4 #(
		.INIT('h8000)
	) name6671 (
		_w17168_,
		_w17173_,
		_w17178_,
		_w17183_,
		_w17184_
	);
	LUT4 #(
		.INIT('h8000)
	) name6672 (
		_w17121_,
		_w17142_,
		_w17163_,
		_w17184_,
		_w17185_
	);
	LUT3 #(
		.INIT('h80)
	) name6673 (
		\wishbone_bd_ram_mem3_reg[18][27]/P0001 ,
		_w11935_,
		_w11963_,
		_w17186_
	);
	LUT3 #(
		.INIT('h80)
	) name6674 (
		\wishbone_bd_ram_mem3_reg[1][27]/P0001 ,
		_w11932_,
		_w11977_,
		_w17187_
	);
	LUT3 #(
		.INIT('h80)
	) name6675 (
		\wishbone_bd_ram_mem3_reg[167][27]/P0001 ,
		_w11930_,
		_w11975_,
		_w17188_
	);
	LUT3 #(
		.INIT('h80)
	) name6676 (
		\wishbone_bd_ram_mem3_reg[250][27]/P0001 ,
		_w11944_,
		_w11952_,
		_w17189_
	);
	LUT4 #(
		.INIT('h0001)
	) name6677 (
		_w17186_,
		_w17187_,
		_w17188_,
		_w17189_,
		_w17190_
	);
	LUT3 #(
		.INIT('h80)
	) name6678 (
		\wishbone_bd_ram_mem3_reg[149][27]/P0001 ,
		_w11933_,
		_w11959_,
		_w17191_
	);
	LUT3 #(
		.INIT('h80)
	) name6679 (
		\wishbone_bd_ram_mem3_reg[21][27]/P0001 ,
		_w11933_,
		_w11935_,
		_w17192_
	);
	LUT3 #(
		.INIT('h80)
	) name6680 (
		\wishbone_bd_ram_mem3_reg[207][27]/P0001 ,
		_w11945_,
		_w11973_,
		_w17193_
	);
	LUT3 #(
		.INIT('h80)
	) name6681 (
		\wishbone_bd_ram_mem3_reg[165][27]/P0001 ,
		_w11930_,
		_w11933_,
		_w17194_
	);
	LUT4 #(
		.INIT('h0001)
	) name6682 (
		_w17191_,
		_w17192_,
		_w17193_,
		_w17194_,
		_w17195_
	);
	LUT3 #(
		.INIT('h80)
	) name6683 (
		\wishbone_bd_ram_mem3_reg[174][27]/P0001 ,
		_w11930_,
		_w11948_,
		_w17196_
	);
	LUT3 #(
		.INIT('h80)
	) name6684 (
		\wishbone_bd_ram_mem3_reg[40][27]/P0001 ,
		_w11957_,
		_w11990_,
		_w17197_
	);
	LUT3 #(
		.INIT('h80)
	) name6685 (
		\wishbone_bd_ram_mem3_reg[236][27]/P0001 ,
		_w11954_,
		_w11982_,
		_w17198_
	);
	LUT3 #(
		.INIT('h80)
	) name6686 (
		\wishbone_bd_ram_mem3_reg[81][27]/P0001 ,
		_w11972_,
		_w11977_,
		_w17199_
	);
	LUT4 #(
		.INIT('h0001)
	) name6687 (
		_w17196_,
		_w17197_,
		_w17198_,
		_w17199_,
		_w17200_
	);
	LUT3 #(
		.INIT('h80)
	) name6688 (
		\wishbone_bd_ram_mem3_reg[157][27]/P0001 ,
		_w11959_,
		_w11966_,
		_w17201_
	);
	LUT3 #(
		.INIT('h80)
	) name6689 (
		\wishbone_bd_ram_mem3_reg[166][27]/P0001 ,
		_w11930_,
		_w11986_,
		_w17202_
	);
	LUT3 #(
		.INIT('h80)
	) name6690 (
		\wishbone_bd_ram_mem3_reg[228][27]/P0001 ,
		_w11929_,
		_w11982_,
		_w17203_
	);
	LUT3 #(
		.INIT('h80)
	) name6691 (
		\wishbone_bd_ram_mem3_reg[28][27]/P0001 ,
		_w11935_,
		_w11954_,
		_w17204_
	);
	LUT4 #(
		.INIT('h0001)
	) name6692 (
		_w17201_,
		_w17202_,
		_w17203_,
		_w17204_,
		_w17205_
	);
	LUT4 #(
		.INIT('h8000)
	) name6693 (
		_w17190_,
		_w17195_,
		_w17200_,
		_w17205_,
		_w17206_
	);
	LUT3 #(
		.INIT('h80)
	) name6694 (
		\wishbone_bd_ram_mem3_reg[206][27]/P0001 ,
		_w11945_,
		_w11948_,
		_w17207_
	);
	LUT3 #(
		.INIT('h80)
	) name6695 (
		\wishbone_bd_ram_mem3_reg[9][27]/P0001 ,
		_w11932_,
		_w11968_,
		_w17208_
	);
	LUT3 #(
		.INIT('h80)
	) name6696 (
		\wishbone_bd_ram_mem3_reg[27][27]/P0001 ,
		_w11935_,
		_w11936_,
		_w17209_
	);
	LUT3 #(
		.INIT('h80)
	) name6697 (
		\wishbone_bd_ram_mem3_reg[95][27]/P0001 ,
		_w11972_,
		_w11973_,
		_w17210_
	);
	LUT4 #(
		.INIT('h0001)
	) name6698 (
		_w17207_,
		_w17208_,
		_w17209_,
		_w17210_,
		_w17211_
	);
	LUT3 #(
		.INIT('h80)
	) name6699 (
		\wishbone_bd_ram_mem3_reg[240][27]/P0001 ,
		_w11941_,
		_w11952_,
		_w17212_
	);
	LUT3 #(
		.INIT('h80)
	) name6700 (
		\wishbone_bd_ram_mem3_reg[97][27]/P0001 ,
		_w11965_,
		_w11977_,
		_w17213_
	);
	LUT3 #(
		.INIT('h80)
	) name6701 (
		\wishbone_bd_ram_mem3_reg[139][27]/P0001 ,
		_w11936_,
		_w11955_,
		_w17214_
	);
	LUT3 #(
		.INIT('h80)
	) name6702 (
		\wishbone_bd_ram_mem3_reg[234][27]/P0001 ,
		_w11944_,
		_w11982_,
		_w17215_
	);
	LUT4 #(
		.INIT('h0001)
	) name6703 (
		_w17212_,
		_w17213_,
		_w17214_,
		_w17215_,
		_w17216_
	);
	LUT3 #(
		.INIT('h80)
	) name6704 (
		\wishbone_bd_ram_mem3_reg[38][27]/P0001 ,
		_w11957_,
		_w11986_,
		_w17217_
	);
	LUT3 #(
		.INIT('h80)
	) name6705 (
		\wishbone_bd_ram_mem3_reg[2][27]/P0001 ,
		_w11932_,
		_w11963_,
		_w17218_
	);
	LUT3 #(
		.INIT('h80)
	) name6706 (
		\wishbone_bd_ram_mem3_reg[115][27]/P0001 ,
		_w11938_,
		_w12012_,
		_w17219_
	);
	LUT3 #(
		.INIT('h80)
	) name6707 (
		\wishbone_bd_ram_mem3_reg[23][27]/P0001 ,
		_w11935_,
		_w11975_,
		_w17220_
	);
	LUT4 #(
		.INIT('h0001)
	) name6708 (
		_w17217_,
		_w17218_,
		_w17219_,
		_w17220_,
		_w17221_
	);
	LUT3 #(
		.INIT('h80)
	) name6709 (
		\wishbone_bd_ram_mem3_reg[163][27]/P0001 ,
		_w11930_,
		_w11938_,
		_w17222_
	);
	LUT3 #(
		.INIT('h80)
	) name6710 (
		\wishbone_bd_ram_mem3_reg[41][27]/P0001 ,
		_w11957_,
		_w11968_,
		_w17223_
	);
	LUT3 #(
		.INIT('h80)
	) name6711 (
		\wishbone_bd_ram_mem3_reg[36][27]/P0001 ,
		_w11929_,
		_w11957_,
		_w17224_
	);
	LUT3 #(
		.INIT('h80)
	) name6712 (
		\wishbone_bd_ram_mem3_reg[71][27]/P0001 ,
		_w11949_,
		_w11975_,
		_w17225_
	);
	LUT4 #(
		.INIT('h0001)
	) name6713 (
		_w17222_,
		_w17223_,
		_w17224_,
		_w17225_,
		_w17226_
	);
	LUT4 #(
		.INIT('h8000)
	) name6714 (
		_w17211_,
		_w17216_,
		_w17221_,
		_w17226_,
		_w17227_
	);
	LUT3 #(
		.INIT('h80)
	) name6715 (
		\wishbone_bd_ram_mem3_reg[253][27]/P0001 ,
		_w11952_,
		_w11966_,
		_w17228_
	);
	LUT3 #(
		.INIT('h80)
	) name6716 (
		\wishbone_bd_ram_mem3_reg[109][27]/P0001 ,
		_w11965_,
		_w11966_,
		_w17229_
	);
	LUT3 #(
		.INIT('h80)
	) name6717 (
		\wishbone_bd_ram_mem3_reg[69][27]/P0001 ,
		_w11933_,
		_w11949_,
		_w17230_
	);
	LUT3 #(
		.INIT('h80)
	) name6718 (
		\wishbone_bd_ram_mem3_reg[199][27]/P0001 ,
		_w11945_,
		_w11975_,
		_w17231_
	);
	LUT4 #(
		.INIT('h0001)
	) name6719 (
		_w17228_,
		_w17229_,
		_w17230_,
		_w17231_,
		_w17232_
	);
	LUT3 #(
		.INIT('h80)
	) name6720 (
		\wishbone_bd_ram_mem3_reg[245][27]/P0001 ,
		_w11933_,
		_w11952_,
		_w17233_
	);
	LUT3 #(
		.INIT('h80)
	) name6721 (
		\wishbone_bd_ram_mem3_reg[146][27]/P0001 ,
		_w11959_,
		_w11963_,
		_w17234_
	);
	LUT3 #(
		.INIT('h80)
	) name6722 (
		\wishbone_bd_ram_mem3_reg[45][27]/P0001 ,
		_w11957_,
		_w11966_,
		_w17235_
	);
	LUT3 #(
		.INIT('h80)
	) name6723 (
		\wishbone_bd_ram_mem3_reg[66][27]/P0001 ,
		_w11949_,
		_w11963_,
		_w17236_
	);
	LUT4 #(
		.INIT('h0001)
	) name6724 (
		_w17233_,
		_w17234_,
		_w17235_,
		_w17236_,
		_w17237_
	);
	LUT3 #(
		.INIT('h80)
	) name6725 (
		\wishbone_bd_ram_mem3_reg[72][27]/P0001 ,
		_w11949_,
		_w11990_,
		_w17238_
	);
	LUT3 #(
		.INIT('h80)
	) name6726 (
		\wishbone_bd_ram_mem3_reg[241][27]/P0001 ,
		_w11952_,
		_w11977_,
		_w17239_
	);
	LUT3 #(
		.INIT('h80)
	) name6727 (
		\wishbone_bd_ram_mem3_reg[56][27]/P0001 ,
		_w11979_,
		_w11990_,
		_w17240_
	);
	LUT3 #(
		.INIT('h80)
	) name6728 (
		\wishbone_bd_ram_mem3_reg[140][27]/P0001 ,
		_w11954_,
		_w11955_,
		_w17241_
	);
	LUT4 #(
		.INIT('h0001)
	) name6729 (
		_w17238_,
		_w17239_,
		_w17240_,
		_w17241_,
		_w17242_
	);
	LUT3 #(
		.INIT('h80)
	) name6730 (
		\wishbone_bd_ram_mem3_reg[57][27]/P0001 ,
		_w11968_,
		_w11979_,
		_w17243_
	);
	LUT3 #(
		.INIT('h80)
	) name6731 (
		\wishbone_bd_ram_mem3_reg[100][27]/P0001 ,
		_w11929_,
		_w11965_,
		_w17244_
	);
	LUT3 #(
		.INIT('h80)
	) name6732 (
		\wishbone_bd_ram_mem3_reg[59][27]/P0001 ,
		_w11936_,
		_w11979_,
		_w17245_
	);
	LUT3 #(
		.INIT('h80)
	) name6733 (
		\wishbone_bd_ram_mem3_reg[10][27]/P0001 ,
		_w11932_,
		_w11944_,
		_w17246_
	);
	LUT4 #(
		.INIT('h0001)
	) name6734 (
		_w17243_,
		_w17244_,
		_w17245_,
		_w17246_,
		_w17247_
	);
	LUT4 #(
		.INIT('h8000)
	) name6735 (
		_w17232_,
		_w17237_,
		_w17242_,
		_w17247_,
		_w17248_
	);
	LUT3 #(
		.INIT('h80)
	) name6736 (
		\wishbone_bd_ram_mem3_reg[106][27]/P0001 ,
		_w11944_,
		_w11965_,
		_w17249_
	);
	LUT3 #(
		.INIT('h80)
	) name6737 (
		\wishbone_bd_ram_mem3_reg[255][27]/P0001 ,
		_w11952_,
		_w11973_,
		_w17250_
	);
	LUT3 #(
		.INIT('h80)
	) name6738 (
		\wishbone_bd_ram_mem3_reg[87][27]/P0001 ,
		_w11972_,
		_w11975_,
		_w17251_
	);
	LUT3 #(
		.INIT('h80)
	) name6739 (
		\wishbone_bd_ram_mem3_reg[15][27]/P0001 ,
		_w11932_,
		_w11973_,
		_w17252_
	);
	LUT4 #(
		.INIT('h0001)
	) name6740 (
		_w17249_,
		_w17250_,
		_w17251_,
		_w17252_,
		_w17253_
	);
	LUT3 #(
		.INIT('h80)
	) name6741 (
		\wishbone_bd_ram_mem3_reg[230][27]/P0001 ,
		_w11982_,
		_w11986_,
		_w17254_
	);
	LUT3 #(
		.INIT('h80)
	) name6742 (
		\wishbone_bd_ram_mem3_reg[170][27]/P0001 ,
		_w11930_,
		_w11944_,
		_w17255_
	);
	LUT3 #(
		.INIT('h80)
	) name6743 (
		\wishbone_bd_ram_mem3_reg[217][27]/P0001 ,
		_w11968_,
		_w11984_,
		_w17256_
	);
	LUT3 #(
		.INIT('h80)
	) name6744 (
		\wishbone_bd_ram_mem3_reg[191][27]/P0001 ,
		_w11942_,
		_w11973_,
		_w17257_
	);
	LUT4 #(
		.INIT('h0001)
	) name6745 (
		_w17254_,
		_w17255_,
		_w17256_,
		_w17257_,
		_w17258_
	);
	LUT3 #(
		.INIT('h80)
	) name6746 (
		\wishbone_bd_ram_mem3_reg[194][27]/P0001 ,
		_w11945_,
		_w11963_,
		_w17259_
	);
	LUT3 #(
		.INIT('h80)
	) name6747 (
		\wishbone_bd_ram_mem3_reg[161][27]/P0001 ,
		_w11930_,
		_w11977_,
		_w17260_
	);
	LUT3 #(
		.INIT('h80)
	) name6748 (
		\wishbone_bd_ram_mem3_reg[14][27]/P0001 ,
		_w11932_,
		_w11948_,
		_w17261_
	);
	LUT3 #(
		.INIT('h80)
	) name6749 (
		\wishbone_bd_ram_mem3_reg[202][27]/P0001 ,
		_w11944_,
		_w11945_,
		_w17262_
	);
	LUT4 #(
		.INIT('h0001)
	) name6750 (
		_w17259_,
		_w17260_,
		_w17261_,
		_w17262_,
		_w17263_
	);
	LUT3 #(
		.INIT('h80)
	) name6751 (
		\wishbone_bd_ram_mem3_reg[22][27]/P0001 ,
		_w11935_,
		_w11986_,
		_w17264_
	);
	LUT3 #(
		.INIT('h80)
	) name6752 (
		\wishbone_bd_ram_mem3_reg[64][27]/P0001 ,
		_w11941_,
		_w11949_,
		_w17265_
	);
	LUT3 #(
		.INIT('h80)
	) name6753 (
		\wishbone_bd_ram_mem3_reg[17][27]/P0001 ,
		_w11935_,
		_w11977_,
		_w17266_
	);
	LUT3 #(
		.INIT('h80)
	) name6754 (
		\wishbone_bd_ram_mem3_reg[33][27]/P0001 ,
		_w11957_,
		_w11977_,
		_w17267_
	);
	LUT4 #(
		.INIT('h0001)
	) name6755 (
		_w17264_,
		_w17265_,
		_w17266_,
		_w17267_,
		_w17268_
	);
	LUT4 #(
		.INIT('h8000)
	) name6756 (
		_w17253_,
		_w17258_,
		_w17263_,
		_w17268_,
		_w17269_
	);
	LUT4 #(
		.INIT('h8000)
	) name6757 (
		_w17206_,
		_w17227_,
		_w17248_,
		_w17269_,
		_w17270_
	);
	LUT3 #(
		.INIT('h80)
	) name6758 (
		\wishbone_bd_ram_mem3_reg[20][27]/P0001 ,
		_w11929_,
		_w11935_,
		_w17271_
	);
	LUT3 #(
		.INIT('h80)
	) name6759 (
		\wishbone_bd_ram_mem3_reg[172][27]/P0001 ,
		_w11930_,
		_w11954_,
		_w17272_
	);
	LUT3 #(
		.INIT('h80)
	) name6760 (
		\wishbone_bd_ram_mem3_reg[218][27]/P0001 ,
		_w11944_,
		_w11984_,
		_w17273_
	);
	LUT3 #(
		.INIT('h80)
	) name6761 (
		\wishbone_bd_ram_mem3_reg[93][27]/P0001 ,
		_w11966_,
		_w11972_,
		_w17274_
	);
	LUT4 #(
		.INIT('h0001)
	) name6762 (
		_w17271_,
		_w17272_,
		_w17273_,
		_w17274_,
		_w17275_
	);
	LUT3 #(
		.INIT('h80)
	) name6763 (
		\wishbone_bd_ram_mem3_reg[125][27]/P0001 ,
		_w11966_,
		_w12012_,
		_w17276_
	);
	LUT3 #(
		.INIT('h80)
	) name6764 (
		\wishbone_bd_ram_mem3_reg[54][27]/P0001 ,
		_w11979_,
		_w11986_,
		_w17277_
	);
	LUT3 #(
		.INIT('h80)
	) name6765 (
		\wishbone_bd_ram_mem3_reg[141][27]/P0001 ,
		_w11955_,
		_w11966_,
		_w17278_
	);
	LUT3 #(
		.INIT('h80)
	) name6766 (
		\wishbone_bd_ram_mem3_reg[178][27]/P0001 ,
		_w11942_,
		_w11963_,
		_w17279_
	);
	LUT4 #(
		.INIT('h0001)
	) name6767 (
		_w17276_,
		_w17277_,
		_w17278_,
		_w17279_,
		_w17280_
	);
	LUT3 #(
		.INIT('h80)
	) name6768 (
		\wishbone_bd_ram_mem3_reg[168][27]/P0001 ,
		_w11930_,
		_w11990_,
		_w17281_
	);
	LUT3 #(
		.INIT('h80)
	) name6769 (
		\wishbone_bd_ram_mem3_reg[254][27]/P0001 ,
		_w11948_,
		_w11952_,
		_w17282_
	);
	LUT3 #(
		.INIT('h80)
	) name6770 (
		\wishbone_bd_ram_mem3_reg[46][27]/P0001 ,
		_w11948_,
		_w11957_,
		_w17283_
	);
	LUT3 #(
		.INIT('h80)
	) name6771 (
		\wishbone_bd_ram_mem3_reg[223][27]/P0001 ,
		_w11973_,
		_w11984_,
		_w17284_
	);
	LUT4 #(
		.INIT('h0001)
	) name6772 (
		_w17281_,
		_w17282_,
		_w17283_,
		_w17284_,
		_w17285_
	);
	LUT3 #(
		.INIT('h80)
	) name6773 (
		\wishbone_bd_ram_mem3_reg[11][27]/P0001 ,
		_w11932_,
		_w11936_,
		_w17286_
	);
	LUT3 #(
		.INIT('h80)
	) name6774 (
		\wishbone_bd_ram_mem3_reg[79][27]/P0001 ,
		_w11949_,
		_w11973_,
		_w17287_
	);
	LUT3 #(
		.INIT('h80)
	) name6775 (
		\wishbone_bd_ram_mem3_reg[137][27]/P0001 ,
		_w11955_,
		_w11968_,
		_w17288_
	);
	LUT3 #(
		.INIT('h80)
	) name6776 (
		\wishbone_bd_ram_mem3_reg[135][27]/P0001 ,
		_w11955_,
		_w11975_,
		_w17289_
	);
	LUT4 #(
		.INIT('h0001)
	) name6777 (
		_w17286_,
		_w17287_,
		_w17288_,
		_w17289_,
		_w17290_
	);
	LUT4 #(
		.INIT('h8000)
	) name6778 (
		_w17275_,
		_w17280_,
		_w17285_,
		_w17290_,
		_w17291_
	);
	LUT3 #(
		.INIT('h80)
	) name6779 (
		\wishbone_bd_ram_mem3_reg[102][27]/P0001 ,
		_w11965_,
		_w11986_,
		_w17292_
	);
	LUT3 #(
		.INIT('h80)
	) name6780 (
		\wishbone_bd_ram_mem3_reg[35][27]/P0001 ,
		_w11938_,
		_w11957_,
		_w17293_
	);
	LUT3 #(
		.INIT('h80)
	) name6781 (
		\wishbone_bd_ram_mem3_reg[29][27]/P0001 ,
		_w11935_,
		_w11966_,
		_w17294_
	);
	LUT3 #(
		.INIT('h80)
	) name6782 (
		\wishbone_bd_ram_mem3_reg[151][27]/P0001 ,
		_w11959_,
		_w11975_,
		_w17295_
	);
	LUT4 #(
		.INIT('h0001)
	) name6783 (
		_w17292_,
		_w17293_,
		_w17294_,
		_w17295_,
		_w17296_
	);
	LUT3 #(
		.INIT('h80)
	) name6784 (
		\wishbone_bd_ram_mem3_reg[144][27]/P0001 ,
		_w11941_,
		_w11959_,
		_w17297_
	);
	LUT3 #(
		.INIT('h80)
	) name6785 (
		\wishbone_bd_ram_mem3_reg[142][27]/P0001 ,
		_w11948_,
		_w11955_,
		_w17298_
	);
	LUT3 #(
		.INIT('h80)
	) name6786 (
		\wishbone_bd_ram_mem3_reg[83][27]/P0001 ,
		_w11938_,
		_w11972_,
		_w17299_
	);
	LUT3 #(
		.INIT('h80)
	) name6787 (
		\wishbone_bd_ram_mem3_reg[76][27]/P0001 ,
		_w11949_,
		_w11954_,
		_w17300_
	);
	LUT4 #(
		.INIT('h0001)
	) name6788 (
		_w17297_,
		_w17298_,
		_w17299_,
		_w17300_,
		_w17301_
	);
	LUT3 #(
		.INIT('h80)
	) name6789 (
		\wishbone_bd_ram_mem3_reg[209][27]/P0001 ,
		_w11977_,
		_w11984_,
		_w17302_
	);
	LUT3 #(
		.INIT('h80)
	) name6790 (
		\wishbone_bd_ram_mem3_reg[158][27]/P0001 ,
		_w11948_,
		_w11959_,
		_w17303_
	);
	LUT3 #(
		.INIT('h80)
	) name6791 (
		\wishbone_bd_ram_mem3_reg[112][27]/P0001 ,
		_w11941_,
		_w12012_,
		_w17304_
	);
	LUT3 #(
		.INIT('h80)
	) name6792 (
		\wishbone_bd_ram_mem3_reg[85][27]/P0001 ,
		_w11933_,
		_w11972_,
		_w17305_
	);
	LUT4 #(
		.INIT('h0001)
	) name6793 (
		_w17302_,
		_w17303_,
		_w17304_,
		_w17305_,
		_w17306_
	);
	LUT3 #(
		.INIT('h80)
	) name6794 (
		\wishbone_bd_ram_mem3_reg[12][27]/P0001 ,
		_w11932_,
		_w11954_,
		_w17307_
	);
	LUT3 #(
		.INIT('h80)
	) name6795 (
		\wishbone_bd_ram_mem3_reg[86][27]/P0001 ,
		_w11972_,
		_w11986_,
		_w17308_
	);
	LUT3 #(
		.INIT('h80)
	) name6796 (
		\wishbone_bd_ram_mem3_reg[215][27]/P0001 ,
		_w11975_,
		_w11984_,
		_w17309_
	);
	LUT3 #(
		.INIT('h80)
	) name6797 (
		\wishbone_bd_ram_mem3_reg[129][27]/P0001 ,
		_w11955_,
		_w11977_,
		_w17310_
	);
	LUT4 #(
		.INIT('h0001)
	) name6798 (
		_w17307_,
		_w17308_,
		_w17309_,
		_w17310_,
		_w17311_
	);
	LUT4 #(
		.INIT('h8000)
	) name6799 (
		_w17296_,
		_w17301_,
		_w17306_,
		_w17311_,
		_w17312_
	);
	LUT3 #(
		.INIT('h80)
	) name6800 (
		\wishbone_bd_ram_mem3_reg[197][27]/P0001 ,
		_w11933_,
		_w11945_,
		_w17313_
	);
	LUT3 #(
		.INIT('h80)
	) name6801 (
		\wishbone_bd_ram_mem3_reg[67][27]/P0001 ,
		_w11938_,
		_w11949_,
		_w17314_
	);
	LUT3 #(
		.INIT('h80)
	) name6802 (
		\wishbone_bd_ram_mem3_reg[114][27]/P0001 ,
		_w11963_,
		_w12012_,
		_w17315_
	);
	LUT3 #(
		.INIT('h80)
	) name6803 (
		\wishbone_bd_ram_mem3_reg[188][27]/P0001 ,
		_w11942_,
		_w11954_,
		_w17316_
	);
	LUT4 #(
		.INIT('h0001)
	) name6804 (
		_w17313_,
		_w17314_,
		_w17315_,
		_w17316_,
		_w17317_
	);
	LUT3 #(
		.INIT('h80)
	) name6805 (
		\wishbone_bd_ram_mem3_reg[145][27]/P0001 ,
		_w11959_,
		_w11977_,
		_w17318_
	);
	LUT3 #(
		.INIT('h80)
	) name6806 (
		\wishbone_bd_ram_mem3_reg[186][27]/P0001 ,
		_w11942_,
		_w11944_,
		_w17319_
	);
	LUT3 #(
		.INIT('h80)
	) name6807 (
		\wishbone_bd_ram_mem3_reg[150][27]/P0001 ,
		_w11959_,
		_w11986_,
		_w17320_
	);
	LUT3 #(
		.INIT('h80)
	) name6808 (
		\wishbone_bd_ram_mem3_reg[211][27]/P0001 ,
		_w11938_,
		_w11984_,
		_w17321_
	);
	LUT4 #(
		.INIT('h0001)
	) name6809 (
		_w17318_,
		_w17319_,
		_w17320_,
		_w17321_,
		_w17322_
	);
	LUT3 #(
		.INIT('h80)
	) name6810 (
		\wishbone_bd_ram_mem3_reg[42][27]/P0001 ,
		_w11944_,
		_w11957_,
		_w17323_
	);
	LUT3 #(
		.INIT('h80)
	) name6811 (
		\wishbone_bd_ram_mem3_reg[48][27]/P0001 ,
		_w11941_,
		_w11979_,
		_w17324_
	);
	LUT3 #(
		.INIT('h80)
	) name6812 (
		\wishbone_bd_ram_mem3_reg[44][27]/P0001 ,
		_w11954_,
		_w11957_,
		_w17325_
	);
	LUT3 #(
		.INIT('h80)
	) name6813 (
		\wishbone_bd_ram_mem3_reg[237][27]/P0001 ,
		_w11966_,
		_w11982_,
		_w17326_
	);
	LUT4 #(
		.INIT('h0001)
	) name6814 (
		_w17323_,
		_w17324_,
		_w17325_,
		_w17326_,
		_w17327_
	);
	LUT3 #(
		.INIT('h80)
	) name6815 (
		\wishbone_bd_ram_mem3_reg[226][27]/P0001 ,
		_w11963_,
		_w11982_,
		_w17328_
	);
	LUT3 #(
		.INIT('h80)
	) name6816 (
		\wishbone_bd_ram_mem3_reg[108][27]/P0001 ,
		_w11954_,
		_w11965_,
		_w17329_
	);
	LUT3 #(
		.INIT('h80)
	) name6817 (
		\wishbone_bd_ram_mem3_reg[246][27]/P0001 ,
		_w11952_,
		_w11986_,
		_w17330_
	);
	LUT3 #(
		.INIT('h80)
	) name6818 (
		\wishbone_bd_ram_mem3_reg[0][27]/P0001 ,
		_w11932_,
		_w11941_,
		_w17331_
	);
	LUT4 #(
		.INIT('h0001)
	) name6819 (
		_w17328_,
		_w17329_,
		_w17330_,
		_w17331_,
		_w17332_
	);
	LUT4 #(
		.INIT('h8000)
	) name6820 (
		_w17317_,
		_w17322_,
		_w17327_,
		_w17332_,
		_w17333_
	);
	LUT3 #(
		.INIT('h80)
	) name6821 (
		\wishbone_bd_ram_mem3_reg[156][27]/P0001 ,
		_w11954_,
		_w11959_,
		_w17334_
	);
	LUT3 #(
		.INIT('h80)
	) name6822 (
		\wishbone_bd_ram_mem3_reg[92][27]/P0001 ,
		_w11954_,
		_w11972_,
		_w17335_
	);
	LUT3 #(
		.INIT('h80)
	) name6823 (
		\wishbone_bd_ram_mem3_reg[90][27]/P0001 ,
		_w11944_,
		_w11972_,
		_w17336_
	);
	LUT3 #(
		.INIT('h80)
	) name6824 (
		\wishbone_bd_ram_mem3_reg[231][27]/P0001 ,
		_w11975_,
		_w11982_,
		_w17337_
	);
	LUT4 #(
		.INIT('h0001)
	) name6825 (
		_w17334_,
		_w17335_,
		_w17336_,
		_w17337_,
		_w17338_
	);
	LUT3 #(
		.INIT('h80)
	) name6826 (
		\wishbone_bd_ram_mem3_reg[251][27]/P0001 ,
		_w11936_,
		_w11952_,
		_w17339_
	);
	LUT3 #(
		.INIT('h80)
	) name6827 (
		\wishbone_bd_ram_mem3_reg[235][27]/P0001 ,
		_w11936_,
		_w11982_,
		_w17340_
	);
	LUT3 #(
		.INIT('h80)
	) name6828 (
		\wishbone_bd_ram_mem3_reg[152][27]/P0001 ,
		_w11959_,
		_w11990_,
		_w17341_
	);
	LUT3 #(
		.INIT('h80)
	) name6829 (
		\wishbone_bd_ram_mem3_reg[224][27]/P0001 ,
		_w11941_,
		_w11982_,
		_w17342_
	);
	LUT4 #(
		.INIT('h0001)
	) name6830 (
		_w17339_,
		_w17340_,
		_w17341_,
		_w17342_,
		_w17343_
	);
	LUT3 #(
		.INIT('h80)
	) name6831 (
		\wishbone_bd_ram_mem3_reg[19][27]/P0001 ,
		_w11935_,
		_w11938_,
		_w17344_
	);
	LUT3 #(
		.INIT('h80)
	) name6832 (
		\wishbone_bd_ram_mem3_reg[229][27]/P0001 ,
		_w11933_,
		_w11982_,
		_w17345_
	);
	LUT3 #(
		.INIT('h80)
	) name6833 (
		\wishbone_bd_ram_mem3_reg[196][27]/P0001 ,
		_w11929_,
		_w11945_,
		_w17346_
	);
	LUT3 #(
		.INIT('h80)
	) name6834 (
		\wishbone_bd_ram_mem3_reg[105][27]/P0001 ,
		_w11965_,
		_w11968_,
		_w17347_
	);
	LUT4 #(
		.INIT('h0001)
	) name6835 (
		_w17344_,
		_w17345_,
		_w17346_,
		_w17347_,
		_w17348_
	);
	LUT3 #(
		.INIT('h80)
	) name6836 (
		\wishbone_bd_ram_mem3_reg[82][27]/P0001 ,
		_w11963_,
		_w11972_,
		_w17349_
	);
	LUT3 #(
		.INIT('h80)
	) name6837 (
		\wishbone_bd_ram_mem3_reg[195][27]/P0001 ,
		_w11938_,
		_w11945_,
		_w17350_
	);
	LUT3 #(
		.INIT('h80)
	) name6838 (
		\wishbone_bd_ram_mem3_reg[50][27]/P0001 ,
		_w11963_,
		_w11979_,
		_w17351_
	);
	LUT3 #(
		.INIT('h80)
	) name6839 (
		\wishbone_bd_ram_mem3_reg[185][27]/P0001 ,
		_w11942_,
		_w11968_,
		_w17352_
	);
	LUT4 #(
		.INIT('h0001)
	) name6840 (
		_w17349_,
		_w17350_,
		_w17351_,
		_w17352_,
		_w17353_
	);
	LUT4 #(
		.INIT('h8000)
	) name6841 (
		_w17338_,
		_w17343_,
		_w17348_,
		_w17353_,
		_w17354_
	);
	LUT4 #(
		.INIT('h8000)
	) name6842 (
		_w17291_,
		_w17312_,
		_w17333_,
		_w17354_,
		_w17355_
	);
	LUT4 #(
		.INIT('h8000)
	) name6843 (
		_w17100_,
		_w17185_,
		_w17270_,
		_w17355_,
		_w17356_
	);
	LUT3 #(
		.INIT('hce)
	) name6844 (
		_w12303_,
		_w17015_,
		_w17356_,
		_w17357_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6845 (
		\wishbone_LatchedTxLength_reg[12]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w17358_
	);
	LUT3 #(
		.INIT('hf4)
	) name6846 (
		_w12301_,
		_w12303_,
		_w17358_,
		_w17359_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6847 (
		\wishbone_LatchedTxLength_reg[13]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w17360_
	);
	LUT3 #(
		.INIT('hf2)
	) name6848 (
		_w12303_,
		_w12668_,
		_w17360_,
		_w17361_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6849 (
		\wishbone_LatchedTxLength_reg[14]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w17362_
	);
	LUT3 #(
		.INIT('hf2)
	) name6850 (
		_w12303_,
		_w13016_,
		_w17362_,
		_w17363_
	);
	LUT4 #(
		.INIT('h1555)
	) name6851 (
		\wishbone_LatchedTxLength_reg[15]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w17364_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6852 (
		\wishbone_LatchedTxLength_reg[15]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w17365_
	);
	LUT2 #(
		.INIT('h1)
	) name6853 (
		wb_rst_i_pad,
		_w17364_,
		_w17366_
	);
	LUT3 #(
		.INIT('hdc)
	) name6854 (
		_w16469_,
		_w17365_,
		_w17366_,
		_w17367_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6855 (
		\wishbone_LatchedTxLength_reg[1]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w17368_
	);
	LUT3 #(
		.INIT('hf2)
	) name6856 (
		_w12303_,
		_w16814_,
		_w17368_,
		_w17369_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6857 (
		\wishbone_LatchedTxLength_reg[2]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w17370_
	);
	LUT3 #(
		.INIT('hf2)
	) name6858 (
		_w12303_,
		_w15775_,
		_w17370_,
		_w17371_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6859 (
		\wishbone_LatchedTxLength_reg[3]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w17372_
	);
	LUT3 #(
		.INIT('h80)
	) name6860 (
		\wishbone_bd_ram_mem2_reg[103][19]/P0001 ,
		_w11965_,
		_w11975_,
		_w17373_
	);
	LUT3 #(
		.INIT('h80)
	) name6861 (
		\wishbone_bd_ram_mem2_reg[223][19]/P0001 ,
		_w11973_,
		_w11984_,
		_w17374_
	);
	LUT3 #(
		.INIT('h80)
	) name6862 (
		\wishbone_bd_ram_mem2_reg[203][19]/P0001 ,
		_w11936_,
		_w11945_,
		_w17375_
	);
	LUT3 #(
		.INIT('h80)
	) name6863 (
		\wishbone_bd_ram_mem2_reg[181][19]/P0001 ,
		_w11933_,
		_w11942_,
		_w17376_
	);
	LUT4 #(
		.INIT('h0001)
	) name6864 (
		_w17373_,
		_w17374_,
		_w17375_,
		_w17376_,
		_w17377_
	);
	LUT3 #(
		.INIT('h80)
	) name6865 (
		\wishbone_bd_ram_mem2_reg[73][19]/P0001 ,
		_w11949_,
		_w11968_,
		_w17378_
	);
	LUT3 #(
		.INIT('h80)
	) name6866 (
		\wishbone_bd_ram_mem2_reg[187][19]/P0001 ,
		_w11936_,
		_w11942_,
		_w17379_
	);
	LUT3 #(
		.INIT('h80)
	) name6867 (
		\wishbone_bd_ram_mem2_reg[26][19]/P0001 ,
		_w11935_,
		_w11944_,
		_w17380_
	);
	LUT3 #(
		.INIT('h80)
	) name6868 (
		\wishbone_bd_ram_mem2_reg[67][19]/P0001 ,
		_w11938_,
		_w11949_,
		_w17381_
	);
	LUT4 #(
		.INIT('h0001)
	) name6869 (
		_w17378_,
		_w17379_,
		_w17380_,
		_w17381_,
		_w17382_
	);
	LUT3 #(
		.INIT('h80)
	) name6870 (
		\wishbone_bd_ram_mem2_reg[193][19]/P0001 ,
		_w11945_,
		_w11977_,
		_w17383_
	);
	LUT3 #(
		.INIT('h80)
	) name6871 (
		\wishbone_bd_ram_mem2_reg[42][19]/P0001 ,
		_w11944_,
		_w11957_,
		_w17384_
	);
	LUT3 #(
		.INIT('h80)
	) name6872 (
		\wishbone_bd_ram_mem2_reg[106][19]/P0001 ,
		_w11944_,
		_w11965_,
		_w17385_
	);
	LUT3 #(
		.INIT('h80)
	) name6873 (
		\wishbone_bd_ram_mem2_reg[15][19]/P0001 ,
		_w11932_,
		_w11973_,
		_w17386_
	);
	LUT4 #(
		.INIT('h0001)
	) name6874 (
		_w17383_,
		_w17384_,
		_w17385_,
		_w17386_,
		_w17387_
	);
	LUT3 #(
		.INIT('h80)
	) name6875 (
		\wishbone_bd_ram_mem2_reg[249][19]/P0001 ,
		_w11952_,
		_w11968_,
		_w17388_
	);
	LUT3 #(
		.INIT('h80)
	) name6876 (
		\wishbone_bd_ram_mem2_reg[32][19]/P0001 ,
		_w11941_,
		_w11957_,
		_w17389_
	);
	LUT3 #(
		.INIT('h80)
	) name6877 (
		\wishbone_bd_ram_mem2_reg[136][19]/P0001 ,
		_w11955_,
		_w11990_,
		_w17390_
	);
	LUT3 #(
		.INIT('h80)
	) name6878 (
		\wishbone_bd_ram_mem2_reg[118][19]/P0001 ,
		_w11986_,
		_w12012_,
		_w17391_
	);
	LUT4 #(
		.INIT('h0001)
	) name6879 (
		_w17388_,
		_w17389_,
		_w17390_,
		_w17391_,
		_w17392_
	);
	LUT4 #(
		.INIT('h8000)
	) name6880 (
		_w17377_,
		_w17382_,
		_w17387_,
		_w17392_,
		_w17393_
	);
	LUT3 #(
		.INIT('h80)
	) name6881 (
		\wishbone_bd_ram_mem2_reg[164][19]/P0001 ,
		_w11929_,
		_w11930_,
		_w17394_
	);
	LUT3 #(
		.INIT('h80)
	) name6882 (
		\wishbone_bd_ram_mem2_reg[56][19]/P0001 ,
		_w11979_,
		_w11990_,
		_w17395_
	);
	LUT3 #(
		.INIT('h80)
	) name6883 (
		\wishbone_bd_ram_mem2_reg[108][19]/P0001 ,
		_w11954_,
		_w11965_,
		_w17396_
	);
	LUT3 #(
		.INIT('h80)
	) name6884 (
		\wishbone_bd_ram_mem2_reg[217][19]/P0001 ,
		_w11968_,
		_w11984_,
		_w17397_
	);
	LUT4 #(
		.INIT('h0001)
	) name6885 (
		_w17394_,
		_w17395_,
		_w17396_,
		_w17397_,
		_w17398_
	);
	LUT3 #(
		.INIT('h80)
	) name6886 (
		\wishbone_bd_ram_mem2_reg[11][19]/P0001 ,
		_w11932_,
		_w11936_,
		_w17399_
	);
	LUT3 #(
		.INIT('h80)
	) name6887 (
		\wishbone_bd_ram_mem2_reg[18][19]/P0001 ,
		_w11935_,
		_w11963_,
		_w17400_
	);
	LUT3 #(
		.INIT('h80)
	) name6888 (
		\wishbone_bd_ram_mem2_reg[237][19]/P0001 ,
		_w11966_,
		_w11982_,
		_w17401_
	);
	LUT3 #(
		.INIT('h80)
	) name6889 (
		\wishbone_bd_ram_mem2_reg[135][19]/P0001 ,
		_w11955_,
		_w11975_,
		_w17402_
	);
	LUT4 #(
		.INIT('h0001)
	) name6890 (
		_w17399_,
		_w17400_,
		_w17401_,
		_w17402_,
		_w17403_
	);
	LUT3 #(
		.INIT('h80)
	) name6891 (
		\wishbone_bd_ram_mem2_reg[37][19]/P0001 ,
		_w11933_,
		_w11957_,
		_w17404_
	);
	LUT3 #(
		.INIT('h80)
	) name6892 (
		\wishbone_bd_ram_mem2_reg[55][19]/P0001 ,
		_w11975_,
		_w11979_,
		_w17405_
	);
	LUT3 #(
		.INIT('h80)
	) name6893 (
		\wishbone_bd_ram_mem2_reg[70][19]/P0001 ,
		_w11949_,
		_w11986_,
		_w17406_
	);
	LUT3 #(
		.INIT('h80)
	) name6894 (
		\wishbone_bd_ram_mem2_reg[170][19]/P0001 ,
		_w11930_,
		_w11944_,
		_w17407_
	);
	LUT4 #(
		.INIT('h0001)
	) name6895 (
		_w17404_,
		_w17405_,
		_w17406_,
		_w17407_,
		_w17408_
	);
	LUT3 #(
		.INIT('h80)
	) name6896 (
		\wishbone_bd_ram_mem2_reg[104][19]/P0001 ,
		_w11965_,
		_w11990_,
		_w17409_
	);
	LUT3 #(
		.INIT('h80)
	) name6897 (
		\wishbone_bd_ram_mem2_reg[156][19]/P0001 ,
		_w11954_,
		_w11959_,
		_w17410_
	);
	LUT3 #(
		.INIT('h80)
	) name6898 (
		\wishbone_bd_ram_mem2_reg[61][19]/P0001 ,
		_w11966_,
		_w11979_,
		_w17411_
	);
	LUT3 #(
		.INIT('h80)
	) name6899 (
		\wishbone_bd_ram_mem2_reg[109][19]/P0001 ,
		_w11965_,
		_w11966_,
		_w17412_
	);
	LUT4 #(
		.INIT('h0001)
	) name6900 (
		_w17409_,
		_w17410_,
		_w17411_,
		_w17412_,
		_w17413_
	);
	LUT4 #(
		.INIT('h8000)
	) name6901 (
		_w17398_,
		_w17403_,
		_w17408_,
		_w17413_,
		_w17414_
	);
	LUT3 #(
		.INIT('h80)
	) name6902 (
		\wishbone_bd_ram_mem2_reg[79][19]/P0001 ,
		_w11949_,
		_w11973_,
		_w17415_
	);
	LUT3 #(
		.INIT('h80)
	) name6903 (
		\wishbone_bd_ram_mem2_reg[91][19]/P0001 ,
		_w11936_,
		_w11972_,
		_w17416_
	);
	LUT3 #(
		.INIT('h80)
	) name6904 (
		\wishbone_bd_ram_mem2_reg[147][19]/P0001 ,
		_w11938_,
		_w11959_,
		_w17417_
	);
	LUT3 #(
		.INIT('h80)
	) name6905 (
		\wishbone_bd_ram_mem2_reg[113][19]/P0001 ,
		_w11977_,
		_w12012_,
		_w17418_
	);
	LUT4 #(
		.INIT('h0001)
	) name6906 (
		_w17415_,
		_w17416_,
		_w17417_,
		_w17418_,
		_w17419_
	);
	LUT3 #(
		.INIT('h80)
	) name6907 (
		\wishbone_bd_ram_mem2_reg[160][19]/P0001 ,
		_w11930_,
		_w11941_,
		_w17420_
	);
	LUT3 #(
		.INIT('h80)
	) name6908 (
		\wishbone_bd_ram_mem2_reg[148][19]/P0001 ,
		_w11929_,
		_w11959_,
		_w17421_
	);
	LUT3 #(
		.INIT('h80)
	) name6909 (
		\wishbone_bd_ram_mem2_reg[23][19]/P0001 ,
		_w11935_,
		_w11975_,
		_w17422_
	);
	LUT3 #(
		.INIT('h80)
	) name6910 (
		\wishbone_bd_ram_mem2_reg[131][19]/P0001 ,
		_w11938_,
		_w11955_,
		_w17423_
	);
	LUT4 #(
		.INIT('h0001)
	) name6911 (
		_w17420_,
		_w17421_,
		_w17422_,
		_w17423_,
		_w17424_
	);
	LUT3 #(
		.INIT('h80)
	) name6912 (
		\wishbone_bd_ram_mem2_reg[52][19]/P0001 ,
		_w11929_,
		_w11979_,
		_w17425_
	);
	LUT3 #(
		.INIT('h80)
	) name6913 (
		\wishbone_bd_ram_mem2_reg[190][19]/P0001 ,
		_w11942_,
		_w11948_,
		_w17426_
	);
	LUT3 #(
		.INIT('h80)
	) name6914 (
		\wishbone_bd_ram_mem2_reg[222][19]/P0001 ,
		_w11948_,
		_w11984_,
		_w17427_
	);
	LUT3 #(
		.INIT('h80)
	) name6915 (
		\wishbone_bd_ram_mem2_reg[122][19]/P0001 ,
		_w11944_,
		_w12012_,
		_w17428_
	);
	LUT4 #(
		.INIT('h0001)
	) name6916 (
		_w17425_,
		_w17426_,
		_w17427_,
		_w17428_,
		_w17429_
	);
	LUT3 #(
		.INIT('h80)
	) name6917 (
		\wishbone_bd_ram_mem2_reg[10][19]/P0001 ,
		_w11932_,
		_w11944_,
		_w17430_
	);
	LUT3 #(
		.INIT('h80)
	) name6918 (
		\wishbone_bd_ram_mem2_reg[74][19]/P0001 ,
		_w11944_,
		_w11949_,
		_w17431_
	);
	LUT3 #(
		.INIT('h80)
	) name6919 (
		\wishbone_bd_ram_mem2_reg[230][19]/P0001 ,
		_w11982_,
		_w11986_,
		_w17432_
	);
	LUT3 #(
		.INIT('h80)
	) name6920 (
		\wishbone_bd_ram_mem2_reg[6][19]/P0001 ,
		_w11932_,
		_w11986_,
		_w17433_
	);
	LUT4 #(
		.INIT('h0001)
	) name6921 (
		_w17430_,
		_w17431_,
		_w17432_,
		_w17433_,
		_w17434_
	);
	LUT4 #(
		.INIT('h8000)
	) name6922 (
		_w17419_,
		_w17424_,
		_w17429_,
		_w17434_,
		_w17435_
	);
	LUT3 #(
		.INIT('h80)
	) name6923 (
		\wishbone_bd_ram_mem2_reg[172][19]/P0001 ,
		_w11930_,
		_w11954_,
		_w17436_
	);
	LUT3 #(
		.INIT('h80)
	) name6924 (
		\wishbone_bd_ram_mem2_reg[212][19]/P0001 ,
		_w11929_,
		_w11984_,
		_w17437_
	);
	LUT3 #(
		.INIT('h80)
	) name6925 (
		\wishbone_bd_ram_mem2_reg[157][19]/P0001 ,
		_w11959_,
		_w11966_,
		_w17438_
	);
	LUT3 #(
		.INIT('h80)
	) name6926 (
		\wishbone_bd_ram_mem2_reg[183][19]/P0001 ,
		_w11942_,
		_w11975_,
		_w17439_
	);
	LUT4 #(
		.INIT('h0001)
	) name6927 (
		_w17436_,
		_w17437_,
		_w17438_,
		_w17439_,
		_w17440_
	);
	LUT3 #(
		.INIT('h80)
	) name6928 (
		\wishbone_bd_ram_mem2_reg[134][19]/P0001 ,
		_w11955_,
		_w11986_,
		_w17441_
	);
	LUT3 #(
		.INIT('h80)
	) name6929 (
		\wishbone_bd_ram_mem2_reg[62][19]/P0001 ,
		_w11948_,
		_w11979_,
		_w17442_
	);
	LUT3 #(
		.INIT('h80)
	) name6930 (
		\wishbone_bd_ram_mem2_reg[102][19]/P0001 ,
		_w11965_,
		_w11986_,
		_w17443_
	);
	LUT3 #(
		.INIT('h80)
	) name6931 (
		\wishbone_bd_ram_mem2_reg[126][19]/P0001 ,
		_w11948_,
		_w12012_,
		_w17444_
	);
	LUT4 #(
		.INIT('h0001)
	) name6932 (
		_w17441_,
		_w17442_,
		_w17443_,
		_w17444_,
		_w17445_
	);
	LUT3 #(
		.INIT('h80)
	) name6933 (
		\wishbone_bd_ram_mem2_reg[252][19]/P0001 ,
		_w11952_,
		_w11954_,
		_w17446_
	);
	LUT3 #(
		.INIT('h80)
	) name6934 (
		\wishbone_bd_ram_mem2_reg[21][19]/P0001 ,
		_w11933_,
		_w11935_,
		_w17447_
	);
	LUT3 #(
		.INIT('h80)
	) name6935 (
		\wishbone_bd_ram_mem2_reg[225][19]/P0001 ,
		_w11977_,
		_w11982_,
		_w17448_
	);
	LUT3 #(
		.INIT('h80)
	) name6936 (
		\wishbone_bd_ram_mem2_reg[205][19]/P0001 ,
		_w11945_,
		_w11966_,
		_w17449_
	);
	LUT4 #(
		.INIT('h0001)
	) name6937 (
		_w17446_,
		_w17447_,
		_w17448_,
		_w17449_,
		_w17450_
	);
	LUT3 #(
		.INIT('h80)
	) name6938 (
		\wishbone_bd_ram_mem2_reg[206][19]/P0001 ,
		_w11945_,
		_w11948_,
		_w17451_
	);
	LUT3 #(
		.INIT('h80)
	) name6939 (
		\wishbone_bd_ram_mem2_reg[215][19]/P0001 ,
		_w11975_,
		_w11984_,
		_w17452_
	);
	LUT3 #(
		.INIT('h80)
	) name6940 (
		\wishbone_bd_ram_mem2_reg[114][19]/P0001 ,
		_w11963_,
		_w12012_,
		_w17453_
	);
	LUT3 #(
		.INIT('h80)
	) name6941 (
		\wishbone_bd_ram_mem2_reg[119][19]/P0001 ,
		_w11975_,
		_w12012_,
		_w17454_
	);
	LUT4 #(
		.INIT('h0001)
	) name6942 (
		_w17451_,
		_w17452_,
		_w17453_,
		_w17454_,
		_w17455_
	);
	LUT4 #(
		.INIT('h8000)
	) name6943 (
		_w17440_,
		_w17445_,
		_w17450_,
		_w17455_,
		_w17456_
	);
	LUT4 #(
		.INIT('h8000)
	) name6944 (
		_w17393_,
		_w17414_,
		_w17435_,
		_w17456_,
		_w17457_
	);
	LUT3 #(
		.INIT('h80)
	) name6945 (
		\wishbone_bd_ram_mem2_reg[151][19]/P0001 ,
		_w11959_,
		_w11975_,
		_w17458_
	);
	LUT3 #(
		.INIT('h80)
	) name6946 (
		\wishbone_bd_ram_mem2_reg[92][19]/P0001 ,
		_w11954_,
		_w11972_,
		_w17459_
	);
	LUT3 #(
		.INIT('h80)
	) name6947 (
		\wishbone_bd_ram_mem2_reg[144][19]/P0001 ,
		_w11941_,
		_w11959_,
		_w17460_
	);
	LUT3 #(
		.INIT('h80)
	) name6948 (
		\wishbone_bd_ram_mem2_reg[5][19]/P0001 ,
		_w11932_,
		_w11933_,
		_w17461_
	);
	LUT4 #(
		.INIT('h0001)
	) name6949 (
		_w17458_,
		_w17459_,
		_w17460_,
		_w17461_,
		_w17462_
	);
	LUT3 #(
		.INIT('h80)
	) name6950 (
		\wishbone_bd_ram_mem2_reg[69][19]/P0001 ,
		_w11933_,
		_w11949_,
		_w17463_
	);
	LUT3 #(
		.INIT('h80)
	) name6951 (
		\wishbone_bd_ram_mem2_reg[87][19]/P0001 ,
		_w11972_,
		_w11975_,
		_w17464_
	);
	LUT3 #(
		.INIT('h80)
	) name6952 (
		\wishbone_bd_ram_mem2_reg[85][19]/P0001 ,
		_w11933_,
		_w11972_,
		_w17465_
	);
	LUT3 #(
		.INIT('h80)
	) name6953 (
		\wishbone_bd_ram_mem2_reg[235][19]/P0001 ,
		_w11936_,
		_w11982_,
		_w17466_
	);
	LUT4 #(
		.INIT('h0001)
	) name6954 (
		_w17463_,
		_w17464_,
		_w17465_,
		_w17466_,
		_w17467_
	);
	LUT3 #(
		.INIT('h80)
	) name6955 (
		\wishbone_bd_ram_mem2_reg[207][19]/P0001 ,
		_w11945_,
		_w11973_,
		_w17468_
	);
	LUT3 #(
		.INIT('h80)
	) name6956 (
		\wishbone_bd_ram_mem2_reg[132][19]/P0001 ,
		_w11929_,
		_w11955_,
		_w17469_
	);
	LUT3 #(
		.INIT('h80)
	) name6957 (
		\wishbone_bd_ram_mem2_reg[159][19]/P0001 ,
		_w11959_,
		_w11973_,
		_w17470_
	);
	LUT3 #(
		.INIT('h80)
	) name6958 (
		\wishbone_bd_ram_mem2_reg[16][19]/P0001 ,
		_w11935_,
		_w11941_,
		_w17471_
	);
	LUT4 #(
		.INIT('h0001)
	) name6959 (
		_w17468_,
		_w17469_,
		_w17470_,
		_w17471_,
		_w17472_
	);
	LUT3 #(
		.INIT('h80)
	) name6960 (
		\wishbone_bd_ram_mem2_reg[150][19]/P0001 ,
		_w11959_,
		_w11986_,
		_w17473_
	);
	LUT3 #(
		.INIT('h80)
	) name6961 (
		\wishbone_bd_ram_mem2_reg[143][19]/P0001 ,
		_w11955_,
		_w11973_,
		_w17474_
	);
	LUT3 #(
		.INIT('h80)
	) name6962 (
		\wishbone_bd_ram_mem2_reg[3][19]/P0001 ,
		_w11932_,
		_w11938_,
		_w17475_
	);
	LUT3 #(
		.INIT('h80)
	) name6963 (
		\wishbone_bd_ram_mem2_reg[227][19]/P0001 ,
		_w11938_,
		_w11982_,
		_w17476_
	);
	LUT4 #(
		.INIT('h0001)
	) name6964 (
		_w17473_,
		_w17474_,
		_w17475_,
		_w17476_,
		_w17477_
	);
	LUT4 #(
		.INIT('h8000)
	) name6965 (
		_w17462_,
		_w17467_,
		_w17472_,
		_w17477_,
		_w17478_
	);
	LUT3 #(
		.INIT('h80)
	) name6966 (
		\wishbone_bd_ram_mem2_reg[89][19]/P0001 ,
		_w11968_,
		_w11972_,
		_w17479_
	);
	LUT3 #(
		.INIT('h80)
	) name6967 (
		\wishbone_bd_ram_mem2_reg[72][19]/P0001 ,
		_w11949_,
		_w11990_,
		_w17480_
	);
	LUT3 #(
		.INIT('h80)
	) name6968 (
		\wishbone_bd_ram_mem2_reg[180][19]/P0001 ,
		_w11929_,
		_w11942_,
		_w17481_
	);
	LUT3 #(
		.INIT('h80)
	) name6969 (
		\wishbone_bd_ram_mem2_reg[248][19]/P0001 ,
		_w11952_,
		_w11990_,
		_w17482_
	);
	LUT4 #(
		.INIT('h0001)
	) name6970 (
		_w17479_,
		_w17480_,
		_w17481_,
		_w17482_,
		_w17483_
	);
	LUT3 #(
		.INIT('h80)
	) name6971 (
		\wishbone_bd_ram_mem2_reg[96][19]/P0001 ,
		_w11941_,
		_w11965_,
		_w17484_
	);
	LUT3 #(
		.INIT('h80)
	) name6972 (
		\wishbone_bd_ram_mem2_reg[121][19]/P0001 ,
		_w11968_,
		_w12012_,
		_w17485_
	);
	LUT3 #(
		.INIT('h80)
	) name6973 (
		\wishbone_bd_ram_mem2_reg[191][19]/P0001 ,
		_w11942_,
		_w11973_,
		_w17486_
	);
	LUT3 #(
		.INIT('h80)
	) name6974 (
		\wishbone_bd_ram_mem2_reg[98][19]/P0001 ,
		_w11963_,
		_w11965_,
		_w17487_
	);
	LUT4 #(
		.INIT('h0001)
	) name6975 (
		_w17484_,
		_w17485_,
		_w17486_,
		_w17487_,
		_w17488_
	);
	LUT3 #(
		.INIT('h80)
	) name6976 (
		\wishbone_bd_ram_mem2_reg[107][19]/P0001 ,
		_w11936_,
		_w11965_,
		_w17489_
	);
	LUT3 #(
		.INIT('h80)
	) name6977 (
		\wishbone_bd_ram_mem2_reg[54][19]/P0001 ,
		_w11979_,
		_w11986_,
		_w17490_
	);
	LUT3 #(
		.INIT('h80)
	) name6978 (
		\wishbone_bd_ram_mem2_reg[64][19]/P0001 ,
		_w11941_,
		_w11949_,
		_w17491_
	);
	LUT3 #(
		.INIT('h80)
	) name6979 (
		\wishbone_bd_ram_mem2_reg[158][19]/P0001 ,
		_w11948_,
		_w11959_,
		_w17492_
	);
	LUT4 #(
		.INIT('h0001)
	) name6980 (
		_w17489_,
		_w17490_,
		_w17491_,
		_w17492_,
		_w17493_
	);
	LUT3 #(
		.INIT('h80)
	) name6981 (
		\wishbone_bd_ram_mem2_reg[161][19]/P0001 ,
		_w11930_,
		_w11977_,
		_w17494_
	);
	LUT3 #(
		.INIT('h80)
	) name6982 (
		\wishbone_bd_ram_mem2_reg[31][19]/P0001 ,
		_w11935_,
		_w11973_,
		_w17495_
	);
	LUT3 #(
		.INIT('h80)
	) name6983 (
		\wishbone_bd_ram_mem2_reg[27][19]/P0001 ,
		_w11935_,
		_w11936_,
		_w17496_
	);
	LUT3 #(
		.INIT('h80)
	) name6984 (
		\wishbone_bd_ram_mem2_reg[210][19]/P0001 ,
		_w11963_,
		_w11984_,
		_w17497_
	);
	LUT4 #(
		.INIT('h0001)
	) name6985 (
		_w17494_,
		_w17495_,
		_w17496_,
		_w17497_,
		_w17498_
	);
	LUT4 #(
		.INIT('h8000)
	) name6986 (
		_w17483_,
		_w17488_,
		_w17493_,
		_w17498_,
		_w17499_
	);
	LUT3 #(
		.INIT('h80)
	) name6987 (
		\wishbone_bd_ram_mem2_reg[176][19]/P0001 ,
		_w11941_,
		_w11942_,
		_w17500_
	);
	LUT3 #(
		.INIT('h80)
	) name6988 (
		\wishbone_bd_ram_mem2_reg[208][19]/P0001 ,
		_w11941_,
		_w11984_,
		_w17501_
	);
	LUT3 #(
		.INIT('h80)
	) name6989 (
		\wishbone_bd_ram_mem2_reg[77][19]/P0001 ,
		_w11949_,
		_w11966_,
		_w17502_
	);
	LUT3 #(
		.INIT('h80)
	) name6990 (
		\wishbone_bd_ram_mem2_reg[182][19]/P0001 ,
		_w11942_,
		_w11986_,
		_w17503_
	);
	LUT4 #(
		.INIT('h0001)
	) name6991 (
		_w17500_,
		_w17501_,
		_w17502_,
		_w17503_,
		_w17504_
	);
	LUT3 #(
		.INIT('h80)
	) name6992 (
		\wishbone_bd_ram_mem2_reg[30][19]/P0001 ,
		_w11935_,
		_w11948_,
		_w17505_
	);
	LUT3 #(
		.INIT('h80)
	) name6993 (
		\wishbone_bd_ram_mem2_reg[36][19]/P0001 ,
		_w11929_,
		_w11957_,
		_w17506_
	);
	LUT3 #(
		.INIT('h80)
	) name6994 (
		\wishbone_bd_ram_mem2_reg[130][19]/P0001 ,
		_w11955_,
		_w11963_,
		_w17507_
	);
	LUT3 #(
		.INIT('h80)
	) name6995 (
		\wishbone_bd_ram_mem2_reg[236][19]/P0001 ,
		_w11954_,
		_w11982_,
		_w17508_
	);
	LUT4 #(
		.INIT('h0001)
	) name6996 (
		_w17505_,
		_w17506_,
		_w17507_,
		_w17508_,
		_w17509_
	);
	LUT3 #(
		.INIT('h80)
	) name6997 (
		\wishbone_bd_ram_mem2_reg[14][19]/P0001 ,
		_w11932_,
		_w11948_,
		_w17510_
	);
	LUT3 #(
		.INIT('h80)
	) name6998 (
		\wishbone_bd_ram_mem2_reg[38][19]/P0001 ,
		_w11957_,
		_w11986_,
		_w17511_
	);
	LUT3 #(
		.INIT('h80)
	) name6999 (
		\wishbone_bd_ram_mem2_reg[138][19]/P0001 ,
		_w11944_,
		_w11955_,
		_w17512_
	);
	LUT3 #(
		.INIT('h80)
	) name7000 (
		\wishbone_bd_ram_mem2_reg[13][19]/P0001 ,
		_w11932_,
		_w11966_,
		_w17513_
	);
	LUT4 #(
		.INIT('h0001)
	) name7001 (
		_w17510_,
		_w17511_,
		_w17512_,
		_w17513_,
		_w17514_
	);
	LUT3 #(
		.INIT('h80)
	) name7002 (
		\wishbone_bd_ram_mem2_reg[49][19]/P0001 ,
		_w11977_,
		_w11979_,
		_w17515_
	);
	LUT3 #(
		.INIT('h80)
	) name7003 (
		\wishbone_bd_ram_mem2_reg[7][19]/P0001 ,
		_w11932_,
		_w11975_,
		_w17516_
	);
	LUT3 #(
		.INIT('h80)
	) name7004 (
		\wishbone_bd_ram_mem2_reg[219][19]/P0001 ,
		_w11936_,
		_w11984_,
		_w17517_
	);
	LUT3 #(
		.INIT('h80)
	) name7005 (
		\wishbone_bd_ram_mem2_reg[245][19]/P0001 ,
		_w11933_,
		_w11952_,
		_w17518_
	);
	LUT4 #(
		.INIT('h0001)
	) name7006 (
		_w17515_,
		_w17516_,
		_w17517_,
		_w17518_,
		_w17519_
	);
	LUT4 #(
		.INIT('h8000)
	) name7007 (
		_w17504_,
		_w17509_,
		_w17514_,
		_w17519_,
		_w17520_
	);
	LUT3 #(
		.INIT('h80)
	) name7008 (
		\wishbone_bd_ram_mem2_reg[39][19]/P0001 ,
		_w11957_,
		_w11975_,
		_w17521_
	);
	LUT3 #(
		.INIT('h80)
	) name7009 (
		\wishbone_bd_ram_mem2_reg[63][19]/P0001 ,
		_w11973_,
		_w11979_,
		_w17522_
	);
	LUT3 #(
		.INIT('h80)
	) name7010 (
		\wishbone_bd_ram_mem2_reg[129][19]/P0001 ,
		_w11955_,
		_w11977_,
		_w17523_
	);
	LUT3 #(
		.INIT('h80)
	) name7011 (
		\wishbone_bd_ram_mem2_reg[201][19]/P0001 ,
		_w11945_,
		_w11968_,
		_w17524_
	);
	LUT4 #(
		.INIT('h0001)
	) name7012 (
		_w17521_,
		_w17522_,
		_w17523_,
		_w17524_,
		_w17525_
	);
	LUT3 #(
		.INIT('h80)
	) name7013 (
		\wishbone_bd_ram_mem2_reg[124][19]/P0001 ,
		_w11954_,
		_w12012_,
		_w17526_
	);
	LUT3 #(
		.INIT('h80)
	) name7014 (
		\wishbone_bd_ram_mem2_reg[28][19]/P0001 ,
		_w11935_,
		_w11954_,
		_w17527_
	);
	LUT3 #(
		.INIT('h80)
	) name7015 (
		\wishbone_bd_ram_mem2_reg[228][19]/P0001 ,
		_w11929_,
		_w11982_,
		_w17528_
	);
	LUT3 #(
		.INIT('h80)
	) name7016 (
		\wishbone_bd_ram_mem2_reg[100][19]/P0001 ,
		_w11929_,
		_w11965_,
		_w17529_
	);
	LUT4 #(
		.INIT('h0001)
	) name7017 (
		_w17526_,
		_w17527_,
		_w17528_,
		_w17529_,
		_w17530_
	);
	LUT3 #(
		.INIT('h80)
	) name7018 (
		\wishbone_bd_ram_mem2_reg[80][19]/P0001 ,
		_w11941_,
		_w11972_,
		_w17531_
	);
	LUT3 #(
		.INIT('h80)
	) name7019 (
		\wishbone_bd_ram_mem2_reg[169][19]/P0001 ,
		_w11930_,
		_w11968_,
		_w17532_
	);
	LUT3 #(
		.INIT('h80)
	) name7020 (
		\wishbone_bd_ram_mem2_reg[229][19]/P0001 ,
		_w11933_,
		_w11982_,
		_w17533_
	);
	LUT3 #(
		.INIT('h80)
	) name7021 (
		\wishbone_bd_ram_mem2_reg[25][19]/P0001 ,
		_w11935_,
		_w11968_,
		_w17534_
	);
	LUT4 #(
		.INIT('h0001)
	) name7022 (
		_w17531_,
		_w17532_,
		_w17533_,
		_w17534_,
		_w17535_
	);
	LUT3 #(
		.INIT('h80)
	) name7023 (
		\wishbone_bd_ram_mem2_reg[20][19]/P0001 ,
		_w11929_,
		_w11935_,
		_w17536_
	);
	LUT3 #(
		.INIT('h80)
	) name7024 (
		\wishbone_bd_ram_mem2_reg[163][19]/P0001 ,
		_w11930_,
		_w11938_,
		_w17537_
	);
	LUT3 #(
		.INIT('h80)
	) name7025 (
		\wishbone_bd_ram_mem2_reg[242][19]/P0001 ,
		_w11952_,
		_w11963_,
		_w17538_
	);
	LUT3 #(
		.INIT('h80)
	) name7026 (
		\wishbone_bd_ram_mem2_reg[60][19]/P0001 ,
		_w11954_,
		_w11979_,
		_w17539_
	);
	LUT4 #(
		.INIT('h0001)
	) name7027 (
		_w17536_,
		_w17537_,
		_w17538_,
		_w17539_,
		_w17540_
	);
	LUT4 #(
		.INIT('h8000)
	) name7028 (
		_w17525_,
		_w17530_,
		_w17535_,
		_w17540_,
		_w17541_
	);
	LUT4 #(
		.INIT('h8000)
	) name7029 (
		_w17478_,
		_w17499_,
		_w17520_,
		_w17541_,
		_w17542_
	);
	LUT3 #(
		.INIT('h80)
	) name7030 (
		\wishbone_bd_ram_mem2_reg[224][19]/P0001 ,
		_w11941_,
		_w11982_,
		_w17543_
	);
	LUT3 #(
		.INIT('h80)
	) name7031 (
		\wishbone_bd_ram_mem2_reg[174][19]/P0001 ,
		_w11930_,
		_w11948_,
		_w17544_
	);
	LUT3 #(
		.INIT('h80)
	) name7032 (
		\wishbone_bd_ram_mem2_reg[202][19]/P0001 ,
		_w11944_,
		_w11945_,
		_w17545_
	);
	LUT3 #(
		.INIT('h80)
	) name7033 (
		\wishbone_bd_ram_mem2_reg[22][19]/P0001 ,
		_w11935_,
		_w11986_,
		_w17546_
	);
	LUT4 #(
		.INIT('h0001)
	) name7034 (
		_w17543_,
		_w17544_,
		_w17545_,
		_w17546_,
		_w17547_
	);
	LUT3 #(
		.INIT('h80)
	) name7035 (
		\wishbone_bd_ram_mem2_reg[189][19]/P0001 ,
		_w11942_,
		_w11966_,
		_w17548_
	);
	LUT3 #(
		.INIT('h80)
	) name7036 (
		\wishbone_bd_ram_mem2_reg[171][19]/P0001 ,
		_w11930_,
		_w11936_,
		_w17549_
	);
	LUT3 #(
		.INIT('h80)
	) name7037 (
		\wishbone_bd_ram_mem2_reg[188][19]/P0001 ,
		_w11942_,
		_w11954_,
		_w17550_
	);
	LUT3 #(
		.INIT('h80)
	) name7038 (
		\wishbone_bd_ram_mem2_reg[45][19]/P0001 ,
		_w11957_,
		_w11966_,
		_w17551_
	);
	LUT4 #(
		.INIT('h0001)
	) name7039 (
		_w17548_,
		_w17549_,
		_w17550_,
		_w17551_,
		_w17552_
	);
	LUT3 #(
		.INIT('h80)
	) name7040 (
		\wishbone_bd_ram_mem2_reg[149][19]/P0001 ,
		_w11933_,
		_w11959_,
		_w17553_
	);
	LUT3 #(
		.INIT('h80)
	) name7041 (
		\wishbone_bd_ram_mem2_reg[200][19]/P0001 ,
		_w11945_,
		_w11990_,
		_w17554_
	);
	LUT3 #(
		.INIT('h80)
	) name7042 (
		\wishbone_bd_ram_mem2_reg[50][19]/P0001 ,
		_w11963_,
		_w11979_,
		_w17555_
	);
	LUT3 #(
		.INIT('h80)
	) name7043 (
		\wishbone_bd_ram_mem2_reg[152][19]/P0001 ,
		_w11959_,
		_w11990_,
		_w17556_
	);
	LUT4 #(
		.INIT('h0001)
	) name7044 (
		_w17553_,
		_w17554_,
		_w17555_,
		_w17556_,
		_w17557_
	);
	LUT3 #(
		.INIT('h80)
	) name7045 (
		\wishbone_bd_ram_mem2_reg[120][19]/P0001 ,
		_w11990_,
		_w12012_,
		_w17558_
	);
	LUT3 #(
		.INIT('h80)
	) name7046 (
		\wishbone_bd_ram_mem2_reg[185][19]/P0001 ,
		_w11942_,
		_w11968_,
		_w17559_
	);
	LUT3 #(
		.INIT('h80)
	) name7047 (
		\wishbone_bd_ram_mem2_reg[101][19]/P0001 ,
		_w11933_,
		_w11965_,
		_w17560_
	);
	LUT3 #(
		.INIT('h80)
	) name7048 (
		\wishbone_bd_ram_mem2_reg[241][19]/P0001 ,
		_w11952_,
		_w11977_,
		_w17561_
	);
	LUT4 #(
		.INIT('h0001)
	) name7049 (
		_w17558_,
		_w17559_,
		_w17560_,
		_w17561_,
		_w17562_
	);
	LUT4 #(
		.INIT('h8000)
	) name7050 (
		_w17547_,
		_w17552_,
		_w17557_,
		_w17562_,
		_w17563_
	);
	LUT3 #(
		.INIT('h80)
	) name7051 (
		\wishbone_bd_ram_mem2_reg[115][19]/P0001 ,
		_w11938_,
		_w12012_,
		_w17564_
	);
	LUT3 #(
		.INIT('h80)
	) name7052 (
		\wishbone_bd_ram_mem2_reg[192][19]/P0001 ,
		_w11941_,
		_w11945_,
		_w17565_
	);
	LUT3 #(
		.INIT('h80)
	) name7053 (
		\wishbone_bd_ram_mem2_reg[197][19]/P0001 ,
		_w11933_,
		_w11945_,
		_w17566_
	);
	LUT3 #(
		.INIT('h80)
	) name7054 (
		\wishbone_bd_ram_mem2_reg[12][19]/P0001 ,
		_w11932_,
		_w11954_,
		_w17567_
	);
	LUT4 #(
		.INIT('h0001)
	) name7055 (
		_w17564_,
		_w17565_,
		_w17566_,
		_w17567_,
		_w17568_
	);
	LUT3 #(
		.INIT('h80)
	) name7056 (
		\wishbone_bd_ram_mem2_reg[46][19]/P0001 ,
		_w11948_,
		_w11957_,
		_w17569_
	);
	LUT3 #(
		.INIT('h80)
	) name7057 (
		\wishbone_bd_ram_mem2_reg[19][19]/P0001 ,
		_w11935_,
		_w11938_,
		_w17570_
	);
	LUT3 #(
		.INIT('h80)
	) name7058 (
		\wishbone_bd_ram_mem2_reg[165][19]/P0001 ,
		_w11930_,
		_w11933_,
		_w17571_
	);
	LUT3 #(
		.INIT('h80)
	) name7059 (
		\wishbone_bd_ram_mem2_reg[218][19]/P0001 ,
		_w11944_,
		_w11984_,
		_w17572_
	);
	LUT4 #(
		.INIT('h0001)
	) name7060 (
		_w17569_,
		_w17570_,
		_w17571_,
		_w17572_,
		_w17573_
	);
	LUT3 #(
		.INIT('h80)
	) name7061 (
		\wishbone_bd_ram_mem2_reg[146][19]/P0001 ,
		_w11959_,
		_w11963_,
		_w17574_
	);
	LUT3 #(
		.INIT('h80)
	) name7062 (
		\wishbone_bd_ram_mem2_reg[179][19]/P0001 ,
		_w11938_,
		_w11942_,
		_w17575_
	);
	LUT3 #(
		.INIT('h80)
	) name7063 (
		\wishbone_bd_ram_mem2_reg[162][19]/P0001 ,
		_w11930_,
		_w11963_,
		_w17576_
	);
	LUT3 #(
		.INIT('h80)
	) name7064 (
		\wishbone_bd_ram_mem2_reg[105][19]/P0001 ,
		_w11965_,
		_w11968_,
		_w17577_
	);
	LUT4 #(
		.INIT('h0001)
	) name7065 (
		_w17574_,
		_w17575_,
		_w17576_,
		_w17577_,
		_w17578_
	);
	LUT3 #(
		.INIT('h80)
	) name7066 (
		\wishbone_bd_ram_mem2_reg[112][19]/P0001 ,
		_w11941_,
		_w12012_,
		_w17579_
	);
	LUT3 #(
		.INIT('h80)
	) name7067 (
		\wishbone_bd_ram_mem2_reg[253][19]/P0001 ,
		_w11952_,
		_w11966_,
		_w17580_
	);
	LUT3 #(
		.INIT('h80)
	) name7068 (
		\wishbone_bd_ram_mem2_reg[226][19]/P0001 ,
		_w11963_,
		_w11982_,
		_w17581_
	);
	LUT3 #(
		.INIT('h80)
	) name7069 (
		\wishbone_bd_ram_mem2_reg[195][19]/P0001 ,
		_w11938_,
		_w11945_,
		_w17582_
	);
	LUT4 #(
		.INIT('h0001)
	) name7070 (
		_w17579_,
		_w17580_,
		_w17581_,
		_w17582_,
		_w17583_
	);
	LUT4 #(
		.INIT('h8000)
	) name7071 (
		_w17568_,
		_w17573_,
		_w17578_,
		_w17583_,
		_w17584_
	);
	LUT3 #(
		.INIT('h80)
	) name7072 (
		\wishbone_bd_ram_mem2_reg[83][19]/P0001 ,
		_w11938_,
		_w11972_,
		_w17585_
	);
	LUT3 #(
		.INIT('h80)
	) name7073 (
		\wishbone_bd_ram_mem2_reg[214][19]/P0001 ,
		_w11984_,
		_w11986_,
		_w17586_
	);
	LUT3 #(
		.INIT('h80)
	) name7074 (
		\wishbone_bd_ram_mem2_reg[220][19]/P0001 ,
		_w11954_,
		_w11984_,
		_w17587_
	);
	LUT3 #(
		.INIT('h80)
	) name7075 (
		\wishbone_bd_ram_mem2_reg[58][19]/P0001 ,
		_w11944_,
		_w11979_,
		_w17588_
	);
	LUT4 #(
		.INIT('h0001)
	) name7076 (
		_w17585_,
		_w17586_,
		_w17587_,
		_w17588_,
		_w17589_
	);
	LUT3 #(
		.INIT('h80)
	) name7077 (
		\wishbone_bd_ram_mem2_reg[51][19]/P0001 ,
		_w11938_,
		_w11979_,
		_w17590_
	);
	LUT3 #(
		.INIT('h80)
	) name7078 (
		\wishbone_bd_ram_mem2_reg[247][19]/P0001 ,
		_w11952_,
		_w11975_,
		_w17591_
	);
	LUT3 #(
		.INIT('h80)
	) name7079 (
		\wishbone_bd_ram_mem2_reg[186][19]/P0001 ,
		_w11942_,
		_w11944_,
		_w17592_
	);
	LUT3 #(
		.INIT('h80)
	) name7080 (
		\wishbone_bd_ram_mem2_reg[233][19]/P0001 ,
		_w11968_,
		_w11982_,
		_w17593_
	);
	LUT4 #(
		.INIT('h0001)
	) name7081 (
		_w17590_,
		_w17591_,
		_w17592_,
		_w17593_,
		_w17594_
	);
	LUT3 #(
		.INIT('h80)
	) name7082 (
		\wishbone_bd_ram_mem2_reg[204][19]/P0001 ,
		_w11945_,
		_w11954_,
		_w17595_
	);
	LUT3 #(
		.INIT('h80)
	) name7083 (
		\wishbone_bd_ram_mem2_reg[213][19]/P0001 ,
		_w11933_,
		_w11984_,
		_w17596_
	);
	LUT3 #(
		.INIT('h80)
	) name7084 (
		\wishbone_bd_ram_mem2_reg[90][19]/P0001 ,
		_w11944_,
		_w11972_,
		_w17597_
	);
	LUT3 #(
		.INIT('h80)
	) name7085 (
		\wishbone_bd_ram_mem2_reg[68][19]/P0001 ,
		_w11929_,
		_w11949_,
		_w17598_
	);
	LUT4 #(
		.INIT('h0001)
	) name7086 (
		_w17595_,
		_w17596_,
		_w17597_,
		_w17598_,
		_w17599_
	);
	LUT3 #(
		.INIT('h80)
	) name7087 (
		\wishbone_bd_ram_mem2_reg[145][19]/P0001 ,
		_w11959_,
		_w11977_,
		_w17600_
	);
	LUT3 #(
		.INIT('h80)
	) name7088 (
		\wishbone_bd_ram_mem2_reg[35][19]/P0001 ,
		_w11938_,
		_w11957_,
		_w17601_
	);
	LUT3 #(
		.INIT('h80)
	) name7089 (
		\wishbone_bd_ram_mem2_reg[94][19]/P0001 ,
		_w11948_,
		_w11972_,
		_w17602_
	);
	LUT3 #(
		.INIT('h80)
	) name7090 (
		\wishbone_bd_ram_mem2_reg[239][19]/P0001 ,
		_w11973_,
		_w11982_,
		_w17603_
	);
	LUT4 #(
		.INIT('h0001)
	) name7091 (
		_w17600_,
		_w17601_,
		_w17602_,
		_w17603_,
		_w17604_
	);
	LUT4 #(
		.INIT('h8000)
	) name7092 (
		_w17589_,
		_w17594_,
		_w17599_,
		_w17604_,
		_w17605_
	);
	LUT3 #(
		.INIT('h80)
	) name7093 (
		\wishbone_bd_ram_mem2_reg[4][19]/P0001 ,
		_w11929_,
		_w11932_,
		_w17606_
	);
	LUT3 #(
		.INIT('h80)
	) name7094 (
		\wishbone_bd_ram_mem2_reg[2][19]/P0001 ,
		_w11932_,
		_w11963_,
		_w17607_
	);
	LUT3 #(
		.INIT('h80)
	) name7095 (
		\wishbone_bd_ram_mem2_reg[246][19]/P0001 ,
		_w11952_,
		_w11986_,
		_w17608_
	);
	LUT3 #(
		.INIT('h80)
	) name7096 (
		\wishbone_bd_ram_mem2_reg[133][19]/P0001 ,
		_w11933_,
		_w11955_,
		_w17609_
	);
	LUT4 #(
		.INIT('h0001)
	) name7097 (
		_w17606_,
		_w17607_,
		_w17608_,
		_w17609_,
		_w17610_
	);
	LUT3 #(
		.INIT('h80)
	) name7098 (
		\wishbone_bd_ram_mem2_reg[84][19]/P0001 ,
		_w11929_,
		_w11972_,
		_w17611_
	);
	LUT3 #(
		.INIT('h80)
	) name7099 (
		\wishbone_bd_ram_mem2_reg[24][19]/P0001 ,
		_w11935_,
		_w11990_,
		_w17612_
	);
	LUT3 #(
		.INIT('h80)
	) name7100 (
		\wishbone_bd_ram_mem2_reg[97][19]/P0001 ,
		_w11965_,
		_w11977_,
		_w17613_
	);
	LUT3 #(
		.INIT('h80)
	) name7101 (
		\wishbone_bd_ram_mem2_reg[1][19]/P0001 ,
		_w11932_,
		_w11977_,
		_w17614_
	);
	LUT4 #(
		.INIT('h0001)
	) name7102 (
		_w17611_,
		_w17612_,
		_w17613_,
		_w17614_,
		_w17615_
	);
	LUT3 #(
		.INIT('h80)
	) name7103 (
		\wishbone_bd_ram_mem2_reg[123][19]/P0001 ,
		_w11936_,
		_w12012_,
		_w17616_
	);
	LUT3 #(
		.INIT('h80)
	) name7104 (
		\wishbone_bd_ram_mem2_reg[88][19]/P0001 ,
		_w11972_,
		_w11990_,
		_w17617_
	);
	LUT3 #(
		.INIT('h80)
	) name7105 (
		\wishbone_bd_ram_mem2_reg[251][19]/P0001 ,
		_w11936_,
		_w11952_,
		_w17618_
	);
	LUT3 #(
		.INIT('h80)
	) name7106 (
		\wishbone_bd_ram_mem2_reg[81][19]/P0001 ,
		_w11972_,
		_w11977_,
		_w17619_
	);
	LUT4 #(
		.INIT('h0001)
	) name7107 (
		_w17616_,
		_w17617_,
		_w17618_,
		_w17619_,
		_w17620_
	);
	LUT3 #(
		.INIT('h80)
	) name7108 (
		\wishbone_bd_ram_mem2_reg[216][19]/P0001 ,
		_w11984_,
		_w11990_,
		_w17621_
	);
	LUT3 #(
		.INIT('h80)
	) name7109 (
		\wishbone_bd_ram_mem2_reg[177][19]/P0001 ,
		_w11942_,
		_w11977_,
		_w17622_
	);
	LUT3 #(
		.INIT('h80)
	) name7110 (
		\wishbone_bd_ram_mem2_reg[175][19]/P0001 ,
		_w11930_,
		_w11973_,
		_w17623_
	);
	LUT3 #(
		.INIT('h80)
	) name7111 (
		\wishbone_bd_ram_mem2_reg[243][19]/P0001 ,
		_w11938_,
		_w11952_,
		_w17624_
	);
	LUT4 #(
		.INIT('h0001)
	) name7112 (
		_w17621_,
		_w17622_,
		_w17623_,
		_w17624_,
		_w17625_
	);
	LUT4 #(
		.INIT('h8000)
	) name7113 (
		_w17610_,
		_w17615_,
		_w17620_,
		_w17625_,
		_w17626_
	);
	LUT4 #(
		.INIT('h8000)
	) name7114 (
		_w17563_,
		_w17584_,
		_w17605_,
		_w17626_,
		_w17627_
	);
	LUT3 #(
		.INIT('h80)
	) name7115 (
		\wishbone_bd_ram_mem2_reg[255][19]/P0001 ,
		_w11952_,
		_w11973_,
		_w17628_
	);
	LUT3 #(
		.INIT('h80)
	) name7116 (
		\wishbone_bd_ram_mem2_reg[155][19]/P0001 ,
		_w11936_,
		_w11959_,
		_w17629_
	);
	LUT3 #(
		.INIT('h80)
	) name7117 (
		\wishbone_bd_ram_mem2_reg[139][19]/P0001 ,
		_w11936_,
		_w11955_,
		_w17630_
	);
	LUT3 #(
		.INIT('h80)
	) name7118 (
		\wishbone_bd_ram_mem2_reg[250][19]/P0001 ,
		_w11944_,
		_w11952_,
		_w17631_
	);
	LUT4 #(
		.INIT('h0001)
	) name7119 (
		_w17628_,
		_w17629_,
		_w17630_,
		_w17631_,
		_w17632_
	);
	LUT3 #(
		.INIT('h80)
	) name7120 (
		\wishbone_bd_ram_mem2_reg[57][19]/P0001 ,
		_w11968_,
		_w11979_,
		_w17633_
	);
	LUT3 #(
		.INIT('h80)
	) name7121 (
		\wishbone_bd_ram_mem2_reg[232][19]/P0001 ,
		_w11982_,
		_w11990_,
		_w17634_
	);
	LUT3 #(
		.INIT('h80)
	) name7122 (
		\wishbone_bd_ram_mem2_reg[34][19]/P0001 ,
		_w11957_,
		_w11963_,
		_w17635_
	);
	LUT3 #(
		.INIT('h80)
	) name7123 (
		\wishbone_bd_ram_mem2_reg[82][19]/P0001 ,
		_w11963_,
		_w11972_,
		_w17636_
	);
	LUT4 #(
		.INIT('h0001)
	) name7124 (
		_w17633_,
		_w17634_,
		_w17635_,
		_w17636_,
		_w17637_
	);
	LUT3 #(
		.INIT('h80)
	) name7125 (
		\wishbone_bd_ram_mem2_reg[154][19]/P0001 ,
		_w11944_,
		_w11959_,
		_w17638_
	);
	LUT3 #(
		.INIT('h80)
	) name7126 (
		\wishbone_bd_ram_mem2_reg[76][19]/P0001 ,
		_w11949_,
		_w11954_,
		_w17639_
	);
	LUT3 #(
		.INIT('h80)
	) name7127 (
		\wishbone_bd_ram_mem2_reg[238][19]/P0001 ,
		_w11948_,
		_w11982_,
		_w17640_
	);
	LUT3 #(
		.INIT('h80)
	) name7128 (
		\wishbone_bd_ram_mem2_reg[8][19]/P0001 ,
		_w11932_,
		_w11990_,
		_w17641_
	);
	LUT4 #(
		.INIT('h0001)
	) name7129 (
		_w17638_,
		_w17639_,
		_w17640_,
		_w17641_,
		_w17642_
	);
	LUT3 #(
		.INIT('h80)
	) name7130 (
		\wishbone_bd_ram_mem2_reg[194][19]/P0001 ,
		_w11945_,
		_w11963_,
		_w17643_
	);
	LUT3 #(
		.INIT('h80)
	) name7131 (
		\wishbone_bd_ram_mem2_reg[44][19]/P0001 ,
		_w11954_,
		_w11957_,
		_w17644_
	);
	LUT3 #(
		.INIT('h80)
	) name7132 (
		\wishbone_bd_ram_mem2_reg[168][19]/P0001 ,
		_w11930_,
		_w11990_,
		_w17645_
	);
	LUT3 #(
		.INIT('h80)
	) name7133 (
		\wishbone_bd_ram_mem2_reg[209][19]/P0001 ,
		_w11977_,
		_w11984_,
		_w17646_
	);
	LUT4 #(
		.INIT('h0001)
	) name7134 (
		_w17643_,
		_w17644_,
		_w17645_,
		_w17646_,
		_w17647_
	);
	LUT4 #(
		.INIT('h8000)
	) name7135 (
		_w17632_,
		_w17637_,
		_w17642_,
		_w17647_,
		_w17648_
	);
	LUT3 #(
		.INIT('h80)
	) name7136 (
		\wishbone_bd_ram_mem2_reg[65][19]/P0001 ,
		_w11949_,
		_w11977_,
		_w17649_
	);
	LUT3 #(
		.INIT('h80)
	) name7137 (
		\wishbone_bd_ram_mem2_reg[234][19]/P0001 ,
		_w11944_,
		_w11982_,
		_w17650_
	);
	LUT3 #(
		.INIT('h80)
	) name7138 (
		\wishbone_bd_ram_mem2_reg[166][19]/P0001 ,
		_w11930_,
		_w11986_,
		_w17651_
	);
	LUT3 #(
		.INIT('h80)
	) name7139 (
		\wishbone_bd_ram_mem2_reg[78][19]/P0001 ,
		_w11948_,
		_w11949_,
		_w17652_
	);
	LUT4 #(
		.INIT('h0001)
	) name7140 (
		_w17649_,
		_w17650_,
		_w17651_,
		_w17652_,
		_w17653_
	);
	LUT3 #(
		.INIT('h80)
	) name7141 (
		\wishbone_bd_ram_mem2_reg[86][19]/P0001 ,
		_w11972_,
		_w11986_,
		_w17654_
	);
	LUT3 #(
		.INIT('h80)
	) name7142 (
		\wishbone_bd_ram_mem2_reg[137][19]/P0001 ,
		_w11955_,
		_w11968_,
		_w17655_
	);
	LUT3 #(
		.INIT('h80)
	) name7143 (
		\wishbone_bd_ram_mem2_reg[66][19]/P0001 ,
		_w11949_,
		_w11963_,
		_w17656_
	);
	LUT3 #(
		.INIT('h80)
	) name7144 (
		\wishbone_bd_ram_mem2_reg[221][19]/P0001 ,
		_w11966_,
		_w11984_,
		_w17657_
	);
	LUT4 #(
		.INIT('h0001)
	) name7145 (
		_w17654_,
		_w17655_,
		_w17656_,
		_w17657_,
		_w17658_
	);
	LUT3 #(
		.INIT('h80)
	) name7146 (
		\wishbone_bd_ram_mem2_reg[95][19]/P0001 ,
		_w11972_,
		_w11973_,
		_w17659_
	);
	LUT3 #(
		.INIT('h80)
	) name7147 (
		\wishbone_bd_ram_mem2_reg[99][19]/P0001 ,
		_w11938_,
		_w11965_,
		_w17660_
	);
	LUT3 #(
		.INIT('h80)
	) name7148 (
		\wishbone_bd_ram_mem2_reg[142][19]/P0001 ,
		_w11948_,
		_w11955_,
		_w17661_
	);
	LUT3 #(
		.INIT('h80)
	) name7149 (
		\wishbone_bd_ram_mem2_reg[153][19]/P0001 ,
		_w11959_,
		_w11968_,
		_w17662_
	);
	LUT4 #(
		.INIT('h0001)
	) name7150 (
		_w17659_,
		_w17660_,
		_w17661_,
		_w17662_,
		_w17663_
	);
	LUT3 #(
		.INIT('h80)
	) name7151 (
		\wishbone_bd_ram_mem2_reg[127][19]/P0001 ,
		_w11973_,
		_w12012_,
		_w17664_
	);
	LUT3 #(
		.INIT('h80)
	) name7152 (
		\wishbone_bd_ram_mem2_reg[244][19]/P0001 ,
		_w11929_,
		_w11952_,
		_w17665_
	);
	LUT3 #(
		.INIT('h80)
	) name7153 (
		\wishbone_bd_ram_mem2_reg[184][19]/P0001 ,
		_w11942_,
		_w11990_,
		_w17666_
	);
	LUT3 #(
		.INIT('h80)
	) name7154 (
		\wishbone_bd_ram_mem2_reg[117][19]/P0001 ,
		_w11933_,
		_w12012_,
		_w17667_
	);
	LUT4 #(
		.INIT('h0001)
	) name7155 (
		_w17664_,
		_w17665_,
		_w17666_,
		_w17667_,
		_w17668_
	);
	LUT4 #(
		.INIT('h8000)
	) name7156 (
		_w17653_,
		_w17658_,
		_w17663_,
		_w17668_,
		_w17669_
	);
	LUT3 #(
		.INIT('h80)
	) name7157 (
		\wishbone_bd_ram_mem2_reg[43][19]/P0001 ,
		_w11936_,
		_w11957_,
		_w17670_
	);
	LUT3 #(
		.INIT('h80)
	) name7158 (
		\wishbone_bd_ram_mem2_reg[231][19]/P0001 ,
		_w11975_,
		_w11982_,
		_w17671_
	);
	LUT3 #(
		.INIT('h80)
	) name7159 (
		\wishbone_bd_ram_mem2_reg[40][19]/P0001 ,
		_w11957_,
		_w11990_,
		_w17672_
	);
	LUT3 #(
		.INIT('h80)
	) name7160 (
		\wishbone_bd_ram_mem2_reg[93][19]/P0001 ,
		_w11966_,
		_w11972_,
		_w17673_
	);
	LUT4 #(
		.INIT('h0001)
	) name7161 (
		_w17670_,
		_w17671_,
		_w17672_,
		_w17673_,
		_w17674_
	);
	LUT3 #(
		.INIT('h80)
	) name7162 (
		\wishbone_bd_ram_mem2_reg[128][19]/P0001 ,
		_w11941_,
		_w11955_,
		_w17675_
	);
	LUT3 #(
		.INIT('h80)
	) name7163 (
		\wishbone_bd_ram_mem2_reg[254][19]/P0001 ,
		_w11948_,
		_w11952_,
		_w17676_
	);
	LUT3 #(
		.INIT('h80)
	) name7164 (
		\wishbone_bd_ram_mem2_reg[196][19]/P0001 ,
		_w11929_,
		_w11945_,
		_w17677_
	);
	LUT3 #(
		.INIT('h80)
	) name7165 (
		\wishbone_bd_ram_mem2_reg[17][19]/P0001 ,
		_w11935_,
		_w11977_,
		_w17678_
	);
	LUT4 #(
		.INIT('h0001)
	) name7166 (
		_w17675_,
		_w17676_,
		_w17677_,
		_w17678_,
		_w17679_
	);
	LUT3 #(
		.INIT('h80)
	) name7167 (
		\wishbone_bd_ram_mem2_reg[173][19]/P0001 ,
		_w11930_,
		_w11966_,
		_w17680_
	);
	LUT3 #(
		.INIT('h80)
	) name7168 (
		\wishbone_bd_ram_mem2_reg[240][19]/P0001 ,
		_w11941_,
		_w11952_,
		_w17681_
	);
	LUT3 #(
		.INIT('h80)
	) name7169 (
		\wishbone_bd_ram_mem2_reg[211][19]/P0001 ,
		_w11938_,
		_w11984_,
		_w17682_
	);
	LUT3 #(
		.INIT('h80)
	) name7170 (
		\wishbone_bd_ram_mem2_reg[116][19]/P0001 ,
		_w11929_,
		_w12012_,
		_w17683_
	);
	LUT4 #(
		.INIT('h0001)
	) name7171 (
		_w17680_,
		_w17681_,
		_w17682_,
		_w17683_,
		_w17684_
	);
	LUT3 #(
		.INIT('h80)
	) name7172 (
		\wishbone_bd_ram_mem2_reg[48][19]/P0001 ,
		_w11941_,
		_w11979_,
		_w17685_
	);
	LUT3 #(
		.INIT('h80)
	) name7173 (
		\wishbone_bd_ram_mem2_reg[141][19]/P0001 ,
		_w11955_,
		_w11966_,
		_w17686_
	);
	LUT3 #(
		.INIT('h80)
	) name7174 (
		\wishbone_bd_ram_mem2_reg[167][19]/P0001 ,
		_w11930_,
		_w11975_,
		_w17687_
	);
	LUT3 #(
		.INIT('h80)
	) name7175 (
		\wishbone_bd_ram_mem2_reg[125][19]/P0001 ,
		_w11966_,
		_w12012_,
		_w17688_
	);
	LUT4 #(
		.INIT('h0001)
	) name7176 (
		_w17685_,
		_w17686_,
		_w17687_,
		_w17688_,
		_w17689_
	);
	LUT4 #(
		.INIT('h8000)
	) name7177 (
		_w17674_,
		_w17679_,
		_w17684_,
		_w17689_,
		_w17690_
	);
	LUT3 #(
		.INIT('h80)
	) name7178 (
		\wishbone_bd_ram_mem2_reg[199][19]/P0001 ,
		_w11945_,
		_w11975_,
		_w17691_
	);
	LUT3 #(
		.INIT('h80)
	) name7179 (
		\wishbone_bd_ram_mem2_reg[71][19]/P0001 ,
		_w11949_,
		_w11975_,
		_w17692_
	);
	LUT3 #(
		.INIT('h80)
	) name7180 (
		\wishbone_bd_ram_mem2_reg[47][19]/P0001 ,
		_w11957_,
		_w11973_,
		_w17693_
	);
	LUT3 #(
		.INIT('h80)
	) name7181 (
		\wishbone_bd_ram_mem2_reg[29][19]/P0001 ,
		_w11935_,
		_w11966_,
		_w17694_
	);
	LUT4 #(
		.INIT('h0001)
	) name7182 (
		_w17691_,
		_w17692_,
		_w17693_,
		_w17694_,
		_w17695_
	);
	LUT3 #(
		.INIT('h80)
	) name7183 (
		\wishbone_bd_ram_mem2_reg[41][19]/P0001 ,
		_w11957_,
		_w11968_,
		_w17696_
	);
	LUT3 #(
		.INIT('h80)
	) name7184 (
		\wishbone_bd_ram_mem2_reg[33][19]/P0001 ,
		_w11957_,
		_w11977_,
		_w17697_
	);
	LUT3 #(
		.INIT('h80)
	) name7185 (
		\wishbone_bd_ram_mem2_reg[198][19]/P0001 ,
		_w11945_,
		_w11986_,
		_w17698_
	);
	LUT3 #(
		.INIT('h80)
	) name7186 (
		\wishbone_bd_ram_mem2_reg[0][19]/P0001 ,
		_w11932_,
		_w11941_,
		_w17699_
	);
	LUT4 #(
		.INIT('h0001)
	) name7187 (
		_w17696_,
		_w17697_,
		_w17698_,
		_w17699_,
		_w17700_
	);
	LUT3 #(
		.INIT('h80)
	) name7188 (
		\wishbone_bd_ram_mem2_reg[178][19]/P0001 ,
		_w11942_,
		_w11963_,
		_w17701_
	);
	LUT3 #(
		.INIT('h80)
	) name7189 (
		\wishbone_bd_ram_mem2_reg[75][19]/P0001 ,
		_w11936_,
		_w11949_,
		_w17702_
	);
	LUT3 #(
		.INIT('h80)
	) name7190 (
		\wishbone_bd_ram_mem2_reg[53][19]/P0001 ,
		_w11933_,
		_w11979_,
		_w17703_
	);
	LUT3 #(
		.INIT('h80)
	) name7191 (
		\wishbone_bd_ram_mem2_reg[111][19]/P0001 ,
		_w11965_,
		_w11973_,
		_w17704_
	);
	LUT4 #(
		.INIT('h0001)
	) name7192 (
		_w17701_,
		_w17702_,
		_w17703_,
		_w17704_,
		_w17705_
	);
	LUT3 #(
		.INIT('h80)
	) name7193 (
		\wishbone_bd_ram_mem2_reg[110][19]/P0001 ,
		_w11948_,
		_w11965_,
		_w17706_
	);
	LUT3 #(
		.INIT('h80)
	) name7194 (
		\wishbone_bd_ram_mem2_reg[59][19]/P0001 ,
		_w11936_,
		_w11979_,
		_w17707_
	);
	LUT3 #(
		.INIT('h80)
	) name7195 (
		\wishbone_bd_ram_mem2_reg[140][19]/P0001 ,
		_w11954_,
		_w11955_,
		_w17708_
	);
	LUT3 #(
		.INIT('h80)
	) name7196 (
		\wishbone_bd_ram_mem2_reg[9][19]/P0001 ,
		_w11932_,
		_w11968_,
		_w17709_
	);
	LUT4 #(
		.INIT('h0001)
	) name7197 (
		_w17706_,
		_w17707_,
		_w17708_,
		_w17709_,
		_w17710_
	);
	LUT4 #(
		.INIT('h8000)
	) name7198 (
		_w17695_,
		_w17700_,
		_w17705_,
		_w17710_,
		_w17711_
	);
	LUT4 #(
		.INIT('h8000)
	) name7199 (
		_w17648_,
		_w17669_,
		_w17690_,
		_w17711_,
		_w17712_
	);
	LUT4 #(
		.INIT('h8000)
	) name7200 (
		_w17457_,
		_w17542_,
		_w17627_,
		_w17712_,
		_w17713_
	);
	LUT3 #(
		.INIT('hce)
	) name7201 (
		_w12303_,
		_w17372_,
		_w17713_,
		_w17714_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name7202 (
		\wishbone_LatchedTxLength_reg[4]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w17715_
	);
	LUT3 #(
		.INIT('hf2)
	) name7203 (
		_w12303_,
		_w14512_,
		_w17715_,
		_w17716_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name7204 (
		\wishbone_LatchedTxLength_reg[5]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w17717_
	);
	LUT3 #(
		.INIT('h80)
	) name7205 (
		\wishbone_bd_ram_mem2_reg[68][21]/P0001 ,
		_w11929_,
		_w11949_,
		_w17718_
	);
	LUT3 #(
		.INIT('h80)
	) name7206 (
		\wishbone_bd_ram_mem2_reg[175][21]/P0001 ,
		_w11930_,
		_w11973_,
		_w17719_
	);
	LUT3 #(
		.INIT('h80)
	) name7207 (
		\wishbone_bd_ram_mem2_reg[37][21]/P0001 ,
		_w11933_,
		_w11957_,
		_w17720_
	);
	LUT3 #(
		.INIT('h80)
	) name7208 (
		\wishbone_bd_ram_mem2_reg[169][21]/P0001 ,
		_w11930_,
		_w11968_,
		_w17721_
	);
	LUT4 #(
		.INIT('h0001)
	) name7209 (
		_w17718_,
		_w17719_,
		_w17720_,
		_w17721_,
		_w17722_
	);
	LUT3 #(
		.INIT('h80)
	) name7210 (
		\wishbone_bd_ram_mem2_reg[101][21]/P0001 ,
		_w11933_,
		_w11965_,
		_w17723_
	);
	LUT3 #(
		.INIT('h80)
	) name7211 (
		\wishbone_bd_ram_mem2_reg[99][21]/P0001 ,
		_w11938_,
		_w11965_,
		_w17724_
	);
	LUT3 #(
		.INIT('h80)
	) name7212 (
		\wishbone_bd_ram_mem2_reg[119][21]/P0001 ,
		_w11975_,
		_w12012_,
		_w17725_
	);
	LUT3 #(
		.INIT('h80)
	) name7213 (
		\wishbone_bd_ram_mem2_reg[145][21]/P0001 ,
		_w11959_,
		_w11977_,
		_w17726_
	);
	LUT4 #(
		.INIT('h0001)
	) name7214 (
		_w17723_,
		_w17724_,
		_w17725_,
		_w17726_,
		_w17727_
	);
	LUT3 #(
		.INIT('h80)
	) name7215 (
		\wishbone_bd_ram_mem2_reg[254][21]/P0001 ,
		_w11948_,
		_w11952_,
		_w17728_
	);
	LUT3 #(
		.INIT('h80)
	) name7216 (
		\wishbone_bd_ram_mem2_reg[183][21]/P0001 ,
		_w11942_,
		_w11975_,
		_w17729_
	);
	LUT3 #(
		.INIT('h80)
	) name7217 (
		\wishbone_bd_ram_mem2_reg[38][21]/P0001 ,
		_w11957_,
		_w11986_,
		_w17730_
	);
	LUT3 #(
		.INIT('h80)
	) name7218 (
		\wishbone_bd_ram_mem2_reg[232][21]/P0001 ,
		_w11982_,
		_w11990_,
		_w17731_
	);
	LUT4 #(
		.INIT('h0001)
	) name7219 (
		_w17728_,
		_w17729_,
		_w17730_,
		_w17731_,
		_w17732_
	);
	LUT3 #(
		.INIT('h80)
	) name7220 (
		\wishbone_bd_ram_mem2_reg[109][21]/P0001 ,
		_w11965_,
		_w11966_,
		_w17733_
	);
	LUT3 #(
		.INIT('h80)
	) name7221 (
		\wishbone_bd_ram_mem2_reg[122][21]/P0001 ,
		_w11944_,
		_w12012_,
		_w17734_
	);
	LUT3 #(
		.INIT('h80)
	) name7222 (
		\wishbone_bd_ram_mem2_reg[28][21]/P0001 ,
		_w11935_,
		_w11954_,
		_w17735_
	);
	LUT3 #(
		.INIT('h80)
	) name7223 (
		\wishbone_bd_ram_mem2_reg[156][21]/P0001 ,
		_w11954_,
		_w11959_,
		_w17736_
	);
	LUT4 #(
		.INIT('h0001)
	) name7224 (
		_w17733_,
		_w17734_,
		_w17735_,
		_w17736_,
		_w17737_
	);
	LUT4 #(
		.INIT('h8000)
	) name7225 (
		_w17722_,
		_w17727_,
		_w17732_,
		_w17737_,
		_w17738_
	);
	LUT3 #(
		.INIT('h80)
	) name7226 (
		\wishbone_bd_ram_mem2_reg[64][21]/P0001 ,
		_w11941_,
		_w11949_,
		_w17739_
	);
	LUT3 #(
		.INIT('h80)
	) name7227 (
		\wishbone_bd_ram_mem2_reg[157][21]/P0001 ,
		_w11959_,
		_w11966_,
		_w17740_
	);
	LUT3 #(
		.INIT('h80)
	) name7228 (
		\wishbone_bd_ram_mem2_reg[144][21]/P0001 ,
		_w11941_,
		_w11959_,
		_w17741_
	);
	LUT3 #(
		.INIT('h80)
	) name7229 (
		\wishbone_bd_ram_mem2_reg[155][21]/P0001 ,
		_w11936_,
		_w11959_,
		_w17742_
	);
	LUT4 #(
		.INIT('h0001)
	) name7230 (
		_w17739_,
		_w17740_,
		_w17741_,
		_w17742_,
		_w17743_
	);
	LUT3 #(
		.INIT('h80)
	) name7231 (
		\wishbone_bd_ram_mem2_reg[23][21]/P0001 ,
		_w11935_,
		_w11975_,
		_w17744_
	);
	LUT3 #(
		.INIT('h80)
	) name7232 (
		\wishbone_bd_ram_mem2_reg[143][21]/P0001 ,
		_w11955_,
		_w11973_,
		_w17745_
	);
	LUT3 #(
		.INIT('h80)
	) name7233 (
		\wishbone_bd_ram_mem2_reg[48][21]/P0001 ,
		_w11941_,
		_w11979_,
		_w17746_
	);
	LUT3 #(
		.INIT('h80)
	) name7234 (
		\wishbone_bd_ram_mem2_reg[9][21]/P0001 ,
		_w11932_,
		_w11968_,
		_w17747_
	);
	LUT4 #(
		.INIT('h0001)
	) name7235 (
		_w17744_,
		_w17745_,
		_w17746_,
		_w17747_,
		_w17748_
	);
	LUT3 #(
		.INIT('h80)
	) name7236 (
		\wishbone_bd_ram_mem2_reg[58][21]/P0001 ,
		_w11944_,
		_w11979_,
		_w17749_
	);
	LUT3 #(
		.INIT('h80)
	) name7237 (
		\wishbone_bd_ram_mem2_reg[198][21]/P0001 ,
		_w11945_,
		_w11986_,
		_w17750_
	);
	LUT3 #(
		.INIT('h80)
	) name7238 (
		\wishbone_bd_ram_mem2_reg[246][21]/P0001 ,
		_w11952_,
		_w11986_,
		_w17751_
	);
	LUT3 #(
		.INIT('h80)
	) name7239 (
		\wishbone_bd_ram_mem2_reg[95][21]/P0001 ,
		_w11972_,
		_w11973_,
		_w17752_
	);
	LUT4 #(
		.INIT('h0001)
	) name7240 (
		_w17749_,
		_w17750_,
		_w17751_,
		_w17752_,
		_w17753_
	);
	LUT3 #(
		.INIT('h80)
	) name7241 (
		\wishbone_bd_ram_mem2_reg[24][21]/P0001 ,
		_w11935_,
		_w11990_,
		_w17754_
	);
	LUT3 #(
		.INIT('h80)
	) name7242 (
		\wishbone_bd_ram_mem2_reg[209][21]/P0001 ,
		_w11977_,
		_w11984_,
		_w17755_
	);
	LUT3 #(
		.INIT('h80)
	) name7243 (
		\wishbone_bd_ram_mem2_reg[149][21]/P0001 ,
		_w11933_,
		_w11959_,
		_w17756_
	);
	LUT3 #(
		.INIT('h80)
	) name7244 (
		\wishbone_bd_ram_mem2_reg[207][21]/P0001 ,
		_w11945_,
		_w11973_,
		_w17757_
	);
	LUT4 #(
		.INIT('h0001)
	) name7245 (
		_w17754_,
		_w17755_,
		_w17756_,
		_w17757_,
		_w17758_
	);
	LUT4 #(
		.INIT('h8000)
	) name7246 (
		_w17743_,
		_w17748_,
		_w17753_,
		_w17758_,
		_w17759_
	);
	LUT3 #(
		.INIT('h80)
	) name7247 (
		\wishbone_bd_ram_mem2_reg[114][21]/P0001 ,
		_w11963_,
		_w12012_,
		_w17760_
	);
	LUT3 #(
		.INIT('h80)
	) name7248 (
		\wishbone_bd_ram_mem2_reg[129][21]/P0001 ,
		_w11955_,
		_w11977_,
		_w17761_
	);
	LUT3 #(
		.INIT('h80)
	) name7249 (
		\wishbone_bd_ram_mem2_reg[70][21]/P0001 ,
		_w11949_,
		_w11986_,
		_w17762_
	);
	LUT3 #(
		.INIT('h80)
	) name7250 (
		\wishbone_bd_ram_mem2_reg[166][21]/P0001 ,
		_w11930_,
		_w11986_,
		_w17763_
	);
	LUT4 #(
		.INIT('h0001)
	) name7251 (
		_w17760_,
		_w17761_,
		_w17762_,
		_w17763_,
		_w17764_
	);
	LUT3 #(
		.INIT('h80)
	) name7252 (
		\wishbone_bd_ram_mem2_reg[65][21]/P0001 ,
		_w11949_,
		_w11977_,
		_w17765_
	);
	LUT3 #(
		.INIT('h80)
	) name7253 (
		\wishbone_bd_ram_mem2_reg[77][21]/P0001 ,
		_w11949_,
		_w11966_,
		_w17766_
	);
	LUT3 #(
		.INIT('h80)
	) name7254 (
		\wishbone_bd_ram_mem2_reg[195][21]/P0001 ,
		_w11938_,
		_w11945_,
		_w17767_
	);
	LUT3 #(
		.INIT('h80)
	) name7255 (
		\wishbone_bd_ram_mem2_reg[192][21]/P0001 ,
		_w11941_,
		_w11945_,
		_w17768_
	);
	LUT4 #(
		.INIT('h0001)
	) name7256 (
		_w17765_,
		_w17766_,
		_w17767_,
		_w17768_,
		_w17769_
	);
	LUT3 #(
		.INIT('h80)
	) name7257 (
		\wishbone_bd_ram_mem2_reg[80][21]/P0001 ,
		_w11941_,
		_w11972_,
		_w17770_
	);
	LUT3 #(
		.INIT('h80)
	) name7258 (
		\wishbone_bd_ram_mem2_reg[210][21]/P0001 ,
		_w11963_,
		_w11984_,
		_w17771_
	);
	LUT3 #(
		.INIT('h80)
	) name7259 (
		\wishbone_bd_ram_mem2_reg[208][21]/P0001 ,
		_w11941_,
		_w11984_,
		_w17772_
	);
	LUT3 #(
		.INIT('h80)
	) name7260 (
		\wishbone_bd_ram_mem2_reg[184][21]/P0001 ,
		_w11942_,
		_w11990_,
		_w17773_
	);
	LUT4 #(
		.INIT('h0001)
	) name7261 (
		_w17770_,
		_w17771_,
		_w17772_,
		_w17773_,
		_w17774_
	);
	LUT3 #(
		.INIT('h80)
	) name7262 (
		\wishbone_bd_ram_mem2_reg[14][21]/P0001 ,
		_w11932_,
		_w11948_,
		_w17775_
	);
	LUT3 #(
		.INIT('h80)
	) name7263 (
		\wishbone_bd_ram_mem2_reg[222][21]/P0001 ,
		_w11948_,
		_w11984_,
		_w17776_
	);
	LUT3 #(
		.INIT('h80)
	) name7264 (
		\wishbone_bd_ram_mem2_reg[40][21]/P0001 ,
		_w11957_,
		_w11990_,
		_w17777_
	);
	LUT3 #(
		.INIT('h80)
	) name7265 (
		\wishbone_bd_ram_mem2_reg[181][21]/P0001 ,
		_w11933_,
		_w11942_,
		_w17778_
	);
	LUT4 #(
		.INIT('h0001)
	) name7266 (
		_w17775_,
		_w17776_,
		_w17777_,
		_w17778_,
		_w17779_
	);
	LUT4 #(
		.INIT('h8000)
	) name7267 (
		_w17764_,
		_w17769_,
		_w17774_,
		_w17779_,
		_w17780_
	);
	LUT3 #(
		.INIT('h80)
	) name7268 (
		\wishbone_bd_ram_mem2_reg[63][21]/P0001 ,
		_w11973_,
		_w11979_,
		_w17781_
	);
	LUT3 #(
		.INIT('h80)
	) name7269 (
		\wishbone_bd_ram_mem2_reg[125][21]/P0001 ,
		_w11966_,
		_w12012_,
		_w17782_
	);
	LUT3 #(
		.INIT('h80)
	) name7270 (
		\wishbone_bd_ram_mem2_reg[104][21]/P0001 ,
		_w11965_,
		_w11990_,
		_w17783_
	);
	LUT3 #(
		.INIT('h80)
	) name7271 (
		\wishbone_bd_ram_mem2_reg[85][21]/P0001 ,
		_w11933_,
		_w11972_,
		_w17784_
	);
	LUT4 #(
		.INIT('h0001)
	) name7272 (
		_w17781_,
		_w17782_,
		_w17783_,
		_w17784_,
		_w17785_
	);
	LUT3 #(
		.INIT('h80)
	) name7273 (
		\wishbone_bd_ram_mem2_reg[81][21]/P0001 ,
		_w11972_,
		_w11977_,
		_w17786_
	);
	LUT3 #(
		.INIT('h80)
	) name7274 (
		\wishbone_bd_ram_mem2_reg[78][21]/P0001 ,
		_w11948_,
		_w11949_,
		_w17787_
	);
	LUT3 #(
		.INIT('h80)
	) name7275 (
		\wishbone_bd_ram_mem2_reg[50][21]/P0001 ,
		_w11963_,
		_w11979_,
		_w17788_
	);
	LUT3 #(
		.INIT('h80)
	) name7276 (
		\wishbone_bd_ram_mem2_reg[127][21]/P0001 ,
		_w11973_,
		_w12012_,
		_w17789_
	);
	LUT4 #(
		.INIT('h0001)
	) name7277 (
		_w17786_,
		_w17787_,
		_w17788_,
		_w17789_,
		_w17790_
	);
	LUT3 #(
		.INIT('h80)
	) name7278 (
		\wishbone_bd_ram_mem2_reg[196][21]/P0001 ,
		_w11929_,
		_w11945_,
		_w17791_
	);
	LUT3 #(
		.INIT('h80)
	) name7279 (
		\wishbone_bd_ram_mem2_reg[27][21]/P0001 ,
		_w11935_,
		_w11936_,
		_w17792_
	);
	LUT3 #(
		.INIT('h80)
	) name7280 (
		\wishbone_bd_ram_mem2_reg[22][21]/P0001 ,
		_w11935_,
		_w11986_,
		_w17793_
	);
	LUT3 #(
		.INIT('h80)
	) name7281 (
		\wishbone_bd_ram_mem2_reg[1][21]/P0001 ,
		_w11932_,
		_w11977_,
		_w17794_
	);
	LUT4 #(
		.INIT('h0001)
	) name7282 (
		_w17791_,
		_w17792_,
		_w17793_,
		_w17794_,
		_w17795_
	);
	LUT3 #(
		.INIT('h80)
	) name7283 (
		\wishbone_bd_ram_mem2_reg[162][21]/P0001 ,
		_w11930_,
		_w11963_,
		_w17796_
	);
	LUT3 #(
		.INIT('h80)
	) name7284 (
		\wishbone_bd_ram_mem2_reg[7][21]/P0001 ,
		_w11932_,
		_w11975_,
		_w17797_
	);
	LUT3 #(
		.INIT('h80)
	) name7285 (
		\wishbone_bd_ram_mem2_reg[151][21]/P0001 ,
		_w11959_,
		_w11975_,
		_w17798_
	);
	LUT3 #(
		.INIT('h80)
	) name7286 (
		\wishbone_bd_ram_mem2_reg[62][21]/P0001 ,
		_w11948_,
		_w11979_,
		_w17799_
	);
	LUT4 #(
		.INIT('h0001)
	) name7287 (
		_w17796_,
		_w17797_,
		_w17798_,
		_w17799_,
		_w17800_
	);
	LUT4 #(
		.INIT('h8000)
	) name7288 (
		_w17785_,
		_w17790_,
		_w17795_,
		_w17800_,
		_w17801_
	);
	LUT4 #(
		.INIT('h8000)
	) name7289 (
		_w17738_,
		_w17759_,
		_w17780_,
		_w17801_,
		_w17802_
	);
	LUT3 #(
		.INIT('h80)
	) name7290 (
		\wishbone_bd_ram_mem2_reg[148][21]/P0001 ,
		_w11929_,
		_w11959_,
		_w17803_
	);
	LUT3 #(
		.INIT('h80)
	) name7291 (
		\wishbone_bd_ram_mem2_reg[193][21]/P0001 ,
		_w11945_,
		_w11977_,
		_w17804_
	);
	LUT3 #(
		.INIT('h80)
	) name7292 (
		\wishbone_bd_ram_mem2_reg[220][21]/P0001 ,
		_w11954_,
		_w11984_,
		_w17805_
	);
	LUT3 #(
		.INIT('h80)
	) name7293 (
		\wishbone_bd_ram_mem2_reg[230][21]/P0001 ,
		_w11982_,
		_w11986_,
		_w17806_
	);
	LUT4 #(
		.INIT('h0001)
	) name7294 (
		_w17803_,
		_w17804_,
		_w17805_,
		_w17806_,
		_w17807_
	);
	LUT3 #(
		.INIT('h80)
	) name7295 (
		\wishbone_bd_ram_mem2_reg[242][21]/P0001 ,
		_w11952_,
		_w11963_,
		_w17808_
	);
	LUT3 #(
		.INIT('h80)
	) name7296 (
		\wishbone_bd_ram_mem2_reg[111][21]/P0001 ,
		_w11965_,
		_w11973_,
		_w17809_
	);
	LUT3 #(
		.INIT('h80)
	) name7297 (
		\wishbone_bd_ram_mem2_reg[2][21]/P0001 ,
		_w11932_,
		_w11963_,
		_w17810_
	);
	LUT3 #(
		.INIT('h80)
	) name7298 (
		\wishbone_bd_ram_mem2_reg[179][21]/P0001 ,
		_w11938_,
		_w11942_,
		_w17811_
	);
	LUT4 #(
		.INIT('h0001)
	) name7299 (
		_w17808_,
		_w17809_,
		_w17810_,
		_w17811_,
		_w17812_
	);
	LUT3 #(
		.INIT('h80)
	) name7300 (
		\wishbone_bd_ram_mem2_reg[168][21]/P0001 ,
		_w11930_,
		_w11990_,
		_w17813_
	);
	LUT3 #(
		.INIT('h80)
	) name7301 (
		\wishbone_bd_ram_mem2_reg[115][21]/P0001 ,
		_w11938_,
		_w12012_,
		_w17814_
	);
	LUT3 #(
		.INIT('h80)
	) name7302 (
		\wishbone_bd_ram_mem2_reg[82][21]/P0001 ,
		_w11963_,
		_w11972_,
		_w17815_
	);
	LUT3 #(
		.INIT('h80)
	) name7303 (
		\wishbone_bd_ram_mem2_reg[177][21]/P0001 ,
		_w11942_,
		_w11977_,
		_w17816_
	);
	LUT4 #(
		.INIT('h0001)
	) name7304 (
		_w17813_,
		_w17814_,
		_w17815_,
		_w17816_,
		_w17817_
	);
	LUT3 #(
		.INIT('h80)
	) name7305 (
		\wishbone_bd_ram_mem2_reg[87][21]/P0001 ,
		_w11972_,
		_w11975_,
		_w17818_
	);
	LUT3 #(
		.INIT('h80)
	) name7306 (
		\wishbone_bd_ram_mem2_reg[141][21]/P0001 ,
		_w11955_,
		_w11966_,
		_w17819_
	);
	LUT3 #(
		.INIT('h80)
	) name7307 (
		\wishbone_bd_ram_mem2_reg[8][21]/P0001 ,
		_w11932_,
		_w11990_,
		_w17820_
	);
	LUT3 #(
		.INIT('h80)
	) name7308 (
		\wishbone_bd_ram_mem2_reg[186][21]/P0001 ,
		_w11942_,
		_w11944_,
		_w17821_
	);
	LUT4 #(
		.INIT('h0001)
	) name7309 (
		_w17818_,
		_w17819_,
		_w17820_,
		_w17821_,
		_w17822_
	);
	LUT4 #(
		.INIT('h8000)
	) name7310 (
		_w17807_,
		_w17812_,
		_w17817_,
		_w17822_,
		_w17823_
	);
	LUT3 #(
		.INIT('h80)
	) name7311 (
		\wishbone_bd_ram_mem2_reg[128][21]/P0001 ,
		_w11941_,
		_w11955_,
		_w17824_
	);
	LUT3 #(
		.INIT('h80)
	) name7312 (
		\wishbone_bd_ram_mem2_reg[255][21]/P0001 ,
		_w11952_,
		_w11973_,
		_w17825_
	);
	LUT3 #(
		.INIT('h80)
	) name7313 (
		\wishbone_bd_ram_mem2_reg[90][21]/P0001 ,
		_w11944_,
		_w11972_,
		_w17826_
	);
	LUT3 #(
		.INIT('h80)
	) name7314 (
		\wishbone_bd_ram_mem2_reg[178][21]/P0001 ,
		_w11942_,
		_w11963_,
		_w17827_
	);
	LUT4 #(
		.INIT('h0001)
	) name7315 (
		_w17824_,
		_w17825_,
		_w17826_,
		_w17827_,
		_w17828_
	);
	LUT3 #(
		.INIT('h80)
	) name7316 (
		\wishbone_bd_ram_mem2_reg[44][21]/P0001 ,
		_w11954_,
		_w11957_,
		_w17829_
	);
	LUT3 #(
		.INIT('h80)
	) name7317 (
		\wishbone_bd_ram_mem2_reg[30][21]/P0001 ,
		_w11935_,
		_w11948_,
		_w17830_
	);
	LUT3 #(
		.INIT('h80)
	) name7318 (
		\wishbone_bd_ram_mem2_reg[171][21]/P0001 ,
		_w11930_,
		_w11936_,
		_w17831_
	);
	LUT3 #(
		.INIT('h80)
	) name7319 (
		\wishbone_bd_ram_mem2_reg[17][21]/P0001 ,
		_w11935_,
		_w11977_,
		_w17832_
	);
	LUT4 #(
		.INIT('h0001)
	) name7320 (
		_w17829_,
		_w17830_,
		_w17831_,
		_w17832_,
		_w17833_
	);
	LUT3 #(
		.INIT('h80)
	) name7321 (
		\wishbone_bd_ram_mem2_reg[212][21]/P0001 ,
		_w11929_,
		_w11984_,
		_w17834_
	);
	LUT3 #(
		.INIT('h80)
	) name7322 (
		\wishbone_bd_ram_mem2_reg[165][21]/P0001 ,
		_w11930_,
		_w11933_,
		_w17835_
	);
	LUT3 #(
		.INIT('h80)
	) name7323 (
		\wishbone_bd_ram_mem2_reg[102][21]/P0001 ,
		_w11965_,
		_w11986_,
		_w17836_
	);
	LUT3 #(
		.INIT('h80)
	) name7324 (
		\wishbone_bd_ram_mem2_reg[213][21]/P0001 ,
		_w11933_,
		_w11984_,
		_w17837_
	);
	LUT4 #(
		.INIT('h0001)
	) name7325 (
		_w17834_,
		_w17835_,
		_w17836_,
		_w17837_,
		_w17838_
	);
	LUT3 #(
		.INIT('h80)
	) name7326 (
		\wishbone_bd_ram_mem2_reg[60][21]/P0001 ,
		_w11954_,
		_w11979_,
		_w17839_
	);
	LUT3 #(
		.INIT('h80)
	) name7327 (
		\wishbone_bd_ram_mem2_reg[238][21]/P0001 ,
		_w11948_,
		_w11982_,
		_w17840_
	);
	LUT3 #(
		.INIT('h80)
	) name7328 (
		\wishbone_bd_ram_mem2_reg[173][21]/P0001 ,
		_w11930_,
		_w11966_,
		_w17841_
	);
	LUT3 #(
		.INIT('h80)
	) name7329 (
		\wishbone_bd_ram_mem2_reg[94][21]/P0001 ,
		_w11948_,
		_w11972_,
		_w17842_
	);
	LUT4 #(
		.INIT('h0001)
	) name7330 (
		_w17839_,
		_w17840_,
		_w17841_,
		_w17842_,
		_w17843_
	);
	LUT4 #(
		.INIT('h8000)
	) name7331 (
		_w17828_,
		_w17833_,
		_w17838_,
		_w17843_,
		_w17844_
	);
	LUT3 #(
		.INIT('h80)
	) name7332 (
		\wishbone_bd_ram_mem2_reg[117][21]/P0001 ,
		_w11933_,
		_w12012_,
		_w17845_
	);
	LUT3 #(
		.INIT('h80)
	) name7333 (
		\wishbone_bd_ram_mem2_reg[100][21]/P0001 ,
		_w11929_,
		_w11965_,
		_w17846_
	);
	LUT3 #(
		.INIT('h80)
	) name7334 (
		\wishbone_bd_ram_mem2_reg[182][21]/P0001 ,
		_w11942_,
		_w11986_,
		_w17847_
	);
	LUT3 #(
		.INIT('h80)
	) name7335 (
		\wishbone_bd_ram_mem2_reg[247][21]/P0001 ,
		_w11952_,
		_w11975_,
		_w17848_
	);
	LUT4 #(
		.INIT('h0001)
	) name7336 (
		_w17845_,
		_w17846_,
		_w17847_,
		_w17848_,
		_w17849_
	);
	LUT3 #(
		.INIT('h80)
	) name7337 (
		\wishbone_bd_ram_mem2_reg[191][21]/P0001 ,
		_w11942_,
		_w11973_,
		_w17850_
	);
	LUT3 #(
		.INIT('h80)
	) name7338 (
		\wishbone_bd_ram_mem2_reg[214][21]/P0001 ,
		_w11984_,
		_w11986_,
		_w17851_
	);
	LUT3 #(
		.INIT('h80)
	) name7339 (
		\wishbone_bd_ram_mem2_reg[120][21]/P0001 ,
		_w11990_,
		_w12012_,
		_w17852_
	);
	LUT3 #(
		.INIT('h80)
	) name7340 (
		\wishbone_bd_ram_mem2_reg[5][21]/P0001 ,
		_w11932_,
		_w11933_,
		_w17853_
	);
	LUT4 #(
		.INIT('h0001)
	) name7341 (
		_w17850_,
		_w17851_,
		_w17852_,
		_w17853_,
		_w17854_
	);
	LUT3 #(
		.INIT('h80)
	) name7342 (
		\wishbone_bd_ram_mem2_reg[237][21]/P0001 ,
		_w11966_,
		_w11982_,
		_w17855_
	);
	LUT3 #(
		.INIT('h80)
	) name7343 (
		\wishbone_bd_ram_mem2_reg[21][21]/P0001 ,
		_w11933_,
		_w11935_,
		_w17856_
	);
	LUT3 #(
		.INIT('h80)
	) name7344 (
		\wishbone_bd_ram_mem2_reg[134][21]/P0001 ,
		_w11955_,
		_w11986_,
		_w17857_
	);
	LUT3 #(
		.INIT('h80)
	) name7345 (
		\wishbone_bd_ram_mem2_reg[211][21]/P0001 ,
		_w11938_,
		_w11984_,
		_w17858_
	);
	LUT4 #(
		.INIT('h0001)
	) name7346 (
		_w17855_,
		_w17856_,
		_w17857_,
		_w17858_,
		_w17859_
	);
	LUT3 #(
		.INIT('h80)
	) name7347 (
		\wishbone_bd_ram_mem2_reg[108][21]/P0001 ,
		_w11954_,
		_w11965_,
		_w17860_
	);
	LUT3 #(
		.INIT('h80)
	) name7348 (
		\wishbone_bd_ram_mem2_reg[190][21]/P0001 ,
		_w11942_,
		_w11948_,
		_w17861_
	);
	LUT3 #(
		.INIT('h80)
	) name7349 (
		\wishbone_bd_ram_mem2_reg[45][21]/P0001 ,
		_w11957_,
		_w11966_,
		_w17862_
	);
	LUT3 #(
		.INIT('h80)
	) name7350 (
		\wishbone_bd_ram_mem2_reg[15][21]/P0001 ,
		_w11932_,
		_w11973_,
		_w17863_
	);
	LUT4 #(
		.INIT('h0001)
	) name7351 (
		_w17860_,
		_w17861_,
		_w17862_,
		_w17863_,
		_w17864_
	);
	LUT4 #(
		.INIT('h8000)
	) name7352 (
		_w17849_,
		_w17854_,
		_w17859_,
		_w17864_,
		_w17865_
	);
	LUT3 #(
		.INIT('h80)
	) name7353 (
		\wishbone_bd_ram_mem2_reg[203][21]/P0001 ,
		_w11936_,
		_w11945_,
		_w17866_
	);
	LUT3 #(
		.INIT('h80)
	) name7354 (
		\wishbone_bd_ram_mem2_reg[229][21]/P0001 ,
		_w11933_,
		_w11982_,
		_w17867_
	);
	LUT3 #(
		.INIT('h80)
	) name7355 (
		\wishbone_bd_ram_mem2_reg[116][21]/P0001 ,
		_w11929_,
		_w12012_,
		_w17868_
	);
	LUT3 #(
		.INIT('h80)
	) name7356 (
		\wishbone_bd_ram_mem2_reg[234][21]/P0001 ,
		_w11944_,
		_w11982_,
		_w17869_
	);
	LUT4 #(
		.INIT('h0001)
	) name7357 (
		_w17866_,
		_w17867_,
		_w17868_,
		_w17869_,
		_w17870_
	);
	LUT3 #(
		.INIT('h80)
	) name7358 (
		\wishbone_bd_ram_mem2_reg[51][21]/P0001 ,
		_w11938_,
		_w11979_,
		_w17871_
	);
	LUT3 #(
		.INIT('h80)
	) name7359 (
		\wishbone_bd_ram_mem2_reg[93][21]/P0001 ,
		_w11966_,
		_w11972_,
		_w17872_
	);
	LUT3 #(
		.INIT('h80)
	) name7360 (
		\wishbone_bd_ram_mem2_reg[226][21]/P0001 ,
		_w11963_,
		_w11982_,
		_w17873_
	);
	LUT3 #(
		.INIT('h80)
	) name7361 (
		\wishbone_bd_ram_mem2_reg[176][21]/P0001 ,
		_w11941_,
		_w11942_,
		_w17874_
	);
	LUT4 #(
		.INIT('h0001)
	) name7362 (
		_w17871_,
		_w17872_,
		_w17873_,
		_w17874_,
		_w17875_
	);
	LUT3 #(
		.INIT('h80)
	) name7363 (
		\wishbone_bd_ram_mem2_reg[121][21]/P0001 ,
		_w11968_,
		_w12012_,
		_w17876_
	);
	LUT3 #(
		.INIT('h80)
	) name7364 (
		\wishbone_bd_ram_mem2_reg[10][21]/P0001 ,
		_w11932_,
		_w11944_,
		_w17877_
	);
	LUT3 #(
		.INIT('h80)
	) name7365 (
		\wishbone_bd_ram_mem2_reg[147][21]/P0001 ,
		_w11938_,
		_w11959_,
		_w17878_
	);
	LUT3 #(
		.INIT('h80)
	) name7366 (
		\wishbone_bd_ram_mem2_reg[206][21]/P0001 ,
		_w11945_,
		_w11948_,
		_w17879_
	);
	LUT4 #(
		.INIT('h0001)
	) name7367 (
		_w17876_,
		_w17877_,
		_w17878_,
		_w17879_,
		_w17880_
	);
	LUT3 #(
		.INIT('h80)
	) name7368 (
		\wishbone_bd_ram_mem2_reg[243][21]/P0001 ,
		_w11938_,
		_w11952_,
		_w17881_
	);
	LUT3 #(
		.INIT('h80)
	) name7369 (
		\wishbone_bd_ram_mem2_reg[248][21]/P0001 ,
		_w11952_,
		_w11990_,
		_w17882_
	);
	LUT3 #(
		.INIT('h80)
	) name7370 (
		\wishbone_bd_ram_mem2_reg[189][21]/P0001 ,
		_w11942_,
		_w11966_,
		_w17883_
	);
	LUT3 #(
		.INIT('h80)
	) name7371 (
		\wishbone_bd_ram_mem2_reg[174][21]/P0001 ,
		_w11930_,
		_w11948_,
		_w17884_
	);
	LUT4 #(
		.INIT('h0001)
	) name7372 (
		_w17881_,
		_w17882_,
		_w17883_,
		_w17884_,
		_w17885_
	);
	LUT4 #(
		.INIT('h8000)
	) name7373 (
		_w17870_,
		_w17875_,
		_w17880_,
		_w17885_,
		_w17886_
	);
	LUT4 #(
		.INIT('h8000)
	) name7374 (
		_w17823_,
		_w17844_,
		_w17865_,
		_w17886_,
		_w17887_
	);
	LUT3 #(
		.INIT('h80)
	) name7375 (
		\wishbone_bd_ram_mem2_reg[42][21]/P0001 ,
		_w11944_,
		_w11957_,
		_w17888_
	);
	LUT3 #(
		.INIT('h80)
	) name7376 (
		\wishbone_bd_ram_mem2_reg[26][21]/P0001 ,
		_w11935_,
		_w11944_,
		_w17889_
	);
	LUT3 #(
		.INIT('h80)
	) name7377 (
		\wishbone_bd_ram_mem2_reg[152][21]/P0001 ,
		_w11959_,
		_w11990_,
		_w17890_
	);
	LUT3 #(
		.INIT('h80)
	) name7378 (
		\wishbone_bd_ram_mem2_reg[233][21]/P0001 ,
		_w11968_,
		_w11982_,
		_w17891_
	);
	LUT4 #(
		.INIT('h0001)
	) name7379 (
		_w17888_,
		_w17889_,
		_w17890_,
		_w17891_,
		_w17892_
	);
	LUT3 #(
		.INIT('h80)
	) name7380 (
		\wishbone_bd_ram_mem2_reg[12][21]/P0001 ,
		_w11932_,
		_w11954_,
		_w17893_
	);
	LUT3 #(
		.INIT('h80)
	) name7381 (
		\wishbone_bd_ram_mem2_reg[20][21]/P0001 ,
		_w11929_,
		_w11935_,
		_w17894_
	);
	LUT3 #(
		.INIT('h80)
	) name7382 (
		\wishbone_bd_ram_mem2_reg[221][21]/P0001 ,
		_w11966_,
		_w11984_,
		_w17895_
	);
	LUT3 #(
		.INIT('h80)
	) name7383 (
		\wishbone_bd_ram_mem2_reg[35][21]/P0001 ,
		_w11938_,
		_w11957_,
		_w17896_
	);
	LUT4 #(
		.INIT('h0001)
	) name7384 (
		_w17893_,
		_w17894_,
		_w17895_,
		_w17896_,
		_w17897_
	);
	LUT3 #(
		.INIT('h80)
	) name7385 (
		\wishbone_bd_ram_mem2_reg[84][21]/P0001 ,
		_w11929_,
		_w11972_,
		_w17898_
	);
	LUT3 #(
		.INIT('h80)
	) name7386 (
		\wishbone_bd_ram_mem2_reg[153][21]/P0001 ,
		_w11959_,
		_w11968_,
		_w17899_
	);
	LUT3 #(
		.INIT('h80)
	) name7387 (
		\wishbone_bd_ram_mem2_reg[106][21]/P0001 ,
		_w11944_,
		_w11965_,
		_w17900_
	);
	LUT3 #(
		.INIT('h80)
	) name7388 (
		\wishbone_bd_ram_mem2_reg[92][21]/P0001 ,
		_w11954_,
		_w11972_,
		_w17901_
	);
	LUT4 #(
		.INIT('h0001)
	) name7389 (
		_w17898_,
		_w17899_,
		_w17900_,
		_w17901_,
		_w17902_
	);
	LUT3 #(
		.INIT('h80)
	) name7390 (
		\wishbone_bd_ram_mem2_reg[160][21]/P0001 ,
		_w11930_,
		_w11941_,
		_w17903_
	);
	LUT3 #(
		.INIT('h80)
	) name7391 (
		\wishbone_bd_ram_mem2_reg[61][21]/P0001 ,
		_w11966_,
		_w11979_,
		_w17904_
	);
	LUT3 #(
		.INIT('h80)
	) name7392 (
		\wishbone_bd_ram_mem2_reg[136][21]/P0001 ,
		_w11955_,
		_w11990_,
		_w17905_
	);
	LUT3 #(
		.INIT('h80)
	) name7393 (
		\wishbone_bd_ram_mem2_reg[41][21]/P0001 ,
		_w11957_,
		_w11968_,
		_w17906_
	);
	LUT4 #(
		.INIT('h0001)
	) name7394 (
		_w17903_,
		_w17904_,
		_w17905_,
		_w17906_,
		_w17907_
	);
	LUT4 #(
		.INIT('h8000)
	) name7395 (
		_w17892_,
		_w17897_,
		_w17902_,
		_w17907_,
		_w17908_
	);
	LUT3 #(
		.INIT('h80)
	) name7396 (
		\wishbone_bd_ram_mem2_reg[201][21]/P0001 ,
		_w11945_,
		_w11968_,
		_w17909_
	);
	LUT3 #(
		.INIT('h80)
	) name7397 (
		\wishbone_bd_ram_mem2_reg[33][21]/P0001 ,
		_w11957_,
		_w11977_,
		_w17910_
	);
	LUT3 #(
		.INIT('h80)
	) name7398 (
		\wishbone_bd_ram_mem2_reg[223][21]/P0001 ,
		_w11973_,
		_w11984_,
		_w17911_
	);
	LUT3 #(
		.INIT('h80)
	) name7399 (
		\wishbone_bd_ram_mem2_reg[72][21]/P0001 ,
		_w11949_,
		_w11990_,
		_w17912_
	);
	LUT4 #(
		.INIT('h0001)
	) name7400 (
		_w17909_,
		_w17910_,
		_w17911_,
		_w17912_,
		_w17913_
	);
	LUT3 #(
		.INIT('h80)
	) name7401 (
		\wishbone_bd_ram_mem2_reg[76][21]/P0001 ,
		_w11949_,
		_w11954_,
		_w17914_
	);
	LUT3 #(
		.INIT('h80)
	) name7402 (
		\wishbone_bd_ram_mem2_reg[75][21]/P0001 ,
		_w11936_,
		_w11949_,
		_w17915_
	);
	LUT3 #(
		.INIT('h80)
	) name7403 (
		\wishbone_bd_ram_mem2_reg[71][21]/P0001 ,
		_w11949_,
		_w11975_,
		_w17916_
	);
	LUT3 #(
		.INIT('h80)
	) name7404 (
		\wishbone_bd_ram_mem2_reg[105][21]/P0001 ,
		_w11965_,
		_w11968_,
		_w17917_
	);
	LUT4 #(
		.INIT('h0001)
	) name7405 (
		_w17914_,
		_w17915_,
		_w17916_,
		_w17917_,
		_w17918_
	);
	LUT3 #(
		.INIT('h80)
	) name7406 (
		\wishbone_bd_ram_mem2_reg[236][21]/P0001 ,
		_w11954_,
		_w11982_,
		_w17919_
	);
	LUT3 #(
		.INIT('h80)
	) name7407 (
		\wishbone_bd_ram_mem2_reg[199][21]/P0001 ,
		_w11945_,
		_w11975_,
		_w17920_
	);
	LUT3 #(
		.INIT('h80)
	) name7408 (
		\wishbone_bd_ram_mem2_reg[66][21]/P0001 ,
		_w11949_,
		_w11963_,
		_w17921_
	);
	LUT3 #(
		.INIT('h80)
	) name7409 (
		\wishbone_bd_ram_mem2_reg[31][21]/P0001 ,
		_w11935_,
		_w11973_,
		_w17922_
	);
	LUT4 #(
		.INIT('h0001)
	) name7410 (
		_w17919_,
		_w17920_,
		_w17921_,
		_w17922_,
		_w17923_
	);
	LUT3 #(
		.INIT('h80)
	) name7411 (
		\wishbone_bd_ram_mem2_reg[188][21]/P0001 ,
		_w11942_,
		_w11954_,
		_w17924_
	);
	LUT3 #(
		.INIT('h80)
	) name7412 (
		\wishbone_bd_ram_mem2_reg[158][21]/P0001 ,
		_w11948_,
		_w11959_,
		_w17925_
	);
	LUT3 #(
		.INIT('h80)
	) name7413 (
		\wishbone_bd_ram_mem2_reg[239][21]/P0001 ,
		_w11973_,
		_w11982_,
		_w17926_
	);
	LUT3 #(
		.INIT('h80)
	) name7414 (
		\wishbone_bd_ram_mem2_reg[91][21]/P0001 ,
		_w11936_,
		_w11972_,
		_w17927_
	);
	LUT4 #(
		.INIT('h0001)
	) name7415 (
		_w17924_,
		_w17925_,
		_w17926_,
		_w17927_,
		_w17928_
	);
	LUT4 #(
		.INIT('h8000)
	) name7416 (
		_w17913_,
		_w17918_,
		_w17923_,
		_w17928_,
		_w17929_
	);
	LUT3 #(
		.INIT('h80)
	) name7417 (
		\wishbone_bd_ram_mem2_reg[240][21]/P0001 ,
		_w11941_,
		_w11952_,
		_w17930_
	);
	LUT3 #(
		.INIT('h80)
	) name7418 (
		\wishbone_bd_ram_mem2_reg[32][21]/P0001 ,
		_w11941_,
		_w11957_,
		_w17931_
	);
	LUT3 #(
		.INIT('h80)
	) name7419 (
		\wishbone_bd_ram_mem2_reg[88][21]/P0001 ,
		_w11972_,
		_w11990_,
		_w17932_
	);
	LUT3 #(
		.INIT('h80)
	) name7420 (
		\wishbone_bd_ram_mem2_reg[205][21]/P0001 ,
		_w11945_,
		_w11966_,
		_w17933_
	);
	LUT4 #(
		.INIT('h0001)
	) name7421 (
		_w17930_,
		_w17931_,
		_w17932_,
		_w17933_,
		_w17934_
	);
	LUT3 #(
		.INIT('h80)
	) name7422 (
		\wishbone_bd_ram_mem2_reg[219][21]/P0001 ,
		_w11936_,
		_w11984_,
		_w17935_
	);
	LUT3 #(
		.INIT('h80)
	) name7423 (
		\wishbone_bd_ram_mem2_reg[103][21]/P0001 ,
		_w11965_,
		_w11975_,
		_w17936_
	);
	LUT3 #(
		.INIT('h80)
	) name7424 (
		\wishbone_bd_ram_mem2_reg[245][21]/P0001 ,
		_w11933_,
		_w11952_,
		_w17937_
	);
	LUT3 #(
		.INIT('h80)
	) name7425 (
		\wishbone_bd_ram_mem2_reg[251][21]/P0001 ,
		_w11936_,
		_w11952_,
		_w17938_
	);
	LUT4 #(
		.INIT('h0001)
	) name7426 (
		_w17935_,
		_w17936_,
		_w17937_,
		_w17938_,
		_w17939_
	);
	LUT3 #(
		.INIT('h80)
	) name7427 (
		\wishbone_bd_ram_mem2_reg[96][21]/P0001 ,
		_w11941_,
		_w11965_,
		_w17940_
	);
	LUT3 #(
		.INIT('h80)
	) name7428 (
		\wishbone_bd_ram_mem2_reg[228][21]/P0001 ,
		_w11929_,
		_w11982_,
		_w17941_
	);
	LUT3 #(
		.INIT('h80)
	) name7429 (
		\wishbone_bd_ram_mem2_reg[18][21]/P0001 ,
		_w11935_,
		_w11963_,
		_w17942_
	);
	LUT3 #(
		.INIT('h80)
	) name7430 (
		\wishbone_bd_ram_mem2_reg[126][21]/P0001 ,
		_w11948_,
		_w12012_,
		_w17943_
	);
	LUT4 #(
		.INIT('h0001)
	) name7431 (
		_w17940_,
		_w17941_,
		_w17942_,
		_w17943_,
		_w17944_
	);
	LUT3 #(
		.INIT('h80)
	) name7432 (
		\wishbone_bd_ram_mem2_reg[161][21]/P0001 ,
		_w11930_,
		_w11977_,
		_w17945_
	);
	LUT3 #(
		.INIT('h80)
	) name7433 (
		\wishbone_bd_ram_mem2_reg[36][21]/P0001 ,
		_w11929_,
		_w11957_,
		_w17946_
	);
	LUT3 #(
		.INIT('h80)
	) name7434 (
		\wishbone_bd_ram_mem2_reg[55][21]/P0001 ,
		_w11975_,
		_w11979_,
		_w17947_
	);
	LUT3 #(
		.INIT('h80)
	) name7435 (
		\wishbone_bd_ram_mem2_reg[215][21]/P0001 ,
		_w11975_,
		_w11984_,
		_w17948_
	);
	LUT4 #(
		.INIT('h0001)
	) name7436 (
		_w17945_,
		_w17946_,
		_w17947_,
		_w17948_,
		_w17949_
	);
	LUT4 #(
		.INIT('h8000)
	) name7437 (
		_w17934_,
		_w17939_,
		_w17944_,
		_w17949_,
		_w17950_
	);
	LUT3 #(
		.INIT('h80)
	) name7438 (
		\wishbone_bd_ram_mem2_reg[118][21]/P0001 ,
		_w11986_,
		_w12012_,
		_w17951_
	);
	LUT3 #(
		.INIT('h80)
	) name7439 (
		\wishbone_bd_ram_mem2_reg[16][21]/P0001 ,
		_w11935_,
		_w11941_,
		_w17952_
	);
	LUT3 #(
		.INIT('h80)
	) name7440 (
		\wishbone_bd_ram_mem2_reg[6][21]/P0001 ,
		_w11932_,
		_w11986_,
		_w17953_
	);
	LUT3 #(
		.INIT('h80)
	) name7441 (
		\wishbone_bd_ram_mem2_reg[139][21]/P0001 ,
		_w11936_,
		_w11955_,
		_w17954_
	);
	LUT4 #(
		.INIT('h0001)
	) name7442 (
		_w17951_,
		_w17952_,
		_w17953_,
		_w17954_,
		_w17955_
	);
	LUT3 #(
		.INIT('h80)
	) name7443 (
		\wishbone_bd_ram_mem2_reg[98][21]/P0001 ,
		_w11963_,
		_w11965_,
		_w17956_
	);
	LUT3 #(
		.INIT('h80)
	) name7444 (
		\wishbone_bd_ram_mem2_reg[200][21]/P0001 ,
		_w11945_,
		_w11990_,
		_w17957_
	);
	LUT3 #(
		.INIT('h80)
	) name7445 (
		\wishbone_bd_ram_mem2_reg[59][21]/P0001 ,
		_w11936_,
		_w11979_,
		_w17958_
	);
	LUT3 #(
		.INIT('h80)
	) name7446 (
		\wishbone_bd_ram_mem2_reg[113][21]/P0001 ,
		_w11977_,
		_w12012_,
		_w17959_
	);
	LUT4 #(
		.INIT('h0001)
	) name7447 (
		_w17956_,
		_w17957_,
		_w17958_,
		_w17959_,
		_w17960_
	);
	LUT3 #(
		.INIT('h80)
	) name7448 (
		\wishbone_bd_ram_mem2_reg[253][21]/P0001 ,
		_w11952_,
		_w11966_,
		_w17961_
	);
	LUT3 #(
		.INIT('h80)
	) name7449 (
		\wishbone_bd_ram_mem2_reg[39][21]/P0001 ,
		_w11957_,
		_w11975_,
		_w17962_
	);
	LUT3 #(
		.INIT('h80)
	) name7450 (
		\wishbone_bd_ram_mem2_reg[194][21]/P0001 ,
		_w11945_,
		_w11963_,
		_w17963_
	);
	LUT3 #(
		.INIT('h80)
	) name7451 (
		\wishbone_bd_ram_mem2_reg[133][21]/P0001 ,
		_w11933_,
		_w11955_,
		_w17964_
	);
	LUT4 #(
		.INIT('h0001)
	) name7452 (
		_w17961_,
		_w17962_,
		_w17963_,
		_w17964_,
		_w17965_
	);
	LUT3 #(
		.INIT('h80)
	) name7453 (
		\wishbone_bd_ram_mem2_reg[97][21]/P0001 ,
		_w11965_,
		_w11977_,
		_w17966_
	);
	LUT3 #(
		.INIT('h80)
	) name7454 (
		\wishbone_bd_ram_mem2_reg[89][21]/P0001 ,
		_w11968_,
		_w11972_,
		_w17967_
	);
	LUT3 #(
		.INIT('h80)
	) name7455 (
		\wishbone_bd_ram_mem2_reg[0][21]/P0001 ,
		_w11932_,
		_w11941_,
		_w17968_
	);
	LUT3 #(
		.INIT('h80)
	) name7456 (
		\wishbone_bd_ram_mem2_reg[107][21]/P0001 ,
		_w11936_,
		_w11965_,
		_w17969_
	);
	LUT4 #(
		.INIT('h0001)
	) name7457 (
		_w17966_,
		_w17967_,
		_w17968_,
		_w17969_,
		_w17970_
	);
	LUT4 #(
		.INIT('h8000)
	) name7458 (
		_w17955_,
		_w17960_,
		_w17965_,
		_w17970_,
		_w17971_
	);
	LUT4 #(
		.INIT('h8000)
	) name7459 (
		_w17908_,
		_w17929_,
		_w17950_,
		_w17971_,
		_w17972_
	);
	LUT3 #(
		.INIT('h80)
	) name7460 (
		\wishbone_bd_ram_mem2_reg[13][21]/P0001 ,
		_w11932_,
		_w11966_,
		_w17973_
	);
	LUT3 #(
		.INIT('h80)
	) name7461 (
		\wishbone_bd_ram_mem2_reg[241][21]/P0001 ,
		_w11952_,
		_w11977_,
		_w17974_
	);
	LUT3 #(
		.INIT('h80)
	) name7462 (
		\wishbone_bd_ram_mem2_reg[167][21]/P0001 ,
		_w11930_,
		_w11975_,
		_w17975_
	);
	LUT3 #(
		.INIT('h80)
	) name7463 (
		\wishbone_bd_ram_mem2_reg[53][21]/P0001 ,
		_w11933_,
		_w11979_,
		_w17976_
	);
	LUT4 #(
		.INIT('h0001)
	) name7464 (
		_w17973_,
		_w17974_,
		_w17975_,
		_w17976_,
		_w17977_
	);
	LUT3 #(
		.INIT('h80)
	) name7465 (
		\wishbone_bd_ram_mem2_reg[135][21]/P0001 ,
		_w11955_,
		_w11975_,
		_w17978_
	);
	LUT3 #(
		.INIT('h80)
	) name7466 (
		\wishbone_bd_ram_mem2_reg[46][21]/P0001 ,
		_w11948_,
		_w11957_,
		_w17979_
	);
	LUT3 #(
		.INIT('h80)
	) name7467 (
		\wishbone_bd_ram_mem2_reg[47][21]/P0001 ,
		_w11957_,
		_w11973_,
		_w17980_
	);
	LUT3 #(
		.INIT('h80)
	) name7468 (
		\wishbone_bd_ram_mem2_reg[132][21]/P0001 ,
		_w11929_,
		_w11955_,
		_w17981_
	);
	LUT4 #(
		.INIT('h0001)
	) name7469 (
		_w17978_,
		_w17979_,
		_w17980_,
		_w17981_,
		_w17982_
	);
	LUT3 #(
		.INIT('h80)
	) name7470 (
		\wishbone_bd_ram_mem2_reg[83][21]/P0001 ,
		_w11938_,
		_w11972_,
		_w17983_
	);
	LUT3 #(
		.INIT('h80)
	) name7471 (
		\wishbone_bd_ram_mem2_reg[252][21]/P0001 ,
		_w11952_,
		_w11954_,
		_w17984_
	);
	LUT3 #(
		.INIT('h80)
	) name7472 (
		\wishbone_bd_ram_mem2_reg[154][21]/P0001 ,
		_w11944_,
		_w11959_,
		_w17985_
	);
	LUT3 #(
		.INIT('h80)
	) name7473 (
		\wishbone_bd_ram_mem2_reg[231][21]/P0001 ,
		_w11975_,
		_w11982_,
		_w17986_
	);
	LUT4 #(
		.INIT('h0001)
	) name7474 (
		_w17983_,
		_w17984_,
		_w17985_,
		_w17986_,
		_w17987_
	);
	LUT3 #(
		.INIT('h80)
	) name7475 (
		\wishbone_bd_ram_mem2_reg[227][21]/P0001 ,
		_w11938_,
		_w11982_,
		_w17988_
	);
	LUT3 #(
		.INIT('h80)
	) name7476 (
		\wishbone_bd_ram_mem2_reg[34][21]/P0001 ,
		_w11957_,
		_w11963_,
		_w17989_
	);
	LUT3 #(
		.INIT('h80)
	) name7477 (
		\wishbone_bd_ram_mem2_reg[11][21]/P0001 ,
		_w11932_,
		_w11936_,
		_w17990_
	);
	LUT3 #(
		.INIT('h80)
	) name7478 (
		\wishbone_bd_ram_mem2_reg[131][21]/P0001 ,
		_w11938_,
		_w11955_,
		_w17991_
	);
	LUT4 #(
		.INIT('h0001)
	) name7479 (
		_w17988_,
		_w17989_,
		_w17990_,
		_w17991_,
		_w17992_
	);
	LUT4 #(
		.INIT('h8000)
	) name7480 (
		_w17977_,
		_w17982_,
		_w17987_,
		_w17992_,
		_w17993_
	);
	LUT3 #(
		.INIT('h80)
	) name7481 (
		\wishbone_bd_ram_mem2_reg[57][21]/P0001 ,
		_w11968_,
		_w11979_,
		_w17994_
	);
	LUT3 #(
		.INIT('h80)
	) name7482 (
		\wishbone_bd_ram_mem2_reg[123][21]/P0001 ,
		_w11936_,
		_w12012_,
		_w17995_
	);
	LUT3 #(
		.INIT('h80)
	) name7483 (
		\wishbone_bd_ram_mem2_reg[3][21]/P0001 ,
		_w11932_,
		_w11938_,
		_w17996_
	);
	LUT3 #(
		.INIT('h80)
	) name7484 (
		\wishbone_bd_ram_mem2_reg[130][21]/P0001 ,
		_w11955_,
		_w11963_,
		_w17997_
	);
	LUT4 #(
		.INIT('h0001)
	) name7485 (
		_w17994_,
		_w17995_,
		_w17996_,
		_w17997_,
		_w17998_
	);
	LUT3 #(
		.INIT('h80)
	) name7486 (
		\wishbone_bd_ram_mem2_reg[224][21]/P0001 ,
		_w11941_,
		_w11982_,
		_w17999_
	);
	LUT3 #(
		.INIT('h80)
	) name7487 (
		\wishbone_bd_ram_mem2_reg[54][21]/P0001 ,
		_w11979_,
		_w11986_,
		_w18000_
	);
	LUT3 #(
		.INIT('h80)
	) name7488 (
		\wishbone_bd_ram_mem2_reg[137][21]/P0001 ,
		_w11955_,
		_w11968_,
		_w18001_
	);
	LUT3 #(
		.INIT('h80)
	) name7489 (
		\wishbone_bd_ram_mem2_reg[172][21]/P0001 ,
		_w11930_,
		_w11954_,
		_w18002_
	);
	LUT4 #(
		.INIT('h0001)
	) name7490 (
		_w17999_,
		_w18000_,
		_w18001_,
		_w18002_,
		_w18003_
	);
	LUT3 #(
		.INIT('h80)
	) name7491 (
		\wishbone_bd_ram_mem2_reg[56][21]/P0001 ,
		_w11979_,
		_w11990_,
		_w18004_
	);
	LUT3 #(
		.INIT('h80)
	) name7492 (
		\wishbone_bd_ram_mem2_reg[150][21]/P0001 ,
		_w11959_,
		_w11986_,
		_w18005_
	);
	LUT3 #(
		.INIT('h80)
	) name7493 (
		\wishbone_bd_ram_mem2_reg[74][21]/P0001 ,
		_w11944_,
		_w11949_,
		_w18006_
	);
	LUT3 #(
		.INIT('h80)
	) name7494 (
		\wishbone_bd_ram_mem2_reg[79][21]/P0001 ,
		_w11949_,
		_w11973_,
		_w18007_
	);
	LUT4 #(
		.INIT('h0001)
	) name7495 (
		_w18004_,
		_w18005_,
		_w18006_,
		_w18007_,
		_w18008_
	);
	LUT3 #(
		.INIT('h80)
	) name7496 (
		\wishbone_bd_ram_mem2_reg[244][21]/P0001 ,
		_w11929_,
		_w11952_,
		_w18009_
	);
	LUT3 #(
		.INIT('h80)
	) name7497 (
		\wishbone_bd_ram_mem2_reg[49][21]/P0001 ,
		_w11977_,
		_w11979_,
		_w18010_
	);
	LUT3 #(
		.INIT('h80)
	) name7498 (
		\wishbone_bd_ram_mem2_reg[217][21]/P0001 ,
		_w11968_,
		_w11984_,
		_w18011_
	);
	LUT3 #(
		.INIT('h80)
	) name7499 (
		\wishbone_bd_ram_mem2_reg[138][21]/P0001 ,
		_w11944_,
		_w11955_,
		_w18012_
	);
	LUT4 #(
		.INIT('h0001)
	) name7500 (
		_w18009_,
		_w18010_,
		_w18011_,
		_w18012_,
		_w18013_
	);
	LUT4 #(
		.INIT('h8000)
	) name7501 (
		_w17998_,
		_w18003_,
		_w18008_,
		_w18013_,
		_w18014_
	);
	LUT3 #(
		.INIT('h80)
	) name7502 (
		\wishbone_bd_ram_mem2_reg[185][21]/P0001 ,
		_w11942_,
		_w11968_,
		_w18015_
	);
	LUT3 #(
		.INIT('h80)
	) name7503 (
		\wishbone_bd_ram_mem2_reg[43][21]/P0001 ,
		_w11936_,
		_w11957_,
		_w18016_
	);
	LUT3 #(
		.INIT('h80)
	) name7504 (
		\wishbone_bd_ram_mem2_reg[69][21]/P0001 ,
		_w11933_,
		_w11949_,
		_w18017_
	);
	LUT3 #(
		.INIT('h80)
	) name7505 (
		\wishbone_bd_ram_mem2_reg[249][21]/P0001 ,
		_w11952_,
		_w11968_,
		_w18018_
	);
	LUT4 #(
		.INIT('h0001)
	) name7506 (
		_w18015_,
		_w18016_,
		_w18017_,
		_w18018_,
		_w18019_
	);
	LUT3 #(
		.INIT('h80)
	) name7507 (
		\wishbone_bd_ram_mem2_reg[29][21]/P0001 ,
		_w11935_,
		_w11966_,
		_w18020_
	);
	LUT3 #(
		.INIT('h80)
	) name7508 (
		\wishbone_bd_ram_mem2_reg[110][21]/P0001 ,
		_w11948_,
		_w11965_,
		_w18021_
	);
	LUT3 #(
		.INIT('h80)
	) name7509 (
		\wishbone_bd_ram_mem2_reg[19][21]/P0001 ,
		_w11935_,
		_w11938_,
		_w18022_
	);
	LUT3 #(
		.INIT('h80)
	) name7510 (
		\wishbone_bd_ram_mem2_reg[204][21]/P0001 ,
		_w11945_,
		_w11954_,
		_w18023_
	);
	LUT4 #(
		.INIT('h0001)
	) name7511 (
		_w18020_,
		_w18021_,
		_w18022_,
		_w18023_,
		_w18024_
	);
	LUT3 #(
		.INIT('h80)
	) name7512 (
		\wishbone_bd_ram_mem2_reg[4][21]/P0001 ,
		_w11929_,
		_w11932_,
		_w18025_
	);
	LUT3 #(
		.INIT('h80)
	) name7513 (
		\wishbone_bd_ram_mem2_reg[202][21]/P0001 ,
		_w11944_,
		_w11945_,
		_w18026_
	);
	LUT3 #(
		.INIT('h80)
	) name7514 (
		\wishbone_bd_ram_mem2_reg[235][21]/P0001 ,
		_w11936_,
		_w11982_,
		_w18027_
	);
	LUT3 #(
		.INIT('h80)
	) name7515 (
		\wishbone_bd_ram_mem2_reg[159][21]/P0001 ,
		_w11959_,
		_w11973_,
		_w18028_
	);
	LUT4 #(
		.INIT('h0001)
	) name7516 (
		_w18025_,
		_w18026_,
		_w18027_,
		_w18028_,
		_w18029_
	);
	LUT3 #(
		.INIT('h80)
	) name7517 (
		\wishbone_bd_ram_mem2_reg[187][21]/P0001 ,
		_w11936_,
		_w11942_,
		_w18030_
	);
	LUT3 #(
		.INIT('h80)
	) name7518 (
		\wishbone_bd_ram_mem2_reg[67][21]/P0001 ,
		_w11938_,
		_w11949_,
		_w18031_
	);
	LUT3 #(
		.INIT('h80)
	) name7519 (
		\wishbone_bd_ram_mem2_reg[73][21]/P0001 ,
		_w11949_,
		_w11968_,
		_w18032_
	);
	LUT3 #(
		.INIT('h80)
	) name7520 (
		\wishbone_bd_ram_mem2_reg[197][21]/P0001 ,
		_w11933_,
		_w11945_,
		_w18033_
	);
	LUT4 #(
		.INIT('h0001)
	) name7521 (
		_w18030_,
		_w18031_,
		_w18032_,
		_w18033_,
		_w18034_
	);
	LUT4 #(
		.INIT('h8000)
	) name7522 (
		_w18019_,
		_w18024_,
		_w18029_,
		_w18034_,
		_w18035_
	);
	LUT3 #(
		.INIT('h80)
	) name7523 (
		\wishbone_bd_ram_mem2_reg[146][21]/P0001 ,
		_w11959_,
		_w11963_,
		_w18036_
	);
	LUT3 #(
		.INIT('h80)
	) name7524 (
		\wishbone_bd_ram_mem2_reg[124][21]/P0001 ,
		_w11954_,
		_w12012_,
		_w18037_
	);
	LUT3 #(
		.INIT('h80)
	) name7525 (
		\wishbone_bd_ram_mem2_reg[164][21]/P0001 ,
		_w11929_,
		_w11930_,
		_w18038_
	);
	LUT3 #(
		.INIT('h80)
	) name7526 (
		\wishbone_bd_ram_mem2_reg[52][21]/P0001 ,
		_w11929_,
		_w11979_,
		_w18039_
	);
	LUT4 #(
		.INIT('h0001)
	) name7527 (
		_w18036_,
		_w18037_,
		_w18038_,
		_w18039_,
		_w18040_
	);
	LUT3 #(
		.INIT('h80)
	) name7528 (
		\wishbone_bd_ram_mem2_reg[216][21]/P0001 ,
		_w11984_,
		_w11990_,
		_w18041_
	);
	LUT3 #(
		.INIT('h80)
	) name7529 (
		\wishbone_bd_ram_mem2_reg[170][21]/P0001 ,
		_w11930_,
		_w11944_,
		_w18042_
	);
	LUT3 #(
		.INIT('h80)
	) name7530 (
		\wishbone_bd_ram_mem2_reg[142][21]/P0001 ,
		_w11948_,
		_w11955_,
		_w18043_
	);
	LUT3 #(
		.INIT('h80)
	) name7531 (
		\wishbone_bd_ram_mem2_reg[140][21]/P0001 ,
		_w11954_,
		_w11955_,
		_w18044_
	);
	LUT4 #(
		.INIT('h0001)
	) name7532 (
		_w18041_,
		_w18042_,
		_w18043_,
		_w18044_,
		_w18045_
	);
	LUT3 #(
		.INIT('h80)
	) name7533 (
		\wishbone_bd_ram_mem2_reg[250][21]/P0001 ,
		_w11944_,
		_w11952_,
		_w18046_
	);
	LUT3 #(
		.INIT('h80)
	) name7534 (
		\wishbone_bd_ram_mem2_reg[225][21]/P0001 ,
		_w11977_,
		_w11982_,
		_w18047_
	);
	LUT3 #(
		.INIT('h80)
	) name7535 (
		\wishbone_bd_ram_mem2_reg[112][21]/P0001 ,
		_w11941_,
		_w12012_,
		_w18048_
	);
	LUT3 #(
		.INIT('h80)
	) name7536 (
		\wishbone_bd_ram_mem2_reg[25][21]/P0001 ,
		_w11935_,
		_w11968_,
		_w18049_
	);
	LUT4 #(
		.INIT('h0001)
	) name7537 (
		_w18046_,
		_w18047_,
		_w18048_,
		_w18049_,
		_w18050_
	);
	LUT3 #(
		.INIT('h80)
	) name7538 (
		\wishbone_bd_ram_mem2_reg[163][21]/P0001 ,
		_w11930_,
		_w11938_,
		_w18051_
	);
	LUT3 #(
		.INIT('h80)
	) name7539 (
		\wishbone_bd_ram_mem2_reg[218][21]/P0001 ,
		_w11944_,
		_w11984_,
		_w18052_
	);
	LUT3 #(
		.INIT('h80)
	) name7540 (
		\wishbone_bd_ram_mem2_reg[180][21]/P0001 ,
		_w11929_,
		_w11942_,
		_w18053_
	);
	LUT3 #(
		.INIT('h80)
	) name7541 (
		\wishbone_bd_ram_mem2_reg[86][21]/P0001 ,
		_w11972_,
		_w11986_,
		_w18054_
	);
	LUT4 #(
		.INIT('h0001)
	) name7542 (
		_w18051_,
		_w18052_,
		_w18053_,
		_w18054_,
		_w18055_
	);
	LUT4 #(
		.INIT('h8000)
	) name7543 (
		_w18040_,
		_w18045_,
		_w18050_,
		_w18055_,
		_w18056_
	);
	LUT4 #(
		.INIT('h8000)
	) name7544 (
		_w17993_,
		_w18014_,
		_w18035_,
		_w18056_,
		_w18057_
	);
	LUT4 #(
		.INIT('h8000)
	) name7545 (
		_w17802_,
		_w17887_,
		_w17972_,
		_w18057_,
		_w18058_
	);
	LUT3 #(
		.INIT('hce)
	) name7546 (
		_w12303_,
		_w17717_,
		_w18058_,
		_w18059_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name7547 (
		\wishbone_LatchedTxLength_reg[7]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w18060_
	);
	LUT3 #(
		.INIT('h80)
	) name7548 (
		\wishbone_bd_ram_mem2_reg[38][23]/P0001 ,
		_w11957_,
		_w11986_,
		_w18061_
	);
	LUT3 #(
		.INIT('h80)
	) name7549 (
		\wishbone_bd_ram_mem2_reg[85][23]/P0001 ,
		_w11933_,
		_w11972_,
		_w18062_
	);
	LUT3 #(
		.INIT('h80)
	) name7550 (
		\wishbone_bd_ram_mem2_reg[50][23]/P0001 ,
		_w11963_,
		_w11979_,
		_w18063_
	);
	LUT3 #(
		.INIT('h80)
	) name7551 (
		\wishbone_bd_ram_mem2_reg[31][23]/P0001 ,
		_w11935_,
		_w11973_,
		_w18064_
	);
	LUT4 #(
		.INIT('h0001)
	) name7552 (
		_w18061_,
		_w18062_,
		_w18063_,
		_w18064_,
		_w18065_
	);
	LUT3 #(
		.INIT('h80)
	) name7553 (
		\wishbone_bd_ram_mem2_reg[139][23]/P0001 ,
		_w11936_,
		_w11955_,
		_w18066_
	);
	LUT3 #(
		.INIT('h80)
	) name7554 (
		\wishbone_bd_ram_mem2_reg[35][23]/P0001 ,
		_w11938_,
		_w11957_,
		_w18067_
	);
	LUT3 #(
		.INIT('h80)
	) name7555 (
		\wishbone_bd_ram_mem2_reg[5][23]/P0001 ,
		_w11932_,
		_w11933_,
		_w18068_
	);
	LUT3 #(
		.INIT('h80)
	) name7556 (
		\wishbone_bd_ram_mem2_reg[199][23]/P0001 ,
		_w11945_,
		_w11975_,
		_w18069_
	);
	LUT4 #(
		.INIT('h0001)
	) name7557 (
		_w18066_,
		_w18067_,
		_w18068_,
		_w18069_,
		_w18070_
	);
	LUT3 #(
		.INIT('h80)
	) name7558 (
		\wishbone_bd_ram_mem2_reg[202][23]/P0001 ,
		_w11944_,
		_w11945_,
		_w18071_
	);
	LUT3 #(
		.INIT('h80)
	) name7559 (
		\wishbone_bd_ram_mem2_reg[191][23]/P0001 ,
		_w11942_,
		_w11973_,
		_w18072_
	);
	LUT3 #(
		.INIT('h80)
	) name7560 (
		\wishbone_bd_ram_mem2_reg[68][23]/P0001 ,
		_w11929_,
		_w11949_,
		_w18073_
	);
	LUT3 #(
		.INIT('h80)
	) name7561 (
		\wishbone_bd_ram_mem2_reg[228][23]/P0001 ,
		_w11929_,
		_w11982_,
		_w18074_
	);
	LUT4 #(
		.INIT('h0001)
	) name7562 (
		_w18071_,
		_w18072_,
		_w18073_,
		_w18074_,
		_w18075_
	);
	LUT3 #(
		.INIT('h80)
	) name7563 (
		\wishbone_bd_ram_mem2_reg[11][23]/P0001 ,
		_w11932_,
		_w11936_,
		_w18076_
	);
	LUT3 #(
		.INIT('h80)
	) name7564 (
		\wishbone_bd_ram_mem2_reg[178][23]/P0001 ,
		_w11942_,
		_w11963_,
		_w18077_
	);
	LUT3 #(
		.INIT('h80)
	) name7565 (
		\wishbone_bd_ram_mem2_reg[210][23]/P0001 ,
		_w11963_,
		_w11984_,
		_w18078_
	);
	LUT3 #(
		.INIT('h80)
	) name7566 (
		\wishbone_bd_ram_mem2_reg[231][23]/P0001 ,
		_w11975_,
		_w11982_,
		_w18079_
	);
	LUT4 #(
		.INIT('h0001)
	) name7567 (
		_w18076_,
		_w18077_,
		_w18078_,
		_w18079_,
		_w18080_
	);
	LUT4 #(
		.INIT('h8000)
	) name7568 (
		_w18065_,
		_w18070_,
		_w18075_,
		_w18080_,
		_w18081_
	);
	LUT3 #(
		.INIT('h80)
	) name7569 (
		\wishbone_bd_ram_mem2_reg[88][23]/P0001 ,
		_w11972_,
		_w11990_,
		_w18082_
	);
	LUT3 #(
		.INIT('h80)
	) name7570 (
		\wishbone_bd_ram_mem2_reg[103][23]/P0001 ,
		_w11965_,
		_w11975_,
		_w18083_
	);
	LUT3 #(
		.INIT('h80)
	) name7571 (
		\wishbone_bd_ram_mem2_reg[61][23]/P0001 ,
		_w11966_,
		_w11979_,
		_w18084_
	);
	LUT3 #(
		.INIT('h80)
	) name7572 (
		\wishbone_bd_ram_mem2_reg[53][23]/P0001 ,
		_w11933_,
		_w11979_,
		_w18085_
	);
	LUT4 #(
		.INIT('h0001)
	) name7573 (
		_w18082_,
		_w18083_,
		_w18084_,
		_w18085_,
		_w18086_
	);
	LUT3 #(
		.INIT('h80)
	) name7574 (
		\wishbone_bd_ram_mem2_reg[249][23]/P0001 ,
		_w11952_,
		_w11968_,
		_w18087_
	);
	LUT3 #(
		.INIT('h80)
	) name7575 (
		\wishbone_bd_ram_mem2_reg[179][23]/P0001 ,
		_w11938_,
		_w11942_,
		_w18088_
	);
	LUT3 #(
		.INIT('h80)
	) name7576 (
		\wishbone_bd_ram_mem2_reg[66][23]/P0001 ,
		_w11949_,
		_w11963_,
		_w18089_
	);
	LUT3 #(
		.INIT('h80)
	) name7577 (
		\wishbone_bd_ram_mem2_reg[180][23]/P0001 ,
		_w11929_,
		_w11942_,
		_w18090_
	);
	LUT4 #(
		.INIT('h0001)
	) name7578 (
		_w18087_,
		_w18088_,
		_w18089_,
		_w18090_,
		_w18091_
	);
	LUT3 #(
		.INIT('h80)
	) name7579 (
		\wishbone_bd_ram_mem2_reg[3][23]/P0001 ,
		_w11932_,
		_w11938_,
		_w18092_
	);
	LUT3 #(
		.INIT('h80)
	) name7580 (
		\wishbone_bd_ram_mem2_reg[194][23]/P0001 ,
		_w11945_,
		_w11963_,
		_w18093_
	);
	LUT3 #(
		.INIT('h80)
	) name7581 (
		\wishbone_bd_ram_mem2_reg[219][23]/P0001 ,
		_w11936_,
		_w11984_,
		_w18094_
	);
	LUT3 #(
		.INIT('h80)
	) name7582 (
		\wishbone_bd_ram_mem2_reg[79][23]/P0001 ,
		_w11949_,
		_w11973_,
		_w18095_
	);
	LUT4 #(
		.INIT('h0001)
	) name7583 (
		_w18092_,
		_w18093_,
		_w18094_,
		_w18095_,
		_w18096_
	);
	LUT3 #(
		.INIT('h80)
	) name7584 (
		\wishbone_bd_ram_mem2_reg[166][23]/P0001 ,
		_w11930_,
		_w11986_,
		_w18097_
	);
	LUT3 #(
		.INIT('h80)
	) name7585 (
		\wishbone_bd_ram_mem2_reg[126][23]/P0001 ,
		_w11948_,
		_w12012_,
		_w18098_
	);
	LUT3 #(
		.INIT('h80)
	) name7586 (
		\wishbone_bd_ram_mem2_reg[153][23]/P0001 ,
		_w11959_,
		_w11968_,
		_w18099_
	);
	LUT3 #(
		.INIT('h80)
	) name7587 (
		\wishbone_bd_ram_mem2_reg[201][23]/P0001 ,
		_w11945_,
		_w11968_,
		_w18100_
	);
	LUT4 #(
		.INIT('h0001)
	) name7588 (
		_w18097_,
		_w18098_,
		_w18099_,
		_w18100_,
		_w18101_
	);
	LUT4 #(
		.INIT('h8000)
	) name7589 (
		_w18086_,
		_w18091_,
		_w18096_,
		_w18101_,
		_w18102_
	);
	LUT3 #(
		.INIT('h80)
	) name7590 (
		\wishbone_bd_ram_mem2_reg[209][23]/P0001 ,
		_w11977_,
		_w11984_,
		_w18103_
	);
	LUT3 #(
		.INIT('h80)
	) name7591 (
		\wishbone_bd_ram_mem2_reg[196][23]/P0001 ,
		_w11929_,
		_w11945_,
		_w18104_
	);
	LUT3 #(
		.INIT('h80)
	) name7592 (
		\wishbone_bd_ram_mem2_reg[10][23]/P0001 ,
		_w11932_,
		_w11944_,
		_w18105_
	);
	LUT3 #(
		.INIT('h80)
	) name7593 (
		\wishbone_bd_ram_mem2_reg[24][23]/P0001 ,
		_w11935_,
		_w11990_,
		_w18106_
	);
	LUT4 #(
		.INIT('h0001)
	) name7594 (
		_w18103_,
		_w18104_,
		_w18105_,
		_w18106_,
		_w18107_
	);
	LUT3 #(
		.INIT('h80)
	) name7595 (
		\wishbone_bd_ram_mem2_reg[175][23]/P0001 ,
		_w11930_,
		_w11973_,
		_w18108_
	);
	LUT3 #(
		.INIT('h80)
	) name7596 (
		\wishbone_bd_ram_mem2_reg[64][23]/P0001 ,
		_w11941_,
		_w11949_,
		_w18109_
	);
	LUT3 #(
		.INIT('h80)
	) name7597 (
		\wishbone_bd_ram_mem2_reg[239][23]/P0001 ,
		_w11973_,
		_w11982_,
		_w18110_
	);
	LUT3 #(
		.INIT('h80)
	) name7598 (
		\wishbone_bd_ram_mem2_reg[118][23]/P0001 ,
		_w11986_,
		_w12012_,
		_w18111_
	);
	LUT4 #(
		.INIT('h0001)
	) name7599 (
		_w18108_,
		_w18109_,
		_w18110_,
		_w18111_,
		_w18112_
	);
	LUT3 #(
		.INIT('h80)
	) name7600 (
		\wishbone_bd_ram_mem2_reg[78][23]/P0001 ,
		_w11948_,
		_w11949_,
		_w18113_
	);
	LUT3 #(
		.INIT('h80)
	) name7601 (
		\wishbone_bd_ram_mem2_reg[207][23]/P0001 ,
		_w11945_,
		_w11973_,
		_w18114_
	);
	LUT3 #(
		.INIT('h80)
	) name7602 (
		\wishbone_bd_ram_mem2_reg[117][23]/P0001 ,
		_w11933_,
		_w12012_,
		_w18115_
	);
	LUT3 #(
		.INIT('h80)
	) name7603 (
		\wishbone_bd_ram_mem2_reg[237][23]/P0001 ,
		_w11966_,
		_w11982_,
		_w18116_
	);
	LUT4 #(
		.INIT('h0001)
	) name7604 (
		_w18113_,
		_w18114_,
		_w18115_,
		_w18116_,
		_w18117_
	);
	LUT3 #(
		.INIT('h80)
	) name7605 (
		\wishbone_bd_ram_mem2_reg[241][23]/P0001 ,
		_w11952_,
		_w11977_,
		_w18118_
	);
	LUT3 #(
		.INIT('h80)
	) name7606 (
		\wishbone_bd_ram_mem2_reg[227][23]/P0001 ,
		_w11938_,
		_w11982_,
		_w18119_
	);
	LUT3 #(
		.INIT('h80)
	) name7607 (
		\wishbone_bd_ram_mem2_reg[9][23]/P0001 ,
		_w11932_,
		_w11968_,
		_w18120_
	);
	LUT3 #(
		.INIT('h80)
	) name7608 (
		\wishbone_bd_ram_mem2_reg[206][23]/P0001 ,
		_w11945_,
		_w11948_,
		_w18121_
	);
	LUT4 #(
		.INIT('h0001)
	) name7609 (
		_w18118_,
		_w18119_,
		_w18120_,
		_w18121_,
		_w18122_
	);
	LUT4 #(
		.INIT('h8000)
	) name7610 (
		_w18107_,
		_w18112_,
		_w18117_,
		_w18122_,
		_w18123_
	);
	LUT3 #(
		.INIT('h80)
	) name7611 (
		\wishbone_bd_ram_mem2_reg[92][23]/P0001 ,
		_w11954_,
		_w11972_,
		_w18124_
	);
	LUT3 #(
		.INIT('h80)
	) name7612 (
		\wishbone_bd_ram_mem2_reg[230][23]/P0001 ,
		_w11982_,
		_w11986_,
		_w18125_
	);
	LUT3 #(
		.INIT('h80)
	) name7613 (
		\wishbone_bd_ram_mem2_reg[182][23]/P0001 ,
		_w11942_,
		_w11986_,
		_w18126_
	);
	LUT3 #(
		.INIT('h80)
	) name7614 (
		\wishbone_bd_ram_mem2_reg[80][23]/P0001 ,
		_w11941_,
		_w11972_,
		_w18127_
	);
	LUT4 #(
		.INIT('h0001)
	) name7615 (
		_w18124_,
		_w18125_,
		_w18126_,
		_w18127_,
		_w18128_
	);
	LUT3 #(
		.INIT('h80)
	) name7616 (
		\wishbone_bd_ram_mem2_reg[213][23]/P0001 ,
		_w11933_,
		_w11984_,
		_w18129_
	);
	LUT3 #(
		.INIT('h80)
	) name7617 (
		\wishbone_bd_ram_mem2_reg[212][23]/P0001 ,
		_w11929_,
		_w11984_,
		_w18130_
	);
	LUT3 #(
		.INIT('h80)
	) name7618 (
		\wishbone_bd_ram_mem2_reg[47][23]/P0001 ,
		_w11957_,
		_w11973_,
		_w18131_
	);
	LUT3 #(
		.INIT('h80)
	) name7619 (
		\wishbone_bd_ram_mem2_reg[1][23]/P0001 ,
		_w11932_,
		_w11977_,
		_w18132_
	);
	LUT4 #(
		.INIT('h0001)
	) name7620 (
		_w18129_,
		_w18130_,
		_w18131_,
		_w18132_,
		_w18133_
	);
	LUT3 #(
		.INIT('h80)
	) name7621 (
		\wishbone_bd_ram_mem2_reg[123][23]/P0001 ,
		_w11936_,
		_w12012_,
		_w18134_
	);
	LUT3 #(
		.INIT('h80)
	) name7622 (
		\wishbone_bd_ram_mem2_reg[149][23]/P0001 ,
		_w11933_,
		_w11959_,
		_w18135_
	);
	LUT3 #(
		.INIT('h80)
	) name7623 (
		\wishbone_bd_ram_mem2_reg[7][23]/P0001 ,
		_w11932_,
		_w11975_,
		_w18136_
	);
	LUT3 #(
		.INIT('h80)
	) name7624 (
		\wishbone_bd_ram_mem2_reg[203][23]/P0001 ,
		_w11936_,
		_w11945_,
		_w18137_
	);
	LUT4 #(
		.INIT('h0001)
	) name7625 (
		_w18134_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18138_
	);
	LUT3 #(
		.INIT('h80)
	) name7626 (
		\wishbone_bd_ram_mem2_reg[97][23]/P0001 ,
		_w11965_,
		_w11977_,
		_w18139_
	);
	LUT3 #(
		.INIT('h80)
	) name7627 (
		\wishbone_bd_ram_mem2_reg[138][23]/P0001 ,
		_w11944_,
		_w11955_,
		_w18140_
	);
	LUT3 #(
		.INIT('h80)
	) name7628 (
		\wishbone_bd_ram_mem2_reg[8][23]/P0001 ,
		_w11932_,
		_w11990_,
		_w18141_
	);
	LUT3 #(
		.INIT('h80)
	) name7629 (
		\wishbone_bd_ram_mem2_reg[62][23]/P0001 ,
		_w11948_,
		_w11979_,
		_w18142_
	);
	LUT4 #(
		.INIT('h0001)
	) name7630 (
		_w18139_,
		_w18140_,
		_w18141_,
		_w18142_,
		_w18143_
	);
	LUT4 #(
		.INIT('h8000)
	) name7631 (
		_w18128_,
		_w18133_,
		_w18138_,
		_w18143_,
		_w18144_
	);
	LUT4 #(
		.INIT('h8000)
	) name7632 (
		_w18081_,
		_w18102_,
		_w18123_,
		_w18144_,
		_w18145_
	);
	LUT3 #(
		.INIT('h80)
	) name7633 (
		\wishbone_bd_ram_mem2_reg[157][23]/P0001 ,
		_w11959_,
		_w11966_,
		_w18146_
	);
	LUT3 #(
		.INIT('h80)
	) name7634 (
		\wishbone_bd_ram_mem2_reg[105][23]/P0001 ,
		_w11965_,
		_w11968_,
		_w18147_
	);
	LUT3 #(
		.INIT('h80)
	) name7635 (
		\wishbone_bd_ram_mem2_reg[220][23]/P0001 ,
		_w11954_,
		_w11984_,
		_w18148_
	);
	LUT3 #(
		.INIT('h80)
	) name7636 (
		\wishbone_bd_ram_mem2_reg[125][23]/P0001 ,
		_w11966_,
		_w12012_,
		_w18149_
	);
	LUT4 #(
		.INIT('h0001)
	) name7637 (
		_w18146_,
		_w18147_,
		_w18148_,
		_w18149_,
		_w18150_
	);
	LUT3 #(
		.INIT('h80)
	) name7638 (
		\wishbone_bd_ram_mem2_reg[243][23]/P0001 ,
		_w11938_,
		_w11952_,
		_w18151_
	);
	LUT3 #(
		.INIT('h80)
	) name7639 (
		\wishbone_bd_ram_mem2_reg[70][23]/P0001 ,
		_w11949_,
		_w11986_,
		_w18152_
	);
	LUT3 #(
		.INIT('h80)
	) name7640 (
		\wishbone_bd_ram_mem2_reg[161][23]/P0001 ,
		_w11930_,
		_w11977_,
		_w18153_
	);
	LUT3 #(
		.INIT('h80)
	) name7641 (
		\wishbone_bd_ram_mem2_reg[29][23]/P0001 ,
		_w11935_,
		_w11966_,
		_w18154_
	);
	LUT4 #(
		.INIT('h0001)
	) name7642 (
		_w18151_,
		_w18152_,
		_w18153_,
		_w18154_,
		_w18155_
	);
	LUT3 #(
		.INIT('h80)
	) name7643 (
		\wishbone_bd_ram_mem2_reg[82][23]/P0001 ,
		_w11963_,
		_w11972_,
		_w18156_
	);
	LUT3 #(
		.INIT('h80)
	) name7644 (
		\wishbone_bd_ram_mem2_reg[55][23]/P0001 ,
		_w11975_,
		_w11979_,
		_w18157_
	);
	LUT3 #(
		.INIT('h80)
	) name7645 (
		\wishbone_bd_ram_mem2_reg[81][23]/P0001 ,
		_w11972_,
		_w11977_,
		_w18158_
	);
	LUT3 #(
		.INIT('h80)
	) name7646 (
		\wishbone_bd_ram_mem2_reg[223][23]/P0001 ,
		_w11973_,
		_w11984_,
		_w18159_
	);
	LUT4 #(
		.INIT('h0001)
	) name7647 (
		_w18156_,
		_w18157_,
		_w18158_,
		_w18159_,
		_w18160_
	);
	LUT3 #(
		.INIT('h80)
	) name7648 (
		\wishbone_bd_ram_mem2_reg[111][23]/P0001 ,
		_w11965_,
		_w11973_,
		_w18161_
	);
	LUT3 #(
		.INIT('h80)
	) name7649 (
		\wishbone_bd_ram_mem2_reg[160][23]/P0001 ,
		_w11930_,
		_w11941_,
		_w18162_
	);
	LUT3 #(
		.INIT('h80)
	) name7650 (
		\wishbone_bd_ram_mem2_reg[192][23]/P0001 ,
		_w11941_,
		_w11945_,
		_w18163_
	);
	LUT3 #(
		.INIT('h80)
	) name7651 (
		\wishbone_bd_ram_mem2_reg[159][23]/P0001 ,
		_w11959_,
		_w11973_,
		_w18164_
	);
	LUT4 #(
		.INIT('h0001)
	) name7652 (
		_w18161_,
		_w18162_,
		_w18163_,
		_w18164_,
		_w18165_
	);
	LUT4 #(
		.INIT('h8000)
	) name7653 (
		_w18150_,
		_w18155_,
		_w18160_,
		_w18165_,
		_w18166_
	);
	LUT3 #(
		.INIT('h80)
	) name7654 (
		\wishbone_bd_ram_mem2_reg[189][23]/P0001 ,
		_w11942_,
		_w11966_,
		_w18167_
	);
	LUT3 #(
		.INIT('h80)
	) name7655 (
		\wishbone_bd_ram_mem2_reg[197][23]/P0001 ,
		_w11933_,
		_w11945_,
		_w18168_
	);
	LUT3 #(
		.INIT('h80)
	) name7656 (
		\wishbone_bd_ram_mem2_reg[72][23]/P0001 ,
		_w11949_,
		_w11990_,
		_w18169_
	);
	LUT3 #(
		.INIT('h80)
	) name7657 (
		\wishbone_bd_ram_mem2_reg[6][23]/P0001 ,
		_w11932_,
		_w11986_,
		_w18170_
	);
	LUT4 #(
		.INIT('h0001)
	) name7658 (
		_w18167_,
		_w18168_,
		_w18169_,
		_w18170_,
		_w18171_
	);
	LUT3 #(
		.INIT('h80)
	) name7659 (
		\wishbone_bd_ram_mem2_reg[43][23]/P0001 ,
		_w11936_,
		_w11957_,
		_w18172_
	);
	LUT3 #(
		.INIT('h80)
	) name7660 (
		\wishbone_bd_ram_mem2_reg[18][23]/P0001 ,
		_w11935_,
		_w11963_,
		_w18173_
	);
	LUT3 #(
		.INIT('h80)
	) name7661 (
		\wishbone_bd_ram_mem2_reg[236][23]/P0001 ,
		_w11954_,
		_w11982_,
		_w18174_
	);
	LUT3 #(
		.INIT('h80)
	) name7662 (
		\wishbone_bd_ram_mem2_reg[102][23]/P0001 ,
		_w11965_,
		_w11986_,
		_w18175_
	);
	LUT4 #(
		.INIT('h0001)
	) name7663 (
		_w18172_,
		_w18173_,
		_w18174_,
		_w18175_,
		_w18176_
	);
	LUT3 #(
		.INIT('h80)
	) name7664 (
		\wishbone_bd_ram_mem2_reg[235][23]/P0001 ,
		_w11936_,
		_w11982_,
		_w18177_
	);
	LUT3 #(
		.INIT('h80)
	) name7665 (
		\wishbone_bd_ram_mem2_reg[112][23]/P0001 ,
		_w11941_,
		_w12012_,
		_w18178_
	);
	LUT3 #(
		.INIT('h80)
	) name7666 (
		\wishbone_bd_ram_mem2_reg[34][23]/P0001 ,
		_w11957_,
		_w11963_,
		_w18179_
	);
	LUT3 #(
		.INIT('h80)
	) name7667 (
		\wishbone_bd_ram_mem2_reg[251][23]/P0001 ,
		_w11936_,
		_w11952_,
		_w18180_
	);
	LUT4 #(
		.INIT('h0001)
	) name7668 (
		_w18177_,
		_w18178_,
		_w18179_,
		_w18180_,
		_w18181_
	);
	LUT3 #(
		.INIT('h80)
	) name7669 (
		\wishbone_bd_ram_mem2_reg[141][23]/P0001 ,
		_w11955_,
		_w11966_,
		_w18182_
	);
	LUT3 #(
		.INIT('h80)
	) name7670 (
		\wishbone_bd_ram_mem2_reg[238][23]/P0001 ,
		_w11948_,
		_w11982_,
		_w18183_
	);
	LUT3 #(
		.INIT('h80)
	) name7671 (
		\wishbone_bd_ram_mem2_reg[114][23]/P0001 ,
		_w11963_,
		_w12012_,
		_w18184_
	);
	LUT3 #(
		.INIT('h80)
	) name7672 (
		\wishbone_bd_ram_mem2_reg[75][23]/P0001 ,
		_w11936_,
		_w11949_,
		_w18185_
	);
	LUT4 #(
		.INIT('h0001)
	) name7673 (
		_w18182_,
		_w18183_,
		_w18184_,
		_w18185_,
		_w18186_
	);
	LUT4 #(
		.INIT('h8000)
	) name7674 (
		_w18171_,
		_w18176_,
		_w18181_,
		_w18186_,
		_w18187_
	);
	LUT3 #(
		.INIT('h80)
	) name7675 (
		\wishbone_bd_ram_mem2_reg[109][23]/P0001 ,
		_w11965_,
		_w11966_,
		_w18188_
	);
	LUT3 #(
		.INIT('h80)
	) name7676 (
		\wishbone_bd_ram_mem2_reg[142][23]/P0001 ,
		_w11948_,
		_w11955_,
		_w18189_
	);
	LUT3 #(
		.INIT('h80)
	) name7677 (
		\wishbone_bd_ram_mem2_reg[104][23]/P0001 ,
		_w11965_,
		_w11990_,
		_w18190_
	);
	LUT3 #(
		.INIT('h80)
	) name7678 (
		\wishbone_bd_ram_mem2_reg[151][23]/P0001 ,
		_w11959_,
		_w11975_,
		_w18191_
	);
	LUT4 #(
		.INIT('h0001)
	) name7679 (
		_w18188_,
		_w18189_,
		_w18190_,
		_w18191_,
		_w18192_
	);
	LUT3 #(
		.INIT('h80)
	) name7680 (
		\wishbone_bd_ram_mem2_reg[211][23]/P0001 ,
		_w11938_,
		_w11984_,
		_w18193_
	);
	LUT3 #(
		.INIT('h80)
	) name7681 (
		\wishbone_bd_ram_mem2_reg[240][23]/P0001 ,
		_w11941_,
		_w11952_,
		_w18194_
	);
	LUT3 #(
		.INIT('h80)
	) name7682 (
		\wishbone_bd_ram_mem2_reg[255][23]/P0001 ,
		_w11952_,
		_w11973_,
		_w18195_
	);
	LUT3 #(
		.INIT('h80)
	) name7683 (
		\wishbone_bd_ram_mem2_reg[135][23]/P0001 ,
		_w11955_,
		_w11975_,
		_w18196_
	);
	LUT4 #(
		.INIT('h0001)
	) name7684 (
		_w18193_,
		_w18194_,
		_w18195_,
		_w18196_,
		_w18197_
	);
	LUT3 #(
		.INIT('h80)
	) name7685 (
		\wishbone_bd_ram_mem2_reg[181][23]/P0001 ,
		_w11933_,
		_w11942_,
		_w18198_
	);
	LUT3 #(
		.INIT('h80)
	) name7686 (
		\wishbone_bd_ram_mem2_reg[144][23]/P0001 ,
		_w11941_,
		_w11959_,
		_w18199_
	);
	LUT3 #(
		.INIT('h80)
	) name7687 (
		\wishbone_bd_ram_mem2_reg[134][23]/P0001 ,
		_w11955_,
		_w11986_,
		_w18200_
	);
	LUT3 #(
		.INIT('h80)
	) name7688 (
		\wishbone_bd_ram_mem2_reg[107][23]/P0001 ,
		_w11936_,
		_w11965_,
		_w18201_
	);
	LUT4 #(
		.INIT('h0001)
	) name7689 (
		_w18198_,
		_w18199_,
		_w18200_,
		_w18201_,
		_w18202_
	);
	LUT3 #(
		.INIT('h80)
	) name7690 (
		\wishbone_bd_ram_mem2_reg[164][23]/P0001 ,
		_w11929_,
		_w11930_,
		_w18203_
	);
	LUT3 #(
		.INIT('h80)
	) name7691 (
		\wishbone_bd_ram_mem2_reg[133][23]/P0001 ,
		_w11933_,
		_w11955_,
		_w18204_
	);
	LUT3 #(
		.INIT('h80)
	) name7692 (
		\wishbone_bd_ram_mem2_reg[163][23]/P0001 ,
		_w11930_,
		_w11938_,
		_w18205_
	);
	LUT3 #(
		.INIT('h80)
	) name7693 (
		\wishbone_bd_ram_mem2_reg[136][23]/P0001 ,
		_w11955_,
		_w11990_,
		_w18206_
	);
	LUT4 #(
		.INIT('h0001)
	) name7694 (
		_w18203_,
		_w18204_,
		_w18205_,
		_w18206_,
		_w18207_
	);
	LUT4 #(
		.INIT('h8000)
	) name7695 (
		_w18192_,
		_w18197_,
		_w18202_,
		_w18207_,
		_w18208_
	);
	LUT3 #(
		.INIT('h80)
	) name7696 (
		\wishbone_bd_ram_mem2_reg[56][23]/P0001 ,
		_w11979_,
		_w11990_,
		_w18209_
	);
	LUT3 #(
		.INIT('h80)
	) name7697 (
		\wishbone_bd_ram_mem2_reg[59][23]/P0001 ,
		_w11936_,
		_w11979_,
		_w18210_
	);
	LUT3 #(
		.INIT('h80)
	) name7698 (
		\wishbone_bd_ram_mem2_reg[129][23]/P0001 ,
		_w11955_,
		_w11977_,
		_w18211_
	);
	LUT3 #(
		.INIT('h80)
	) name7699 (
		\wishbone_bd_ram_mem2_reg[245][23]/P0001 ,
		_w11933_,
		_w11952_,
		_w18212_
	);
	LUT4 #(
		.INIT('h0001)
	) name7700 (
		_w18209_,
		_w18210_,
		_w18211_,
		_w18212_,
		_w18213_
	);
	LUT3 #(
		.INIT('h80)
	) name7701 (
		\wishbone_bd_ram_mem2_reg[54][23]/P0001 ,
		_w11979_,
		_w11986_,
		_w18214_
	);
	LUT3 #(
		.INIT('h80)
	) name7702 (
		\wishbone_bd_ram_mem2_reg[234][23]/P0001 ,
		_w11944_,
		_w11982_,
		_w18215_
	);
	LUT3 #(
		.INIT('h80)
	) name7703 (
		\wishbone_bd_ram_mem2_reg[222][23]/P0001 ,
		_w11948_,
		_w11984_,
		_w18216_
	);
	LUT3 #(
		.INIT('h80)
	) name7704 (
		\wishbone_bd_ram_mem2_reg[73][23]/P0001 ,
		_w11949_,
		_w11968_,
		_w18217_
	);
	LUT4 #(
		.INIT('h0001)
	) name7705 (
		_w18214_,
		_w18215_,
		_w18216_,
		_w18217_,
		_w18218_
	);
	LUT3 #(
		.INIT('h80)
	) name7706 (
		\wishbone_bd_ram_mem2_reg[140][23]/P0001 ,
		_w11954_,
		_w11955_,
		_w18219_
	);
	LUT3 #(
		.INIT('h80)
	) name7707 (
		\wishbone_bd_ram_mem2_reg[87][23]/P0001 ,
		_w11972_,
		_w11975_,
		_w18220_
	);
	LUT3 #(
		.INIT('h80)
	) name7708 (
		\wishbone_bd_ram_mem2_reg[51][23]/P0001 ,
		_w11938_,
		_w11979_,
		_w18221_
	);
	LUT3 #(
		.INIT('h80)
	) name7709 (
		\wishbone_bd_ram_mem2_reg[250][23]/P0001 ,
		_w11944_,
		_w11952_,
		_w18222_
	);
	LUT4 #(
		.INIT('h0001)
	) name7710 (
		_w18219_,
		_w18220_,
		_w18221_,
		_w18222_,
		_w18223_
	);
	LUT3 #(
		.INIT('h80)
	) name7711 (
		\wishbone_bd_ram_mem2_reg[242][23]/P0001 ,
		_w11952_,
		_w11963_,
		_w18224_
	);
	LUT3 #(
		.INIT('h80)
	) name7712 (
		\wishbone_bd_ram_mem2_reg[214][23]/P0001 ,
		_w11984_,
		_w11986_,
		_w18225_
	);
	LUT3 #(
		.INIT('h80)
	) name7713 (
		\wishbone_bd_ram_mem2_reg[20][23]/P0001 ,
		_w11929_,
		_w11935_,
		_w18226_
	);
	LUT3 #(
		.INIT('h80)
	) name7714 (
		\wishbone_bd_ram_mem2_reg[65][23]/P0001 ,
		_w11949_,
		_w11977_,
		_w18227_
	);
	LUT4 #(
		.INIT('h0001)
	) name7715 (
		_w18224_,
		_w18225_,
		_w18226_,
		_w18227_,
		_w18228_
	);
	LUT4 #(
		.INIT('h8000)
	) name7716 (
		_w18213_,
		_w18218_,
		_w18223_,
		_w18228_,
		_w18229_
	);
	LUT4 #(
		.INIT('h8000)
	) name7717 (
		_w18166_,
		_w18187_,
		_w18208_,
		_w18229_,
		_w18230_
	);
	LUT3 #(
		.INIT('h80)
	) name7718 (
		\wishbone_bd_ram_mem2_reg[2][23]/P0001 ,
		_w11932_,
		_w11963_,
		_w18231_
	);
	LUT3 #(
		.INIT('h80)
	) name7719 (
		\wishbone_bd_ram_mem2_reg[42][23]/P0001 ,
		_w11944_,
		_w11957_,
		_w18232_
	);
	LUT3 #(
		.INIT('h80)
	) name7720 (
		\wishbone_bd_ram_mem2_reg[218][23]/P0001 ,
		_w11944_,
		_w11984_,
		_w18233_
	);
	LUT3 #(
		.INIT('h80)
	) name7721 (
		\wishbone_bd_ram_mem2_reg[158][23]/P0001 ,
		_w11948_,
		_w11959_,
		_w18234_
	);
	LUT4 #(
		.INIT('h0001)
	) name7722 (
		_w18231_,
		_w18232_,
		_w18233_,
		_w18234_,
		_w18235_
	);
	LUT3 #(
		.INIT('h80)
	) name7723 (
		\wishbone_bd_ram_mem2_reg[12][23]/P0001 ,
		_w11932_,
		_w11954_,
		_w18236_
	);
	LUT3 #(
		.INIT('h80)
	) name7724 (
		\wishbone_bd_ram_mem2_reg[30][23]/P0001 ,
		_w11935_,
		_w11948_,
		_w18237_
	);
	LUT3 #(
		.INIT('h80)
	) name7725 (
		\wishbone_bd_ram_mem2_reg[221][23]/P0001 ,
		_w11966_,
		_w11984_,
		_w18238_
	);
	LUT3 #(
		.INIT('h80)
	) name7726 (
		\wishbone_bd_ram_mem2_reg[188][23]/P0001 ,
		_w11942_,
		_w11954_,
		_w18239_
	);
	LUT4 #(
		.INIT('h0001)
	) name7727 (
		_w18236_,
		_w18237_,
		_w18238_,
		_w18239_,
		_w18240_
	);
	LUT3 #(
		.INIT('h80)
	) name7728 (
		\wishbone_bd_ram_mem2_reg[98][23]/P0001 ,
		_w11963_,
		_w11965_,
		_w18241_
	);
	LUT3 #(
		.INIT('h80)
	) name7729 (
		\wishbone_bd_ram_mem2_reg[27][23]/P0001 ,
		_w11935_,
		_w11936_,
		_w18242_
	);
	LUT3 #(
		.INIT('h80)
	) name7730 (
		\wishbone_bd_ram_mem2_reg[205][23]/P0001 ,
		_w11945_,
		_w11966_,
		_w18243_
	);
	LUT3 #(
		.INIT('h80)
	) name7731 (
		\wishbone_bd_ram_mem2_reg[71][23]/P0001 ,
		_w11949_,
		_w11975_,
		_w18244_
	);
	LUT4 #(
		.INIT('h0001)
	) name7732 (
		_w18241_,
		_w18242_,
		_w18243_,
		_w18244_,
		_w18245_
	);
	LUT3 #(
		.INIT('h80)
	) name7733 (
		\wishbone_bd_ram_mem2_reg[40][23]/P0001 ,
		_w11957_,
		_w11990_,
		_w18246_
	);
	LUT3 #(
		.INIT('h80)
	) name7734 (
		\wishbone_bd_ram_mem2_reg[21][23]/P0001 ,
		_w11933_,
		_w11935_,
		_w18247_
	);
	LUT3 #(
		.INIT('h80)
	) name7735 (
		\wishbone_bd_ram_mem2_reg[101][23]/P0001 ,
		_w11933_,
		_w11965_,
		_w18248_
	);
	LUT3 #(
		.INIT('h80)
	) name7736 (
		\wishbone_bd_ram_mem2_reg[147][23]/P0001 ,
		_w11938_,
		_w11959_,
		_w18249_
	);
	LUT4 #(
		.INIT('h0001)
	) name7737 (
		_w18246_,
		_w18247_,
		_w18248_,
		_w18249_,
		_w18250_
	);
	LUT4 #(
		.INIT('h8000)
	) name7738 (
		_w18235_,
		_w18240_,
		_w18245_,
		_w18250_,
		_w18251_
	);
	LUT3 #(
		.INIT('h80)
	) name7739 (
		\wishbone_bd_ram_mem2_reg[233][23]/P0001 ,
		_w11968_,
		_w11982_,
		_w18252_
	);
	LUT3 #(
		.INIT('h80)
	) name7740 (
		\wishbone_bd_ram_mem2_reg[37][23]/P0001 ,
		_w11933_,
		_w11957_,
		_w18253_
	);
	LUT3 #(
		.INIT('h80)
	) name7741 (
		\wishbone_bd_ram_mem2_reg[177][23]/P0001 ,
		_w11942_,
		_w11977_,
		_w18254_
	);
	LUT3 #(
		.INIT('h80)
	) name7742 (
		\wishbone_bd_ram_mem2_reg[174][23]/P0001 ,
		_w11930_,
		_w11948_,
		_w18255_
	);
	LUT4 #(
		.INIT('h0001)
	) name7743 (
		_w18252_,
		_w18253_,
		_w18254_,
		_w18255_,
		_w18256_
	);
	LUT3 #(
		.INIT('h80)
	) name7744 (
		\wishbone_bd_ram_mem2_reg[94][23]/P0001 ,
		_w11948_,
		_w11972_,
		_w18257_
	);
	LUT3 #(
		.INIT('h80)
	) name7745 (
		\wishbone_bd_ram_mem2_reg[176][23]/P0001 ,
		_w11941_,
		_w11942_,
		_w18258_
	);
	LUT3 #(
		.INIT('h80)
	) name7746 (
		\wishbone_bd_ram_mem2_reg[172][23]/P0001 ,
		_w11930_,
		_w11954_,
		_w18259_
	);
	LUT3 #(
		.INIT('h80)
	) name7747 (
		\wishbone_bd_ram_mem2_reg[193][23]/P0001 ,
		_w11945_,
		_w11977_,
		_w18260_
	);
	LUT4 #(
		.INIT('h0001)
	) name7748 (
		_w18257_,
		_w18258_,
		_w18259_,
		_w18260_,
		_w18261_
	);
	LUT3 #(
		.INIT('h80)
	) name7749 (
		\wishbone_bd_ram_mem2_reg[67][23]/P0001 ,
		_w11938_,
		_w11949_,
		_w18262_
	);
	LUT3 #(
		.INIT('h80)
	) name7750 (
		\wishbone_bd_ram_mem2_reg[121][23]/P0001 ,
		_w11968_,
		_w12012_,
		_w18263_
	);
	LUT3 #(
		.INIT('h80)
	) name7751 (
		\wishbone_bd_ram_mem2_reg[48][23]/P0001 ,
		_w11941_,
		_w11979_,
		_w18264_
	);
	LUT3 #(
		.INIT('h80)
	) name7752 (
		\wishbone_bd_ram_mem2_reg[169][23]/P0001 ,
		_w11930_,
		_w11968_,
		_w18265_
	);
	LUT4 #(
		.INIT('h0001)
	) name7753 (
		_w18262_,
		_w18263_,
		_w18264_,
		_w18265_,
		_w18266_
	);
	LUT3 #(
		.INIT('h80)
	) name7754 (
		\wishbone_bd_ram_mem2_reg[99][23]/P0001 ,
		_w11938_,
		_w11965_,
		_w18267_
	);
	LUT3 #(
		.INIT('h80)
	) name7755 (
		\wishbone_bd_ram_mem2_reg[186][23]/P0001 ,
		_w11942_,
		_w11944_,
		_w18268_
	);
	LUT3 #(
		.INIT('h80)
	) name7756 (
		\wishbone_bd_ram_mem2_reg[195][23]/P0001 ,
		_w11938_,
		_w11945_,
		_w18269_
	);
	LUT3 #(
		.INIT('h80)
	) name7757 (
		\wishbone_bd_ram_mem2_reg[76][23]/P0001 ,
		_w11949_,
		_w11954_,
		_w18270_
	);
	LUT4 #(
		.INIT('h0001)
	) name7758 (
		_w18267_,
		_w18268_,
		_w18269_,
		_w18270_,
		_w18271_
	);
	LUT4 #(
		.INIT('h8000)
	) name7759 (
		_w18256_,
		_w18261_,
		_w18266_,
		_w18271_,
		_w18272_
	);
	LUT3 #(
		.INIT('h80)
	) name7760 (
		\wishbone_bd_ram_mem2_reg[217][23]/P0001 ,
		_w11968_,
		_w11984_,
		_w18273_
	);
	LUT3 #(
		.INIT('h80)
	) name7761 (
		\wishbone_bd_ram_mem2_reg[162][23]/P0001 ,
		_w11930_,
		_w11963_,
		_w18274_
	);
	LUT3 #(
		.INIT('h80)
	) name7762 (
		\wishbone_bd_ram_mem2_reg[4][23]/P0001 ,
		_w11929_,
		_w11932_,
		_w18275_
	);
	LUT3 #(
		.INIT('h80)
	) name7763 (
		\wishbone_bd_ram_mem2_reg[106][23]/P0001 ,
		_w11944_,
		_w11965_,
		_w18276_
	);
	LUT4 #(
		.INIT('h0001)
	) name7764 (
		_w18273_,
		_w18274_,
		_w18275_,
		_w18276_,
		_w18277_
	);
	LUT3 #(
		.INIT('h80)
	) name7765 (
		\wishbone_bd_ram_mem2_reg[246][23]/P0001 ,
		_w11952_,
		_w11986_,
		_w18278_
	);
	LUT3 #(
		.INIT('h80)
	) name7766 (
		\wishbone_bd_ram_mem2_reg[156][23]/P0001 ,
		_w11954_,
		_w11959_,
		_w18279_
	);
	LUT3 #(
		.INIT('h80)
	) name7767 (
		\wishbone_bd_ram_mem2_reg[74][23]/P0001 ,
		_w11944_,
		_w11949_,
		_w18280_
	);
	LUT3 #(
		.INIT('h80)
	) name7768 (
		\wishbone_bd_ram_mem2_reg[91][23]/P0001 ,
		_w11936_,
		_w11972_,
		_w18281_
	);
	LUT4 #(
		.INIT('h0001)
	) name7769 (
		_w18278_,
		_w18279_,
		_w18280_,
		_w18281_,
		_w18282_
	);
	LUT3 #(
		.INIT('h80)
	) name7770 (
		\wishbone_bd_ram_mem2_reg[95][23]/P0001 ,
		_w11972_,
		_w11973_,
		_w18283_
	);
	LUT3 #(
		.INIT('h80)
	) name7771 (
		\wishbone_bd_ram_mem2_reg[232][23]/P0001 ,
		_w11982_,
		_w11990_,
		_w18284_
	);
	LUT3 #(
		.INIT('h80)
	) name7772 (
		\wishbone_bd_ram_mem2_reg[13][23]/P0001 ,
		_w11932_,
		_w11966_,
		_w18285_
	);
	LUT3 #(
		.INIT('h80)
	) name7773 (
		\wishbone_bd_ram_mem2_reg[173][23]/P0001 ,
		_w11930_,
		_w11966_,
		_w18286_
	);
	LUT4 #(
		.INIT('h0001)
	) name7774 (
		_w18283_,
		_w18284_,
		_w18285_,
		_w18286_,
		_w18287_
	);
	LUT3 #(
		.INIT('h80)
	) name7775 (
		\wishbone_bd_ram_mem2_reg[26][23]/P0001 ,
		_w11935_,
		_w11944_,
		_w18288_
	);
	LUT3 #(
		.INIT('h80)
	) name7776 (
		\wishbone_bd_ram_mem2_reg[150][23]/P0001 ,
		_w11959_,
		_w11986_,
		_w18289_
	);
	LUT3 #(
		.INIT('h80)
	) name7777 (
		\wishbone_bd_ram_mem2_reg[22][23]/P0001 ,
		_w11935_,
		_w11986_,
		_w18290_
	);
	LUT3 #(
		.INIT('h80)
	) name7778 (
		\wishbone_bd_ram_mem2_reg[168][23]/P0001 ,
		_w11930_,
		_w11990_,
		_w18291_
	);
	LUT4 #(
		.INIT('h0001)
	) name7779 (
		_w18288_,
		_w18289_,
		_w18290_,
		_w18291_,
		_w18292_
	);
	LUT4 #(
		.INIT('h8000)
	) name7780 (
		_w18277_,
		_w18282_,
		_w18287_,
		_w18292_,
		_w18293_
	);
	LUT3 #(
		.INIT('h80)
	) name7781 (
		\wishbone_bd_ram_mem2_reg[127][23]/P0001 ,
		_w11973_,
		_w12012_,
		_w18294_
	);
	LUT3 #(
		.INIT('h80)
	) name7782 (
		\wishbone_bd_ram_mem2_reg[224][23]/P0001 ,
		_w11941_,
		_w11982_,
		_w18295_
	);
	LUT3 #(
		.INIT('h80)
	) name7783 (
		\wishbone_bd_ram_mem2_reg[229][23]/P0001 ,
		_w11933_,
		_w11982_,
		_w18296_
	);
	LUT3 #(
		.INIT('h80)
	) name7784 (
		\wishbone_bd_ram_mem2_reg[225][23]/P0001 ,
		_w11977_,
		_w11982_,
		_w18297_
	);
	LUT4 #(
		.INIT('h0001)
	) name7785 (
		_w18294_,
		_w18295_,
		_w18296_,
		_w18297_,
		_w18298_
	);
	LUT3 #(
		.INIT('h80)
	) name7786 (
		\wishbone_bd_ram_mem2_reg[58][23]/P0001 ,
		_w11944_,
		_w11979_,
		_w18299_
	);
	LUT3 #(
		.INIT('h80)
	) name7787 (
		\wishbone_bd_ram_mem2_reg[200][23]/P0001 ,
		_w11945_,
		_w11990_,
		_w18300_
	);
	LUT3 #(
		.INIT('h80)
	) name7788 (
		\wishbone_bd_ram_mem2_reg[254][23]/P0001 ,
		_w11948_,
		_w11952_,
		_w18301_
	);
	LUT3 #(
		.INIT('h80)
	) name7789 (
		\wishbone_bd_ram_mem2_reg[204][23]/P0001 ,
		_w11945_,
		_w11954_,
		_w18302_
	);
	LUT4 #(
		.INIT('h0001)
	) name7790 (
		_w18299_,
		_w18300_,
		_w18301_,
		_w18302_,
		_w18303_
	);
	LUT3 #(
		.INIT('h80)
	) name7791 (
		\wishbone_bd_ram_mem2_reg[252][23]/P0001 ,
		_w11952_,
		_w11954_,
		_w18304_
	);
	LUT3 #(
		.INIT('h80)
	) name7792 (
		\wishbone_bd_ram_mem2_reg[77][23]/P0001 ,
		_w11949_,
		_w11966_,
		_w18305_
	);
	LUT3 #(
		.INIT('h80)
	) name7793 (
		\wishbone_bd_ram_mem2_reg[116][23]/P0001 ,
		_w11929_,
		_w12012_,
		_w18306_
	);
	LUT3 #(
		.INIT('h80)
	) name7794 (
		\wishbone_bd_ram_mem2_reg[23][23]/P0001 ,
		_w11935_,
		_w11975_,
		_w18307_
	);
	LUT4 #(
		.INIT('h0001)
	) name7795 (
		_w18304_,
		_w18305_,
		_w18306_,
		_w18307_,
		_w18308_
	);
	LUT3 #(
		.INIT('h80)
	) name7796 (
		\wishbone_bd_ram_mem2_reg[83][23]/P0001 ,
		_w11938_,
		_w11972_,
		_w18309_
	);
	LUT3 #(
		.INIT('h80)
	) name7797 (
		\wishbone_bd_ram_mem2_reg[69][23]/P0001 ,
		_w11933_,
		_w11949_,
		_w18310_
	);
	LUT3 #(
		.INIT('h80)
	) name7798 (
		\wishbone_bd_ram_mem2_reg[119][23]/P0001 ,
		_w11975_,
		_w12012_,
		_w18311_
	);
	LUT3 #(
		.INIT('h80)
	) name7799 (
		\wishbone_bd_ram_mem2_reg[146][23]/P0001 ,
		_w11959_,
		_w11963_,
		_w18312_
	);
	LUT4 #(
		.INIT('h0001)
	) name7800 (
		_w18309_,
		_w18310_,
		_w18311_,
		_w18312_,
		_w18313_
	);
	LUT4 #(
		.INIT('h8000)
	) name7801 (
		_w18298_,
		_w18303_,
		_w18308_,
		_w18313_,
		_w18314_
	);
	LUT4 #(
		.INIT('h8000)
	) name7802 (
		_w18251_,
		_w18272_,
		_w18293_,
		_w18314_,
		_w18315_
	);
	LUT3 #(
		.INIT('h80)
	) name7803 (
		\wishbone_bd_ram_mem2_reg[0][23]/P0001 ,
		_w11932_,
		_w11941_,
		_w18316_
	);
	LUT3 #(
		.INIT('h80)
	) name7804 (
		\wishbone_bd_ram_mem2_reg[122][23]/P0001 ,
		_w11944_,
		_w12012_,
		_w18317_
	);
	LUT3 #(
		.INIT('h80)
	) name7805 (
		\wishbone_bd_ram_mem2_reg[46][23]/P0001 ,
		_w11948_,
		_w11957_,
		_w18318_
	);
	LUT3 #(
		.INIT('h80)
	) name7806 (
		\wishbone_bd_ram_mem2_reg[155][23]/P0001 ,
		_w11936_,
		_w11959_,
		_w18319_
	);
	LUT4 #(
		.INIT('h0001)
	) name7807 (
		_w18316_,
		_w18317_,
		_w18318_,
		_w18319_,
		_w18320_
	);
	LUT3 #(
		.INIT('h80)
	) name7808 (
		\wishbone_bd_ram_mem2_reg[57][23]/P0001 ,
		_w11968_,
		_w11979_,
		_w18321_
	);
	LUT3 #(
		.INIT('h80)
	) name7809 (
		\wishbone_bd_ram_mem2_reg[28][23]/P0001 ,
		_w11935_,
		_w11954_,
		_w18322_
	);
	LUT3 #(
		.INIT('h80)
	) name7810 (
		\wishbone_bd_ram_mem2_reg[148][23]/P0001 ,
		_w11929_,
		_w11959_,
		_w18323_
	);
	LUT3 #(
		.INIT('h80)
	) name7811 (
		\wishbone_bd_ram_mem2_reg[190][23]/P0001 ,
		_w11942_,
		_w11948_,
		_w18324_
	);
	LUT4 #(
		.INIT('h0001)
	) name7812 (
		_w18321_,
		_w18322_,
		_w18323_,
		_w18324_,
		_w18325_
	);
	LUT3 #(
		.INIT('h80)
	) name7813 (
		\wishbone_bd_ram_mem2_reg[63][23]/P0001 ,
		_w11973_,
		_w11979_,
		_w18326_
	);
	LUT3 #(
		.INIT('h80)
	) name7814 (
		\wishbone_bd_ram_mem2_reg[253][23]/P0001 ,
		_w11952_,
		_w11966_,
		_w18327_
	);
	LUT3 #(
		.INIT('h80)
	) name7815 (
		\wishbone_bd_ram_mem2_reg[36][23]/P0001 ,
		_w11929_,
		_w11957_,
		_w18328_
	);
	LUT3 #(
		.INIT('h80)
	) name7816 (
		\wishbone_bd_ram_mem2_reg[113][23]/P0001 ,
		_w11977_,
		_w12012_,
		_w18329_
	);
	LUT4 #(
		.INIT('h0001)
	) name7817 (
		_w18326_,
		_w18327_,
		_w18328_,
		_w18329_,
		_w18330_
	);
	LUT3 #(
		.INIT('h80)
	) name7818 (
		\wishbone_bd_ram_mem2_reg[132][23]/P0001 ,
		_w11929_,
		_w11955_,
		_w18331_
	);
	LUT3 #(
		.INIT('h80)
	) name7819 (
		\wishbone_bd_ram_mem2_reg[17][23]/P0001 ,
		_w11935_,
		_w11977_,
		_w18332_
	);
	LUT3 #(
		.INIT('h80)
	) name7820 (
		\wishbone_bd_ram_mem2_reg[208][23]/P0001 ,
		_w11941_,
		_w11984_,
		_w18333_
	);
	LUT3 #(
		.INIT('h80)
	) name7821 (
		\wishbone_bd_ram_mem2_reg[49][23]/P0001 ,
		_w11977_,
		_w11979_,
		_w18334_
	);
	LUT4 #(
		.INIT('h0001)
	) name7822 (
		_w18331_,
		_w18332_,
		_w18333_,
		_w18334_,
		_w18335_
	);
	LUT4 #(
		.INIT('h8000)
	) name7823 (
		_w18320_,
		_w18325_,
		_w18330_,
		_w18335_,
		_w18336_
	);
	LUT3 #(
		.INIT('h80)
	) name7824 (
		\wishbone_bd_ram_mem2_reg[120][23]/P0001 ,
		_w11990_,
		_w12012_,
		_w18337_
	);
	LUT3 #(
		.INIT('h80)
	) name7825 (
		\wishbone_bd_ram_mem2_reg[115][23]/P0001 ,
		_w11938_,
		_w12012_,
		_w18338_
	);
	LUT3 #(
		.INIT('h80)
	) name7826 (
		\wishbone_bd_ram_mem2_reg[84][23]/P0001 ,
		_w11929_,
		_w11972_,
		_w18339_
	);
	LUT3 #(
		.INIT('h80)
	) name7827 (
		\wishbone_bd_ram_mem2_reg[16][23]/P0001 ,
		_w11935_,
		_w11941_,
		_w18340_
	);
	LUT4 #(
		.INIT('h0001)
	) name7828 (
		_w18337_,
		_w18338_,
		_w18339_,
		_w18340_,
		_w18341_
	);
	LUT3 #(
		.INIT('h80)
	) name7829 (
		\wishbone_bd_ram_mem2_reg[143][23]/P0001 ,
		_w11955_,
		_w11973_,
		_w18342_
	);
	LUT3 #(
		.INIT('h80)
	) name7830 (
		\wishbone_bd_ram_mem2_reg[152][23]/P0001 ,
		_w11959_,
		_w11990_,
		_w18343_
	);
	LUT3 #(
		.INIT('h80)
	) name7831 (
		\wishbone_bd_ram_mem2_reg[25][23]/P0001 ,
		_w11935_,
		_w11968_,
		_w18344_
	);
	LUT3 #(
		.INIT('h80)
	) name7832 (
		\wishbone_bd_ram_mem2_reg[32][23]/P0001 ,
		_w11941_,
		_w11957_,
		_w18345_
	);
	LUT4 #(
		.INIT('h0001)
	) name7833 (
		_w18342_,
		_w18343_,
		_w18344_,
		_w18345_,
		_w18346_
	);
	LUT3 #(
		.INIT('h80)
	) name7834 (
		\wishbone_bd_ram_mem2_reg[247][23]/P0001 ,
		_w11952_,
		_w11975_,
		_w18347_
	);
	LUT3 #(
		.INIT('h80)
	) name7835 (
		\wishbone_bd_ram_mem2_reg[154][23]/P0001 ,
		_w11944_,
		_w11959_,
		_w18348_
	);
	LUT3 #(
		.INIT('h80)
	) name7836 (
		\wishbone_bd_ram_mem2_reg[93][23]/P0001 ,
		_w11966_,
		_w11972_,
		_w18349_
	);
	LUT3 #(
		.INIT('h80)
	) name7837 (
		\wishbone_bd_ram_mem2_reg[39][23]/P0001 ,
		_w11957_,
		_w11975_,
		_w18350_
	);
	LUT4 #(
		.INIT('h0001)
	) name7838 (
		_w18347_,
		_w18348_,
		_w18349_,
		_w18350_,
		_w18351_
	);
	LUT3 #(
		.INIT('h80)
	) name7839 (
		\wishbone_bd_ram_mem2_reg[33][23]/P0001 ,
		_w11957_,
		_w11977_,
		_w18352_
	);
	LUT3 #(
		.INIT('h80)
	) name7840 (
		\wishbone_bd_ram_mem2_reg[131][23]/P0001 ,
		_w11938_,
		_w11955_,
		_w18353_
	);
	LUT3 #(
		.INIT('h80)
	) name7841 (
		\wishbone_bd_ram_mem2_reg[248][23]/P0001 ,
		_w11952_,
		_w11990_,
		_w18354_
	);
	LUT3 #(
		.INIT('h80)
	) name7842 (
		\wishbone_bd_ram_mem2_reg[15][23]/P0001 ,
		_w11932_,
		_w11973_,
		_w18355_
	);
	LUT4 #(
		.INIT('h0001)
	) name7843 (
		_w18352_,
		_w18353_,
		_w18354_,
		_w18355_,
		_w18356_
	);
	LUT4 #(
		.INIT('h8000)
	) name7844 (
		_w18341_,
		_w18346_,
		_w18351_,
		_w18356_,
		_w18357_
	);
	LUT3 #(
		.INIT('h80)
	) name7845 (
		\wishbone_bd_ram_mem2_reg[170][23]/P0001 ,
		_w11930_,
		_w11944_,
		_w18358_
	);
	LUT3 #(
		.INIT('h80)
	) name7846 (
		\wishbone_bd_ram_mem2_reg[44][23]/P0001 ,
		_w11954_,
		_w11957_,
		_w18359_
	);
	LUT3 #(
		.INIT('h80)
	) name7847 (
		\wishbone_bd_ram_mem2_reg[90][23]/P0001 ,
		_w11944_,
		_w11972_,
		_w18360_
	);
	LUT3 #(
		.INIT('h80)
	) name7848 (
		\wishbone_bd_ram_mem2_reg[198][23]/P0001 ,
		_w11945_,
		_w11986_,
		_w18361_
	);
	LUT4 #(
		.INIT('h0001)
	) name7849 (
		_w18358_,
		_w18359_,
		_w18360_,
		_w18361_,
		_w18362_
	);
	LUT3 #(
		.INIT('h80)
	) name7850 (
		\wishbone_bd_ram_mem2_reg[128][23]/P0001 ,
		_w11941_,
		_w11955_,
		_w18363_
	);
	LUT3 #(
		.INIT('h80)
	) name7851 (
		\wishbone_bd_ram_mem2_reg[184][23]/P0001 ,
		_w11942_,
		_w11990_,
		_w18364_
	);
	LUT3 #(
		.INIT('h80)
	) name7852 (
		\wishbone_bd_ram_mem2_reg[19][23]/P0001 ,
		_w11935_,
		_w11938_,
		_w18365_
	);
	LUT3 #(
		.INIT('h80)
	) name7853 (
		\wishbone_bd_ram_mem2_reg[244][23]/P0001 ,
		_w11929_,
		_w11952_,
		_w18366_
	);
	LUT4 #(
		.INIT('h0001)
	) name7854 (
		_w18363_,
		_w18364_,
		_w18365_,
		_w18366_,
		_w18367_
	);
	LUT3 #(
		.INIT('h80)
	) name7855 (
		\wishbone_bd_ram_mem2_reg[96][23]/P0001 ,
		_w11941_,
		_w11965_,
		_w18368_
	);
	LUT3 #(
		.INIT('h80)
	) name7856 (
		\wishbone_bd_ram_mem2_reg[14][23]/P0001 ,
		_w11932_,
		_w11948_,
		_w18369_
	);
	LUT3 #(
		.INIT('h80)
	) name7857 (
		\wishbone_bd_ram_mem2_reg[89][23]/P0001 ,
		_w11968_,
		_w11972_,
		_w18370_
	);
	LUT3 #(
		.INIT('h80)
	) name7858 (
		\wishbone_bd_ram_mem2_reg[100][23]/P0001 ,
		_w11929_,
		_w11965_,
		_w18371_
	);
	LUT4 #(
		.INIT('h0001)
	) name7859 (
		_w18368_,
		_w18369_,
		_w18370_,
		_w18371_,
		_w18372_
	);
	LUT3 #(
		.INIT('h80)
	) name7860 (
		\wishbone_bd_ram_mem2_reg[216][23]/P0001 ,
		_w11984_,
		_w11990_,
		_w18373_
	);
	LUT3 #(
		.INIT('h80)
	) name7861 (
		\wishbone_bd_ram_mem2_reg[86][23]/P0001 ,
		_w11972_,
		_w11986_,
		_w18374_
	);
	LUT3 #(
		.INIT('h80)
	) name7862 (
		\wishbone_bd_ram_mem2_reg[215][23]/P0001 ,
		_w11975_,
		_w11984_,
		_w18375_
	);
	LUT3 #(
		.INIT('h80)
	) name7863 (
		\wishbone_bd_ram_mem2_reg[145][23]/P0001 ,
		_w11959_,
		_w11977_,
		_w18376_
	);
	LUT4 #(
		.INIT('h0001)
	) name7864 (
		_w18373_,
		_w18374_,
		_w18375_,
		_w18376_,
		_w18377_
	);
	LUT4 #(
		.INIT('h8000)
	) name7865 (
		_w18362_,
		_w18367_,
		_w18372_,
		_w18377_,
		_w18378_
	);
	LUT3 #(
		.INIT('h80)
	) name7866 (
		\wishbone_bd_ram_mem2_reg[52][23]/P0001 ,
		_w11929_,
		_w11979_,
		_w18379_
	);
	LUT3 #(
		.INIT('h80)
	) name7867 (
		\wishbone_bd_ram_mem2_reg[137][23]/P0001 ,
		_w11955_,
		_w11968_,
		_w18380_
	);
	LUT3 #(
		.INIT('h80)
	) name7868 (
		\wishbone_bd_ram_mem2_reg[108][23]/P0001 ,
		_w11954_,
		_w11965_,
		_w18381_
	);
	LUT3 #(
		.INIT('h80)
	) name7869 (
		\wishbone_bd_ram_mem2_reg[60][23]/P0001 ,
		_w11954_,
		_w11979_,
		_w18382_
	);
	LUT4 #(
		.INIT('h0001)
	) name7870 (
		_w18379_,
		_w18380_,
		_w18381_,
		_w18382_,
		_w18383_
	);
	LUT3 #(
		.INIT('h80)
	) name7871 (
		\wishbone_bd_ram_mem2_reg[187][23]/P0001 ,
		_w11936_,
		_w11942_,
		_w18384_
	);
	LUT3 #(
		.INIT('h80)
	) name7872 (
		\wishbone_bd_ram_mem2_reg[185][23]/P0001 ,
		_w11942_,
		_w11968_,
		_w18385_
	);
	LUT3 #(
		.INIT('h80)
	) name7873 (
		\wishbone_bd_ram_mem2_reg[167][23]/P0001 ,
		_w11930_,
		_w11975_,
		_w18386_
	);
	LUT3 #(
		.INIT('h80)
	) name7874 (
		\wishbone_bd_ram_mem2_reg[130][23]/P0001 ,
		_w11955_,
		_w11963_,
		_w18387_
	);
	LUT4 #(
		.INIT('h0001)
	) name7875 (
		_w18384_,
		_w18385_,
		_w18386_,
		_w18387_,
		_w18388_
	);
	LUT3 #(
		.INIT('h80)
	) name7876 (
		\wishbone_bd_ram_mem2_reg[41][23]/P0001 ,
		_w11957_,
		_w11968_,
		_w18389_
	);
	LUT3 #(
		.INIT('h80)
	) name7877 (
		\wishbone_bd_ram_mem2_reg[226][23]/P0001 ,
		_w11963_,
		_w11982_,
		_w18390_
	);
	LUT3 #(
		.INIT('h80)
	) name7878 (
		\wishbone_bd_ram_mem2_reg[165][23]/P0001 ,
		_w11930_,
		_w11933_,
		_w18391_
	);
	LUT3 #(
		.INIT('h80)
	) name7879 (
		\wishbone_bd_ram_mem2_reg[124][23]/P0001 ,
		_w11954_,
		_w12012_,
		_w18392_
	);
	LUT4 #(
		.INIT('h0001)
	) name7880 (
		_w18389_,
		_w18390_,
		_w18391_,
		_w18392_,
		_w18393_
	);
	LUT3 #(
		.INIT('h80)
	) name7881 (
		\wishbone_bd_ram_mem2_reg[45][23]/P0001 ,
		_w11957_,
		_w11966_,
		_w18394_
	);
	LUT3 #(
		.INIT('h80)
	) name7882 (
		\wishbone_bd_ram_mem2_reg[110][23]/P0001 ,
		_w11948_,
		_w11965_,
		_w18395_
	);
	LUT3 #(
		.INIT('h80)
	) name7883 (
		\wishbone_bd_ram_mem2_reg[183][23]/P0001 ,
		_w11942_,
		_w11975_,
		_w18396_
	);
	LUT3 #(
		.INIT('h80)
	) name7884 (
		\wishbone_bd_ram_mem2_reg[171][23]/P0001 ,
		_w11930_,
		_w11936_,
		_w18397_
	);
	LUT4 #(
		.INIT('h0001)
	) name7885 (
		_w18394_,
		_w18395_,
		_w18396_,
		_w18397_,
		_w18398_
	);
	LUT4 #(
		.INIT('h8000)
	) name7886 (
		_w18383_,
		_w18388_,
		_w18393_,
		_w18398_,
		_w18399_
	);
	LUT4 #(
		.INIT('h8000)
	) name7887 (
		_w18336_,
		_w18357_,
		_w18378_,
		_w18399_,
		_w18400_
	);
	LUT4 #(
		.INIT('h8000)
	) name7888 (
		_w18145_,
		_w18230_,
		_w18315_,
		_w18400_,
		_w18401_
	);
	LUT3 #(
		.INIT('hce)
	) name7889 (
		_w12303_,
		_w18060_,
		_w18401_,
		_w18402_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name7890 (
		\wishbone_LatchedTxLength_reg[8]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w18403_
	);
	LUT3 #(
		.INIT('hf2)
	) name7891 (
		_w12303_,
		_w13397_,
		_w18403_,
		_w18404_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name7892 (
		\wishbone_LatchedTxLength_reg[6]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w18405_
	);
	LUT3 #(
		.INIT('h80)
	) name7893 (
		\wishbone_bd_ram_mem2_reg[86][22]/P0001 ,
		_w11972_,
		_w11986_,
		_w18406_
	);
	LUT3 #(
		.INIT('h80)
	) name7894 (
		\wishbone_bd_ram_mem2_reg[79][22]/P0001 ,
		_w11949_,
		_w11973_,
		_w18407_
	);
	LUT3 #(
		.INIT('h80)
	) name7895 (
		\wishbone_bd_ram_mem2_reg[52][22]/P0001 ,
		_w11929_,
		_w11979_,
		_w18408_
	);
	LUT3 #(
		.INIT('h80)
	) name7896 (
		\wishbone_bd_ram_mem2_reg[74][22]/P0001 ,
		_w11944_,
		_w11949_,
		_w18409_
	);
	LUT4 #(
		.INIT('h0001)
	) name7897 (
		_w18406_,
		_w18407_,
		_w18408_,
		_w18409_,
		_w18410_
	);
	LUT3 #(
		.INIT('h80)
	) name7898 (
		\wishbone_bd_ram_mem2_reg[202][22]/P0001 ,
		_w11944_,
		_w11945_,
		_w18411_
	);
	LUT3 #(
		.INIT('h80)
	) name7899 (
		\wishbone_bd_ram_mem2_reg[228][22]/P0001 ,
		_w11929_,
		_w11982_,
		_w18412_
	);
	LUT3 #(
		.INIT('h80)
	) name7900 (
		\wishbone_bd_ram_mem2_reg[64][22]/P0001 ,
		_w11941_,
		_w11949_,
		_w18413_
	);
	LUT3 #(
		.INIT('h80)
	) name7901 (
		\wishbone_bd_ram_mem2_reg[247][22]/P0001 ,
		_w11952_,
		_w11975_,
		_w18414_
	);
	LUT4 #(
		.INIT('h0001)
	) name7902 (
		_w18411_,
		_w18412_,
		_w18413_,
		_w18414_,
		_w18415_
	);
	LUT3 #(
		.INIT('h80)
	) name7903 (
		\wishbone_bd_ram_mem2_reg[133][22]/P0001 ,
		_w11933_,
		_w11955_,
		_w18416_
	);
	LUT3 #(
		.INIT('h80)
	) name7904 (
		\wishbone_bd_ram_mem2_reg[204][22]/P0001 ,
		_w11945_,
		_w11954_,
		_w18417_
	);
	LUT3 #(
		.INIT('h80)
	) name7905 (
		\wishbone_bd_ram_mem2_reg[135][22]/P0001 ,
		_w11955_,
		_w11975_,
		_w18418_
	);
	LUT3 #(
		.INIT('h80)
	) name7906 (
		\wishbone_bd_ram_mem2_reg[111][22]/P0001 ,
		_w11965_,
		_w11973_,
		_w18419_
	);
	LUT4 #(
		.INIT('h0001)
	) name7907 (
		_w18416_,
		_w18417_,
		_w18418_,
		_w18419_,
		_w18420_
	);
	LUT3 #(
		.INIT('h80)
	) name7908 (
		\wishbone_bd_ram_mem2_reg[32][22]/P0001 ,
		_w11941_,
		_w11957_,
		_w18421_
	);
	LUT3 #(
		.INIT('h80)
	) name7909 (
		\wishbone_bd_ram_mem2_reg[194][22]/P0001 ,
		_w11945_,
		_w11963_,
		_w18422_
	);
	LUT3 #(
		.INIT('h80)
	) name7910 (
		\wishbone_bd_ram_mem2_reg[51][22]/P0001 ,
		_w11938_,
		_w11979_,
		_w18423_
	);
	LUT3 #(
		.INIT('h80)
	) name7911 (
		\wishbone_bd_ram_mem2_reg[180][22]/P0001 ,
		_w11929_,
		_w11942_,
		_w18424_
	);
	LUT4 #(
		.INIT('h0001)
	) name7912 (
		_w18421_,
		_w18422_,
		_w18423_,
		_w18424_,
		_w18425_
	);
	LUT4 #(
		.INIT('h8000)
	) name7913 (
		_w18410_,
		_w18415_,
		_w18420_,
		_w18425_,
		_w18426_
	);
	LUT3 #(
		.INIT('h80)
	) name7914 (
		\wishbone_bd_ram_mem2_reg[42][22]/P0001 ,
		_w11944_,
		_w11957_,
		_w18427_
	);
	LUT3 #(
		.INIT('h80)
	) name7915 (
		\wishbone_bd_ram_mem2_reg[107][22]/P0001 ,
		_w11936_,
		_w11965_,
		_w18428_
	);
	LUT3 #(
		.INIT('h80)
	) name7916 (
		\wishbone_bd_ram_mem2_reg[2][22]/P0001 ,
		_w11932_,
		_w11963_,
		_w18429_
	);
	LUT3 #(
		.INIT('h80)
	) name7917 (
		\wishbone_bd_ram_mem2_reg[138][22]/P0001 ,
		_w11944_,
		_w11955_,
		_w18430_
	);
	LUT4 #(
		.INIT('h0001)
	) name7918 (
		_w18427_,
		_w18428_,
		_w18429_,
		_w18430_,
		_w18431_
	);
	LUT3 #(
		.INIT('h80)
	) name7919 (
		\wishbone_bd_ram_mem2_reg[248][22]/P0001 ,
		_w11952_,
		_w11990_,
		_w18432_
	);
	LUT3 #(
		.INIT('h80)
	) name7920 (
		\wishbone_bd_ram_mem2_reg[164][22]/P0001 ,
		_w11929_,
		_w11930_,
		_w18433_
	);
	LUT3 #(
		.INIT('h80)
	) name7921 (
		\wishbone_bd_ram_mem2_reg[251][22]/P0001 ,
		_w11936_,
		_w11952_,
		_w18434_
	);
	LUT3 #(
		.INIT('h80)
	) name7922 (
		\wishbone_bd_ram_mem2_reg[50][22]/P0001 ,
		_w11963_,
		_w11979_,
		_w18435_
	);
	LUT4 #(
		.INIT('h0001)
	) name7923 (
		_w18432_,
		_w18433_,
		_w18434_,
		_w18435_,
		_w18436_
	);
	LUT3 #(
		.INIT('h80)
	) name7924 (
		\wishbone_bd_ram_mem2_reg[174][22]/P0001 ,
		_w11930_,
		_w11948_,
		_w18437_
	);
	LUT3 #(
		.INIT('h80)
	) name7925 (
		\wishbone_bd_ram_mem2_reg[165][22]/P0001 ,
		_w11930_,
		_w11933_,
		_w18438_
	);
	LUT3 #(
		.INIT('h80)
	) name7926 (
		\wishbone_bd_ram_mem2_reg[226][22]/P0001 ,
		_w11963_,
		_w11982_,
		_w18439_
	);
	LUT3 #(
		.INIT('h80)
	) name7927 (
		\wishbone_bd_ram_mem2_reg[243][22]/P0001 ,
		_w11938_,
		_w11952_,
		_w18440_
	);
	LUT4 #(
		.INIT('h0001)
	) name7928 (
		_w18437_,
		_w18438_,
		_w18439_,
		_w18440_,
		_w18441_
	);
	LUT3 #(
		.INIT('h80)
	) name7929 (
		\wishbone_bd_ram_mem2_reg[30][22]/P0001 ,
		_w11935_,
		_w11948_,
		_w18442_
	);
	LUT3 #(
		.INIT('h80)
	) name7930 (
		\wishbone_bd_ram_mem2_reg[212][22]/P0001 ,
		_w11929_,
		_w11984_,
		_w18443_
	);
	LUT3 #(
		.INIT('h80)
	) name7931 (
		\wishbone_bd_ram_mem2_reg[146][22]/P0001 ,
		_w11959_,
		_w11963_,
		_w18444_
	);
	LUT3 #(
		.INIT('h80)
	) name7932 (
		\wishbone_bd_ram_mem2_reg[206][22]/P0001 ,
		_w11945_,
		_w11948_,
		_w18445_
	);
	LUT4 #(
		.INIT('h0001)
	) name7933 (
		_w18442_,
		_w18443_,
		_w18444_,
		_w18445_,
		_w18446_
	);
	LUT4 #(
		.INIT('h8000)
	) name7934 (
		_w18431_,
		_w18436_,
		_w18441_,
		_w18446_,
		_w18447_
	);
	LUT3 #(
		.INIT('h80)
	) name7935 (
		\wishbone_bd_ram_mem2_reg[140][22]/P0001 ,
		_w11954_,
		_w11955_,
		_w18448_
	);
	LUT3 #(
		.INIT('h80)
	) name7936 (
		\wishbone_bd_ram_mem2_reg[59][22]/P0001 ,
		_w11936_,
		_w11979_,
		_w18449_
	);
	LUT3 #(
		.INIT('h80)
	) name7937 (
		\wishbone_bd_ram_mem2_reg[176][22]/P0001 ,
		_w11941_,
		_w11942_,
		_w18450_
	);
	LUT3 #(
		.INIT('h80)
	) name7938 (
		\wishbone_bd_ram_mem2_reg[67][22]/P0001 ,
		_w11938_,
		_w11949_,
		_w18451_
	);
	LUT4 #(
		.INIT('h0001)
	) name7939 (
		_w18448_,
		_w18449_,
		_w18450_,
		_w18451_,
		_w18452_
	);
	LUT3 #(
		.INIT('h80)
	) name7940 (
		\wishbone_bd_ram_mem2_reg[106][22]/P0001 ,
		_w11944_,
		_w11965_,
		_w18453_
	);
	LUT3 #(
		.INIT('h80)
	) name7941 (
		\wishbone_bd_ram_mem2_reg[85][22]/P0001 ,
		_w11933_,
		_w11972_,
		_w18454_
	);
	LUT3 #(
		.INIT('h80)
	) name7942 (
		\wishbone_bd_ram_mem2_reg[221][22]/P0001 ,
		_w11966_,
		_w11984_,
		_w18455_
	);
	LUT3 #(
		.INIT('h80)
	) name7943 (
		\wishbone_bd_ram_mem2_reg[128][22]/P0001 ,
		_w11941_,
		_w11955_,
		_w18456_
	);
	LUT4 #(
		.INIT('h0001)
	) name7944 (
		_w18453_,
		_w18454_,
		_w18455_,
		_w18456_,
		_w18457_
	);
	LUT3 #(
		.INIT('h80)
	) name7945 (
		\wishbone_bd_ram_mem2_reg[104][22]/P0001 ,
		_w11965_,
		_w11990_,
		_w18458_
	);
	LUT3 #(
		.INIT('h80)
	) name7946 (
		\wishbone_bd_ram_mem2_reg[41][22]/P0001 ,
		_w11957_,
		_w11968_,
		_w18459_
	);
	LUT3 #(
		.INIT('h80)
	) name7947 (
		\wishbone_bd_ram_mem2_reg[63][22]/P0001 ,
		_w11973_,
		_w11979_,
		_w18460_
	);
	LUT3 #(
		.INIT('h80)
	) name7948 (
		\wishbone_bd_ram_mem2_reg[210][22]/P0001 ,
		_w11963_,
		_w11984_,
		_w18461_
	);
	LUT4 #(
		.INIT('h0001)
	) name7949 (
		_w18458_,
		_w18459_,
		_w18460_,
		_w18461_,
		_w18462_
	);
	LUT3 #(
		.INIT('h80)
	) name7950 (
		\wishbone_bd_ram_mem2_reg[222][22]/P0001 ,
		_w11948_,
		_w11984_,
		_w18463_
	);
	LUT3 #(
		.INIT('h80)
	) name7951 (
		\wishbone_bd_ram_mem2_reg[254][22]/P0001 ,
		_w11948_,
		_w11952_,
		_w18464_
	);
	LUT3 #(
		.INIT('h80)
	) name7952 (
		\wishbone_bd_ram_mem2_reg[148][22]/P0001 ,
		_w11929_,
		_w11959_,
		_w18465_
	);
	LUT3 #(
		.INIT('h80)
	) name7953 (
		\wishbone_bd_ram_mem2_reg[239][22]/P0001 ,
		_w11973_,
		_w11982_,
		_w18466_
	);
	LUT4 #(
		.INIT('h0001)
	) name7954 (
		_w18463_,
		_w18464_,
		_w18465_,
		_w18466_,
		_w18467_
	);
	LUT4 #(
		.INIT('h8000)
	) name7955 (
		_w18452_,
		_w18457_,
		_w18462_,
		_w18467_,
		_w18468_
	);
	LUT3 #(
		.INIT('h80)
	) name7956 (
		\wishbone_bd_ram_mem2_reg[116][22]/P0001 ,
		_w11929_,
		_w12012_,
		_w18469_
	);
	LUT3 #(
		.INIT('h80)
	) name7957 (
		\wishbone_bd_ram_mem2_reg[144][22]/P0001 ,
		_w11941_,
		_w11959_,
		_w18470_
	);
	LUT3 #(
		.INIT('h80)
	) name7958 (
		\wishbone_bd_ram_mem2_reg[80][22]/P0001 ,
		_w11941_,
		_w11972_,
		_w18471_
	);
	LUT3 #(
		.INIT('h80)
	) name7959 (
		\wishbone_bd_ram_mem2_reg[108][22]/P0001 ,
		_w11954_,
		_w11965_,
		_w18472_
	);
	LUT4 #(
		.INIT('h0001)
	) name7960 (
		_w18469_,
		_w18470_,
		_w18471_,
		_w18472_,
		_w18473_
	);
	LUT3 #(
		.INIT('h80)
	) name7961 (
		\wishbone_bd_ram_mem2_reg[214][22]/P0001 ,
		_w11984_,
		_w11986_,
		_w18474_
	);
	LUT3 #(
		.INIT('h80)
	) name7962 (
		\wishbone_bd_ram_mem2_reg[173][22]/P0001 ,
		_w11930_,
		_w11966_,
		_w18475_
	);
	LUT3 #(
		.INIT('h80)
	) name7963 (
		\wishbone_bd_ram_mem2_reg[60][22]/P0001 ,
		_w11954_,
		_w11979_,
		_w18476_
	);
	LUT3 #(
		.INIT('h80)
	) name7964 (
		\wishbone_bd_ram_mem2_reg[5][22]/P0001 ,
		_w11932_,
		_w11933_,
		_w18477_
	);
	LUT4 #(
		.INIT('h0001)
	) name7965 (
		_w18474_,
		_w18475_,
		_w18476_,
		_w18477_,
		_w18478_
	);
	LUT3 #(
		.INIT('h80)
	) name7966 (
		\wishbone_bd_ram_mem2_reg[97][22]/P0001 ,
		_w11965_,
		_w11977_,
		_w18479_
	);
	LUT3 #(
		.INIT('h80)
	) name7967 (
		\wishbone_bd_ram_mem2_reg[141][22]/P0001 ,
		_w11955_,
		_w11966_,
		_w18480_
	);
	LUT3 #(
		.INIT('h80)
	) name7968 (
		\wishbone_bd_ram_mem2_reg[58][22]/P0001 ,
		_w11944_,
		_w11979_,
		_w18481_
	);
	LUT3 #(
		.INIT('h80)
	) name7969 (
		\wishbone_bd_ram_mem2_reg[0][22]/P0001 ,
		_w11932_,
		_w11941_,
		_w18482_
	);
	LUT4 #(
		.INIT('h0001)
	) name7970 (
		_w18479_,
		_w18480_,
		_w18481_,
		_w18482_,
		_w18483_
	);
	LUT3 #(
		.INIT('h80)
	) name7971 (
		\wishbone_bd_ram_mem2_reg[76][22]/P0001 ,
		_w11949_,
		_w11954_,
		_w18484_
	);
	LUT3 #(
		.INIT('h80)
	) name7972 (
		\wishbone_bd_ram_mem2_reg[14][22]/P0001 ,
		_w11932_,
		_w11948_,
		_w18485_
	);
	LUT3 #(
		.INIT('h80)
	) name7973 (
		\wishbone_bd_ram_mem2_reg[57][22]/P0001 ,
		_w11968_,
		_w11979_,
		_w18486_
	);
	LUT3 #(
		.INIT('h80)
	) name7974 (
		\wishbone_bd_ram_mem2_reg[153][22]/P0001 ,
		_w11959_,
		_w11968_,
		_w18487_
	);
	LUT4 #(
		.INIT('h0001)
	) name7975 (
		_w18484_,
		_w18485_,
		_w18486_,
		_w18487_,
		_w18488_
	);
	LUT4 #(
		.INIT('h8000)
	) name7976 (
		_w18473_,
		_w18478_,
		_w18483_,
		_w18488_,
		_w18489_
	);
	LUT4 #(
		.INIT('h8000)
	) name7977 (
		_w18426_,
		_w18447_,
		_w18468_,
		_w18489_,
		_w18490_
	);
	LUT3 #(
		.INIT('h80)
	) name7978 (
		\wishbone_bd_ram_mem2_reg[160][22]/P0001 ,
		_w11930_,
		_w11941_,
		_w18491_
	);
	LUT3 #(
		.INIT('h80)
	) name7979 (
		\wishbone_bd_ram_mem2_reg[23][22]/P0001 ,
		_w11935_,
		_w11975_,
		_w18492_
	);
	LUT3 #(
		.INIT('h80)
	) name7980 (
		\wishbone_bd_ram_mem2_reg[191][22]/P0001 ,
		_w11942_,
		_w11973_,
		_w18493_
	);
	LUT3 #(
		.INIT('h80)
	) name7981 (
		\wishbone_bd_ram_mem2_reg[98][22]/P0001 ,
		_w11963_,
		_w11965_,
		_w18494_
	);
	LUT4 #(
		.INIT('h0001)
	) name7982 (
		_w18491_,
		_w18492_,
		_w18493_,
		_w18494_,
		_w18495_
	);
	LUT3 #(
		.INIT('h80)
	) name7983 (
		\wishbone_bd_ram_mem2_reg[200][22]/P0001 ,
		_w11945_,
		_w11990_,
		_w18496_
	);
	LUT3 #(
		.INIT('h80)
	) name7984 (
		\wishbone_bd_ram_mem2_reg[139][22]/P0001 ,
		_w11936_,
		_w11955_,
		_w18497_
	);
	LUT3 #(
		.INIT('h80)
	) name7985 (
		\wishbone_bd_ram_mem2_reg[61][22]/P0001 ,
		_w11966_,
		_w11979_,
		_w18498_
	);
	LUT3 #(
		.INIT('h80)
	) name7986 (
		\wishbone_bd_ram_mem2_reg[17][22]/P0001 ,
		_w11935_,
		_w11977_,
		_w18499_
	);
	LUT4 #(
		.INIT('h0001)
	) name7987 (
		_w18496_,
		_w18497_,
		_w18498_,
		_w18499_,
		_w18500_
	);
	LUT3 #(
		.INIT('h80)
	) name7988 (
		\wishbone_bd_ram_mem2_reg[112][22]/P0001 ,
		_w11941_,
		_w12012_,
		_w18501_
	);
	LUT3 #(
		.INIT('h80)
	) name7989 (
		\wishbone_bd_ram_mem2_reg[169][22]/P0001 ,
		_w11930_,
		_w11968_,
		_w18502_
	);
	LUT3 #(
		.INIT('h80)
	) name7990 (
		\wishbone_bd_ram_mem2_reg[105][22]/P0001 ,
		_w11965_,
		_w11968_,
		_w18503_
	);
	LUT3 #(
		.INIT('h80)
	) name7991 (
		\wishbone_bd_ram_mem2_reg[220][22]/P0001 ,
		_w11954_,
		_w11984_,
		_w18504_
	);
	LUT4 #(
		.INIT('h0001)
	) name7992 (
		_w18501_,
		_w18502_,
		_w18503_,
		_w18504_,
		_w18505_
	);
	LUT3 #(
		.INIT('h80)
	) name7993 (
		\wishbone_bd_ram_mem2_reg[75][22]/P0001 ,
		_w11936_,
		_w11949_,
		_w18506_
	);
	LUT3 #(
		.INIT('h80)
	) name7994 (
		\wishbone_bd_ram_mem2_reg[157][22]/P0001 ,
		_w11959_,
		_w11966_,
		_w18507_
	);
	LUT3 #(
		.INIT('h80)
	) name7995 (
		\wishbone_bd_ram_mem2_reg[145][22]/P0001 ,
		_w11959_,
		_w11977_,
		_w18508_
	);
	LUT3 #(
		.INIT('h80)
	) name7996 (
		\wishbone_bd_ram_mem2_reg[237][22]/P0001 ,
		_w11966_,
		_w11982_,
		_w18509_
	);
	LUT4 #(
		.INIT('h0001)
	) name7997 (
		_w18506_,
		_w18507_,
		_w18508_,
		_w18509_,
		_w18510_
	);
	LUT4 #(
		.INIT('h8000)
	) name7998 (
		_w18495_,
		_w18500_,
		_w18505_,
		_w18510_,
		_w18511_
	);
	LUT3 #(
		.INIT('h80)
	) name7999 (
		\wishbone_bd_ram_mem2_reg[56][22]/P0001 ,
		_w11979_,
		_w11990_,
		_w18512_
	);
	LUT3 #(
		.INIT('h80)
	) name8000 (
		\wishbone_bd_ram_mem2_reg[127][22]/P0001 ,
		_w11973_,
		_w12012_,
		_w18513_
	);
	LUT3 #(
		.INIT('h80)
	) name8001 (
		\wishbone_bd_ram_mem2_reg[49][22]/P0001 ,
		_w11977_,
		_w11979_,
		_w18514_
	);
	LUT3 #(
		.INIT('h80)
	) name8002 (
		\wishbone_bd_ram_mem2_reg[15][22]/P0001 ,
		_w11932_,
		_w11973_,
		_w18515_
	);
	LUT4 #(
		.INIT('h0001)
	) name8003 (
		_w18512_,
		_w18513_,
		_w18514_,
		_w18515_,
		_w18516_
	);
	LUT3 #(
		.INIT('h80)
	) name8004 (
		\wishbone_bd_ram_mem2_reg[189][22]/P0001 ,
		_w11942_,
		_w11966_,
		_w18517_
	);
	LUT3 #(
		.INIT('h80)
	) name8005 (
		\wishbone_bd_ram_mem2_reg[166][22]/P0001 ,
		_w11930_,
		_w11986_,
		_w18518_
	);
	LUT3 #(
		.INIT('h80)
	) name8006 (
		\wishbone_bd_ram_mem2_reg[44][22]/P0001 ,
		_w11954_,
		_w11957_,
		_w18519_
	);
	LUT3 #(
		.INIT('h80)
	) name8007 (
		\wishbone_bd_ram_mem2_reg[121][22]/P0001 ,
		_w11968_,
		_w12012_,
		_w18520_
	);
	LUT4 #(
		.INIT('h0001)
	) name8008 (
		_w18517_,
		_w18518_,
		_w18519_,
		_w18520_,
		_w18521_
	);
	LUT3 #(
		.INIT('h80)
	) name8009 (
		\wishbone_bd_ram_mem2_reg[38][22]/P0001 ,
		_w11957_,
		_w11986_,
		_w18522_
	);
	LUT3 #(
		.INIT('h80)
	) name8010 (
		\wishbone_bd_ram_mem2_reg[234][22]/P0001 ,
		_w11944_,
		_w11982_,
		_w18523_
	);
	LUT3 #(
		.INIT('h80)
	) name8011 (
		\wishbone_bd_ram_mem2_reg[20][22]/P0001 ,
		_w11929_,
		_w11935_,
		_w18524_
	);
	LUT3 #(
		.INIT('h80)
	) name8012 (
		\wishbone_bd_ram_mem2_reg[45][22]/P0001 ,
		_w11957_,
		_w11966_,
		_w18525_
	);
	LUT4 #(
		.INIT('h0001)
	) name8013 (
		_w18522_,
		_w18523_,
		_w18524_,
		_w18525_,
		_w18526_
	);
	LUT3 #(
		.INIT('h80)
	) name8014 (
		\wishbone_bd_ram_mem2_reg[156][22]/P0001 ,
		_w11954_,
		_w11959_,
		_w18527_
	);
	LUT3 #(
		.INIT('h80)
	) name8015 (
		\wishbone_bd_ram_mem2_reg[252][22]/P0001 ,
		_w11952_,
		_w11954_,
		_w18528_
	);
	LUT3 #(
		.INIT('h80)
	) name8016 (
		\wishbone_bd_ram_mem2_reg[175][22]/P0001 ,
		_w11930_,
		_w11973_,
		_w18529_
	);
	LUT3 #(
		.INIT('h80)
	) name8017 (
		\wishbone_bd_ram_mem2_reg[53][22]/P0001 ,
		_w11933_,
		_w11979_,
		_w18530_
	);
	LUT4 #(
		.INIT('h0001)
	) name8018 (
		_w18527_,
		_w18528_,
		_w18529_,
		_w18530_,
		_w18531_
	);
	LUT4 #(
		.INIT('h8000)
	) name8019 (
		_w18516_,
		_w18521_,
		_w18526_,
		_w18531_,
		_w18532_
	);
	LUT3 #(
		.INIT('h80)
	) name8020 (
		\wishbone_bd_ram_mem2_reg[35][22]/P0001 ,
		_w11938_,
		_w11957_,
		_w18533_
	);
	LUT3 #(
		.INIT('h80)
	) name8021 (
		\wishbone_bd_ram_mem2_reg[184][22]/P0001 ,
		_w11942_,
		_w11990_,
		_w18534_
	);
	LUT3 #(
		.INIT('h80)
	) name8022 (
		\wishbone_bd_ram_mem2_reg[16][22]/P0001 ,
		_w11935_,
		_w11941_,
		_w18535_
	);
	LUT3 #(
		.INIT('h80)
	) name8023 (
		\wishbone_bd_ram_mem2_reg[130][22]/P0001 ,
		_w11955_,
		_w11963_,
		_w18536_
	);
	LUT4 #(
		.INIT('h0001)
	) name8024 (
		_w18533_,
		_w18534_,
		_w18535_,
		_w18536_,
		_w18537_
	);
	LUT3 #(
		.INIT('h80)
	) name8025 (
		\wishbone_bd_ram_mem2_reg[244][22]/P0001 ,
		_w11929_,
		_w11952_,
		_w18538_
	);
	LUT3 #(
		.INIT('h80)
	) name8026 (
		\wishbone_bd_ram_mem2_reg[215][22]/P0001 ,
		_w11975_,
		_w11984_,
		_w18539_
	);
	LUT3 #(
		.INIT('h80)
	) name8027 (
		\wishbone_bd_ram_mem2_reg[217][22]/P0001 ,
		_w11968_,
		_w11984_,
		_w18540_
	);
	LUT3 #(
		.INIT('h80)
	) name8028 (
		\wishbone_bd_ram_mem2_reg[34][22]/P0001 ,
		_w11957_,
		_w11963_,
		_w18541_
	);
	LUT4 #(
		.INIT('h0001)
	) name8029 (
		_w18538_,
		_w18539_,
		_w18540_,
		_w18541_,
		_w18542_
	);
	LUT3 #(
		.INIT('h80)
	) name8030 (
		\wishbone_bd_ram_mem2_reg[207][22]/P0001 ,
		_w11945_,
		_w11973_,
		_w18543_
	);
	LUT3 #(
		.INIT('h80)
	) name8031 (
		\wishbone_bd_ram_mem2_reg[26][22]/P0001 ,
		_w11935_,
		_w11944_,
		_w18544_
	);
	LUT3 #(
		.INIT('h80)
	) name8032 (
		\wishbone_bd_ram_mem2_reg[154][22]/P0001 ,
		_w11944_,
		_w11959_,
		_w18545_
	);
	LUT3 #(
		.INIT('h80)
	) name8033 (
		\wishbone_bd_ram_mem2_reg[113][22]/P0001 ,
		_w11977_,
		_w12012_,
		_w18546_
	);
	LUT4 #(
		.INIT('h0001)
	) name8034 (
		_w18543_,
		_w18544_,
		_w18545_,
		_w18546_,
		_w18547_
	);
	LUT3 #(
		.INIT('h80)
	) name8035 (
		\wishbone_bd_ram_mem2_reg[143][22]/P0001 ,
		_w11955_,
		_w11973_,
		_w18548_
	);
	LUT3 #(
		.INIT('h80)
	) name8036 (
		\wishbone_bd_ram_mem2_reg[96][22]/P0001 ,
		_w11941_,
		_w11965_,
		_w18549_
	);
	LUT3 #(
		.INIT('h80)
	) name8037 (
		\wishbone_bd_ram_mem2_reg[136][22]/P0001 ,
		_w11955_,
		_w11990_,
		_w18550_
	);
	LUT3 #(
		.INIT('h80)
	) name8038 (
		\wishbone_bd_ram_mem2_reg[137][22]/P0001 ,
		_w11955_,
		_w11968_,
		_w18551_
	);
	LUT4 #(
		.INIT('h0001)
	) name8039 (
		_w18548_,
		_w18549_,
		_w18550_,
		_w18551_,
		_w18552_
	);
	LUT4 #(
		.INIT('h8000)
	) name8040 (
		_w18537_,
		_w18542_,
		_w18547_,
		_w18552_,
		_w18553_
	);
	LUT3 #(
		.INIT('h80)
	) name8041 (
		\wishbone_bd_ram_mem2_reg[18][22]/P0001 ,
		_w11935_,
		_w11963_,
		_w18554_
	);
	LUT3 #(
		.INIT('h80)
	) name8042 (
		\wishbone_bd_ram_mem2_reg[55][22]/P0001 ,
		_w11975_,
		_w11979_,
		_w18555_
	);
	LUT3 #(
		.INIT('h80)
	) name8043 (
		\wishbone_bd_ram_mem2_reg[77][22]/P0001 ,
		_w11949_,
		_w11966_,
		_w18556_
	);
	LUT3 #(
		.INIT('h80)
	) name8044 (
		\wishbone_bd_ram_mem2_reg[66][22]/P0001 ,
		_w11949_,
		_w11963_,
		_w18557_
	);
	LUT4 #(
		.INIT('h0001)
	) name8045 (
		_w18554_,
		_w18555_,
		_w18556_,
		_w18557_,
		_w18558_
	);
	LUT3 #(
		.INIT('h80)
	) name8046 (
		\wishbone_bd_ram_mem2_reg[100][22]/P0001 ,
		_w11929_,
		_w11965_,
		_w18559_
	);
	LUT3 #(
		.INIT('h80)
	) name8047 (
		\wishbone_bd_ram_mem2_reg[246][22]/P0001 ,
		_w11952_,
		_w11986_,
		_w18560_
	);
	LUT3 #(
		.INIT('h80)
	) name8048 (
		\wishbone_bd_ram_mem2_reg[10][22]/P0001 ,
		_w11932_,
		_w11944_,
		_w18561_
	);
	LUT3 #(
		.INIT('h80)
	) name8049 (
		\wishbone_bd_ram_mem2_reg[31][22]/P0001 ,
		_w11935_,
		_w11973_,
		_w18562_
	);
	LUT4 #(
		.INIT('h0001)
	) name8050 (
		_w18559_,
		_w18560_,
		_w18561_,
		_w18562_,
		_w18563_
	);
	LUT3 #(
		.INIT('h80)
	) name8051 (
		\wishbone_bd_ram_mem2_reg[203][22]/P0001 ,
		_w11936_,
		_w11945_,
		_w18564_
	);
	LUT3 #(
		.INIT('h80)
	) name8052 (
		\wishbone_bd_ram_mem2_reg[232][22]/P0001 ,
		_w11982_,
		_w11990_,
		_w18565_
	);
	LUT3 #(
		.INIT('h80)
	) name8053 (
		\wishbone_bd_ram_mem2_reg[159][22]/P0001 ,
		_w11959_,
		_w11973_,
		_w18566_
	);
	LUT3 #(
		.INIT('h80)
	) name8054 (
		\wishbone_bd_ram_mem2_reg[233][22]/P0001 ,
		_w11968_,
		_w11982_,
		_w18567_
	);
	LUT4 #(
		.INIT('h0001)
	) name8055 (
		_w18564_,
		_w18565_,
		_w18566_,
		_w18567_,
		_w18568_
	);
	LUT3 #(
		.INIT('h80)
	) name8056 (
		\wishbone_bd_ram_mem2_reg[114][22]/P0001 ,
		_w11963_,
		_w12012_,
		_w18569_
	);
	LUT3 #(
		.INIT('h80)
	) name8057 (
		\wishbone_bd_ram_mem2_reg[208][22]/P0001 ,
		_w11941_,
		_w11984_,
		_w18570_
	);
	LUT3 #(
		.INIT('h80)
	) name8058 (
		\wishbone_bd_ram_mem2_reg[95][22]/P0001 ,
		_w11972_,
		_w11973_,
		_w18571_
	);
	LUT3 #(
		.INIT('h80)
	) name8059 (
		\wishbone_bd_ram_mem2_reg[24][22]/P0001 ,
		_w11935_,
		_w11990_,
		_w18572_
	);
	LUT4 #(
		.INIT('h0001)
	) name8060 (
		_w18569_,
		_w18570_,
		_w18571_,
		_w18572_,
		_w18573_
	);
	LUT4 #(
		.INIT('h8000)
	) name8061 (
		_w18558_,
		_w18563_,
		_w18568_,
		_w18573_,
		_w18574_
	);
	LUT4 #(
		.INIT('h8000)
	) name8062 (
		_w18511_,
		_w18532_,
		_w18553_,
		_w18574_,
		_w18575_
	);
	LUT3 #(
		.INIT('h80)
	) name8063 (
		\wishbone_bd_ram_mem2_reg[4][22]/P0001 ,
		_w11929_,
		_w11932_,
		_w18576_
	);
	LUT3 #(
		.INIT('h80)
	) name8064 (
		\wishbone_bd_ram_mem2_reg[21][22]/P0001 ,
		_w11933_,
		_w11935_,
		_w18577_
	);
	LUT3 #(
		.INIT('h80)
	) name8065 (
		\wishbone_bd_ram_mem2_reg[167][22]/P0001 ,
		_w11930_,
		_w11975_,
		_w18578_
	);
	LUT3 #(
		.INIT('h80)
	) name8066 (
		\wishbone_bd_ram_mem2_reg[181][22]/P0001 ,
		_w11933_,
		_w11942_,
		_w18579_
	);
	LUT4 #(
		.INIT('h0001)
	) name8067 (
		_w18576_,
		_w18577_,
		_w18578_,
		_w18579_,
		_w18580_
	);
	LUT3 #(
		.INIT('h80)
	) name8068 (
		\wishbone_bd_ram_mem2_reg[149][22]/P0001 ,
		_w11933_,
		_w11959_,
		_w18581_
	);
	LUT3 #(
		.INIT('h80)
	) name8069 (
		\wishbone_bd_ram_mem2_reg[1][22]/P0001 ,
		_w11932_,
		_w11977_,
		_w18582_
	);
	LUT3 #(
		.INIT('h80)
	) name8070 (
		\wishbone_bd_ram_mem2_reg[201][22]/P0001 ,
		_w11945_,
		_w11968_,
		_w18583_
	);
	LUT3 #(
		.INIT('h80)
	) name8071 (
		\wishbone_bd_ram_mem2_reg[117][22]/P0001 ,
		_w11933_,
		_w12012_,
		_w18584_
	);
	LUT4 #(
		.INIT('h0001)
	) name8072 (
		_w18581_,
		_w18582_,
		_w18583_,
		_w18584_,
		_w18585_
	);
	LUT3 #(
		.INIT('h80)
	) name8073 (
		\wishbone_bd_ram_mem2_reg[72][22]/P0001 ,
		_w11949_,
		_w11990_,
		_w18586_
	);
	LUT3 #(
		.INIT('h80)
	) name8074 (
		\wishbone_bd_ram_mem2_reg[9][22]/P0001 ,
		_w11932_,
		_w11968_,
		_w18587_
	);
	LUT3 #(
		.INIT('h80)
	) name8075 (
		\wishbone_bd_ram_mem2_reg[90][22]/P0001 ,
		_w11944_,
		_w11972_,
		_w18588_
	);
	LUT3 #(
		.INIT('h80)
	) name8076 (
		\wishbone_bd_ram_mem2_reg[168][22]/P0001 ,
		_w11930_,
		_w11990_,
		_w18589_
	);
	LUT4 #(
		.INIT('h0001)
	) name8077 (
		_w18586_,
		_w18587_,
		_w18588_,
		_w18589_,
		_w18590_
	);
	LUT3 #(
		.INIT('h80)
	) name8078 (
		\wishbone_bd_ram_mem2_reg[47][22]/P0001 ,
		_w11957_,
		_w11973_,
		_w18591_
	);
	LUT3 #(
		.INIT('h80)
	) name8079 (
		\wishbone_bd_ram_mem2_reg[125][22]/P0001 ,
		_w11966_,
		_w12012_,
		_w18592_
	);
	LUT3 #(
		.INIT('h80)
	) name8080 (
		\wishbone_bd_ram_mem2_reg[216][22]/P0001 ,
		_w11984_,
		_w11990_,
		_w18593_
	);
	LUT3 #(
		.INIT('h80)
	) name8081 (
		\wishbone_bd_ram_mem2_reg[19][22]/P0001 ,
		_w11935_,
		_w11938_,
		_w18594_
	);
	LUT4 #(
		.INIT('h0001)
	) name8082 (
		_w18591_,
		_w18592_,
		_w18593_,
		_w18594_,
		_w18595_
	);
	LUT4 #(
		.INIT('h8000)
	) name8083 (
		_w18580_,
		_w18585_,
		_w18590_,
		_w18595_,
		_w18596_
	);
	LUT3 #(
		.INIT('h80)
	) name8084 (
		\wishbone_bd_ram_mem2_reg[250][22]/P0001 ,
		_w11944_,
		_w11952_,
		_w18597_
	);
	LUT3 #(
		.INIT('h80)
	) name8085 (
		\wishbone_bd_ram_mem2_reg[12][22]/P0001 ,
		_w11932_,
		_w11954_,
		_w18598_
	);
	LUT3 #(
		.INIT('h80)
	) name8086 (
		\wishbone_bd_ram_mem2_reg[27][22]/P0001 ,
		_w11935_,
		_w11936_,
		_w18599_
	);
	LUT3 #(
		.INIT('h80)
	) name8087 (
		\wishbone_bd_ram_mem2_reg[88][22]/P0001 ,
		_w11972_,
		_w11990_,
		_w18600_
	);
	LUT4 #(
		.INIT('h0001)
	) name8088 (
		_w18597_,
		_w18598_,
		_w18599_,
		_w18600_,
		_w18601_
	);
	LUT3 #(
		.INIT('h80)
	) name8089 (
		\wishbone_bd_ram_mem2_reg[187][22]/P0001 ,
		_w11936_,
		_w11942_,
		_w18602_
	);
	LUT3 #(
		.INIT('h80)
	) name8090 (
		\wishbone_bd_ram_mem2_reg[172][22]/P0001 ,
		_w11930_,
		_w11954_,
		_w18603_
	);
	LUT3 #(
		.INIT('h80)
	) name8091 (
		\wishbone_bd_ram_mem2_reg[109][22]/P0001 ,
		_w11965_,
		_w11966_,
		_w18604_
	);
	LUT3 #(
		.INIT('h80)
	) name8092 (
		\wishbone_bd_ram_mem2_reg[82][22]/P0001 ,
		_w11963_,
		_w11972_,
		_w18605_
	);
	LUT4 #(
		.INIT('h0001)
	) name8093 (
		_w18602_,
		_w18603_,
		_w18604_,
		_w18605_,
		_w18606_
	);
	LUT3 #(
		.INIT('h80)
	) name8094 (
		\wishbone_bd_ram_mem2_reg[131][22]/P0001 ,
		_w11938_,
		_w11955_,
		_w18607_
	);
	LUT3 #(
		.INIT('h80)
	) name8095 (
		\wishbone_bd_ram_mem2_reg[68][22]/P0001 ,
		_w11929_,
		_w11949_,
		_w18608_
	);
	LUT3 #(
		.INIT('h80)
	) name8096 (
		\wishbone_bd_ram_mem2_reg[196][22]/P0001 ,
		_w11929_,
		_w11945_,
		_w18609_
	);
	LUT3 #(
		.INIT('h80)
	) name8097 (
		\wishbone_bd_ram_mem2_reg[115][22]/P0001 ,
		_w11938_,
		_w12012_,
		_w18610_
	);
	LUT4 #(
		.INIT('h0001)
	) name8098 (
		_w18607_,
		_w18608_,
		_w18609_,
		_w18610_,
		_w18611_
	);
	LUT3 #(
		.INIT('h80)
	) name8099 (
		\wishbone_bd_ram_mem2_reg[11][22]/P0001 ,
		_w11932_,
		_w11936_,
		_w18612_
	);
	LUT3 #(
		.INIT('h80)
	) name8100 (
		\wishbone_bd_ram_mem2_reg[147][22]/P0001 ,
		_w11938_,
		_w11959_,
		_w18613_
	);
	LUT3 #(
		.INIT('h80)
	) name8101 (
		\wishbone_bd_ram_mem2_reg[36][22]/P0001 ,
		_w11929_,
		_w11957_,
		_w18614_
	);
	LUT3 #(
		.INIT('h80)
	) name8102 (
		\wishbone_bd_ram_mem2_reg[87][22]/P0001 ,
		_w11972_,
		_w11975_,
		_w18615_
	);
	LUT4 #(
		.INIT('h0001)
	) name8103 (
		_w18612_,
		_w18613_,
		_w18614_,
		_w18615_,
		_w18616_
	);
	LUT4 #(
		.INIT('h8000)
	) name8104 (
		_w18601_,
		_w18606_,
		_w18611_,
		_w18616_,
		_w18617_
	);
	LUT3 #(
		.INIT('h80)
	) name8105 (
		\wishbone_bd_ram_mem2_reg[190][22]/P0001 ,
		_w11942_,
		_w11948_,
		_w18618_
	);
	LUT3 #(
		.INIT('h80)
	) name8106 (
		\wishbone_bd_ram_mem2_reg[22][22]/P0001 ,
		_w11935_,
		_w11986_,
		_w18619_
	);
	LUT3 #(
		.INIT('h80)
	) name8107 (
		\wishbone_bd_ram_mem2_reg[89][22]/P0001 ,
		_w11968_,
		_w11972_,
		_w18620_
	);
	LUT3 #(
		.INIT('h80)
	) name8108 (
		\wishbone_bd_ram_mem2_reg[197][22]/P0001 ,
		_w11933_,
		_w11945_,
		_w18621_
	);
	LUT4 #(
		.INIT('h0001)
	) name8109 (
		_w18618_,
		_w18619_,
		_w18620_,
		_w18621_,
		_w18622_
	);
	LUT3 #(
		.INIT('h80)
	) name8110 (
		\wishbone_bd_ram_mem2_reg[94][22]/P0001 ,
		_w11948_,
		_w11972_,
		_w18623_
	);
	LUT3 #(
		.INIT('h80)
	) name8111 (
		\wishbone_bd_ram_mem2_reg[177][22]/P0001 ,
		_w11942_,
		_w11977_,
		_w18624_
	);
	LUT3 #(
		.INIT('h80)
	) name8112 (
		\wishbone_bd_ram_mem2_reg[155][22]/P0001 ,
		_w11936_,
		_w11959_,
		_w18625_
	);
	LUT3 #(
		.INIT('h80)
	) name8113 (
		\wishbone_bd_ram_mem2_reg[48][22]/P0001 ,
		_w11941_,
		_w11979_,
		_w18626_
	);
	LUT4 #(
		.INIT('h0001)
	) name8114 (
		_w18623_,
		_w18624_,
		_w18625_,
		_w18626_,
		_w18627_
	);
	LUT3 #(
		.INIT('h80)
	) name8115 (
		\wishbone_bd_ram_mem2_reg[69][22]/P0001 ,
		_w11933_,
		_w11949_,
		_w18628_
	);
	LUT3 #(
		.INIT('h80)
	) name8116 (
		\wishbone_bd_ram_mem2_reg[188][22]/P0001 ,
		_w11942_,
		_w11954_,
		_w18629_
	);
	LUT3 #(
		.INIT('h80)
	) name8117 (
		\wishbone_bd_ram_mem2_reg[118][22]/P0001 ,
		_w11986_,
		_w12012_,
		_w18630_
	);
	LUT3 #(
		.INIT('h80)
	) name8118 (
		\wishbone_bd_ram_mem2_reg[161][22]/P0001 ,
		_w11930_,
		_w11977_,
		_w18631_
	);
	LUT4 #(
		.INIT('h0001)
	) name8119 (
		_w18628_,
		_w18629_,
		_w18630_,
		_w18631_,
		_w18632_
	);
	LUT3 #(
		.INIT('h80)
	) name8120 (
		\wishbone_bd_ram_mem2_reg[39][22]/P0001 ,
		_w11957_,
		_w11975_,
		_w18633_
	);
	LUT3 #(
		.INIT('h80)
	) name8121 (
		\wishbone_bd_ram_mem2_reg[142][22]/P0001 ,
		_w11948_,
		_w11955_,
		_w18634_
	);
	LUT3 #(
		.INIT('h80)
	) name8122 (
		\wishbone_bd_ram_mem2_reg[122][22]/P0001 ,
		_w11944_,
		_w12012_,
		_w18635_
	);
	LUT3 #(
		.INIT('h80)
	) name8123 (
		\wishbone_bd_ram_mem2_reg[83][22]/P0001 ,
		_w11938_,
		_w11972_,
		_w18636_
	);
	LUT4 #(
		.INIT('h0001)
	) name8124 (
		_w18633_,
		_w18634_,
		_w18635_,
		_w18636_,
		_w18637_
	);
	LUT4 #(
		.INIT('h8000)
	) name8125 (
		_w18622_,
		_w18627_,
		_w18632_,
		_w18637_,
		_w18638_
	);
	LUT3 #(
		.INIT('h80)
	) name8126 (
		\wishbone_bd_ram_mem2_reg[179][22]/P0001 ,
		_w11938_,
		_w11942_,
		_w18639_
	);
	LUT3 #(
		.INIT('h80)
	) name8127 (
		\wishbone_bd_ram_mem2_reg[126][22]/P0001 ,
		_w11948_,
		_w12012_,
		_w18640_
	);
	LUT3 #(
		.INIT('h80)
	) name8128 (
		\wishbone_bd_ram_mem2_reg[7][22]/P0001 ,
		_w11932_,
		_w11975_,
		_w18641_
	);
	LUT3 #(
		.INIT('h80)
	) name8129 (
		\wishbone_bd_ram_mem2_reg[209][22]/P0001 ,
		_w11977_,
		_w11984_,
		_w18642_
	);
	LUT4 #(
		.INIT('h0001)
	) name8130 (
		_w18639_,
		_w18640_,
		_w18641_,
		_w18642_,
		_w18643_
	);
	LUT3 #(
		.INIT('h80)
	) name8131 (
		\wishbone_bd_ram_mem2_reg[120][22]/P0001 ,
		_w11990_,
		_w12012_,
		_w18644_
	);
	LUT3 #(
		.INIT('h80)
	) name8132 (
		\wishbone_bd_ram_mem2_reg[242][22]/P0001 ,
		_w11952_,
		_w11963_,
		_w18645_
	);
	LUT3 #(
		.INIT('h80)
	) name8133 (
		\wishbone_bd_ram_mem2_reg[249][22]/P0001 ,
		_w11952_,
		_w11968_,
		_w18646_
	);
	LUT3 #(
		.INIT('h80)
	) name8134 (
		\wishbone_bd_ram_mem2_reg[223][22]/P0001 ,
		_w11973_,
		_w11984_,
		_w18647_
	);
	LUT4 #(
		.INIT('h0001)
	) name8135 (
		_w18644_,
		_w18645_,
		_w18646_,
		_w18647_,
		_w18648_
	);
	LUT3 #(
		.INIT('h80)
	) name8136 (
		\wishbone_bd_ram_mem2_reg[240][22]/P0001 ,
		_w11941_,
		_w11952_,
		_w18649_
	);
	LUT3 #(
		.INIT('h80)
	) name8137 (
		\wishbone_bd_ram_mem2_reg[29][22]/P0001 ,
		_w11935_,
		_w11966_,
		_w18650_
	);
	LUT3 #(
		.INIT('h80)
	) name8138 (
		\wishbone_bd_ram_mem2_reg[25][22]/P0001 ,
		_w11935_,
		_w11968_,
		_w18651_
	);
	LUT3 #(
		.INIT('h80)
	) name8139 (
		\wishbone_bd_ram_mem2_reg[124][22]/P0001 ,
		_w11954_,
		_w12012_,
		_w18652_
	);
	LUT4 #(
		.INIT('h0001)
	) name8140 (
		_w18649_,
		_w18650_,
		_w18651_,
		_w18652_,
		_w18653_
	);
	LUT3 #(
		.INIT('h80)
	) name8141 (
		\wishbone_bd_ram_mem2_reg[253][22]/P0001 ,
		_w11952_,
		_w11966_,
		_w18654_
	);
	LUT3 #(
		.INIT('h80)
	) name8142 (
		\wishbone_bd_ram_mem2_reg[84][22]/P0001 ,
		_w11929_,
		_w11972_,
		_w18655_
	);
	LUT3 #(
		.INIT('h80)
	) name8143 (
		\wishbone_bd_ram_mem2_reg[8][22]/P0001 ,
		_w11932_,
		_w11990_,
		_w18656_
	);
	LUT3 #(
		.INIT('h80)
	) name8144 (
		\wishbone_bd_ram_mem2_reg[37][22]/P0001 ,
		_w11933_,
		_w11957_,
		_w18657_
	);
	LUT4 #(
		.INIT('h0001)
	) name8145 (
		_w18654_,
		_w18655_,
		_w18656_,
		_w18657_,
		_w18658_
	);
	LUT4 #(
		.INIT('h8000)
	) name8146 (
		_w18643_,
		_w18648_,
		_w18653_,
		_w18658_,
		_w18659_
	);
	LUT4 #(
		.INIT('h8000)
	) name8147 (
		_w18596_,
		_w18617_,
		_w18638_,
		_w18659_,
		_w18660_
	);
	LUT3 #(
		.INIT('h80)
	) name8148 (
		\wishbone_bd_ram_mem2_reg[70][22]/P0001 ,
		_w11949_,
		_w11986_,
		_w18661_
	);
	LUT3 #(
		.INIT('h80)
	) name8149 (
		\wishbone_bd_ram_mem2_reg[129][22]/P0001 ,
		_w11955_,
		_w11977_,
		_w18662_
	);
	LUT3 #(
		.INIT('h80)
	) name8150 (
		\wishbone_bd_ram_mem2_reg[54][22]/P0001 ,
		_w11979_,
		_w11986_,
		_w18663_
	);
	LUT3 #(
		.INIT('h80)
	) name8151 (
		\wishbone_bd_ram_mem2_reg[73][22]/P0001 ,
		_w11949_,
		_w11968_,
		_w18664_
	);
	LUT4 #(
		.INIT('h0001)
	) name8152 (
		_w18661_,
		_w18662_,
		_w18663_,
		_w18664_,
		_w18665_
	);
	LUT3 #(
		.INIT('h80)
	) name8153 (
		\wishbone_bd_ram_mem2_reg[170][22]/P0001 ,
		_w11930_,
		_w11944_,
		_w18666_
	);
	LUT3 #(
		.INIT('h80)
	) name8154 (
		\wishbone_bd_ram_mem2_reg[152][22]/P0001 ,
		_w11959_,
		_w11990_,
		_w18667_
	);
	LUT3 #(
		.INIT('h80)
	) name8155 (
		\wishbone_bd_ram_mem2_reg[62][22]/P0001 ,
		_w11948_,
		_w11979_,
		_w18668_
	);
	LUT3 #(
		.INIT('h80)
	) name8156 (
		\wishbone_bd_ram_mem2_reg[229][22]/P0001 ,
		_w11933_,
		_w11982_,
		_w18669_
	);
	LUT4 #(
		.INIT('h0001)
	) name8157 (
		_w18666_,
		_w18667_,
		_w18668_,
		_w18669_,
		_w18670_
	);
	LUT3 #(
		.INIT('h80)
	) name8158 (
		\wishbone_bd_ram_mem2_reg[81][22]/P0001 ,
		_w11972_,
		_w11977_,
		_w18671_
	);
	LUT3 #(
		.INIT('h80)
	) name8159 (
		\wishbone_bd_ram_mem2_reg[238][22]/P0001 ,
		_w11948_,
		_w11982_,
		_w18672_
	);
	LUT3 #(
		.INIT('h80)
	) name8160 (
		\wishbone_bd_ram_mem2_reg[28][22]/P0001 ,
		_w11935_,
		_w11954_,
		_w18673_
	);
	LUT3 #(
		.INIT('h80)
	) name8161 (
		\wishbone_bd_ram_mem2_reg[183][22]/P0001 ,
		_w11942_,
		_w11975_,
		_w18674_
	);
	LUT4 #(
		.INIT('h0001)
	) name8162 (
		_w18671_,
		_w18672_,
		_w18673_,
		_w18674_,
		_w18675_
	);
	LUT3 #(
		.INIT('h80)
	) name8163 (
		\wishbone_bd_ram_mem2_reg[163][22]/P0001 ,
		_w11930_,
		_w11938_,
		_w18676_
	);
	LUT3 #(
		.INIT('h80)
	) name8164 (
		\wishbone_bd_ram_mem2_reg[255][22]/P0001 ,
		_w11952_,
		_w11973_,
		_w18677_
	);
	LUT3 #(
		.INIT('h80)
	) name8165 (
		\wishbone_bd_ram_mem2_reg[99][22]/P0001 ,
		_w11938_,
		_w11965_,
		_w18678_
	);
	LUT3 #(
		.INIT('h80)
	) name8166 (
		\wishbone_bd_ram_mem2_reg[119][22]/P0001 ,
		_w11975_,
		_w12012_,
		_w18679_
	);
	LUT4 #(
		.INIT('h0001)
	) name8167 (
		_w18676_,
		_w18677_,
		_w18678_,
		_w18679_,
		_w18680_
	);
	LUT4 #(
		.INIT('h8000)
	) name8168 (
		_w18665_,
		_w18670_,
		_w18675_,
		_w18680_,
		_w18681_
	);
	LUT3 #(
		.INIT('h80)
	) name8169 (
		\wishbone_bd_ram_mem2_reg[151][22]/P0001 ,
		_w11959_,
		_w11975_,
		_w18682_
	);
	LUT3 #(
		.INIT('h80)
	) name8170 (
		\wishbone_bd_ram_mem2_reg[6][22]/P0001 ,
		_w11932_,
		_w11986_,
		_w18683_
	);
	LUT3 #(
		.INIT('h80)
	) name8171 (
		\wishbone_bd_ram_mem2_reg[230][22]/P0001 ,
		_w11982_,
		_w11986_,
		_w18684_
	);
	LUT3 #(
		.INIT('h80)
	) name8172 (
		\wishbone_bd_ram_mem2_reg[102][22]/P0001 ,
		_w11965_,
		_w11986_,
		_w18685_
	);
	LUT4 #(
		.INIT('h0001)
	) name8173 (
		_w18682_,
		_w18683_,
		_w18684_,
		_w18685_,
		_w18686_
	);
	LUT3 #(
		.INIT('h80)
	) name8174 (
		\wishbone_bd_ram_mem2_reg[192][22]/P0001 ,
		_w11941_,
		_w11945_,
		_w18687_
	);
	LUT3 #(
		.INIT('h80)
	) name8175 (
		\wishbone_bd_ram_mem2_reg[134][22]/P0001 ,
		_w11955_,
		_w11986_,
		_w18688_
	);
	LUT3 #(
		.INIT('h80)
	) name8176 (
		\wishbone_bd_ram_mem2_reg[225][22]/P0001 ,
		_w11977_,
		_w11982_,
		_w18689_
	);
	LUT3 #(
		.INIT('h80)
	) name8177 (
		\wishbone_bd_ram_mem2_reg[91][22]/P0001 ,
		_w11936_,
		_w11972_,
		_w18690_
	);
	LUT4 #(
		.INIT('h0001)
	) name8178 (
		_w18687_,
		_w18688_,
		_w18689_,
		_w18690_,
		_w18691_
	);
	LUT3 #(
		.INIT('h80)
	) name8179 (
		\wishbone_bd_ram_mem2_reg[224][22]/P0001 ,
		_w11941_,
		_w11982_,
		_w18692_
	);
	LUT3 #(
		.INIT('h80)
	) name8180 (
		\wishbone_bd_ram_mem2_reg[186][22]/P0001 ,
		_w11942_,
		_w11944_,
		_w18693_
	);
	LUT3 #(
		.INIT('h80)
	) name8181 (
		\wishbone_bd_ram_mem2_reg[193][22]/P0001 ,
		_w11945_,
		_w11977_,
		_w18694_
	);
	LUT3 #(
		.INIT('h80)
	) name8182 (
		\wishbone_bd_ram_mem2_reg[78][22]/P0001 ,
		_w11948_,
		_w11949_,
		_w18695_
	);
	LUT4 #(
		.INIT('h0001)
	) name8183 (
		_w18692_,
		_w18693_,
		_w18694_,
		_w18695_,
		_w18696_
	);
	LUT3 #(
		.INIT('h80)
	) name8184 (
		\wishbone_bd_ram_mem2_reg[40][22]/P0001 ,
		_w11957_,
		_w11990_,
		_w18697_
	);
	LUT3 #(
		.INIT('h80)
	) name8185 (
		\wishbone_bd_ram_mem2_reg[65][22]/P0001 ,
		_w11949_,
		_w11977_,
		_w18698_
	);
	LUT3 #(
		.INIT('h80)
	) name8186 (
		\wishbone_bd_ram_mem2_reg[213][22]/P0001 ,
		_w11933_,
		_w11984_,
		_w18699_
	);
	LUT3 #(
		.INIT('h80)
	) name8187 (
		\wishbone_bd_ram_mem2_reg[71][22]/P0001 ,
		_w11949_,
		_w11975_,
		_w18700_
	);
	LUT4 #(
		.INIT('h0001)
	) name8188 (
		_w18697_,
		_w18698_,
		_w18699_,
		_w18700_,
		_w18701_
	);
	LUT4 #(
		.INIT('h8000)
	) name8189 (
		_w18686_,
		_w18691_,
		_w18696_,
		_w18701_,
		_w18702_
	);
	LUT3 #(
		.INIT('h80)
	) name8190 (
		\wishbone_bd_ram_mem2_reg[199][22]/P0001 ,
		_w11945_,
		_w11975_,
		_w18703_
	);
	LUT3 #(
		.INIT('h80)
	) name8191 (
		\wishbone_bd_ram_mem2_reg[235][22]/P0001 ,
		_w11936_,
		_w11982_,
		_w18704_
	);
	LUT3 #(
		.INIT('h80)
	) name8192 (
		\wishbone_bd_ram_mem2_reg[185][22]/P0001 ,
		_w11942_,
		_w11968_,
		_w18705_
	);
	LUT3 #(
		.INIT('h80)
	) name8193 (
		\wishbone_bd_ram_mem2_reg[241][22]/P0001 ,
		_w11952_,
		_w11977_,
		_w18706_
	);
	LUT4 #(
		.INIT('h0001)
	) name8194 (
		_w18703_,
		_w18704_,
		_w18705_,
		_w18706_,
		_w18707_
	);
	LUT3 #(
		.INIT('h80)
	) name8195 (
		\wishbone_bd_ram_mem2_reg[92][22]/P0001 ,
		_w11954_,
		_w11972_,
		_w18708_
	);
	LUT3 #(
		.INIT('h80)
	) name8196 (
		\wishbone_bd_ram_mem2_reg[195][22]/P0001 ,
		_w11938_,
		_w11945_,
		_w18709_
	);
	LUT3 #(
		.INIT('h80)
	) name8197 (
		\wishbone_bd_ram_mem2_reg[150][22]/P0001 ,
		_w11959_,
		_w11986_,
		_w18710_
	);
	LUT3 #(
		.INIT('h80)
	) name8198 (
		\wishbone_bd_ram_mem2_reg[211][22]/P0001 ,
		_w11938_,
		_w11984_,
		_w18711_
	);
	LUT4 #(
		.INIT('h0001)
	) name8199 (
		_w18708_,
		_w18709_,
		_w18710_,
		_w18711_,
		_w18712_
	);
	LUT3 #(
		.INIT('h80)
	) name8200 (
		\wishbone_bd_ram_mem2_reg[13][22]/P0001 ,
		_w11932_,
		_w11966_,
		_w18713_
	);
	LUT3 #(
		.INIT('h80)
	) name8201 (
		\wishbone_bd_ram_mem2_reg[101][22]/P0001 ,
		_w11933_,
		_w11965_,
		_w18714_
	);
	LUT3 #(
		.INIT('h80)
	) name8202 (
		\wishbone_bd_ram_mem2_reg[43][22]/P0001 ,
		_w11936_,
		_w11957_,
		_w18715_
	);
	LUT3 #(
		.INIT('h80)
	) name8203 (
		\wishbone_bd_ram_mem2_reg[110][22]/P0001 ,
		_w11948_,
		_w11965_,
		_w18716_
	);
	LUT4 #(
		.INIT('h0001)
	) name8204 (
		_w18713_,
		_w18714_,
		_w18715_,
		_w18716_,
		_w18717_
	);
	LUT3 #(
		.INIT('h80)
	) name8205 (
		\wishbone_bd_ram_mem2_reg[227][22]/P0001 ,
		_w11938_,
		_w11982_,
		_w18718_
	);
	LUT3 #(
		.INIT('h80)
	) name8206 (
		\wishbone_bd_ram_mem2_reg[182][22]/P0001 ,
		_w11942_,
		_w11986_,
		_w18719_
	);
	LUT3 #(
		.INIT('h80)
	) name8207 (
		\wishbone_bd_ram_mem2_reg[219][22]/P0001 ,
		_w11936_,
		_w11984_,
		_w18720_
	);
	LUT3 #(
		.INIT('h80)
	) name8208 (
		\wishbone_bd_ram_mem2_reg[3][22]/P0001 ,
		_w11932_,
		_w11938_,
		_w18721_
	);
	LUT4 #(
		.INIT('h0001)
	) name8209 (
		_w18718_,
		_w18719_,
		_w18720_,
		_w18721_,
		_w18722_
	);
	LUT4 #(
		.INIT('h8000)
	) name8210 (
		_w18707_,
		_w18712_,
		_w18717_,
		_w18722_,
		_w18723_
	);
	LUT3 #(
		.INIT('h80)
	) name8211 (
		\wishbone_bd_ram_mem2_reg[231][22]/P0001 ,
		_w11975_,
		_w11982_,
		_w18724_
	);
	LUT3 #(
		.INIT('h80)
	) name8212 (
		\wishbone_bd_ram_mem2_reg[123][22]/P0001 ,
		_w11936_,
		_w12012_,
		_w18725_
	);
	LUT3 #(
		.INIT('h80)
	) name8213 (
		\wishbone_bd_ram_mem2_reg[171][22]/P0001 ,
		_w11930_,
		_w11936_,
		_w18726_
	);
	LUT3 #(
		.INIT('h80)
	) name8214 (
		\wishbone_bd_ram_mem2_reg[103][22]/P0001 ,
		_w11965_,
		_w11975_,
		_w18727_
	);
	LUT4 #(
		.INIT('h0001)
	) name8215 (
		_w18724_,
		_w18725_,
		_w18726_,
		_w18727_,
		_w18728_
	);
	LUT3 #(
		.INIT('h80)
	) name8216 (
		\wishbone_bd_ram_mem2_reg[245][22]/P0001 ,
		_w11933_,
		_w11952_,
		_w18729_
	);
	LUT3 #(
		.INIT('h80)
	) name8217 (
		\wishbone_bd_ram_mem2_reg[236][22]/P0001 ,
		_w11954_,
		_w11982_,
		_w18730_
	);
	LUT3 #(
		.INIT('h80)
	) name8218 (
		\wishbone_bd_ram_mem2_reg[218][22]/P0001 ,
		_w11944_,
		_w11984_,
		_w18731_
	);
	LUT3 #(
		.INIT('h80)
	) name8219 (
		\wishbone_bd_ram_mem2_reg[162][22]/P0001 ,
		_w11930_,
		_w11963_,
		_w18732_
	);
	LUT4 #(
		.INIT('h0001)
	) name8220 (
		_w18729_,
		_w18730_,
		_w18731_,
		_w18732_,
		_w18733_
	);
	LUT3 #(
		.INIT('h80)
	) name8221 (
		\wishbone_bd_ram_mem2_reg[46][22]/P0001 ,
		_w11948_,
		_w11957_,
		_w18734_
	);
	LUT3 #(
		.INIT('h80)
	) name8222 (
		\wishbone_bd_ram_mem2_reg[178][22]/P0001 ,
		_w11942_,
		_w11963_,
		_w18735_
	);
	LUT3 #(
		.INIT('h80)
	) name8223 (
		\wishbone_bd_ram_mem2_reg[198][22]/P0001 ,
		_w11945_,
		_w11986_,
		_w18736_
	);
	LUT3 #(
		.INIT('h80)
	) name8224 (
		\wishbone_bd_ram_mem2_reg[132][22]/P0001 ,
		_w11929_,
		_w11955_,
		_w18737_
	);
	LUT4 #(
		.INIT('h0001)
	) name8225 (
		_w18734_,
		_w18735_,
		_w18736_,
		_w18737_,
		_w18738_
	);
	LUT3 #(
		.INIT('h80)
	) name8226 (
		\wishbone_bd_ram_mem2_reg[93][22]/P0001 ,
		_w11966_,
		_w11972_,
		_w18739_
	);
	LUT3 #(
		.INIT('h80)
	) name8227 (
		\wishbone_bd_ram_mem2_reg[158][22]/P0001 ,
		_w11948_,
		_w11959_,
		_w18740_
	);
	LUT3 #(
		.INIT('h80)
	) name8228 (
		\wishbone_bd_ram_mem2_reg[33][22]/P0001 ,
		_w11957_,
		_w11977_,
		_w18741_
	);
	LUT3 #(
		.INIT('h80)
	) name8229 (
		\wishbone_bd_ram_mem2_reg[205][22]/P0001 ,
		_w11945_,
		_w11966_,
		_w18742_
	);
	LUT4 #(
		.INIT('h0001)
	) name8230 (
		_w18739_,
		_w18740_,
		_w18741_,
		_w18742_,
		_w18743_
	);
	LUT4 #(
		.INIT('h8000)
	) name8231 (
		_w18728_,
		_w18733_,
		_w18738_,
		_w18743_,
		_w18744_
	);
	LUT4 #(
		.INIT('h8000)
	) name8232 (
		_w18681_,
		_w18702_,
		_w18723_,
		_w18744_,
		_w18745_
	);
	LUT4 #(
		.INIT('h8000)
	) name8233 (
		_w18490_,
		_w18575_,
		_w18660_,
		_w18745_,
		_w18746_
	);
	LUT3 #(
		.INIT('hce)
	) name8234 (
		_w12303_,
		_w18405_,
		_w18746_,
		_w18747_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name8235 (
		\wishbone_LatchedTxLength_reg[9]/NET0131 ,
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w18748_
	);
	LUT3 #(
		.INIT('hf2)
	) name8236 (
		_w12303_,
		_w15222_,
		_w18748_,
		_w18749_
	);
	LUT4 #(
		.INIT('h0001)
	) name8237 (
		\wb_sel_i[0]_pad ,
		\wb_sel_i[1]_pad ,
		\wb_sel_i[2]_pad ,
		\wb_sel_i[3]_pad ,
		_w18750_
	);
	LUT4 #(
		.INIT('h1000)
	) name8238 (
		\wb_adr_i[10]_pad ,
		\wb_adr_i[11]_pad ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w18751_
	);
	LUT3 #(
		.INIT('h10)
	) name8239 (
		wb_we_i_pad,
		_w18750_,
		_w18751_,
		_w18752_
	);
	LUT4 #(
		.INIT('h0001)
	) name8240 (
		\wb_adr_i[6]_pad ,
		\wb_adr_i[7]_pad ,
		\wb_adr_i[8]_pad ,
		\wb_adr_i[9]_pad ,
		_w18753_
	);
	LUT4 #(
		.INIT('h0040)
	) name8241 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w18754_
	);
	LUT2 #(
		.INIT('h8)
	) name8242 (
		_w18753_,
		_w18754_,
		_w18755_
	);
	LUT3 #(
		.INIT('h80)
	) name8243 (
		\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 ,
		_w18753_,
		_w18754_,
		_w18756_
	);
	LUT3 #(
		.INIT('h02)
	) name8244 (
		\wb_adr_i[6]_pad ,
		\wb_adr_i[7]_pad ,
		\wb_adr_i[9]_pad ,
		_w18757_
	);
	LUT2 #(
		.INIT('h1)
	) name8245 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[8]_pad ,
		_w18758_
	);
	LUT3 #(
		.INIT('h02)
	) name8246 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w18759_
	);
	LUT4 #(
		.INIT('h0008)
	) name8247 (
		\ethreg1_RXHASH0_2_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w18760_
	);
	LUT3 #(
		.INIT('h80)
	) name8248 (
		_w18757_,
		_w18758_,
		_w18760_,
		_w18761_
	);
	LUT2 #(
		.INIT('h2)
	) name8249 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[8]_pad ,
		_w18762_
	);
	LUT4 #(
		.INIT('h0008)
	) name8250 (
		\ethreg1_RXHASH1_2_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w18763_
	);
	LUT3 #(
		.INIT('h80)
	) name8251 (
		_w18757_,
		_w18762_,
		_w18763_,
		_w18764_
	);
	LUT3 #(
		.INIT('h01)
	) name8252 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w18765_
	);
	LUT4 #(
		.INIT('h0002)
	) name8253 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w18766_
	);
	LUT3 #(
		.INIT('h80)
	) name8254 (
		_w18757_,
		_w18758_,
		_w18766_,
		_w18767_
	);
	LUT4 #(
		.INIT('h0002)
	) name8255 (
		_w18752_,
		_w18761_,
		_w18764_,
		_w18767_,
		_w18768_
	);
	LUT3 #(
		.INIT('h8a)
	) name8256 (
		_w18752_,
		_w18756_,
		_w18768_,
		_w18769_
	);
	LUT3 #(
		.INIT('h45)
	) name8257 (
		wb_rst_i_pad,
		_w18756_,
		_w18768_,
		_w18770_
	);
	LUT3 #(
		.INIT('hdc)
	) name8258 (
		_w18058_,
		_w18769_,
		_w18770_,
		_w18771_
	);
	LUT3 #(
		.INIT('h80)
	) name8259 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		_w18753_,
		_w18754_,
		_w18772_
	);
	LUT4 #(
		.INIT('h0008)
	) name8260 (
		\ethreg1_RXHASH0_2_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w18773_
	);
	LUT3 #(
		.INIT('h80)
	) name8261 (
		_w18757_,
		_w18758_,
		_w18773_,
		_w18774_
	);
	LUT4 #(
		.INIT('h0008)
	) name8262 (
		\ethreg1_RXHASH1_2_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w18775_
	);
	LUT3 #(
		.INIT('h80)
	) name8263 (
		_w18757_,
		_w18762_,
		_w18775_,
		_w18776_
	);
	LUT4 #(
		.INIT('h0002)
	) name8264 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w18777_
	);
	LUT3 #(
		.INIT('h80)
	) name8265 (
		_w18757_,
		_w18758_,
		_w18777_,
		_w18778_
	);
	LUT4 #(
		.INIT('h0002)
	) name8266 (
		_w18752_,
		_w18774_,
		_w18776_,
		_w18778_,
		_w18779_
	);
	LUT3 #(
		.INIT('h8a)
	) name8267 (
		_w18752_,
		_w18772_,
		_w18779_,
		_w18780_
	);
	LUT3 #(
		.INIT('h45)
	) name8268 (
		wb_rst_i_pad,
		_w18772_,
		_w18779_,
		_w18781_
	);
	LUT3 #(
		.INIT('hdc)
	) name8269 (
		_w18746_,
		_w18780_,
		_w18781_,
		_w18782_
	);
	LUT4 #(
		.INIT('h0002)
	) name8270 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w18783_
	);
	LUT3 #(
		.INIT('h80)
	) name8271 (
		_w18757_,
		_w18762_,
		_w18783_,
		_w18784_
	);
	LUT4 #(
		.INIT('h0004)
	) name8272 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[6]_pad ,
		\wb_adr_i[8]_pad ,
		_w18785_
	);
	LUT4 #(
		.INIT('h0008)
	) name8273 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[5]_pad ,
		\wb_adr_i[7]_pad ,
		\wb_adr_i[9]_pad ,
		_w18786_
	);
	LUT3 #(
		.INIT('h80)
	) name8274 (
		\ethreg1_MIIRX_DATA_DataOut_reg[12]/NET0131 ,
		_w18785_,
		_w18786_,
		_w18787_
	);
	LUT4 #(
		.INIT('h0008)
	) name8275 (
		\ethreg1_RXHASH0_1_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w18788_
	);
	LUT3 #(
		.INIT('h80)
	) name8276 (
		_w18757_,
		_w18758_,
		_w18788_,
		_w18789_
	);
	LUT4 #(
		.INIT('h0008)
	) name8277 (
		\ethreg1_RXHASH1_1_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w18790_
	);
	LUT3 #(
		.INIT('h80)
	) name8278 (
		_w18757_,
		_w18762_,
		_w18790_,
		_w18791_
	);
	LUT4 #(
		.INIT('h0001)
	) name8279 (
		_w18784_,
		_w18787_,
		_w18789_,
		_w18791_,
		_w18792_
	);
	LUT4 #(
		.INIT('h0002)
	) name8280 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w18793_
	);
	LUT3 #(
		.INIT('h04)
	) name8281 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w18794_
	);
	LUT4 #(
		.INIT('h0020)
	) name8282 (
		\ethreg1_TXCTRL_1_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w18795_
	);
	LUT4 #(
		.INIT('h777f)
	) name8283 (
		_w18757_,
		_w18758_,
		_w18793_,
		_w18795_,
		_w18796_
	);
	LUT2 #(
		.INIT('h8)
	) name8284 (
		_w18752_,
		_w18796_,
		_w18797_
	);
	LUT4 #(
		.INIT('h0004)
	) name8285 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[5]_pad ,
		\wb_adr_i[7]_pad ,
		\wb_adr_i[9]_pad ,
		_w18798_
	);
	LUT3 #(
		.INIT('h80)
	) name8286 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[4]/NET0131 ,
		_w18785_,
		_w18798_,
		_w18799_
	);
	LUT4 #(
		.INIT('h0001)
	) name8287 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[5]_pad ,
		\wb_adr_i[7]_pad ,
		\wb_adr_i[9]_pad ,
		_w18800_
	);
	LUT4 #(
		.INIT('h0001)
	) name8288 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[6]_pad ,
		\wb_adr_i[8]_pad ,
		_w18801_
	);
	LUT2 #(
		.INIT('h8)
	) name8289 (
		_w18800_,
		_w18801_,
		_w18802_
	);
	LUT3 #(
		.INIT('h80)
	) name8290 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		_w18800_,
		_w18801_,
		_w18803_
	);
	LUT3 #(
		.INIT('h80)
	) name8291 (
		\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 ,
		_w18753_,
		_w18754_,
		_w18804_
	);
	LUT4 #(
		.INIT('h0008)
	) name8292 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[6]_pad ,
		\wb_adr_i[8]_pad ,
		_w18805_
	);
	LUT3 #(
		.INIT('h80)
	) name8293 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[4]/NET0131 ,
		_w18798_,
		_w18805_,
		_w18806_
	);
	LUT4 #(
		.INIT('h0001)
	) name8294 (
		_w18799_,
		_w18803_,
		_w18804_,
		_w18806_,
		_w18807_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name8295 (
		_w18752_,
		_w18792_,
		_w18796_,
		_w18807_,
		_w18808_
	);
	LUT3 #(
		.INIT('h80)
	) name8296 (
		\wishbone_bd_ram_mem1_reg[43][12]/P0001 ,
		_w11936_,
		_w11957_,
		_w18809_
	);
	LUT3 #(
		.INIT('h80)
	) name8297 (
		\wishbone_bd_ram_mem1_reg[135][12]/P0001 ,
		_w11955_,
		_w11975_,
		_w18810_
	);
	LUT3 #(
		.INIT('h80)
	) name8298 (
		\wishbone_bd_ram_mem1_reg[103][12]/P0001 ,
		_w11965_,
		_w11975_,
		_w18811_
	);
	LUT3 #(
		.INIT('h80)
	) name8299 (
		\wishbone_bd_ram_mem1_reg[219][12]/P0001 ,
		_w11936_,
		_w11984_,
		_w18812_
	);
	LUT4 #(
		.INIT('h0001)
	) name8300 (
		_w18809_,
		_w18810_,
		_w18811_,
		_w18812_,
		_w18813_
	);
	LUT3 #(
		.INIT('h80)
	) name8301 (
		\wishbone_bd_ram_mem1_reg[82][12]/P0001 ,
		_w11963_,
		_w11972_,
		_w18814_
	);
	LUT3 #(
		.INIT('h80)
	) name8302 (
		\wishbone_bd_ram_mem1_reg[55][12]/P0001 ,
		_w11975_,
		_w11979_,
		_w18815_
	);
	LUT3 #(
		.INIT('h80)
	) name8303 (
		\wishbone_bd_ram_mem1_reg[205][12]/P0001 ,
		_w11945_,
		_w11966_,
		_w18816_
	);
	LUT3 #(
		.INIT('h80)
	) name8304 (
		\wishbone_bd_ram_mem1_reg[175][12]/P0001 ,
		_w11930_,
		_w11973_,
		_w18817_
	);
	LUT4 #(
		.INIT('h0001)
	) name8305 (
		_w18814_,
		_w18815_,
		_w18816_,
		_w18817_,
		_w18818_
	);
	LUT3 #(
		.INIT('h80)
	) name8306 (
		\wishbone_bd_ram_mem1_reg[252][12]/P0001 ,
		_w11952_,
		_w11954_,
		_w18819_
	);
	LUT3 #(
		.INIT('h80)
	) name8307 (
		\wishbone_bd_ram_mem1_reg[180][12]/P0001 ,
		_w11929_,
		_w11942_,
		_w18820_
	);
	LUT3 #(
		.INIT('h80)
	) name8308 (
		\wishbone_bd_ram_mem1_reg[1][12]/P0001 ,
		_w11932_,
		_w11977_,
		_w18821_
	);
	LUT3 #(
		.INIT('h80)
	) name8309 (
		\wishbone_bd_ram_mem1_reg[31][12]/P0001 ,
		_w11935_,
		_w11973_,
		_w18822_
	);
	LUT4 #(
		.INIT('h0001)
	) name8310 (
		_w18819_,
		_w18820_,
		_w18821_,
		_w18822_,
		_w18823_
	);
	LUT3 #(
		.INIT('h80)
	) name8311 (
		\wishbone_bd_ram_mem1_reg[112][12]/P0001 ,
		_w11941_,
		_w12012_,
		_w18824_
	);
	LUT3 #(
		.INIT('h80)
	) name8312 (
		\wishbone_bd_ram_mem1_reg[249][12]/P0001 ,
		_w11952_,
		_w11968_,
		_w18825_
	);
	LUT3 #(
		.INIT('h80)
	) name8313 (
		\wishbone_bd_ram_mem1_reg[201][12]/P0001 ,
		_w11945_,
		_w11968_,
		_w18826_
	);
	LUT3 #(
		.INIT('h80)
	) name8314 (
		\wishbone_bd_ram_mem1_reg[47][12]/P0001 ,
		_w11957_,
		_w11973_,
		_w18827_
	);
	LUT4 #(
		.INIT('h0001)
	) name8315 (
		_w18824_,
		_w18825_,
		_w18826_,
		_w18827_,
		_w18828_
	);
	LUT4 #(
		.INIT('h8000)
	) name8316 (
		_w18813_,
		_w18818_,
		_w18823_,
		_w18828_,
		_w18829_
	);
	LUT3 #(
		.INIT('h80)
	) name8317 (
		\wishbone_bd_ram_mem1_reg[118][12]/P0001 ,
		_w11986_,
		_w12012_,
		_w18830_
	);
	LUT3 #(
		.INIT('h80)
	) name8318 (
		\wishbone_bd_ram_mem1_reg[231][12]/P0001 ,
		_w11975_,
		_w11982_,
		_w18831_
	);
	LUT3 #(
		.INIT('h80)
	) name8319 (
		\wishbone_bd_ram_mem1_reg[121][12]/P0001 ,
		_w11968_,
		_w12012_,
		_w18832_
	);
	LUT3 #(
		.INIT('h80)
	) name8320 (
		\wishbone_bd_ram_mem1_reg[229][12]/P0001 ,
		_w11933_,
		_w11982_,
		_w18833_
	);
	LUT4 #(
		.INIT('h0001)
	) name8321 (
		_w18830_,
		_w18831_,
		_w18832_,
		_w18833_,
		_w18834_
	);
	LUT3 #(
		.INIT('h80)
	) name8322 (
		\wishbone_bd_ram_mem1_reg[193][12]/P0001 ,
		_w11945_,
		_w11977_,
		_w18835_
	);
	LUT3 #(
		.INIT('h80)
	) name8323 (
		\wishbone_bd_ram_mem1_reg[126][12]/P0001 ,
		_w11948_,
		_w12012_,
		_w18836_
	);
	LUT3 #(
		.INIT('h80)
	) name8324 (
		\wishbone_bd_ram_mem1_reg[35][12]/P0001 ,
		_w11938_,
		_w11957_,
		_w18837_
	);
	LUT3 #(
		.INIT('h80)
	) name8325 (
		\wishbone_bd_ram_mem1_reg[191][12]/P0001 ,
		_w11942_,
		_w11973_,
		_w18838_
	);
	LUT4 #(
		.INIT('h0001)
	) name8326 (
		_w18835_,
		_w18836_,
		_w18837_,
		_w18838_,
		_w18839_
	);
	LUT3 #(
		.INIT('h80)
	) name8327 (
		\wishbone_bd_ram_mem1_reg[104][12]/P0001 ,
		_w11965_,
		_w11990_,
		_w18840_
	);
	LUT3 #(
		.INIT('h80)
	) name8328 (
		\wishbone_bd_ram_mem1_reg[248][12]/P0001 ,
		_w11952_,
		_w11990_,
		_w18841_
	);
	LUT3 #(
		.INIT('h80)
	) name8329 (
		\wishbone_bd_ram_mem1_reg[241][12]/P0001 ,
		_w11952_,
		_w11977_,
		_w18842_
	);
	LUT3 #(
		.INIT('h80)
	) name8330 (
		\wishbone_bd_ram_mem1_reg[127][12]/P0001 ,
		_w11973_,
		_w12012_,
		_w18843_
	);
	LUT4 #(
		.INIT('h0001)
	) name8331 (
		_w18840_,
		_w18841_,
		_w18842_,
		_w18843_,
		_w18844_
	);
	LUT3 #(
		.INIT('h80)
	) name8332 (
		\wishbone_bd_ram_mem1_reg[144][12]/P0001 ,
		_w11941_,
		_w11959_,
		_w18845_
	);
	LUT3 #(
		.INIT('h80)
	) name8333 (
		\wishbone_bd_ram_mem1_reg[49][12]/P0001 ,
		_w11977_,
		_w11979_,
		_w18846_
	);
	LUT3 #(
		.INIT('h80)
	) name8334 (
		\wishbone_bd_ram_mem1_reg[220][12]/P0001 ,
		_w11954_,
		_w11984_,
		_w18847_
	);
	LUT3 #(
		.INIT('h80)
	) name8335 (
		\wishbone_bd_ram_mem1_reg[210][12]/P0001 ,
		_w11963_,
		_w11984_,
		_w18848_
	);
	LUT4 #(
		.INIT('h0001)
	) name8336 (
		_w18845_,
		_w18846_,
		_w18847_,
		_w18848_,
		_w18849_
	);
	LUT4 #(
		.INIT('h8000)
	) name8337 (
		_w18834_,
		_w18839_,
		_w18844_,
		_w18849_,
		_w18850_
	);
	LUT3 #(
		.INIT('h80)
	) name8338 (
		\wishbone_bd_ram_mem1_reg[8][12]/P0001 ,
		_w11932_,
		_w11990_,
		_w18851_
	);
	LUT3 #(
		.INIT('h80)
	) name8339 (
		\wishbone_bd_ram_mem1_reg[245][12]/P0001 ,
		_w11933_,
		_w11952_,
		_w18852_
	);
	LUT3 #(
		.INIT('h80)
	) name8340 (
		\wishbone_bd_ram_mem1_reg[105][12]/P0001 ,
		_w11965_,
		_w11968_,
		_w18853_
	);
	LUT3 #(
		.INIT('h80)
	) name8341 (
		\wishbone_bd_ram_mem1_reg[106][12]/P0001 ,
		_w11944_,
		_w11965_,
		_w18854_
	);
	LUT4 #(
		.INIT('h0001)
	) name8342 (
		_w18851_,
		_w18852_,
		_w18853_,
		_w18854_,
		_w18855_
	);
	LUT3 #(
		.INIT('h80)
	) name8343 (
		\wishbone_bd_ram_mem1_reg[243][12]/P0001 ,
		_w11938_,
		_w11952_,
		_w18856_
	);
	LUT3 #(
		.INIT('h80)
	) name8344 (
		\wishbone_bd_ram_mem1_reg[96][12]/P0001 ,
		_w11941_,
		_w11965_,
		_w18857_
	);
	LUT3 #(
		.INIT('h80)
	) name8345 (
		\wishbone_bd_ram_mem1_reg[239][12]/P0001 ,
		_w11973_,
		_w11982_,
		_w18858_
	);
	LUT3 #(
		.INIT('h80)
	) name8346 (
		\wishbone_bd_ram_mem1_reg[7][12]/P0001 ,
		_w11932_,
		_w11975_,
		_w18859_
	);
	LUT4 #(
		.INIT('h0001)
	) name8347 (
		_w18856_,
		_w18857_,
		_w18858_,
		_w18859_,
		_w18860_
	);
	LUT3 #(
		.INIT('h80)
	) name8348 (
		\wishbone_bd_ram_mem1_reg[230][12]/P0001 ,
		_w11982_,
		_w11986_,
		_w18861_
	);
	LUT3 #(
		.INIT('h80)
	) name8349 (
		\wishbone_bd_ram_mem1_reg[158][12]/P0001 ,
		_w11948_,
		_w11959_,
		_w18862_
	);
	LUT3 #(
		.INIT('h80)
	) name8350 (
		\wishbone_bd_ram_mem1_reg[187][12]/P0001 ,
		_w11936_,
		_w11942_,
		_w18863_
	);
	LUT3 #(
		.INIT('h80)
	) name8351 (
		\wishbone_bd_ram_mem1_reg[54][12]/P0001 ,
		_w11979_,
		_w11986_,
		_w18864_
	);
	LUT4 #(
		.INIT('h0001)
	) name8352 (
		_w18861_,
		_w18862_,
		_w18863_,
		_w18864_,
		_w18865_
	);
	LUT3 #(
		.INIT('h80)
	) name8353 (
		\wishbone_bd_ram_mem1_reg[129][12]/P0001 ,
		_w11955_,
		_w11977_,
		_w18866_
	);
	LUT3 #(
		.INIT('h80)
	) name8354 (
		\wishbone_bd_ram_mem1_reg[215][12]/P0001 ,
		_w11975_,
		_w11984_,
		_w18867_
	);
	LUT3 #(
		.INIT('h80)
	) name8355 (
		\wishbone_bd_ram_mem1_reg[52][12]/P0001 ,
		_w11929_,
		_w11979_,
		_w18868_
	);
	LUT3 #(
		.INIT('h80)
	) name8356 (
		\wishbone_bd_ram_mem1_reg[147][12]/P0001 ,
		_w11938_,
		_w11959_,
		_w18869_
	);
	LUT4 #(
		.INIT('h0001)
	) name8357 (
		_w18866_,
		_w18867_,
		_w18868_,
		_w18869_,
		_w18870_
	);
	LUT4 #(
		.INIT('h8000)
	) name8358 (
		_w18855_,
		_w18860_,
		_w18865_,
		_w18870_,
		_w18871_
	);
	LUT3 #(
		.INIT('h80)
	) name8359 (
		\wishbone_bd_ram_mem1_reg[216][12]/P0001 ,
		_w11984_,
		_w11990_,
		_w18872_
	);
	LUT3 #(
		.INIT('h80)
	) name8360 (
		\wishbone_bd_ram_mem1_reg[174][12]/P0001 ,
		_w11930_,
		_w11948_,
		_w18873_
	);
	LUT3 #(
		.INIT('h80)
	) name8361 (
		\wishbone_bd_ram_mem1_reg[77][12]/P0001 ,
		_w11949_,
		_w11966_,
		_w18874_
	);
	LUT3 #(
		.INIT('h80)
	) name8362 (
		\wishbone_bd_ram_mem1_reg[120][12]/P0001 ,
		_w11990_,
		_w12012_,
		_w18875_
	);
	LUT4 #(
		.INIT('h0001)
	) name8363 (
		_w18872_,
		_w18873_,
		_w18874_,
		_w18875_,
		_w18876_
	);
	LUT3 #(
		.INIT('h80)
	) name8364 (
		\wishbone_bd_ram_mem1_reg[227][12]/P0001 ,
		_w11938_,
		_w11982_,
		_w18877_
	);
	LUT3 #(
		.INIT('h80)
	) name8365 (
		\wishbone_bd_ram_mem1_reg[199][12]/P0001 ,
		_w11945_,
		_w11975_,
		_w18878_
	);
	LUT3 #(
		.INIT('h80)
	) name8366 (
		\wishbone_bd_ram_mem1_reg[244][12]/P0001 ,
		_w11929_,
		_w11952_,
		_w18879_
	);
	LUT3 #(
		.INIT('h80)
	) name8367 (
		\wishbone_bd_ram_mem1_reg[26][12]/P0001 ,
		_w11935_,
		_w11944_,
		_w18880_
	);
	LUT4 #(
		.INIT('h0001)
	) name8368 (
		_w18877_,
		_w18878_,
		_w18879_,
		_w18880_,
		_w18881_
	);
	LUT3 #(
		.INIT('h80)
	) name8369 (
		\wishbone_bd_ram_mem1_reg[155][12]/P0001 ,
		_w11936_,
		_w11959_,
		_w18882_
	);
	LUT3 #(
		.INIT('h80)
	) name8370 (
		\wishbone_bd_ram_mem1_reg[27][12]/P0001 ,
		_w11935_,
		_w11936_,
		_w18883_
	);
	LUT3 #(
		.INIT('h80)
	) name8371 (
		\wishbone_bd_ram_mem1_reg[111][12]/P0001 ,
		_w11965_,
		_w11973_,
		_w18884_
	);
	LUT3 #(
		.INIT('h80)
	) name8372 (
		\wishbone_bd_ram_mem1_reg[225][12]/P0001 ,
		_w11977_,
		_w11982_,
		_w18885_
	);
	LUT4 #(
		.INIT('h0001)
	) name8373 (
		_w18882_,
		_w18883_,
		_w18884_,
		_w18885_,
		_w18886_
	);
	LUT3 #(
		.INIT('h80)
	) name8374 (
		\wishbone_bd_ram_mem1_reg[217][12]/P0001 ,
		_w11968_,
		_w11984_,
		_w18887_
	);
	LUT3 #(
		.INIT('h80)
	) name8375 (
		\wishbone_bd_ram_mem1_reg[234][12]/P0001 ,
		_w11944_,
		_w11982_,
		_w18888_
	);
	LUT3 #(
		.INIT('h80)
	) name8376 (
		\wishbone_bd_ram_mem1_reg[5][12]/P0001 ,
		_w11932_,
		_w11933_,
		_w18889_
	);
	LUT3 #(
		.INIT('h80)
	) name8377 (
		\wishbone_bd_ram_mem1_reg[62][12]/P0001 ,
		_w11948_,
		_w11979_,
		_w18890_
	);
	LUT4 #(
		.INIT('h0001)
	) name8378 (
		_w18887_,
		_w18888_,
		_w18889_,
		_w18890_,
		_w18891_
	);
	LUT4 #(
		.INIT('h8000)
	) name8379 (
		_w18876_,
		_w18881_,
		_w18886_,
		_w18891_,
		_w18892_
	);
	LUT4 #(
		.INIT('h8000)
	) name8380 (
		_w18829_,
		_w18850_,
		_w18871_,
		_w18892_,
		_w18893_
	);
	LUT3 #(
		.INIT('h80)
	) name8381 (
		\wishbone_bd_ram_mem1_reg[33][12]/P0001 ,
		_w11957_,
		_w11977_,
		_w18894_
	);
	LUT3 #(
		.INIT('h80)
	) name8382 (
		\wishbone_bd_ram_mem1_reg[238][12]/P0001 ,
		_w11948_,
		_w11982_,
		_w18895_
	);
	LUT3 #(
		.INIT('h80)
	) name8383 (
		\wishbone_bd_ram_mem1_reg[153][12]/P0001 ,
		_w11959_,
		_w11968_,
		_w18896_
	);
	LUT3 #(
		.INIT('h80)
	) name8384 (
		\wishbone_bd_ram_mem1_reg[24][12]/P0001 ,
		_w11935_,
		_w11990_,
		_w18897_
	);
	LUT4 #(
		.INIT('h0001)
	) name8385 (
		_w18894_,
		_w18895_,
		_w18896_,
		_w18897_,
		_w18898_
	);
	LUT3 #(
		.INIT('h80)
	) name8386 (
		\wishbone_bd_ram_mem1_reg[212][12]/P0001 ,
		_w11929_,
		_w11984_,
		_w18899_
	);
	LUT3 #(
		.INIT('h80)
	) name8387 (
		\wishbone_bd_ram_mem1_reg[59][12]/P0001 ,
		_w11936_,
		_w11979_,
		_w18900_
	);
	LUT3 #(
		.INIT('h80)
	) name8388 (
		\wishbone_bd_ram_mem1_reg[85][12]/P0001 ,
		_w11933_,
		_w11972_,
		_w18901_
	);
	LUT3 #(
		.INIT('h80)
	) name8389 (
		\wishbone_bd_ram_mem1_reg[90][12]/P0001 ,
		_w11944_,
		_w11972_,
		_w18902_
	);
	LUT4 #(
		.INIT('h0001)
	) name8390 (
		_w18899_,
		_w18900_,
		_w18901_,
		_w18902_,
		_w18903_
	);
	LUT3 #(
		.INIT('h80)
	) name8391 (
		\wishbone_bd_ram_mem1_reg[139][12]/P0001 ,
		_w11936_,
		_w11955_,
		_w18904_
	);
	LUT3 #(
		.INIT('h80)
	) name8392 (
		\wishbone_bd_ram_mem1_reg[97][12]/P0001 ,
		_w11965_,
		_w11977_,
		_w18905_
	);
	LUT3 #(
		.INIT('h80)
	) name8393 (
		\wishbone_bd_ram_mem1_reg[232][12]/P0001 ,
		_w11982_,
		_w11990_,
		_w18906_
	);
	LUT3 #(
		.INIT('h80)
	) name8394 (
		\wishbone_bd_ram_mem1_reg[223][12]/P0001 ,
		_w11973_,
		_w11984_,
		_w18907_
	);
	LUT4 #(
		.INIT('h0001)
	) name8395 (
		_w18904_,
		_w18905_,
		_w18906_,
		_w18907_,
		_w18908_
	);
	LUT3 #(
		.INIT('h80)
	) name8396 (
		\wishbone_bd_ram_mem1_reg[165][12]/P0001 ,
		_w11930_,
		_w11933_,
		_w18909_
	);
	LUT3 #(
		.INIT('h80)
	) name8397 (
		\wishbone_bd_ram_mem1_reg[146][12]/P0001 ,
		_w11959_,
		_w11963_,
		_w18910_
	);
	LUT3 #(
		.INIT('h80)
	) name8398 (
		\wishbone_bd_ram_mem1_reg[128][12]/P0001 ,
		_w11941_,
		_w11955_,
		_w18911_
	);
	LUT3 #(
		.INIT('h80)
	) name8399 (
		\wishbone_bd_ram_mem1_reg[28][12]/P0001 ,
		_w11935_,
		_w11954_,
		_w18912_
	);
	LUT4 #(
		.INIT('h0001)
	) name8400 (
		_w18909_,
		_w18910_,
		_w18911_,
		_w18912_,
		_w18913_
	);
	LUT4 #(
		.INIT('h8000)
	) name8401 (
		_w18898_,
		_w18903_,
		_w18908_,
		_w18913_,
		_w18914_
	);
	LUT3 #(
		.INIT('h80)
	) name8402 (
		\wishbone_bd_ram_mem1_reg[236][12]/P0001 ,
		_w11954_,
		_w11982_,
		_w18915_
	);
	LUT3 #(
		.INIT('h80)
	) name8403 (
		\wishbone_bd_ram_mem1_reg[86][12]/P0001 ,
		_w11972_,
		_w11986_,
		_w18916_
	);
	LUT3 #(
		.INIT('h80)
	) name8404 (
		\wishbone_bd_ram_mem1_reg[161][12]/P0001 ,
		_w11930_,
		_w11977_,
		_w18917_
	);
	LUT3 #(
		.INIT('h80)
	) name8405 (
		\wishbone_bd_ram_mem1_reg[117][12]/P0001 ,
		_w11933_,
		_w12012_,
		_w18918_
	);
	LUT4 #(
		.INIT('h0001)
	) name8406 (
		_w18915_,
		_w18916_,
		_w18917_,
		_w18918_,
		_w18919_
	);
	LUT3 #(
		.INIT('h80)
	) name8407 (
		\wishbone_bd_ram_mem1_reg[17][12]/P0001 ,
		_w11935_,
		_w11977_,
		_w18920_
	);
	LUT3 #(
		.INIT('h80)
	) name8408 (
		\wishbone_bd_ram_mem1_reg[95][12]/P0001 ,
		_w11972_,
		_w11973_,
		_w18921_
	);
	LUT3 #(
		.INIT('h80)
	) name8409 (
		\wishbone_bd_ram_mem1_reg[189][12]/P0001 ,
		_w11942_,
		_w11966_,
		_w18922_
	);
	LUT3 #(
		.INIT('h80)
	) name8410 (
		\wishbone_bd_ram_mem1_reg[145][12]/P0001 ,
		_w11959_,
		_w11977_,
		_w18923_
	);
	LUT4 #(
		.INIT('h0001)
	) name8411 (
		_w18920_,
		_w18921_,
		_w18922_,
		_w18923_,
		_w18924_
	);
	LUT3 #(
		.INIT('h80)
	) name8412 (
		\wishbone_bd_ram_mem1_reg[13][12]/P0001 ,
		_w11932_,
		_w11966_,
		_w18925_
	);
	LUT3 #(
		.INIT('h80)
	) name8413 (
		\wishbone_bd_ram_mem1_reg[83][12]/P0001 ,
		_w11938_,
		_w11972_,
		_w18926_
	);
	LUT3 #(
		.INIT('h80)
	) name8414 (
		\wishbone_bd_ram_mem1_reg[125][12]/P0001 ,
		_w11966_,
		_w12012_,
		_w18927_
	);
	LUT3 #(
		.INIT('h80)
	) name8415 (
		\wishbone_bd_ram_mem1_reg[22][12]/P0001 ,
		_w11935_,
		_w11986_,
		_w18928_
	);
	LUT4 #(
		.INIT('h0001)
	) name8416 (
		_w18925_,
		_w18926_,
		_w18927_,
		_w18928_,
		_w18929_
	);
	LUT3 #(
		.INIT('h80)
	) name8417 (
		\wishbone_bd_ram_mem1_reg[211][12]/P0001 ,
		_w11938_,
		_w11984_,
		_w18930_
	);
	LUT3 #(
		.INIT('h80)
	) name8418 (
		\wishbone_bd_ram_mem1_reg[194][12]/P0001 ,
		_w11945_,
		_w11963_,
		_w18931_
	);
	LUT3 #(
		.INIT('h80)
	) name8419 (
		\wishbone_bd_ram_mem1_reg[166][12]/P0001 ,
		_w11930_,
		_w11986_,
		_w18932_
	);
	LUT3 #(
		.INIT('h80)
	) name8420 (
		\wishbone_bd_ram_mem1_reg[208][12]/P0001 ,
		_w11941_,
		_w11984_,
		_w18933_
	);
	LUT4 #(
		.INIT('h0001)
	) name8421 (
		_w18930_,
		_w18931_,
		_w18932_,
		_w18933_,
		_w18934_
	);
	LUT4 #(
		.INIT('h8000)
	) name8422 (
		_w18919_,
		_w18924_,
		_w18929_,
		_w18934_,
		_w18935_
	);
	LUT3 #(
		.INIT('h80)
	) name8423 (
		\wishbone_bd_ram_mem1_reg[76][12]/P0001 ,
		_w11949_,
		_w11954_,
		_w18936_
	);
	LUT3 #(
		.INIT('h80)
	) name8424 (
		\wishbone_bd_ram_mem1_reg[233][12]/P0001 ,
		_w11968_,
		_w11982_,
		_w18937_
	);
	LUT3 #(
		.INIT('h80)
	) name8425 (
		\wishbone_bd_ram_mem1_reg[200][12]/P0001 ,
		_w11945_,
		_w11990_,
		_w18938_
	);
	LUT3 #(
		.INIT('h80)
	) name8426 (
		\wishbone_bd_ram_mem1_reg[242][12]/P0001 ,
		_w11952_,
		_w11963_,
		_w18939_
	);
	LUT4 #(
		.INIT('h0001)
	) name8427 (
		_w18936_,
		_w18937_,
		_w18938_,
		_w18939_,
		_w18940_
	);
	LUT3 #(
		.INIT('h80)
	) name8428 (
		\wishbone_bd_ram_mem1_reg[141][12]/P0001 ,
		_w11955_,
		_w11966_,
		_w18941_
	);
	LUT3 #(
		.INIT('h80)
	) name8429 (
		\wishbone_bd_ram_mem1_reg[169][12]/P0001 ,
		_w11930_,
		_w11968_,
		_w18942_
	);
	LUT3 #(
		.INIT('h80)
	) name8430 (
		\wishbone_bd_ram_mem1_reg[4][12]/P0001 ,
		_w11929_,
		_w11932_,
		_w18943_
	);
	LUT3 #(
		.INIT('h80)
	) name8431 (
		\wishbone_bd_ram_mem1_reg[78][12]/P0001 ,
		_w11948_,
		_w11949_,
		_w18944_
	);
	LUT4 #(
		.INIT('h0001)
	) name8432 (
		_w18941_,
		_w18942_,
		_w18943_,
		_w18944_,
		_w18945_
	);
	LUT3 #(
		.INIT('h80)
	) name8433 (
		\wishbone_bd_ram_mem1_reg[218][12]/P0001 ,
		_w11944_,
		_w11984_,
		_w18946_
	);
	LUT3 #(
		.INIT('h80)
	) name8434 (
		\wishbone_bd_ram_mem1_reg[57][12]/P0001 ,
		_w11968_,
		_w11979_,
		_w18947_
	);
	LUT3 #(
		.INIT('h80)
	) name8435 (
		\wishbone_bd_ram_mem1_reg[134][12]/P0001 ,
		_w11955_,
		_w11986_,
		_w18948_
	);
	LUT3 #(
		.INIT('h80)
	) name8436 (
		\wishbone_bd_ram_mem1_reg[183][12]/P0001 ,
		_w11942_,
		_w11975_,
		_w18949_
	);
	LUT4 #(
		.INIT('h0001)
	) name8437 (
		_w18946_,
		_w18947_,
		_w18948_,
		_w18949_,
		_w18950_
	);
	LUT3 #(
		.INIT('h80)
	) name8438 (
		\wishbone_bd_ram_mem1_reg[247][12]/P0001 ,
		_w11952_,
		_w11975_,
		_w18951_
	);
	LUT3 #(
		.INIT('h80)
	) name8439 (
		\wishbone_bd_ram_mem1_reg[240][12]/P0001 ,
		_w11941_,
		_w11952_,
		_w18952_
	);
	LUT3 #(
		.INIT('h80)
	) name8440 (
		\wishbone_bd_ram_mem1_reg[6][12]/P0001 ,
		_w11932_,
		_w11986_,
		_w18953_
	);
	LUT3 #(
		.INIT('h80)
	) name8441 (
		\wishbone_bd_ram_mem1_reg[81][12]/P0001 ,
		_w11972_,
		_w11977_,
		_w18954_
	);
	LUT4 #(
		.INIT('h0001)
	) name8442 (
		_w18951_,
		_w18952_,
		_w18953_,
		_w18954_,
		_w18955_
	);
	LUT4 #(
		.INIT('h8000)
	) name8443 (
		_w18940_,
		_w18945_,
		_w18950_,
		_w18955_,
		_w18956_
	);
	LUT3 #(
		.INIT('h80)
	) name8444 (
		\wishbone_bd_ram_mem1_reg[20][12]/P0001 ,
		_w11929_,
		_w11935_,
		_w18957_
	);
	LUT3 #(
		.INIT('h80)
	) name8445 (
		\wishbone_bd_ram_mem1_reg[123][12]/P0001 ,
		_w11936_,
		_w12012_,
		_w18958_
	);
	LUT3 #(
		.INIT('h80)
	) name8446 (
		\wishbone_bd_ram_mem1_reg[63][12]/P0001 ,
		_w11973_,
		_w11979_,
		_w18959_
	);
	LUT3 #(
		.INIT('h80)
	) name8447 (
		\wishbone_bd_ram_mem1_reg[196][12]/P0001 ,
		_w11929_,
		_w11945_,
		_w18960_
	);
	LUT4 #(
		.INIT('h0001)
	) name8448 (
		_w18957_,
		_w18958_,
		_w18959_,
		_w18960_,
		_w18961_
	);
	LUT3 #(
		.INIT('h80)
	) name8449 (
		\wishbone_bd_ram_mem1_reg[250][12]/P0001 ,
		_w11944_,
		_w11952_,
		_w18962_
	);
	LUT3 #(
		.INIT('h80)
	) name8450 (
		\wishbone_bd_ram_mem1_reg[23][12]/P0001 ,
		_w11935_,
		_w11975_,
		_w18963_
	);
	LUT3 #(
		.INIT('h80)
	) name8451 (
		\wishbone_bd_ram_mem1_reg[66][12]/P0001 ,
		_w11949_,
		_w11963_,
		_w18964_
	);
	LUT3 #(
		.INIT('h80)
	) name8452 (
		\wishbone_bd_ram_mem1_reg[116][12]/P0001 ,
		_w11929_,
		_w12012_,
		_w18965_
	);
	LUT4 #(
		.INIT('h0001)
	) name8453 (
		_w18962_,
		_w18963_,
		_w18964_,
		_w18965_,
		_w18966_
	);
	LUT3 #(
		.INIT('h80)
	) name8454 (
		\wishbone_bd_ram_mem1_reg[235][12]/P0001 ,
		_w11936_,
		_w11982_,
		_w18967_
	);
	LUT3 #(
		.INIT('h80)
	) name8455 (
		\wishbone_bd_ram_mem1_reg[124][12]/P0001 ,
		_w11954_,
		_w12012_,
		_w18968_
	);
	LUT3 #(
		.INIT('h80)
	) name8456 (
		\wishbone_bd_ram_mem1_reg[110][12]/P0001 ,
		_w11948_,
		_w11965_,
		_w18969_
	);
	LUT3 #(
		.INIT('h80)
	) name8457 (
		\wishbone_bd_ram_mem1_reg[181][12]/P0001 ,
		_w11933_,
		_w11942_,
		_w18970_
	);
	LUT4 #(
		.INIT('h0001)
	) name8458 (
		_w18967_,
		_w18968_,
		_w18969_,
		_w18970_,
		_w18971_
	);
	LUT3 #(
		.INIT('h80)
	) name8459 (
		\wishbone_bd_ram_mem1_reg[38][12]/P0001 ,
		_w11957_,
		_w11986_,
		_w18972_
	);
	LUT3 #(
		.INIT('h80)
	) name8460 (
		\wishbone_bd_ram_mem1_reg[202][12]/P0001 ,
		_w11944_,
		_w11945_,
		_w18973_
	);
	LUT3 #(
		.INIT('h80)
	) name8461 (
		\wishbone_bd_ram_mem1_reg[131][12]/P0001 ,
		_w11938_,
		_w11955_,
		_w18974_
	);
	LUT3 #(
		.INIT('h80)
	) name8462 (
		\wishbone_bd_ram_mem1_reg[29][12]/P0001 ,
		_w11935_,
		_w11966_,
		_w18975_
	);
	LUT4 #(
		.INIT('h0001)
	) name8463 (
		_w18972_,
		_w18973_,
		_w18974_,
		_w18975_,
		_w18976_
	);
	LUT4 #(
		.INIT('h8000)
	) name8464 (
		_w18961_,
		_w18966_,
		_w18971_,
		_w18976_,
		_w18977_
	);
	LUT4 #(
		.INIT('h8000)
	) name8465 (
		_w18914_,
		_w18935_,
		_w18956_,
		_w18977_,
		_w18978_
	);
	LUT3 #(
		.INIT('h80)
	) name8466 (
		\wishbone_bd_ram_mem1_reg[108][12]/P0001 ,
		_w11954_,
		_w11965_,
		_w18979_
	);
	LUT3 #(
		.INIT('h80)
	) name8467 (
		\wishbone_bd_ram_mem1_reg[69][12]/P0001 ,
		_w11933_,
		_w11949_,
		_w18980_
	);
	LUT3 #(
		.INIT('h80)
	) name8468 (
		\wishbone_bd_ram_mem1_reg[41][12]/P0001 ,
		_w11957_,
		_w11968_,
		_w18981_
	);
	LUT3 #(
		.INIT('h80)
	) name8469 (
		\wishbone_bd_ram_mem1_reg[207][12]/P0001 ,
		_w11945_,
		_w11973_,
		_w18982_
	);
	LUT4 #(
		.INIT('h0001)
	) name8470 (
		_w18979_,
		_w18980_,
		_w18981_,
		_w18982_,
		_w18983_
	);
	LUT3 #(
		.INIT('h80)
	) name8471 (
		\wishbone_bd_ram_mem1_reg[177][12]/P0001 ,
		_w11942_,
		_w11977_,
		_w18984_
	);
	LUT3 #(
		.INIT('h80)
	) name8472 (
		\wishbone_bd_ram_mem1_reg[89][12]/P0001 ,
		_w11968_,
		_w11972_,
		_w18985_
	);
	LUT3 #(
		.INIT('h80)
	) name8473 (
		\wishbone_bd_ram_mem1_reg[154][12]/P0001 ,
		_w11944_,
		_w11959_,
		_w18986_
	);
	LUT3 #(
		.INIT('h80)
	) name8474 (
		\wishbone_bd_ram_mem1_reg[101][12]/P0001 ,
		_w11933_,
		_w11965_,
		_w18987_
	);
	LUT4 #(
		.INIT('h0001)
	) name8475 (
		_w18984_,
		_w18985_,
		_w18986_,
		_w18987_,
		_w18988_
	);
	LUT3 #(
		.INIT('h80)
	) name8476 (
		\wishbone_bd_ram_mem1_reg[164][12]/P0001 ,
		_w11929_,
		_w11930_,
		_w18989_
	);
	LUT3 #(
		.INIT('h80)
	) name8477 (
		\wishbone_bd_ram_mem1_reg[149][12]/P0001 ,
		_w11933_,
		_w11959_,
		_w18990_
	);
	LUT3 #(
		.INIT('h80)
	) name8478 (
		\wishbone_bd_ram_mem1_reg[58][12]/P0001 ,
		_w11944_,
		_w11979_,
		_w18991_
	);
	LUT3 #(
		.INIT('h80)
	) name8479 (
		\wishbone_bd_ram_mem1_reg[162][12]/P0001 ,
		_w11930_,
		_w11963_,
		_w18992_
	);
	LUT4 #(
		.INIT('h0001)
	) name8480 (
		_w18989_,
		_w18990_,
		_w18991_,
		_w18992_,
		_w18993_
	);
	LUT3 #(
		.INIT('h80)
	) name8481 (
		\wishbone_bd_ram_mem1_reg[60][12]/P0001 ,
		_w11954_,
		_w11979_,
		_w18994_
	);
	LUT3 #(
		.INIT('h80)
	) name8482 (
		\wishbone_bd_ram_mem1_reg[18][12]/P0001 ,
		_w11935_,
		_w11963_,
		_w18995_
	);
	LUT3 #(
		.INIT('h80)
	) name8483 (
		\wishbone_bd_ram_mem1_reg[10][12]/P0001 ,
		_w11932_,
		_w11944_,
		_w18996_
	);
	LUT3 #(
		.INIT('h80)
	) name8484 (
		\wishbone_bd_ram_mem1_reg[206][12]/P0001 ,
		_w11945_,
		_w11948_,
		_w18997_
	);
	LUT4 #(
		.INIT('h0001)
	) name8485 (
		_w18994_,
		_w18995_,
		_w18996_,
		_w18997_,
		_w18998_
	);
	LUT4 #(
		.INIT('h8000)
	) name8486 (
		_w18983_,
		_w18988_,
		_w18993_,
		_w18998_,
		_w18999_
	);
	LUT3 #(
		.INIT('h80)
	) name8487 (
		\wishbone_bd_ram_mem1_reg[142][12]/P0001 ,
		_w11948_,
		_w11955_,
		_w19000_
	);
	LUT3 #(
		.INIT('h80)
	) name8488 (
		\wishbone_bd_ram_mem1_reg[204][12]/P0001 ,
		_w11945_,
		_w11954_,
		_w19001_
	);
	LUT3 #(
		.INIT('h80)
	) name8489 (
		\wishbone_bd_ram_mem1_reg[12][12]/P0001 ,
		_w11932_,
		_w11954_,
		_w19002_
	);
	LUT3 #(
		.INIT('h80)
	) name8490 (
		\wishbone_bd_ram_mem1_reg[143][12]/P0001 ,
		_w11955_,
		_w11973_,
		_w19003_
	);
	LUT4 #(
		.INIT('h0001)
	) name8491 (
		_w19000_,
		_w19001_,
		_w19002_,
		_w19003_,
		_w19004_
	);
	LUT3 #(
		.INIT('h80)
	) name8492 (
		\wishbone_bd_ram_mem1_reg[190][12]/P0001 ,
		_w11942_,
		_w11948_,
		_w19005_
	);
	LUT3 #(
		.INIT('h80)
	) name8493 (
		\wishbone_bd_ram_mem1_reg[198][12]/P0001 ,
		_w11945_,
		_w11986_,
		_w19006_
	);
	LUT3 #(
		.INIT('h80)
	) name8494 (
		\wishbone_bd_ram_mem1_reg[122][12]/P0001 ,
		_w11944_,
		_w12012_,
		_w19007_
	);
	LUT3 #(
		.INIT('h80)
	) name8495 (
		\wishbone_bd_ram_mem1_reg[92][12]/P0001 ,
		_w11954_,
		_w11972_,
		_w19008_
	);
	LUT4 #(
		.INIT('h0001)
	) name8496 (
		_w19005_,
		_w19006_,
		_w19007_,
		_w19008_,
		_w19009_
	);
	LUT3 #(
		.INIT('h80)
	) name8497 (
		\wishbone_bd_ram_mem1_reg[119][12]/P0001 ,
		_w11975_,
		_w12012_,
		_w19010_
	);
	LUT3 #(
		.INIT('h80)
	) name8498 (
		\wishbone_bd_ram_mem1_reg[64][12]/P0001 ,
		_w11941_,
		_w11949_,
		_w19011_
	);
	LUT3 #(
		.INIT('h80)
	) name8499 (
		\wishbone_bd_ram_mem1_reg[25][12]/P0001 ,
		_w11935_,
		_w11968_,
		_w19012_
	);
	LUT3 #(
		.INIT('h80)
	) name8500 (
		\wishbone_bd_ram_mem1_reg[188][12]/P0001 ,
		_w11942_,
		_w11954_,
		_w19013_
	);
	LUT4 #(
		.INIT('h0001)
	) name8501 (
		_w19010_,
		_w19011_,
		_w19012_,
		_w19013_,
		_w19014_
	);
	LUT3 #(
		.INIT('h80)
	) name8502 (
		\wishbone_bd_ram_mem1_reg[132][12]/P0001 ,
		_w11929_,
		_w11955_,
		_w19015_
	);
	LUT3 #(
		.INIT('h80)
	) name8503 (
		\wishbone_bd_ram_mem1_reg[167][12]/P0001 ,
		_w11930_,
		_w11975_,
		_w19016_
	);
	LUT3 #(
		.INIT('h80)
	) name8504 (
		\wishbone_bd_ram_mem1_reg[19][12]/P0001 ,
		_w11935_,
		_w11938_,
		_w19017_
	);
	LUT3 #(
		.INIT('h80)
	) name8505 (
		\wishbone_bd_ram_mem1_reg[115][12]/P0001 ,
		_w11938_,
		_w12012_,
		_w19018_
	);
	LUT4 #(
		.INIT('h0001)
	) name8506 (
		_w19015_,
		_w19016_,
		_w19017_,
		_w19018_,
		_w19019_
	);
	LUT4 #(
		.INIT('h8000)
	) name8507 (
		_w19004_,
		_w19009_,
		_w19014_,
		_w19019_,
		_w19020_
	);
	LUT3 #(
		.INIT('h80)
	) name8508 (
		\wishbone_bd_ram_mem1_reg[14][12]/P0001 ,
		_w11932_,
		_w11948_,
		_w19021_
	);
	LUT3 #(
		.INIT('h80)
	) name8509 (
		\wishbone_bd_ram_mem1_reg[163][12]/P0001 ,
		_w11930_,
		_w11938_,
		_w19022_
	);
	LUT3 #(
		.INIT('h80)
	) name8510 (
		\wishbone_bd_ram_mem1_reg[173][12]/P0001 ,
		_w11930_,
		_w11966_,
		_w19023_
	);
	LUT3 #(
		.INIT('h80)
	) name8511 (
		\wishbone_bd_ram_mem1_reg[192][12]/P0001 ,
		_w11941_,
		_w11945_,
		_w19024_
	);
	LUT4 #(
		.INIT('h0001)
	) name8512 (
		_w19021_,
		_w19022_,
		_w19023_,
		_w19024_,
		_w19025_
	);
	LUT3 #(
		.INIT('h80)
	) name8513 (
		\wishbone_bd_ram_mem1_reg[70][12]/P0001 ,
		_w11949_,
		_w11986_,
		_w19026_
	);
	LUT3 #(
		.INIT('h80)
	) name8514 (
		\wishbone_bd_ram_mem1_reg[148][12]/P0001 ,
		_w11929_,
		_w11959_,
		_w19027_
	);
	LUT3 #(
		.INIT('h80)
	) name8515 (
		\wishbone_bd_ram_mem1_reg[138][12]/P0001 ,
		_w11944_,
		_w11955_,
		_w19028_
	);
	LUT3 #(
		.INIT('h80)
	) name8516 (
		\wishbone_bd_ram_mem1_reg[109][12]/P0001 ,
		_w11965_,
		_w11966_,
		_w19029_
	);
	LUT4 #(
		.INIT('h0001)
	) name8517 (
		_w19026_,
		_w19027_,
		_w19028_,
		_w19029_,
		_w19030_
	);
	LUT3 #(
		.INIT('h80)
	) name8518 (
		\wishbone_bd_ram_mem1_reg[209][12]/P0001 ,
		_w11977_,
		_w11984_,
		_w19031_
	);
	LUT3 #(
		.INIT('h80)
	) name8519 (
		\wishbone_bd_ram_mem1_reg[176][12]/P0001 ,
		_w11941_,
		_w11942_,
		_w19032_
	);
	LUT3 #(
		.INIT('h80)
	) name8520 (
		\wishbone_bd_ram_mem1_reg[65][12]/P0001 ,
		_w11949_,
		_w11977_,
		_w19033_
	);
	LUT3 #(
		.INIT('h80)
	) name8521 (
		\wishbone_bd_ram_mem1_reg[151][12]/P0001 ,
		_w11959_,
		_w11975_,
		_w19034_
	);
	LUT4 #(
		.INIT('h0001)
	) name8522 (
		_w19031_,
		_w19032_,
		_w19033_,
		_w19034_,
		_w19035_
	);
	LUT3 #(
		.INIT('h80)
	) name8523 (
		\wishbone_bd_ram_mem1_reg[185][12]/P0001 ,
		_w11942_,
		_w11968_,
		_w19036_
	);
	LUT3 #(
		.INIT('h80)
	) name8524 (
		\wishbone_bd_ram_mem1_reg[36][12]/P0001 ,
		_w11929_,
		_w11957_,
		_w19037_
	);
	LUT3 #(
		.INIT('h80)
	) name8525 (
		\wishbone_bd_ram_mem1_reg[73][12]/P0001 ,
		_w11949_,
		_w11968_,
		_w19038_
	);
	LUT3 #(
		.INIT('h80)
	) name8526 (
		\wishbone_bd_ram_mem1_reg[136][12]/P0001 ,
		_w11955_,
		_w11990_,
		_w19039_
	);
	LUT4 #(
		.INIT('h0001)
	) name8527 (
		_w19036_,
		_w19037_,
		_w19038_,
		_w19039_,
		_w19040_
	);
	LUT4 #(
		.INIT('h8000)
	) name8528 (
		_w19025_,
		_w19030_,
		_w19035_,
		_w19040_,
		_w19041_
	);
	LUT3 #(
		.INIT('h80)
	) name8529 (
		\wishbone_bd_ram_mem1_reg[224][12]/P0001 ,
		_w11941_,
		_w11982_,
		_w19042_
	);
	LUT3 #(
		.INIT('h80)
	) name8530 (
		\wishbone_bd_ram_mem1_reg[182][12]/P0001 ,
		_w11942_,
		_w11986_,
		_w19043_
	);
	LUT3 #(
		.INIT('h80)
	) name8531 (
		\wishbone_bd_ram_mem1_reg[0][12]/P0001 ,
		_w11932_,
		_w11941_,
		_w19044_
	);
	LUT3 #(
		.INIT('h80)
	) name8532 (
		\wishbone_bd_ram_mem1_reg[32][12]/P0001 ,
		_w11941_,
		_w11957_,
		_w19045_
	);
	LUT4 #(
		.INIT('h0001)
	) name8533 (
		_w19042_,
		_w19043_,
		_w19044_,
		_w19045_,
		_w19046_
	);
	LUT3 #(
		.INIT('h80)
	) name8534 (
		\wishbone_bd_ram_mem1_reg[56][12]/P0001 ,
		_w11979_,
		_w11990_,
		_w19047_
	);
	LUT3 #(
		.INIT('h80)
	) name8535 (
		\wishbone_bd_ram_mem1_reg[179][12]/P0001 ,
		_w11938_,
		_w11942_,
		_w19048_
	);
	LUT3 #(
		.INIT('h80)
	) name8536 (
		\wishbone_bd_ram_mem1_reg[255][12]/P0001 ,
		_w11952_,
		_w11973_,
		_w19049_
	);
	LUT3 #(
		.INIT('h80)
	) name8537 (
		\wishbone_bd_ram_mem1_reg[37][12]/P0001 ,
		_w11933_,
		_w11957_,
		_w19050_
	);
	LUT4 #(
		.INIT('h0001)
	) name8538 (
		_w19047_,
		_w19048_,
		_w19049_,
		_w19050_,
		_w19051_
	);
	LUT3 #(
		.INIT('h80)
	) name8539 (
		\wishbone_bd_ram_mem1_reg[45][12]/P0001 ,
		_w11957_,
		_w11966_,
		_w19052_
	);
	LUT3 #(
		.INIT('h80)
	) name8540 (
		\wishbone_bd_ram_mem1_reg[170][12]/P0001 ,
		_w11930_,
		_w11944_,
		_w19053_
	);
	LUT3 #(
		.INIT('h80)
	) name8541 (
		\wishbone_bd_ram_mem1_reg[94][12]/P0001 ,
		_w11948_,
		_w11972_,
		_w19054_
	);
	LUT3 #(
		.INIT('h80)
	) name8542 (
		\wishbone_bd_ram_mem1_reg[74][12]/P0001 ,
		_w11944_,
		_w11949_,
		_w19055_
	);
	LUT4 #(
		.INIT('h0001)
	) name8543 (
		_w19052_,
		_w19053_,
		_w19054_,
		_w19055_,
		_w19056_
	);
	LUT3 #(
		.INIT('h80)
	) name8544 (
		\wishbone_bd_ram_mem1_reg[178][12]/P0001 ,
		_w11942_,
		_w11963_,
		_w19057_
	);
	LUT3 #(
		.INIT('h80)
	) name8545 (
		\wishbone_bd_ram_mem1_reg[30][12]/P0001 ,
		_w11935_,
		_w11948_,
		_w19058_
	);
	LUT3 #(
		.INIT('h80)
	) name8546 (
		\wishbone_bd_ram_mem1_reg[171][12]/P0001 ,
		_w11930_,
		_w11936_,
		_w19059_
	);
	LUT3 #(
		.INIT('h80)
	) name8547 (
		\wishbone_bd_ram_mem1_reg[160][12]/P0001 ,
		_w11930_,
		_w11941_,
		_w19060_
	);
	LUT4 #(
		.INIT('h0001)
	) name8548 (
		_w19057_,
		_w19058_,
		_w19059_,
		_w19060_,
		_w19061_
	);
	LUT4 #(
		.INIT('h8000)
	) name8549 (
		_w19046_,
		_w19051_,
		_w19056_,
		_w19061_,
		_w19062_
	);
	LUT4 #(
		.INIT('h8000)
	) name8550 (
		_w18999_,
		_w19020_,
		_w19041_,
		_w19062_,
		_w19063_
	);
	LUT3 #(
		.INIT('h80)
	) name8551 (
		\wishbone_bd_ram_mem1_reg[98][12]/P0001 ,
		_w11963_,
		_w11965_,
		_w19064_
	);
	LUT3 #(
		.INIT('h80)
	) name8552 (
		\wishbone_bd_ram_mem1_reg[130][12]/P0001 ,
		_w11955_,
		_w11963_,
		_w19065_
	);
	LUT3 #(
		.INIT('h80)
	) name8553 (
		\wishbone_bd_ram_mem1_reg[100][12]/P0001 ,
		_w11929_,
		_w11965_,
		_w19066_
	);
	LUT3 #(
		.INIT('h80)
	) name8554 (
		\wishbone_bd_ram_mem1_reg[99][12]/P0001 ,
		_w11938_,
		_w11965_,
		_w19067_
	);
	LUT4 #(
		.INIT('h0001)
	) name8555 (
		_w19064_,
		_w19065_,
		_w19066_,
		_w19067_,
		_w19068_
	);
	LUT3 #(
		.INIT('h80)
	) name8556 (
		\wishbone_bd_ram_mem1_reg[3][12]/P0001 ,
		_w11932_,
		_w11938_,
		_w19069_
	);
	LUT3 #(
		.INIT('h80)
	) name8557 (
		\wishbone_bd_ram_mem1_reg[159][12]/P0001 ,
		_w11959_,
		_w11973_,
		_w19070_
	);
	LUT3 #(
		.INIT('h80)
	) name8558 (
		\wishbone_bd_ram_mem1_reg[156][12]/P0001 ,
		_w11954_,
		_w11959_,
		_w19071_
	);
	LUT3 #(
		.INIT('h80)
	) name8559 (
		\wishbone_bd_ram_mem1_reg[251][12]/P0001 ,
		_w11936_,
		_w11952_,
		_w19072_
	);
	LUT4 #(
		.INIT('h0001)
	) name8560 (
		_w19069_,
		_w19070_,
		_w19071_,
		_w19072_,
		_w19073_
	);
	LUT3 #(
		.INIT('h80)
	) name8561 (
		\wishbone_bd_ram_mem1_reg[172][12]/P0001 ,
		_w11930_,
		_w11954_,
		_w19074_
	);
	LUT3 #(
		.INIT('h80)
	) name8562 (
		\wishbone_bd_ram_mem1_reg[213][12]/P0001 ,
		_w11933_,
		_w11984_,
		_w19075_
	);
	LUT3 #(
		.INIT('h80)
	) name8563 (
		\wishbone_bd_ram_mem1_reg[150][12]/P0001 ,
		_w11959_,
		_w11986_,
		_w19076_
	);
	LUT3 #(
		.INIT('h80)
	) name8564 (
		\wishbone_bd_ram_mem1_reg[157][12]/P0001 ,
		_w11959_,
		_w11966_,
		_w19077_
	);
	LUT4 #(
		.INIT('h0001)
	) name8565 (
		_w19074_,
		_w19075_,
		_w19076_,
		_w19077_,
		_w19078_
	);
	LUT3 #(
		.INIT('h80)
	) name8566 (
		\wishbone_bd_ram_mem1_reg[71][12]/P0001 ,
		_w11949_,
		_w11975_,
		_w19079_
	);
	LUT3 #(
		.INIT('h80)
	) name8567 (
		\wishbone_bd_ram_mem1_reg[2][12]/P0001 ,
		_w11932_,
		_w11963_,
		_w19080_
	);
	LUT3 #(
		.INIT('h80)
	) name8568 (
		\wishbone_bd_ram_mem1_reg[168][12]/P0001 ,
		_w11930_,
		_w11990_,
		_w19081_
	);
	LUT3 #(
		.INIT('h80)
	) name8569 (
		\wishbone_bd_ram_mem1_reg[203][12]/P0001 ,
		_w11936_,
		_w11945_,
		_w19082_
	);
	LUT4 #(
		.INIT('h0001)
	) name8570 (
		_w19079_,
		_w19080_,
		_w19081_,
		_w19082_,
		_w19083_
	);
	LUT4 #(
		.INIT('h8000)
	) name8571 (
		_w19068_,
		_w19073_,
		_w19078_,
		_w19083_,
		_w19084_
	);
	LUT3 #(
		.INIT('h80)
	) name8572 (
		\wishbone_bd_ram_mem1_reg[80][12]/P0001 ,
		_w11941_,
		_w11972_,
		_w19085_
	);
	LUT3 #(
		.INIT('h80)
	) name8573 (
		\wishbone_bd_ram_mem1_reg[91][12]/P0001 ,
		_w11936_,
		_w11972_,
		_w19086_
	);
	LUT3 #(
		.INIT('h80)
	) name8574 (
		\wishbone_bd_ram_mem1_reg[102][12]/P0001 ,
		_w11965_,
		_w11986_,
		_w19087_
	);
	LUT3 #(
		.INIT('h80)
	) name8575 (
		\wishbone_bd_ram_mem1_reg[67][12]/P0001 ,
		_w11938_,
		_w11949_,
		_w19088_
	);
	LUT4 #(
		.INIT('h0001)
	) name8576 (
		_w19085_,
		_w19086_,
		_w19087_,
		_w19088_,
		_w19089_
	);
	LUT3 #(
		.INIT('h80)
	) name8577 (
		\wishbone_bd_ram_mem1_reg[72][12]/P0001 ,
		_w11949_,
		_w11990_,
		_w19090_
	);
	LUT3 #(
		.INIT('h80)
	) name8578 (
		\wishbone_bd_ram_mem1_reg[184][12]/P0001 ,
		_w11942_,
		_w11990_,
		_w19091_
	);
	LUT3 #(
		.INIT('h80)
	) name8579 (
		\wishbone_bd_ram_mem1_reg[11][12]/P0001 ,
		_w11932_,
		_w11936_,
		_w19092_
	);
	LUT3 #(
		.INIT('h80)
	) name8580 (
		\wishbone_bd_ram_mem1_reg[214][12]/P0001 ,
		_w11984_,
		_w11986_,
		_w19093_
	);
	LUT4 #(
		.INIT('h0001)
	) name8581 (
		_w19090_,
		_w19091_,
		_w19092_,
		_w19093_,
		_w19094_
	);
	LUT3 #(
		.INIT('h80)
	) name8582 (
		\wishbone_bd_ram_mem1_reg[133][12]/P0001 ,
		_w11933_,
		_w11955_,
		_w19095_
	);
	LUT3 #(
		.INIT('h80)
	) name8583 (
		\wishbone_bd_ram_mem1_reg[221][12]/P0001 ,
		_w11966_,
		_w11984_,
		_w19096_
	);
	LUT3 #(
		.INIT('h80)
	) name8584 (
		\wishbone_bd_ram_mem1_reg[226][12]/P0001 ,
		_w11963_,
		_w11982_,
		_w19097_
	);
	LUT3 #(
		.INIT('h80)
	) name8585 (
		\wishbone_bd_ram_mem1_reg[88][12]/P0001 ,
		_w11972_,
		_w11990_,
		_w19098_
	);
	LUT4 #(
		.INIT('h0001)
	) name8586 (
		_w19095_,
		_w19096_,
		_w19097_,
		_w19098_,
		_w19099_
	);
	LUT3 #(
		.INIT('h80)
	) name8587 (
		\wishbone_bd_ram_mem1_reg[50][12]/P0001 ,
		_w11963_,
		_w11979_,
		_w19100_
	);
	LUT3 #(
		.INIT('h80)
	) name8588 (
		\wishbone_bd_ram_mem1_reg[61][12]/P0001 ,
		_w11966_,
		_w11979_,
		_w19101_
	);
	LUT3 #(
		.INIT('h80)
	) name8589 (
		\wishbone_bd_ram_mem1_reg[53][12]/P0001 ,
		_w11933_,
		_w11979_,
		_w19102_
	);
	LUT3 #(
		.INIT('h80)
	) name8590 (
		\wishbone_bd_ram_mem1_reg[246][12]/P0001 ,
		_w11952_,
		_w11986_,
		_w19103_
	);
	LUT4 #(
		.INIT('h0001)
	) name8591 (
		_w19100_,
		_w19101_,
		_w19102_,
		_w19103_,
		_w19104_
	);
	LUT4 #(
		.INIT('h8000)
	) name8592 (
		_w19089_,
		_w19094_,
		_w19099_,
		_w19104_,
		_w19105_
	);
	LUT3 #(
		.INIT('h80)
	) name8593 (
		\wishbone_bd_ram_mem1_reg[34][12]/P0001 ,
		_w11957_,
		_w11963_,
		_w19106_
	);
	LUT3 #(
		.INIT('h80)
	) name8594 (
		\wishbone_bd_ram_mem1_reg[21][12]/P0001 ,
		_w11933_,
		_w11935_,
		_w19107_
	);
	LUT3 #(
		.INIT('h80)
	) name8595 (
		\wishbone_bd_ram_mem1_reg[140][12]/P0001 ,
		_w11954_,
		_w11955_,
		_w19108_
	);
	LUT3 #(
		.INIT('h80)
	) name8596 (
		\wishbone_bd_ram_mem1_reg[75][12]/P0001 ,
		_w11936_,
		_w11949_,
		_w19109_
	);
	LUT4 #(
		.INIT('h0001)
	) name8597 (
		_w19106_,
		_w19107_,
		_w19108_,
		_w19109_,
		_w19110_
	);
	LUT3 #(
		.INIT('h80)
	) name8598 (
		\wishbone_bd_ram_mem1_reg[39][12]/P0001 ,
		_w11957_,
		_w11975_,
		_w19111_
	);
	LUT3 #(
		.INIT('h80)
	) name8599 (
		\wishbone_bd_ram_mem1_reg[152][12]/P0001 ,
		_w11959_,
		_w11990_,
		_w19112_
	);
	LUT3 #(
		.INIT('h80)
	) name8600 (
		\wishbone_bd_ram_mem1_reg[195][12]/P0001 ,
		_w11938_,
		_w11945_,
		_w19113_
	);
	LUT3 #(
		.INIT('h80)
	) name8601 (
		\wishbone_bd_ram_mem1_reg[113][12]/P0001 ,
		_w11977_,
		_w12012_,
		_w19114_
	);
	LUT4 #(
		.INIT('h0001)
	) name8602 (
		_w19111_,
		_w19112_,
		_w19113_,
		_w19114_,
		_w19115_
	);
	LUT3 #(
		.INIT('h80)
	) name8603 (
		\wishbone_bd_ram_mem1_reg[68][12]/P0001 ,
		_w11929_,
		_w11949_,
		_w19116_
	);
	LUT3 #(
		.INIT('h80)
	) name8604 (
		\wishbone_bd_ram_mem1_reg[15][12]/P0001 ,
		_w11932_,
		_w11973_,
		_w19117_
	);
	LUT3 #(
		.INIT('h80)
	) name8605 (
		\wishbone_bd_ram_mem1_reg[42][12]/P0001 ,
		_w11944_,
		_w11957_,
		_w19118_
	);
	LUT3 #(
		.INIT('h80)
	) name8606 (
		\wishbone_bd_ram_mem1_reg[46][12]/P0001 ,
		_w11948_,
		_w11957_,
		_w19119_
	);
	LUT4 #(
		.INIT('h0001)
	) name8607 (
		_w19116_,
		_w19117_,
		_w19118_,
		_w19119_,
		_w19120_
	);
	LUT3 #(
		.INIT('h80)
	) name8608 (
		\wishbone_bd_ram_mem1_reg[137][12]/P0001 ,
		_w11955_,
		_w11968_,
		_w19121_
	);
	LUT3 #(
		.INIT('h80)
	) name8609 (
		\wishbone_bd_ram_mem1_reg[197][12]/P0001 ,
		_w11933_,
		_w11945_,
		_w19122_
	);
	LUT3 #(
		.INIT('h80)
	) name8610 (
		\wishbone_bd_ram_mem1_reg[253][12]/P0001 ,
		_w11952_,
		_w11966_,
		_w19123_
	);
	LUT3 #(
		.INIT('h80)
	) name8611 (
		\wishbone_bd_ram_mem1_reg[44][12]/P0001 ,
		_w11954_,
		_w11957_,
		_w19124_
	);
	LUT4 #(
		.INIT('h0001)
	) name8612 (
		_w19121_,
		_w19122_,
		_w19123_,
		_w19124_,
		_w19125_
	);
	LUT4 #(
		.INIT('h8000)
	) name8613 (
		_w19110_,
		_w19115_,
		_w19120_,
		_w19125_,
		_w19126_
	);
	LUT3 #(
		.INIT('h80)
	) name8614 (
		\wishbone_bd_ram_mem1_reg[9][12]/P0001 ,
		_w11932_,
		_w11968_,
		_w19127_
	);
	LUT3 #(
		.INIT('h80)
	) name8615 (
		\wishbone_bd_ram_mem1_reg[228][12]/P0001 ,
		_w11929_,
		_w11982_,
		_w19128_
	);
	LUT3 #(
		.INIT('h80)
	) name8616 (
		\wishbone_bd_ram_mem1_reg[79][12]/P0001 ,
		_w11949_,
		_w11973_,
		_w19129_
	);
	LUT3 #(
		.INIT('h80)
	) name8617 (
		\wishbone_bd_ram_mem1_reg[40][12]/P0001 ,
		_w11957_,
		_w11990_,
		_w19130_
	);
	LUT4 #(
		.INIT('h0001)
	) name8618 (
		_w19127_,
		_w19128_,
		_w19129_,
		_w19130_,
		_w19131_
	);
	LUT3 #(
		.INIT('h80)
	) name8619 (
		\wishbone_bd_ram_mem1_reg[87][12]/P0001 ,
		_w11972_,
		_w11975_,
		_w19132_
	);
	LUT3 #(
		.INIT('h80)
	) name8620 (
		\wishbone_bd_ram_mem1_reg[84][12]/P0001 ,
		_w11929_,
		_w11972_,
		_w19133_
	);
	LUT3 #(
		.INIT('h80)
	) name8621 (
		\wishbone_bd_ram_mem1_reg[186][12]/P0001 ,
		_w11942_,
		_w11944_,
		_w19134_
	);
	LUT3 #(
		.INIT('h80)
	) name8622 (
		\wishbone_bd_ram_mem1_reg[114][12]/P0001 ,
		_w11963_,
		_w12012_,
		_w19135_
	);
	LUT4 #(
		.INIT('h0001)
	) name8623 (
		_w19132_,
		_w19133_,
		_w19134_,
		_w19135_,
		_w19136_
	);
	LUT3 #(
		.INIT('h80)
	) name8624 (
		\wishbone_bd_ram_mem1_reg[51][12]/P0001 ,
		_w11938_,
		_w11979_,
		_w19137_
	);
	LUT3 #(
		.INIT('h80)
	) name8625 (
		\wishbone_bd_ram_mem1_reg[93][12]/P0001 ,
		_w11966_,
		_w11972_,
		_w19138_
	);
	LUT3 #(
		.INIT('h80)
	) name8626 (
		\wishbone_bd_ram_mem1_reg[254][12]/P0001 ,
		_w11948_,
		_w11952_,
		_w19139_
	);
	LUT3 #(
		.INIT('h80)
	) name8627 (
		\wishbone_bd_ram_mem1_reg[222][12]/P0001 ,
		_w11948_,
		_w11984_,
		_w19140_
	);
	LUT4 #(
		.INIT('h0001)
	) name8628 (
		_w19137_,
		_w19138_,
		_w19139_,
		_w19140_,
		_w19141_
	);
	LUT3 #(
		.INIT('h80)
	) name8629 (
		\wishbone_bd_ram_mem1_reg[48][12]/P0001 ,
		_w11941_,
		_w11979_,
		_w19142_
	);
	LUT3 #(
		.INIT('h80)
	) name8630 (
		\wishbone_bd_ram_mem1_reg[237][12]/P0001 ,
		_w11966_,
		_w11982_,
		_w19143_
	);
	LUT3 #(
		.INIT('h80)
	) name8631 (
		\wishbone_bd_ram_mem1_reg[107][12]/P0001 ,
		_w11936_,
		_w11965_,
		_w19144_
	);
	LUT3 #(
		.INIT('h80)
	) name8632 (
		\wishbone_bd_ram_mem1_reg[16][12]/P0001 ,
		_w11935_,
		_w11941_,
		_w19145_
	);
	LUT4 #(
		.INIT('h0001)
	) name8633 (
		_w19142_,
		_w19143_,
		_w19144_,
		_w19145_,
		_w19146_
	);
	LUT4 #(
		.INIT('h8000)
	) name8634 (
		_w19131_,
		_w19136_,
		_w19141_,
		_w19146_,
		_w19147_
	);
	LUT4 #(
		.INIT('h8000)
	) name8635 (
		_w19084_,
		_w19105_,
		_w19126_,
		_w19147_,
		_w19148_
	);
	LUT4 #(
		.INIT('h8000)
	) name8636 (
		_w18893_,
		_w18978_,
		_w19063_,
		_w19148_,
		_w19149_
	);
	LUT4 #(
		.INIT('h1555)
	) name8637 (
		wb_rst_i_pad,
		_w18792_,
		_w18797_,
		_w18807_,
		_w19150_
	);
	LUT3 #(
		.INIT('hba)
	) name8638 (
		_w18808_,
		_w19149_,
		_w19150_,
		_w19151_
	);
	LUT3 #(
		.INIT('h70)
	) name8639 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_TxLength_reg[3]/NET0131 ,
		_w19152_
	);
	LUT2 #(
		.INIT('h4)
	) name8640 (
		_w12302_,
		_w19152_,
		_w19153_
	);
	LUT4 #(
		.INIT('hfe00)
	) name8641 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		\wishbone_TxLength_reg[2]/NET0131 ,
		\wishbone_TxLength_reg[3]/NET0131 ,
		_w19154_
	);
	LUT4 #(
		.INIT('haaa2)
	) name8642 (
		_w12304_,
		_w14519_,
		_w14521_,
		_w19154_,
		_w19155_
	);
	LUT3 #(
		.INIT('h70)
	) name8643 (
		_w12312_,
		_w12317_,
		_w19155_,
		_w19156_
	);
	LUT2 #(
		.INIT('h1)
	) name8644 (
		\wishbone_TxLength_reg[1]/NET0131 ,
		\wishbone_TxLength_reg[2]/NET0131 ,
		_w19157_
	);
	LUT4 #(
		.INIT('h0013)
	) name8645 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[2]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w19158_
	);
	LUT4 #(
		.INIT('hddde)
	) name8646 (
		\wishbone_TxLength_reg[3]/NET0131 ,
		_w14519_,
		_w19157_,
		_w19158_,
		_w19159_
	);
	LUT2 #(
		.INIT('h4)
	) name8647 (
		_w12302_,
		_w19159_,
		_w19160_
	);
	LUT3 #(
		.INIT('h15)
	) name8648 (
		_w19153_,
		_w19156_,
		_w19160_,
		_w19161_
	);
	LUT3 #(
		.INIT('h2f)
	) name8649 (
		_w12303_,
		_w17713_,
		_w19161_,
		_w19162_
	);
	LUT3 #(
		.INIT('h70)
	) name8650 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_TxLength_reg[6]/NET0131 ,
		_w19163_
	);
	LUT4 #(
		.INIT('hd111)
	) name8651 (
		\wishbone_TxLength_reg[6]/NET0131 ,
		_w12304_,
		_w12312_,
		_w12317_,
		_w19164_
	);
	LUT4 #(
		.INIT('h0001)
	) name8652 (
		\wishbone_TxLength_reg[2]/NET0131 ,
		\wishbone_TxLength_reg[3]/NET0131 ,
		\wishbone_TxLength_reg[4]/NET0131 ,
		\wishbone_TxLength_reg[5]/NET0131 ,
		_w19165_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name8653 (
		\wishbone_TxLength_reg[4]/NET0131 ,
		\wishbone_TxLength_reg[5]/NET0131 ,
		\wishbone_TxLength_reg[6]/NET0131 ,
		_w12308_,
		_w19166_
	);
	LUT3 #(
		.INIT('h08)
	) name8654 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		\wishbone_TxLength_reg[6]/NET0131 ,
		_w19167_
	);
	LUT2 #(
		.INIT('h2)
	) name8655 (
		_w14517_,
		_w19167_,
		_w19168_
	);
	LUT4 #(
		.INIT('h50f3)
	) name8656 (
		_w14516_,
		_w14524_,
		_w19166_,
		_w19168_,
		_w19169_
	);
	LUT3 #(
		.INIT('h10)
	) name8657 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[5]/NET0131 ,
		\wishbone_TxLength_reg[6]/NET0131 ,
		_w19170_
	);
	LUT2 #(
		.INIT('h8)
	) name8658 (
		_w14527_,
		_w19170_,
		_w19171_
	);
	LUT3 #(
		.INIT('h80)
	) name8659 (
		\wishbone_TxLength_reg[6]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w19172_
	);
	LUT4 #(
		.INIT('h1000)
	) name8660 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w19173_
	);
	LUT3 #(
		.INIT('h13)
	) name8661 (
		_w19165_,
		_w19172_,
		_w19173_,
		_w19174_
	);
	LUT4 #(
		.INIT('h90c0)
	) name8662 (
		\wishbone_TxLength_reg[5]/NET0131 ,
		\wishbone_TxLength_reg[6]/NET0131 ,
		_w14526_,
		_w14527_,
		_w19175_
	);
	LUT4 #(
		.INIT('h0054)
	) name8663 (
		_w19163_,
		_w19171_,
		_w19174_,
		_w19175_,
		_w19176_
	);
	LUT4 #(
		.INIT('h0111)
	) name8664 (
		_w12302_,
		_w19164_,
		_w19169_,
		_w19176_,
		_w19177_
	);
	LUT3 #(
		.INIT('hf2)
	) name8665 (
		_w12303_,
		_w18746_,
		_w19177_,
		_w19178_
	);
	LUT4 #(
		.INIT('h70f0)
	) name8666 (
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w19179_
	);
	LUT4 #(
		.INIT('h4000)
	) name8667 (
		wb_rst_i_pad,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w19180_
	);
	LUT3 #(
		.INIT('hdc)
	) name8668 (
		_w14151_,
		_w19179_,
		_w19180_,
		_w19181_
	);
	LUT3 #(
		.INIT('h70)
	) name8669 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		_w19182_
	);
	LUT2 #(
		.INIT('h4)
	) name8670 (
		_w15303_,
		_w19182_,
		_w19183_
	);
	LUT3 #(
		.INIT('h80)
	) name8671 (
		\wishbone_bd_ram_mem0_reg[153][0]/P0001 ,
		_w11959_,
		_w11968_,
		_w19184_
	);
	LUT3 #(
		.INIT('h80)
	) name8672 (
		\wishbone_bd_ram_mem0_reg[174][0]/P0001 ,
		_w11930_,
		_w11948_,
		_w19185_
	);
	LUT3 #(
		.INIT('h80)
	) name8673 (
		\wishbone_bd_ram_mem0_reg[166][0]/P0001 ,
		_w11930_,
		_w11986_,
		_w19186_
	);
	LUT3 #(
		.INIT('h80)
	) name8674 (
		\wishbone_bd_ram_mem0_reg[150][0]/P0001 ,
		_w11959_,
		_w11986_,
		_w19187_
	);
	LUT4 #(
		.INIT('h0001)
	) name8675 (
		_w19184_,
		_w19185_,
		_w19186_,
		_w19187_,
		_w19188_
	);
	LUT3 #(
		.INIT('h80)
	) name8676 (
		\wishbone_bd_ram_mem0_reg[159][0]/P0001 ,
		_w11959_,
		_w11973_,
		_w19189_
	);
	LUT3 #(
		.INIT('h80)
	) name8677 (
		\wishbone_bd_ram_mem0_reg[25][0]/P0001 ,
		_w11935_,
		_w11968_,
		_w19190_
	);
	LUT3 #(
		.INIT('h80)
	) name8678 (
		\wishbone_bd_ram_mem0_reg[26][0]/P0001 ,
		_w11935_,
		_w11944_,
		_w19191_
	);
	LUT3 #(
		.INIT('h80)
	) name8679 (
		\wishbone_bd_ram_mem0_reg[146][0]/P0001 ,
		_w11959_,
		_w11963_,
		_w19192_
	);
	LUT4 #(
		.INIT('h0001)
	) name8680 (
		_w19189_,
		_w19190_,
		_w19191_,
		_w19192_,
		_w19193_
	);
	LUT3 #(
		.INIT('h80)
	) name8681 (
		\wishbone_bd_ram_mem0_reg[14][0]/P0001 ,
		_w11932_,
		_w11948_,
		_w19194_
	);
	LUT3 #(
		.INIT('h80)
	) name8682 (
		\wishbone_bd_ram_mem0_reg[189][0]/P0001 ,
		_w11942_,
		_w11966_,
		_w19195_
	);
	LUT3 #(
		.INIT('h80)
	) name8683 (
		\wishbone_bd_ram_mem0_reg[3][0]/P0001 ,
		_w11932_,
		_w11938_,
		_w19196_
	);
	LUT3 #(
		.INIT('h80)
	) name8684 (
		\wishbone_bd_ram_mem0_reg[194][0]/P0001 ,
		_w11945_,
		_w11963_,
		_w19197_
	);
	LUT4 #(
		.INIT('h0001)
	) name8685 (
		_w19194_,
		_w19195_,
		_w19196_,
		_w19197_,
		_w19198_
	);
	LUT3 #(
		.INIT('h80)
	) name8686 (
		\wishbone_bd_ram_mem0_reg[101][0]/P0001 ,
		_w11933_,
		_w11965_,
		_w19199_
	);
	LUT3 #(
		.INIT('h80)
	) name8687 (
		\wishbone_bd_ram_mem0_reg[238][0]/P0001 ,
		_w11948_,
		_w11982_,
		_w19200_
	);
	LUT3 #(
		.INIT('h80)
	) name8688 (
		\wishbone_bd_ram_mem0_reg[115][0]/P0001 ,
		_w11938_,
		_w12012_,
		_w19201_
	);
	LUT3 #(
		.INIT('h80)
	) name8689 (
		\wishbone_bd_ram_mem0_reg[164][0]/P0001 ,
		_w11929_,
		_w11930_,
		_w19202_
	);
	LUT4 #(
		.INIT('h0001)
	) name8690 (
		_w19199_,
		_w19200_,
		_w19201_,
		_w19202_,
		_w19203_
	);
	LUT4 #(
		.INIT('h8000)
	) name8691 (
		_w19188_,
		_w19193_,
		_w19198_,
		_w19203_,
		_w19204_
	);
	LUT3 #(
		.INIT('h80)
	) name8692 (
		\wishbone_bd_ram_mem0_reg[114][0]/P0001 ,
		_w11963_,
		_w12012_,
		_w19205_
	);
	LUT3 #(
		.INIT('h80)
	) name8693 (
		\wishbone_bd_ram_mem0_reg[79][0]/P0001 ,
		_w11949_,
		_w11973_,
		_w19206_
	);
	LUT3 #(
		.INIT('h80)
	) name8694 (
		\wishbone_bd_ram_mem0_reg[151][0]/P0001 ,
		_w11959_,
		_w11975_,
		_w19207_
	);
	LUT3 #(
		.INIT('h80)
	) name8695 (
		\wishbone_bd_ram_mem0_reg[112][0]/P0001 ,
		_w11941_,
		_w12012_,
		_w19208_
	);
	LUT4 #(
		.INIT('h0001)
	) name8696 (
		_w19205_,
		_w19206_,
		_w19207_,
		_w19208_,
		_w19209_
	);
	LUT3 #(
		.INIT('h80)
	) name8697 (
		\wishbone_bd_ram_mem0_reg[228][0]/P0001 ,
		_w11929_,
		_w11982_,
		_w19210_
	);
	LUT3 #(
		.INIT('h80)
	) name8698 (
		\wishbone_bd_ram_mem0_reg[0][0]/P0001 ,
		_w11932_,
		_w11941_,
		_w19211_
	);
	LUT3 #(
		.INIT('h80)
	) name8699 (
		\wishbone_bd_ram_mem0_reg[184][0]/P0001 ,
		_w11942_,
		_w11990_,
		_w19212_
	);
	LUT3 #(
		.INIT('h80)
	) name8700 (
		\wishbone_bd_ram_mem0_reg[30][0]/P0001 ,
		_w11935_,
		_w11948_,
		_w19213_
	);
	LUT4 #(
		.INIT('h0001)
	) name8701 (
		_w19210_,
		_w19211_,
		_w19212_,
		_w19213_,
		_w19214_
	);
	LUT3 #(
		.INIT('h80)
	) name8702 (
		\wishbone_bd_ram_mem0_reg[103][0]/P0001 ,
		_w11965_,
		_w11975_,
		_w19215_
	);
	LUT3 #(
		.INIT('h80)
	) name8703 (
		\wishbone_bd_ram_mem0_reg[7][0]/P0001 ,
		_w11932_,
		_w11975_,
		_w19216_
	);
	LUT3 #(
		.INIT('h80)
	) name8704 (
		\wishbone_bd_ram_mem0_reg[45][0]/P0001 ,
		_w11957_,
		_w11966_,
		_w19217_
	);
	LUT3 #(
		.INIT('h80)
	) name8705 (
		\wishbone_bd_ram_mem0_reg[39][0]/P0001 ,
		_w11957_,
		_w11975_,
		_w19218_
	);
	LUT4 #(
		.INIT('h0001)
	) name8706 (
		_w19215_,
		_w19216_,
		_w19217_,
		_w19218_,
		_w19219_
	);
	LUT3 #(
		.INIT('h80)
	) name8707 (
		\wishbone_bd_ram_mem0_reg[126][0]/P0001 ,
		_w11948_,
		_w12012_,
		_w19220_
	);
	LUT3 #(
		.INIT('h80)
	) name8708 (
		\wishbone_bd_ram_mem0_reg[47][0]/P0001 ,
		_w11957_,
		_w11973_,
		_w19221_
	);
	LUT3 #(
		.INIT('h80)
	) name8709 (
		\wishbone_bd_ram_mem0_reg[58][0]/P0001 ,
		_w11944_,
		_w11979_,
		_w19222_
	);
	LUT3 #(
		.INIT('h80)
	) name8710 (
		\wishbone_bd_ram_mem0_reg[196][0]/P0001 ,
		_w11929_,
		_w11945_,
		_w19223_
	);
	LUT4 #(
		.INIT('h0001)
	) name8711 (
		_w19220_,
		_w19221_,
		_w19222_,
		_w19223_,
		_w19224_
	);
	LUT4 #(
		.INIT('h8000)
	) name8712 (
		_w19209_,
		_w19214_,
		_w19219_,
		_w19224_,
		_w19225_
	);
	LUT3 #(
		.INIT('h80)
	) name8713 (
		\wishbone_bd_ram_mem0_reg[205][0]/P0001 ,
		_w11945_,
		_w11966_,
		_w19226_
	);
	LUT3 #(
		.INIT('h80)
	) name8714 (
		\wishbone_bd_ram_mem0_reg[207][0]/P0001 ,
		_w11945_,
		_w11973_,
		_w19227_
	);
	LUT3 #(
		.INIT('h80)
	) name8715 (
		\wishbone_bd_ram_mem0_reg[110][0]/P0001 ,
		_w11948_,
		_w11965_,
		_w19228_
	);
	LUT3 #(
		.INIT('h80)
	) name8716 (
		\wishbone_bd_ram_mem0_reg[149][0]/P0001 ,
		_w11933_,
		_w11959_,
		_w19229_
	);
	LUT4 #(
		.INIT('h0001)
	) name8717 (
		_w19226_,
		_w19227_,
		_w19228_,
		_w19229_,
		_w19230_
	);
	LUT3 #(
		.INIT('h80)
	) name8718 (
		\wishbone_bd_ram_mem0_reg[236][0]/P0001 ,
		_w11954_,
		_w11982_,
		_w19231_
	);
	LUT3 #(
		.INIT('h80)
	) name8719 (
		\wishbone_bd_ram_mem0_reg[113][0]/P0001 ,
		_w11977_,
		_w12012_,
		_w19232_
	);
	LUT3 #(
		.INIT('h80)
	) name8720 (
		\wishbone_bd_ram_mem0_reg[109][0]/P0001 ,
		_w11965_,
		_w11966_,
		_w19233_
	);
	LUT3 #(
		.INIT('h80)
	) name8721 (
		\wishbone_bd_ram_mem0_reg[127][0]/P0001 ,
		_w11973_,
		_w12012_,
		_w19234_
	);
	LUT4 #(
		.INIT('h0001)
	) name8722 (
		_w19231_,
		_w19232_,
		_w19233_,
		_w19234_,
		_w19235_
	);
	LUT3 #(
		.INIT('h80)
	) name8723 (
		\wishbone_bd_ram_mem0_reg[171][0]/P0001 ,
		_w11930_,
		_w11936_,
		_w19236_
	);
	LUT3 #(
		.INIT('h80)
	) name8724 (
		\wishbone_bd_ram_mem0_reg[22][0]/P0001 ,
		_w11935_,
		_w11986_,
		_w19237_
	);
	LUT3 #(
		.INIT('h80)
	) name8725 (
		\wishbone_bd_ram_mem0_reg[132][0]/P0001 ,
		_w11929_,
		_w11955_,
		_w19238_
	);
	LUT3 #(
		.INIT('h80)
	) name8726 (
		\wishbone_bd_ram_mem0_reg[165][0]/P0001 ,
		_w11930_,
		_w11933_,
		_w19239_
	);
	LUT4 #(
		.INIT('h0001)
	) name8727 (
		_w19236_,
		_w19237_,
		_w19238_,
		_w19239_,
		_w19240_
	);
	LUT3 #(
		.INIT('h80)
	) name8728 (
		\wishbone_bd_ram_mem0_reg[241][0]/P0001 ,
		_w11952_,
		_w11977_,
		_w19241_
	);
	LUT3 #(
		.INIT('h80)
	) name8729 (
		\wishbone_bd_ram_mem0_reg[186][0]/P0001 ,
		_w11942_,
		_w11944_,
		_w19242_
	);
	LUT3 #(
		.INIT('h80)
	) name8730 (
		\wishbone_bd_ram_mem0_reg[119][0]/P0001 ,
		_w11975_,
		_w12012_,
		_w19243_
	);
	LUT3 #(
		.INIT('h80)
	) name8731 (
		\wishbone_bd_ram_mem0_reg[48][0]/P0001 ,
		_w11941_,
		_w11979_,
		_w19244_
	);
	LUT4 #(
		.INIT('h0001)
	) name8732 (
		_w19241_,
		_w19242_,
		_w19243_,
		_w19244_,
		_w19245_
	);
	LUT4 #(
		.INIT('h8000)
	) name8733 (
		_w19230_,
		_w19235_,
		_w19240_,
		_w19245_,
		_w19246_
	);
	LUT3 #(
		.INIT('h80)
	) name8734 (
		\wishbone_bd_ram_mem0_reg[155][0]/P0001 ,
		_w11936_,
		_w11959_,
		_w19247_
	);
	LUT3 #(
		.INIT('h80)
	) name8735 (
		\wishbone_bd_ram_mem0_reg[62][0]/P0001 ,
		_w11948_,
		_w11979_,
		_w19248_
	);
	LUT3 #(
		.INIT('h80)
	) name8736 (
		\wishbone_bd_ram_mem0_reg[148][0]/P0001 ,
		_w11929_,
		_w11959_,
		_w19249_
	);
	LUT3 #(
		.INIT('h80)
	) name8737 (
		\wishbone_bd_ram_mem0_reg[89][0]/P0001 ,
		_w11968_,
		_w11972_,
		_w19250_
	);
	LUT4 #(
		.INIT('h0001)
	) name8738 (
		_w19247_,
		_w19248_,
		_w19249_,
		_w19250_,
		_w19251_
	);
	LUT3 #(
		.INIT('h80)
	) name8739 (
		\wishbone_bd_ram_mem0_reg[213][0]/P0001 ,
		_w11933_,
		_w11984_,
		_w19252_
	);
	LUT3 #(
		.INIT('h80)
	) name8740 (
		\wishbone_bd_ram_mem0_reg[212][0]/P0001 ,
		_w11929_,
		_w11984_,
		_w19253_
	);
	LUT3 #(
		.INIT('h80)
	) name8741 (
		\wishbone_bd_ram_mem0_reg[84][0]/P0001 ,
		_w11929_,
		_w11972_,
		_w19254_
	);
	LUT3 #(
		.INIT('h80)
	) name8742 (
		\wishbone_bd_ram_mem0_reg[1][0]/P0001 ,
		_w11932_,
		_w11977_,
		_w19255_
	);
	LUT4 #(
		.INIT('h0001)
	) name8743 (
		_w19252_,
		_w19253_,
		_w19254_,
		_w19255_,
		_w19256_
	);
	LUT3 #(
		.INIT('h80)
	) name8744 (
		\wishbone_bd_ram_mem0_reg[252][0]/P0001 ,
		_w11952_,
		_w11954_,
		_w19257_
	);
	LUT3 #(
		.INIT('h80)
	) name8745 (
		\wishbone_bd_ram_mem0_reg[96][0]/P0001 ,
		_w11941_,
		_w11965_,
		_w19258_
	);
	LUT3 #(
		.INIT('h80)
	) name8746 (
		\wishbone_bd_ram_mem0_reg[123][0]/P0001 ,
		_w11936_,
		_w12012_,
		_w19259_
	);
	LUT3 #(
		.INIT('h80)
	) name8747 (
		\wishbone_bd_ram_mem0_reg[102][0]/P0001 ,
		_w11965_,
		_w11986_,
		_w19260_
	);
	LUT4 #(
		.INIT('h0001)
	) name8748 (
		_w19257_,
		_w19258_,
		_w19259_,
		_w19260_,
		_w19261_
	);
	LUT3 #(
		.INIT('h80)
	) name8749 (
		\wishbone_bd_ram_mem0_reg[41][0]/P0001 ,
		_w11957_,
		_w11968_,
		_w19262_
	);
	LUT3 #(
		.INIT('h80)
	) name8750 (
		\wishbone_bd_ram_mem0_reg[46][0]/P0001 ,
		_w11948_,
		_w11957_,
		_w19263_
	);
	LUT3 #(
		.INIT('h80)
	) name8751 (
		\wishbone_bd_ram_mem0_reg[61][0]/P0001 ,
		_w11966_,
		_w11979_,
		_w19264_
	);
	LUT3 #(
		.INIT('h80)
	) name8752 (
		\wishbone_bd_ram_mem0_reg[230][0]/P0001 ,
		_w11982_,
		_w11986_,
		_w19265_
	);
	LUT4 #(
		.INIT('h0001)
	) name8753 (
		_w19262_,
		_w19263_,
		_w19264_,
		_w19265_,
		_w19266_
	);
	LUT4 #(
		.INIT('h8000)
	) name8754 (
		_w19251_,
		_w19256_,
		_w19261_,
		_w19266_,
		_w19267_
	);
	LUT4 #(
		.INIT('h8000)
	) name8755 (
		_w19204_,
		_w19225_,
		_w19246_,
		_w19267_,
		_w19268_
	);
	LUT3 #(
		.INIT('h80)
	) name8756 (
		\wishbone_bd_ram_mem0_reg[68][0]/P0001 ,
		_w11929_,
		_w11949_,
		_w19269_
	);
	LUT3 #(
		.INIT('h80)
	) name8757 (
		\wishbone_bd_ram_mem0_reg[31][0]/P0001 ,
		_w11935_,
		_w11973_,
		_w19270_
	);
	LUT3 #(
		.INIT('h80)
	) name8758 (
		\wishbone_bd_ram_mem0_reg[209][0]/P0001 ,
		_w11977_,
		_w11984_,
		_w19271_
	);
	LUT3 #(
		.INIT('h80)
	) name8759 (
		\wishbone_bd_ram_mem0_reg[179][0]/P0001 ,
		_w11938_,
		_w11942_,
		_w19272_
	);
	LUT4 #(
		.INIT('h0001)
	) name8760 (
		_w19269_,
		_w19270_,
		_w19271_,
		_w19272_,
		_w19273_
	);
	LUT3 #(
		.INIT('h80)
	) name8761 (
		\wishbone_bd_ram_mem0_reg[223][0]/P0001 ,
		_w11973_,
		_w11984_,
		_w19274_
	);
	LUT3 #(
		.INIT('h80)
	) name8762 (
		\wishbone_bd_ram_mem0_reg[66][0]/P0001 ,
		_w11949_,
		_w11963_,
		_w19275_
	);
	LUT3 #(
		.INIT('h80)
	) name8763 (
		\wishbone_bd_ram_mem0_reg[12][0]/P0001 ,
		_w11932_,
		_w11954_,
		_w19276_
	);
	LUT3 #(
		.INIT('h80)
	) name8764 (
		\wishbone_bd_ram_mem0_reg[211][0]/P0001 ,
		_w11938_,
		_w11984_,
		_w19277_
	);
	LUT4 #(
		.INIT('h0001)
	) name8765 (
		_w19274_,
		_w19275_,
		_w19276_,
		_w19277_,
		_w19278_
	);
	LUT3 #(
		.INIT('h80)
	) name8766 (
		\wishbone_bd_ram_mem0_reg[91][0]/P0001 ,
		_w11936_,
		_w11972_,
		_w19279_
	);
	LUT3 #(
		.INIT('h80)
	) name8767 (
		\wishbone_bd_ram_mem0_reg[133][0]/P0001 ,
		_w11933_,
		_w11955_,
		_w19280_
	);
	LUT3 #(
		.INIT('h80)
	) name8768 (
		\wishbone_bd_ram_mem0_reg[234][0]/P0001 ,
		_w11944_,
		_w11982_,
		_w19281_
	);
	LUT3 #(
		.INIT('h80)
	) name8769 (
		\wishbone_bd_ram_mem0_reg[42][0]/P0001 ,
		_w11944_,
		_w11957_,
		_w19282_
	);
	LUT4 #(
		.INIT('h0001)
	) name8770 (
		_w19279_,
		_w19280_,
		_w19281_,
		_w19282_,
		_w19283_
	);
	LUT3 #(
		.INIT('h80)
	) name8771 (
		\wishbone_bd_ram_mem0_reg[237][0]/P0001 ,
		_w11966_,
		_w11982_,
		_w19284_
	);
	LUT3 #(
		.INIT('h80)
	) name8772 (
		\wishbone_bd_ram_mem0_reg[135][0]/P0001 ,
		_w11955_,
		_w11975_,
		_w19285_
	);
	LUT3 #(
		.INIT('h80)
	) name8773 (
		\wishbone_bd_ram_mem0_reg[192][0]/P0001 ,
		_w11941_,
		_w11945_,
		_w19286_
	);
	LUT3 #(
		.INIT('h80)
	) name8774 (
		\wishbone_bd_ram_mem0_reg[198][0]/P0001 ,
		_w11945_,
		_w11986_,
		_w19287_
	);
	LUT4 #(
		.INIT('h0001)
	) name8775 (
		_w19284_,
		_w19285_,
		_w19286_,
		_w19287_,
		_w19288_
	);
	LUT4 #(
		.INIT('h8000)
	) name8776 (
		_w19273_,
		_w19278_,
		_w19283_,
		_w19288_,
		_w19289_
	);
	LUT3 #(
		.INIT('h80)
	) name8777 (
		\wishbone_bd_ram_mem0_reg[183][0]/P0001 ,
		_w11942_,
		_w11975_,
		_w19290_
	);
	LUT3 #(
		.INIT('h80)
	) name8778 (
		\wishbone_bd_ram_mem0_reg[60][0]/P0001 ,
		_w11954_,
		_w11979_,
		_w19291_
	);
	LUT3 #(
		.INIT('h80)
	) name8779 (
		\wishbone_bd_ram_mem0_reg[86][0]/P0001 ,
		_w11972_,
		_w11986_,
		_w19292_
	);
	LUT3 #(
		.INIT('h80)
	) name8780 (
		\wishbone_bd_ram_mem0_reg[6][0]/P0001 ,
		_w11932_,
		_w11986_,
		_w19293_
	);
	LUT4 #(
		.INIT('h0001)
	) name8781 (
		_w19290_,
		_w19291_,
		_w19292_,
		_w19293_,
		_w19294_
	);
	LUT3 #(
		.INIT('h80)
	) name8782 (
		\wishbone_bd_ram_mem0_reg[185][0]/P0001 ,
		_w11942_,
		_w11968_,
		_w19295_
	);
	LUT3 #(
		.INIT('h80)
	) name8783 (
		\wishbone_bd_ram_mem0_reg[130][0]/P0001 ,
		_w11955_,
		_w11963_,
		_w19296_
	);
	LUT3 #(
		.INIT('h80)
	) name8784 (
		\wishbone_bd_ram_mem0_reg[235][0]/P0001 ,
		_w11936_,
		_w11982_,
		_w19297_
	);
	LUT3 #(
		.INIT('h80)
	) name8785 (
		\wishbone_bd_ram_mem0_reg[21][0]/P0001 ,
		_w11933_,
		_w11935_,
		_w19298_
	);
	LUT4 #(
		.INIT('h0001)
	) name8786 (
		_w19295_,
		_w19296_,
		_w19297_,
		_w19298_,
		_w19299_
	);
	LUT3 #(
		.INIT('h80)
	) name8787 (
		\wishbone_bd_ram_mem0_reg[175][0]/P0001 ,
		_w11930_,
		_w11973_,
		_w19300_
	);
	LUT3 #(
		.INIT('h80)
	) name8788 (
		\wishbone_bd_ram_mem0_reg[36][0]/P0001 ,
		_w11929_,
		_w11957_,
		_w19301_
	);
	LUT3 #(
		.INIT('h80)
	) name8789 (
		\wishbone_bd_ram_mem0_reg[247][0]/P0001 ,
		_w11952_,
		_w11975_,
		_w19302_
	);
	LUT3 #(
		.INIT('h80)
	) name8790 (
		\wishbone_bd_ram_mem0_reg[215][0]/P0001 ,
		_w11975_,
		_w11984_,
		_w19303_
	);
	LUT4 #(
		.INIT('h0001)
	) name8791 (
		_w19300_,
		_w19301_,
		_w19302_,
		_w19303_,
		_w19304_
	);
	LUT3 #(
		.INIT('h80)
	) name8792 (
		\wishbone_bd_ram_mem0_reg[197][0]/P0001 ,
		_w11933_,
		_w11945_,
		_w19305_
	);
	LUT3 #(
		.INIT('h80)
	) name8793 (
		\wishbone_bd_ram_mem0_reg[122][0]/P0001 ,
		_w11944_,
		_w12012_,
		_w19306_
	);
	LUT3 #(
		.INIT('h80)
	) name8794 (
		\wishbone_bd_ram_mem0_reg[244][0]/P0001 ,
		_w11929_,
		_w11952_,
		_w19307_
	);
	LUT3 #(
		.INIT('h80)
	) name8795 (
		\wishbone_bd_ram_mem0_reg[93][0]/P0001 ,
		_w11966_,
		_w11972_,
		_w19308_
	);
	LUT4 #(
		.INIT('h0001)
	) name8796 (
		_w19305_,
		_w19306_,
		_w19307_,
		_w19308_,
		_w19309_
	);
	LUT4 #(
		.INIT('h8000)
	) name8797 (
		_w19294_,
		_w19299_,
		_w19304_,
		_w19309_,
		_w19310_
	);
	LUT3 #(
		.INIT('h80)
	) name8798 (
		\wishbone_bd_ram_mem0_reg[195][0]/P0001 ,
		_w11938_,
		_w11945_,
		_w19311_
	);
	LUT3 #(
		.INIT('h80)
	) name8799 (
		\wishbone_bd_ram_mem0_reg[226][0]/P0001 ,
		_w11963_,
		_w11982_,
		_w19312_
	);
	LUT3 #(
		.INIT('h80)
	) name8800 (
		\wishbone_bd_ram_mem0_reg[24][0]/P0001 ,
		_w11935_,
		_w11990_,
		_w19313_
	);
	LUT3 #(
		.INIT('h80)
	) name8801 (
		\wishbone_bd_ram_mem0_reg[8][0]/P0001 ,
		_w11932_,
		_w11990_,
		_w19314_
	);
	LUT4 #(
		.INIT('h0001)
	) name8802 (
		_w19311_,
		_w19312_,
		_w19313_,
		_w19314_,
		_w19315_
	);
	LUT3 #(
		.INIT('h80)
	) name8803 (
		\wishbone_bd_ram_mem0_reg[199][0]/P0001 ,
		_w11945_,
		_w11975_,
		_w19316_
	);
	LUT3 #(
		.INIT('h80)
	) name8804 (
		\wishbone_bd_ram_mem0_reg[250][0]/P0001 ,
		_w11944_,
		_w11952_,
		_w19317_
	);
	LUT3 #(
		.INIT('h80)
	) name8805 (
		\wishbone_bd_ram_mem0_reg[5][0]/P0001 ,
		_w11932_,
		_w11933_,
		_w19318_
	);
	LUT3 #(
		.INIT('h80)
	) name8806 (
		\wishbone_bd_ram_mem0_reg[9][0]/P0001 ,
		_w11932_,
		_w11968_,
		_w19319_
	);
	LUT4 #(
		.INIT('h0001)
	) name8807 (
		_w19316_,
		_w19317_,
		_w19318_,
		_w19319_,
		_w19320_
	);
	LUT3 #(
		.INIT('h80)
	) name8808 (
		\wishbone_bd_ram_mem0_reg[214][0]/P0001 ,
		_w11984_,
		_w11986_,
		_w19321_
	);
	LUT3 #(
		.INIT('h80)
	) name8809 (
		\wishbone_bd_ram_mem0_reg[203][0]/P0001 ,
		_w11936_,
		_w11945_,
		_w19322_
	);
	LUT3 #(
		.INIT('h80)
	) name8810 (
		\wishbone_bd_ram_mem0_reg[232][0]/P0001 ,
		_w11982_,
		_w11990_,
		_w19323_
	);
	LUT3 #(
		.INIT('h80)
	) name8811 (
		\wishbone_bd_ram_mem0_reg[140][0]/P0001 ,
		_w11954_,
		_w11955_,
		_w19324_
	);
	LUT4 #(
		.INIT('h0001)
	) name8812 (
		_w19321_,
		_w19322_,
		_w19323_,
		_w19324_,
		_w19325_
	);
	LUT3 #(
		.INIT('h80)
	) name8813 (
		\wishbone_bd_ram_mem0_reg[64][0]/P0001 ,
		_w11941_,
		_w11949_,
		_w19326_
	);
	LUT3 #(
		.INIT('h80)
	) name8814 (
		\wishbone_bd_ram_mem0_reg[222][0]/P0001 ,
		_w11948_,
		_w11984_,
		_w19327_
	);
	LUT3 #(
		.INIT('h80)
	) name8815 (
		\wishbone_bd_ram_mem0_reg[10][0]/P0001 ,
		_w11932_,
		_w11944_,
		_w19328_
	);
	LUT3 #(
		.INIT('h80)
	) name8816 (
		\wishbone_bd_ram_mem0_reg[28][0]/P0001 ,
		_w11935_,
		_w11954_,
		_w19329_
	);
	LUT4 #(
		.INIT('h0001)
	) name8817 (
		_w19326_,
		_w19327_,
		_w19328_,
		_w19329_,
		_w19330_
	);
	LUT4 #(
		.INIT('h8000)
	) name8818 (
		_w19315_,
		_w19320_,
		_w19325_,
		_w19330_,
		_w19331_
	);
	LUT3 #(
		.INIT('h80)
	) name8819 (
		\wishbone_bd_ram_mem0_reg[144][0]/P0001 ,
		_w11941_,
		_w11959_,
		_w19332_
	);
	LUT3 #(
		.INIT('h80)
	) name8820 (
		\wishbone_bd_ram_mem0_reg[188][0]/P0001 ,
		_w11942_,
		_w11954_,
		_w19333_
	);
	LUT3 #(
		.INIT('h80)
	) name8821 (
		\wishbone_bd_ram_mem0_reg[249][0]/P0001 ,
		_w11952_,
		_w11968_,
		_w19334_
	);
	LUT3 #(
		.INIT('h80)
	) name8822 (
		\wishbone_bd_ram_mem0_reg[251][0]/P0001 ,
		_w11936_,
		_w11952_,
		_w19335_
	);
	LUT4 #(
		.INIT('h0001)
	) name8823 (
		_w19332_,
		_w19333_,
		_w19334_,
		_w19335_,
		_w19336_
	);
	LUT3 #(
		.INIT('h80)
	) name8824 (
		\wishbone_bd_ram_mem0_reg[87][0]/P0001 ,
		_w11972_,
		_w11975_,
		_w19337_
	);
	LUT3 #(
		.INIT('h80)
	) name8825 (
		\wishbone_bd_ram_mem0_reg[82][0]/P0001 ,
		_w11963_,
		_w11972_,
		_w19338_
	);
	LUT3 #(
		.INIT('h80)
	) name8826 (
		\wishbone_bd_ram_mem0_reg[11][0]/P0001 ,
		_w11932_,
		_w11936_,
		_w19339_
	);
	LUT3 #(
		.INIT('h80)
	) name8827 (
		\wishbone_bd_ram_mem0_reg[81][0]/P0001 ,
		_w11972_,
		_w11977_,
		_w19340_
	);
	LUT4 #(
		.INIT('h0001)
	) name8828 (
		_w19337_,
		_w19338_,
		_w19339_,
		_w19340_,
		_w19341_
	);
	LUT3 #(
		.INIT('h80)
	) name8829 (
		\wishbone_bd_ram_mem0_reg[160][0]/P0001 ,
		_w11930_,
		_w11941_,
		_w19342_
	);
	LUT3 #(
		.INIT('h80)
	) name8830 (
		\wishbone_bd_ram_mem0_reg[32][0]/P0001 ,
		_w11941_,
		_w11957_,
		_w19343_
	);
	LUT3 #(
		.INIT('h80)
	) name8831 (
		\wishbone_bd_ram_mem0_reg[169][0]/P0001 ,
		_w11930_,
		_w11968_,
		_w19344_
	);
	LUT3 #(
		.INIT('h80)
	) name8832 (
		\wishbone_bd_ram_mem0_reg[216][0]/P0001 ,
		_w11984_,
		_w11990_,
		_w19345_
	);
	LUT4 #(
		.INIT('h0001)
	) name8833 (
		_w19342_,
		_w19343_,
		_w19344_,
		_w19345_,
		_w19346_
	);
	LUT3 #(
		.INIT('h80)
	) name8834 (
		\wishbone_bd_ram_mem0_reg[18][0]/P0001 ,
		_w11935_,
		_w11963_,
		_w19347_
	);
	LUT3 #(
		.INIT('h80)
	) name8835 (
		\wishbone_bd_ram_mem0_reg[111][0]/P0001 ,
		_w11965_,
		_w11973_,
		_w19348_
	);
	LUT3 #(
		.INIT('h80)
	) name8836 (
		\wishbone_bd_ram_mem0_reg[242][0]/P0001 ,
		_w11952_,
		_w11963_,
		_w19349_
	);
	LUT3 #(
		.INIT('h80)
	) name8837 (
		\wishbone_bd_ram_mem0_reg[78][0]/P0001 ,
		_w11948_,
		_w11949_,
		_w19350_
	);
	LUT4 #(
		.INIT('h0001)
	) name8838 (
		_w19347_,
		_w19348_,
		_w19349_,
		_w19350_,
		_w19351_
	);
	LUT4 #(
		.INIT('h8000)
	) name8839 (
		_w19336_,
		_w19341_,
		_w19346_,
		_w19351_,
		_w19352_
	);
	LUT4 #(
		.INIT('h8000)
	) name8840 (
		_w19289_,
		_w19310_,
		_w19331_,
		_w19352_,
		_w19353_
	);
	LUT3 #(
		.INIT('h80)
	) name8841 (
		\wishbone_bd_ram_mem0_reg[57][0]/P0001 ,
		_w11968_,
		_w11979_,
		_w19354_
	);
	LUT3 #(
		.INIT('h80)
	) name8842 (
		\wishbone_bd_ram_mem0_reg[177][0]/P0001 ,
		_w11942_,
		_w11977_,
		_w19355_
	);
	LUT3 #(
		.INIT('h80)
	) name8843 (
		\wishbone_bd_ram_mem0_reg[163][0]/P0001 ,
		_w11930_,
		_w11938_,
		_w19356_
	);
	LUT3 #(
		.INIT('h80)
	) name8844 (
		\wishbone_bd_ram_mem0_reg[190][0]/P0001 ,
		_w11942_,
		_w11948_,
		_w19357_
	);
	LUT4 #(
		.INIT('h0001)
	) name8845 (
		_w19354_,
		_w19355_,
		_w19356_,
		_w19357_,
		_w19358_
	);
	LUT3 #(
		.INIT('h80)
	) name8846 (
		\wishbone_bd_ram_mem0_reg[243][0]/P0001 ,
		_w11938_,
		_w11952_,
		_w19359_
	);
	LUT3 #(
		.INIT('h80)
	) name8847 (
		\wishbone_bd_ram_mem0_reg[191][0]/P0001 ,
		_w11942_,
		_w11973_,
		_w19360_
	);
	LUT3 #(
		.INIT('h80)
	) name8848 (
		\wishbone_bd_ram_mem0_reg[217][0]/P0001 ,
		_w11968_,
		_w11984_,
		_w19361_
	);
	LUT3 #(
		.INIT('h80)
	) name8849 (
		\wishbone_bd_ram_mem0_reg[229][0]/P0001 ,
		_w11933_,
		_w11982_,
		_w19362_
	);
	LUT4 #(
		.INIT('h0001)
	) name8850 (
		_w19359_,
		_w19360_,
		_w19361_,
		_w19362_,
		_w19363_
	);
	LUT3 #(
		.INIT('h80)
	) name8851 (
		\wishbone_bd_ram_mem0_reg[231][0]/P0001 ,
		_w11975_,
		_w11982_,
		_w19364_
	);
	LUT3 #(
		.INIT('h80)
	) name8852 (
		\wishbone_bd_ram_mem0_reg[77][0]/P0001 ,
		_w11949_,
		_w11966_,
		_w19365_
	);
	LUT3 #(
		.INIT('h80)
	) name8853 (
		\wishbone_bd_ram_mem0_reg[37][0]/P0001 ,
		_w11933_,
		_w11957_,
		_w19366_
	);
	LUT3 #(
		.INIT('h80)
	) name8854 (
		\wishbone_bd_ram_mem0_reg[181][0]/P0001 ,
		_w11933_,
		_w11942_,
		_w19367_
	);
	LUT4 #(
		.INIT('h0001)
	) name8855 (
		_w19364_,
		_w19365_,
		_w19366_,
		_w19367_,
		_w19368_
	);
	LUT3 #(
		.INIT('h80)
	) name8856 (
		\wishbone_bd_ram_mem0_reg[120][0]/P0001 ,
		_w11990_,
		_w12012_,
		_w19369_
	);
	LUT3 #(
		.INIT('h80)
	) name8857 (
		\wishbone_bd_ram_mem0_reg[17][0]/P0001 ,
		_w11935_,
		_w11977_,
		_w19370_
	);
	LUT3 #(
		.INIT('h80)
	) name8858 (
		\wishbone_bd_ram_mem0_reg[225][0]/P0001 ,
		_w11977_,
		_w11982_,
		_w19371_
	);
	LUT3 #(
		.INIT('h80)
	) name8859 (
		\wishbone_bd_ram_mem0_reg[219][0]/P0001 ,
		_w11936_,
		_w11984_,
		_w19372_
	);
	LUT4 #(
		.INIT('h0001)
	) name8860 (
		_w19369_,
		_w19370_,
		_w19371_,
		_w19372_,
		_w19373_
	);
	LUT4 #(
		.INIT('h8000)
	) name8861 (
		_w19358_,
		_w19363_,
		_w19368_,
		_w19373_,
		_w19374_
	);
	LUT3 #(
		.INIT('h80)
	) name8862 (
		\wishbone_bd_ram_mem0_reg[227][0]/P0001 ,
		_w11938_,
		_w11982_,
		_w19375_
	);
	LUT3 #(
		.INIT('h80)
	) name8863 (
		\wishbone_bd_ram_mem0_reg[106][0]/P0001 ,
		_w11944_,
		_w11965_,
		_w19376_
	);
	LUT3 #(
		.INIT('h80)
	) name8864 (
		\wishbone_bd_ram_mem0_reg[161][0]/P0001 ,
		_w11930_,
		_w11977_,
		_w19377_
	);
	LUT3 #(
		.INIT('h80)
	) name8865 (
		\wishbone_bd_ram_mem0_reg[85][0]/P0001 ,
		_w11933_,
		_w11972_,
		_w19378_
	);
	LUT4 #(
		.INIT('h0001)
	) name8866 (
		_w19375_,
		_w19376_,
		_w19377_,
		_w19378_,
		_w19379_
	);
	LUT3 #(
		.INIT('h80)
	) name8867 (
		\wishbone_bd_ram_mem0_reg[75][0]/P0001 ,
		_w11936_,
		_w11949_,
		_w19380_
	);
	LUT3 #(
		.INIT('h80)
	) name8868 (
		\wishbone_bd_ram_mem0_reg[168][0]/P0001 ,
		_w11930_,
		_w11990_,
		_w19381_
	);
	LUT3 #(
		.INIT('h80)
	) name8869 (
		\wishbone_bd_ram_mem0_reg[240][0]/P0001 ,
		_w11941_,
		_w11952_,
		_w19382_
	);
	LUT3 #(
		.INIT('h80)
	) name8870 (
		\wishbone_bd_ram_mem0_reg[152][0]/P0001 ,
		_w11959_,
		_w11990_,
		_w19383_
	);
	LUT4 #(
		.INIT('h0001)
	) name8871 (
		_w19380_,
		_w19381_,
		_w19382_,
		_w19383_,
		_w19384_
	);
	LUT3 #(
		.INIT('h80)
	) name8872 (
		\wishbone_bd_ram_mem0_reg[90][0]/P0001 ,
		_w11944_,
		_w11972_,
		_w19385_
	);
	LUT3 #(
		.INIT('h80)
	) name8873 (
		\wishbone_bd_ram_mem0_reg[128][0]/P0001 ,
		_w11941_,
		_w11955_,
		_w19386_
	);
	LUT3 #(
		.INIT('h80)
	) name8874 (
		\wishbone_bd_ram_mem0_reg[187][0]/P0001 ,
		_w11936_,
		_w11942_,
		_w19387_
	);
	LUT3 #(
		.INIT('h80)
	) name8875 (
		\wishbone_bd_ram_mem0_reg[248][0]/P0001 ,
		_w11952_,
		_w11990_,
		_w19388_
	);
	LUT4 #(
		.INIT('h0001)
	) name8876 (
		_w19385_,
		_w19386_,
		_w19387_,
		_w19388_,
		_w19389_
	);
	LUT3 #(
		.INIT('h80)
	) name8877 (
		\wishbone_bd_ram_mem0_reg[202][0]/P0001 ,
		_w11944_,
		_w11945_,
		_w19390_
	);
	LUT3 #(
		.INIT('h80)
	) name8878 (
		\wishbone_bd_ram_mem0_reg[23][0]/P0001 ,
		_w11935_,
		_w11975_,
		_w19391_
	);
	LUT3 #(
		.INIT('h80)
	) name8879 (
		\wishbone_bd_ram_mem0_reg[208][0]/P0001 ,
		_w11941_,
		_w11984_,
		_w19392_
	);
	LUT3 #(
		.INIT('h80)
	) name8880 (
		\wishbone_bd_ram_mem0_reg[76][0]/P0001 ,
		_w11949_,
		_w11954_,
		_w19393_
	);
	LUT4 #(
		.INIT('h0001)
	) name8881 (
		_w19390_,
		_w19391_,
		_w19392_,
		_w19393_,
		_w19394_
	);
	LUT4 #(
		.INIT('h8000)
	) name8882 (
		_w19379_,
		_w19384_,
		_w19389_,
		_w19394_,
		_w19395_
	);
	LUT3 #(
		.INIT('h80)
	) name8883 (
		\wishbone_bd_ram_mem0_reg[246][0]/P0001 ,
		_w11952_,
		_w11986_,
		_w19396_
	);
	LUT3 #(
		.INIT('h80)
	) name8884 (
		\wishbone_bd_ram_mem0_reg[193][0]/P0001 ,
		_w11945_,
		_w11977_,
		_w19397_
	);
	LUT3 #(
		.INIT('h80)
	) name8885 (
		\wishbone_bd_ram_mem0_reg[50][0]/P0001 ,
		_w11963_,
		_w11979_,
		_w19398_
	);
	LUT3 #(
		.INIT('h80)
	) name8886 (
		\wishbone_bd_ram_mem0_reg[38][0]/P0001 ,
		_w11957_,
		_w11986_,
		_w19399_
	);
	LUT4 #(
		.INIT('h0001)
	) name8887 (
		_w19396_,
		_w19397_,
		_w19398_,
		_w19399_,
		_w19400_
	);
	LUT3 #(
		.INIT('h80)
	) name8888 (
		\wishbone_bd_ram_mem0_reg[147][0]/P0001 ,
		_w11938_,
		_w11959_,
		_w19401_
	);
	LUT3 #(
		.INIT('h80)
	) name8889 (
		\wishbone_bd_ram_mem0_reg[49][0]/P0001 ,
		_w11977_,
		_w11979_,
		_w19402_
	);
	LUT3 #(
		.INIT('h80)
	) name8890 (
		\wishbone_bd_ram_mem0_reg[94][0]/P0001 ,
		_w11948_,
		_w11972_,
		_w19403_
	);
	LUT3 #(
		.INIT('h80)
	) name8891 (
		\wishbone_bd_ram_mem0_reg[74][0]/P0001 ,
		_w11944_,
		_w11949_,
		_w19404_
	);
	LUT4 #(
		.INIT('h0001)
	) name8892 (
		_w19401_,
		_w19402_,
		_w19403_,
		_w19404_,
		_w19405_
	);
	LUT3 #(
		.INIT('h80)
	) name8893 (
		\wishbone_bd_ram_mem0_reg[33][0]/P0001 ,
		_w11957_,
		_w11977_,
		_w19406_
	);
	LUT3 #(
		.INIT('h80)
	) name8894 (
		\wishbone_bd_ram_mem0_reg[134][0]/P0001 ,
		_w11955_,
		_w11986_,
		_w19407_
	);
	LUT3 #(
		.INIT('h80)
	) name8895 (
		\wishbone_bd_ram_mem0_reg[180][0]/P0001 ,
		_w11929_,
		_w11942_,
		_w19408_
	);
	LUT3 #(
		.INIT('h80)
	) name8896 (
		\wishbone_bd_ram_mem0_reg[98][0]/P0001 ,
		_w11963_,
		_w11965_,
		_w19409_
	);
	LUT4 #(
		.INIT('h0001)
	) name8897 (
		_w19406_,
		_w19407_,
		_w19408_,
		_w19409_,
		_w19410_
	);
	LUT3 #(
		.INIT('h80)
	) name8898 (
		\wishbone_bd_ram_mem0_reg[121][0]/P0001 ,
		_w11968_,
		_w12012_,
		_w19411_
	);
	LUT3 #(
		.INIT('h80)
	) name8899 (
		\wishbone_bd_ram_mem0_reg[162][0]/P0001 ,
		_w11930_,
		_w11963_,
		_w19412_
	);
	LUT3 #(
		.INIT('h80)
	) name8900 (
		\wishbone_bd_ram_mem0_reg[210][0]/P0001 ,
		_w11963_,
		_w11984_,
		_w19413_
	);
	LUT3 #(
		.INIT('h80)
	) name8901 (
		\wishbone_bd_ram_mem0_reg[176][0]/P0001 ,
		_w11941_,
		_w11942_,
		_w19414_
	);
	LUT4 #(
		.INIT('h0001)
	) name8902 (
		_w19411_,
		_w19412_,
		_w19413_,
		_w19414_,
		_w19415_
	);
	LUT4 #(
		.INIT('h8000)
	) name8903 (
		_w19400_,
		_w19405_,
		_w19410_,
		_w19415_,
		_w19416_
	);
	LUT3 #(
		.INIT('h80)
	) name8904 (
		\wishbone_bd_ram_mem0_reg[200][0]/P0001 ,
		_w11945_,
		_w11990_,
		_w19417_
	);
	LUT3 #(
		.INIT('h80)
	) name8905 (
		\wishbone_bd_ram_mem0_reg[125][0]/P0001 ,
		_w11966_,
		_w12012_,
		_w19418_
	);
	LUT3 #(
		.INIT('h80)
	) name8906 (
		\wishbone_bd_ram_mem0_reg[124][0]/P0001 ,
		_w11954_,
		_w12012_,
		_w19419_
	);
	LUT3 #(
		.INIT('h80)
	) name8907 (
		\wishbone_bd_ram_mem0_reg[15][0]/P0001 ,
		_w11932_,
		_w11973_,
		_w19420_
	);
	LUT4 #(
		.INIT('h0001)
	) name8908 (
		_w19417_,
		_w19418_,
		_w19419_,
		_w19420_,
		_w19421_
	);
	LUT3 #(
		.INIT('h80)
	) name8909 (
		\wishbone_bd_ram_mem0_reg[44][0]/P0001 ,
		_w11954_,
		_w11957_,
		_w19422_
	);
	LUT3 #(
		.INIT('h80)
	) name8910 (
		\wishbone_bd_ram_mem0_reg[118][0]/P0001 ,
		_w11986_,
		_w12012_,
		_w19423_
	);
	LUT3 #(
		.INIT('h80)
	) name8911 (
		\wishbone_bd_ram_mem0_reg[137][0]/P0001 ,
		_w11955_,
		_w11968_,
		_w19424_
	);
	LUT3 #(
		.INIT('h80)
	) name8912 (
		\wishbone_bd_ram_mem0_reg[43][0]/P0001 ,
		_w11936_,
		_w11957_,
		_w19425_
	);
	LUT4 #(
		.INIT('h0001)
	) name8913 (
		_w19422_,
		_w19423_,
		_w19424_,
		_w19425_,
		_w19426_
	);
	LUT3 #(
		.INIT('h80)
	) name8914 (
		\wishbone_bd_ram_mem0_reg[55][0]/P0001 ,
		_w11975_,
		_w11979_,
		_w19427_
	);
	LUT3 #(
		.INIT('h80)
	) name8915 (
		\wishbone_bd_ram_mem0_reg[131][0]/P0001 ,
		_w11938_,
		_w11955_,
		_w19428_
	);
	LUT3 #(
		.INIT('h80)
	) name8916 (
		\wishbone_bd_ram_mem0_reg[233][0]/P0001 ,
		_w11968_,
		_w11982_,
		_w19429_
	);
	LUT3 #(
		.INIT('h80)
	) name8917 (
		\wishbone_bd_ram_mem0_reg[158][0]/P0001 ,
		_w11948_,
		_w11959_,
		_w19430_
	);
	LUT4 #(
		.INIT('h0001)
	) name8918 (
		_w19427_,
		_w19428_,
		_w19429_,
		_w19430_,
		_w19431_
	);
	LUT3 #(
		.INIT('h80)
	) name8919 (
		\wishbone_bd_ram_mem0_reg[63][0]/P0001 ,
		_w11973_,
		_w11979_,
		_w19432_
	);
	LUT3 #(
		.INIT('h80)
	) name8920 (
		\wishbone_bd_ram_mem0_reg[69][0]/P0001 ,
		_w11933_,
		_w11949_,
		_w19433_
	);
	LUT3 #(
		.INIT('h80)
	) name8921 (
		\wishbone_bd_ram_mem0_reg[40][0]/P0001 ,
		_w11957_,
		_w11990_,
		_w19434_
	);
	LUT3 #(
		.INIT('h80)
	) name8922 (
		\wishbone_bd_ram_mem0_reg[16][0]/P0001 ,
		_w11935_,
		_w11941_,
		_w19435_
	);
	LUT4 #(
		.INIT('h0001)
	) name8923 (
		_w19432_,
		_w19433_,
		_w19434_,
		_w19435_,
		_w19436_
	);
	LUT4 #(
		.INIT('h8000)
	) name8924 (
		_w19421_,
		_w19426_,
		_w19431_,
		_w19436_,
		_w19437_
	);
	LUT4 #(
		.INIT('h8000)
	) name8925 (
		_w19374_,
		_w19395_,
		_w19416_,
		_w19437_,
		_w19438_
	);
	LUT3 #(
		.INIT('h80)
	) name8926 (
		\wishbone_bd_ram_mem0_reg[20][0]/P0001 ,
		_w11929_,
		_w11935_,
		_w19439_
	);
	LUT3 #(
		.INIT('h80)
	) name8927 (
		\wishbone_bd_ram_mem0_reg[178][0]/P0001 ,
		_w11942_,
		_w11963_,
		_w19440_
	);
	LUT3 #(
		.INIT('h80)
	) name8928 (
		\wishbone_bd_ram_mem0_reg[139][0]/P0001 ,
		_w11936_,
		_w11955_,
		_w19441_
	);
	LUT3 #(
		.INIT('h80)
	) name8929 (
		\wishbone_bd_ram_mem0_reg[206][0]/P0001 ,
		_w11945_,
		_w11948_,
		_w19442_
	);
	LUT4 #(
		.INIT('h0001)
	) name8930 (
		_w19439_,
		_w19440_,
		_w19441_,
		_w19442_,
		_w19443_
	);
	LUT3 #(
		.INIT('h80)
	) name8931 (
		\wishbone_bd_ram_mem0_reg[255][0]/P0001 ,
		_w11952_,
		_w11973_,
		_w19444_
	);
	LUT3 #(
		.INIT('h80)
	) name8932 (
		\wishbone_bd_ram_mem0_reg[138][0]/P0001 ,
		_w11944_,
		_w11955_,
		_w19445_
	);
	LUT3 #(
		.INIT('h80)
	) name8933 (
		\wishbone_bd_ram_mem0_reg[104][0]/P0001 ,
		_w11965_,
		_w11990_,
		_w19446_
	);
	LUT3 #(
		.INIT('h80)
	) name8934 (
		\wishbone_bd_ram_mem0_reg[167][0]/P0001 ,
		_w11930_,
		_w11975_,
		_w19447_
	);
	LUT4 #(
		.INIT('h0001)
	) name8935 (
		_w19444_,
		_w19445_,
		_w19446_,
		_w19447_,
		_w19448_
	);
	LUT3 #(
		.INIT('h80)
	) name8936 (
		\wishbone_bd_ram_mem0_reg[218][0]/P0001 ,
		_w11944_,
		_w11984_,
		_w19449_
	);
	LUT3 #(
		.INIT('h80)
	) name8937 (
		\wishbone_bd_ram_mem0_reg[239][0]/P0001 ,
		_w11973_,
		_w11982_,
		_w19450_
	);
	LUT3 #(
		.INIT('h80)
	) name8938 (
		\wishbone_bd_ram_mem0_reg[92][0]/P0001 ,
		_w11954_,
		_w11972_,
		_w19451_
	);
	LUT3 #(
		.INIT('h80)
	) name8939 (
		\wishbone_bd_ram_mem0_reg[173][0]/P0001 ,
		_w11930_,
		_w11966_,
		_w19452_
	);
	LUT4 #(
		.INIT('h0001)
	) name8940 (
		_w19449_,
		_w19450_,
		_w19451_,
		_w19452_,
		_w19453_
	);
	LUT3 #(
		.INIT('h80)
	) name8941 (
		\wishbone_bd_ram_mem0_reg[129][0]/P0001 ,
		_w11955_,
		_w11977_,
		_w19454_
	);
	LUT3 #(
		.INIT('h80)
	) name8942 (
		\wishbone_bd_ram_mem0_reg[56][0]/P0001 ,
		_w11979_,
		_w11990_,
		_w19455_
	);
	LUT3 #(
		.INIT('h80)
	) name8943 (
		\wishbone_bd_ram_mem0_reg[19][0]/P0001 ,
		_w11935_,
		_w11938_,
		_w19456_
	);
	LUT3 #(
		.INIT('h80)
	) name8944 (
		\wishbone_bd_ram_mem0_reg[108][0]/P0001 ,
		_w11954_,
		_w11965_,
		_w19457_
	);
	LUT4 #(
		.INIT('h0001)
	) name8945 (
		_w19454_,
		_w19455_,
		_w19456_,
		_w19457_,
		_w19458_
	);
	LUT4 #(
		.INIT('h8000)
	) name8946 (
		_w19443_,
		_w19448_,
		_w19453_,
		_w19458_,
		_w19459_
	);
	LUT3 #(
		.INIT('h80)
	) name8947 (
		\wishbone_bd_ram_mem0_reg[52][0]/P0001 ,
		_w11929_,
		_w11979_,
		_w19460_
	);
	LUT3 #(
		.INIT('h80)
	) name8948 (
		\wishbone_bd_ram_mem0_reg[201][0]/P0001 ,
		_w11945_,
		_w11968_,
		_w19461_
	);
	LUT3 #(
		.INIT('h80)
	) name8949 (
		\wishbone_bd_ram_mem0_reg[4][0]/P0001 ,
		_w11929_,
		_w11932_,
		_w19462_
	);
	LUT3 #(
		.INIT('h80)
	) name8950 (
		\wishbone_bd_ram_mem0_reg[107][0]/P0001 ,
		_w11936_,
		_w11965_,
		_w19463_
	);
	LUT4 #(
		.INIT('h0001)
	) name8951 (
		_w19460_,
		_w19461_,
		_w19462_,
		_w19463_,
		_w19464_
	);
	LUT3 #(
		.INIT('h80)
	) name8952 (
		\wishbone_bd_ram_mem0_reg[141][0]/P0001 ,
		_w11955_,
		_w11966_,
		_w19465_
	);
	LUT3 #(
		.INIT('h80)
	) name8953 (
		\wishbone_bd_ram_mem0_reg[105][0]/P0001 ,
		_w11965_,
		_w11968_,
		_w19466_
	);
	LUT3 #(
		.INIT('h80)
	) name8954 (
		\wishbone_bd_ram_mem0_reg[59][0]/P0001 ,
		_w11936_,
		_w11979_,
		_w19467_
	);
	LUT3 #(
		.INIT('h80)
	) name8955 (
		\wishbone_bd_ram_mem0_reg[51][0]/P0001 ,
		_w11938_,
		_w11979_,
		_w19468_
	);
	LUT4 #(
		.INIT('h0001)
	) name8956 (
		_w19465_,
		_w19466_,
		_w19467_,
		_w19468_,
		_w19469_
	);
	LUT3 #(
		.INIT('h80)
	) name8957 (
		\wishbone_bd_ram_mem0_reg[34][0]/P0001 ,
		_w11957_,
		_w11963_,
		_w19470_
	);
	LUT3 #(
		.INIT('h80)
	) name8958 (
		\wishbone_bd_ram_mem0_reg[70][0]/P0001 ,
		_w11949_,
		_w11986_,
		_w19471_
	);
	LUT3 #(
		.INIT('h80)
	) name8959 (
		\wishbone_bd_ram_mem0_reg[73][0]/P0001 ,
		_w11949_,
		_w11968_,
		_w19472_
	);
	LUT3 #(
		.INIT('h80)
	) name8960 (
		\wishbone_bd_ram_mem0_reg[157][0]/P0001 ,
		_w11959_,
		_w11966_,
		_w19473_
	);
	LUT4 #(
		.INIT('h0001)
	) name8961 (
		_w19470_,
		_w19471_,
		_w19472_,
		_w19473_,
		_w19474_
	);
	LUT3 #(
		.INIT('h80)
	) name8962 (
		\wishbone_bd_ram_mem0_reg[88][0]/P0001 ,
		_w11972_,
		_w11990_,
		_w19475_
	);
	LUT3 #(
		.INIT('h80)
	) name8963 (
		\wishbone_bd_ram_mem0_reg[204][0]/P0001 ,
		_w11945_,
		_w11954_,
		_w19476_
	);
	LUT3 #(
		.INIT('h80)
	) name8964 (
		\wishbone_bd_ram_mem0_reg[54][0]/P0001 ,
		_w11979_,
		_w11986_,
		_w19477_
	);
	LUT3 #(
		.INIT('h80)
	) name8965 (
		\wishbone_bd_ram_mem0_reg[117][0]/P0001 ,
		_w11933_,
		_w12012_,
		_w19478_
	);
	LUT4 #(
		.INIT('h0001)
	) name8966 (
		_w19475_,
		_w19476_,
		_w19477_,
		_w19478_,
		_w19479_
	);
	LUT4 #(
		.INIT('h8000)
	) name8967 (
		_w19464_,
		_w19469_,
		_w19474_,
		_w19479_,
		_w19480_
	);
	LUT3 #(
		.INIT('h80)
	) name8968 (
		\wishbone_bd_ram_mem0_reg[95][0]/P0001 ,
		_w11972_,
		_w11973_,
		_w19481_
	);
	LUT3 #(
		.INIT('h80)
	) name8969 (
		\wishbone_bd_ram_mem0_reg[156][0]/P0001 ,
		_w11954_,
		_w11959_,
		_w19482_
	);
	LUT3 #(
		.INIT('h80)
	) name8970 (
		\wishbone_bd_ram_mem0_reg[72][0]/P0001 ,
		_w11949_,
		_w11990_,
		_w19483_
	);
	LUT3 #(
		.INIT('h80)
	) name8971 (
		\wishbone_bd_ram_mem0_reg[142][0]/P0001 ,
		_w11948_,
		_w11955_,
		_w19484_
	);
	LUT4 #(
		.INIT('h0001)
	) name8972 (
		_w19481_,
		_w19482_,
		_w19483_,
		_w19484_,
		_w19485_
	);
	LUT3 #(
		.INIT('h80)
	) name8973 (
		\wishbone_bd_ram_mem0_reg[224][0]/P0001 ,
		_w11941_,
		_w11982_,
		_w19486_
	);
	LUT3 #(
		.INIT('h80)
	) name8974 (
		\wishbone_bd_ram_mem0_reg[53][0]/P0001 ,
		_w11933_,
		_w11979_,
		_w19487_
	);
	LUT3 #(
		.INIT('h80)
	) name8975 (
		\wishbone_bd_ram_mem0_reg[253][0]/P0001 ,
		_w11952_,
		_w11966_,
		_w19488_
	);
	LUT3 #(
		.INIT('h80)
	) name8976 (
		\wishbone_bd_ram_mem0_reg[170][0]/P0001 ,
		_w11930_,
		_w11944_,
		_w19489_
	);
	LUT4 #(
		.INIT('h0001)
	) name8977 (
		_w19486_,
		_w19487_,
		_w19488_,
		_w19489_,
		_w19490_
	);
	LUT3 #(
		.INIT('h80)
	) name8978 (
		\wishbone_bd_ram_mem0_reg[182][0]/P0001 ,
		_w11942_,
		_w11986_,
		_w19491_
	);
	LUT3 #(
		.INIT('h80)
	) name8979 (
		\wishbone_bd_ram_mem0_reg[99][0]/P0001 ,
		_w11938_,
		_w11965_,
		_w19492_
	);
	LUT3 #(
		.INIT('h80)
	) name8980 (
		\wishbone_bd_ram_mem0_reg[67][0]/P0001 ,
		_w11938_,
		_w11949_,
		_w19493_
	);
	LUT3 #(
		.INIT('h80)
	) name8981 (
		\wishbone_bd_ram_mem0_reg[116][0]/P0001 ,
		_w11929_,
		_w12012_,
		_w19494_
	);
	LUT4 #(
		.INIT('h0001)
	) name8982 (
		_w19491_,
		_w19492_,
		_w19493_,
		_w19494_,
		_w19495_
	);
	LUT3 #(
		.INIT('h80)
	) name8983 (
		\wishbone_bd_ram_mem0_reg[97][0]/P0001 ,
		_w11965_,
		_w11977_,
		_w19496_
	);
	LUT3 #(
		.INIT('h80)
	) name8984 (
		\wishbone_bd_ram_mem0_reg[65][0]/P0001 ,
		_w11949_,
		_w11977_,
		_w19497_
	);
	LUT3 #(
		.INIT('h80)
	) name8985 (
		\wishbone_bd_ram_mem0_reg[245][0]/P0001 ,
		_w11933_,
		_w11952_,
		_w19498_
	);
	LUT3 #(
		.INIT('h80)
	) name8986 (
		\wishbone_bd_ram_mem0_reg[2][0]/P0001 ,
		_w11932_,
		_w11963_,
		_w19499_
	);
	LUT4 #(
		.INIT('h0001)
	) name8987 (
		_w19496_,
		_w19497_,
		_w19498_,
		_w19499_,
		_w19500_
	);
	LUT4 #(
		.INIT('h8000)
	) name8988 (
		_w19485_,
		_w19490_,
		_w19495_,
		_w19500_,
		_w19501_
	);
	LUT3 #(
		.INIT('h80)
	) name8989 (
		\wishbone_bd_ram_mem0_reg[143][0]/P0001 ,
		_w11955_,
		_w11973_,
		_w19502_
	);
	LUT3 #(
		.INIT('h80)
	) name8990 (
		\wishbone_bd_ram_mem0_reg[254][0]/P0001 ,
		_w11948_,
		_w11952_,
		_w19503_
	);
	LUT3 #(
		.INIT('h80)
	) name8991 (
		\wishbone_bd_ram_mem0_reg[27][0]/P0001 ,
		_w11935_,
		_w11936_,
		_w19504_
	);
	LUT3 #(
		.INIT('h80)
	) name8992 (
		\wishbone_bd_ram_mem0_reg[29][0]/P0001 ,
		_w11935_,
		_w11966_,
		_w19505_
	);
	LUT4 #(
		.INIT('h0001)
	) name8993 (
		_w19502_,
		_w19503_,
		_w19504_,
		_w19505_,
		_w19506_
	);
	LUT3 #(
		.INIT('h80)
	) name8994 (
		\wishbone_bd_ram_mem0_reg[221][0]/P0001 ,
		_w11966_,
		_w11984_,
		_w19507_
	);
	LUT3 #(
		.INIT('h80)
	) name8995 (
		\wishbone_bd_ram_mem0_reg[220][0]/P0001 ,
		_w11954_,
		_w11984_,
		_w19508_
	);
	LUT3 #(
		.INIT('h80)
	) name8996 (
		\wishbone_bd_ram_mem0_reg[136][0]/P0001 ,
		_w11955_,
		_w11990_,
		_w19509_
	);
	LUT3 #(
		.INIT('h80)
	) name8997 (
		\wishbone_bd_ram_mem0_reg[145][0]/P0001 ,
		_w11959_,
		_w11977_,
		_w19510_
	);
	LUT4 #(
		.INIT('h0001)
	) name8998 (
		_w19507_,
		_w19508_,
		_w19509_,
		_w19510_,
		_w19511_
	);
	LUT3 #(
		.INIT('h80)
	) name8999 (
		\wishbone_bd_ram_mem0_reg[172][0]/P0001 ,
		_w11930_,
		_w11954_,
		_w19512_
	);
	LUT3 #(
		.INIT('h80)
	) name9000 (
		\wishbone_bd_ram_mem0_reg[100][0]/P0001 ,
		_w11929_,
		_w11965_,
		_w19513_
	);
	LUT3 #(
		.INIT('h80)
	) name9001 (
		\wishbone_bd_ram_mem0_reg[71][0]/P0001 ,
		_w11949_,
		_w11975_,
		_w19514_
	);
	LUT3 #(
		.INIT('h80)
	) name9002 (
		\wishbone_bd_ram_mem0_reg[35][0]/P0001 ,
		_w11938_,
		_w11957_,
		_w19515_
	);
	LUT4 #(
		.INIT('h0001)
	) name9003 (
		_w19512_,
		_w19513_,
		_w19514_,
		_w19515_,
		_w19516_
	);
	LUT3 #(
		.INIT('h80)
	) name9004 (
		\wishbone_bd_ram_mem0_reg[154][0]/P0001 ,
		_w11944_,
		_w11959_,
		_w19517_
	);
	LUT3 #(
		.INIT('h80)
	) name9005 (
		\wishbone_bd_ram_mem0_reg[83][0]/P0001 ,
		_w11938_,
		_w11972_,
		_w19518_
	);
	LUT3 #(
		.INIT('h80)
	) name9006 (
		\wishbone_bd_ram_mem0_reg[13][0]/P0001 ,
		_w11932_,
		_w11966_,
		_w19519_
	);
	LUT3 #(
		.INIT('h80)
	) name9007 (
		\wishbone_bd_ram_mem0_reg[80][0]/P0001 ,
		_w11941_,
		_w11972_,
		_w19520_
	);
	LUT4 #(
		.INIT('h0001)
	) name9008 (
		_w19517_,
		_w19518_,
		_w19519_,
		_w19520_,
		_w19521_
	);
	LUT4 #(
		.INIT('h8000)
	) name9009 (
		_w19506_,
		_w19511_,
		_w19516_,
		_w19521_,
		_w19522_
	);
	LUT4 #(
		.INIT('h8000)
	) name9010 (
		_w19459_,
		_w19480_,
		_w19501_,
		_w19522_,
		_w19523_
	);
	LUT4 #(
		.INIT('h8000)
	) name9011 (
		_w19268_,
		_w19353_,
		_w19438_,
		_w19523_,
		_w19524_
	);
	LUT3 #(
		.INIT('hce)
	) name9012 (
		_w19180_,
		_w19183_,
		_w19524_,
		_w19525_
	);
	LUT4 #(
		.INIT('h70f0)
	) name9013 (
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w19526_
	);
	LUT3 #(
		.INIT('hf2)
	) name9014 (
		_w19180_,
		_w19524_,
		_w19526_,
		_w19527_
	);
	LUT3 #(
		.INIT('h70)
	) name9015 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w19528_
	);
	LUT2 #(
		.INIT('h4)
	) name9016 (
		_w15303_,
		_w19528_,
		_w19529_
	);
	LUT3 #(
		.INIT('hf4)
	) name9017 (
		_w14151_,
		_w19180_,
		_w19529_,
		_w19530_
	);
	LUT3 #(
		.INIT('h80)
	) name9018 (
		\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 ,
		_w18753_,
		_w18754_,
		_w19531_
	);
	LUT4 #(
		.INIT('h0008)
	) name9019 (
		\ethreg1_RXHASH0_2_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19532_
	);
	LUT3 #(
		.INIT('h80)
	) name9020 (
		_w18757_,
		_w18758_,
		_w19532_,
		_w19533_
	);
	LUT4 #(
		.INIT('h0008)
	) name9021 (
		\ethreg1_RXHASH1_2_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19534_
	);
	LUT3 #(
		.INIT('h80)
	) name9022 (
		_w18757_,
		_w18762_,
		_w19534_,
		_w19535_
	);
	LUT4 #(
		.INIT('h0002)
	) name9023 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19536_
	);
	LUT3 #(
		.INIT('h80)
	) name9024 (
		_w18757_,
		_w18758_,
		_w19536_,
		_w19537_
	);
	LUT4 #(
		.INIT('h0002)
	) name9025 (
		_w18752_,
		_w19533_,
		_w19535_,
		_w19537_,
		_w19538_
	);
	LUT3 #(
		.INIT('h8a)
	) name9026 (
		_w18752_,
		_w19531_,
		_w19538_,
		_w19539_
	);
	LUT3 #(
		.INIT('h45)
	) name9027 (
		wb_rst_i_pad,
		_w19531_,
		_w19538_,
		_w19540_
	);
	LUT3 #(
		.INIT('hdc)
	) name9028 (
		_w18401_,
		_w19539_,
		_w19540_,
		_w19541_
	);
	LUT3 #(
		.INIT('h80)
	) name9029 (
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		_w18753_,
		_w18754_,
		_w19542_
	);
	LUT4 #(
		.INIT('h0008)
	) name9030 (
		\ethreg1_RXHASH0_3_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19543_
	);
	LUT3 #(
		.INIT('h80)
	) name9031 (
		_w18757_,
		_w18758_,
		_w19543_,
		_w19544_
	);
	LUT4 #(
		.INIT('h0008)
	) name9032 (
		\ethreg1_RXHASH1_3_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19545_
	);
	LUT3 #(
		.INIT('h80)
	) name9033 (
		_w18757_,
		_w18762_,
		_w19545_,
		_w19546_
	);
	LUT4 #(
		.INIT('h0002)
	) name9034 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19547_
	);
	LUT3 #(
		.INIT('h80)
	) name9035 (
		_w18757_,
		_w18758_,
		_w19547_,
		_w19548_
	);
	LUT4 #(
		.INIT('h0002)
	) name9036 (
		_w18752_,
		_w19544_,
		_w19546_,
		_w19548_,
		_w19549_
	);
	LUT3 #(
		.INIT('h8a)
	) name9037 (
		_w18752_,
		_w19542_,
		_w19549_,
		_w19550_
	);
	LUT3 #(
		.INIT('h45)
	) name9038 (
		wb_rst_i_pad,
		_w19542_,
		_w19549_,
		_w19551_
	);
	LUT3 #(
		.INIT('hdc)
	) name9039 (
		_w13397_,
		_w19550_,
		_w19551_,
		_w19552_
	);
	LUT3 #(
		.INIT('h80)
	) name9040 (
		\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 ,
		_w18753_,
		_w18754_,
		_w19553_
	);
	LUT4 #(
		.INIT('h0008)
	) name9041 (
		\ethreg1_RXHASH0_3_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19554_
	);
	LUT3 #(
		.INIT('h80)
	) name9042 (
		_w18757_,
		_w18758_,
		_w19554_,
		_w19555_
	);
	LUT4 #(
		.INIT('h0008)
	) name9043 (
		\ethreg1_RXHASH1_3_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19556_
	);
	LUT3 #(
		.INIT('h80)
	) name9044 (
		_w18757_,
		_w18762_,
		_w19556_,
		_w19557_
	);
	LUT4 #(
		.INIT('h0002)
	) name9045 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19558_
	);
	LUT3 #(
		.INIT('h80)
	) name9046 (
		_w18757_,
		_w18758_,
		_w19558_,
		_w19559_
	);
	LUT4 #(
		.INIT('h0002)
	) name9047 (
		_w18752_,
		_w19555_,
		_w19557_,
		_w19559_,
		_w19560_
	);
	LUT3 #(
		.INIT('h8a)
	) name9048 (
		_w18752_,
		_w19553_,
		_w19560_,
		_w19561_
	);
	LUT3 #(
		.INIT('h45)
	) name9049 (
		wb_rst_i_pad,
		_w19553_,
		_w19560_,
		_w19562_
	);
	LUT3 #(
		.INIT('hdc)
	) name9050 (
		_w15222_,
		_w19561_,
		_w19562_,
		_w19563_
	);
	LUT3 #(
		.INIT('h80)
	) name9051 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		_w18753_,
		_w18754_,
		_w19564_
	);
	LUT4 #(
		.INIT('h0008)
	) name9052 (
		\ethreg1_RXHASH0_3_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19565_
	);
	LUT3 #(
		.INIT('h80)
	) name9053 (
		_w18757_,
		_w18758_,
		_w19565_,
		_w19566_
	);
	LUT4 #(
		.INIT('h0008)
	) name9054 (
		\ethreg1_RXHASH1_3_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19567_
	);
	LUT3 #(
		.INIT('h80)
	) name9055 (
		_w18757_,
		_w18762_,
		_w19567_,
		_w19568_
	);
	LUT4 #(
		.INIT('h0002)
	) name9056 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19569_
	);
	LUT3 #(
		.INIT('h80)
	) name9057 (
		_w18757_,
		_w18758_,
		_w19569_,
		_w19570_
	);
	LUT4 #(
		.INIT('h0002)
	) name9058 (
		_w18752_,
		_w19566_,
		_w19568_,
		_w19570_,
		_w19571_
	);
	LUT3 #(
		.INIT('h8a)
	) name9059 (
		_w18752_,
		_w19564_,
		_w19571_,
		_w19572_
	);
	LUT3 #(
		.INIT('h45)
	) name9060 (
		wb_rst_i_pad,
		_w19564_,
		_w19571_,
		_w19573_
	);
	LUT3 #(
		.INIT('hdc)
	) name9061 (
		_w14872_,
		_w19572_,
		_w19573_,
		_w19574_
	);
	LUT3 #(
		.INIT('h80)
	) name9062 (
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		_w18753_,
		_w18754_,
		_w19575_
	);
	LUT4 #(
		.INIT('h0008)
	) name9063 (
		\ethreg1_RXHASH0_3_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19576_
	);
	LUT3 #(
		.INIT('h80)
	) name9064 (
		_w18757_,
		_w18758_,
		_w19576_,
		_w19577_
	);
	LUT4 #(
		.INIT('h0008)
	) name9065 (
		\ethreg1_RXHASH1_3_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19578_
	);
	LUT3 #(
		.INIT('h80)
	) name9066 (
		_w18757_,
		_w18762_,
		_w19578_,
		_w19579_
	);
	LUT4 #(
		.INIT('h0002)
	) name9067 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19580_
	);
	LUT3 #(
		.INIT('h80)
	) name9068 (
		_w18757_,
		_w18758_,
		_w19580_,
		_w19581_
	);
	LUT4 #(
		.INIT('h0002)
	) name9069 (
		_w18752_,
		_w19577_,
		_w19579_,
		_w19581_,
		_w19582_
	);
	LUT3 #(
		.INIT('h8a)
	) name9070 (
		_w18752_,
		_w19575_,
		_w19582_,
		_w19583_
	);
	LUT3 #(
		.INIT('h45)
	) name9071 (
		wb_rst_i_pad,
		_w19575_,
		_w19582_,
		_w19584_
	);
	LUT3 #(
		.INIT('hdc)
	) name9072 (
		_w17356_,
		_w19583_,
		_w19584_,
		_w19585_
	);
	LUT3 #(
		.INIT('h80)
	) name9073 (
		\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 ,
		_w18753_,
		_w18754_,
		_w19586_
	);
	LUT4 #(
		.INIT('h0008)
	) name9074 (
		\ethreg1_RXHASH0_3_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19587_
	);
	LUT3 #(
		.INIT('h80)
	) name9075 (
		_w18757_,
		_w18758_,
		_w19587_,
		_w19588_
	);
	LUT4 #(
		.INIT('h0008)
	) name9076 (
		\ethreg1_RXHASH1_3_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19589_
	);
	LUT3 #(
		.INIT('h80)
	) name9077 (
		_w18757_,
		_w18762_,
		_w19589_,
		_w19590_
	);
	LUT4 #(
		.INIT('h0002)
	) name9078 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19591_
	);
	LUT3 #(
		.INIT('h80)
	) name9079 (
		_w18757_,
		_w18758_,
		_w19591_,
		_w19592_
	);
	LUT4 #(
		.INIT('h0002)
	) name9080 (
		_w18752_,
		_w19588_,
		_w19590_,
		_w19592_,
		_w19593_
	);
	LUT3 #(
		.INIT('h8a)
	) name9081 (
		_w18752_,
		_w19586_,
		_w19593_,
		_w19594_
	);
	LUT3 #(
		.INIT('h45)
	) name9082 (
		wb_rst_i_pad,
		_w19586_,
		_w19593_,
		_w19595_
	);
	LUT3 #(
		.INIT('hdc)
	) name9083 (
		_w12301_,
		_w19594_,
		_w19595_,
		_w19596_
	);
	LUT3 #(
		.INIT('h80)
	) name9084 (
		\ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131 ,
		_w18753_,
		_w18754_,
		_w19597_
	);
	LUT4 #(
		.INIT('h0008)
	) name9085 (
		\ethreg1_RXHASH0_3_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19598_
	);
	LUT3 #(
		.INIT('h80)
	) name9086 (
		_w18757_,
		_w18758_,
		_w19598_,
		_w19599_
	);
	LUT4 #(
		.INIT('h0008)
	) name9087 (
		\ethreg1_RXHASH1_3_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19600_
	);
	LUT3 #(
		.INIT('h80)
	) name9088 (
		_w18757_,
		_w18762_,
		_w19600_,
		_w19601_
	);
	LUT4 #(
		.INIT('h0002)
	) name9089 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19602_
	);
	LUT3 #(
		.INIT('h80)
	) name9090 (
		_w18757_,
		_w18758_,
		_w19602_,
		_w19603_
	);
	LUT4 #(
		.INIT('h0002)
	) name9091 (
		_w18752_,
		_w19599_,
		_w19601_,
		_w19603_,
		_w19604_
	);
	LUT3 #(
		.INIT('h8a)
	) name9092 (
		_w18752_,
		_w19597_,
		_w19604_,
		_w19605_
	);
	LUT3 #(
		.INIT('h45)
	) name9093 (
		wb_rst_i_pad,
		_w19597_,
		_w19604_,
		_w19606_
	);
	LUT3 #(
		.INIT('hdc)
	) name9094 (
		_w12668_,
		_w19605_,
		_w19606_,
		_w19607_
	);
	LUT3 #(
		.INIT('h20)
	) name9095 (
		m_wb_we_o_pad,
		_w11890_,
		_w11900_,
		_w19608_
	);
	LUT2 #(
		.INIT('hd)
	) name9096 (
		_w11906_,
		_w19608_,
		_w19609_
	);
	LUT3 #(
		.INIT('h80)
	) name9097 (
		\ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131 ,
		_w18753_,
		_w18754_,
		_w19610_
	);
	LUT4 #(
		.INIT('h0008)
	) name9098 (
		\ethreg1_RXHASH0_3_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19611_
	);
	LUT3 #(
		.INIT('h80)
	) name9099 (
		_w18757_,
		_w18758_,
		_w19611_,
		_w19612_
	);
	LUT4 #(
		.INIT('h0008)
	) name9100 (
		\ethreg1_RXHASH1_3_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19613_
	);
	LUT3 #(
		.INIT('h80)
	) name9101 (
		_w18757_,
		_w18762_,
		_w19613_,
		_w19614_
	);
	LUT4 #(
		.INIT('h0002)
	) name9102 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19615_
	);
	LUT3 #(
		.INIT('h80)
	) name9103 (
		_w18757_,
		_w18758_,
		_w19615_,
		_w19616_
	);
	LUT4 #(
		.INIT('h0002)
	) name9104 (
		_w18752_,
		_w19612_,
		_w19614_,
		_w19616_,
		_w19617_
	);
	LUT3 #(
		.INIT('h8a)
	) name9105 (
		_w18752_,
		_w19610_,
		_w19617_,
		_w19618_
	);
	LUT3 #(
		.INIT('h45)
	) name9106 (
		wb_rst_i_pad,
		_w19610_,
		_w19617_,
		_w19619_
	);
	LUT3 #(
		.INIT('hdc)
	) name9107 (
		_w13016_,
		_w19618_,
		_w19619_,
		_w19620_
	);
	LUT3 #(
		.INIT('h80)
	) name9108 (
		\ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131 ,
		_w18753_,
		_w18754_,
		_w19621_
	);
	LUT4 #(
		.INIT('h0008)
	) name9109 (
		\ethreg1_RXHASH0_3_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19622_
	);
	LUT3 #(
		.INIT('h80)
	) name9110 (
		_w18757_,
		_w18758_,
		_w19622_,
		_w19623_
	);
	LUT4 #(
		.INIT('h0008)
	) name9111 (
		\ethreg1_RXHASH1_3_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19624_
	);
	LUT3 #(
		.INIT('h80)
	) name9112 (
		_w18757_,
		_w18762_,
		_w19624_,
		_w19625_
	);
	LUT4 #(
		.INIT('h0002)
	) name9113 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19626_
	);
	LUT3 #(
		.INIT('h80)
	) name9114 (
		_w18757_,
		_w18758_,
		_w19626_,
		_w19627_
	);
	LUT4 #(
		.INIT('h0002)
	) name9115 (
		_w18752_,
		_w19623_,
		_w19625_,
		_w19627_,
		_w19628_
	);
	LUT3 #(
		.INIT('h8a)
	) name9116 (
		_w18752_,
		_w19621_,
		_w19628_,
		_w19629_
	);
	LUT3 #(
		.INIT('h45)
	) name9117 (
		wb_rst_i_pad,
		_w19621_,
		_w19628_,
		_w19630_
	);
	LUT3 #(
		.INIT('hdc)
	) name9118 (
		_w16469_,
		_w19629_,
		_w19630_,
		_w19631_
	);
	LUT4 #(
		.INIT('h0008)
	) name9119 (
		\ethreg1_RXHASH1_0_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19632_
	);
	LUT3 #(
		.INIT('h80)
	) name9120 (
		_w18757_,
		_w18762_,
		_w19632_,
		_w19633_
	);
	LUT4 #(
		.INIT('h0002)
	) name9121 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19634_
	);
	LUT3 #(
		.INIT('h80)
	) name9122 (
		_w18757_,
		_w18758_,
		_w19634_,
		_w19635_
	);
	LUT3 #(
		.INIT('h80)
	) name9123 (
		\ethreg1_MIIRX_DATA_DataOut_reg[3]/NET0131 ,
		_w18785_,
		_w18786_,
		_w19636_
	);
	LUT3 #(
		.INIT('h80)
	) name9124 (
		\ethreg1_MODER_0_DataOut_reg[3]/NET0131 ,
		_w18800_,
		_w18801_,
		_w19637_
	);
	LUT4 #(
		.INIT('h0001)
	) name9125 (
		_w19633_,
		_w19635_,
		_w19636_,
		_w19637_,
		_w19638_
	);
	LUT3 #(
		.INIT('h80)
	) name9126 (
		\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 ,
		_w18753_,
		_w18754_,
		_w19639_
	);
	LUT2 #(
		.INIT('h8)
	) name9127 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		_w19640_
	);
	LUT4 #(
		.INIT('h0080)
	) name9128 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19641_
	);
	LUT2 #(
		.INIT('h8)
	) name9129 (
		_w18753_,
		_w19641_,
		_w19642_
	);
	LUT3 #(
		.INIT('h80)
	) name9130 (
		\ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131 ,
		_w18753_,
		_w19641_,
		_w19643_
	);
	LUT2 #(
		.INIT('h1)
	) name9131 (
		_w19639_,
		_w19643_,
		_w19644_
	);
	LUT2 #(
		.INIT('h8)
	) name9132 (
		_w19638_,
		_w19644_,
		_w19645_
	);
	LUT4 #(
		.INIT('h0002)
	) name9133 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[6]_pad ,
		\wb_adr_i[8]_pad ,
		_w19646_
	);
	LUT3 #(
		.INIT('h80)
	) name9134 (
		\ethreg1_irq_rxe_reg/NET0131 ,
		_w18800_,
		_w19646_,
		_w19647_
	);
	LUT4 #(
		.INIT('h0020)
	) name9135 (
		\ethreg1_TXCTRL_0_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19648_
	);
	LUT3 #(
		.INIT('h80)
	) name9136 (
		_w18757_,
		_w18758_,
		_w19648_,
		_w19649_
	);
	LUT3 #(
		.INIT('h80)
	) name9137 (
		\ethreg1_IPGR1_0_DataOut_reg[3]/NET0131 ,
		_w18785_,
		_w18800_,
		_w19650_
	);
	LUT3 #(
		.INIT('h80)
	) name9138 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[3]/NET0131 ,
		_w18785_,
		_w18798_,
		_w19651_
	);
	LUT4 #(
		.INIT('h0001)
	) name9139 (
		_w19647_,
		_w19649_,
		_w19650_,
		_w19651_,
		_w19652_
	);
	LUT4 #(
		.INIT('h0002)
	) name9140 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19653_
	);
	LUT3 #(
		.INIT('h80)
	) name9141 (
		_w18757_,
		_w18762_,
		_w19653_,
		_w19654_
	);
	LUT4 #(
		.INIT('h0002)
	) name9142 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[5]_pad ,
		\wb_adr_i[7]_pad ,
		\wb_adr_i[9]_pad ,
		_w19655_
	);
	LUT3 #(
		.INIT('h80)
	) name9143 (
		\ethreg1_INT_MASK_0_DataOut_reg[3]/NET0131 ,
		_w18801_,
		_w19655_,
		_w19656_
	);
	LUT3 #(
		.INIT('h80)
	) name9144 (
		\ethreg1_IPGR2_0_DataOut_reg[3]/NET0131 ,
		_w18800_,
		_w18805_,
		_w19657_
	);
	LUT3 #(
		.INIT('h80)
	) name9145 (
		\ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131 ,
		_w18786_,
		_w18801_,
		_w19658_
	);
	LUT4 #(
		.INIT('h0001)
	) name9146 (
		_w19654_,
		_w19656_,
		_w19657_,
		_w19658_,
		_w19659_
	);
	LUT3 #(
		.INIT('h80)
	) name9147 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[3]/NET0131 ,
		_w18798_,
		_w18801_,
		_w19660_
	);
	LUT3 #(
		.INIT('h80)
	) name9148 (
		\ethreg1_IPGT_0_DataOut_reg[3]/NET0131 ,
		_w19646_,
		_w19655_,
		_w19661_
	);
	LUT3 #(
		.INIT('h80)
	) name9149 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[3]/NET0131 ,
		_w18798_,
		_w18805_,
		_w19662_
	);
	LUT4 #(
		.INIT('h0008)
	) name9150 (
		\ethreg1_RXHASH0_0_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w19663_
	);
	LUT3 #(
		.INIT('h80)
	) name9151 (
		_w18757_,
		_w18758_,
		_w19663_,
		_w19664_
	);
	LUT4 #(
		.INIT('h0001)
	) name9152 (
		_w19660_,
		_w19661_,
		_w19662_,
		_w19664_,
		_w19665_
	);
	LUT4 #(
		.INIT('h8000)
	) name9153 (
		_w18752_,
		_w19652_,
		_w19659_,
		_w19665_,
		_w19666_
	);
	LUT3 #(
		.INIT('h2a)
	) name9154 (
		_w18752_,
		_w19645_,
		_w19666_,
		_w19667_
	);
	LUT3 #(
		.INIT('h80)
	) name9155 (
		\wishbone_bd_ram_mem0_reg[209][3]/P0001 ,
		_w11977_,
		_w11984_,
		_w19668_
	);
	LUT3 #(
		.INIT('h80)
	) name9156 (
		\wishbone_bd_ram_mem0_reg[12][3]/P0001 ,
		_w11932_,
		_w11954_,
		_w19669_
	);
	LUT3 #(
		.INIT('h80)
	) name9157 (
		\wishbone_bd_ram_mem0_reg[37][3]/P0001 ,
		_w11933_,
		_w11957_,
		_w19670_
	);
	LUT3 #(
		.INIT('h80)
	) name9158 (
		\wishbone_bd_ram_mem0_reg[162][3]/P0001 ,
		_w11930_,
		_w11963_,
		_w19671_
	);
	LUT4 #(
		.INIT('h0001)
	) name9159 (
		_w19668_,
		_w19669_,
		_w19670_,
		_w19671_,
		_w19672_
	);
	LUT3 #(
		.INIT('h80)
	) name9160 (
		\wishbone_bd_ram_mem0_reg[94][3]/P0001 ,
		_w11948_,
		_w11972_,
		_w19673_
	);
	LUT3 #(
		.INIT('h80)
	) name9161 (
		\wishbone_bd_ram_mem0_reg[97][3]/P0001 ,
		_w11965_,
		_w11977_,
		_w19674_
	);
	LUT3 #(
		.INIT('h80)
	) name9162 (
		\wishbone_bd_ram_mem0_reg[128][3]/P0001 ,
		_w11941_,
		_w11955_,
		_w19675_
	);
	LUT3 #(
		.INIT('h80)
	) name9163 (
		\wishbone_bd_ram_mem0_reg[175][3]/P0001 ,
		_w11930_,
		_w11973_,
		_w19676_
	);
	LUT4 #(
		.INIT('h0001)
	) name9164 (
		_w19673_,
		_w19674_,
		_w19675_,
		_w19676_,
		_w19677_
	);
	LUT3 #(
		.INIT('h80)
	) name9165 (
		\wishbone_bd_ram_mem0_reg[187][3]/P0001 ,
		_w11936_,
		_w11942_,
		_w19678_
	);
	LUT3 #(
		.INIT('h80)
	) name9166 (
		\wishbone_bd_ram_mem0_reg[197][3]/P0001 ,
		_w11933_,
		_w11945_,
		_w19679_
	);
	LUT3 #(
		.INIT('h80)
	) name9167 (
		\wishbone_bd_ram_mem0_reg[102][3]/P0001 ,
		_w11965_,
		_w11986_,
		_w19680_
	);
	LUT3 #(
		.INIT('h80)
	) name9168 (
		\wishbone_bd_ram_mem0_reg[228][3]/P0001 ,
		_w11929_,
		_w11982_,
		_w19681_
	);
	LUT4 #(
		.INIT('h0001)
	) name9169 (
		_w19678_,
		_w19679_,
		_w19680_,
		_w19681_,
		_w19682_
	);
	LUT3 #(
		.INIT('h80)
	) name9170 (
		\wishbone_bd_ram_mem0_reg[11][3]/P0001 ,
		_w11932_,
		_w11936_,
		_w19683_
	);
	LUT3 #(
		.INIT('h80)
	) name9171 (
		\wishbone_bd_ram_mem0_reg[246][3]/P0001 ,
		_w11952_,
		_w11986_,
		_w19684_
	);
	LUT3 #(
		.INIT('h80)
	) name9172 (
		\wishbone_bd_ram_mem0_reg[115][3]/P0001 ,
		_w11938_,
		_w12012_,
		_w19685_
	);
	LUT3 #(
		.INIT('h80)
	) name9173 (
		\wishbone_bd_ram_mem0_reg[156][3]/P0001 ,
		_w11954_,
		_w11959_,
		_w19686_
	);
	LUT4 #(
		.INIT('h0001)
	) name9174 (
		_w19683_,
		_w19684_,
		_w19685_,
		_w19686_,
		_w19687_
	);
	LUT4 #(
		.INIT('h8000)
	) name9175 (
		_w19672_,
		_w19677_,
		_w19682_,
		_w19687_,
		_w19688_
	);
	LUT3 #(
		.INIT('h80)
	) name9176 (
		\wishbone_bd_ram_mem0_reg[144][3]/P0001 ,
		_w11941_,
		_w11959_,
		_w19689_
	);
	LUT3 #(
		.INIT('h80)
	) name9177 (
		\wishbone_bd_ram_mem0_reg[153][3]/P0001 ,
		_w11959_,
		_w11968_,
		_w19690_
	);
	LUT3 #(
		.INIT('h80)
	) name9178 (
		\wishbone_bd_ram_mem0_reg[3][3]/P0001 ,
		_w11932_,
		_w11938_,
		_w19691_
	);
	LUT3 #(
		.INIT('h80)
	) name9179 (
		\wishbone_bd_ram_mem0_reg[122][3]/P0001 ,
		_w11944_,
		_w12012_,
		_w19692_
	);
	LUT4 #(
		.INIT('h0001)
	) name9180 (
		_w19689_,
		_w19690_,
		_w19691_,
		_w19692_,
		_w19693_
	);
	LUT3 #(
		.INIT('h80)
	) name9181 (
		\wishbone_bd_ram_mem0_reg[225][3]/P0001 ,
		_w11977_,
		_w11982_,
		_w19694_
	);
	LUT3 #(
		.INIT('h80)
	) name9182 (
		\wishbone_bd_ram_mem0_reg[179][3]/P0001 ,
		_w11938_,
		_w11942_,
		_w19695_
	);
	LUT3 #(
		.INIT('h80)
	) name9183 (
		\wishbone_bd_ram_mem0_reg[216][3]/P0001 ,
		_w11984_,
		_w11990_,
		_w19696_
	);
	LUT3 #(
		.INIT('h80)
	) name9184 (
		\wishbone_bd_ram_mem0_reg[30][3]/P0001 ,
		_w11935_,
		_w11948_,
		_w19697_
	);
	LUT4 #(
		.INIT('h0001)
	) name9185 (
		_w19694_,
		_w19695_,
		_w19696_,
		_w19697_,
		_w19698_
	);
	LUT3 #(
		.INIT('h80)
	) name9186 (
		\wishbone_bd_ram_mem0_reg[43][3]/P0001 ,
		_w11936_,
		_w11957_,
		_w19699_
	);
	LUT3 #(
		.INIT('h80)
	) name9187 (
		\wishbone_bd_ram_mem0_reg[194][3]/P0001 ,
		_w11945_,
		_w11963_,
		_w19700_
	);
	LUT3 #(
		.INIT('h80)
	) name9188 (
		\wishbone_bd_ram_mem0_reg[229][3]/P0001 ,
		_w11933_,
		_w11982_,
		_w19701_
	);
	LUT3 #(
		.INIT('h80)
	) name9189 (
		\wishbone_bd_ram_mem0_reg[21][3]/P0001 ,
		_w11933_,
		_w11935_,
		_w19702_
	);
	LUT4 #(
		.INIT('h0001)
	) name9190 (
		_w19699_,
		_w19700_,
		_w19701_,
		_w19702_,
		_w19703_
	);
	LUT3 #(
		.INIT('h80)
	) name9191 (
		\wishbone_bd_ram_mem0_reg[14][3]/P0001 ,
		_w11932_,
		_w11948_,
		_w19704_
	);
	LUT3 #(
		.INIT('h80)
	) name9192 (
		\wishbone_bd_ram_mem0_reg[49][3]/P0001 ,
		_w11977_,
		_w11979_,
		_w19705_
	);
	LUT3 #(
		.INIT('h80)
	) name9193 (
		\wishbone_bd_ram_mem0_reg[231][3]/P0001 ,
		_w11975_,
		_w11982_,
		_w19706_
	);
	LUT3 #(
		.INIT('h80)
	) name9194 (
		\wishbone_bd_ram_mem0_reg[226][3]/P0001 ,
		_w11963_,
		_w11982_,
		_w19707_
	);
	LUT4 #(
		.INIT('h0001)
	) name9195 (
		_w19704_,
		_w19705_,
		_w19706_,
		_w19707_,
		_w19708_
	);
	LUT4 #(
		.INIT('h8000)
	) name9196 (
		_w19693_,
		_w19698_,
		_w19703_,
		_w19708_,
		_w19709_
	);
	LUT3 #(
		.INIT('h80)
	) name9197 (
		\wishbone_bd_ram_mem0_reg[247][3]/P0001 ,
		_w11952_,
		_w11975_,
		_w19710_
	);
	LUT3 #(
		.INIT('h80)
	) name9198 (
		\wishbone_bd_ram_mem0_reg[93][3]/P0001 ,
		_w11966_,
		_w11972_,
		_w19711_
	);
	LUT3 #(
		.INIT('h80)
	) name9199 (
		\wishbone_bd_ram_mem0_reg[48][3]/P0001 ,
		_w11941_,
		_w11979_,
		_w19712_
	);
	LUT3 #(
		.INIT('h80)
	) name9200 (
		\wishbone_bd_ram_mem0_reg[96][3]/P0001 ,
		_w11941_,
		_w11965_,
		_w19713_
	);
	LUT4 #(
		.INIT('h0001)
	) name9201 (
		_w19710_,
		_w19711_,
		_w19712_,
		_w19713_,
		_w19714_
	);
	LUT3 #(
		.INIT('h80)
	) name9202 (
		\wishbone_bd_ram_mem0_reg[211][3]/P0001 ,
		_w11938_,
		_w11984_,
		_w19715_
	);
	LUT3 #(
		.INIT('h80)
	) name9203 (
		\wishbone_bd_ram_mem0_reg[106][3]/P0001 ,
		_w11944_,
		_w11965_,
		_w19716_
	);
	LUT3 #(
		.INIT('h80)
	) name9204 (
		\wishbone_bd_ram_mem0_reg[190][3]/P0001 ,
		_w11942_,
		_w11948_,
		_w19717_
	);
	LUT3 #(
		.INIT('h80)
	) name9205 (
		\wishbone_bd_ram_mem0_reg[108][3]/P0001 ,
		_w11954_,
		_w11965_,
		_w19718_
	);
	LUT4 #(
		.INIT('h0001)
	) name9206 (
		_w19715_,
		_w19716_,
		_w19717_,
		_w19718_,
		_w19719_
	);
	LUT3 #(
		.INIT('h80)
	) name9207 (
		\wishbone_bd_ram_mem0_reg[180][3]/P0001 ,
		_w11929_,
		_w11942_,
		_w19720_
	);
	LUT3 #(
		.INIT('h80)
	) name9208 (
		\wishbone_bd_ram_mem0_reg[109][3]/P0001 ,
		_w11965_,
		_w11966_,
		_w19721_
	);
	LUT3 #(
		.INIT('h80)
	) name9209 (
		\wishbone_bd_ram_mem0_reg[117][3]/P0001 ,
		_w11933_,
		_w12012_,
		_w19722_
	);
	LUT3 #(
		.INIT('h80)
	) name9210 (
		\wishbone_bd_ram_mem0_reg[184][3]/P0001 ,
		_w11942_,
		_w11990_,
		_w19723_
	);
	LUT4 #(
		.INIT('h0001)
	) name9211 (
		_w19720_,
		_w19721_,
		_w19722_,
		_w19723_,
		_w19724_
	);
	LUT3 #(
		.INIT('h80)
	) name9212 (
		\wishbone_bd_ram_mem0_reg[111][3]/P0001 ,
		_w11965_,
		_w11973_,
		_w19725_
	);
	LUT3 #(
		.INIT('h80)
	) name9213 (
		\wishbone_bd_ram_mem0_reg[215][3]/P0001 ,
		_w11975_,
		_w11984_,
		_w19726_
	);
	LUT3 #(
		.INIT('h80)
	) name9214 (
		\wishbone_bd_ram_mem0_reg[119][3]/P0001 ,
		_w11975_,
		_w12012_,
		_w19727_
	);
	LUT3 #(
		.INIT('h80)
	) name9215 (
		\wishbone_bd_ram_mem0_reg[181][3]/P0001 ,
		_w11933_,
		_w11942_,
		_w19728_
	);
	LUT4 #(
		.INIT('h0001)
	) name9216 (
		_w19725_,
		_w19726_,
		_w19727_,
		_w19728_,
		_w19729_
	);
	LUT4 #(
		.INIT('h8000)
	) name9217 (
		_w19714_,
		_w19719_,
		_w19724_,
		_w19729_,
		_w19730_
	);
	LUT3 #(
		.INIT('h80)
	) name9218 (
		\wishbone_bd_ram_mem0_reg[137][3]/P0001 ,
		_w11955_,
		_w11968_,
		_w19731_
	);
	LUT3 #(
		.INIT('h80)
	) name9219 (
		\wishbone_bd_ram_mem0_reg[174][3]/P0001 ,
		_w11930_,
		_w11948_,
		_w19732_
	);
	LUT3 #(
		.INIT('h80)
	) name9220 (
		\wishbone_bd_ram_mem0_reg[164][3]/P0001 ,
		_w11929_,
		_w11930_,
		_w19733_
	);
	LUT3 #(
		.INIT('h80)
	) name9221 (
		\wishbone_bd_ram_mem0_reg[146][3]/P0001 ,
		_w11959_,
		_w11963_,
		_w19734_
	);
	LUT4 #(
		.INIT('h0001)
	) name9222 (
		_w19731_,
		_w19732_,
		_w19733_,
		_w19734_,
		_w19735_
	);
	LUT3 #(
		.INIT('h80)
	) name9223 (
		\wishbone_bd_ram_mem0_reg[239][3]/P0001 ,
		_w11973_,
		_w11982_,
		_w19736_
	);
	LUT3 #(
		.INIT('h80)
	) name9224 (
		\wishbone_bd_ram_mem0_reg[223][3]/P0001 ,
		_w11973_,
		_w11984_,
		_w19737_
	);
	LUT3 #(
		.INIT('h80)
	) name9225 (
		\wishbone_bd_ram_mem0_reg[149][3]/P0001 ,
		_w11933_,
		_w11959_,
		_w19738_
	);
	LUT3 #(
		.INIT('h80)
	) name9226 (
		\wishbone_bd_ram_mem0_reg[4][3]/P0001 ,
		_w11929_,
		_w11932_,
		_w19739_
	);
	LUT4 #(
		.INIT('h0001)
	) name9227 (
		_w19736_,
		_w19737_,
		_w19738_,
		_w19739_,
		_w19740_
	);
	LUT3 #(
		.INIT('h80)
	) name9228 (
		\wishbone_bd_ram_mem0_reg[133][3]/P0001 ,
		_w11933_,
		_w11955_,
		_w19741_
	);
	LUT3 #(
		.INIT('h80)
	) name9229 (
		\wishbone_bd_ram_mem0_reg[157][3]/P0001 ,
		_w11959_,
		_w11966_,
		_w19742_
	);
	LUT3 #(
		.INIT('h80)
	) name9230 (
		\wishbone_bd_ram_mem0_reg[123][3]/P0001 ,
		_w11936_,
		_w12012_,
		_w19743_
	);
	LUT3 #(
		.INIT('h80)
	) name9231 (
		\wishbone_bd_ram_mem0_reg[38][3]/P0001 ,
		_w11957_,
		_w11986_,
		_w19744_
	);
	LUT4 #(
		.INIT('h0001)
	) name9232 (
		_w19741_,
		_w19742_,
		_w19743_,
		_w19744_,
		_w19745_
	);
	LUT3 #(
		.INIT('h80)
	) name9233 (
		\wishbone_bd_ram_mem0_reg[105][3]/P0001 ,
		_w11965_,
		_w11968_,
		_w19746_
	);
	LUT3 #(
		.INIT('h80)
	) name9234 (
		\wishbone_bd_ram_mem0_reg[74][3]/P0001 ,
		_w11944_,
		_w11949_,
		_w19747_
	);
	LUT3 #(
		.INIT('h80)
	) name9235 (
		\wishbone_bd_ram_mem0_reg[44][3]/P0001 ,
		_w11954_,
		_w11957_,
		_w19748_
	);
	LUT3 #(
		.INIT('h80)
	) name9236 (
		\wishbone_bd_ram_mem0_reg[120][3]/P0001 ,
		_w11990_,
		_w12012_,
		_w19749_
	);
	LUT4 #(
		.INIT('h0001)
	) name9237 (
		_w19746_,
		_w19747_,
		_w19748_,
		_w19749_,
		_w19750_
	);
	LUT4 #(
		.INIT('h8000)
	) name9238 (
		_w19735_,
		_w19740_,
		_w19745_,
		_w19750_,
		_w19751_
	);
	LUT4 #(
		.INIT('h8000)
	) name9239 (
		_w19688_,
		_w19709_,
		_w19730_,
		_w19751_,
		_w19752_
	);
	LUT3 #(
		.INIT('h80)
	) name9240 (
		\wishbone_bd_ram_mem0_reg[148][3]/P0001 ,
		_w11929_,
		_w11959_,
		_w19753_
	);
	LUT3 #(
		.INIT('h80)
	) name9241 (
		\wishbone_bd_ram_mem0_reg[202][3]/P0001 ,
		_w11944_,
		_w11945_,
		_w19754_
	);
	LUT3 #(
		.INIT('h80)
	) name9242 (
		\wishbone_bd_ram_mem0_reg[244][3]/P0001 ,
		_w11929_,
		_w11952_,
		_w19755_
	);
	LUT3 #(
		.INIT('h80)
	) name9243 (
		\wishbone_bd_ram_mem0_reg[125][3]/P0001 ,
		_w11966_,
		_w12012_,
		_w19756_
	);
	LUT4 #(
		.INIT('h0001)
	) name9244 (
		_w19753_,
		_w19754_,
		_w19755_,
		_w19756_,
		_w19757_
	);
	LUT3 #(
		.INIT('h80)
	) name9245 (
		\wishbone_bd_ram_mem0_reg[212][3]/P0001 ,
		_w11929_,
		_w11984_,
		_w19758_
	);
	LUT3 #(
		.INIT('h80)
	) name9246 (
		\wishbone_bd_ram_mem0_reg[241][3]/P0001 ,
		_w11952_,
		_w11977_,
		_w19759_
	);
	LUT3 #(
		.INIT('h80)
	) name9247 (
		\wishbone_bd_ram_mem0_reg[85][3]/P0001 ,
		_w11933_,
		_w11972_,
		_w19760_
	);
	LUT3 #(
		.INIT('h80)
	) name9248 (
		\wishbone_bd_ram_mem0_reg[65][3]/P0001 ,
		_w11949_,
		_w11977_,
		_w19761_
	);
	LUT4 #(
		.INIT('h0001)
	) name9249 (
		_w19758_,
		_w19759_,
		_w19760_,
		_w19761_,
		_w19762_
	);
	LUT3 #(
		.INIT('h80)
	) name9250 (
		\wishbone_bd_ram_mem0_reg[186][3]/P0001 ,
		_w11942_,
		_w11944_,
		_w19763_
	);
	LUT3 #(
		.INIT('h80)
	) name9251 (
		\wishbone_bd_ram_mem0_reg[101][3]/P0001 ,
		_w11933_,
		_w11965_,
		_w19764_
	);
	LUT3 #(
		.INIT('h80)
	) name9252 (
		\wishbone_bd_ram_mem0_reg[210][3]/P0001 ,
		_w11963_,
		_w11984_,
		_w19765_
	);
	LUT3 #(
		.INIT('h80)
	) name9253 (
		\wishbone_bd_ram_mem0_reg[140][3]/P0001 ,
		_w11954_,
		_w11955_,
		_w19766_
	);
	LUT4 #(
		.INIT('h0001)
	) name9254 (
		_w19763_,
		_w19764_,
		_w19765_,
		_w19766_,
		_w19767_
	);
	LUT3 #(
		.INIT('h80)
	) name9255 (
		\wishbone_bd_ram_mem0_reg[87][3]/P0001 ,
		_w11972_,
		_w11975_,
		_w19768_
	);
	LUT3 #(
		.INIT('h80)
	) name9256 (
		\wishbone_bd_ram_mem0_reg[135][3]/P0001 ,
		_w11955_,
		_w11975_,
		_w19769_
	);
	LUT3 #(
		.INIT('h80)
	) name9257 (
		\wishbone_bd_ram_mem0_reg[98][3]/P0001 ,
		_w11963_,
		_w11965_,
		_w19770_
	);
	LUT3 #(
		.INIT('h80)
	) name9258 (
		\wishbone_bd_ram_mem0_reg[198][3]/P0001 ,
		_w11945_,
		_w11986_,
		_w19771_
	);
	LUT4 #(
		.INIT('h0001)
	) name9259 (
		_w19768_,
		_w19769_,
		_w19770_,
		_w19771_,
		_w19772_
	);
	LUT4 #(
		.INIT('h8000)
	) name9260 (
		_w19757_,
		_w19762_,
		_w19767_,
		_w19772_,
		_w19773_
	);
	LUT3 #(
		.INIT('h80)
	) name9261 (
		\wishbone_bd_ram_mem0_reg[86][3]/P0001 ,
		_w11972_,
		_w11986_,
		_w19774_
	);
	LUT3 #(
		.INIT('h80)
	) name9262 (
		\wishbone_bd_ram_mem0_reg[236][3]/P0001 ,
		_w11954_,
		_w11982_,
		_w19775_
	);
	LUT3 #(
		.INIT('h80)
	) name9263 (
		\wishbone_bd_ram_mem0_reg[160][3]/P0001 ,
		_w11930_,
		_w11941_,
		_w19776_
	);
	LUT3 #(
		.INIT('h80)
	) name9264 (
		\wishbone_bd_ram_mem0_reg[32][3]/P0001 ,
		_w11941_,
		_w11957_,
		_w19777_
	);
	LUT4 #(
		.INIT('h0001)
	) name9265 (
		_w19774_,
		_w19775_,
		_w19776_,
		_w19777_,
		_w19778_
	);
	LUT3 #(
		.INIT('h80)
	) name9266 (
		\wishbone_bd_ram_mem0_reg[17][3]/P0001 ,
		_w11935_,
		_w11977_,
		_w19779_
	);
	LUT3 #(
		.INIT('h80)
	) name9267 (
		\wishbone_bd_ram_mem0_reg[57][3]/P0001 ,
		_w11968_,
		_w11979_,
		_w19780_
	);
	LUT3 #(
		.INIT('h80)
	) name9268 (
		\wishbone_bd_ram_mem0_reg[40][3]/P0001 ,
		_w11957_,
		_w11990_,
		_w19781_
	);
	LUT3 #(
		.INIT('h80)
	) name9269 (
		\wishbone_bd_ram_mem0_reg[182][3]/P0001 ,
		_w11942_,
		_w11986_,
		_w19782_
	);
	LUT4 #(
		.INIT('h0001)
	) name9270 (
		_w19779_,
		_w19780_,
		_w19781_,
		_w19782_,
		_w19783_
	);
	LUT3 #(
		.INIT('h80)
	) name9271 (
		\wishbone_bd_ram_mem0_reg[9][3]/P0001 ,
		_w11932_,
		_w11968_,
		_w19784_
	);
	LUT3 #(
		.INIT('h80)
	) name9272 (
		\wishbone_bd_ram_mem0_reg[92][3]/P0001 ,
		_w11954_,
		_w11972_,
		_w19785_
	);
	LUT3 #(
		.INIT('h80)
	) name9273 (
		\wishbone_bd_ram_mem0_reg[39][3]/P0001 ,
		_w11957_,
		_w11975_,
		_w19786_
	);
	LUT3 #(
		.INIT('h80)
	) name9274 (
		\wishbone_bd_ram_mem0_reg[28][3]/P0001 ,
		_w11935_,
		_w11954_,
		_w19787_
	);
	LUT4 #(
		.INIT('h0001)
	) name9275 (
		_w19784_,
		_w19785_,
		_w19786_,
		_w19787_,
		_w19788_
	);
	LUT3 #(
		.INIT('h80)
	) name9276 (
		\wishbone_bd_ram_mem0_reg[189][3]/P0001 ,
		_w11942_,
		_w11966_,
		_w19789_
	);
	LUT3 #(
		.INIT('h80)
	) name9277 (
		\wishbone_bd_ram_mem0_reg[248][3]/P0001 ,
		_w11952_,
		_w11990_,
		_w19790_
	);
	LUT3 #(
		.INIT('h80)
	) name9278 (
		\wishbone_bd_ram_mem0_reg[79][3]/P0001 ,
		_w11949_,
		_w11973_,
		_w19791_
	);
	LUT3 #(
		.INIT('h80)
	) name9279 (
		\wishbone_bd_ram_mem0_reg[167][3]/P0001 ,
		_w11930_,
		_w11975_,
		_w19792_
	);
	LUT4 #(
		.INIT('h0001)
	) name9280 (
		_w19789_,
		_w19790_,
		_w19791_,
		_w19792_,
		_w19793_
	);
	LUT4 #(
		.INIT('h8000)
	) name9281 (
		_w19778_,
		_w19783_,
		_w19788_,
		_w19793_,
		_w19794_
	);
	LUT3 #(
		.INIT('h80)
	) name9282 (
		\wishbone_bd_ram_mem0_reg[76][3]/P0001 ,
		_w11949_,
		_w11954_,
		_w19795_
	);
	LUT3 #(
		.INIT('h80)
	) name9283 (
		\wishbone_bd_ram_mem0_reg[196][3]/P0001 ,
		_w11929_,
		_w11945_,
		_w19796_
	);
	LUT3 #(
		.INIT('h80)
	) name9284 (
		\wishbone_bd_ram_mem0_reg[151][3]/P0001 ,
		_w11959_,
		_w11975_,
		_w19797_
	);
	LUT3 #(
		.INIT('h80)
	) name9285 (
		\wishbone_bd_ram_mem0_reg[185][3]/P0001 ,
		_w11942_,
		_w11968_,
		_w19798_
	);
	LUT4 #(
		.INIT('h0001)
	) name9286 (
		_w19795_,
		_w19796_,
		_w19797_,
		_w19798_,
		_w19799_
	);
	LUT3 #(
		.INIT('h80)
	) name9287 (
		\wishbone_bd_ram_mem0_reg[199][3]/P0001 ,
		_w11945_,
		_w11975_,
		_w19800_
	);
	LUT3 #(
		.INIT('h80)
	) name9288 (
		\wishbone_bd_ram_mem0_reg[83][3]/P0001 ,
		_w11938_,
		_w11972_,
		_w19801_
	);
	LUT3 #(
		.INIT('h80)
	) name9289 (
		\wishbone_bd_ram_mem0_reg[5][3]/P0001 ,
		_w11932_,
		_w11933_,
		_w19802_
	);
	LUT3 #(
		.INIT('h80)
	) name9290 (
		\wishbone_bd_ram_mem0_reg[78][3]/P0001 ,
		_w11948_,
		_w11949_,
		_w19803_
	);
	LUT4 #(
		.INIT('h0001)
	) name9291 (
		_w19800_,
		_w19801_,
		_w19802_,
		_w19803_,
		_w19804_
	);
	LUT3 #(
		.INIT('h80)
	) name9292 (
		\wishbone_bd_ram_mem0_reg[221][3]/P0001 ,
		_w11966_,
		_w11984_,
		_w19805_
	);
	LUT3 #(
		.INIT('h80)
	) name9293 (
		\wishbone_bd_ram_mem0_reg[64][3]/P0001 ,
		_w11941_,
		_w11949_,
		_w19806_
	);
	LUT3 #(
		.INIT('h80)
	) name9294 (
		\wishbone_bd_ram_mem0_reg[139][3]/P0001 ,
		_w11936_,
		_w11955_,
		_w19807_
	);
	LUT3 #(
		.INIT('h80)
	) name9295 (
		\wishbone_bd_ram_mem0_reg[243][3]/P0001 ,
		_w11938_,
		_w11952_,
		_w19808_
	);
	LUT4 #(
		.INIT('h0001)
	) name9296 (
		_w19805_,
		_w19806_,
		_w19807_,
		_w19808_,
		_w19809_
	);
	LUT3 #(
		.INIT('h80)
	) name9297 (
		\wishbone_bd_ram_mem0_reg[59][3]/P0001 ,
		_w11936_,
		_w11979_,
		_w19810_
	);
	LUT3 #(
		.INIT('h80)
	) name9298 (
		\wishbone_bd_ram_mem0_reg[249][3]/P0001 ,
		_w11952_,
		_w11968_,
		_w19811_
	);
	LUT3 #(
		.INIT('h80)
	) name9299 (
		\wishbone_bd_ram_mem0_reg[8][3]/P0001 ,
		_w11932_,
		_w11990_,
		_w19812_
	);
	LUT3 #(
		.INIT('h80)
	) name9300 (
		\wishbone_bd_ram_mem0_reg[81][3]/P0001 ,
		_w11972_,
		_w11977_,
		_w19813_
	);
	LUT4 #(
		.INIT('h0001)
	) name9301 (
		_w19810_,
		_w19811_,
		_w19812_,
		_w19813_,
		_w19814_
	);
	LUT4 #(
		.INIT('h8000)
	) name9302 (
		_w19799_,
		_w19804_,
		_w19809_,
		_w19814_,
		_w19815_
	);
	LUT3 #(
		.INIT('h80)
	) name9303 (
		\wishbone_bd_ram_mem0_reg[131][3]/P0001 ,
		_w11938_,
		_w11955_,
		_w19816_
	);
	LUT3 #(
		.INIT('h80)
	) name9304 (
		\wishbone_bd_ram_mem0_reg[155][3]/P0001 ,
		_w11936_,
		_w11959_,
		_w19817_
	);
	LUT3 #(
		.INIT('h80)
	) name9305 (
		\wishbone_bd_ram_mem0_reg[222][3]/P0001 ,
		_w11948_,
		_w11984_,
		_w19818_
	);
	LUT3 #(
		.INIT('h80)
	) name9306 (
		\wishbone_bd_ram_mem0_reg[46][3]/P0001 ,
		_w11948_,
		_w11957_,
		_w19819_
	);
	LUT4 #(
		.INIT('h0001)
	) name9307 (
		_w19816_,
		_w19817_,
		_w19818_,
		_w19819_,
		_w19820_
	);
	LUT3 #(
		.INIT('h80)
	) name9308 (
		\wishbone_bd_ram_mem0_reg[150][3]/P0001 ,
		_w11959_,
		_w11986_,
		_w19821_
	);
	LUT3 #(
		.INIT('h80)
	) name9309 (
		\wishbone_bd_ram_mem0_reg[207][3]/P0001 ,
		_w11945_,
		_w11973_,
		_w19822_
	);
	LUT3 #(
		.INIT('h80)
	) name9310 (
		\wishbone_bd_ram_mem0_reg[7][3]/P0001 ,
		_w11932_,
		_w11975_,
		_w19823_
	);
	LUT3 #(
		.INIT('h80)
	) name9311 (
		\wishbone_bd_ram_mem0_reg[142][3]/P0001 ,
		_w11948_,
		_w11955_,
		_w19824_
	);
	LUT4 #(
		.INIT('h0001)
	) name9312 (
		_w19821_,
		_w19822_,
		_w19823_,
		_w19824_,
		_w19825_
	);
	LUT3 #(
		.INIT('h80)
	) name9313 (
		\wishbone_bd_ram_mem0_reg[235][3]/P0001 ,
		_w11936_,
		_w11982_,
		_w19826_
	);
	LUT3 #(
		.INIT('h80)
	) name9314 (
		\wishbone_bd_ram_mem0_reg[99][3]/P0001 ,
		_w11938_,
		_w11965_,
		_w19827_
	);
	LUT3 #(
		.INIT('h80)
	) name9315 (
		\wishbone_bd_ram_mem0_reg[147][3]/P0001 ,
		_w11938_,
		_w11959_,
		_w19828_
	);
	LUT3 #(
		.INIT('h80)
	) name9316 (
		\wishbone_bd_ram_mem0_reg[206][3]/P0001 ,
		_w11945_,
		_w11948_,
		_w19829_
	);
	LUT4 #(
		.INIT('h0001)
	) name9317 (
		_w19826_,
		_w19827_,
		_w19828_,
		_w19829_,
		_w19830_
	);
	LUT3 #(
		.INIT('h80)
	) name9318 (
		\wishbone_bd_ram_mem0_reg[242][3]/P0001 ,
		_w11952_,
		_w11963_,
		_w19831_
	);
	LUT3 #(
		.INIT('h80)
	) name9319 (
		\wishbone_bd_ram_mem0_reg[238][3]/P0001 ,
		_w11948_,
		_w11982_,
		_w19832_
	);
	LUT3 #(
		.INIT('h80)
	) name9320 (
		\wishbone_bd_ram_mem0_reg[130][3]/P0001 ,
		_w11955_,
		_w11963_,
		_w19833_
	);
	LUT3 #(
		.INIT('h80)
	) name9321 (
		\wishbone_bd_ram_mem0_reg[141][3]/P0001 ,
		_w11955_,
		_w11966_,
		_w19834_
	);
	LUT4 #(
		.INIT('h0001)
	) name9322 (
		_w19831_,
		_w19832_,
		_w19833_,
		_w19834_,
		_w19835_
	);
	LUT4 #(
		.INIT('h8000)
	) name9323 (
		_w19820_,
		_w19825_,
		_w19830_,
		_w19835_,
		_w19836_
	);
	LUT4 #(
		.INIT('h8000)
	) name9324 (
		_w19773_,
		_w19794_,
		_w19815_,
		_w19836_,
		_w19837_
	);
	LUT3 #(
		.INIT('h80)
	) name9325 (
		\wishbone_bd_ram_mem0_reg[2][3]/P0001 ,
		_w11932_,
		_w11963_,
		_w19838_
	);
	LUT3 #(
		.INIT('h80)
	) name9326 (
		\wishbone_bd_ram_mem0_reg[69][3]/P0001 ,
		_w11933_,
		_w11949_,
		_w19839_
	);
	LUT3 #(
		.INIT('h80)
	) name9327 (
		\wishbone_bd_ram_mem0_reg[152][3]/P0001 ,
		_w11959_,
		_w11990_,
		_w19840_
	);
	LUT3 #(
		.INIT('h80)
	) name9328 (
		\wishbone_bd_ram_mem0_reg[253][3]/P0001 ,
		_w11952_,
		_w11966_,
		_w19841_
	);
	LUT4 #(
		.INIT('h0001)
	) name9329 (
		_w19838_,
		_w19839_,
		_w19840_,
		_w19841_,
		_w19842_
	);
	LUT3 #(
		.INIT('h80)
	) name9330 (
		\wishbone_bd_ram_mem0_reg[29][3]/P0001 ,
		_w11935_,
		_w11966_,
		_w19843_
	);
	LUT3 #(
		.INIT('h80)
	) name9331 (
		\wishbone_bd_ram_mem0_reg[72][3]/P0001 ,
		_w11949_,
		_w11990_,
		_w19844_
	);
	LUT3 #(
		.INIT('h80)
	) name9332 (
		\wishbone_bd_ram_mem0_reg[250][3]/P0001 ,
		_w11944_,
		_w11952_,
		_w19845_
	);
	LUT3 #(
		.INIT('h80)
	) name9333 (
		\wishbone_bd_ram_mem0_reg[71][3]/P0001 ,
		_w11949_,
		_w11975_,
		_w19846_
	);
	LUT4 #(
		.INIT('h0001)
	) name9334 (
		_w19843_,
		_w19844_,
		_w19845_,
		_w19846_,
		_w19847_
	);
	LUT3 #(
		.INIT('h80)
	) name9335 (
		\wishbone_bd_ram_mem0_reg[84][3]/P0001 ,
		_w11929_,
		_w11972_,
		_w19848_
	);
	LUT3 #(
		.INIT('h80)
	) name9336 (
		\wishbone_bd_ram_mem0_reg[50][3]/P0001 ,
		_w11963_,
		_w11979_,
		_w19849_
	);
	LUT3 #(
		.INIT('h80)
	) name9337 (
		\wishbone_bd_ram_mem0_reg[68][3]/P0001 ,
		_w11929_,
		_w11949_,
		_w19850_
	);
	LUT3 #(
		.INIT('h80)
	) name9338 (
		\wishbone_bd_ram_mem0_reg[219][3]/P0001 ,
		_w11936_,
		_w11984_,
		_w19851_
	);
	LUT4 #(
		.INIT('h0001)
	) name9339 (
		_w19848_,
		_w19849_,
		_w19850_,
		_w19851_,
		_w19852_
	);
	LUT3 #(
		.INIT('h80)
	) name9340 (
		\wishbone_bd_ram_mem0_reg[161][3]/P0001 ,
		_w11930_,
		_w11977_,
		_w19853_
	);
	LUT3 #(
		.INIT('h80)
	) name9341 (
		\wishbone_bd_ram_mem0_reg[95][3]/P0001 ,
		_w11972_,
		_w11973_,
		_w19854_
	);
	LUT3 #(
		.INIT('h80)
	) name9342 (
		\wishbone_bd_ram_mem0_reg[132][3]/P0001 ,
		_w11929_,
		_w11955_,
		_w19855_
	);
	LUT3 #(
		.INIT('h80)
	) name9343 (
		\wishbone_bd_ram_mem0_reg[41][3]/P0001 ,
		_w11957_,
		_w11968_,
		_w19856_
	);
	LUT4 #(
		.INIT('h0001)
	) name9344 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w19857_
	);
	LUT4 #(
		.INIT('h8000)
	) name9345 (
		_w19842_,
		_w19847_,
		_w19852_,
		_w19857_,
		_w19858_
	);
	LUT3 #(
		.INIT('h80)
	) name9346 (
		\wishbone_bd_ram_mem0_reg[227][3]/P0001 ,
		_w11938_,
		_w11982_,
		_w19859_
	);
	LUT3 #(
		.INIT('h80)
	) name9347 (
		\wishbone_bd_ram_mem0_reg[33][3]/P0001 ,
		_w11957_,
		_w11977_,
		_w19860_
	);
	LUT3 #(
		.INIT('h80)
	) name9348 (
		\wishbone_bd_ram_mem0_reg[13][3]/P0001 ,
		_w11932_,
		_w11966_,
		_w19861_
	);
	LUT3 #(
		.INIT('h80)
	) name9349 (
		\wishbone_bd_ram_mem0_reg[177][3]/P0001 ,
		_w11942_,
		_w11977_,
		_w19862_
	);
	LUT4 #(
		.INIT('h0001)
	) name9350 (
		_w19859_,
		_w19860_,
		_w19861_,
		_w19862_,
		_w19863_
	);
	LUT3 #(
		.INIT('h80)
	) name9351 (
		\wishbone_bd_ram_mem0_reg[201][3]/P0001 ,
		_w11945_,
		_w11968_,
		_w19864_
	);
	LUT3 #(
		.INIT('h80)
	) name9352 (
		\wishbone_bd_ram_mem0_reg[195][3]/P0001 ,
		_w11938_,
		_w11945_,
		_w19865_
	);
	LUT3 #(
		.INIT('h80)
	) name9353 (
		\wishbone_bd_ram_mem0_reg[188][3]/P0001 ,
		_w11942_,
		_w11954_,
		_w19866_
	);
	LUT3 #(
		.INIT('h80)
	) name9354 (
		\wishbone_bd_ram_mem0_reg[165][3]/P0001 ,
		_w11930_,
		_w11933_,
		_w19867_
	);
	LUT4 #(
		.INIT('h0001)
	) name9355 (
		_w19864_,
		_w19865_,
		_w19866_,
		_w19867_,
		_w19868_
	);
	LUT3 #(
		.INIT('h80)
	) name9356 (
		\wishbone_bd_ram_mem0_reg[60][3]/P0001 ,
		_w11954_,
		_w11979_,
		_w19869_
	);
	LUT3 #(
		.INIT('h80)
	) name9357 (
		\wishbone_bd_ram_mem0_reg[18][3]/P0001 ,
		_w11935_,
		_w11963_,
		_w19870_
	);
	LUT3 #(
		.INIT('h80)
	) name9358 (
		\wishbone_bd_ram_mem0_reg[25][3]/P0001 ,
		_w11935_,
		_w11968_,
		_w19871_
	);
	LUT3 #(
		.INIT('h80)
	) name9359 (
		\wishbone_bd_ram_mem0_reg[124][3]/P0001 ,
		_w11954_,
		_w12012_,
		_w19872_
	);
	LUT4 #(
		.INIT('h0001)
	) name9360 (
		_w19869_,
		_w19870_,
		_w19871_,
		_w19872_,
		_w19873_
	);
	LUT3 #(
		.INIT('h80)
	) name9361 (
		\wishbone_bd_ram_mem0_reg[10][3]/P0001 ,
		_w11932_,
		_w11944_,
		_w19874_
	);
	LUT3 #(
		.INIT('h80)
	) name9362 (
		\wishbone_bd_ram_mem0_reg[23][3]/P0001 ,
		_w11935_,
		_w11975_,
		_w19875_
	);
	LUT3 #(
		.INIT('h80)
	) name9363 (
		\wishbone_bd_ram_mem0_reg[22][3]/P0001 ,
		_w11935_,
		_w11986_,
		_w19876_
	);
	LUT3 #(
		.INIT('h80)
	) name9364 (
		\wishbone_bd_ram_mem0_reg[134][3]/P0001 ,
		_w11955_,
		_w11986_,
		_w19877_
	);
	LUT4 #(
		.INIT('h0001)
	) name9365 (
		_w19874_,
		_w19875_,
		_w19876_,
		_w19877_,
		_w19878_
	);
	LUT4 #(
		.INIT('h8000)
	) name9366 (
		_w19863_,
		_w19868_,
		_w19873_,
		_w19878_,
		_w19879_
	);
	LUT3 #(
		.INIT('h80)
	) name9367 (
		\wishbone_bd_ram_mem0_reg[254][3]/P0001 ,
		_w11948_,
		_w11952_,
		_w19880_
	);
	LUT3 #(
		.INIT('h80)
	) name9368 (
		\wishbone_bd_ram_mem0_reg[6][3]/P0001 ,
		_w11932_,
		_w11986_,
		_w19881_
	);
	LUT3 #(
		.INIT('h80)
	) name9369 (
		\wishbone_bd_ram_mem0_reg[88][3]/P0001 ,
		_w11972_,
		_w11990_,
		_w19882_
	);
	LUT3 #(
		.INIT('h80)
	) name9370 (
		\wishbone_bd_ram_mem0_reg[203][3]/P0001 ,
		_w11936_,
		_w11945_,
		_w19883_
	);
	LUT4 #(
		.INIT('h0001)
	) name9371 (
		_w19880_,
		_w19881_,
		_w19882_,
		_w19883_,
		_w19884_
	);
	LUT3 #(
		.INIT('h80)
	) name9372 (
		\wishbone_bd_ram_mem0_reg[163][3]/P0001 ,
		_w11930_,
		_w11938_,
		_w19885_
	);
	LUT3 #(
		.INIT('h80)
	) name9373 (
		\wishbone_bd_ram_mem0_reg[103][3]/P0001 ,
		_w11965_,
		_w11975_,
		_w19886_
	);
	LUT3 #(
		.INIT('h80)
	) name9374 (
		\wishbone_bd_ram_mem0_reg[100][3]/P0001 ,
		_w11929_,
		_w11965_,
		_w19887_
	);
	LUT3 #(
		.INIT('h80)
	) name9375 (
		\wishbone_bd_ram_mem0_reg[159][3]/P0001 ,
		_w11959_,
		_w11973_,
		_w19888_
	);
	LUT4 #(
		.INIT('h0001)
	) name9376 (
		_w19885_,
		_w19886_,
		_w19887_,
		_w19888_,
		_w19889_
	);
	LUT3 #(
		.INIT('h80)
	) name9377 (
		\wishbone_bd_ram_mem0_reg[104][3]/P0001 ,
		_w11965_,
		_w11990_,
		_w19890_
	);
	LUT3 #(
		.INIT('h80)
	) name9378 (
		\wishbone_bd_ram_mem0_reg[176][3]/P0001 ,
		_w11941_,
		_w11942_,
		_w19891_
	);
	LUT3 #(
		.INIT('h80)
	) name9379 (
		\wishbone_bd_ram_mem0_reg[80][3]/P0001 ,
		_w11941_,
		_w11972_,
		_w19892_
	);
	LUT3 #(
		.INIT('h80)
	) name9380 (
		\wishbone_bd_ram_mem0_reg[200][3]/P0001 ,
		_w11945_,
		_w11990_,
		_w19893_
	);
	LUT4 #(
		.INIT('h0001)
	) name9381 (
		_w19890_,
		_w19891_,
		_w19892_,
		_w19893_,
		_w19894_
	);
	LUT3 #(
		.INIT('h80)
	) name9382 (
		\wishbone_bd_ram_mem0_reg[26][3]/P0001 ,
		_w11935_,
		_w11944_,
		_w19895_
	);
	LUT3 #(
		.INIT('h80)
	) name9383 (
		\wishbone_bd_ram_mem0_reg[218][3]/P0001 ,
		_w11944_,
		_w11984_,
		_w19896_
	);
	LUT3 #(
		.INIT('h80)
	) name9384 (
		\wishbone_bd_ram_mem0_reg[82][3]/P0001 ,
		_w11963_,
		_w11972_,
		_w19897_
	);
	LUT3 #(
		.INIT('h80)
	) name9385 (
		\wishbone_bd_ram_mem0_reg[19][3]/P0001 ,
		_w11935_,
		_w11938_,
		_w19898_
	);
	LUT4 #(
		.INIT('h0001)
	) name9386 (
		_w19895_,
		_w19896_,
		_w19897_,
		_w19898_,
		_w19899_
	);
	LUT4 #(
		.INIT('h8000)
	) name9387 (
		_w19884_,
		_w19889_,
		_w19894_,
		_w19899_,
		_w19900_
	);
	LUT3 #(
		.INIT('h80)
	) name9388 (
		\wishbone_bd_ram_mem0_reg[205][3]/P0001 ,
		_w11945_,
		_w11966_,
		_w19901_
	);
	LUT3 #(
		.INIT('h80)
	) name9389 (
		\wishbone_bd_ram_mem0_reg[255][3]/P0001 ,
		_w11952_,
		_w11973_,
		_w19902_
	);
	LUT3 #(
		.INIT('h80)
	) name9390 (
		\wishbone_bd_ram_mem0_reg[45][3]/P0001 ,
		_w11957_,
		_w11966_,
		_w19903_
	);
	LUT3 #(
		.INIT('h80)
	) name9391 (
		\wishbone_bd_ram_mem0_reg[15][3]/P0001 ,
		_w11932_,
		_w11973_,
		_w19904_
	);
	LUT4 #(
		.INIT('h0001)
	) name9392 (
		_w19901_,
		_w19902_,
		_w19903_,
		_w19904_,
		_w19905_
	);
	LUT3 #(
		.INIT('h80)
	) name9393 (
		\wishbone_bd_ram_mem0_reg[192][3]/P0001 ,
		_w11941_,
		_w11945_,
		_w19906_
	);
	LUT3 #(
		.INIT('h80)
	) name9394 (
		\wishbone_bd_ram_mem0_reg[126][3]/P0001 ,
		_w11948_,
		_w12012_,
		_w19907_
	);
	LUT3 #(
		.INIT('h80)
	) name9395 (
		\wishbone_bd_ram_mem0_reg[240][3]/P0001 ,
		_w11941_,
		_w11952_,
		_w19908_
	);
	LUT3 #(
		.INIT('h80)
	) name9396 (
		\wishbone_bd_ram_mem0_reg[113][3]/P0001 ,
		_w11977_,
		_w12012_,
		_w19909_
	);
	LUT4 #(
		.INIT('h0001)
	) name9397 (
		_w19906_,
		_w19907_,
		_w19908_,
		_w19909_,
		_w19910_
	);
	LUT3 #(
		.INIT('h80)
	) name9398 (
		\wishbone_bd_ram_mem0_reg[252][3]/P0001 ,
		_w11952_,
		_w11954_,
		_w19911_
	);
	LUT3 #(
		.INIT('h80)
	) name9399 (
		\wishbone_bd_ram_mem0_reg[34][3]/P0001 ,
		_w11957_,
		_w11963_,
		_w19912_
	);
	LUT3 #(
		.INIT('h80)
	) name9400 (
		\wishbone_bd_ram_mem0_reg[73][3]/P0001 ,
		_w11949_,
		_w11968_,
		_w19913_
	);
	LUT3 #(
		.INIT('h80)
	) name9401 (
		\wishbone_bd_ram_mem0_reg[234][3]/P0001 ,
		_w11944_,
		_w11982_,
		_w19914_
	);
	LUT4 #(
		.INIT('h0001)
	) name9402 (
		_w19911_,
		_w19912_,
		_w19913_,
		_w19914_,
		_w19915_
	);
	LUT3 #(
		.INIT('h80)
	) name9403 (
		\wishbone_bd_ram_mem0_reg[35][3]/P0001 ,
		_w11938_,
		_w11957_,
		_w19916_
	);
	LUT3 #(
		.INIT('h80)
	) name9404 (
		\wishbone_bd_ram_mem0_reg[62][3]/P0001 ,
		_w11948_,
		_w11979_,
		_w19917_
	);
	LUT3 #(
		.INIT('h80)
	) name9405 (
		\wishbone_bd_ram_mem0_reg[67][3]/P0001 ,
		_w11938_,
		_w11949_,
		_w19918_
	);
	LUT3 #(
		.INIT('h80)
	) name9406 (
		\wishbone_bd_ram_mem0_reg[16][3]/P0001 ,
		_w11935_,
		_w11941_,
		_w19919_
	);
	LUT4 #(
		.INIT('h0001)
	) name9407 (
		_w19916_,
		_w19917_,
		_w19918_,
		_w19919_,
		_w19920_
	);
	LUT4 #(
		.INIT('h8000)
	) name9408 (
		_w19905_,
		_w19910_,
		_w19915_,
		_w19920_,
		_w19921_
	);
	LUT4 #(
		.INIT('h8000)
	) name9409 (
		_w19858_,
		_w19879_,
		_w19900_,
		_w19921_,
		_w19922_
	);
	LUT3 #(
		.INIT('h80)
	) name9410 (
		\wishbone_bd_ram_mem0_reg[20][3]/P0001 ,
		_w11929_,
		_w11935_,
		_w19923_
	);
	LUT3 #(
		.INIT('h80)
	) name9411 (
		\wishbone_bd_ram_mem0_reg[112][3]/P0001 ,
		_w11941_,
		_w12012_,
		_w19924_
	);
	LUT3 #(
		.INIT('h80)
	) name9412 (
		\wishbone_bd_ram_mem0_reg[208][3]/P0001 ,
		_w11941_,
		_w11984_,
		_w19925_
	);
	LUT3 #(
		.INIT('h80)
	) name9413 (
		\wishbone_bd_ram_mem0_reg[169][3]/P0001 ,
		_w11930_,
		_w11968_,
		_w19926_
	);
	LUT4 #(
		.INIT('h0001)
	) name9414 (
		_w19923_,
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_
	);
	LUT3 #(
		.INIT('h80)
	) name9415 (
		\wishbone_bd_ram_mem0_reg[121][3]/P0001 ,
		_w11968_,
		_w12012_,
		_w19928_
	);
	LUT3 #(
		.INIT('h80)
	) name9416 (
		\wishbone_bd_ram_mem0_reg[138][3]/P0001 ,
		_w11944_,
		_w11955_,
		_w19929_
	);
	LUT3 #(
		.INIT('h80)
	) name9417 (
		\wishbone_bd_ram_mem0_reg[47][3]/P0001 ,
		_w11957_,
		_w11973_,
		_w19930_
	);
	LUT3 #(
		.INIT('h80)
	) name9418 (
		\wishbone_bd_ram_mem0_reg[251][3]/P0001 ,
		_w11936_,
		_w11952_,
		_w19931_
	);
	LUT4 #(
		.INIT('h0001)
	) name9419 (
		_w19928_,
		_w19929_,
		_w19930_,
		_w19931_,
		_w19932_
	);
	LUT3 #(
		.INIT('h80)
	) name9420 (
		\wishbone_bd_ram_mem0_reg[214][3]/P0001 ,
		_w11984_,
		_w11986_,
		_w19933_
	);
	LUT3 #(
		.INIT('h80)
	) name9421 (
		\wishbone_bd_ram_mem0_reg[213][3]/P0001 ,
		_w11933_,
		_w11984_,
		_w19934_
	);
	LUT3 #(
		.INIT('h80)
	) name9422 (
		\wishbone_bd_ram_mem0_reg[51][3]/P0001 ,
		_w11938_,
		_w11979_,
		_w19935_
	);
	LUT3 #(
		.INIT('h80)
	) name9423 (
		\wishbone_bd_ram_mem0_reg[220][3]/P0001 ,
		_w11954_,
		_w11984_,
		_w19936_
	);
	LUT4 #(
		.INIT('h0001)
	) name9424 (
		_w19933_,
		_w19934_,
		_w19935_,
		_w19936_,
		_w19937_
	);
	LUT3 #(
		.INIT('h80)
	) name9425 (
		\wishbone_bd_ram_mem0_reg[55][3]/P0001 ,
		_w11975_,
		_w11979_,
		_w19938_
	);
	LUT3 #(
		.INIT('h80)
	) name9426 (
		\wishbone_bd_ram_mem0_reg[24][3]/P0001 ,
		_w11935_,
		_w11990_,
		_w19939_
	);
	LUT3 #(
		.INIT('h80)
	) name9427 (
		\wishbone_bd_ram_mem0_reg[168][3]/P0001 ,
		_w11930_,
		_w11990_,
		_w19940_
	);
	LUT3 #(
		.INIT('h80)
	) name9428 (
		\wishbone_bd_ram_mem0_reg[118][3]/P0001 ,
		_w11986_,
		_w12012_,
		_w19941_
	);
	LUT4 #(
		.INIT('h0001)
	) name9429 (
		_w19938_,
		_w19939_,
		_w19940_,
		_w19941_,
		_w19942_
	);
	LUT4 #(
		.INIT('h8000)
	) name9430 (
		_w19927_,
		_w19932_,
		_w19937_,
		_w19942_,
		_w19943_
	);
	LUT3 #(
		.INIT('h80)
	) name9431 (
		\wishbone_bd_ram_mem0_reg[90][3]/P0001 ,
		_w11944_,
		_w11972_,
		_w19944_
	);
	LUT3 #(
		.INIT('h80)
	) name9432 (
		\wishbone_bd_ram_mem0_reg[75][3]/P0001 ,
		_w11936_,
		_w11949_,
		_w19945_
	);
	LUT3 #(
		.INIT('h80)
	) name9433 (
		\wishbone_bd_ram_mem0_reg[61][3]/P0001 ,
		_w11966_,
		_w11979_,
		_w19946_
	);
	LUT3 #(
		.INIT('h80)
	) name9434 (
		\wishbone_bd_ram_mem0_reg[171][3]/P0001 ,
		_w11930_,
		_w11936_,
		_w19947_
	);
	LUT4 #(
		.INIT('h0001)
	) name9435 (
		_w19944_,
		_w19945_,
		_w19946_,
		_w19947_,
		_w19948_
	);
	LUT3 #(
		.INIT('h80)
	) name9436 (
		\wishbone_bd_ram_mem0_reg[89][3]/P0001 ,
		_w11968_,
		_w11972_,
		_w19949_
	);
	LUT3 #(
		.INIT('h80)
	) name9437 (
		\wishbone_bd_ram_mem0_reg[54][3]/P0001 ,
		_w11979_,
		_w11986_,
		_w19950_
	);
	LUT3 #(
		.INIT('h80)
	) name9438 (
		\wishbone_bd_ram_mem0_reg[31][3]/P0001 ,
		_w11935_,
		_w11973_,
		_w19951_
	);
	LUT3 #(
		.INIT('h80)
	) name9439 (
		\wishbone_bd_ram_mem0_reg[172][3]/P0001 ,
		_w11930_,
		_w11954_,
		_w19952_
	);
	LUT4 #(
		.INIT('h0001)
	) name9440 (
		_w19949_,
		_w19950_,
		_w19951_,
		_w19952_,
		_w19953_
	);
	LUT3 #(
		.INIT('h80)
	) name9441 (
		\wishbone_bd_ram_mem0_reg[114][3]/P0001 ,
		_w11963_,
		_w12012_,
		_w19954_
	);
	LUT3 #(
		.INIT('h80)
	) name9442 (
		\wishbone_bd_ram_mem0_reg[237][3]/P0001 ,
		_w11966_,
		_w11982_,
		_w19955_
	);
	LUT3 #(
		.INIT('h80)
	) name9443 (
		\wishbone_bd_ram_mem0_reg[158][3]/P0001 ,
		_w11948_,
		_w11959_,
		_w19956_
	);
	LUT3 #(
		.INIT('h80)
	) name9444 (
		\wishbone_bd_ram_mem0_reg[173][3]/P0001 ,
		_w11930_,
		_w11966_,
		_w19957_
	);
	LUT4 #(
		.INIT('h0001)
	) name9445 (
		_w19954_,
		_w19955_,
		_w19956_,
		_w19957_,
		_w19958_
	);
	LUT3 #(
		.INIT('h80)
	) name9446 (
		\wishbone_bd_ram_mem0_reg[27][3]/P0001 ,
		_w11935_,
		_w11936_,
		_w19959_
	);
	LUT3 #(
		.INIT('h80)
	) name9447 (
		\wishbone_bd_ram_mem0_reg[166][3]/P0001 ,
		_w11930_,
		_w11986_,
		_w19960_
	);
	LUT3 #(
		.INIT('h80)
	) name9448 (
		\wishbone_bd_ram_mem0_reg[53][3]/P0001 ,
		_w11933_,
		_w11979_,
		_w19961_
	);
	LUT3 #(
		.INIT('h80)
	) name9449 (
		\wishbone_bd_ram_mem0_reg[129][3]/P0001 ,
		_w11955_,
		_w11977_,
		_w19962_
	);
	LUT4 #(
		.INIT('h0001)
	) name9450 (
		_w19959_,
		_w19960_,
		_w19961_,
		_w19962_,
		_w19963_
	);
	LUT4 #(
		.INIT('h8000)
	) name9451 (
		_w19948_,
		_w19953_,
		_w19958_,
		_w19963_,
		_w19964_
	);
	LUT3 #(
		.INIT('h80)
	) name9452 (
		\wishbone_bd_ram_mem0_reg[178][3]/P0001 ,
		_w11942_,
		_w11963_,
		_w19965_
	);
	LUT3 #(
		.INIT('h80)
	) name9453 (
		\wishbone_bd_ram_mem0_reg[170][3]/P0001 ,
		_w11930_,
		_w11944_,
		_w19966_
	);
	LUT3 #(
		.INIT('h80)
	) name9454 (
		\wishbone_bd_ram_mem0_reg[191][3]/P0001 ,
		_w11942_,
		_w11973_,
		_w19967_
	);
	LUT3 #(
		.INIT('h80)
	) name9455 (
		\wishbone_bd_ram_mem0_reg[91][3]/P0001 ,
		_w11936_,
		_w11972_,
		_w19968_
	);
	LUT4 #(
		.INIT('h0001)
	) name9456 (
		_w19965_,
		_w19966_,
		_w19967_,
		_w19968_,
		_w19969_
	);
	LUT3 #(
		.INIT('h80)
	) name9457 (
		\wishbone_bd_ram_mem0_reg[145][3]/P0001 ,
		_w11959_,
		_w11977_,
		_w19970_
	);
	LUT3 #(
		.INIT('h80)
	) name9458 (
		\wishbone_bd_ram_mem0_reg[110][3]/P0001 ,
		_w11948_,
		_w11965_,
		_w19971_
	);
	LUT3 #(
		.INIT('h80)
	) name9459 (
		\wishbone_bd_ram_mem0_reg[116][3]/P0001 ,
		_w11929_,
		_w12012_,
		_w19972_
	);
	LUT3 #(
		.INIT('h80)
	) name9460 (
		\wishbone_bd_ram_mem0_reg[204][3]/P0001 ,
		_w11945_,
		_w11954_,
		_w19973_
	);
	LUT4 #(
		.INIT('h0001)
	) name9461 (
		_w19970_,
		_w19971_,
		_w19972_,
		_w19973_,
		_w19974_
	);
	LUT3 #(
		.INIT('h80)
	) name9462 (
		\wishbone_bd_ram_mem0_reg[1][3]/P0001 ,
		_w11932_,
		_w11977_,
		_w19975_
	);
	LUT3 #(
		.INIT('h80)
	) name9463 (
		\wishbone_bd_ram_mem0_reg[66][3]/P0001 ,
		_w11949_,
		_w11963_,
		_w19976_
	);
	LUT3 #(
		.INIT('h80)
	) name9464 (
		\wishbone_bd_ram_mem0_reg[52][3]/P0001 ,
		_w11929_,
		_w11979_,
		_w19977_
	);
	LUT3 #(
		.INIT('h80)
	) name9465 (
		\wishbone_bd_ram_mem0_reg[232][3]/P0001 ,
		_w11982_,
		_w11990_,
		_w19978_
	);
	LUT4 #(
		.INIT('h0001)
	) name9466 (
		_w19975_,
		_w19976_,
		_w19977_,
		_w19978_,
		_w19979_
	);
	LUT3 #(
		.INIT('h80)
	) name9467 (
		\wishbone_bd_ram_mem0_reg[127][3]/P0001 ,
		_w11973_,
		_w12012_,
		_w19980_
	);
	LUT3 #(
		.INIT('h80)
	) name9468 (
		\wishbone_bd_ram_mem0_reg[107][3]/P0001 ,
		_w11936_,
		_w11965_,
		_w19981_
	);
	LUT3 #(
		.INIT('h80)
	) name9469 (
		\wishbone_bd_ram_mem0_reg[233][3]/P0001 ,
		_w11968_,
		_w11982_,
		_w19982_
	);
	LUT3 #(
		.INIT('h80)
	) name9470 (
		\wishbone_bd_ram_mem0_reg[0][3]/P0001 ,
		_w11932_,
		_w11941_,
		_w19983_
	);
	LUT4 #(
		.INIT('h0001)
	) name9471 (
		_w19980_,
		_w19981_,
		_w19982_,
		_w19983_,
		_w19984_
	);
	LUT4 #(
		.INIT('h8000)
	) name9472 (
		_w19969_,
		_w19974_,
		_w19979_,
		_w19984_,
		_w19985_
	);
	LUT3 #(
		.INIT('h80)
	) name9473 (
		\wishbone_bd_ram_mem0_reg[143][3]/P0001 ,
		_w11955_,
		_w11973_,
		_w19986_
	);
	LUT3 #(
		.INIT('h80)
	) name9474 (
		\wishbone_bd_ram_mem0_reg[63][3]/P0001 ,
		_w11973_,
		_w11979_,
		_w19987_
	);
	LUT3 #(
		.INIT('h80)
	) name9475 (
		\wishbone_bd_ram_mem0_reg[77][3]/P0001 ,
		_w11949_,
		_w11966_,
		_w19988_
	);
	LUT3 #(
		.INIT('h80)
	) name9476 (
		\wishbone_bd_ram_mem0_reg[230][3]/P0001 ,
		_w11982_,
		_w11986_,
		_w19989_
	);
	LUT4 #(
		.INIT('h0001)
	) name9477 (
		_w19986_,
		_w19987_,
		_w19988_,
		_w19989_,
		_w19990_
	);
	LUT3 #(
		.INIT('h80)
	) name9478 (
		\wishbone_bd_ram_mem0_reg[70][3]/P0001 ,
		_w11949_,
		_w11986_,
		_w19991_
	);
	LUT3 #(
		.INIT('h80)
	) name9479 (
		\wishbone_bd_ram_mem0_reg[58][3]/P0001 ,
		_w11944_,
		_w11979_,
		_w19992_
	);
	LUT3 #(
		.INIT('h80)
	) name9480 (
		\wishbone_bd_ram_mem0_reg[136][3]/P0001 ,
		_w11955_,
		_w11990_,
		_w19993_
	);
	LUT3 #(
		.INIT('h80)
	) name9481 (
		\wishbone_bd_ram_mem0_reg[224][3]/P0001 ,
		_w11941_,
		_w11982_,
		_w19994_
	);
	LUT4 #(
		.INIT('h0001)
	) name9482 (
		_w19991_,
		_w19992_,
		_w19993_,
		_w19994_,
		_w19995_
	);
	LUT3 #(
		.INIT('h80)
	) name9483 (
		\wishbone_bd_ram_mem0_reg[36][3]/P0001 ,
		_w11929_,
		_w11957_,
		_w19996_
	);
	LUT3 #(
		.INIT('h80)
	) name9484 (
		\wishbone_bd_ram_mem0_reg[245][3]/P0001 ,
		_w11933_,
		_w11952_,
		_w19997_
	);
	LUT3 #(
		.INIT('h80)
	) name9485 (
		\wishbone_bd_ram_mem0_reg[56][3]/P0001 ,
		_w11979_,
		_w11990_,
		_w19998_
	);
	LUT3 #(
		.INIT('h80)
	) name9486 (
		\wishbone_bd_ram_mem0_reg[193][3]/P0001 ,
		_w11945_,
		_w11977_,
		_w19999_
	);
	LUT4 #(
		.INIT('h0001)
	) name9487 (
		_w19996_,
		_w19997_,
		_w19998_,
		_w19999_,
		_w20000_
	);
	LUT3 #(
		.INIT('h80)
	) name9488 (
		\wishbone_bd_ram_mem0_reg[217][3]/P0001 ,
		_w11968_,
		_w11984_,
		_w20001_
	);
	LUT3 #(
		.INIT('h80)
	) name9489 (
		\wishbone_bd_ram_mem0_reg[154][3]/P0001 ,
		_w11944_,
		_w11959_,
		_w20002_
	);
	LUT3 #(
		.INIT('h80)
	) name9490 (
		\wishbone_bd_ram_mem0_reg[42][3]/P0001 ,
		_w11944_,
		_w11957_,
		_w20003_
	);
	LUT3 #(
		.INIT('h80)
	) name9491 (
		\wishbone_bd_ram_mem0_reg[183][3]/P0001 ,
		_w11942_,
		_w11975_,
		_w20004_
	);
	LUT4 #(
		.INIT('h0001)
	) name9492 (
		_w20001_,
		_w20002_,
		_w20003_,
		_w20004_,
		_w20005_
	);
	LUT4 #(
		.INIT('h8000)
	) name9493 (
		_w19990_,
		_w19995_,
		_w20000_,
		_w20005_,
		_w20006_
	);
	LUT4 #(
		.INIT('h8000)
	) name9494 (
		_w19943_,
		_w19964_,
		_w19985_,
		_w20006_,
		_w20007_
	);
	LUT4 #(
		.INIT('h8000)
	) name9495 (
		_w19752_,
		_w19837_,
		_w19922_,
		_w20007_,
		_w20008_
	);
	LUT3 #(
		.INIT('h15)
	) name9496 (
		wb_rst_i_pad,
		_w19645_,
		_w19666_,
		_w20009_
	);
	LUT3 #(
		.INIT('hba)
	) name9497 (
		_w19667_,
		_w20008_,
		_w20009_,
		_w20010_
	);
	LUT3 #(
		.INIT('h80)
	) name9498 (
		\ethreg1_IPGR2_0_DataOut_reg[4]/NET0131 ,
		_w18800_,
		_w18805_,
		_w20011_
	);
	LUT3 #(
		.INIT('h80)
	) name9499 (
		\ethreg1_MIIRX_DATA_DataOut_reg[4]/NET0131 ,
		_w18785_,
		_w18786_,
		_w20012_
	);
	LUT3 #(
		.INIT('h80)
	) name9500 (
		\ethreg1_MODER_0_DataOut_reg[4]/NET0131 ,
		_w18800_,
		_w18801_,
		_w20013_
	);
	LUT4 #(
		.INIT('h0008)
	) name9501 (
		\ethreg1_RXHASH0_0_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w20014_
	);
	LUT3 #(
		.INIT('h80)
	) name9502 (
		_w18757_,
		_w18758_,
		_w20014_,
		_w20015_
	);
	LUT4 #(
		.INIT('h0001)
	) name9503 (
		_w20011_,
		_w20012_,
		_w20013_,
		_w20015_,
		_w20016_
	);
	LUT3 #(
		.INIT('h80)
	) name9504 (
		\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 ,
		_w18753_,
		_w18754_,
		_w20017_
	);
	LUT3 #(
		.INIT('h80)
	) name9505 (
		\ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131 ,
		_w18753_,
		_w19641_,
		_w20018_
	);
	LUT2 #(
		.INIT('h1)
	) name9506 (
		_w20017_,
		_w20018_,
		_w20019_
	);
	LUT2 #(
		.INIT('h8)
	) name9507 (
		_w20016_,
		_w20019_,
		_w20020_
	);
	LUT3 #(
		.INIT('h80)
	) name9508 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[4]/NET0131 ,
		_w18798_,
		_w18805_,
		_w20021_
	);
	LUT3 #(
		.INIT('h80)
	) name9509 (
		\ethreg1_IPGR1_0_DataOut_reg[4]/NET0131 ,
		_w18785_,
		_w18800_,
		_w20022_
	);
	LUT3 #(
		.INIT('h80)
	) name9510 (
		\ethreg1_IPGT_0_DataOut_reg[4]/NET0131 ,
		_w19646_,
		_w19655_,
		_w20023_
	);
	LUT3 #(
		.INIT('h80)
	) name9511 (
		\ethreg1_INT_MASK_0_DataOut_reg[4]/NET0131 ,
		_w18801_,
		_w19655_,
		_w20024_
	);
	LUT4 #(
		.INIT('h0001)
	) name9512 (
		_w20021_,
		_w20022_,
		_w20023_,
		_w20024_,
		_w20025_
	);
	LUT4 #(
		.INIT('h0008)
	) name9513 (
		\ethreg1_RXHASH1_0_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w20026_
	);
	LUT3 #(
		.INIT('h80)
	) name9514 (
		_w18757_,
		_w18762_,
		_w20026_,
		_w20027_
	);
	LUT4 #(
		.INIT('h0002)
	) name9515 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w20028_
	);
	LUT3 #(
		.INIT('h80)
	) name9516 (
		_w18757_,
		_w18758_,
		_w20028_,
		_w20029_
	);
	LUT4 #(
		.INIT('h0002)
	) name9517 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w20030_
	);
	LUT3 #(
		.INIT('h80)
	) name9518 (
		_w18757_,
		_w18762_,
		_w20030_,
		_w20031_
	);
	LUT3 #(
		.INIT('h80)
	) name9519 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[4]/NET0131 ,
		_w18798_,
		_w18801_,
		_w20032_
	);
	LUT4 #(
		.INIT('h0001)
	) name9520 (
		_w20027_,
		_w20029_,
		_w20031_,
		_w20032_,
		_w20033_
	);
	LUT4 #(
		.INIT('h0020)
	) name9521 (
		\ethreg1_TXCTRL_0_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w20034_
	);
	LUT3 #(
		.INIT('h80)
	) name9522 (
		_w18757_,
		_w18758_,
		_w20034_,
		_w20035_
	);
	LUT3 #(
		.INIT('h80)
	) name9523 (
		\ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131 ,
		_w18786_,
		_w18801_,
		_w20036_
	);
	LUT3 #(
		.INIT('h80)
	) name9524 (
		\ethreg1_irq_busy_reg/NET0131 ,
		_w18800_,
		_w19646_,
		_w20037_
	);
	LUT3 #(
		.INIT('h80)
	) name9525 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[4]/NET0131 ,
		_w18785_,
		_w18798_,
		_w20038_
	);
	LUT4 #(
		.INIT('h0001)
	) name9526 (
		_w20035_,
		_w20036_,
		_w20037_,
		_w20038_,
		_w20039_
	);
	LUT4 #(
		.INIT('h8000)
	) name9527 (
		_w18752_,
		_w20025_,
		_w20033_,
		_w20039_,
		_w20040_
	);
	LUT3 #(
		.INIT('h2a)
	) name9528 (
		_w18752_,
		_w20020_,
		_w20040_,
		_w20041_
	);
	LUT3 #(
		.INIT('h80)
	) name9529 (
		\wishbone_bd_ram_mem0_reg[61][4]/P0001 ,
		_w11966_,
		_w11979_,
		_w20042_
	);
	LUT3 #(
		.INIT('h80)
	) name9530 (
		\wishbone_bd_ram_mem0_reg[72][4]/P0001 ,
		_w11949_,
		_w11990_,
		_w20043_
	);
	LUT3 #(
		.INIT('h80)
	) name9531 (
		\wishbone_bd_ram_mem0_reg[9][4]/P0001 ,
		_w11932_,
		_w11968_,
		_w20044_
	);
	LUT3 #(
		.INIT('h80)
	) name9532 (
		\wishbone_bd_ram_mem0_reg[35][4]/P0001 ,
		_w11938_,
		_w11957_,
		_w20045_
	);
	LUT4 #(
		.INIT('h0001)
	) name9533 (
		_w20042_,
		_w20043_,
		_w20044_,
		_w20045_,
		_w20046_
	);
	LUT3 #(
		.INIT('h80)
	) name9534 (
		\wishbone_bd_ram_mem0_reg[54][4]/P0001 ,
		_w11979_,
		_w11986_,
		_w20047_
	);
	LUT3 #(
		.INIT('h80)
	) name9535 (
		\wishbone_bd_ram_mem0_reg[87][4]/P0001 ,
		_w11972_,
		_w11975_,
		_w20048_
	);
	LUT3 #(
		.INIT('h80)
	) name9536 (
		\wishbone_bd_ram_mem0_reg[119][4]/P0001 ,
		_w11975_,
		_w12012_,
		_w20049_
	);
	LUT3 #(
		.INIT('h80)
	) name9537 (
		\wishbone_bd_ram_mem0_reg[37][4]/P0001 ,
		_w11933_,
		_w11957_,
		_w20050_
	);
	LUT4 #(
		.INIT('h0001)
	) name9538 (
		_w20047_,
		_w20048_,
		_w20049_,
		_w20050_,
		_w20051_
	);
	LUT3 #(
		.INIT('h80)
	) name9539 (
		\wishbone_bd_ram_mem0_reg[48][4]/P0001 ,
		_w11941_,
		_w11979_,
		_w20052_
	);
	LUT3 #(
		.INIT('h80)
	) name9540 (
		\wishbone_bd_ram_mem0_reg[95][4]/P0001 ,
		_w11972_,
		_w11973_,
		_w20053_
	);
	LUT3 #(
		.INIT('h80)
	) name9541 (
		\wishbone_bd_ram_mem0_reg[62][4]/P0001 ,
		_w11948_,
		_w11979_,
		_w20054_
	);
	LUT3 #(
		.INIT('h80)
	) name9542 (
		\wishbone_bd_ram_mem0_reg[139][4]/P0001 ,
		_w11936_,
		_w11955_,
		_w20055_
	);
	LUT4 #(
		.INIT('h0001)
	) name9543 (
		_w20052_,
		_w20053_,
		_w20054_,
		_w20055_,
		_w20056_
	);
	LUT3 #(
		.INIT('h80)
	) name9544 (
		\wishbone_bd_ram_mem0_reg[22][4]/P0001 ,
		_w11935_,
		_w11986_,
		_w20057_
	);
	LUT3 #(
		.INIT('h80)
	) name9545 (
		\wishbone_bd_ram_mem0_reg[187][4]/P0001 ,
		_w11936_,
		_w11942_,
		_w20058_
	);
	LUT3 #(
		.INIT('h80)
	) name9546 (
		\wishbone_bd_ram_mem0_reg[25][4]/P0001 ,
		_w11935_,
		_w11968_,
		_w20059_
	);
	LUT3 #(
		.INIT('h80)
	) name9547 (
		\wishbone_bd_ram_mem0_reg[146][4]/P0001 ,
		_w11959_,
		_w11963_,
		_w20060_
	);
	LUT4 #(
		.INIT('h0001)
	) name9548 (
		_w20057_,
		_w20058_,
		_w20059_,
		_w20060_,
		_w20061_
	);
	LUT4 #(
		.INIT('h8000)
	) name9549 (
		_w20046_,
		_w20051_,
		_w20056_,
		_w20061_,
		_w20062_
	);
	LUT3 #(
		.INIT('h80)
	) name9550 (
		\wishbone_bd_ram_mem0_reg[145][4]/P0001 ,
		_w11959_,
		_w11977_,
		_w20063_
	);
	LUT3 #(
		.INIT('h80)
	) name9551 (
		\wishbone_bd_ram_mem0_reg[107][4]/P0001 ,
		_w11936_,
		_w11965_,
		_w20064_
	);
	LUT3 #(
		.INIT('h80)
	) name9552 (
		\wishbone_bd_ram_mem0_reg[106][4]/P0001 ,
		_w11944_,
		_w11965_,
		_w20065_
	);
	LUT3 #(
		.INIT('h80)
	) name9553 (
		\wishbone_bd_ram_mem0_reg[129][4]/P0001 ,
		_w11955_,
		_w11977_,
		_w20066_
	);
	LUT4 #(
		.INIT('h0001)
	) name9554 (
		_w20063_,
		_w20064_,
		_w20065_,
		_w20066_,
		_w20067_
	);
	LUT3 #(
		.INIT('h80)
	) name9555 (
		\wishbone_bd_ram_mem0_reg[226][4]/P0001 ,
		_w11963_,
		_w11982_,
		_w20068_
	);
	LUT3 #(
		.INIT('h80)
	) name9556 (
		\wishbone_bd_ram_mem0_reg[243][4]/P0001 ,
		_w11938_,
		_w11952_,
		_w20069_
	);
	LUT3 #(
		.INIT('h80)
	) name9557 (
		\wishbone_bd_ram_mem0_reg[36][4]/P0001 ,
		_w11929_,
		_w11957_,
		_w20070_
	);
	LUT3 #(
		.INIT('h80)
	) name9558 (
		\wishbone_bd_ram_mem0_reg[17][4]/P0001 ,
		_w11935_,
		_w11977_,
		_w20071_
	);
	LUT4 #(
		.INIT('h0001)
	) name9559 (
		_w20068_,
		_w20069_,
		_w20070_,
		_w20071_,
		_w20072_
	);
	LUT3 #(
		.INIT('h80)
	) name9560 (
		\wishbone_bd_ram_mem0_reg[231][4]/P0001 ,
		_w11975_,
		_w11982_,
		_w20073_
	);
	LUT3 #(
		.INIT('h80)
	) name9561 (
		\wishbone_bd_ram_mem0_reg[253][4]/P0001 ,
		_w11952_,
		_w11966_,
		_w20074_
	);
	LUT3 #(
		.INIT('h80)
	) name9562 (
		\wishbone_bd_ram_mem0_reg[225][4]/P0001 ,
		_w11977_,
		_w11982_,
		_w20075_
	);
	LUT3 #(
		.INIT('h80)
	) name9563 (
		\wishbone_bd_ram_mem0_reg[5][4]/P0001 ,
		_w11932_,
		_w11933_,
		_w20076_
	);
	LUT4 #(
		.INIT('h0001)
	) name9564 (
		_w20073_,
		_w20074_,
		_w20075_,
		_w20076_,
		_w20077_
	);
	LUT3 #(
		.INIT('h80)
	) name9565 (
		\wishbone_bd_ram_mem0_reg[12][4]/P0001 ,
		_w11932_,
		_w11954_,
		_w20078_
	);
	LUT3 #(
		.INIT('h80)
	) name9566 (
		\wishbone_bd_ram_mem0_reg[244][4]/P0001 ,
		_w11929_,
		_w11952_,
		_w20079_
	);
	LUT3 #(
		.INIT('h80)
	) name9567 (
		\wishbone_bd_ram_mem0_reg[143][4]/P0001 ,
		_w11955_,
		_w11973_,
		_w20080_
	);
	LUT3 #(
		.INIT('h80)
	) name9568 (
		\wishbone_bd_ram_mem0_reg[97][4]/P0001 ,
		_w11965_,
		_w11977_,
		_w20081_
	);
	LUT4 #(
		.INIT('h0001)
	) name9569 (
		_w20078_,
		_w20079_,
		_w20080_,
		_w20081_,
		_w20082_
	);
	LUT4 #(
		.INIT('h8000)
	) name9570 (
		_w20067_,
		_w20072_,
		_w20077_,
		_w20082_,
		_w20083_
	);
	LUT3 #(
		.INIT('h80)
	) name9571 (
		\wishbone_bd_ram_mem0_reg[179][4]/P0001 ,
		_w11938_,
		_w11942_,
		_w20084_
	);
	LUT3 #(
		.INIT('h80)
	) name9572 (
		\wishbone_bd_ram_mem0_reg[184][4]/P0001 ,
		_w11942_,
		_w11990_,
		_w20085_
	);
	LUT3 #(
		.INIT('h80)
	) name9573 (
		\wishbone_bd_ram_mem0_reg[237][4]/P0001 ,
		_w11966_,
		_w11982_,
		_w20086_
	);
	LUT3 #(
		.INIT('h80)
	) name9574 (
		\wishbone_bd_ram_mem0_reg[21][4]/P0001 ,
		_w11933_,
		_w11935_,
		_w20087_
	);
	LUT4 #(
		.INIT('h0001)
	) name9575 (
		_w20084_,
		_w20085_,
		_w20086_,
		_w20087_,
		_w20088_
	);
	LUT3 #(
		.INIT('h80)
	) name9576 (
		\wishbone_bd_ram_mem0_reg[236][4]/P0001 ,
		_w11954_,
		_w11982_,
		_w20089_
	);
	LUT3 #(
		.INIT('h80)
	) name9577 (
		\wishbone_bd_ram_mem0_reg[157][4]/P0001 ,
		_w11959_,
		_w11966_,
		_w20090_
	);
	LUT3 #(
		.INIT('h80)
	) name9578 (
		\wishbone_bd_ram_mem0_reg[111][4]/P0001 ,
		_w11965_,
		_w11973_,
		_w20091_
	);
	LUT3 #(
		.INIT('h80)
	) name9579 (
		\wishbone_bd_ram_mem0_reg[49][4]/P0001 ,
		_w11977_,
		_w11979_,
		_w20092_
	);
	LUT4 #(
		.INIT('h0001)
	) name9580 (
		_w20089_,
		_w20090_,
		_w20091_,
		_w20092_,
		_w20093_
	);
	LUT3 #(
		.INIT('h80)
	) name9581 (
		\wishbone_bd_ram_mem0_reg[86][4]/P0001 ,
		_w11972_,
		_w11986_,
		_w20094_
	);
	LUT3 #(
		.INIT('h80)
	) name9582 (
		\wishbone_bd_ram_mem0_reg[14][4]/P0001 ,
		_w11932_,
		_w11948_,
		_w20095_
	);
	LUT3 #(
		.INIT('h80)
	) name9583 (
		\wishbone_bd_ram_mem0_reg[116][4]/P0001 ,
		_w11929_,
		_w12012_,
		_w20096_
	);
	LUT3 #(
		.INIT('h80)
	) name9584 (
		\wishbone_bd_ram_mem0_reg[186][4]/P0001 ,
		_w11942_,
		_w11944_,
		_w20097_
	);
	LUT4 #(
		.INIT('h0001)
	) name9585 (
		_w20094_,
		_w20095_,
		_w20096_,
		_w20097_,
		_w20098_
	);
	LUT3 #(
		.INIT('h80)
	) name9586 (
		\wishbone_bd_ram_mem0_reg[165][4]/P0001 ,
		_w11930_,
		_w11933_,
		_w20099_
	);
	LUT3 #(
		.INIT('h80)
	) name9587 (
		\wishbone_bd_ram_mem0_reg[147][4]/P0001 ,
		_w11938_,
		_w11959_,
		_w20100_
	);
	LUT3 #(
		.INIT('h80)
	) name9588 (
		\wishbone_bd_ram_mem0_reg[38][4]/P0001 ,
		_w11957_,
		_w11986_,
		_w20101_
	);
	LUT3 #(
		.INIT('h80)
	) name9589 (
		\wishbone_bd_ram_mem0_reg[233][4]/P0001 ,
		_w11968_,
		_w11982_,
		_w20102_
	);
	LUT4 #(
		.INIT('h0001)
	) name9590 (
		_w20099_,
		_w20100_,
		_w20101_,
		_w20102_,
		_w20103_
	);
	LUT4 #(
		.INIT('h8000)
	) name9591 (
		_w20088_,
		_w20093_,
		_w20098_,
		_w20103_,
		_w20104_
	);
	LUT3 #(
		.INIT('h80)
	) name9592 (
		\wishbone_bd_ram_mem0_reg[55][4]/P0001 ,
		_w11975_,
		_w11979_,
		_w20105_
	);
	LUT3 #(
		.INIT('h80)
	) name9593 (
		\wishbone_bd_ram_mem0_reg[77][4]/P0001 ,
		_w11949_,
		_w11966_,
		_w20106_
	);
	LUT3 #(
		.INIT('h80)
	) name9594 (
		\wishbone_bd_ram_mem0_reg[153][4]/P0001 ,
		_w11959_,
		_w11968_,
		_w20107_
	);
	LUT3 #(
		.INIT('h80)
	) name9595 (
		\wishbone_bd_ram_mem0_reg[192][4]/P0001 ,
		_w11941_,
		_w11945_,
		_w20108_
	);
	LUT4 #(
		.INIT('h0001)
	) name9596 (
		_w20105_,
		_w20106_,
		_w20107_,
		_w20108_,
		_w20109_
	);
	LUT3 #(
		.INIT('h80)
	) name9597 (
		\wishbone_bd_ram_mem0_reg[215][4]/P0001 ,
		_w11975_,
		_w11984_,
		_w20110_
	);
	LUT3 #(
		.INIT('h80)
	) name9598 (
		\wishbone_bd_ram_mem0_reg[175][4]/P0001 ,
		_w11930_,
		_w11973_,
		_w20111_
	);
	LUT3 #(
		.INIT('h80)
	) name9599 (
		\wishbone_bd_ram_mem0_reg[60][4]/P0001 ,
		_w11954_,
		_w11979_,
		_w20112_
	);
	LUT3 #(
		.INIT('h80)
	) name9600 (
		\wishbone_bd_ram_mem0_reg[193][4]/P0001 ,
		_w11945_,
		_w11977_,
		_w20113_
	);
	LUT4 #(
		.INIT('h0001)
	) name9601 (
		_w20110_,
		_w20111_,
		_w20112_,
		_w20113_,
		_w20114_
	);
	LUT3 #(
		.INIT('h80)
	) name9602 (
		\wishbone_bd_ram_mem0_reg[196][4]/P0001 ,
		_w11929_,
		_w11945_,
		_w20115_
	);
	LUT3 #(
		.INIT('h80)
	) name9603 (
		\wishbone_bd_ram_mem0_reg[135][4]/P0001 ,
		_w11955_,
		_w11975_,
		_w20116_
	);
	LUT3 #(
		.INIT('h80)
	) name9604 (
		\wishbone_bd_ram_mem0_reg[82][4]/P0001 ,
		_w11963_,
		_w11972_,
		_w20117_
	);
	LUT3 #(
		.INIT('h80)
	) name9605 (
		\wishbone_bd_ram_mem0_reg[166][4]/P0001 ,
		_w11930_,
		_w11986_,
		_w20118_
	);
	LUT4 #(
		.INIT('h0001)
	) name9606 (
		_w20115_,
		_w20116_,
		_w20117_,
		_w20118_,
		_w20119_
	);
	LUT3 #(
		.INIT('h80)
	) name9607 (
		\wishbone_bd_ram_mem0_reg[51][4]/P0001 ,
		_w11938_,
		_w11979_,
		_w20120_
	);
	LUT3 #(
		.INIT('h80)
	) name9608 (
		\wishbone_bd_ram_mem0_reg[206][4]/P0001 ,
		_w11945_,
		_w11948_,
		_w20121_
	);
	LUT3 #(
		.INIT('h80)
	) name9609 (
		\wishbone_bd_ram_mem0_reg[173][4]/P0001 ,
		_w11930_,
		_w11966_,
		_w20122_
	);
	LUT3 #(
		.INIT('h80)
	) name9610 (
		\wishbone_bd_ram_mem0_reg[39][4]/P0001 ,
		_w11957_,
		_w11975_,
		_w20123_
	);
	LUT4 #(
		.INIT('h0001)
	) name9611 (
		_w20120_,
		_w20121_,
		_w20122_,
		_w20123_,
		_w20124_
	);
	LUT4 #(
		.INIT('h8000)
	) name9612 (
		_w20109_,
		_w20114_,
		_w20119_,
		_w20124_,
		_w20125_
	);
	LUT4 #(
		.INIT('h8000)
	) name9613 (
		_w20062_,
		_w20083_,
		_w20104_,
		_w20125_,
		_w20126_
	);
	LUT3 #(
		.INIT('h80)
	) name9614 (
		\wishbone_bd_ram_mem0_reg[141][4]/P0001 ,
		_w11955_,
		_w11966_,
		_w20127_
	);
	LUT3 #(
		.INIT('h80)
	) name9615 (
		\wishbone_bd_ram_mem0_reg[133][4]/P0001 ,
		_w11933_,
		_w11955_,
		_w20128_
	);
	LUT3 #(
		.INIT('h80)
	) name9616 (
		\wishbone_bd_ram_mem0_reg[199][4]/P0001 ,
		_w11945_,
		_w11975_,
		_w20129_
	);
	LUT3 #(
		.INIT('h80)
	) name9617 (
		\wishbone_bd_ram_mem0_reg[120][4]/P0001 ,
		_w11990_,
		_w12012_,
		_w20130_
	);
	LUT4 #(
		.INIT('h0001)
	) name9618 (
		_w20127_,
		_w20128_,
		_w20129_,
		_w20130_,
		_w20131_
	);
	LUT3 #(
		.INIT('h80)
	) name9619 (
		\wishbone_bd_ram_mem0_reg[58][4]/P0001 ,
		_w11944_,
		_w11979_,
		_w20132_
	);
	LUT3 #(
		.INIT('h80)
	) name9620 (
		\wishbone_bd_ram_mem0_reg[101][4]/P0001 ,
		_w11933_,
		_w11965_,
		_w20133_
	);
	LUT3 #(
		.INIT('h80)
	) name9621 (
		\wishbone_bd_ram_mem0_reg[4][4]/P0001 ,
		_w11929_,
		_w11932_,
		_w20134_
	);
	LUT3 #(
		.INIT('h80)
	) name9622 (
		\wishbone_bd_ram_mem0_reg[209][4]/P0001 ,
		_w11977_,
		_w11984_,
		_w20135_
	);
	LUT4 #(
		.INIT('h0001)
	) name9623 (
		_w20132_,
		_w20133_,
		_w20134_,
		_w20135_,
		_w20136_
	);
	LUT3 #(
		.INIT('h80)
	) name9624 (
		\wishbone_bd_ram_mem0_reg[241][4]/P0001 ,
		_w11952_,
		_w11977_,
		_w20137_
	);
	LUT3 #(
		.INIT('h80)
	) name9625 (
		\wishbone_bd_ram_mem0_reg[208][4]/P0001 ,
		_w11941_,
		_w11984_,
		_w20138_
	);
	LUT3 #(
		.INIT('h80)
	) name9626 (
		\wishbone_bd_ram_mem0_reg[93][4]/P0001 ,
		_w11966_,
		_w11972_,
		_w20139_
	);
	LUT3 #(
		.INIT('h80)
	) name9627 (
		\wishbone_bd_ram_mem0_reg[98][4]/P0001 ,
		_w11963_,
		_w11965_,
		_w20140_
	);
	LUT4 #(
		.INIT('h0001)
	) name9628 (
		_w20137_,
		_w20138_,
		_w20139_,
		_w20140_,
		_w20141_
	);
	LUT3 #(
		.INIT('h80)
	) name9629 (
		\wishbone_bd_ram_mem0_reg[228][4]/P0001 ,
		_w11929_,
		_w11982_,
		_w20142_
	);
	LUT3 #(
		.INIT('h80)
	) name9630 (
		\wishbone_bd_ram_mem0_reg[118][4]/P0001 ,
		_w11986_,
		_w12012_,
		_w20143_
	);
	LUT3 #(
		.INIT('h80)
	) name9631 (
		\wishbone_bd_ram_mem0_reg[164][4]/P0001 ,
		_w11929_,
		_w11930_,
		_w20144_
	);
	LUT3 #(
		.INIT('h80)
	) name9632 (
		\wishbone_bd_ram_mem0_reg[202][4]/P0001 ,
		_w11944_,
		_w11945_,
		_w20145_
	);
	LUT4 #(
		.INIT('h0001)
	) name9633 (
		_w20142_,
		_w20143_,
		_w20144_,
		_w20145_,
		_w20146_
	);
	LUT4 #(
		.INIT('h8000)
	) name9634 (
		_w20131_,
		_w20136_,
		_w20141_,
		_w20146_,
		_w20147_
	);
	LUT3 #(
		.INIT('h80)
	) name9635 (
		\wishbone_bd_ram_mem0_reg[156][4]/P0001 ,
		_w11954_,
		_w11959_,
		_w20148_
	);
	LUT3 #(
		.INIT('h80)
	) name9636 (
		\wishbone_bd_ram_mem0_reg[66][4]/P0001 ,
		_w11949_,
		_w11963_,
		_w20149_
	);
	LUT3 #(
		.INIT('h80)
	) name9637 (
		\wishbone_bd_ram_mem0_reg[171][4]/P0001 ,
		_w11930_,
		_w11936_,
		_w20150_
	);
	LUT3 #(
		.INIT('h80)
	) name9638 (
		\wishbone_bd_ram_mem0_reg[182][4]/P0001 ,
		_w11942_,
		_w11986_,
		_w20151_
	);
	LUT4 #(
		.INIT('h0001)
	) name9639 (
		_w20148_,
		_w20149_,
		_w20150_,
		_w20151_,
		_w20152_
	);
	LUT3 #(
		.INIT('h80)
	) name9640 (
		\wishbone_bd_ram_mem0_reg[0][4]/P0001 ,
		_w11932_,
		_w11941_,
		_w20153_
	);
	LUT3 #(
		.INIT('h80)
	) name9641 (
		\wishbone_bd_ram_mem0_reg[161][4]/P0001 ,
		_w11930_,
		_w11977_,
		_w20154_
	);
	LUT3 #(
		.INIT('h80)
	) name9642 (
		\wishbone_bd_ram_mem0_reg[212][4]/P0001 ,
		_w11929_,
		_w11984_,
		_w20155_
	);
	LUT3 #(
		.INIT('h80)
	) name9643 (
		\wishbone_bd_ram_mem0_reg[108][4]/P0001 ,
		_w11954_,
		_w11965_,
		_w20156_
	);
	LUT4 #(
		.INIT('h0001)
	) name9644 (
		_w20153_,
		_w20154_,
		_w20155_,
		_w20156_,
		_w20157_
	);
	LUT3 #(
		.INIT('h80)
	) name9645 (
		\wishbone_bd_ram_mem0_reg[1][4]/P0001 ,
		_w11932_,
		_w11977_,
		_w20158_
	);
	LUT3 #(
		.INIT('h80)
	) name9646 (
		\wishbone_bd_ram_mem0_reg[188][4]/P0001 ,
		_w11942_,
		_w11954_,
		_w20159_
	);
	LUT3 #(
		.INIT('h80)
	) name9647 (
		\wishbone_bd_ram_mem0_reg[246][4]/P0001 ,
		_w11952_,
		_w11986_,
		_w20160_
	);
	LUT3 #(
		.INIT('h80)
	) name9648 (
		\wishbone_bd_ram_mem0_reg[6][4]/P0001 ,
		_w11932_,
		_w11986_,
		_w20161_
	);
	LUT4 #(
		.INIT('h0001)
	) name9649 (
		_w20158_,
		_w20159_,
		_w20160_,
		_w20161_,
		_w20162_
	);
	LUT3 #(
		.INIT('h80)
	) name9650 (
		\wishbone_bd_ram_mem0_reg[3][4]/P0001 ,
		_w11932_,
		_w11938_,
		_w20163_
	);
	LUT3 #(
		.INIT('h80)
	) name9651 (
		\wishbone_bd_ram_mem0_reg[83][4]/P0001 ,
		_w11938_,
		_w11972_,
		_w20164_
	);
	LUT3 #(
		.INIT('h80)
	) name9652 (
		\wishbone_bd_ram_mem0_reg[242][4]/P0001 ,
		_w11952_,
		_w11963_,
		_w20165_
	);
	LUT3 #(
		.INIT('h80)
	) name9653 (
		\wishbone_bd_ram_mem0_reg[234][4]/P0001 ,
		_w11944_,
		_w11982_,
		_w20166_
	);
	LUT4 #(
		.INIT('h0001)
	) name9654 (
		_w20163_,
		_w20164_,
		_w20165_,
		_w20166_,
		_w20167_
	);
	LUT4 #(
		.INIT('h8000)
	) name9655 (
		_w20152_,
		_w20157_,
		_w20162_,
		_w20167_,
		_w20168_
	);
	LUT3 #(
		.INIT('h80)
	) name9656 (
		\wishbone_bd_ram_mem0_reg[240][4]/P0001 ,
		_w11941_,
		_w11952_,
		_w20169_
	);
	LUT3 #(
		.INIT('h80)
	) name9657 (
		\wishbone_bd_ram_mem0_reg[10][4]/P0001 ,
		_w11932_,
		_w11944_,
		_w20170_
	);
	LUT3 #(
		.INIT('h80)
	) name9658 (
		\wishbone_bd_ram_mem0_reg[130][4]/P0001 ,
		_w11955_,
		_w11963_,
		_w20171_
	);
	LUT3 #(
		.INIT('h80)
	) name9659 (
		\wishbone_bd_ram_mem0_reg[43][4]/P0001 ,
		_w11936_,
		_w11957_,
		_w20172_
	);
	LUT4 #(
		.INIT('h0001)
	) name9660 (
		_w20169_,
		_w20170_,
		_w20171_,
		_w20172_,
		_w20173_
	);
	LUT3 #(
		.INIT('h80)
	) name9661 (
		\wishbone_bd_ram_mem0_reg[203][4]/P0001 ,
		_w11936_,
		_w11945_,
		_w20174_
	);
	LUT3 #(
		.INIT('h80)
	) name9662 (
		\wishbone_bd_ram_mem0_reg[252][4]/P0001 ,
		_w11952_,
		_w11954_,
		_w20175_
	);
	LUT3 #(
		.INIT('h80)
	) name9663 (
		\wishbone_bd_ram_mem0_reg[65][4]/P0001 ,
		_w11949_,
		_w11977_,
		_w20176_
	);
	LUT3 #(
		.INIT('h80)
	) name9664 (
		\wishbone_bd_ram_mem0_reg[103][4]/P0001 ,
		_w11965_,
		_w11975_,
		_w20177_
	);
	LUT4 #(
		.INIT('h0001)
	) name9665 (
		_w20174_,
		_w20175_,
		_w20176_,
		_w20177_,
		_w20178_
	);
	LUT3 #(
		.INIT('h80)
	) name9666 (
		\wishbone_bd_ram_mem0_reg[207][4]/P0001 ,
		_w11945_,
		_w11973_,
		_w20179_
	);
	LUT3 #(
		.INIT('h80)
	) name9667 (
		\wishbone_bd_ram_mem0_reg[104][4]/P0001 ,
		_w11965_,
		_w11990_,
		_w20180_
	);
	LUT3 #(
		.INIT('h80)
	) name9668 (
		\wishbone_bd_ram_mem0_reg[63][4]/P0001 ,
		_w11973_,
		_w11979_,
		_w20181_
	);
	LUT3 #(
		.INIT('h80)
	) name9669 (
		\wishbone_bd_ram_mem0_reg[127][4]/P0001 ,
		_w11973_,
		_w12012_,
		_w20182_
	);
	LUT4 #(
		.INIT('h0001)
	) name9670 (
		_w20179_,
		_w20180_,
		_w20181_,
		_w20182_,
		_w20183_
	);
	LUT3 #(
		.INIT('h80)
	) name9671 (
		\wishbone_bd_ram_mem0_reg[177][4]/P0001 ,
		_w11942_,
		_w11977_,
		_w20184_
	);
	LUT3 #(
		.INIT('h80)
	) name9672 (
		\wishbone_bd_ram_mem0_reg[251][4]/P0001 ,
		_w11936_,
		_w11952_,
		_w20185_
	);
	LUT3 #(
		.INIT('h80)
	) name9673 (
		\wishbone_bd_ram_mem0_reg[134][4]/P0001 ,
		_w11955_,
		_w11986_,
		_w20186_
	);
	LUT3 #(
		.INIT('h80)
	) name9674 (
		\wishbone_bd_ram_mem0_reg[110][4]/P0001 ,
		_w11948_,
		_w11965_,
		_w20187_
	);
	LUT4 #(
		.INIT('h0001)
	) name9675 (
		_w20184_,
		_w20185_,
		_w20186_,
		_w20187_,
		_w20188_
	);
	LUT4 #(
		.INIT('h8000)
	) name9676 (
		_w20173_,
		_w20178_,
		_w20183_,
		_w20188_,
		_w20189_
	);
	LUT3 #(
		.INIT('h80)
	) name9677 (
		\wishbone_bd_ram_mem0_reg[88][4]/P0001 ,
		_w11972_,
		_w11990_,
		_w20190_
	);
	LUT3 #(
		.INIT('h80)
	) name9678 (
		\wishbone_bd_ram_mem0_reg[172][4]/P0001 ,
		_w11930_,
		_w11954_,
		_w20191_
	);
	LUT3 #(
		.INIT('h80)
	) name9679 (
		\wishbone_bd_ram_mem0_reg[94][4]/P0001 ,
		_w11948_,
		_w11972_,
		_w20192_
	);
	LUT3 #(
		.INIT('h80)
	) name9680 (
		\wishbone_bd_ram_mem0_reg[213][4]/P0001 ,
		_w11933_,
		_w11984_,
		_w20193_
	);
	LUT4 #(
		.INIT('h0001)
	) name9681 (
		_w20190_,
		_w20191_,
		_w20192_,
		_w20193_,
		_w20194_
	);
	LUT3 #(
		.INIT('h80)
	) name9682 (
		\wishbone_bd_ram_mem0_reg[100][4]/P0001 ,
		_w11929_,
		_w11965_,
		_w20195_
	);
	LUT3 #(
		.INIT('h80)
	) name9683 (
		\wishbone_bd_ram_mem0_reg[168][4]/P0001 ,
		_w11930_,
		_w11990_,
		_w20196_
	);
	LUT3 #(
		.INIT('h80)
	) name9684 (
		\wishbone_bd_ram_mem0_reg[23][4]/P0001 ,
		_w11935_,
		_w11975_,
		_w20197_
	);
	LUT3 #(
		.INIT('h80)
	) name9685 (
		\wishbone_bd_ram_mem0_reg[137][4]/P0001 ,
		_w11955_,
		_w11968_,
		_w20198_
	);
	LUT4 #(
		.INIT('h0001)
	) name9686 (
		_w20195_,
		_w20196_,
		_w20197_,
		_w20198_,
		_w20199_
	);
	LUT3 #(
		.INIT('h80)
	) name9687 (
		\wishbone_bd_ram_mem0_reg[33][4]/P0001 ,
		_w11957_,
		_w11977_,
		_w20200_
	);
	LUT3 #(
		.INIT('h80)
	) name9688 (
		\wishbone_bd_ram_mem0_reg[123][4]/P0001 ,
		_w11936_,
		_w12012_,
		_w20201_
	);
	LUT3 #(
		.INIT('h80)
	) name9689 (
		\wishbone_bd_ram_mem0_reg[28][4]/P0001 ,
		_w11935_,
		_w11954_,
		_w20202_
	);
	LUT3 #(
		.INIT('h80)
	) name9690 (
		\wishbone_bd_ram_mem0_reg[201][4]/P0001 ,
		_w11945_,
		_w11968_,
		_w20203_
	);
	LUT4 #(
		.INIT('h0001)
	) name9691 (
		_w20200_,
		_w20201_,
		_w20202_,
		_w20203_,
		_w20204_
	);
	LUT3 #(
		.INIT('h80)
	) name9692 (
		\wishbone_bd_ram_mem0_reg[140][4]/P0001 ,
		_w11954_,
		_w11955_,
		_w20205_
	);
	LUT3 #(
		.INIT('h80)
	) name9693 (
		\wishbone_bd_ram_mem0_reg[249][4]/P0001 ,
		_w11952_,
		_w11968_,
		_w20206_
	);
	LUT3 #(
		.INIT('h80)
	) name9694 (
		\wishbone_bd_ram_mem0_reg[189][4]/P0001 ,
		_w11942_,
		_w11966_,
		_w20207_
	);
	LUT3 #(
		.INIT('h80)
	) name9695 (
		\wishbone_bd_ram_mem0_reg[34][4]/P0001 ,
		_w11957_,
		_w11963_,
		_w20208_
	);
	LUT4 #(
		.INIT('h0001)
	) name9696 (
		_w20205_,
		_w20206_,
		_w20207_,
		_w20208_,
		_w20209_
	);
	LUT4 #(
		.INIT('h8000)
	) name9697 (
		_w20194_,
		_w20199_,
		_w20204_,
		_w20209_,
		_w20210_
	);
	LUT4 #(
		.INIT('h8000)
	) name9698 (
		_w20147_,
		_w20168_,
		_w20189_,
		_w20210_,
		_w20211_
	);
	LUT3 #(
		.INIT('h80)
	) name9699 (
		\wishbone_bd_ram_mem0_reg[13][4]/P0001 ,
		_w11932_,
		_w11966_,
		_w20212_
	);
	LUT3 #(
		.INIT('h80)
	) name9700 (
		\wishbone_bd_ram_mem0_reg[114][4]/P0001 ,
		_w11963_,
		_w12012_,
		_w20213_
	);
	LUT3 #(
		.INIT('h80)
	) name9701 (
		\wishbone_bd_ram_mem0_reg[142][4]/P0001 ,
		_w11948_,
		_w11955_,
		_w20214_
	);
	LUT3 #(
		.INIT('h80)
	) name9702 (
		\wishbone_bd_ram_mem0_reg[178][4]/P0001 ,
		_w11942_,
		_w11963_,
		_w20215_
	);
	LUT4 #(
		.INIT('h0001)
	) name9703 (
		_w20212_,
		_w20213_,
		_w20214_,
		_w20215_,
		_w20216_
	);
	LUT3 #(
		.INIT('h80)
	) name9704 (
		\wishbone_bd_ram_mem0_reg[64][4]/P0001 ,
		_w11941_,
		_w11949_,
		_w20217_
	);
	LUT3 #(
		.INIT('h80)
	) name9705 (
		\wishbone_bd_ram_mem0_reg[113][4]/P0001 ,
		_w11977_,
		_w12012_,
		_w20218_
	);
	LUT3 #(
		.INIT('h80)
	) name9706 (
		\wishbone_bd_ram_mem0_reg[227][4]/P0001 ,
		_w11938_,
		_w11982_,
		_w20219_
	);
	LUT3 #(
		.INIT('h80)
	) name9707 (
		\wishbone_bd_ram_mem0_reg[105][4]/P0001 ,
		_w11965_,
		_w11968_,
		_w20220_
	);
	LUT4 #(
		.INIT('h0001)
	) name9708 (
		_w20217_,
		_w20218_,
		_w20219_,
		_w20220_,
		_w20221_
	);
	LUT3 #(
		.INIT('h80)
	) name9709 (
		\wishbone_bd_ram_mem0_reg[125][4]/P0001 ,
		_w11966_,
		_w12012_,
		_w20222_
	);
	LUT3 #(
		.INIT('h80)
	) name9710 (
		\wishbone_bd_ram_mem0_reg[30][4]/P0001 ,
		_w11935_,
		_w11948_,
		_w20223_
	);
	LUT3 #(
		.INIT('h80)
	) name9711 (
		\wishbone_bd_ram_mem0_reg[220][4]/P0001 ,
		_w11954_,
		_w11984_,
		_w20224_
	);
	LUT3 #(
		.INIT('h80)
	) name9712 (
		\wishbone_bd_ram_mem0_reg[218][4]/P0001 ,
		_w11944_,
		_w11984_,
		_w20225_
	);
	LUT4 #(
		.INIT('h0001)
	) name9713 (
		_w20222_,
		_w20223_,
		_w20224_,
		_w20225_,
		_w20226_
	);
	LUT3 #(
		.INIT('h80)
	) name9714 (
		\wishbone_bd_ram_mem0_reg[56][4]/P0001 ,
		_w11979_,
		_w11990_,
		_w20227_
	);
	LUT3 #(
		.INIT('h80)
	) name9715 (
		\wishbone_bd_ram_mem0_reg[84][4]/P0001 ,
		_w11929_,
		_w11972_,
		_w20228_
	);
	LUT3 #(
		.INIT('h80)
	) name9716 (
		\wishbone_bd_ram_mem0_reg[232][4]/P0001 ,
		_w11982_,
		_w11990_,
		_w20229_
	);
	LUT3 #(
		.INIT('h80)
	) name9717 (
		\wishbone_bd_ram_mem0_reg[159][4]/P0001 ,
		_w11959_,
		_w11973_,
		_w20230_
	);
	LUT4 #(
		.INIT('h0001)
	) name9718 (
		_w20227_,
		_w20228_,
		_w20229_,
		_w20230_,
		_w20231_
	);
	LUT4 #(
		.INIT('h8000)
	) name9719 (
		_w20216_,
		_w20221_,
		_w20226_,
		_w20231_,
		_w20232_
	);
	LUT3 #(
		.INIT('h80)
	) name9720 (
		\wishbone_bd_ram_mem0_reg[229][4]/P0001 ,
		_w11933_,
		_w11982_,
		_w20233_
	);
	LUT3 #(
		.INIT('h80)
	) name9721 (
		\wishbone_bd_ram_mem0_reg[52][4]/P0001 ,
		_w11929_,
		_w11979_,
		_w20234_
	);
	LUT3 #(
		.INIT('h80)
	) name9722 (
		\wishbone_bd_ram_mem0_reg[126][4]/P0001 ,
		_w11948_,
		_w12012_,
		_w20235_
	);
	LUT3 #(
		.INIT('h80)
	) name9723 (
		\wishbone_bd_ram_mem0_reg[89][4]/P0001 ,
		_w11968_,
		_w11972_,
		_w20236_
	);
	LUT4 #(
		.INIT('h0001)
	) name9724 (
		_w20233_,
		_w20234_,
		_w20235_,
		_w20236_,
		_w20237_
	);
	LUT3 #(
		.INIT('h80)
	) name9725 (
		\wishbone_bd_ram_mem0_reg[254][4]/P0001 ,
		_w11948_,
		_w11952_,
		_w20238_
	);
	LUT3 #(
		.INIT('h80)
	) name9726 (
		\wishbone_bd_ram_mem0_reg[91][4]/P0001 ,
		_w11936_,
		_w11972_,
		_w20239_
	);
	LUT3 #(
		.INIT('h80)
	) name9727 (
		\wishbone_bd_ram_mem0_reg[222][4]/P0001 ,
		_w11948_,
		_w11984_,
		_w20240_
	);
	LUT3 #(
		.INIT('h80)
	) name9728 (
		\wishbone_bd_ram_mem0_reg[154][4]/P0001 ,
		_w11944_,
		_w11959_,
		_w20241_
	);
	LUT4 #(
		.INIT('h0001)
	) name9729 (
		_w20238_,
		_w20239_,
		_w20240_,
		_w20241_,
		_w20242_
	);
	LUT3 #(
		.INIT('h80)
	) name9730 (
		\wishbone_bd_ram_mem0_reg[69][4]/P0001 ,
		_w11933_,
		_w11949_,
		_w20243_
	);
	LUT3 #(
		.INIT('h80)
	) name9731 (
		\wishbone_bd_ram_mem0_reg[42][4]/P0001 ,
		_w11944_,
		_w11957_,
		_w20244_
	);
	LUT3 #(
		.INIT('h80)
	) name9732 (
		\wishbone_bd_ram_mem0_reg[7][4]/P0001 ,
		_w11932_,
		_w11975_,
		_w20245_
	);
	LUT3 #(
		.INIT('h80)
	) name9733 (
		\wishbone_bd_ram_mem0_reg[19][4]/P0001 ,
		_w11935_,
		_w11938_,
		_w20246_
	);
	LUT4 #(
		.INIT('h0001)
	) name9734 (
		_w20243_,
		_w20244_,
		_w20245_,
		_w20246_,
		_w20247_
	);
	LUT3 #(
		.INIT('h80)
	) name9735 (
		\wishbone_bd_ram_mem0_reg[219][4]/P0001 ,
		_w11936_,
		_w11984_,
		_w20248_
	);
	LUT3 #(
		.INIT('h80)
	) name9736 (
		\wishbone_bd_ram_mem0_reg[31][4]/P0001 ,
		_w11935_,
		_w11973_,
		_w20249_
	);
	LUT3 #(
		.INIT('h80)
	) name9737 (
		\wishbone_bd_ram_mem0_reg[248][4]/P0001 ,
		_w11952_,
		_w11990_,
		_w20250_
	);
	LUT3 #(
		.INIT('h80)
	) name9738 (
		\wishbone_bd_ram_mem0_reg[81][4]/P0001 ,
		_w11972_,
		_w11977_,
		_w20251_
	);
	LUT4 #(
		.INIT('h0001)
	) name9739 (
		_w20248_,
		_w20249_,
		_w20250_,
		_w20251_,
		_w20252_
	);
	LUT4 #(
		.INIT('h8000)
	) name9740 (
		_w20237_,
		_w20242_,
		_w20247_,
		_w20252_,
		_w20253_
	);
	LUT3 #(
		.INIT('h80)
	) name9741 (
		\wishbone_bd_ram_mem0_reg[194][4]/P0001 ,
		_w11945_,
		_w11963_,
		_w20254_
	);
	LUT3 #(
		.INIT('h80)
	) name9742 (
		\wishbone_bd_ram_mem0_reg[132][4]/P0001 ,
		_w11929_,
		_w11955_,
		_w20255_
	);
	LUT3 #(
		.INIT('h80)
	) name9743 (
		\wishbone_bd_ram_mem0_reg[2][4]/P0001 ,
		_w11932_,
		_w11963_,
		_w20256_
	);
	LUT3 #(
		.INIT('h80)
	) name9744 (
		\wishbone_bd_ram_mem0_reg[255][4]/P0001 ,
		_w11952_,
		_w11973_,
		_w20257_
	);
	LUT4 #(
		.INIT('h0001)
	) name9745 (
		_w20254_,
		_w20255_,
		_w20256_,
		_w20257_,
		_w20258_
	);
	LUT3 #(
		.INIT('h80)
	) name9746 (
		\wishbone_bd_ram_mem0_reg[221][4]/P0001 ,
		_w11966_,
		_w11984_,
		_w20259_
	);
	LUT3 #(
		.INIT('h80)
	) name9747 (
		\wishbone_bd_ram_mem0_reg[180][4]/P0001 ,
		_w11929_,
		_w11942_,
		_w20260_
	);
	LUT3 #(
		.INIT('h80)
	) name9748 (
		\wishbone_bd_ram_mem0_reg[76][4]/P0001 ,
		_w11949_,
		_w11954_,
		_w20261_
	);
	LUT3 #(
		.INIT('h80)
	) name9749 (
		\wishbone_bd_ram_mem0_reg[74][4]/P0001 ,
		_w11944_,
		_w11949_,
		_w20262_
	);
	LUT4 #(
		.INIT('h0001)
	) name9750 (
		_w20259_,
		_w20260_,
		_w20261_,
		_w20262_,
		_w20263_
	);
	LUT3 #(
		.INIT('h80)
	) name9751 (
		\wishbone_bd_ram_mem0_reg[50][4]/P0001 ,
		_w11963_,
		_w11979_,
		_w20264_
	);
	LUT3 #(
		.INIT('h80)
	) name9752 (
		\wishbone_bd_ram_mem0_reg[92][4]/P0001 ,
		_w11954_,
		_w11972_,
		_w20265_
	);
	LUT3 #(
		.INIT('h80)
	) name9753 (
		\wishbone_bd_ram_mem0_reg[96][4]/P0001 ,
		_w11941_,
		_w11965_,
		_w20266_
	);
	LUT3 #(
		.INIT('h80)
	) name9754 (
		\wishbone_bd_ram_mem0_reg[224][4]/P0001 ,
		_w11941_,
		_w11982_,
		_w20267_
	);
	LUT4 #(
		.INIT('h0001)
	) name9755 (
		_w20264_,
		_w20265_,
		_w20266_,
		_w20267_,
		_w20268_
	);
	LUT3 #(
		.INIT('h80)
	) name9756 (
		\wishbone_bd_ram_mem0_reg[29][4]/P0001 ,
		_w11935_,
		_w11966_,
		_w20269_
	);
	LUT3 #(
		.INIT('h80)
	) name9757 (
		\wishbone_bd_ram_mem0_reg[136][4]/P0001 ,
		_w11955_,
		_w11990_,
		_w20270_
	);
	LUT3 #(
		.INIT('h80)
	) name9758 (
		\wishbone_bd_ram_mem0_reg[162][4]/P0001 ,
		_w11930_,
		_w11963_,
		_w20271_
	);
	LUT3 #(
		.INIT('h80)
	) name9759 (
		\wishbone_bd_ram_mem0_reg[75][4]/P0001 ,
		_w11936_,
		_w11949_,
		_w20272_
	);
	LUT4 #(
		.INIT('h0001)
	) name9760 (
		_w20269_,
		_w20270_,
		_w20271_,
		_w20272_,
		_w20273_
	);
	LUT4 #(
		.INIT('h8000)
	) name9761 (
		_w20258_,
		_w20263_,
		_w20268_,
		_w20273_,
		_w20274_
	);
	LUT3 #(
		.INIT('h80)
	) name9762 (
		\wishbone_bd_ram_mem0_reg[185][4]/P0001 ,
		_w11942_,
		_w11968_,
		_w20275_
	);
	LUT3 #(
		.INIT('h80)
	) name9763 (
		\wishbone_bd_ram_mem0_reg[197][4]/P0001 ,
		_w11933_,
		_w11945_,
		_w20276_
	);
	LUT3 #(
		.INIT('h80)
	) name9764 (
		\wishbone_bd_ram_mem0_reg[169][4]/P0001 ,
		_w11930_,
		_w11968_,
		_w20277_
	);
	LUT3 #(
		.INIT('h80)
	) name9765 (
		\wishbone_bd_ram_mem0_reg[73][4]/P0001 ,
		_w11949_,
		_w11968_,
		_w20278_
	);
	LUT4 #(
		.INIT('h0001)
	) name9766 (
		_w20275_,
		_w20276_,
		_w20277_,
		_w20278_,
		_w20279_
	);
	LUT3 #(
		.INIT('h80)
	) name9767 (
		\wishbone_bd_ram_mem0_reg[57][4]/P0001 ,
		_w11968_,
		_w11979_,
		_w20280_
	);
	LUT3 #(
		.INIT('h80)
	) name9768 (
		\wishbone_bd_ram_mem0_reg[79][4]/P0001 ,
		_w11949_,
		_w11973_,
		_w20281_
	);
	LUT3 #(
		.INIT('h80)
	) name9769 (
		\wishbone_bd_ram_mem0_reg[163][4]/P0001 ,
		_w11930_,
		_w11938_,
		_w20282_
	);
	LUT3 #(
		.INIT('h80)
	) name9770 (
		\wishbone_bd_ram_mem0_reg[211][4]/P0001 ,
		_w11938_,
		_w11984_,
		_w20283_
	);
	LUT4 #(
		.INIT('h0001)
	) name9771 (
		_w20280_,
		_w20281_,
		_w20282_,
		_w20283_,
		_w20284_
	);
	LUT3 #(
		.INIT('h80)
	) name9772 (
		\wishbone_bd_ram_mem0_reg[190][4]/P0001 ,
		_w11942_,
		_w11948_,
		_w20285_
	);
	LUT3 #(
		.INIT('h80)
	) name9773 (
		\wishbone_bd_ram_mem0_reg[18][4]/P0001 ,
		_w11935_,
		_w11963_,
		_w20286_
	);
	LUT3 #(
		.INIT('h80)
	) name9774 (
		\wishbone_bd_ram_mem0_reg[217][4]/P0001 ,
		_w11968_,
		_w11984_,
		_w20287_
	);
	LUT3 #(
		.INIT('h80)
	) name9775 (
		\wishbone_bd_ram_mem0_reg[205][4]/P0001 ,
		_w11945_,
		_w11966_,
		_w20288_
	);
	LUT4 #(
		.INIT('h0001)
	) name9776 (
		_w20285_,
		_w20286_,
		_w20287_,
		_w20288_,
		_w20289_
	);
	LUT3 #(
		.INIT('h80)
	) name9777 (
		\wishbone_bd_ram_mem0_reg[15][4]/P0001 ,
		_w11932_,
		_w11973_,
		_w20290_
	);
	LUT3 #(
		.INIT('h80)
	) name9778 (
		\wishbone_bd_ram_mem0_reg[78][4]/P0001 ,
		_w11948_,
		_w11949_,
		_w20291_
	);
	LUT3 #(
		.INIT('h80)
	) name9779 (
		\wishbone_bd_ram_mem0_reg[204][4]/P0001 ,
		_w11945_,
		_w11954_,
		_w20292_
	);
	LUT3 #(
		.INIT('h80)
	) name9780 (
		\wishbone_bd_ram_mem0_reg[24][4]/P0001 ,
		_w11935_,
		_w11990_,
		_w20293_
	);
	LUT4 #(
		.INIT('h0001)
	) name9781 (
		_w20290_,
		_w20291_,
		_w20292_,
		_w20293_,
		_w20294_
	);
	LUT4 #(
		.INIT('h8000)
	) name9782 (
		_w20279_,
		_w20284_,
		_w20289_,
		_w20294_,
		_w20295_
	);
	LUT4 #(
		.INIT('h8000)
	) name9783 (
		_w20232_,
		_w20253_,
		_w20274_,
		_w20295_,
		_w20296_
	);
	LUT3 #(
		.INIT('h80)
	) name9784 (
		\wishbone_bd_ram_mem0_reg[80][4]/P0001 ,
		_w11941_,
		_w11972_,
		_w20297_
	);
	LUT3 #(
		.INIT('h80)
	) name9785 (
		\wishbone_bd_ram_mem0_reg[53][4]/P0001 ,
		_w11933_,
		_w11979_,
		_w20298_
	);
	LUT3 #(
		.INIT('h80)
	) name9786 (
		\wishbone_bd_ram_mem0_reg[59][4]/P0001 ,
		_w11936_,
		_w11979_,
		_w20299_
	);
	LUT3 #(
		.INIT('h80)
	) name9787 (
		\wishbone_bd_ram_mem0_reg[150][4]/P0001 ,
		_w11959_,
		_w11986_,
		_w20300_
	);
	LUT4 #(
		.INIT('h0001)
	) name9788 (
		_w20297_,
		_w20298_,
		_w20299_,
		_w20300_,
		_w20301_
	);
	LUT3 #(
		.INIT('h80)
	) name9789 (
		\wishbone_bd_ram_mem0_reg[230][4]/P0001 ,
		_w11982_,
		_w11986_,
		_w20302_
	);
	LUT3 #(
		.INIT('h80)
	) name9790 (
		\wishbone_bd_ram_mem0_reg[45][4]/P0001 ,
		_w11957_,
		_w11966_,
		_w20303_
	);
	LUT3 #(
		.INIT('h80)
	) name9791 (
		\wishbone_bd_ram_mem0_reg[160][4]/P0001 ,
		_w11930_,
		_w11941_,
		_w20304_
	);
	LUT3 #(
		.INIT('h80)
	) name9792 (
		\wishbone_bd_ram_mem0_reg[41][4]/P0001 ,
		_w11957_,
		_w11968_,
		_w20305_
	);
	LUT4 #(
		.INIT('h0001)
	) name9793 (
		_w20302_,
		_w20303_,
		_w20304_,
		_w20305_,
		_w20306_
	);
	LUT3 #(
		.INIT('h80)
	) name9794 (
		\wishbone_bd_ram_mem0_reg[117][4]/P0001 ,
		_w11933_,
		_w12012_,
		_w20307_
	);
	LUT3 #(
		.INIT('h80)
	) name9795 (
		\wishbone_bd_ram_mem0_reg[70][4]/P0001 ,
		_w11949_,
		_w11986_,
		_w20308_
	);
	LUT3 #(
		.INIT('h80)
	) name9796 (
		\wishbone_bd_ram_mem0_reg[115][4]/P0001 ,
		_w11938_,
		_w12012_,
		_w20309_
	);
	LUT3 #(
		.INIT('h80)
	) name9797 (
		\wishbone_bd_ram_mem0_reg[183][4]/P0001 ,
		_w11942_,
		_w11975_,
		_w20310_
	);
	LUT4 #(
		.INIT('h0001)
	) name9798 (
		_w20307_,
		_w20308_,
		_w20309_,
		_w20310_,
		_w20311_
	);
	LUT3 #(
		.INIT('h80)
	) name9799 (
		\wishbone_bd_ram_mem0_reg[109][4]/P0001 ,
		_w11965_,
		_w11966_,
		_w20312_
	);
	LUT3 #(
		.INIT('h80)
	) name9800 (
		\wishbone_bd_ram_mem0_reg[170][4]/P0001 ,
		_w11930_,
		_w11944_,
		_w20313_
	);
	LUT3 #(
		.INIT('h80)
	) name9801 (
		\wishbone_bd_ram_mem0_reg[32][4]/P0001 ,
		_w11941_,
		_w11957_,
		_w20314_
	);
	LUT3 #(
		.INIT('h80)
	) name9802 (
		\wishbone_bd_ram_mem0_reg[128][4]/P0001 ,
		_w11941_,
		_w11955_,
		_w20315_
	);
	LUT4 #(
		.INIT('h0001)
	) name9803 (
		_w20312_,
		_w20313_,
		_w20314_,
		_w20315_,
		_w20316_
	);
	LUT4 #(
		.INIT('h8000)
	) name9804 (
		_w20301_,
		_w20306_,
		_w20311_,
		_w20316_,
		_w20317_
	);
	LUT3 #(
		.INIT('h80)
	) name9805 (
		\wishbone_bd_ram_mem0_reg[47][4]/P0001 ,
		_w11957_,
		_w11973_,
		_w20318_
	);
	LUT3 #(
		.INIT('h80)
	) name9806 (
		\wishbone_bd_ram_mem0_reg[181][4]/P0001 ,
		_w11933_,
		_w11942_,
		_w20319_
	);
	LUT3 #(
		.INIT('h80)
	) name9807 (
		\wishbone_bd_ram_mem0_reg[20][4]/P0001 ,
		_w11929_,
		_w11935_,
		_w20320_
	);
	LUT3 #(
		.INIT('h80)
	) name9808 (
		\wishbone_bd_ram_mem0_reg[155][4]/P0001 ,
		_w11936_,
		_w11959_,
		_w20321_
	);
	LUT4 #(
		.INIT('h0001)
	) name9809 (
		_w20318_,
		_w20319_,
		_w20320_,
		_w20321_,
		_w20322_
	);
	LUT3 #(
		.INIT('h80)
	) name9810 (
		\wishbone_bd_ram_mem0_reg[148][4]/P0001 ,
		_w11929_,
		_w11959_,
		_w20323_
	);
	LUT3 #(
		.INIT('h80)
	) name9811 (
		\wishbone_bd_ram_mem0_reg[167][4]/P0001 ,
		_w11930_,
		_w11975_,
		_w20324_
	);
	LUT3 #(
		.INIT('h80)
	) name9812 (
		\wishbone_bd_ram_mem0_reg[216][4]/P0001 ,
		_w11984_,
		_w11990_,
		_w20325_
	);
	LUT3 #(
		.INIT('h80)
	) name9813 (
		\wishbone_bd_ram_mem0_reg[11][4]/P0001 ,
		_w11932_,
		_w11936_,
		_w20326_
	);
	LUT4 #(
		.INIT('h0001)
	) name9814 (
		_w20323_,
		_w20324_,
		_w20325_,
		_w20326_,
		_w20327_
	);
	LUT3 #(
		.INIT('h80)
	) name9815 (
		\wishbone_bd_ram_mem0_reg[68][4]/P0001 ,
		_w11929_,
		_w11949_,
		_w20328_
	);
	LUT3 #(
		.INIT('h80)
	) name9816 (
		\wishbone_bd_ram_mem0_reg[198][4]/P0001 ,
		_w11945_,
		_w11986_,
		_w20329_
	);
	LUT3 #(
		.INIT('h80)
	) name9817 (
		\wishbone_bd_ram_mem0_reg[176][4]/P0001 ,
		_w11941_,
		_w11942_,
		_w20330_
	);
	LUT3 #(
		.INIT('h80)
	) name9818 (
		\wishbone_bd_ram_mem0_reg[26][4]/P0001 ,
		_w11935_,
		_w11944_,
		_w20331_
	);
	LUT4 #(
		.INIT('h0001)
	) name9819 (
		_w20328_,
		_w20329_,
		_w20330_,
		_w20331_,
		_w20332_
	);
	LUT3 #(
		.INIT('h80)
	) name9820 (
		\wishbone_bd_ram_mem0_reg[40][4]/P0001 ,
		_w11957_,
		_w11990_,
		_w20333_
	);
	LUT3 #(
		.INIT('h80)
	) name9821 (
		\wishbone_bd_ram_mem0_reg[149][4]/P0001 ,
		_w11933_,
		_w11959_,
		_w20334_
	);
	LUT3 #(
		.INIT('h80)
	) name9822 (
		\wishbone_bd_ram_mem0_reg[250][4]/P0001 ,
		_w11944_,
		_w11952_,
		_w20335_
	);
	LUT3 #(
		.INIT('h80)
	) name9823 (
		\wishbone_bd_ram_mem0_reg[138][4]/P0001 ,
		_w11944_,
		_w11955_,
		_w20336_
	);
	LUT4 #(
		.INIT('h0001)
	) name9824 (
		_w20333_,
		_w20334_,
		_w20335_,
		_w20336_,
		_w20337_
	);
	LUT4 #(
		.INIT('h8000)
	) name9825 (
		_w20322_,
		_w20327_,
		_w20332_,
		_w20337_,
		_w20338_
	);
	LUT3 #(
		.INIT('h80)
	) name9826 (
		\wishbone_bd_ram_mem0_reg[223][4]/P0001 ,
		_w11973_,
		_w11984_,
		_w20339_
	);
	LUT3 #(
		.INIT('h80)
	) name9827 (
		\wishbone_bd_ram_mem0_reg[27][4]/P0001 ,
		_w11935_,
		_w11936_,
		_w20340_
	);
	LUT3 #(
		.INIT('h80)
	) name9828 (
		\wishbone_bd_ram_mem0_reg[247][4]/P0001 ,
		_w11952_,
		_w11975_,
		_w20341_
	);
	LUT3 #(
		.INIT('h80)
	) name9829 (
		\wishbone_bd_ram_mem0_reg[152][4]/P0001 ,
		_w11959_,
		_w11990_,
		_w20342_
	);
	LUT4 #(
		.INIT('h0001)
	) name9830 (
		_w20339_,
		_w20340_,
		_w20341_,
		_w20342_,
		_w20343_
	);
	LUT3 #(
		.INIT('h80)
	) name9831 (
		\wishbone_bd_ram_mem0_reg[90][4]/P0001 ,
		_w11944_,
		_w11972_,
		_w20344_
	);
	LUT3 #(
		.INIT('h80)
	) name9832 (
		\wishbone_bd_ram_mem0_reg[210][4]/P0001 ,
		_w11963_,
		_w11984_,
		_w20345_
	);
	LUT3 #(
		.INIT('h80)
	) name9833 (
		\wishbone_bd_ram_mem0_reg[71][4]/P0001 ,
		_w11949_,
		_w11975_,
		_w20346_
	);
	LUT3 #(
		.INIT('h80)
	) name9834 (
		\wishbone_bd_ram_mem0_reg[191][4]/P0001 ,
		_w11942_,
		_w11973_,
		_w20347_
	);
	LUT4 #(
		.INIT('h0001)
	) name9835 (
		_w20344_,
		_w20345_,
		_w20346_,
		_w20347_,
		_w20348_
	);
	LUT3 #(
		.INIT('h80)
	) name9836 (
		\wishbone_bd_ram_mem0_reg[121][4]/P0001 ,
		_w11968_,
		_w12012_,
		_w20349_
	);
	LUT3 #(
		.INIT('h80)
	) name9837 (
		\wishbone_bd_ram_mem0_reg[214][4]/P0001 ,
		_w11984_,
		_w11986_,
		_w20350_
	);
	LUT3 #(
		.INIT('h80)
	) name9838 (
		\wishbone_bd_ram_mem0_reg[67][4]/P0001 ,
		_w11938_,
		_w11949_,
		_w20351_
	);
	LUT3 #(
		.INIT('h80)
	) name9839 (
		\wishbone_bd_ram_mem0_reg[124][4]/P0001 ,
		_w11954_,
		_w12012_,
		_w20352_
	);
	LUT4 #(
		.INIT('h0001)
	) name9840 (
		_w20349_,
		_w20350_,
		_w20351_,
		_w20352_,
		_w20353_
	);
	LUT3 #(
		.INIT('h80)
	) name9841 (
		\wishbone_bd_ram_mem0_reg[239][4]/P0001 ,
		_w11973_,
		_w11982_,
		_w20354_
	);
	LUT3 #(
		.INIT('h80)
	) name9842 (
		\wishbone_bd_ram_mem0_reg[174][4]/P0001 ,
		_w11930_,
		_w11948_,
		_w20355_
	);
	LUT3 #(
		.INIT('h80)
	) name9843 (
		\wishbone_bd_ram_mem0_reg[245][4]/P0001 ,
		_w11933_,
		_w11952_,
		_w20356_
	);
	LUT3 #(
		.INIT('h80)
	) name9844 (
		\wishbone_bd_ram_mem0_reg[16][4]/P0001 ,
		_w11935_,
		_w11941_,
		_w20357_
	);
	LUT4 #(
		.INIT('h0001)
	) name9845 (
		_w20354_,
		_w20355_,
		_w20356_,
		_w20357_,
		_w20358_
	);
	LUT4 #(
		.INIT('h8000)
	) name9846 (
		_w20343_,
		_w20348_,
		_w20353_,
		_w20358_,
		_w20359_
	);
	LUT3 #(
		.INIT('h80)
	) name9847 (
		\wishbone_bd_ram_mem0_reg[151][4]/P0001 ,
		_w11959_,
		_w11975_,
		_w20360_
	);
	LUT3 #(
		.INIT('h80)
	) name9848 (
		\wishbone_bd_ram_mem0_reg[131][4]/P0001 ,
		_w11938_,
		_w11955_,
		_w20361_
	);
	LUT3 #(
		.INIT('h80)
	) name9849 (
		\wishbone_bd_ram_mem0_reg[144][4]/P0001 ,
		_w11941_,
		_w11959_,
		_w20362_
	);
	LUT3 #(
		.INIT('h80)
	) name9850 (
		\wishbone_bd_ram_mem0_reg[102][4]/P0001 ,
		_w11965_,
		_w11986_,
		_w20363_
	);
	LUT4 #(
		.INIT('h0001)
	) name9851 (
		_w20360_,
		_w20361_,
		_w20362_,
		_w20363_,
		_w20364_
	);
	LUT3 #(
		.INIT('h80)
	) name9852 (
		\wishbone_bd_ram_mem0_reg[238][4]/P0001 ,
		_w11948_,
		_w11982_,
		_w20365_
	);
	LUT3 #(
		.INIT('h80)
	) name9853 (
		\wishbone_bd_ram_mem0_reg[200][4]/P0001 ,
		_w11945_,
		_w11990_,
		_w20366_
	);
	LUT3 #(
		.INIT('h80)
	) name9854 (
		\wishbone_bd_ram_mem0_reg[122][4]/P0001 ,
		_w11944_,
		_w12012_,
		_w20367_
	);
	LUT3 #(
		.INIT('h80)
	) name9855 (
		\wishbone_bd_ram_mem0_reg[235][4]/P0001 ,
		_w11936_,
		_w11982_,
		_w20368_
	);
	LUT4 #(
		.INIT('h0001)
	) name9856 (
		_w20365_,
		_w20366_,
		_w20367_,
		_w20368_,
		_w20369_
	);
	LUT3 #(
		.INIT('h80)
	) name9857 (
		\wishbone_bd_ram_mem0_reg[46][4]/P0001 ,
		_w11948_,
		_w11957_,
		_w20370_
	);
	LUT3 #(
		.INIT('h80)
	) name9858 (
		\wishbone_bd_ram_mem0_reg[44][4]/P0001 ,
		_w11954_,
		_w11957_,
		_w20371_
	);
	LUT3 #(
		.INIT('h80)
	) name9859 (
		\wishbone_bd_ram_mem0_reg[195][4]/P0001 ,
		_w11938_,
		_w11945_,
		_w20372_
	);
	LUT3 #(
		.INIT('h80)
	) name9860 (
		\wishbone_bd_ram_mem0_reg[112][4]/P0001 ,
		_w11941_,
		_w12012_,
		_w20373_
	);
	LUT4 #(
		.INIT('h0001)
	) name9861 (
		_w20370_,
		_w20371_,
		_w20372_,
		_w20373_,
		_w20374_
	);
	LUT3 #(
		.INIT('h80)
	) name9862 (
		\wishbone_bd_ram_mem0_reg[99][4]/P0001 ,
		_w11938_,
		_w11965_,
		_w20375_
	);
	LUT3 #(
		.INIT('h80)
	) name9863 (
		\wishbone_bd_ram_mem0_reg[158][4]/P0001 ,
		_w11948_,
		_w11959_,
		_w20376_
	);
	LUT3 #(
		.INIT('h80)
	) name9864 (
		\wishbone_bd_ram_mem0_reg[8][4]/P0001 ,
		_w11932_,
		_w11990_,
		_w20377_
	);
	LUT3 #(
		.INIT('h80)
	) name9865 (
		\wishbone_bd_ram_mem0_reg[85][4]/P0001 ,
		_w11933_,
		_w11972_,
		_w20378_
	);
	LUT4 #(
		.INIT('h0001)
	) name9866 (
		_w20375_,
		_w20376_,
		_w20377_,
		_w20378_,
		_w20379_
	);
	LUT4 #(
		.INIT('h8000)
	) name9867 (
		_w20364_,
		_w20369_,
		_w20374_,
		_w20379_,
		_w20380_
	);
	LUT4 #(
		.INIT('h8000)
	) name9868 (
		_w20317_,
		_w20338_,
		_w20359_,
		_w20380_,
		_w20381_
	);
	LUT4 #(
		.INIT('h8000)
	) name9869 (
		_w20126_,
		_w20211_,
		_w20296_,
		_w20381_,
		_w20382_
	);
	LUT3 #(
		.INIT('h15)
	) name9870 (
		wb_rst_i_pad,
		_w20020_,
		_w20040_,
		_w20383_
	);
	LUT3 #(
		.INIT('hba)
	) name9871 (
		_w20041_,
		_w20382_,
		_w20383_,
		_w20384_
	);
	LUT3 #(
		.INIT('h80)
	) name9872 (
		\ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131 ,
		_w18753_,
		_w19641_,
		_w20385_
	);
	LUT3 #(
		.INIT('h80)
	) name9873 (
		\ethreg1_irq_txc_reg/NET0131 ,
		_w18800_,
		_w19646_,
		_w20386_
	);
	LUT3 #(
		.INIT('h80)
	) name9874 (
		\ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131 ,
		_w18786_,
		_w18801_,
		_w20387_
	);
	LUT3 #(
		.INIT('h80)
	) name9875 (
		\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 ,
		_w18753_,
		_w18754_,
		_w20388_
	);
	LUT3 #(
		.INIT('h80)
	) name9876 (
		\ethreg1_MIIRX_DATA_DataOut_reg[5]/NET0131 ,
		_w18785_,
		_w18786_,
		_w20389_
	);
	LUT4 #(
		.INIT('h0001)
	) name9877 (
		_w20386_,
		_w20387_,
		_w20388_,
		_w20389_,
		_w20390_
	);
	LUT2 #(
		.INIT('h4)
	) name9878 (
		_w20385_,
		_w20390_,
		_w20391_
	);
	LUT3 #(
		.INIT('h80)
	) name9879 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[5]/NET0131 ,
		_w18798_,
		_w18805_,
		_w20392_
	);
	LUT4 #(
		.INIT('h0002)
	) name9880 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w20393_
	);
	LUT3 #(
		.INIT('h80)
	) name9881 (
		_w18757_,
		_w18762_,
		_w20393_,
		_w20394_
	);
	LUT4 #(
		.INIT('h0008)
	) name9882 (
		\ethreg1_RXHASH1_0_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w20395_
	);
	LUT3 #(
		.INIT('h80)
	) name9883 (
		_w18757_,
		_w18762_,
		_w20395_,
		_w20396_
	);
	LUT3 #(
		.INIT('h80)
	) name9884 (
		\ethreg1_IPGR1_0_DataOut_reg[5]/NET0131 ,
		_w18785_,
		_w18800_,
		_w20397_
	);
	LUT4 #(
		.INIT('h0001)
	) name9885 (
		_w20392_,
		_w20394_,
		_w20396_,
		_w20397_,
		_w20398_
	);
	LUT4 #(
		.INIT('h0008)
	) name9886 (
		\ethreg1_RXHASH0_0_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w20399_
	);
	LUT3 #(
		.INIT('h80)
	) name9887 (
		_w18757_,
		_w18758_,
		_w20399_,
		_w20400_
	);
	LUT3 #(
		.INIT('h80)
	) name9888 (
		\ethreg1_INT_MASK_0_DataOut_reg[5]/NET0131 ,
		_w18801_,
		_w19655_,
		_w20401_
	);
	LUT3 #(
		.INIT('h80)
	) name9889 (
		\ethreg1_IPGT_0_DataOut_reg[5]/NET0131 ,
		_w19646_,
		_w19655_,
		_w20402_
	);
	LUT3 #(
		.INIT('h80)
	) name9890 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[5]/NET0131 ,
		_w18798_,
		_w18801_,
		_w20403_
	);
	LUT4 #(
		.INIT('h0001)
	) name9891 (
		_w20400_,
		_w20401_,
		_w20402_,
		_w20403_,
		_w20404_
	);
	LUT3 #(
		.INIT('h80)
	) name9892 (
		\ethreg1_MODER_0_DataOut_reg[5]/NET0131 ,
		_w18800_,
		_w18801_,
		_w20405_
	);
	LUT4 #(
		.INIT('h0002)
	) name9893 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w20406_
	);
	LUT3 #(
		.INIT('h80)
	) name9894 (
		_w18757_,
		_w18758_,
		_w20406_,
		_w20407_
	);
	LUT4 #(
		.INIT('h0020)
	) name9895 (
		\ethreg1_TXCTRL_0_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w20408_
	);
	LUT3 #(
		.INIT('h80)
	) name9896 (
		_w18757_,
		_w18758_,
		_w20408_,
		_w20409_
	);
	LUT3 #(
		.INIT('h80)
	) name9897 (
		\ethreg1_IPGR2_0_DataOut_reg[5]/NET0131 ,
		_w18800_,
		_w18805_,
		_w20410_
	);
	LUT4 #(
		.INIT('h0001)
	) name9898 (
		_w20405_,
		_w20407_,
		_w20409_,
		_w20410_,
		_w20411_
	);
	LUT4 #(
		.INIT('h8000)
	) name9899 (
		_w18752_,
		_w20398_,
		_w20404_,
		_w20411_,
		_w20412_
	);
	LUT3 #(
		.INIT('h2a)
	) name9900 (
		_w18752_,
		_w20391_,
		_w20412_,
		_w20413_
	);
	LUT3 #(
		.INIT('h80)
	) name9901 (
		\wishbone_bd_ram_mem0_reg[80][5]/P0001 ,
		_w11941_,
		_w11972_,
		_w20414_
	);
	LUT3 #(
		.INIT('h80)
	) name9902 (
		\wishbone_bd_ram_mem0_reg[37][5]/P0001 ,
		_w11933_,
		_w11957_,
		_w20415_
	);
	LUT3 #(
		.INIT('h80)
	) name9903 (
		\wishbone_bd_ram_mem0_reg[18][5]/P0001 ,
		_w11935_,
		_w11963_,
		_w20416_
	);
	LUT3 #(
		.INIT('h80)
	) name9904 (
		\wishbone_bd_ram_mem0_reg[73][5]/P0001 ,
		_w11949_,
		_w11968_,
		_w20417_
	);
	LUT4 #(
		.INIT('h0001)
	) name9905 (
		_w20414_,
		_w20415_,
		_w20416_,
		_w20417_,
		_w20418_
	);
	LUT3 #(
		.INIT('h80)
	) name9906 (
		\wishbone_bd_ram_mem0_reg[241][5]/P0001 ,
		_w11952_,
		_w11977_,
		_w20419_
	);
	LUT3 #(
		.INIT('h80)
	) name9907 (
		\wishbone_bd_ram_mem0_reg[193][5]/P0001 ,
		_w11945_,
		_w11977_,
		_w20420_
	);
	LUT3 #(
		.INIT('h80)
	) name9908 (
		\wishbone_bd_ram_mem0_reg[141][5]/P0001 ,
		_w11955_,
		_w11966_,
		_w20421_
	);
	LUT3 #(
		.INIT('h80)
	) name9909 (
		\wishbone_bd_ram_mem0_reg[203][5]/P0001 ,
		_w11936_,
		_w11945_,
		_w20422_
	);
	LUT4 #(
		.INIT('h0001)
	) name9910 (
		_w20419_,
		_w20420_,
		_w20421_,
		_w20422_,
		_w20423_
	);
	LUT3 #(
		.INIT('h80)
	) name9911 (
		\wishbone_bd_ram_mem0_reg[187][5]/P0001 ,
		_w11936_,
		_w11942_,
		_w20424_
	);
	LUT3 #(
		.INIT('h80)
	) name9912 (
		\wishbone_bd_ram_mem0_reg[170][5]/P0001 ,
		_w11930_,
		_w11944_,
		_w20425_
	);
	LUT3 #(
		.INIT('h80)
	) name9913 (
		\wishbone_bd_ram_mem0_reg[29][5]/P0001 ,
		_w11935_,
		_w11966_,
		_w20426_
	);
	LUT3 #(
		.INIT('h80)
	) name9914 (
		\wishbone_bd_ram_mem0_reg[210][5]/P0001 ,
		_w11963_,
		_w11984_,
		_w20427_
	);
	LUT4 #(
		.INIT('h0001)
	) name9915 (
		_w20424_,
		_w20425_,
		_w20426_,
		_w20427_,
		_w20428_
	);
	LUT3 #(
		.INIT('h80)
	) name9916 (
		\wishbone_bd_ram_mem0_reg[159][5]/P0001 ,
		_w11959_,
		_w11973_,
		_w20429_
	);
	LUT3 #(
		.INIT('h80)
	) name9917 (
		\wishbone_bd_ram_mem0_reg[248][5]/P0001 ,
		_w11952_,
		_w11990_,
		_w20430_
	);
	LUT3 #(
		.INIT('h80)
	) name9918 (
		\wishbone_bd_ram_mem0_reg[48][5]/P0001 ,
		_w11941_,
		_w11979_,
		_w20431_
	);
	LUT3 #(
		.INIT('h80)
	) name9919 (
		\wishbone_bd_ram_mem0_reg[121][5]/P0001 ,
		_w11968_,
		_w12012_,
		_w20432_
	);
	LUT4 #(
		.INIT('h0001)
	) name9920 (
		_w20429_,
		_w20430_,
		_w20431_,
		_w20432_,
		_w20433_
	);
	LUT4 #(
		.INIT('h8000)
	) name9921 (
		_w20418_,
		_w20423_,
		_w20428_,
		_w20433_,
		_w20434_
	);
	LUT3 #(
		.INIT('h80)
	) name9922 (
		\wishbone_bd_ram_mem0_reg[23][5]/P0001 ,
		_w11935_,
		_w11975_,
		_w20435_
	);
	LUT3 #(
		.INIT('h80)
	) name9923 (
		\wishbone_bd_ram_mem0_reg[145][5]/P0001 ,
		_w11959_,
		_w11977_,
		_w20436_
	);
	LUT3 #(
		.INIT('h80)
	) name9924 (
		\wishbone_bd_ram_mem0_reg[44][5]/P0001 ,
		_w11954_,
		_w11957_,
		_w20437_
	);
	LUT3 #(
		.INIT('h80)
	) name9925 (
		\wishbone_bd_ram_mem0_reg[136][5]/P0001 ,
		_w11955_,
		_w11990_,
		_w20438_
	);
	LUT4 #(
		.INIT('h0001)
	) name9926 (
		_w20435_,
		_w20436_,
		_w20437_,
		_w20438_,
		_w20439_
	);
	LUT3 #(
		.INIT('h80)
	) name9927 (
		\wishbone_bd_ram_mem0_reg[201][5]/P0001 ,
		_w11945_,
		_w11968_,
		_w20440_
	);
	LUT3 #(
		.INIT('h80)
	) name9928 (
		\wishbone_bd_ram_mem0_reg[183][5]/P0001 ,
		_w11942_,
		_w11975_,
		_w20441_
	);
	LUT3 #(
		.INIT('h80)
	) name9929 (
		\wishbone_bd_ram_mem0_reg[76][5]/P0001 ,
		_w11949_,
		_w11954_,
		_w20442_
	);
	LUT3 #(
		.INIT('h80)
	) name9930 (
		\wishbone_bd_ram_mem0_reg[43][5]/P0001 ,
		_w11936_,
		_w11957_,
		_w20443_
	);
	LUT4 #(
		.INIT('h0001)
	) name9931 (
		_w20440_,
		_w20441_,
		_w20442_,
		_w20443_,
		_w20444_
	);
	LUT3 #(
		.INIT('h80)
	) name9932 (
		\wishbone_bd_ram_mem0_reg[236][5]/P0001 ,
		_w11954_,
		_w11982_,
		_w20445_
	);
	LUT3 #(
		.INIT('h80)
	) name9933 (
		\wishbone_bd_ram_mem0_reg[207][5]/P0001 ,
		_w11945_,
		_w11973_,
		_w20446_
	);
	LUT3 #(
		.INIT('h80)
	) name9934 (
		\wishbone_bd_ram_mem0_reg[227][5]/P0001 ,
		_w11938_,
		_w11982_,
		_w20447_
	);
	LUT3 #(
		.INIT('h80)
	) name9935 (
		\wishbone_bd_ram_mem0_reg[138][5]/P0001 ,
		_w11944_,
		_w11955_,
		_w20448_
	);
	LUT4 #(
		.INIT('h0001)
	) name9936 (
		_w20445_,
		_w20446_,
		_w20447_,
		_w20448_,
		_w20449_
	);
	LUT3 #(
		.INIT('h80)
	) name9937 (
		\wishbone_bd_ram_mem0_reg[13][5]/P0001 ,
		_w11932_,
		_w11966_,
		_w20450_
	);
	LUT3 #(
		.INIT('h80)
	) name9938 (
		\wishbone_bd_ram_mem0_reg[74][5]/P0001 ,
		_w11944_,
		_w11949_,
		_w20451_
	);
	LUT3 #(
		.INIT('h80)
	) name9939 (
		\wishbone_bd_ram_mem0_reg[125][5]/P0001 ,
		_w11966_,
		_w12012_,
		_w20452_
	);
	LUT3 #(
		.INIT('h80)
	) name9940 (
		\wishbone_bd_ram_mem0_reg[216][5]/P0001 ,
		_w11984_,
		_w11990_,
		_w20453_
	);
	LUT4 #(
		.INIT('h0001)
	) name9941 (
		_w20450_,
		_w20451_,
		_w20452_,
		_w20453_,
		_w20454_
	);
	LUT4 #(
		.INIT('h8000)
	) name9942 (
		_w20439_,
		_w20444_,
		_w20449_,
		_w20454_,
		_w20455_
	);
	LUT3 #(
		.INIT('h80)
	) name9943 (
		\wishbone_bd_ram_mem0_reg[243][5]/P0001 ,
		_w11938_,
		_w11952_,
		_w20456_
	);
	LUT3 #(
		.INIT('h80)
	) name9944 (
		\wishbone_bd_ram_mem0_reg[99][5]/P0001 ,
		_w11938_,
		_w11965_,
		_w20457_
	);
	LUT3 #(
		.INIT('h80)
	) name9945 (
		\wishbone_bd_ram_mem0_reg[93][5]/P0001 ,
		_w11966_,
		_w11972_,
		_w20458_
	);
	LUT3 #(
		.INIT('h80)
	) name9946 (
		\wishbone_bd_ram_mem0_reg[65][5]/P0001 ,
		_w11949_,
		_w11977_,
		_w20459_
	);
	LUT4 #(
		.INIT('h0001)
	) name9947 (
		_w20456_,
		_w20457_,
		_w20458_,
		_w20459_,
		_w20460_
	);
	LUT3 #(
		.INIT('h80)
	) name9948 (
		\wishbone_bd_ram_mem0_reg[220][5]/P0001 ,
		_w11954_,
		_w11984_,
		_w20461_
	);
	LUT3 #(
		.INIT('h80)
	) name9949 (
		\wishbone_bd_ram_mem0_reg[245][5]/P0001 ,
		_w11933_,
		_w11952_,
		_w20462_
	);
	LUT3 #(
		.INIT('h80)
	) name9950 (
		\wishbone_bd_ram_mem0_reg[214][5]/P0001 ,
		_w11984_,
		_w11986_,
		_w20463_
	);
	LUT3 #(
		.INIT('h80)
	) name9951 (
		\wishbone_bd_ram_mem0_reg[108][5]/P0001 ,
		_w11954_,
		_w11965_,
		_w20464_
	);
	LUT4 #(
		.INIT('h0001)
	) name9952 (
		_w20461_,
		_w20462_,
		_w20463_,
		_w20464_,
		_w20465_
	);
	LUT3 #(
		.INIT('h80)
	) name9953 (
		\wishbone_bd_ram_mem0_reg[153][5]/P0001 ,
		_w11959_,
		_w11968_,
		_w20466_
	);
	LUT3 #(
		.INIT('h80)
	) name9954 (
		\wishbone_bd_ram_mem0_reg[70][5]/P0001 ,
		_w11949_,
		_w11986_,
		_w20467_
	);
	LUT3 #(
		.INIT('h80)
	) name9955 (
		\wishbone_bd_ram_mem0_reg[167][5]/P0001 ,
		_w11930_,
		_w11975_,
		_w20468_
	);
	LUT3 #(
		.INIT('h80)
	) name9956 (
		\wishbone_bd_ram_mem0_reg[132][5]/P0001 ,
		_w11929_,
		_w11955_,
		_w20469_
	);
	LUT4 #(
		.INIT('h0001)
	) name9957 (
		_w20466_,
		_w20467_,
		_w20468_,
		_w20469_,
		_w20470_
	);
	LUT3 #(
		.INIT('h80)
	) name9958 (
		\wishbone_bd_ram_mem0_reg[111][5]/P0001 ,
		_w11965_,
		_w11973_,
		_w20471_
	);
	LUT3 #(
		.INIT('h80)
	) name9959 (
		\wishbone_bd_ram_mem0_reg[229][5]/P0001 ,
		_w11933_,
		_w11982_,
		_w20472_
	);
	LUT3 #(
		.INIT('h80)
	) name9960 (
		\wishbone_bd_ram_mem0_reg[164][5]/P0001 ,
		_w11929_,
		_w11930_,
		_w20473_
	);
	LUT3 #(
		.INIT('h80)
	) name9961 (
		\wishbone_bd_ram_mem0_reg[225][5]/P0001 ,
		_w11977_,
		_w11982_,
		_w20474_
	);
	LUT4 #(
		.INIT('h0001)
	) name9962 (
		_w20471_,
		_w20472_,
		_w20473_,
		_w20474_,
		_w20475_
	);
	LUT4 #(
		.INIT('h8000)
	) name9963 (
		_w20460_,
		_w20465_,
		_w20470_,
		_w20475_,
		_w20476_
	);
	LUT3 #(
		.INIT('h80)
	) name9964 (
		\wishbone_bd_ram_mem0_reg[208][5]/P0001 ,
		_w11941_,
		_w11984_,
		_w20477_
	);
	LUT3 #(
		.INIT('h80)
	) name9965 (
		\wishbone_bd_ram_mem0_reg[102][5]/P0001 ,
		_w11965_,
		_w11986_,
		_w20478_
	);
	LUT3 #(
		.INIT('h80)
	) name9966 (
		\wishbone_bd_ram_mem0_reg[174][5]/P0001 ,
		_w11930_,
		_w11948_,
		_w20479_
	);
	LUT3 #(
		.INIT('h80)
	) name9967 (
		\wishbone_bd_ram_mem0_reg[231][5]/P0001 ,
		_w11975_,
		_w11982_,
		_w20480_
	);
	LUT4 #(
		.INIT('h0001)
	) name9968 (
		_w20477_,
		_w20478_,
		_w20479_,
		_w20480_,
		_w20481_
	);
	LUT3 #(
		.INIT('h80)
	) name9969 (
		\wishbone_bd_ram_mem0_reg[206][5]/P0001 ,
		_w11945_,
		_w11948_,
		_w20482_
	);
	LUT3 #(
		.INIT('h80)
	) name9970 (
		\wishbone_bd_ram_mem0_reg[204][5]/P0001 ,
		_w11945_,
		_w11954_,
		_w20483_
	);
	LUT3 #(
		.INIT('h80)
	) name9971 (
		\wishbone_bd_ram_mem0_reg[20][5]/P0001 ,
		_w11929_,
		_w11935_,
		_w20484_
	);
	LUT3 #(
		.INIT('h80)
	) name9972 (
		\wishbone_bd_ram_mem0_reg[4][5]/P0001 ,
		_w11929_,
		_w11932_,
		_w20485_
	);
	LUT4 #(
		.INIT('h0001)
	) name9973 (
		_w20482_,
		_w20483_,
		_w20484_,
		_w20485_,
		_w20486_
	);
	LUT3 #(
		.INIT('h80)
	) name9974 (
		\wishbone_bd_ram_mem0_reg[186][5]/P0001 ,
		_w11942_,
		_w11944_,
		_w20487_
	);
	LUT3 #(
		.INIT('h80)
	) name9975 (
		\wishbone_bd_ram_mem0_reg[26][5]/P0001 ,
		_w11935_,
		_w11944_,
		_w20488_
	);
	LUT3 #(
		.INIT('h80)
	) name9976 (
		\wishbone_bd_ram_mem0_reg[134][5]/P0001 ,
		_w11955_,
		_w11986_,
		_w20489_
	);
	LUT3 #(
		.INIT('h80)
	) name9977 (
		\wishbone_bd_ram_mem0_reg[38][5]/P0001 ,
		_w11957_,
		_w11986_,
		_w20490_
	);
	LUT4 #(
		.INIT('h0001)
	) name9978 (
		_w20487_,
		_w20488_,
		_w20489_,
		_w20490_,
		_w20491_
	);
	LUT3 #(
		.INIT('h80)
	) name9979 (
		\wishbone_bd_ram_mem0_reg[171][5]/P0001 ,
		_w11930_,
		_w11936_,
		_w20492_
	);
	LUT3 #(
		.INIT('h80)
	) name9980 (
		\wishbone_bd_ram_mem0_reg[35][5]/P0001 ,
		_w11938_,
		_w11957_,
		_w20493_
	);
	LUT3 #(
		.INIT('h80)
	) name9981 (
		\wishbone_bd_ram_mem0_reg[3][5]/P0001 ,
		_w11932_,
		_w11938_,
		_w20494_
	);
	LUT3 #(
		.INIT('h80)
	) name9982 (
		\wishbone_bd_ram_mem0_reg[88][5]/P0001 ,
		_w11972_,
		_w11990_,
		_w20495_
	);
	LUT4 #(
		.INIT('h0001)
	) name9983 (
		_w20492_,
		_w20493_,
		_w20494_,
		_w20495_,
		_w20496_
	);
	LUT4 #(
		.INIT('h8000)
	) name9984 (
		_w20481_,
		_w20486_,
		_w20491_,
		_w20496_,
		_w20497_
	);
	LUT4 #(
		.INIT('h8000)
	) name9985 (
		_w20434_,
		_w20455_,
		_w20476_,
		_w20497_,
		_w20498_
	);
	LUT3 #(
		.INIT('h80)
	) name9986 (
		\wishbone_bd_ram_mem0_reg[57][5]/P0001 ,
		_w11968_,
		_w11979_,
		_w20499_
	);
	LUT3 #(
		.INIT('h80)
	) name9987 (
		\wishbone_bd_ram_mem0_reg[198][5]/P0001 ,
		_w11945_,
		_w11986_,
		_w20500_
	);
	LUT3 #(
		.INIT('h80)
	) name9988 (
		\wishbone_bd_ram_mem0_reg[242][5]/P0001 ,
		_w11952_,
		_w11963_,
		_w20501_
	);
	LUT3 #(
		.INIT('h80)
	) name9989 (
		\wishbone_bd_ram_mem0_reg[180][5]/P0001 ,
		_w11929_,
		_w11942_,
		_w20502_
	);
	LUT4 #(
		.INIT('h0001)
	) name9990 (
		_w20499_,
		_w20500_,
		_w20501_,
		_w20502_,
		_w20503_
	);
	LUT3 #(
		.INIT('h80)
	) name9991 (
		\wishbone_bd_ram_mem0_reg[127][5]/P0001 ,
		_w11973_,
		_w12012_,
		_w20504_
	);
	LUT3 #(
		.INIT('h80)
	) name9992 (
		\wishbone_bd_ram_mem0_reg[232][5]/P0001 ,
		_w11982_,
		_w11990_,
		_w20505_
	);
	LUT3 #(
		.INIT('h80)
	) name9993 (
		\wishbone_bd_ram_mem0_reg[56][5]/P0001 ,
		_w11979_,
		_w11990_,
		_w20506_
	);
	LUT3 #(
		.INIT('h80)
	) name9994 (
		\wishbone_bd_ram_mem0_reg[1][5]/P0001 ,
		_w11932_,
		_w11977_,
		_w20507_
	);
	LUT4 #(
		.INIT('h0001)
	) name9995 (
		_w20504_,
		_w20505_,
		_w20506_,
		_w20507_,
		_w20508_
	);
	LUT3 #(
		.INIT('h80)
	) name9996 (
		\wishbone_bd_ram_mem0_reg[237][5]/P0001 ,
		_w11966_,
		_w11982_,
		_w20509_
	);
	LUT3 #(
		.INIT('h80)
	) name9997 (
		\wishbone_bd_ram_mem0_reg[100][5]/P0001 ,
		_w11929_,
		_w11965_,
		_w20510_
	);
	LUT3 #(
		.INIT('h80)
	) name9998 (
		\wishbone_bd_ram_mem0_reg[154][5]/P0001 ,
		_w11944_,
		_w11959_,
		_w20511_
	);
	LUT3 #(
		.INIT('h80)
	) name9999 (
		\wishbone_bd_ram_mem0_reg[173][5]/P0001 ,
		_w11930_,
		_w11966_,
		_w20512_
	);
	LUT4 #(
		.INIT('h0001)
	) name10000 (
		_w20509_,
		_w20510_,
		_w20511_,
		_w20512_,
		_w20513_
	);
	LUT3 #(
		.INIT('h80)
	) name10001 (
		\wishbone_bd_ram_mem0_reg[91][5]/P0001 ,
		_w11936_,
		_w11972_,
		_w20514_
	);
	LUT3 #(
		.INIT('h80)
	) name10002 (
		\wishbone_bd_ram_mem0_reg[49][5]/P0001 ,
		_w11977_,
		_w11979_,
		_w20515_
	);
	LUT3 #(
		.INIT('h80)
	) name10003 (
		\wishbone_bd_ram_mem0_reg[98][5]/P0001 ,
		_w11963_,
		_w11965_,
		_w20516_
	);
	LUT3 #(
		.INIT('h80)
	) name10004 (
		\wishbone_bd_ram_mem0_reg[105][5]/P0001 ,
		_w11965_,
		_w11968_,
		_w20517_
	);
	LUT4 #(
		.INIT('h0001)
	) name10005 (
		_w20514_,
		_w20515_,
		_w20516_,
		_w20517_,
		_w20518_
	);
	LUT4 #(
		.INIT('h8000)
	) name10006 (
		_w20503_,
		_w20508_,
		_w20513_,
		_w20518_,
		_w20519_
	);
	LUT3 #(
		.INIT('h80)
	) name10007 (
		\wishbone_bd_ram_mem0_reg[61][5]/P0001 ,
		_w11966_,
		_w11979_,
		_w20520_
	);
	LUT3 #(
		.INIT('h80)
	) name10008 (
		\wishbone_bd_ram_mem0_reg[200][5]/P0001 ,
		_w11945_,
		_w11990_,
		_w20521_
	);
	LUT3 #(
		.INIT('h80)
	) name10009 (
		\wishbone_bd_ram_mem0_reg[149][5]/P0001 ,
		_w11933_,
		_w11959_,
		_w20522_
	);
	LUT3 #(
		.INIT('h80)
	) name10010 (
		\wishbone_bd_ram_mem0_reg[32][5]/P0001 ,
		_w11941_,
		_w11957_,
		_w20523_
	);
	LUT4 #(
		.INIT('h0001)
	) name10011 (
		_w20520_,
		_w20521_,
		_w20522_,
		_w20523_,
		_w20524_
	);
	LUT3 #(
		.INIT('h80)
	) name10012 (
		\wishbone_bd_ram_mem0_reg[30][5]/P0001 ,
		_w11935_,
		_w11948_,
		_w20525_
	);
	LUT3 #(
		.INIT('h80)
	) name10013 (
		\wishbone_bd_ram_mem0_reg[60][5]/P0001 ,
		_w11954_,
		_w11979_,
		_w20526_
	);
	LUT3 #(
		.INIT('h80)
	) name10014 (
		\wishbone_bd_ram_mem0_reg[33][5]/P0001 ,
		_w11957_,
		_w11977_,
		_w20527_
	);
	LUT3 #(
		.INIT('h80)
	) name10015 (
		\wishbone_bd_ram_mem0_reg[95][5]/P0001 ,
		_w11972_,
		_w11973_,
		_w20528_
	);
	LUT4 #(
		.INIT('h0001)
	) name10016 (
		_w20525_,
		_w20526_,
		_w20527_,
		_w20528_,
		_w20529_
	);
	LUT3 #(
		.INIT('h80)
	) name10017 (
		\wishbone_bd_ram_mem0_reg[50][5]/P0001 ,
		_w11963_,
		_w11979_,
		_w20530_
	);
	LUT3 #(
		.INIT('h80)
	) name10018 (
		\wishbone_bd_ram_mem0_reg[94][5]/P0001 ,
		_w11948_,
		_w11972_,
		_w20531_
	);
	LUT3 #(
		.INIT('h80)
	) name10019 (
		\wishbone_bd_ram_mem0_reg[39][5]/P0001 ,
		_w11957_,
		_w11975_,
		_w20532_
	);
	LUT3 #(
		.INIT('h80)
	) name10020 (
		\wishbone_bd_ram_mem0_reg[51][5]/P0001 ,
		_w11938_,
		_w11979_,
		_w20533_
	);
	LUT4 #(
		.INIT('h0001)
	) name10021 (
		_w20530_,
		_w20531_,
		_w20532_,
		_w20533_,
		_w20534_
	);
	LUT3 #(
		.INIT('h80)
	) name10022 (
		\wishbone_bd_ram_mem0_reg[166][5]/P0001 ,
		_w11930_,
		_w11986_,
		_w20535_
	);
	LUT3 #(
		.INIT('h80)
	) name10023 (
		\wishbone_bd_ram_mem0_reg[246][5]/P0001 ,
		_w11952_,
		_w11986_,
		_w20536_
	);
	LUT3 #(
		.INIT('h80)
	) name10024 (
		\wishbone_bd_ram_mem0_reg[175][5]/P0001 ,
		_w11930_,
		_w11973_,
		_w20537_
	);
	LUT3 #(
		.INIT('h80)
	) name10025 (
		\wishbone_bd_ram_mem0_reg[150][5]/P0001 ,
		_w11959_,
		_w11986_,
		_w20538_
	);
	LUT4 #(
		.INIT('h0001)
	) name10026 (
		_w20535_,
		_w20536_,
		_w20537_,
		_w20538_,
		_w20539_
	);
	LUT4 #(
		.INIT('h8000)
	) name10027 (
		_w20524_,
		_w20529_,
		_w20534_,
		_w20539_,
		_w20540_
	);
	LUT3 #(
		.INIT('h80)
	) name10028 (
		\wishbone_bd_ram_mem0_reg[14][5]/P0001 ,
		_w11932_,
		_w11948_,
		_w20541_
	);
	LUT3 #(
		.INIT('h80)
	) name10029 (
		\wishbone_bd_ram_mem0_reg[169][5]/P0001 ,
		_w11930_,
		_w11968_,
		_w20542_
	);
	LUT3 #(
		.INIT('h80)
	) name10030 (
		\wishbone_bd_ram_mem0_reg[143][5]/P0001 ,
		_w11955_,
		_w11973_,
		_w20543_
	);
	LUT3 #(
		.INIT('h80)
	) name10031 (
		\wishbone_bd_ram_mem0_reg[185][5]/P0001 ,
		_w11942_,
		_w11968_,
		_w20544_
	);
	LUT4 #(
		.INIT('h0001)
	) name10032 (
		_w20541_,
		_w20542_,
		_w20543_,
		_w20544_,
		_w20545_
	);
	LUT3 #(
		.INIT('h80)
	) name10033 (
		\wishbone_bd_ram_mem0_reg[106][5]/P0001 ,
		_w11944_,
		_w11965_,
		_w20546_
	);
	LUT3 #(
		.INIT('h80)
	) name10034 (
		\wishbone_bd_ram_mem0_reg[215][5]/P0001 ,
		_w11975_,
		_w11984_,
		_w20547_
	);
	LUT3 #(
		.INIT('h80)
	) name10035 (
		\wishbone_bd_ram_mem0_reg[12][5]/P0001 ,
		_w11932_,
		_w11954_,
		_w20548_
	);
	LUT3 #(
		.INIT('h80)
	) name10036 (
		\wishbone_bd_ram_mem0_reg[118][5]/P0001 ,
		_w11986_,
		_w12012_,
		_w20549_
	);
	LUT4 #(
		.INIT('h0001)
	) name10037 (
		_w20546_,
		_w20547_,
		_w20548_,
		_w20549_,
		_w20550_
	);
	LUT3 #(
		.INIT('h80)
	) name10038 (
		\wishbone_bd_ram_mem0_reg[15][5]/P0001 ,
		_w11932_,
		_w11973_,
		_w20551_
	);
	LUT3 #(
		.INIT('h80)
	) name10039 (
		\wishbone_bd_ram_mem0_reg[131][5]/P0001 ,
		_w11938_,
		_w11955_,
		_w20552_
	);
	LUT3 #(
		.INIT('h80)
	) name10040 (
		\wishbone_bd_ram_mem0_reg[172][5]/P0001 ,
		_w11930_,
		_w11954_,
		_w20553_
	);
	LUT3 #(
		.INIT('h80)
	) name10041 (
		\wishbone_bd_ram_mem0_reg[209][5]/P0001 ,
		_w11977_,
		_w11984_,
		_w20554_
	);
	LUT4 #(
		.INIT('h0001)
	) name10042 (
		_w20551_,
		_w20552_,
		_w20553_,
		_w20554_,
		_w20555_
	);
	LUT3 #(
		.INIT('h80)
	) name10043 (
		\wishbone_bd_ram_mem0_reg[120][5]/P0001 ,
		_w11990_,
		_w12012_,
		_w20556_
	);
	LUT3 #(
		.INIT('h80)
	) name10044 (
		\wishbone_bd_ram_mem0_reg[239][5]/P0001 ,
		_w11973_,
		_w11982_,
		_w20557_
	);
	LUT3 #(
		.INIT('h80)
	) name10045 (
		\wishbone_bd_ram_mem0_reg[116][5]/P0001 ,
		_w11929_,
		_w12012_,
		_w20558_
	);
	LUT3 #(
		.INIT('h80)
	) name10046 (
		\wishbone_bd_ram_mem0_reg[122][5]/P0001 ,
		_w11944_,
		_w12012_,
		_w20559_
	);
	LUT4 #(
		.INIT('h0001)
	) name10047 (
		_w20556_,
		_w20557_,
		_w20558_,
		_w20559_,
		_w20560_
	);
	LUT4 #(
		.INIT('h8000)
	) name10048 (
		_w20545_,
		_w20550_,
		_w20555_,
		_w20560_,
		_w20561_
	);
	LUT3 #(
		.INIT('h80)
	) name10049 (
		\wishbone_bd_ram_mem0_reg[64][5]/P0001 ,
		_w11941_,
		_w11949_,
		_w20562_
	);
	LUT3 #(
		.INIT('h80)
	) name10050 (
		\wishbone_bd_ram_mem0_reg[71][5]/P0001 ,
		_w11949_,
		_w11975_,
		_w20563_
	);
	LUT3 #(
		.INIT('h80)
	) name10051 (
		\wishbone_bd_ram_mem0_reg[195][5]/P0001 ,
		_w11938_,
		_w11945_,
		_w20564_
	);
	LUT3 #(
		.INIT('h80)
	) name10052 (
		\wishbone_bd_ram_mem0_reg[41][5]/P0001 ,
		_w11957_,
		_w11968_,
		_w20565_
	);
	LUT4 #(
		.INIT('h0001)
	) name10053 (
		_w20562_,
		_w20563_,
		_w20564_,
		_w20565_,
		_w20566_
	);
	LUT3 #(
		.INIT('h80)
	) name10054 (
		\wishbone_bd_ram_mem0_reg[123][5]/P0001 ,
		_w11936_,
		_w12012_,
		_w20567_
	);
	LUT3 #(
		.INIT('h80)
	) name10055 (
		\wishbone_bd_ram_mem0_reg[181][5]/P0001 ,
		_w11933_,
		_w11942_,
		_w20568_
	);
	LUT3 #(
		.INIT('h80)
	) name10056 (
		\wishbone_bd_ram_mem0_reg[28][5]/P0001 ,
		_w11935_,
		_w11954_,
		_w20569_
	);
	LUT3 #(
		.INIT('h80)
	) name10057 (
		\wishbone_bd_ram_mem0_reg[218][5]/P0001 ,
		_w11944_,
		_w11984_,
		_w20570_
	);
	LUT4 #(
		.INIT('h0001)
	) name10058 (
		_w20567_,
		_w20568_,
		_w20569_,
		_w20570_,
		_w20571_
	);
	LUT3 #(
		.INIT('h80)
	) name10059 (
		\wishbone_bd_ram_mem0_reg[247][5]/P0001 ,
		_w11952_,
		_w11975_,
		_w20572_
	);
	LUT3 #(
		.INIT('h80)
	) name10060 (
		\wishbone_bd_ram_mem0_reg[197][5]/P0001 ,
		_w11933_,
		_w11945_,
		_w20573_
	);
	LUT3 #(
		.INIT('h80)
	) name10061 (
		\wishbone_bd_ram_mem0_reg[55][5]/P0001 ,
		_w11975_,
		_w11979_,
		_w20574_
	);
	LUT3 #(
		.INIT('h80)
	) name10062 (
		\wishbone_bd_ram_mem0_reg[194][5]/P0001 ,
		_w11945_,
		_w11963_,
		_w20575_
	);
	LUT4 #(
		.INIT('h0001)
	) name10063 (
		_w20572_,
		_w20573_,
		_w20574_,
		_w20575_,
		_w20576_
	);
	LUT3 #(
		.INIT('h80)
	) name10064 (
		\wishbone_bd_ram_mem0_reg[211][5]/P0001 ,
		_w11938_,
		_w11984_,
		_w20577_
	);
	LUT3 #(
		.INIT('h80)
	) name10065 (
		\wishbone_bd_ram_mem0_reg[189][5]/P0001 ,
		_w11942_,
		_w11966_,
		_w20578_
	);
	LUT3 #(
		.INIT('h80)
	) name10066 (
		\wishbone_bd_ram_mem0_reg[146][5]/P0001 ,
		_w11959_,
		_w11963_,
		_w20579_
	);
	LUT3 #(
		.INIT('h80)
	) name10067 (
		\wishbone_bd_ram_mem0_reg[157][5]/P0001 ,
		_w11959_,
		_w11966_,
		_w20580_
	);
	LUT4 #(
		.INIT('h0001)
	) name10068 (
		_w20577_,
		_w20578_,
		_w20579_,
		_w20580_,
		_w20581_
	);
	LUT4 #(
		.INIT('h8000)
	) name10069 (
		_w20566_,
		_w20571_,
		_w20576_,
		_w20581_,
		_w20582_
	);
	LUT4 #(
		.INIT('h8000)
	) name10070 (
		_w20519_,
		_w20540_,
		_w20561_,
		_w20582_,
		_w20583_
	);
	LUT3 #(
		.INIT('h80)
	) name10071 (
		\wishbone_bd_ram_mem0_reg[52][5]/P0001 ,
		_w11929_,
		_w11979_,
		_w20584_
	);
	LUT3 #(
		.INIT('h80)
	) name10072 (
		\wishbone_bd_ram_mem0_reg[8][5]/P0001 ,
		_w11932_,
		_w11990_,
		_w20585_
	);
	LUT3 #(
		.INIT('h80)
	) name10073 (
		\wishbone_bd_ram_mem0_reg[101][5]/P0001 ,
		_w11933_,
		_w11965_,
		_w20586_
	);
	LUT3 #(
		.INIT('h80)
	) name10074 (
		\wishbone_bd_ram_mem0_reg[217][5]/P0001 ,
		_w11968_,
		_w11984_,
		_w20587_
	);
	LUT4 #(
		.INIT('h0001)
	) name10075 (
		_w20584_,
		_w20585_,
		_w20586_,
		_w20587_,
		_w20588_
	);
	LUT3 #(
		.INIT('h80)
	) name10076 (
		\wishbone_bd_ram_mem0_reg[84][5]/P0001 ,
		_w11929_,
		_w11972_,
		_w20589_
	);
	LUT3 #(
		.INIT('h80)
	) name10077 (
		\wishbone_bd_ram_mem0_reg[17][5]/P0001 ,
		_w11935_,
		_w11977_,
		_w20590_
	);
	LUT3 #(
		.INIT('h80)
	) name10078 (
		\wishbone_bd_ram_mem0_reg[252][5]/P0001 ,
		_w11952_,
		_w11954_,
		_w20591_
	);
	LUT3 #(
		.INIT('h80)
	) name10079 (
		\wishbone_bd_ram_mem0_reg[155][5]/P0001 ,
		_w11936_,
		_w11959_,
		_w20592_
	);
	LUT4 #(
		.INIT('h0001)
	) name10080 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20592_,
		_w20593_
	);
	LUT3 #(
		.INIT('h80)
	) name10081 (
		\wishbone_bd_ram_mem0_reg[89][5]/P0001 ,
		_w11968_,
		_w11972_,
		_w20594_
	);
	LUT3 #(
		.INIT('h80)
	) name10082 (
		\wishbone_bd_ram_mem0_reg[2][5]/P0001 ,
		_w11932_,
		_w11963_,
		_w20595_
	);
	LUT3 #(
		.INIT('h80)
	) name10083 (
		\wishbone_bd_ram_mem0_reg[212][5]/P0001 ,
		_w11929_,
		_w11984_,
		_w20596_
	);
	LUT3 #(
		.INIT('h80)
	) name10084 (
		\wishbone_bd_ram_mem0_reg[86][5]/P0001 ,
		_w11972_,
		_w11986_,
		_w20597_
	);
	LUT4 #(
		.INIT('h0001)
	) name10085 (
		_w20594_,
		_w20595_,
		_w20596_,
		_w20597_,
		_w20598_
	);
	LUT3 #(
		.INIT('h80)
	) name10086 (
		\wishbone_bd_ram_mem0_reg[77][5]/P0001 ,
		_w11949_,
		_w11966_,
		_w20599_
	);
	LUT3 #(
		.INIT('h80)
	) name10087 (
		\wishbone_bd_ram_mem0_reg[182][5]/P0001 ,
		_w11942_,
		_w11986_,
		_w20600_
	);
	LUT3 #(
		.INIT('h80)
	) name10088 (
		\wishbone_bd_ram_mem0_reg[158][5]/P0001 ,
		_w11948_,
		_w11959_,
		_w20601_
	);
	LUT3 #(
		.INIT('h80)
	) name10089 (
		\wishbone_bd_ram_mem0_reg[7][5]/P0001 ,
		_w11932_,
		_w11975_,
		_w20602_
	);
	LUT4 #(
		.INIT('h0001)
	) name10090 (
		_w20599_,
		_w20600_,
		_w20601_,
		_w20602_,
		_w20603_
	);
	LUT4 #(
		.INIT('h8000)
	) name10091 (
		_w20588_,
		_w20593_,
		_w20598_,
		_w20603_,
		_w20604_
	);
	LUT3 #(
		.INIT('h80)
	) name10092 (
		\wishbone_bd_ram_mem0_reg[219][5]/P0001 ,
		_w11936_,
		_w11984_,
		_w20605_
	);
	LUT3 #(
		.INIT('h80)
	) name10093 (
		\wishbone_bd_ram_mem0_reg[0][5]/P0001 ,
		_w11932_,
		_w11941_,
		_w20606_
	);
	LUT3 #(
		.INIT('h80)
	) name10094 (
		\wishbone_bd_ram_mem0_reg[79][5]/P0001 ,
		_w11949_,
		_w11973_,
		_w20607_
	);
	LUT3 #(
		.INIT('h80)
	) name10095 (
		\wishbone_bd_ram_mem0_reg[156][5]/P0001 ,
		_w11954_,
		_w11959_,
		_w20608_
	);
	LUT4 #(
		.INIT('h0001)
	) name10096 (
		_w20605_,
		_w20606_,
		_w20607_,
		_w20608_,
		_w20609_
	);
	LUT3 #(
		.INIT('h80)
	) name10097 (
		\wishbone_bd_ram_mem0_reg[250][5]/P0001 ,
		_w11944_,
		_w11952_,
		_w20610_
	);
	LUT3 #(
		.INIT('h80)
	) name10098 (
		\wishbone_bd_ram_mem0_reg[184][5]/P0001 ,
		_w11942_,
		_w11990_,
		_w20611_
	);
	LUT3 #(
		.INIT('h80)
	) name10099 (
		\wishbone_bd_ram_mem0_reg[16][5]/P0001 ,
		_w11935_,
		_w11941_,
		_w20612_
	);
	LUT3 #(
		.INIT('h80)
	) name10100 (
		\wishbone_bd_ram_mem0_reg[176][5]/P0001 ,
		_w11941_,
		_w11942_,
		_w20613_
	);
	LUT4 #(
		.INIT('h0001)
	) name10101 (
		_w20610_,
		_w20611_,
		_w20612_,
		_w20613_,
		_w20614_
	);
	LUT3 #(
		.INIT('h80)
	) name10102 (
		\wishbone_bd_ram_mem0_reg[47][5]/P0001 ,
		_w11957_,
		_w11973_,
		_w20615_
	);
	LUT3 #(
		.INIT('h80)
	) name10103 (
		\wishbone_bd_ram_mem0_reg[40][5]/P0001 ,
		_w11957_,
		_w11990_,
		_w20616_
	);
	LUT3 #(
		.INIT('h80)
	) name10104 (
		\wishbone_bd_ram_mem0_reg[115][5]/P0001 ,
		_w11938_,
		_w12012_,
		_w20617_
	);
	LUT3 #(
		.INIT('h80)
	) name10105 (
		\wishbone_bd_ram_mem0_reg[22][5]/P0001 ,
		_w11935_,
		_w11986_,
		_w20618_
	);
	LUT4 #(
		.INIT('h0001)
	) name10106 (
		_w20615_,
		_w20616_,
		_w20617_,
		_w20618_,
		_w20619_
	);
	LUT3 #(
		.INIT('h80)
	) name10107 (
		\wishbone_bd_ram_mem0_reg[66][5]/P0001 ,
		_w11949_,
		_w11963_,
		_w20620_
	);
	LUT3 #(
		.INIT('h80)
	) name10108 (
		\wishbone_bd_ram_mem0_reg[163][5]/P0001 ,
		_w11930_,
		_w11938_,
		_w20621_
	);
	LUT3 #(
		.INIT('h80)
	) name10109 (
		\wishbone_bd_ram_mem0_reg[83][5]/P0001 ,
		_w11938_,
		_w11972_,
		_w20622_
	);
	LUT3 #(
		.INIT('h80)
	) name10110 (
		\wishbone_bd_ram_mem0_reg[152][5]/P0001 ,
		_w11959_,
		_w11990_,
		_w20623_
	);
	LUT4 #(
		.INIT('h0001)
	) name10111 (
		_w20620_,
		_w20621_,
		_w20622_,
		_w20623_,
		_w20624_
	);
	LUT4 #(
		.INIT('h8000)
	) name10112 (
		_w20609_,
		_w20614_,
		_w20619_,
		_w20624_,
		_w20625_
	);
	LUT3 #(
		.INIT('h80)
	) name10113 (
		\wishbone_bd_ram_mem0_reg[253][5]/P0001 ,
		_w11952_,
		_w11966_,
		_w20626_
	);
	LUT3 #(
		.INIT('h80)
	) name10114 (
		\wishbone_bd_ram_mem0_reg[109][5]/P0001 ,
		_w11965_,
		_w11966_,
		_w20627_
	);
	LUT3 #(
		.INIT('h80)
	) name10115 (
		\wishbone_bd_ram_mem0_reg[72][5]/P0001 ,
		_w11949_,
		_w11990_,
		_w20628_
	);
	LUT3 #(
		.INIT('h80)
	) name10116 (
		\wishbone_bd_ram_mem0_reg[199][5]/P0001 ,
		_w11945_,
		_w11975_,
		_w20629_
	);
	LUT4 #(
		.INIT('h0001)
	) name10117 (
		_w20626_,
		_w20627_,
		_w20628_,
		_w20629_,
		_w20630_
	);
	LUT3 #(
		.INIT('h80)
	) name10118 (
		\wishbone_bd_ram_mem0_reg[213][5]/P0001 ,
		_w11933_,
		_w11984_,
		_w20631_
	);
	LUT3 #(
		.INIT('h80)
	) name10119 (
		\wishbone_bd_ram_mem0_reg[130][5]/P0001 ,
		_w11955_,
		_w11963_,
		_w20632_
	);
	LUT3 #(
		.INIT('h80)
	) name10120 (
		\wishbone_bd_ram_mem0_reg[54][5]/P0001 ,
		_w11979_,
		_w11986_,
		_w20633_
	);
	LUT3 #(
		.INIT('h80)
	) name10121 (
		\wishbone_bd_ram_mem0_reg[36][5]/P0001 ,
		_w11929_,
		_w11957_,
		_w20634_
	);
	LUT4 #(
		.INIT('h0001)
	) name10122 (
		_w20631_,
		_w20632_,
		_w20633_,
		_w20634_,
		_w20635_
	);
	LUT3 #(
		.INIT('h80)
	) name10123 (
		\wishbone_bd_ram_mem0_reg[234][5]/P0001 ,
		_w11944_,
		_w11982_,
		_w20636_
	);
	LUT3 #(
		.INIT('h80)
	) name10124 (
		\wishbone_bd_ram_mem0_reg[124][5]/P0001 ,
		_w11954_,
		_w12012_,
		_w20637_
	);
	LUT3 #(
		.INIT('h80)
	) name10125 (
		\wishbone_bd_ram_mem0_reg[34][5]/P0001 ,
		_w11957_,
		_w11963_,
		_w20638_
	);
	LUT3 #(
		.INIT('h80)
	) name10126 (
		\wishbone_bd_ram_mem0_reg[196][5]/P0001 ,
		_w11929_,
		_w11945_,
		_w20639_
	);
	LUT4 #(
		.INIT('h0001)
	) name10127 (
		_w20636_,
		_w20637_,
		_w20638_,
		_w20639_,
		_w20640_
	);
	LUT3 #(
		.INIT('h80)
	) name10128 (
		\wishbone_bd_ram_mem0_reg[160][5]/P0001 ,
		_w11930_,
		_w11941_,
		_w20641_
	);
	LUT3 #(
		.INIT('h80)
	) name10129 (
		\wishbone_bd_ram_mem0_reg[117][5]/P0001 ,
		_w11933_,
		_w12012_,
		_w20642_
	);
	LUT3 #(
		.INIT('h80)
	) name10130 (
		\wishbone_bd_ram_mem0_reg[137][5]/P0001 ,
		_w11955_,
		_w11968_,
		_w20643_
	);
	LUT3 #(
		.INIT('h80)
	) name10131 (
		\wishbone_bd_ram_mem0_reg[147][5]/P0001 ,
		_w11938_,
		_w11959_,
		_w20644_
	);
	LUT4 #(
		.INIT('h0001)
	) name10132 (
		_w20641_,
		_w20642_,
		_w20643_,
		_w20644_,
		_w20645_
	);
	LUT4 #(
		.INIT('h8000)
	) name10133 (
		_w20630_,
		_w20635_,
		_w20640_,
		_w20645_,
		_w20646_
	);
	LUT3 #(
		.INIT('h80)
	) name10134 (
		\wishbone_bd_ram_mem0_reg[126][5]/P0001 ,
		_w11948_,
		_w12012_,
		_w20647_
	);
	LUT3 #(
		.INIT('h80)
	) name10135 (
		\wishbone_bd_ram_mem0_reg[191][5]/P0001 ,
		_w11942_,
		_w11973_,
		_w20648_
	);
	LUT3 #(
		.INIT('h80)
	) name10136 (
		\wishbone_bd_ram_mem0_reg[45][5]/P0001 ,
		_w11957_,
		_w11966_,
		_w20649_
	);
	LUT3 #(
		.INIT('h80)
	) name10137 (
		\wishbone_bd_ram_mem0_reg[19][5]/P0001 ,
		_w11935_,
		_w11938_,
		_w20650_
	);
	LUT4 #(
		.INIT('h0001)
	) name10138 (
		_w20647_,
		_w20648_,
		_w20649_,
		_w20650_,
		_w20651_
	);
	LUT3 #(
		.INIT('h80)
	) name10139 (
		\wishbone_bd_ram_mem0_reg[230][5]/P0001 ,
		_w11982_,
		_w11986_,
		_w20652_
	);
	LUT3 #(
		.INIT('h80)
	) name10140 (
		\wishbone_bd_ram_mem0_reg[205][5]/P0001 ,
		_w11945_,
		_w11966_,
		_w20653_
	);
	LUT3 #(
		.INIT('h80)
	) name10141 (
		\wishbone_bd_ram_mem0_reg[240][5]/P0001 ,
		_w11941_,
		_w11952_,
		_w20654_
	);
	LUT3 #(
		.INIT('h80)
	) name10142 (
		\wishbone_bd_ram_mem0_reg[255][5]/P0001 ,
		_w11952_,
		_w11973_,
		_w20655_
	);
	LUT4 #(
		.INIT('h0001)
	) name10143 (
		_w20652_,
		_w20653_,
		_w20654_,
		_w20655_,
		_w20656_
	);
	LUT3 #(
		.INIT('h80)
	) name10144 (
		\wishbone_bd_ram_mem0_reg[233][5]/P0001 ,
		_w11968_,
		_w11982_,
		_w20657_
	);
	LUT3 #(
		.INIT('h80)
	) name10145 (
		\wishbone_bd_ram_mem0_reg[161][5]/P0001 ,
		_w11930_,
		_w11977_,
		_w20658_
	);
	LUT3 #(
		.INIT('h80)
	) name10146 (
		\wishbone_bd_ram_mem0_reg[6][5]/P0001 ,
		_w11932_,
		_w11986_,
		_w20659_
	);
	LUT3 #(
		.INIT('h80)
	) name10147 (
		\wishbone_bd_ram_mem0_reg[188][5]/P0001 ,
		_w11942_,
		_w11954_,
		_w20660_
	);
	LUT4 #(
		.INIT('h0001)
	) name10148 (
		_w20657_,
		_w20658_,
		_w20659_,
		_w20660_,
		_w20661_
	);
	LUT3 #(
		.INIT('h80)
	) name10149 (
		\wishbone_bd_ram_mem0_reg[119][5]/P0001 ,
		_w11975_,
		_w12012_,
		_w20662_
	);
	LUT3 #(
		.INIT('h80)
	) name10150 (
		\wishbone_bd_ram_mem0_reg[148][5]/P0001 ,
		_w11929_,
		_w11959_,
		_w20663_
	);
	LUT3 #(
		.INIT('h80)
	) name10151 (
		\wishbone_bd_ram_mem0_reg[21][5]/P0001 ,
		_w11933_,
		_w11935_,
		_w20664_
	);
	LUT3 #(
		.INIT('h80)
	) name10152 (
		\wishbone_bd_ram_mem0_reg[68][5]/P0001 ,
		_w11929_,
		_w11949_,
		_w20665_
	);
	LUT4 #(
		.INIT('h0001)
	) name10153 (
		_w20662_,
		_w20663_,
		_w20664_,
		_w20665_,
		_w20666_
	);
	LUT4 #(
		.INIT('h8000)
	) name10154 (
		_w20651_,
		_w20656_,
		_w20661_,
		_w20666_,
		_w20667_
	);
	LUT4 #(
		.INIT('h8000)
	) name10155 (
		_w20604_,
		_w20625_,
		_w20646_,
		_w20667_,
		_w20668_
	);
	LUT3 #(
		.INIT('h80)
	) name10156 (
		\wishbone_bd_ram_mem0_reg[62][5]/P0001 ,
		_w11948_,
		_w11979_,
		_w20669_
	);
	LUT3 #(
		.INIT('h80)
	) name10157 (
		\wishbone_bd_ram_mem0_reg[112][5]/P0001 ,
		_w11941_,
		_w12012_,
		_w20670_
	);
	LUT3 #(
		.INIT('h80)
	) name10158 (
		\wishbone_bd_ram_mem0_reg[92][5]/P0001 ,
		_w11954_,
		_w11972_,
		_w20671_
	);
	LUT3 #(
		.INIT('h80)
	) name10159 (
		\wishbone_bd_ram_mem0_reg[168][5]/P0001 ,
		_w11930_,
		_w11990_,
		_w20672_
	);
	LUT4 #(
		.INIT('h0001)
	) name10160 (
		_w20669_,
		_w20670_,
		_w20671_,
		_w20672_,
		_w20673_
	);
	LUT3 #(
		.INIT('h80)
	) name10161 (
		\wishbone_bd_ram_mem0_reg[107][5]/P0001 ,
		_w11936_,
		_w11965_,
		_w20674_
	);
	LUT3 #(
		.INIT('h80)
	) name10162 (
		\wishbone_bd_ram_mem0_reg[165][5]/P0001 ,
		_w11930_,
		_w11933_,
		_w20675_
	);
	LUT3 #(
		.INIT('h80)
	) name10163 (
		\wishbone_bd_ram_mem0_reg[128][5]/P0001 ,
		_w11941_,
		_w11955_,
		_w20676_
	);
	LUT3 #(
		.INIT('h80)
	) name10164 (
		\wishbone_bd_ram_mem0_reg[254][5]/P0001 ,
		_w11948_,
		_w11952_,
		_w20677_
	);
	LUT4 #(
		.INIT('h0001)
	) name10165 (
		_w20674_,
		_w20675_,
		_w20676_,
		_w20677_,
		_w20678_
	);
	LUT3 #(
		.INIT('h80)
	) name10166 (
		\wishbone_bd_ram_mem0_reg[81][5]/P0001 ,
		_w11972_,
		_w11977_,
		_w20679_
	);
	LUT3 #(
		.INIT('h80)
	) name10167 (
		\wishbone_bd_ram_mem0_reg[178][5]/P0001 ,
		_w11942_,
		_w11963_,
		_w20680_
	);
	LUT3 #(
		.INIT('h80)
	) name10168 (
		\wishbone_bd_ram_mem0_reg[11][5]/P0001 ,
		_w11932_,
		_w11936_,
		_w20681_
	);
	LUT3 #(
		.INIT('h80)
	) name10169 (
		\wishbone_bd_ram_mem0_reg[5][5]/P0001 ,
		_w11932_,
		_w11933_,
		_w20682_
	);
	LUT4 #(
		.INIT('h0001)
	) name10170 (
		_w20679_,
		_w20680_,
		_w20681_,
		_w20682_,
		_w20683_
	);
	LUT3 #(
		.INIT('h80)
	) name10171 (
		\wishbone_bd_ram_mem0_reg[46][5]/P0001 ,
		_w11948_,
		_w11957_,
		_w20684_
	);
	LUT3 #(
		.INIT('h80)
	) name10172 (
		\wishbone_bd_ram_mem0_reg[24][5]/P0001 ,
		_w11935_,
		_w11990_,
		_w20685_
	);
	LUT3 #(
		.INIT('h80)
	) name10173 (
		\wishbone_bd_ram_mem0_reg[59][5]/P0001 ,
		_w11936_,
		_w11979_,
		_w20686_
	);
	LUT3 #(
		.INIT('h80)
	) name10174 (
		\wishbone_bd_ram_mem0_reg[135][5]/P0001 ,
		_w11955_,
		_w11975_,
		_w20687_
	);
	LUT4 #(
		.INIT('h0001)
	) name10175 (
		_w20684_,
		_w20685_,
		_w20686_,
		_w20687_,
		_w20688_
	);
	LUT4 #(
		.INIT('h8000)
	) name10176 (
		_w20673_,
		_w20678_,
		_w20683_,
		_w20688_,
		_w20689_
	);
	LUT3 #(
		.INIT('h80)
	) name10177 (
		\wishbone_bd_ram_mem0_reg[192][5]/P0001 ,
		_w11941_,
		_w11945_,
		_w20690_
	);
	LUT3 #(
		.INIT('h80)
	) name10178 (
		\wishbone_bd_ram_mem0_reg[25][5]/P0001 ,
		_w11935_,
		_w11968_,
		_w20691_
	);
	LUT3 #(
		.INIT('h80)
	) name10179 (
		\wishbone_bd_ram_mem0_reg[226][5]/P0001 ,
		_w11963_,
		_w11982_,
		_w20692_
	);
	LUT3 #(
		.INIT('h80)
	) name10180 (
		\wishbone_bd_ram_mem0_reg[144][5]/P0001 ,
		_w11941_,
		_w11959_,
		_w20693_
	);
	LUT4 #(
		.INIT('h0001)
	) name10181 (
		_w20690_,
		_w20691_,
		_w20692_,
		_w20693_,
		_w20694_
	);
	LUT3 #(
		.INIT('h80)
	) name10182 (
		\wishbone_bd_ram_mem0_reg[151][5]/P0001 ,
		_w11959_,
		_w11975_,
		_w20695_
	);
	LUT3 #(
		.INIT('h80)
	) name10183 (
		\wishbone_bd_ram_mem0_reg[129][5]/P0001 ,
		_w11955_,
		_w11977_,
		_w20696_
	);
	LUT3 #(
		.INIT('h80)
	) name10184 (
		\wishbone_bd_ram_mem0_reg[31][5]/P0001 ,
		_w11935_,
		_w11973_,
		_w20697_
	);
	LUT3 #(
		.INIT('h80)
	) name10185 (
		\wishbone_bd_ram_mem0_reg[75][5]/P0001 ,
		_w11936_,
		_w11949_,
		_w20698_
	);
	LUT4 #(
		.INIT('h0001)
	) name10186 (
		_w20695_,
		_w20696_,
		_w20697_,
		_w20698_,
		_w20699_
	);
	LUT3 #(
		.INIT('h80)
	) name10187 (
		\wishbone_bd_ram_mem0_reg[114][5]/P0001 ,
		_w11963_,
		_w12012_,
		_w20700_
	);
	LUT3 #(
		.INIT('h80)
	) name10188 (
		\wishbone_bd_ram_mem0_reg[228][5]/P0001 ,
		_w11929_,
		_w11982_,
		_w20701_
	);
	LUT3 #(
		.INIT('h80)
	) name10189 (
		\wishbone_bd_ram_mem0_reg[110][5]/P0001 ,
		_w11948_,
		_w11965_,
		_w20702_
	);
	LUT3 #(
		.INIT('h80)
	) name10190 (
		\wishbone_bd_ram_mem0_reg[78][5]/P0001 ,
		_w11948_,
		_w11949_,
		_w20703_
	);
	LUT4 #(
		.INIT('h0001)
	) name10191 (
		_w20700_,
		_w20701_,
		_w20702_,
		_w20703_,
		_w20704_
	);
	LUT3 #(
		.INIT('h80)
	) name10192 (
		\wishbone_bd_ram_mem0_reg[224][5]/P0001 ,
		_w11941_,
		_w11982_,
		_w20705_
	);
	LUT3 #(
		.INIT('h80)
	) name10193 (
		\wishbone_bd_ram_mem0_reg[85][5]/P0001 ,
		_w11933_,
		_w11972_,
		_w20706_
	);
	LUT3 #(
		.INIT('h80)
	) name10194 (
		\wishbone_bd_ram_mem0_reg[67][5]/P0001 ,
		_w11938_,
		_w11949_,
		_w20707_
	);
	LUT3 #(
		.INIT('h80)
	) name10195 (
		\wishbone_bd_ram_mem0_reg[142][5]/P0001 ,
		_w11948_,
		_w11955_,
		_w20708_
	);
	LUT4 #(
		.INIT('h0001)
	) name10196 (
		_w20705_,
		_w20706_,
		_w20707_,
		_w20708_,
		_w20709_
	);
	LUT4 #(
		.INIT('h8000)
	) name10197 (
		_w20694_,
		_w20699_,
		_w20704_,
		_w20709_,
		_w20710_
	);
	LUT3 #(
		.INIT('h80)
	) name10198 (
		\wishbone_bd_ram_mem0_reg[140][5]/P0001 ,
		_w11954_,
		_w11955_,
		_w20711_
	);
	LUT3 #(
		.INIT('h80)
	) name10199 (
		\wishbone_bd_ram_mem0_reg[69][5]/P0001 ,
		_w11933_,
		_w11949_,
		_w20712_
	);
	LUT3 #(
		.INIT('h80)
	) name10200 (
		\wishbone_bd_ram_mem0_reg[244][5]/P0001 ,
		_w11929_,
		_w11952_,
		_w20713_
	);
	LUT3 #(
		.INIT('h80)
	) name10201 (
		\wishbone_bd_ram_mem0_reg[202][5]/P0001 ,
		_w11944_,
		_w11945_,
		_w20714_
	);
	LUT4 #(
		.INIT('h0001)
	) name10202 (
		_w20711_,
		_w20712_,
		_w20713_,
		_w20714_,
		_w20715_
	);
	LUT3 #(
		.INIT('h80)
	) name10203 (
		\wishbone_bd_ram_mem0_reg[177][5]/P0001 ,
		_w11942_,
		_w11977_,
		_w20716_
	);
	LUT3 #(
		.INIT('h80)
	) name10204 (
		\wishbone_bd_ram_mem0_reg[133][5]/P0001 ,
		_w11933_,
		_w11955_,
		_w20717_
	);
	LUT3 #(
		.INIT('h80)
	) name10205 (
		\wishbone_bd_ram_mem0_reg[87][5]/P0001 ,
		_w11972_,
		_w11975_,
		_w20718_
	);
	LUT3 #(
		.INIT('h80)
	) name10206 (
		\wishbone_bd_ram_mem0_reg[179][5]/P0001 ,
		_w11938_,
		_w11942_,
		_w20719_
	);
	LUT4 #(
		.INIT('h0001)
	) name10207 (
		_w20716_,
		_w20717_,
		_w20718_,
		_w20719_,
		_w20720_
	);
	LUT3 #(
		.INIT('h80)
	) name10208 (
		\wishbone_bd_ram_mem0_reg[42][5]/P0001 ,
		_w11944_,
		_w11957_,
		_w20721_
	);
	LUT3 #(
		.INIT('h80)
	) name10209 (
		\wishbone_bd_ram_mem0_reg[10][5]/P0001 ,
		_w11932_,
		_w11944_,
		_w20722_
	);
	LUT3 #(
		.INIT('h80)
	) name10210 (
		\wishbone_bd_ram_mem0_reg[27][5]/P0001 ,
		_w11935_,
		_w11936_,
		_w20723_
	);
	LUT3 #(
		.INIT('h80)
	) name10211 (
		\wishbone_bd_ram_mem0_reg[162][5]/P0001 ,
		_w11930_,
		_w11963_,
		_w20724_
	);
	LUT4 #(
		.INIT('h0001)
	) name10212 (
		_w20721_,
		_w20722_,
		_w20723_,
		_w20724_,
		_w20725_
	);
	LUT3 #(
		.INIT('h80)
	) name10213 (
		\wishbone_bd_ram_mem0_reg[190][5]/P0001 ,
		_w11942_,
		_w11948_,
		_w20726_
	);
	LUT3 #(
		.INIT('h80)
	) name10214 (
		\wishbone_bd_ram_mem0_reg[103][5]/P0001 ,
		_w11965_,
		_w11975_,
		_w20727_
	);
	LUT3 #(
		.INIT('h80)
	) name10215 (
		\wishbone_bd_ram_mem0_reg[221][5]/P0001 ,
		_w11966_,
		_w11984_,
		_w20728_
	);
	LUT3 #(
		.INIT('h80)
	) name10216 (
		\wishbone_bd_ram_mem0_reg[9][5]/P0001 ,
		_w11932_,
		_w11968_,
		_w20729_
	);
	LUT4 #(
		.INIT('h0001)
	) name10217 (
		_w20726_,
		_w20727_,
		_w20728_,
		_w20729_,
		_w20730_
	);
	LUT4 #(
		.INIT('h8000)
	) name10218 (
		_w20715_,
		_w20720_,
		_w20725_,
		_w20730_,
		_w20731_
	);
	LUT3 #(
		.INIT('h80)
	) name10219 (
		\wishbone_bd_ram_mem0_reg[104][5]/P0001 ,
		_w11965_,
		_w11990_,
		_w20732_
	);
	LUT3 #(
		.INIT('h80)
	) name10220 (
		\wishbone_bd_ram_mem0_reg[63][5]/P0001 ,
		_w11973_,
		_w11979_,
		_w20733_
	);
	LUT3 #(
		.INIT('h80)
	) name10221 (
		\wishbone_bd_ram_mem0_reg[90][5]/P0001 ,
		_w11944_,
		_w11972_,
		_w20734_
	);
	LUT3 #(
		.INIT('h80)
	) name10222 (
		\wishbone_bd_ram_mem0_reg[96][5]/P0001 ,
		_w11941_,
		_w11965_,
		_w20735_
	);
	LUT4 #(
		.INIT('h0001)
	) name10223 (
		_w20732_,
		_w20733_,
		_w20734_,
		_w20735_,
		_w20736_
	);
	LUT3 #(
		.INIT('h80)
	) name10224 (
		\wishbone_bd_ram_mem0_reg[251][5]/P0001 ,
		_w11936_,
		_w11952_,
		_w20737_
	);
	LUT3 #(
		.INIT('h80)
	) name10225 (
		\wishbone_bd_ram_mem0_reg[235][5]/P0001 ,
		_w11936_,
		_w11982_,
		_w20738_
	);
	LUT3 #(
		.INIT('h80)
	) name10226 (
		\wishbone_bd_ram_mem0_reg[53][5]/P0001 ,
		_w11933_,
		_w11979_,
		_w20739_
	);
	LUT3 #(
		.INIT('h80)
	) name10227 (
		\wishbone_bd_ram_mem0_reg[223][5]/P0001 ,
		_w11973_,
		_w11984_,
		_w20740_
	);
	LUT4 #(
		.INIT('h0001)
	) name10228 (
		_w20737_,
		_w20738_,
		_w20739_,
		_w20740_,
		_w20741_
	);
	LUT3 #(
		.INIT('h80)
	) name10229 (
		\wishbone_bd_ram_mem0_reg[249][5]/P0001 ,
		_w11952_,
		_w11968_,
		_w20742_
	);
	LUT3 #(
		.INIT('h80)
	) name10230 (
		\wishbone_bd_ram_mem0_reg[238][5]/P0001 ,
		_w11948_,
		_w11982_,
		_w20743_
	);
	LUT3 #(
		.INIT('h80)
	) name10231 (
		\wishbone_bd_ram_mem0_reg[139][5]/P0001 ,
		_w11936_,
		_w11955_,
		_w20744_
	);
	LUT3 #(
		.INIT('h80)
	) name10232 (
		\wishbone_bd_ram_mem0_reg[97][5]/P0001 ,
		_w11965_,
		_w11977_,
		_w20745_
	);
	LUT4 #(
		.INIT('h0001)
	) name10233 (
		_w20742_,
		_w20743_,
		_w20744_,
		_w20745_,
		_w20746_
	);
	LUT3 #(
		.INIT('h80)
	) name10234 (
		\wishbone_bd_ram_mem0_reg[82][5]/P0001 ,
		_w11963_,
		_w11972_,
		_w20747_
	);
	LUT3 #(
		.INIT('h80)
	) name10235 (
		\wishbone_bd_ram_mem0_reg[222][5]/P0001 ,
		_w11948_,
		_w11984_,
		_w20748_
	);
	LUT3 #(
		.INIT('h80)
	) name10236 (
		\wishbone_bd_ram_mem0_reg[58][5]/P0001 ,
		_w11944_,
		_w11979_,
		_w20749_
	);
	LUT3 #(
		.INIT('h80)
	) name10237 (
		\wishbone_bd_ram_mem0_reg[113][5]/P0001 ,
		_w11977_,
		_w12012_,
		_w20750_
	);
	LUT4 #(
		.INIT('h0001)
	) name10238 (
		_w20747_,
		_w20748_,
		_w20749_,
		_w20750_,
		_w20751_
	);
	LUT4 #(
		.INIT('h8000)
	) name10239 (
		_w20736_,
		_w20741_,
		_w20746_,
		_w20751_,
		_w20752_
	);
	LUT4 #(
		.INIT('h8000)
	) name10240 (
		_w20689_,
		_w20710_,
		_w20731_,
		_w20752_,
		_w20753_
	);
	LUT4 #(
		.INIT('h8000)
	) name10241 (
		_w20498_,
		_w20583_,
		_w20668_,
		_w20753_,
		_w20754_
	);
	LUT3 #(
		.INIT('h15)
	) name10242 (
		wb_rst_i_pad,
		_w20391_,
		_w20412_,
		_w20755_
	);
	LUT3 #(
		.INIT('hba)
	) name10243 (
		_w20413_,
		_w20754_,
		_w20755_,
		_w20756_
	);
	LUT4 #(
		.INIT('h0002)
	) name10244 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w20757_
	);
	LUT3 #(
		.INIT('h80)
	) name10245 (
		_w18757_,
		_w18758_,
		_w20757_,
		_w20758_
	);
	LUT3 #(
		.INIT('h80)
	) name10246 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131 ,
		_w18798_,
		_w18801_,
		_w20759_
	);
	LUT3 #(
		.INIT('h80)
	) name10247 (
		\ethreg1_MIIRX_DATA_DataOut_reg[7]/NET0131 ,
		_w18785_,
		_w18786_,
		_w20760_
	);
	LUT4 #(
		.INIT('h0008)
	) name10248 (
		\ethreg1_RXHASH0_0_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w20761_
	);
	LUT3 #(
		.INIT('h80)
	) name10249 (
		_w18757_,
		_w18758_,
		_w20761_,
		_w20762_
	);
	LUT4 #(
		.INIT('h0001)
	) name10250 (
		_w20758_,
		_w20759_,
		_w20760_,
		_w20762_,
		_w20763_
	);
	LUT3 #(
		.INIT('h80)
	) name10251 (
		\ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131 ,
		_w18786_,
		_w18801_,
		_w20764_
	);
	LUT3 #(
		.INIT('h80)
	) name10252 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		_w18800_,
		_w18801_,
		_w20765_
	);
	LUT2 #(
		.INIT('h1)
	) name10253 (
		_w20764_,
		_w20765_,
		_w20766_
	);
	LUT3 #(
		.INIT('h02)
	) name10254 (
		_w18752_,
		_w20764_,
		_w20765_,
		_w20767_
	);
	LUT3 #(
		.INIT('h80)
	) name10255 (
		\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 ,
		_w18753_,
		_w18754_,
		_w20768_
	);
	LUT4 #(
		.INIT('h0008)
	) name10256 (
		\ethreg1_RXHASH1_0_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w20769_
	);
	LUT4 #(
		.INIT('h0002)
	) name10257 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w20770_
	);
	LUT4 #(
		.INIT('h777f)
	) name10258 (
		_w18757_,
		_w18762_,
		_w20769_,
		_w20770_,
		_w20771_
	);
	LUT4 #(
		.INIT('h0020)
	) name10259 (
		\ethreg1_TXCTRL_0_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w20772_
	);
	LUT3 #(
		.INIT('h80)
	) name10260 (
		_w18757_,
		_w18758_,
		_w20772_,
		_w20773_
	);
	LUT3 #(
		.INIT('h80)
	) name10261 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[7]/NET0131 ,
		_w18798_,
		_w18805_,
		_w20774_
	);
	LUT4 #(
		.INIT('h0004)
	) name10262 (
		_w20768_,
		_w20771_,
		_w20773_,
		_w20774_,
		_w20775_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10263 (
		_w18752_,
		_w20763_,
		_w20766_,
		_w20775_,
		_w20776_
	);
	LUT3 #(
		.INIT('h80)
	) name10264 (
		\wishbone_bd_ram_mem0_reg[49][7]/P0001 ,
		_w11977_,
		_w11979_,
		_w20777_
	);
	LUT3 #(
		.INIT('h80)
	) name10265 (
		\wishbone_bd_ram_mem0_reg[69][7]/P0001 ,
		_w11933_,
		_w11949_,
		_w20778_
	);
	LUT3 #(
		.INIT('h80)
	) name10266 (
		\wishbone_bd_ram_mem0_reg[21][7]/P0001 ,
		_w11933_,
		_w11935_,
		_w20779_
	);
	LUT3 #(
		.INIT('h80)
	) name10267 (
		\wishbone_bd_ram_mem0_reg[105][7]/P0001 ,
		_w11965_,
		_w11968_,
		_w20780_
	);
	LUT4 #(
		.INIT('h0001)
	) name10268 (
		_w20777_,
		_w20778_,
		_w20779_,
		_w20780_,
		_w20781_
	);
	LUT3 #(
		.INIT('h80)
	) name10269 (
		\wishbone_bd_ram_mem0_reg[222][7]/P0001 ,
		_w11948_,
		_w11984_,
		_w20782_
	);
	LUT3 #(
		.INIT('h80)
	) name10270 (
		\wishbone_bd_ram_mem0_reg[193][7]/P0001 ,
		_w11945_,
		_w11977_,
		_w20783_
	);
	LUT3 #(
		.INIT('h80)
	) name10271 (
		\wishbone_bd_ram_mem0_reg[85][7]/P0001 ,
		_w11933_,
		_w11972_,
		_w20784_
	);
	LUT3 #(
		.INIT('h80)
	) name10272 (
		\wishbone_bd_ram_mem0_reg[242][7]/P0001 ,
		_w11952_,
		_w11963_,
		_w20785_
	);
	LUT4 #(
		.INIT('h0001)
	) name10273 (
		_w20782_,
		_w20783_,
		_w20784_,
		_w20785_,
		_w20786_
	);
	LUT3 #(
		.INIT('h80)
	) name10274 (
		\wishbone_bd_ram_mem0_reg[240][7]/P0001 ,
		_w11941_,
		_w11952_,
		_w20787_
	);
	LUT3 #(
		.INIT('h80)
	) name10275 (
		\wishbone_bd_ram_mem0_reg[183][7]/P0001 ,
		_w11942_,
		_w11975_,
		_w20788_
	);
	LUT3 #(
		.INIT('h80)
	) name10276 (
		\wishbone_bd_ram_mem0_reg[118][7]/P0001 ,
		_w11986_,
		_w12012_,
		_w20789_
	);
	LUT3 #(
		.INIT('h80)
	) name10277 (
		\wishbone_bd_ram_mem0_reg[213][7]/P0001 ,
		_w11933_,
		_w11984_,
		_w20790_
	);
	LUT4 #(
		.INIT('h0001)
	) name10278 (
		_w20787_,
		_w20788_,
		_w20789_,
		_w20790_,
		_w20791_
	);
	LUT3 #(
		.INIT('h80)
	) name10279 (
		\wishbone_bd_ram_mem0_reg[116][7]/P0001 ,
		_w11929_,
		_w12012_,
		_w20792_
	);
	LUT3 #(
		.INIT('h80)
	) name10280 (
		\wishbone_bd_ram_mem0_reg[248][7]/P0001 ,
		_w11952_,
		_w11990_,
		_w20793_
	);
	LUT3 #(
		.INIT('h80)
	) name10281 (
		\wishbone_bd_ram_mem0_reg[28][7]/P0001 ,
		_w11935_,
		_w11954_,
		_w20794_
	);
	LUT3 #(
		.INIT('h80)
	) name10282 (
		\wishbone_bd_ram_mem0_reg[144][7]/P0001 ,
		_w11941_,
		_w11959_,
		_w20795_
	);
	LUT4 #(
		.INIT('h0001)
	) name10283 (
		_w20792_,
		_w20793_,
		_w20794_,
		_w20795_,
		_w20796_
	);
	LUT4 #(
		.INIT('h8000)
	) name10284 (
		_w20781_,
		_w20786_,
		_w20791_,
		_w20796_,
		_w20797_
	);
	LUT3 #(
		.INIT('h80)
	) name10285 (
		\wishbone_bd_ram_mem0_reg[156][7]/P0001 ,
		_w11954_,
		_w11959_,
		_w20798_
	);
	LUT3 #(
		.INIT('h80)
	) name10286 (
		\wishbone_bd_ram_mem0_reg[153][7]/P0001 ,
		_w11959_,
		_w11968_,
		_w20799_
	);
	LUT3 #(
		.INIT('h80)
	) name10287 (
		\wishbone_bd_ram_mem0_reg[44][7]/P0001 ,
		_w11954_,
		_w11957_,
		_w20800_
	);
	LUT3 #(
		.INIT('h80)
	) name10288 (
		\wishbone_bd_ram_mem0_reg[59][7]/P0001 ,
		_w11936_,
		_w11979_,
		_w20801_
	);
	LUT4 #(
		.INIT('h0001)
	) name10289 (
		_w20798_,
		_w20799_,
		_w20800_,
		_w20801_,
		_w20802_
	);
	LUT3 #(
		.INIT('h80)
	) name10290 (
		\wishbone_bd_ram_mem0_reg[176][7]/P0001 ,
		_w11941_,
		_w11942_,
		_w20803_
	);
	LUT3 #(
		.INIT('h80)
	) name10291 (
		\wishbone_bd_ram_mem0_reg[235][7]/P0001 ,
		_w11936_,
		_w11982_,
		_w20804_
	);
	LUT3 #(
		.INIT('h80)
	) name10292 (
		\wishbone_bd_ram_mem0_reg[163][7]/P0001 ,
		_w11930_,
		_w11938_,
		_w20805_
	);
	LUT3 #(
		.INIT('h80)
	) name10293 (
		\wishbone_bd_ram_mem0_reg[9][7]/P0001 ,
		_w11932_,
		_w11968_,
		_w20806_
	);
	LUT4 #(
		.INIT('h0001)
	) name10294 (
		_w20803_,
		_w20804_,
		_w20805_,
		_w20806_,
		_w20807_
	);
	LUT3 #(
		.INIT('h80)
	) name10295 (
		\wishbone_bd_ram_mem0_reg[166][7]/P0001 ,
		_w11930_,
		_w11986_,
		_w20808_
	);
	LUT3 #(
		.INIT('h80)
	) name10296 (
		\wishbone_bd_ram_mem0_reg[251][7]/P0001 ,
		_w11936_,
		_w11952_,
		_w20809_
	);
	LUT3 #(
		.INIT('h80)
	) name10297 (
		\wishbone_bd_ram_mem0_reg[178][7]/P0001 ,
		_w11942_,
		_w11963_,
		_w20810_
	);
	LUT3 #(
		.INIT('h80)
	) name10298 (
		\wishbone_bd_ram_mem0_reg[37][7]/P0001 ,
		_w11933_,
		_w11957_,
		_w20811_
	);
	LUT4 #(
		.INIT('h0001)
	) name10299 (
		_w20808_,
		_w20809_,
		_w20810_,
		_w20811_,
		_w20812_
	);
	LUT3 #(
		.INIT('h80)
	) name10300 (
		\wishbone_bd_ram_mem0_reg[17][7]/P0001 ,
		_w11935_,
		_w11977_,
		_w20813_
	);
	LUT3 #(
		.INIT('h80)
	) name10301 (
		\wishbone_bd_ram_mem0_reg[170][7]/P0001 ,
		_w11930_,
		_w11944_,
		_w20814_
	);
	LUT3 #(
		.INIT('h80)
	) name10302 (
		\wishbone_bd_ram_mem0_reg[192][7]/P0001 ,
		_w11941_,
		_w11945_,
		_w20815_
	);
	LUT3 #(
		.INIT('h80)
	) name10303 (
		\wishbone_bd_ram_mem0_reg[207][7]/P0001 ,
		_w11945_,
		_w11973_,
		_w20816_
	);
	LUT4 #(
		.INIT('h0001)
	) name10304 (
		_w20813_,
		_w20814_,
		_w20815_,
		_w20816_,
		_w20817_
	);
	LUT4 #(
		.INIT('h8000)
	) name10305 (
		_w20802_,
		_w20807_,
		_w20812_,
		_w20817_,
		_w20818_
	);
	LUT3 #(
		.INIT('h80)
	) name10306 (
		\wishbone_bd_ram_mem0_reg[244][7]/P0001 ,
		_w11929_,
		_w11952_,
		_w20819_
	);
	LUT3 #(
		.INIT('h80)
	) name10307 (
		\wishbone_bd_ram_mem0_reg[101][7]/P0001 ,
		_w11933_,
		_w11965_,
		_w20820_
	);
	LUT3 #(
		.INIT('h80)
	) name10308 (
		\wishbone_bd_ram_mem0_reg[169][7]/P0001 ,
		_w11930_,
		_w11968_,
		_w20821_
	);
	LUT3 #(
		.INIT('h80)
	) name10309 (
		\wishbone_bd_ram_mem0_reg[104][7]/P0001 ,
		_w11965_,
		_w11990_,
		_w20822_
	);
	LUT4 #(
		.INIT('h0001)
	) name10310 (
		_w20819_,
		_w20820_,
		_w20821_,
		_w20822_,
		_w20823_
	);
	LUT3 #(
		.INIT('h80)
	) name10311 (
		\wishbone_bd_ram_mem0_reg[161][7]/P0001 ,
		_w11930_,
		_w11977_,
		_w20824_
	);
	LUT3 #(
		.INIT('h80)
	) name10312 (
		\wishbone_bd_ram_mem0_reg[173][7]/P0001 ,
		_w11930_,
		_w11966_,
		_w20825_
	);
	LUT3 #(
		.INIT('h80)
	) name10313 (
		\wishbone_bd_ram_mem0_reg[233][7]/P0001 ,
		_w11968_,
		_w11982_,
		_w20826_
	);
	LUT3 #(
		.INIT('h80)
	) name10314 (
		\wishbone_bd_ram_mem0_reg[98][7]/P0001 ,
		_w11963_,
		_w11965_,
		_w20827_
	);
	LUT4 #(
		.INIT('h0001)
	) name10315 (
		_w20824_,
		_w20825_,
		_w20826_,
		_w20827_,
		_w20828_
	);
	LUT3 #(
		.INIT('h80)
	) name10316 (
		\wishbone_bd_ram_mem0_reg[243][7]/P0001 ,
		_w11938_,
		_w11952_,
		_w20829_
	);
	LUT3 #(
		.INIT('h80)
	) name10317 (
		\wishbone_bd_ram_mem0_reg[19][7]/P0001 ,
		_w11935_,
		_w11938_,
		_w20830_
	);
	LUT3 #(
		.INIT('h80)
	) name10318 (
		\wishbone_bd_ram_mem0_reg[190][7]/P0001 ,
		_w11942_,
		_w11948_,
		_w20831_
	);
	LUT3 #(
		.INIT('h80)
	) name10319 (
		\wishbone_bd_ram_mem0_reg[188][7]/P0001 ,
		_w11942_,
		_w11954_,
		_w20832_
	);
	LUT4 #(
		.INIT('h0001)
	) name10320 (
		_w20829_,
		_w20830_,
		_w20831_,
		_w20832_,
		_w20833_
	);
	LUT3 #(
		.INIT('h80)
	) name10321 (
		\wishbone_bd_ram_mem0_reg[112][7]/P0001 ,
		_w11941_,
		_w12012_,
		_w20834_
	);
	LUT3 #(
		.INIT('h80)
	) name10322 (
		\wishbone_bd_ram_mem0_reg[252][7]/P0001 ,
		_w11952_,
		_w11954_,
		_w20835_
	);
	LUT3 #(
		.INIT('h80)
	) name10323 (
		\wishbone_bd_ram_mem0_reg[60][7]/P0001 ,
		_w11954_,
		_w11979_,
		_w20836_
	);
	LUT3 #(
		.INIT('h80)
	) name10324 (
		\wishbone_bd_ram_mem0_reg[181][7]/P0001 ,
		_w11933_,
		_w11942_,
		_w20837_
	);
	LUT4 #(
		.INIT('h0001)
	) name10325 (
		_w20834_,
		_w20835_,
		_w20836_,
		_w20837_,
		_w20838_
	);
	LUT4 #(
		.INIT('h8000)
	) name10326 (
		_w20823_,
		_w20828_,
		_w20833_,
		_w20838_,
		_w20839_
	);
	LUT3 #(
		.INIT('h80)
	) name10327 (
		\wishbone_bd_ram_mem0_reg[218][7]/P0001 ,
		_w11944_,
		_w11984_,
		_w20840_
	);
	LUT3 #(
		.INIT('h80)
	) name10328 (
		\wishbone_bd_ram_mem0_reg[130][7]/P0001 ,
		_w11955_,
		_w11963_,
		_w20841_
	);
	LUT3 #(
		.INIT('h80)
	) name10329 (
		\wishbone_bd_ram_mem0_reg[79][7]/P0001 ,
		_w11949_,
		_w11973_,
		_w20842_
	);
	LUT3 #(
		.INIT('h80)
	) name10330 (
		\wishbone_bd_ram_mem0_reg[189][7]/P0001 ,
		_w11942_,
		_w11966_,
		_w20843_
	);
	LUT4 #(
		.INIT('h0001)
	) name10331 (
		_w20840_,
		_w20841_,
		_w20842_,
		_w20843_,
		_w20844_
	);
	LUT3 #(
		.INIT('h80)
	) name10332 (
		\wishbone_bd_ram_mem0_reg[91][7]/P0001 ,
		_w11936_,
		_w11972_,
		_w20845_
	);
	LUT3 #(
		.INIT('h80)
	) name10333 (
		\wishbone_bd_ram_mem0_reg[72][7]/P0001 ,
		_w11949_,
		_w11990_,
		_w20846_
	);
	LUT3 #(
		.INIT('h80)
	) name10334 (
		\wishbone_bd_ram_mem0_reg[149][7]/P0001 ,
		_w11933_,
		_w11959_,
		_w20847_
	);
	LUT3 #(
		.INIT('h80)
	) name10335 (
		\wishbone_bd_ram_mem0_reg[24][7]/P0001 ,
		_w11935_,
		_w11990_,
		_w20848_
	);
	LUT4 #(
		.INIT('h0001)
	) name10336 (
		_w20845_,
		_w20846_,
		_w20847_,
		_w20848_,
		_w20849_
	);
	LUT3 #(
		.INIT('h80)
	) name10337 (
		\wishbone_bd_ram_mem0_reg[22][7]/P0001 ,
		_w11935_,
		_w11986_,
		_w20850_
	);
	LUT3 #(
		.INIT('h80)
	) name10338 (
		\wishbone_bd_ram_mem0_reg[34][7]/P0001 ,
		_w11957_,
		_w11963_,
		_w20851_
	);
	LUT3 #(
		.INIT('h80)
	) name10339 (
		\wishbone_bd_ram_mem0_reg[136][7]/P0001 ,
		_w11955_,
		_w11990_,
		_w20852_
	);
	LUT3 #(
		.INIT('h80)
	) name10340 (
		\wishbone_bd_ram_mem0_reg[39][7]/P0001 ,
		_w11957_,
		_w11975_,
		_w20853_
	);
	LUT4 #(
		.INIT('h0001)
	) name10341 (
		_w20850_,
		_w20851_,
		_w20852_,
		_w20853_,
		_w20854_
	);
	LUT3 #(
		.INIT('h80)
	) name10342 (
		\wishbone_bd_ram_mem0_reg[172][7]/P0001 ,
		_w11930_,
		_w11954_,
		_w20855_
	);
	LUT3 #(
		.INIT('h80)
	) name10343 (
		\wishbone_bd_ram_mem0_reg[55][7]/P0001 ,
		_w11975_,
		_w11979_,
		_w20856_
	);
	LUT3 #(
		.INIT('h80)
	) name10344 (
		\wishbone_bd_ram_mem0_reg[95][7]/P0001 ,
		_w11972_,
		_w11973_,
		_w20857_
	);
	LUT3 #(
		.INIT('h80)
	) name10345 (
		\wishbone_bd_ram_mem0_reg[180][7]/P0001 ,
		_w11929_,
		_w11942_,
		_w20858_
	);
	LUT4 #(
		.INIT('h0001)
	) name10346 (
		_w20855_,
		_w20856_,
		_w20857_,
		_w20858_,
		_w20859_
	);
	LUT4 #(
		.INIT('h8000)
	) name10347 (
		_w20844_,
		_w20849_,
		_w20854_,
		_w20859_,
		_w20860_
	);
	LUT4 #(
		.INIT('h8000)
	) name10348 (
		_w20797_,
		_w20818_,
		_w20839_,
		_w20860_,
		_w20861_
	);
	LUT3 #(
		.INIT('h80)
	) name10349 (
		\wishbone_bd_ram_mem0_reg[61][7]/P0001 ,
		_w11966_,
		_w11979_,
		_w20862_
	);
	LUT3 #(
		.INIT('h80)
	) name10350 (
		\wishbone_bd_ram_mem0_reg[124][7]/P0001 ,
		_w11954_,
		_w12012_,
		_w20863_
	);
	LUT3 #(
		.INIT('h80)
	) name10351 (
		\wishbone_bd_ram_mem0_reg[247][7]/P0001 ,
		_w11952_,
		_w11975_,
		_w20864_
	);
	LUT3 #(
		.INIT('h80)
	) name10352 (
		\wishbone_bd_ram_mem0_reg[212][7]/P0001 ,
		_w11929_,
		_w11984_,
		_w20865_
	);
	LUT4 #(
		.INIT('h0001)
	) name10353 (
		_w20862_,
		_w20863_,
		_w20864_,
		_w20865_,
		_w20866_
	);
	LUT3 #(
		.INIT('h80)
	) name10354 (
		\wishbone_bd_ram_mem0_reg[255][7]/P0001 ,
		_w11952_,
		_w11973_,
		_w20867_
	);
	LUT3 #(
		.INIT('h80)
	) name10355 (
		\wishbone_bd_ram_mem0_reg[237][7]/P0001 ,
		_w11966_,
		_w11982_,
		_w20868_
	);
	LUT3 #(
		.INIT('h80)
	) name10356 (
		\wishbone_bd_ram_mem0_reg[128][7]/P0001 ,
		_w11941_,
		_w11955_,
		_w20869_
	);
	LUT3 #(
		.INIT('h80)
	) name10357 (
		\wishbone_bd_ram_mem0_reg[5][7]/P0001 ,
		_w11932_,
		_w11933_,
		_w20870_
	);
	LUT4 #(
		.INIT('h0001)
	) name10358 (
		_w20867_,
		_w20868_,
		_w20869_,
		_w20870_,
		_w20871_
	);
	LUT3 #(
		.INIT('h80)
	) name10359 (
		\wishbone_bd_ram_mem0_reg[196][7]/P0001 ,
		_w11929_,
		_w11945_,
		_w20872_
	);
	LUT3 #(
		.INIT('h80)
	) name10360 (
		\wishbone_bd_ram_mem0_reg[82][7]/P0001 ,
		_w11963_,
		_w11972_,
		_w20873_
	);
	LUT3 #(
		.INIT('h80)
	) name10361 (
		\wishbone_bd_ram_mem0_reg[253][7]/P0001 ,
		_w11952_,
		_w11966_,
		_w20874_
	);
	LUT3 #(
		.INIT('h80)
	) name10362 (
		\wishbone_bd_ram_mem0_reg[211][7]/P0001 ,
		_w11938_,
		_w11984_,
		_w20875_
	);
	LUT4 #(
		.INIT('h0001)
	) name10363 (
		_w20872_,
		_w20873_,
		_w20874_,
		_w20875_,
		_w20876_
	);
	LUT3 #(
		.INIT('h80)
	) name10364 (
		\wishbone_bd_ram_mem0_reg[70][7]/P0001 ,
		_w11949_,
		_w11986_,
		_w20877_
	);
	LUT3 #(
		.INIT('h80)
	) name10365 (
		\wishbone_bd_ram_mem0_reg[141][7]/P0001 ,
		_w11955_,
		_w11966_,
		_w20878_
	);
	LUT3 #(
		.INIT('h80)
	) name10366 (
		\wishbone_bd_ram_mem0_reg[108][7]/P0001 ,
		_w11954_,
		_w11965_,
		_w20879_
	);
	LUT3 #(
		.INIT('h80)
	) name10367 (
		\wishbone_bd_ram_mem0_reg[186][7]/P0001 ,
		_w11942_,
		_w11944_,
		_w20880_
	);
	LUT4 #(
		.INIT('h0001)
	) name10368 (
		_w20877_,
		_w20878_,
		_w20879_,
		_w20880_,
		_w20881_
	);
	LUT4 #(
		.INIT('h8000)
	) name10369 (
		_w20866_,
		_w20871_,
		_w20876_,
		_w20881_,
		_w20882_
	);
	LUT3 #(
		.INIT('h80)
	) name10370 (
		\wishbone_bd_ram_mem0_reg[57][7]/P0001 ,
		_w11968_,
		_w11979_,
		_w20883_
	);
	LUT3 #(
		.INIT('h80)
	) name10371 (
		\wishbone_bd_ram_mem0_reg[179][7]/P0001 ,
		_w11938_,
		_w11942_,
		_w20884_
	);
	LUT3 #(
		.INIT('h80)
	) name10372 (
		\wishbone_bd_ram_mem0_reg[42][7]/P0001 ,
		_w11944_,
		_w11957_,
		_w20885_
	);
	LUT3 #(
		.INIT('h80)
	) name10373 (
		\wishbone_bd_ram_mem0_reg[31][7]/P0001 ,
		_w11935_,
		_w11973_,
		_w20886_
	);
	LUT4 #(
		.INIT('h0001)
	) name10374 (
		_w20883_,
		_w20884_,
		_w20885_,
		_w20886_,
		_w20887_
	);
	LUT3 #(
		.INIT('h80)
	) name10375 (
		\wishbone_bd_ram_mem0_reg[8][7]/P0001 ,
		_w11932_,
		_w11990_,
		_w20888_
	);
	LUT3 #(
		.INIT('h80)
	) name10376 (
		\wishbone_bd_ram_mem0_reg[80][7]/P0001 ,
		_w11941_,
		_w11972_,
		_w20889_
	);
	LUT3 #(
		.INIT('h80)
	) name10377 (
		\wishbone_bd_ram_mem0_reg[230][7]/P0001 ,
		_w11982_,
		_w11986_,
		_w20890_
	);
	LUT3 #(
		.INIT('h80)
	) name10378 (
		\wishbone_bd_ram_mem0_reg[64][7]/P0001 ,
		_w11941_,
		_w11949_,
		_w20891_
	);
	LUT4 #(
		.INIT('h0001)
	) name10379 (
		_w20888_,
		_w20889_,
		_w20890_,
		_w20891_,
		_w20892_
	);
	LUT3 #(
		.INIT('h80)
	) name10380 (
		\wishbone_bd_ram_mem0_reg[16][7]/P0001 ,
		_w11935_,
		_w11941_,
		_w20893_
	);
	LUT3 #(
		.INIT('h80)
	) name10381 (
		\wishbone_bd_ram_mem0_reg[219][7]/P0001 ,
		_w11936_,
		_w11984_,
		_w20894_
	);
	LUT3 #(
		.INIT('h80)
	) name10382 (
		\wishbone_bd_ram_mem0_reg[38][7]/P0001 ,
		_w11957_,
		_w11986_,
		_w20895_
	);
	LUT3 #(
		.INIT('h80)
	) name10383 (
		\wishbone_bd_ram_mem0_reg[23][7]/P0001 ,
		_w11935_,
		_w11975_,
		_w20896_
	);
	LUT4 #(
		.INIT('h0001)
	) name10384 (
		_w20893_,
		_w20894_,
		_w20895_,
		_w20896_,
		_w20897_
	);
	LUT3 #(
		.INIT('h80)
	) name10385 (
		\wishbone_bd_ram_mem0_reg[107][7]/P0001 ,
		_w11936_,
		_w11965_,
		_w20898_
	);
	LUT3 #(
		.INIT('h80)
	) name10386 (
		\wishbone_bd_ram_mem0_reg[246][7]/P0001 ,
		_w11952_,
		_w11986_,
		_w20899_
	);
	LUT3 #(
		.INIT('h80)
	) name10387 (
		\wishbone_bd_ram_mem0_reg[77][7]/P0001 ,
		_w11949_,
		_w11966_,
		_w20900_
	);
	LUT3 #(
		.INIT('h80)
	) name10388 (
		\wishbone_bd_ram_mem0_reg[109][7]/P0001 ,
		_w11965_,
		_w11966_,
		_w20901_
	);
	LUT4 #(
		.INIT('h0001)
	) name10389 (
		_w20898_,
		_w20899_,
		_w20900_,
		_w20901_,
		_w20902_
	);
	LUT4 #(
		.INIT('h8000)
	) name10390 (
		_w20887_,
		_w20892_,
		_w20897_,
		_w20902_,
		_w20903_
	);
	LUT3 #(
		.INIT('h80)
	) name10391 (
		\wishbone_bd_ram_mem0_reg[7][7]/P0001 ,
		_w11932_,
		_w11975_,
		_w20904_
	);
	LUT3 #(
		.INIT('h80)
	) name10392 (
		\wishbone_bd_ram_mem0_reg[158][7]/P0001 ,
		_w11948_,
		_w11959_,
		_w20905_
	);
	LUT3 #(
		.INIT('h80)
	) name10393 (
		\wishbone_bd_ram_mem0_reg[102][7]/P0001 ,
		_w11965_,
		_w11986_,
		_w20906_
	);
	LUT3 #(
		.INIT('h80)
	) name10394 (
		\wishbone_bd_ram_mem0_reg[114][7]/P0001 ,
		_w11963_,
		_w12012_,
		_w20907_
	);
	LUT4 #(
		.INIT('h0001)
	) name10395 (
		_w20904_,
		_w20905_,
		_w20906_,
		_w20907_,
		_w20908_
	);
	LUT3 #(
		.INIT('h80)
	) name10396 (
		\wishbone_bd_ram_mem0_reg[191][7]/P0001 ,
		_w11942_,
		_w11973_,
		_w20909_
	);
	LUT3 #(
		.INIT('h80)
	) name10397 (
		\wishbone_bd_ram_mem0_reg[92][7]/P0001 ,
		_w11954_,
		_w11972_,
		_w20910_
	);
	LUT3 #(
		.INIT('h80)
	) name10398 (
		\wishbone_bd_ram_mem0_reg[30][7]/P0001 ,
		_w11935_,
		_w11948_,
		_w20911_
	);
	LUT3 #(
		.INIT('h80)
	) name10399 (
		\wishbone_bd_ram_mem0_reg[26][7]/P0001 ,
		_w11935_,
		_w11944_,
		_w20912_
	);
	LUT4 #(
		.INIT('h0001)
	) name10400 (
		_w20909_,
		_w20910_,
		_w20911_,
		_w20912_,
		_w20913_
	);
	LUT3 #(
		.INIT('h80)
	) name10401 (
		\wishbone_bd_ram_mem0_reg[221][7]/P0001 ,
		_w11966_,
		_w11984_,
		_w20914_
	);
	LUT3 #(
		.INIT('h80)
	) name10402 (
		\wishbone_bd_ram_mem0_reg[131][7]/P0001 ,
		_w11938_,
		_w11955_,
		_w20915_
	);
	LUT3 #(
		.INIT('h80)
	) name10403 (
		\wishbone_bd_ram_mem0_reg[210][7]/P0001 ,
		_w11963_,
		_w11984_,
		_w20916_
	);
	LUT3 #(
		.INIT('h80)
	) name10404 (
		\wishbone_bd_ram_mem0_reg[223][7]/P0001 ,
		_w11973_,
		_w11984_,
		_w20917_
	);
	LUT4 #(
		.INIT('h0001)
	) name10405 (
		_w20914_,
		_w20915_,
		_w20916_,
		_w20917_,
		_w20918_
	);
	LUT3 #(
		.INIT('h80)
	) name10406 (
		\wishbone_bd_ram_mem0_reg[151][7]/P0001 ,
		_w11959_,
		_w11975_,
		_w20919_
	);
	LUT3 #(
		.INIT('h80)
	) name10407 (
		\wishbone_bd_ram_mem0_reg[227][7]/P0001 ,
		_w11938_,
		_w11982_,
		_w20920_
	);
	LUT3 #(
		.INIT('h80)
	) name10408 (
		\wishbone_bd_ram_mem0_reg[122][7]/P0001 ,
		_w11944_,
		_w12012_,
		_w20921_
	);
	LUT3 #(
		.INIT('h80)
	) name10409 (
		\wishbone_bd_ram_mem0_reg[117][7]/P0001 ,
		_w11933_,
		_w12012_,
		_w20922_
	);
	LUT4 #(
		.INIT('h0001)
	) name10410 (
		_w20919_,
		_w20920_,
		_w20921_,
		_w20922_,
		_w20923_
	);
	LUT4 #(
		.INIT('h8000)
	) name10411 (
		_w20908_,
		_w20913_,
		_w20918_,
		_w20923_,
		_w20924_
	);
	LUT3 #(
		.INIT('h80)
	) name10412 (
		\wishbone_bd_ram_mem0_reg[3][7]/P0001 ,
		_w11932_,
		_w11938_,
		_w20925_
	);
	LUT3 #(
		.INIT('h80)
	) name10413 (
		\wishbone_bd_ram_mem0_reg[10][7]/P0001 ,
		_w11932_,
		_w11944_,
		_w20926_
	);
	LUT3 #(
		.INIT('h80)
	) name10414 (
		\wishbone_bd_ram_mem0_reg[198][7]/P0001 ,
		_w11945_,
		_w11986_,
		_w20927_
	);
	LUT3 #(
		.INIT('h80)
	) name10415 (
		\wishbone_bd_ram_mem0_reg[232][7]/P0001 ,
		_w11982_,
		_w11990_,
		_w20928_
	);
	LUT4 #(
		.INIT('h0001)
	) name10416 (
		_w20925_,
		_w20926_,
		_w20927_,
		_w20928_,
		_w20929_
	);
	LUT3 #(
		.INIT('h80)
	) name10417 (
		\wishbone_bd_ram_mem0_reg[150][7]/P0001 ,
		_w11959_,
		_w11986_,
		_w20930_
	);
	LUT3 #(
		.INIT('h80)
	) name10418 (
		\wishbone_bd_ram_mem0_reg[245][7]/P0001 ,
		_w11933_,
		_w11952_,
		_w20931_
	);
	LUT3 #(
		.INIT('h80)
	) name10419 (
		\wishbone_bd_ram_mem0_reg[74][7]/P0001 ,
		_w11944_,
		_w11949_,
		_w20932_
	);
	LUT3 #(
		.INIT('h80)
	) name10420 (
		\wishbone_bd_ram_mem0_reg[138][7]/P0001 ,
		_w11944_,
		_w11955_,
		_w20933_
	);
	LUT4 #(
		.INIT('h0001)
	) name10421 (
		_w20930_,
		_w20931_,
		_w20932_,
		_w20933_,
		_w20934_
	);
	LUT3 #(
		.INIT('h80)
	) name10422 (
		\wishbone_bd_ram_mem0_reg[224][7]/P0001 ,
		_w11941_,
		_w11982_,
		_w20935_
	);
	LUT3 #(
		.INIT('h80)
	) name10423 (
		\wishbone_bd_ram_mem0_reg[152][7]/P0001 ,
		_w11959_,
		_w11990_,
		_w20936_
	);
	LUT3 #(
		.INIT('h80)
	) name10424 (
		\wishbone_bd_ram_mem0_reg[35][7]/P0001 ,
		_w11938_,
		_w11957_,
		_w20937_
	);
	LUT3 #(
		.INIT('h80)
	) name10425 (
		\wishbone_bd_ram_mem0_reg[238][7]/P0001 ,
		_w11948_,
		_w11982_,
		_w20938_
	);
	LUT4 #(
		.INIT('h0001)
	) name10426 (
		_w20935_,
		_w20936_,
		_w20937_,
		_w20938_,
		_w20939_
	);
	LUT3 #(
		.INIT('h80)
	) name10427 (
		\wishbone_bd_ram_mem0_reg[120][7]/P0001 ,
		_w11990_,
		_w12012_,
		_w20940_
	);
	LUT3 #(
		.INIT('h80)
	) name10428 (
		\wishbone_bd_ram_mem0_reg[206][7]/P0001 ,
		_w11945_,
		_w11948_,
		_w20941_
	);
	LUT3 #(
		.INIT('h80)
	) name10429 (
		\wishbone_bd_ram_mem0_reg[13][7]/P0001 ,
		_w11932_,
		_w11966_,
		_w20942_
	);
	LUT3 #(
		.INIT('h80)
	) name10430 (
		\wishbone_bd_ram_mem0_reg[119][7]/P0001 ,
		_w11975_,
		_w12012_,
		_w20943_
	);
	LUT4 #(
		.INIT('h0001)
	) name10431 (
		_w20940_,
		_w20941_,
		_w20942_,
		_w20943_,
		_w20944_
	);
	LUT4 #(
		.INIT('h8000)
	) name10432 (
		_w20929_,
		_w20934_,
		_w20939_,
		_w20944_,
		_w20945_
	);
	LUT4 #(
		.INIT('h8000)
	) name10433 (
		_w20882_,
		_w20903_,
		_w20924_,
		_w20945_,
		_w20946_
	);
	LUT3 #(
		.INIT('h80)
	) name10434 (
		\wishbone_bd_ram_mem0_reg[29][7]/P0001 ,
		_w11935_,
		_w11966_,
		_w20947_
	);
	LUT3 #(
		.INIT('h80)
	) name10435 (
		\wishbone_bd_ram_mem0_reg[0][7]/P0001 ,
		_w11932_,
		_w11941_,
		_w20948_
	);
	LUT3 #(
		.INIT('h80)
	) name10436 (
		\wishbone_bd_ram_mem0_reg[99][7]/P0001 ,
		_w11938_,
		_w11965_,
		_w20949_
	);
	LUT3 #(
		.INIT('h80)
	) name10437 (
		\wishbone_bd_ram_mem0_reg[239][7]/P0001 ,
		_w11973_,
		_w11982_,
		_w20950_
	);
	LUT4 #(
		.INIT('h0001)
	) name10438 (
		_w20947_,
		_w20948_,
		_w20949_,
		_w20950_,
		_w20951_
	);
	LUT3 #(
		.INIT('h80)
	) name10439 (
		\wishbone_bd_ram_mem0_reg[160][7]/P0001 ,
		_w11930_,
		_w11941_,
		_w20952_
	);
	LUT3 #(
		.INIT('h80)
	) name10440 (
		\wishbone_bd_ram_mem0_reg[2][7]/P0001 ,
		_w11932_,
		_w11963_,
		_w20953_
	);
	LUT3 #(
		.INIT('h80)
	) name10441 (
		\wishbone_bd_ram_mem0_reg[254][7]/P0001 ,
		_w11948_,
		_w11952_,
		_w20954_
	);
	LUT3 #(
		.INIT('h80)
	) name10442 (
		\wishbone_bd_ram_mem0_reg[155][7]/P0001 ,
		_w11936_,
		_w11959_,
		_w20955_
	);
	LUT4 #(
		.INIT('h0001)
	) name10443 (
		_w20952_,
		_w20953_,
		_w20954_,
		_w20955_,
		_w20956_
	);
	LUT3 #(
		.INIT('h80)
	) name10444 (
		\wishbone_bd_ram_mem0_reg[217][7]/P0001 ,
		_w11968_,
		_w11984_,
		_w20957_
	);
	LUT3 #(
		.INIT('h80)
	) name10445 (
		\wishbone_bd_ram_mem0_reg[1][7]/P0001 ,
		_w11932_,
		_w11977_,
		_w20958_
	);
	LUT3 #(
		.INIT('h80)
	) name10446 (
		\wishbone_bd_ram_mem0_reg[84][7]/P0001 ,
		_w11929_,
		_w11972_,
		_w20959_
	);
	LUT3 #(
		.INIT('h80)
	) name10447 (
		\wishbone_bd_ram_mem0_reg[214][7]/P0001 ,
		_w11984_,
		_w11986_,
		_w20960_
	);
	LUT4 #(
		.INIT('h0001)
	) name10448 (
		_w20957_,
		_w20958_,
		_w20959_,
		_w20960_,
		_w20961_
	);
	LUT3 #(
		.INIT('h80)
	) name10449 (
		\wishbone_bd_ram_mem0_reg[62][7]/P0001 ,
		_w11948_,
		_w11979_,
		_w20962_
	);
	LUT3 #(
		.INIT('h80)
	) name10450 (
		\wishbone_bd_ram_mem0_reg[182][7]/P0001 ,
		_w11942_,
		_w11986_,
		_w20963_
	);
	LUT3 #(
		.INIT('h80)
	) name10451 (
		\wishbone_bd_ram_mem0_reg[94][7]/P0001 ,
		_w11948_,
		_w11972_,
		_w20964_
	);
	LUT3 #(
		.INIT('h80)
	) name10452 (
		\wishbone_bd_ram_mem0_reg[41][7]/P0001 ,
		_w11957_,
		_w11968_,
		_w20965_
	);
	LUT4 #(
		.INIT('h0001)
	) name10453 (
		_w20962_,
		_w20963_,
		_w20964_,
		_w20965_,
		_w20966_
	);
	LUT4 #(
		.INIT('h8000)
	) name10454 (
		_w20951_,
		_w20956_,
		_w20961_,
		_w20966_,
		_w20967_
	);
	LUT3 #(
		.INIT('h80)
	) name10455 (
		\wishbone_bd_ram_mem0_reg[201][7]/P0001 ,
		_w11945_,
		_w11968_,
		_w20968_
	);
	LUT3 #(
		.INIT('h80)
	) name10456 (
		\wishbone_bd_ram_mem0_reg[33][7]/P0001 ,
		_w11957_,
		_w11977_,
		_w20969_
	);
	LUT3 #(
		.INIT('h80)
	) name10457 (
		\wishbone_bd_ram_mem0_reg[52][7]/P0001 ,
		_w11929_,
		_w11979_,
		_w20970_
	);
	LUT3 #(
		.INIT('h80)
	) name10458 (
		\wishbone_bd_ram_mem0_reg[78][7]/P0001 ,
		_w11948_,
		_w11949_,
		_w20971_
	);
	LUT4 #(
		.INIT('h0001)
	) name10459 (
		_w20968_,
		_w20969_,
		_w20970_,
		_w20971_,
		_w20972_
	);
	LUT3 #(
		.INIT('h80)
	) name10460 (
		\wishbone_bd_ram_mem0_reg[226][7]/P0001 ,
		_w11963_,
		_w11982_,
		_w20973_
	);
	LUT3 #(
		.INIT('h80)
	) name10461 (
		\wishbone_bd_ram_mem0_reg[215][7]/P0001 ,
		_w11975_,
		_w11984_,
		_w20974_
	);
	LUT3 #(
		.INIT('h80)
	) name10462 (
		\wishbone_bd_ram_mem0_reg[184][7]/P0001 ,
		_w11942_,
		_w11990_,
		_w20975_
	);
	LUT3 #(
		.INIT('h80)
	) name10463 (
		\wishbone_bd_ram_mem0_reg[83][7]/P0001 ,
		_w11938_,
		_w11972_,
		_w20976_
	);
	LUT4 #(
		.INIT('h0001)
	) name10464 (
		_w20973_,
		_w20974_,
		_w20975_,
		_w20976_,
		_w20977_
	);
	LUT3 #(
		.INIT('h80)
	) name10465 (
		\wishbone_bd_ram_mem0_reg[171][7]/P0001 ,
		_w11930_,
		_w11936_,
		_w20978_
	);
	LUT3 #(
		.INIT('h80)
	) name10466 (
		\wishbone_bd_ram_mem0_reg[65][7]/P0001 ,
		_w11949_,
		_w11977_,
		_w20979_
	);
	LUT3 #(
		.INIT('h80)
	) name10467 (
		\wishbone_bd_ram_mem0_reg[14][7]/P0001 ,
		_w11932_,
		_w11948_,
		_w20980_
	);
	LUT3 #(
		.INIT('h80)
	) name10468 (
		\wishbone_bd_ram_mem0_reg[25][7]/P0001 ,
		_w11935_,
		_w11968_,
		_w20981_
	);
	LUT4 #(
		.INIT('h0001)
	) name10469 (
		_w20978_,
		_w20979_,
		_w20980_,
		_w20981_,
		_w20982_
	);
	LUT3 #(
		.INIT('h80)
	) name10470 (
		\wishbone_bd_ram_mem0_reg[66][7]/P0001 ,
		_w11949_,
		_w11963_,
		_w20983_
	);
	LUT3 #(
		.INIT('h80)
	) name10471 (
		\wishbone_bd_ram_mem0_reg[46][7]/P0001 ,
		_w11948_,
		_w11957_,
		_w20984_
	);
	LUT3 #(
		.INIT('h80)
	) name10472 (
		\wishbone_bd_ram_mem0_reg[159][7]/P0001 ,
		_w11959_,
		_w11973_,
		_w20985_
	);
	LUT3 #(
		.INIT('h80)
	) name10473 (
		\wishbone_bd_ram_mem0_reg[89][7]/P0001 ,
		_w11968_,
		_w11972_,
		_w20986_
	);
	LUT4 #(
		.INIT('h0001)
	) name10474 (
		_w20983_,
		_w20984_,
		_w20985_,
		_w20986_,
		_w20987_
	);
	LUT4 #(
		.INIT('h8000)
	) name10475 (
		_w20972_,
		_w20977_,
		_w20982_,
		_w20987_,
		_w20988_
	);
	LUT3 #(
		.INIT('h80)
	) name10476 (
		\wishbone_bd_ram_mem0_reg[250][7]/P0001 ,
		_w11944_,
		_w11952_,
		_w20989_
	);
	LUT3 #(
		.INIT('h80)
	) name10477 (
		\wishbone_bd_ram_mem0_reg[51][7]/P0001 ,
		_w11938_,
		_w11979_,
		_w20990_
	);
	LUT3 #(
		.INIT('h80)
	) name10478 (
		\wishbone_bd_ram_mem0_reg[209][7]/P0001 ,
		_w11977_,
		_w11984_,
		_w20991_
	);
	LUT3 #(
		.INIT('h80)
	) name10479 (
		\wishbone_bd_ram_mem0_reg[127][7]/P0001 ,
		_w11973_,
		_w12012_,
		_w20992_
	);
	LUT4 #(
		.INIT('h0001)
	) name10480 (
		_w20989_,
		_w20990_,
		_w20991_,
		_w20992_,
		_w20993_
	);
	LUT3 #(
		.INIT('h80)
	) name10481 (
		\wishbone_bd_ram_mem0_reg[87][7]/P0001 ,
		_w11972_,
		_w11975_,
		_w20994_
	);
	LUT3 #(
		.INIT('h80)
	) name10482 (
		\wishbone_bd_ram_mem0_reg[103][7]/P0001 ,
		_w11965_,
		_w11975_,
		_w20995_
	);
	LUT3 #(
		.INIT('h80)
	) name10483 (
		\wishbone_bd_ram_mem0_reg[234][7]/P0001 ,
		_w11944_,
		_w11982_,
		_w20996_
	);
	LUT3 #(
		.INIT('h80)
	) name10484 (
		\wishbone_bd_ram_mem0_reg[81][7]/P0001 ,
		_w11972_,
		_w11977_,
		_w20997_
	);
	LUT4 #(
		.INIT('h0001)
	) name10485 (
		_w20994_,
		_w20995_,
		_w20996_,
		_w20997_,
		_w20998_
	);
	LUT3 #(
		.INIT('h80)
	) name10486 (
		\wishbone_bd_ram_mem0_reg[88][7]/P0001 ,
		_w11972_,
		_w11990_,
		_w20999_
	);
	LUT3 #(
		.INIT('h80)
	) name10487 (
		\wishbone_bd_ram_mem0_reg[133][7]/P0001 ,
		_w11933_,
		_w11955_,
		_w21000_
	);
	LUT3 #(
		.INIT('h80)
	) name10488 (
		\wishbone_bd_ram_mem0_reg[20][7]/P0001 ,
		_w11929_,
		_w11935_,
		_w21001_
	);
	LUT3 #(
		.INIT('h80)
	) name10489 (
		\wishbone_bd_ram_mem0_reg[204][7]/P0001 ,
		_w11945_,
		_w11954_,
		_w21002_
	);
	LUT4 #(
		.INIT('h0001)
	) name10490 (
		_w20999_,
		_w21000_,
		_w21001_,
		_w21002_,
		_w21003_
	);
	LUT3 #(
		.INIT('h80)
	) name10491 (
		\wishbone_bd_ram_mem0_reg[140][7]/P0001 ,
		_w11954_,
		_w11955_,
		_w21004_
	);
	LUT3 #(
		.INIT('h80)
	) name10492 (
		\wishbone_bd_ram_mem0_reg[137][7]/P0001 ,
		_w11955_,
		_w11968_,
		_w21005_
	);
	LUT3 #(
		.INIT('h80)
	) name10493 (
		\wishbone_bd_ram_mem0_reg[123][7]/P0001 ,
		_w11936_,
		_w12012_,
		_w21006_
	);
	LUT3 #(
		.INIT('h80)
	) name10494 (
		\wishbone_bd_ram_mem0_reg[76][7]/P0001 ,
		_w11949_,
		_w11954_,
		_w21007_
	);
	LUT4 #(
		.INIT('h0001)
	) name10495 (
		_w21004_,
		_w21005_,
		_w21006_,
		_w21007_,
		_w21008_
	);
	LUT4 #(
		.INIT('h8000)
	) name10496 (
		_w20993_,
		_w20998_,
		_w21003_,
		_w21008_,
		_w21009_
	);
	LUT3 #(
		.INIT('h80)
	) name10497 (
		\wishbone_bd_ram_mem0_reg[126][7]/P0001 ,
		_w11948_,
		_w12012_,
		_w21010_
	);
	LUT3 #(
		.INIT('h80)
	) name10498 (
		\wishbone_bd_ram_mem0_reg[174][7]/P0001 ,
		_w11930_,
		_w11948_,
		_w21011_
	);
	LUT3 #(
		.INIT('h80)
	) name10499 (
		\wishbone_bd_ram_mem0_reg[63][7]/P0001 ,
		_w11973_,
		_w11979_,
		_w21012_
	);
	LUT3 #(
		.INIT('h80)
	) name10500 (
		\wishbone_bd_ram_mem0_reg[115][7]/P0001 ,
		_w11938_,
		_w12012_,
		_w21013_
	);
	LUT4 #(
		.INIT('h0001)
	) name10501 (
		_w21010_,
		_w21011_,
		_w21012_,
		_w21013_,
		_w21014_
	);
	LUT3 #(
		.INIT('h80)
	) name10502 (
		\wishbone_bd_ram_mem0_reg[231][7]/P0001 ,
		_w11975_,
		_w11982_,
		_w21015_
	);
	LUT3 #(
		.INIT('h80)
	) name10503 (
		\wishbone_bd_ram_mem0_reg[205][7]/P0001 ,
		_w11945_,
		_w11966_,
		_w21016_
	);
	LUT3 #(
		.INIT('h80)
	) name10504 (
		\wishbone_bd_ram_mem0_reg[187][7]/P0001 ,
		_w11936_,
		_w11942_,
		_w21017_
	);
	LUT3 #(
		.INIT('h80)
	) name10505 (
		\wishbone_bd_ram_mem0_reg[113][7]/P0001 ,
		_w11977_,
		_w12012_,
		_w21018_
	);
	LUT4 #(
		.INIT('h0001)
	) name10506 (
		_w21015_,
		_w21016_,
		_w21017_,
		_w21018_,
		_w21019_
	);
	LUT3 #(
		.INIT('h80)
	) name10507 (
		\wishbone_bd_ram_mem0_reg[139][7]/P0001 ,
		_w11936_,
		_w11955_,
		_w21020_
	);
	LUT3 #(
		.INIT('h80)
	) name10508 (
		\wishbone_bd_ram_mem0_reg[157][7]/P0001 ,
		_w11959_,
		_w11966_,
		_w21021_
	);
	LUT3 #(
		.INIT('h80)
	) name10509 (
		\wishbone_bd_ram_mem0_reg[15][7]/P0001 ,
		_w11932_,
		_w11973_,
		_w21022_
	);
	LUT3 #(
		.INIT('h80)
	) name10510 (
		\wishbone_bd_ram_mem0_reg[132][7]/P0001 ,
		_w11929_,
		_w11955_,
		_w21023_
	);
	LUT4 #(
		.INIT('h0001)
	) name10511 (
		_w21020_,
		_w21021_,
		_w21022_,
		_w21023_,
		_w21024_
	);
	LUT3 #(
		.INIT('h80)
	) name10512 (
		\wishbone_bd_ram_mem0_reg[147][7]/P0001 ,
		_w11938_,
		_w11959_,
		_w21025_
	);
	LUT3 #(
		.INIT('h80)
	) name10513 (
		\wishbone_bd_ram_mem0_reg[75][7]/P0001 ,
		_w11936_,
		_w11949_,
		_w21026_
	);
	LUT3 #(
		.INIT('h80)
	) name10514 (
		\wishbone_bd_ram_mem0_reg[18][7]/P0001 ,
		_w11935_,
		_w11963_,
		_w21027_
	);
	LUT3 #(
		.INIT('h80)
	) name10515 (
		\wishbone_bd_ram_mem0_reg[40][7]/P0001 ,
		_w11957_,
		_w11990_,
		_w21028_
	);
	LUT4 #(
		.INIT('h0001)
	) name10516 (
		_w21025_,
		_w21026_,
		_w21027_,
		_w21028_,
		_w21029_
	);
	LUT4 #(
		.INIT('h8000)
	) name10517 (
		_w21014_,
		_w21019_,
		_w21024_,
		_w21029_,
		_w21030_
	);
	LUT4 #(
		.INIT('h8000)
	) name10518 (
		_w20967_,
		_w20988_,
		_w21009_,
		_w21030_,
		_w21031_
	);
	LUT3 #(
		.INIT('h80)
	) name10519 (
		\wishbone_bd_ram_mem0_reg[135][7]/P0001 ,
		_w11955_,
		_w11975_,
		_w21032_
	);
	LUT3 #(
		.INIT('h80)
	) name10520 (
		\wishbone_bd_ram_mem0_reg[111][7]/P0001 ,
		_w11965_,
		_w11973_,
		_w21033_
	);
	LUT3 #(
		.INIT('h80)
	) name10521 (
		\wishbone_bd_ram_mem0_reg[134][7]/P0001 ,
		_w11955_,
		_w11986_,
		_w21034_
	);
	LUT3 #(
		.INIT('h80)
	) name10522 (
		\wishbone_bd_ram_mem0_reg[165][7]/P0001 ,
		_w11930_,
		_w11933_,
		_w21035_
	);
	LUT4 #(
		.INIT('h0001)
	) name10523 (
		_w21032_,
		_w21033_,
		_w21034_,
		_w21035_,
		_w21036_
	);
	LUT3 #(
		.INIT('h80)
	) name10524 (
		\wishbone_bd_ram_mem0_reg[90][7]/P0001 ,
		_w11944_,
		_w11972_,
		_w21037_
	);
	LUT3 #(
		.INIT('h80)
	) name10525 (
		\wishbone_bd_ram_mem0_reg[100][7]/P0001 ,
		_w11929_,
		_w11965_,
		_w21038_
	);
	LUT3 #(
		.INIT('h80)
	) name10526 (
		\wishbone_bd_ram_mem0_reg[47][7]/P0001 ,
		_w11957_,
		_w11973_,
		_w21039_
	);
	LUT3 #(
		.INIT('h80)
	) name10527 (
		\wishbone_bd_ram_mem0_reg[249][7]/P0001 ,
		_w11952_,
		_w11968_,
		_w21040_
	);
	LUT4 #(
		.INIT('h0001)
	) name10528 (
		_w21037_,
		_w21038_,
		_w21039_,
		_w21040_,
		_w21041_
	);
	LUT3 #(
		.INIT('h80)
	) name10529 (
		\wishbone_bd_ram_mem0_reg[162][7]/P0001 ,
		_w11930_,
		_w11963_,
		_w21042_
	);
	LUT3 #(
		.INIT('h80)
	) name10530 (
		\wishbone_bd_ram_mem0_reg[225][7]/P0001 ,
		_w11977_,
		_w11982_,
		_w21043_
	);
	LUT3 #(
		.INIT('h80)
	) name10531 (
		\wishbone_bd_ram_mem0_reg[6][7]/P0001 ,
		_w11932_,
		_w11986_,
		_w21044_
	);
	LUT3 #(
		.INIT('h80)
	) name10532 (
		\wishbone_bd_ram_mem0_reg[220][7]/P0001 ,
		_w11954_,
		_w11984_,
		_w21045_
	);
	LUT4 #(
		.INIT('h0001)
	) name10533 (
		_w21042_,
		_w21043_,
		_w21044_,
		_w21045_,
		_w21046_
	);
	LUT3 #(
		.INIT('h80)
	) name10534 (
		\wishbone_bd_ram_mem0_reg[73][7]/P0001 ,
		_w11949_,
		_w11968_,
		_w21047_
	);
	LUT3 #(
		.INIT('h80)
	) name10535 (
		\wishbone_bd_ram_mem0_reg[4][7]/P0001 ,
		_w11929_,
		_w11932_,
		_w21048_
	);
	LUT3 #(
		.INIT('h80)
	) name10536 (
		\wishbone_bd_ram_mem0_reg[129][7]/P0001 ,
		_w11955_,
		_w11977_,
		_w21049_
	);
	LUT3 #(
		.INIT('h80)
	) name10537 (
		\wishbone_bd_ram_mem0_reg[56][7]/P0001 ,
		_w11979_,
		_w11990_,
		_w21050_
	);
	LUT4 #(
		.INIT('h0001)
	) name10538 (
		_w21047_,
		_w21048_,
		_w21049_,
		_w21050_,
		_w21051_
	);
	LUT4 #(
		.INIT('h8000)
	) name10539 (
		_w21036_,
		_w21041_,
		_w21046_,
		_w21051_,
		_w21052_
	);
	LUT3 #(
		.INIT('h80)
	) name10540 (
		\wishbone_bd_ram_mem0_reg[145][7]/P0001 ,
		_w11959_,
		_w11977_,
		_w21053_
	);
	LUT3 #(
		.INIT('h80)
	) name10541 (
		\wishbone_bd_ram_mem0_reg[11][7]/P0001 ,
		_w11932_,
		_w11936_,
		_w21054_
	);
	LUT3 #(
		.INIT('h80)
	) name10542 (
		\wishbone_bd_ram_mem0_reg[148][7]/P0001 ,
		_w11929_,
		_w11959_,
		_w21055_
	);
	LUT3 #(
		.INIT('h80)
	) name10543 (
		\wishbone_bd_ram_mem0_reg[121][7]/P0001 ,
		_w11968_,
		_w12012_,
		_w21056_
	);
	LUT4 #(
		.INIT('h0001)
	) name10544 (
		_w21053_,
		_w21054_,
		_w21055_,
		_w21056_,
		_w21057_
	);
	LUT3 #(
		.INIT('h80)
	) name10545 (
		\wishbone_bd_ram_mem0_reg[125][7]/P0001 ,
		_w11966_,
		_w12012_,
		_w21058_
	);
	LUT3 #(
		.INIT('h80)
	) name10546 (
		\wishbone_bd_ram_mem0_reg[54][7]/P0001 ,
		_w11979_,
		_w11986_,
		_w21059_
	);
	LUT3 #(
		.INIT('h80)
	) name10547 (
		\wishbone_bd_ram_mem0_reg[32][7]/P0001 ,
		_w11941_,
		_w11957_,
		_w21060_
	);
	LUT3 #(
		.INIT('h80)
	) name10548 (
		\wishbone_bd_ram_mem0_reg[96][7]/P0001 ,
		_w11941_,
		_w11965_,
		_w21061_
	);
	LUT4 #(
		.INIT('h0001)
	) name10549 (
		_w21058_,
		_w21059_,
		_w21060_,
		_w21061_,
		_w21062_
	);
	LUT3 #(
		.INIT('h80)
	) name10550 (
		\wishbone_bd_ram_mem0_reg[185][7]/P0001 ,
		_w11942_,
		_w11968_,
		_w21063_
	);
	LUT3 #(
		.INIT('h80)
	) name10551 (
		\wishbone_bd_ram_mem0_reg[241][7]/P0001 ,
		_w11952_,
		_w11977_,
		_w21064_
	);
	LUT3 #(
		.INIT('h80)
	) name10552 (
		\wishbone_bd_ram_mem0_reg[93][7]/P0001 ,
		_w11966_,
		_w11972_,
		_w21065_
	);
	LUT3 #(
		.INIT('h80)
	) name10553 (
		\wishbone_bd_ram_mem0_reg[58][7]/P0001 ,
		_w11944_,
		_w11979_,
		_w21066_
	);
	LUT4 #(
		.INIT('h0001)
	) name10554 (
		_w21063_,
		_w21064_,
		_w21065_,
		_w21066_,
		_w21067_
	);
	LUT3 #(
		.INIT('h80)
	) name10555 (
		\wishbone_bd_ram_mem0_reg[27][7]/P0001 ,
		_w11935_,
		_w11936_,
		_w21068_
	);
	LUT3 #(
		.INIT('h80)
	) name10556 (
		\wishbone_bd_ram_mem0_reg[164][7]/P0001 ,
		_w11929_,
		_w11930_,
		_w21069_
	);
	LUT3 #(
		.INIT('h80)
	) name10557 (
		\wishbone_bd_ram_mem0_reg[216][7]/P0001 ,
		_w11984_,
		_w11990_,
		_w21070_
	);
	LUT3 #(
		.INIT('h80)
	) name10558 (
		\wishbone_bd_ram_mem0_reg[168][7]/P0001 ,
		_w11930_,
		_w11990_,
		_w21071_
	);
	LUT4 #(
		.INIT('h0001)
	) name10559 (
		_w21068_,
		_w21069_,
		_w21070_,
		_w21071_,
		_w21072_
	);
	LUT4 #(
		.INIT('h8000)
	) name10560 (
		_w21057_,
		_w21062_,
		_w21067_,
		_w21072_,
		_w21073_
	);
	LUT3 #(
		.INIT('h80)
	) name10561 (
		\wishbone_bd_ram_mem0_reg[203][7]/P0001 ,
		_w11936_,
		_w11945_,
		_w21074_
	);
	LUT3 #(
		.INIT('h80)
	) name10562 (
		\wishbone_bd_ram_mem0_reg[68][7]/P0001 ,
		_w11929_,
		_w11949_,
		_w21075_
	);
	LUT3 #(
		.INIT('h80)
	) name10563 (
		\wishbone_bd_ram_mem0_reg[197][7]/P0001 ,
		_w11933_,
		_w11945_,
		_w21076_
	);
	LUT3 #(
		.INIT('h80)
	) name10564 (
		\wishbone_bd_ram_mem0_reg[228][7]/P0001 ,
		_w11929_,
		_w11982_,
		_w21077_
	);
	LUT4 #(
		.INIT('h0001)
	) name10565 (
		_w21074_,
		_w21075_,
		_w21076_,
		_w21077_,
		_w21078_
	);
	LUT3 #(
		.INIT('h80)
	) name10566 (
		\wishbone_bd_ram_mem0_reg[143][7]/P0001 ,
		_w11955_,
		_w11973_,
		_w21079_
	);
	LUT3 #(
		.INIT('h80)
	) name10567 (
		\wishbone_bd_ram_mem0_reg[110][7]/P0001 ,
		_w11948_,
		_w11965_,
		_w21080_
	);
	LUT3 #(
		.INIT('h80)
	) name10568 (
		\wishbone_bd_ram_mem0_reg[167][7]/P0001 ,
		_w11930_,
		_w11975_,
		_w21081_
	);
	LUT3 #(
		.INIT('h80)
	) name10569 (
		\wishbone_bd_ram_mem0_reg[200][7]/P0001 ,
		_w11945_,
		_w11990_,
		_w21082_
	);
	LUT4 #(
		.INIT('h0001)
	) name10570 (
		_w21079_,
		_w21080_,
		_w21081_,
		_w21082_,
		_w21083_
	);
	LUT3 #(
		.INIT('h80)
	) name10571 (
		\wishbone_bd_ram_mem0_reg[50][7]/P0001 ,
		_w11963_,
		_w11979_,
		_w21084_
	);
	LUT3 #(
		.INIT('h80)
	) name10572 (
		\wishbone_bd_ram_mem0_reg[97][7]/P0001 ,
		_w11965_,
		_w11977_,
		_w21085_
	);
	LUT3 #(
		.INIT('h80)
	) name10573 (
		\wishbone_bd_ram_mem0_reg[175][7]/P0001 ,
		_w11930_,
		_w11973_,
		_w21086_
	);
	LUT3 #(
		.INIT('h80)
	) name10574 (
		\wishbone_bd_ram_mem0_reg[195][7]/P0001 ,
		_w11938_,
		_w11945_,
		_w21087_
	);
	LUT4 #(
		.INIT('h0001)
	) name10575 (
		_w21084_,
		_w21085_,
		_w21086_,
		_w21087_,
		_w21088_
	);
	LUT3 #(
		.INIT('h80)
	) name10576 (
		\wishbone_bd_ram_mem0_reg[229][7]/P0001 ,
		_w11933_,
		_w11982_,
		_w21089_
	);
	LUT3 #(
		.INIT('h80)
	) name10577 (
		\wishbone_bd_ram_mem0_reg[86][7]/P0001 ,
		_w11972_,
		_w11986_,
		_w21090_
	);
	LUT3 #(
		.INIT('h80)
	) name10578 (
		\wishbone_bd_ram_mem0_reg[208][7]/P0001 ,
		_w11941_,
		_w11984_,
		_w21091_
	);
	LUT3 #(
		.INIT('h80)
	) name10579 (
		\wishbone_bd_ram_mem0_reg[67][7]/P0001 ,
		_w11938_,
		_w11949_,
		_w21092_
	);
	LUT4 #(
		.INIT('h0001)
	) name10580 (
		_w21089_,
		_w21090_,
		_w21091_,
		_w21092_,
		_w21093_
	);
	LUT4 #(
		.INIT('h8000)
	) name10581 (
		_w21078_,
		_w21083_,
		_w21088_,
		_w21093_,
		_w21094_
	);
	LUT3 #(
		.INIT('h80)
	) name10582 (
		\wishbone_bd_ram_mem0_reg[146][7]/P0001 ,
		_w11959_,
		_w11963_,
		_w21095_
	);
	LUT3 #(
		.INIT('h80)
	) name10583 (
		\wishbone_bd_ram_mem0_reg[45][7]/P0001 ,
		_w11957_,
		_w11966_,
		_w21096_
	);
	LUT3 #(
		.INIT('h80)
	) name10584 (
		\wishbone_bd_ram_mem0_reg[106][7]/P0001 ,
		_w11944_,
		_w11965_,
		_w21097_
	);
	LUT3 #(
		.INIT('h80)
	) name10585 (
		\wishbone_bd_ram_mem0_reg[177][7]/P0001 ,
		_w11942_,
		_w11977_,
		_w21098_
	);
	LUT4 #(
		.INIT('h0001)
	) name10586 (
		_w21095_,
		_w21096_,
		_w21097_,
		_w21098_,
		_w21099_
	);
	LUT3 #(
		.INIT('h80)
	) name10587 (
		\wishbone_bd_ram_mem0_reg[48][7]/P0001 ,
		_w11941_,
		_w11979_,
		_w21100_
	);
	LUT3 #(
		.INIT('h80)
	) name10588 (
		\wishbone_bd_ram_mem0_reg[43][7]/P0001 ,
		_w11936_,
		_w11957_,
		_w21101_
	);
	LUT3 #(
		.INIT('h80)
	) name10589 (
		\wishbone_bd_ram_mem0_reg[142][7]/P0001 ,
		_w11948_,
		_w11955_,
		_w21102_
	);
	LUT3 #(
		.INIT('h80)
	) name10590 (
		\wishbone_bd_ram_mem0_reg[199][7]/P0001 ,
		_w11945_,
		_w11975_,
		_w21103_
	);
	LUT4 #(
		.INIT('h0001)
	) name10591 (
		_w21100_,
		_w21101_,
		_w21102_,
		_w21103_,
		_w21104_
	);
	LUT3 #(
		.INIT('h80)
	) name10592 (
		\wishbone_bd_ram_mem0_reg[36][7]/P0001 ,
		_w11929_,
		_w11957_,
		_w21105_
	);
	LUT3 #(
		.INIT('h80)
	) name10593 (
		\wishbone_bd_ram_mem0_reg[194][7]/P0001 ,
		_w11945_,
		_w11963_,
		_w21106_
	);
	LUT3 #(
		.INIT('h80)
	) name10594 (
		\wishbone_bd_ram_mem0_reg[202][7]/P0001 ,
		_w11944_,
		_w11945_,
		_w21107_
	);
	LUT3 #(
		.INIT('h80)
	) name10595 (
		\wishbone_bd_ram_mem0_reg[71][7]/P0001 ,
		_w11949_,
		_w11975_,
		_w21108_
	);
	LUT4 #(
		.INIT('h0001)
	) name10596 (
		_w21105_,
		_w21106_,
		_w21107_,
		_w21108_,
		_w21109_
	);
	LUT3 #(
		.INIT('h80)
	) name10597 (
		\wishbone_bd_ram_mem0_reg[53][7]/P0001 ,
		_w11933_,
		_w11979_,
		_w21110_
	);
	LUT3 #(
		.INIT('h80)
	) name10598 (
		\wishbone_bd_ram_mem0_reg[154][7]/P0001 ,
		_w11944_,
		_w11959_,
		_w21111_
	);
	LUT3 #(
		.INIT('h80)
	) name10599 (
		\wishbone_bd_ram_mem0_reg[12][7]/P0001 ,
		_w11932_,
		_w11954_,
		_w21112_
	);
	LUT3 #(
		.INIT('h80)
	) name10600 (
		\wishbone_bd_ram_mem0_reg[236][7]/P0001 ,
		_w11954_,
		_w11982_,
		_w21113_
	);
	LUT4 #(
		.INIT('h0001)
	) name10601 (
		_w21110_,
		_w21111_,
		_w21112_,
		_w21113_,
		_w21114_
	);
	LUT4 #(
		.INIT('h8000)
	) name10602 (
		_w21099_,
		_w21104_,
		_w21109_,
		_w21114_,
		_w21115_
	);
	LUT4 #(
		.INIT('h8000)
	) name10603 (
		_w21052_,
		_w21073_,
		_w21094_,
		_w21115_,
		_w21116_
	);
	LUT4 #(
		.INIT('h8000)
	) name10604 (
		_w20861_,
		_w20946_,
		_w21031_,
		_w21116_,
		_w21117_
	);
	LUT4 #(
		.INIT('h1555)
	) name10605 (
		wb_rst_i_pad,
		_w20763_,
		_w20767_,
		_w20775_,
		_w21118_
	);
	LUT3 #(
		.INIT('hba)
	) name10606 (
		_w20776_,
		_w21117_,
		_w21118_,
		_w21119_
	);
	LUT4 #(
		.INIT('h0002)
	) name10607 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21120_
	);
	LUT3 #(
		.INIT('h80)
	) name10608 (
		_w18757_,
		_w18758_,
		_w21120_,
		_w21121_
	);
	LUT3 #(
		.INIT('h80)
	) name10609 (
		\ethreg1_MODER_1_DataOut_reg[0]/NET0131 ,
		_w18800_,
		_w18801_,
		_w21122_
	);
	LUT3 #(
		.INIT('h80)
	) name10610 (
		\ethreg1_MIIRX_DATA_DataOut_reg[8]/NET0131 ,
		_w18785_,
		_w18786_,
		_w21123_
	);
	LUT4 #(
		.INIT('h0008)
	) name10611 (
		\ethreg1_RXHASH0_1_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21124_
	);
	LUT3 #(
		.INIT('h80)
	) name10612 (
		_w18757_,
		_w18758_,
		_w21124_,
		_w21125_
	);
	LUT4 #(
		.INIT('h0001)
	) name10613 (
		_w21121_,
		_w21122_,
		_w21123_,
		_w21125_,
		_w21126_
	);
	LUT3 #(
		.INIT('h80)
	) name10614 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[0]/NET0131 ,
		_w18798_,
		_w18805_,
		_w21127_
	);
	LUT3 #(
		.INIT('h80)
	) name10615 (
		\ethreg1_MIIMODER_1_DataOut_reg[0]/NET0131 ,
		_w18786_,
		_w18801_,
		_w21128_
	);
	LUT2 #(
		.INIT('h1)
	) name10616 (
		_w21127_,
		_w21128_,
		_w21129_
	);
	LUT3 #(
		.INIT('h02)
	) name10617 (
		_w18752_,
		_w21127_,
		_w21128_,
		_w21130_
	);
	LUT3 #(
		.INIT('h80)
	) name10618 (
		\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 ,
		_w18753_,
		_w18754_,
		_w21131_
	);
	LUT4 #(
		.INIT('h0008)
	) name10619 (
		\ethreg1_RXHASH1_1_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21132_
	);
	LUT4 #(
		.INIT('h0002)
	) name10620 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21133_
	);
	LUT4 #(
		.INIT('h777f)
	) name10621 (
		_w18757_,
		_w18762_,
		_w21132_,
		_w21133_,
		_w21134_
	);
	LUT4 #(
		.INIT('h0020)
	) name10622 (
		\ethreg1_TXCTRL_1_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21135_
	);
	LUT3 #(
		.INIT('h80)
	) name10623 (
		_w18757_,
		_w18758_,
		_w21135_,
		_w21136_
	);
	LUT3 #(
		.INIT('h80)
	) name10624 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[0]/NET0131 ,
		_w18785_,
		_w18798_,
		_w21137_
	);
	LUT4 #(
		.INIT('h0004)
	) name10625 (
		_w21131_,
		_w21134_,
		_w21136_,
		_w21137_,
		_w21138_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10626 (
		_w18752_,
		_w21126_,
		_w21129_,
		_w21138_,
		_w21139_
	);
	LUT3 #(
		.INIT('h80)
	) name10627 (
		\wishbone_bd_ram_mem1_reg[239][8]/P0001 ,
		_w11973_,
		_w11982_,
		_w21140_
	);
	LUT3 #(
		.INIT('h80)
	) name10628 (
		\wishbone_bd_ram_mem1_reg[33][8]/P0001 ,
		_w11957_,
		_w11977_,
		_w21141_
	);
	LUT3 #(
		.INIT('h80)
	) name10629 (
		\wishbone_bd_ram_mem1_reg[72][8]/P0001 ,
		_w11949_,
		_w11990_,
		_w21142_
	);
	LUT3 #(
		.INIT('h80)
	) name10630 (
		\wishbone_bd_ram_mem1_reg[223][8]/P0001 ,
		_w11973_,
		_w11984_,
		_w21143_
	);
	LUT4 #(
		.INIT('h0001)
	) name10631 (
		_w21140_,
		_w21141_,
		_w21142_,
		_w21143_,
		_w21144_
	);
	LUT3 #(
		.INIT('h80)
	) name10632 (
		\wishbone_bd_ram_mem1_reg[92][8]/P0001 ,
		_w11954_,
		_w11972_,
		_w21145_
	);
	LUT3 #(
		.INIT('h80)
	) name10633 (
		\wishbone_bd_ram_mem1_reg[232][8]/P0001 ,
		_w11982_,
		_w11990_,
		_w21146_
	);
	LUT3 #(
		.INIT('h80)
	) name10634 (
		\wishbone_bd_ram_mem1_reg[118][8]/P0001 ,
		_w11986_,
		_w12012_,
		_w21147_
	);
	LUT3 #(
		.INIT('h80)
	) name10635 (
		\wishbone_bd_ram_mem1_reg[4][8]/P0001 ,
		_w11929_,
		_w11932_,
		_w21148_
	);
	LUT4 #(
		.INIT('h0001)
	) name10636 (
		_w21145_,
		_w21146_,
		_w21147_,
		_w21148_,
		_w21149_
	);
	LUT3 #(
		.INIT('h80)
	) name10637 (
		\wishbone_bd_ram_mem1_reg[190][8]/P0001 ,
		_w11942_,
		_w11948_,
		_w21150_
	);
	LUT3 #(
		.INIT('h80)
	) name10638 (
		\wishbone_bd_ram_mem1_reg[43][8]/P0001 ,
		_w11936_,
		_w11957_,
		_w21151_
	);
	LUT3 #(
		.INIT('h80)
	) name10639 (
		\wishbone_bd_ram_mem1_reg[57][8]/P0001 ,
		_w11968_,
		_w11979_,
		_w21152_
	);
	LUT3 #(
		.INIT('h80)
	) name10640 (
		\wishbone_bd_ram_mem1_reg[188][8]/P0001 ,
		_w11942_,
		_w11954_,
		_w21153_
	);
	LUT4 #(
		.INIT('h0001)
	) name10641 (
		_w21150_,
		_w21151_,
		_w21152_,
		_w21153_,
		_w21154_
	);
	LUT3 #(
		.INIT('h80)
	) name10642 (
		\wishbone_bd_ram_mem1_reg[35][8]/P0001 ,
		_w11938_,
		_w11957_,
		_w21155_
	);
	LUT3 #(
		.INIT('h80)
	) name10643 (
		\wishbone_bd_ram_mem1_reg[226][8]/P0001 ,
		_w11963_,
		_w11982_,
		_w21156_
	);
	LUT3 #(
		.INIT('h80)
	) name10644 (
		\wishbone_bd_ram_mem1_reg[66][8]/P0001 ,
		_w11949_,
		_w11963_,
		_w21157_
	);
	LUT3 #(
		.INIT('h80)
	) name10645 (
		\wishbone_bd_ram_mem1_reg[89][8]/P0001 ,
		_w11968_,
		_w11972_,
		_w21158_
	);
	LUT4 #(
		.INIT('h0001)
	) name10646 (
		_w21155_,
		_w21156_,
		_w21157_,
		_w21158_,
		_w21159_
	);
	LUT4 #(
		.INIT('h8000)
	) name10647 (
		_w21144_,
		_w21149_,
		_w21154_,
		_w21159_,
		_w21160_
	);
	LUT3 #(
		.INIT('h80)
	) name10648 (
		\wishbone_bd_ram_mem1_reg[145][8]/P0001 ,
		_w11959_,
		_w11977_,
		_w21161_
	);
	LUT3 #(
		.INIT('h80)
	) name10649 (
		\wishbone_bd_ram_mem1_reg[174][8]/P0001 ,
		_w11930_,
		_w11948_,
		_w21162_
	);
	LUT3 #(
		.INIT('h80)
	) name10650 (
		\wishbone_bd_ram_mem1_reg[42][8]/P0001 ,
		_w11944_,
		_w11957_,
		_w21163_
	);
	LUT3 #(
		.INIT('h80)
	) name10651 (
		\wishbone_bd_ram_mem1_reg[117][8]/P0001 ,
		_w11933_,
		_w12012_,
		_w21164_
	);
	LUT4 #(
		.INIT('h0001)
	) name10652 (
		_w21161_,
		_w21162_,
		_w21163_,
		_w21164_,
		_w21165_
	);
	LUT3 #(
		.INIT('h80)
	) name10653 (
		\wishbone_bd_ram_mem1_reg[229][8]/P0001 ,
		_w11933_,
		_w11982_,
		_w21166_
	);
	LUT3 #(
		.INIT('h80)
	) name10654 (
		\wishbone_bd_ram_mem1_reg[127][8]/P0001 ,
		_w11973_,
		_w12012_,
		_w21167_
	);
	LUT3 #(
		.INIT('h80)
	) name10655 (
		\wishbone_bd_ram_mem1_reg[46][8]/P0001 ,
		_w11948_,
		_w11957_,
		_w21168_
	);
	LUT3 #(
		.INIT('h80)
	) name10656 (
		\wishbone_bd_ram_mem1_reg[44][8]/P0001 ,
		_w11954_,
		_w11957_,
		_w21169_
	);
	LUT4 #(
		.INIT('h0001)
	) name10657 (
		_w21166_,
		_w21167_,
		_w21168_,
		_w21169_,
		_w21170_
	);
	LUT3 #(
		.INIT('h80)
	) name10658 (
		\wishbone_bd_ram_mem1_reg[180][8]/P0001 ,
		_w11929_,
		_w11942_,
		_w21171_
	);
	LUT3 #(
		.INIT('h80)
	) name10659 (
		\wishbone_bd_ram_mem1_reg[178][8]/P0001 ,
		_w11942_,
		_w11963_,
		_w21172_
	);
	LUT3 #(
		.INIT('h80)
	) name10660 (
		\wishbone_bd_ram_mem1_reg[252][8]/P0001 ,
		_w11952_,
		_w11954_,
		_w21173_
	);
	LUT3 #(
		.INIT('h80)
	) name10661 (
		\wishbone_bd_ram_mem1_reg[5][8]/P0001 ,
		_w11932_,
		_w11933_,
		_w21174_
	);
	LUT4 #(
		.INIT('h0001)
	) name10662 (
		_w21171_,
		_w21172_,
		_w21173_,
		_w21174_,
		_w21175_
	);
	LUT3 #(
		.INIT('h80)
	) name10663 (
		\wishbone_bd_ram_mem1_reg[18][8]/P0001 ,
		_w11935_,
		_w11963_,
		_w21176_
	);
	LUT3 #(
		.INIT('h80)
	) name10664 (
		\wishbone_bd_ram_mem1_reg[211][8]/P0001 ,
		_w11938_,
		_w11984_,
		_w21177_
	);
	LUT3 #(
		.INIT('h80)
	) name10665 (
		\wishbone_bd_ram_mem1_reg[171][8]/P0001 ,
		_w11930_,
		_w11936_,
		_w21178_
	);
	LUT3 #(
		.INIT('h80)
	) name10666 (
		\wishbone_bd_ram_mem1_reg[48][8]/P0001 ,
		_w11941_,
		_w11979_,
		_w21179_
	);
	LUT4 #(
		.INIT('h0001)
	) name10667 (
		_w21176_,
		_w21177_,
		_w21178_,
		_w21179_,
		_w21180_
	);
	LUT4 #(
		.INIT('h8000)
	) name10668 (
		_w21165_,
		_w21170_,
		_w21175_,
		_w21180_,
		_w21181_
	);
	LUT3 #(
		.INIT('h80)
	) name10669 (
		\wishbone_bd_ram_mem1_reg[255][8]/P0001 ,
		_w11952_,
		_w11973_,
		_w21182_
	);
	LUT3 #(
		.INIT('h80)
	) name10670 (
		\wishbone_bd_ram_mem1_reg[111][8]/P0001 ,
		_w11965_,
		_w11973_,
		_w21183_
	);
	LUT3 #(
		.INIT('h80)
	) name10671 (
		\wishbone_bd_ram_mem1_reg[210][8]/P0001 ,
		_w11963_,
		_w11984_,
		_w21184_
	);
	LUT3 #(
		.INIT('h80)
	) name10672 (
		\wishbone_bd_ram_mem1_reg[19][8]/P0001 ,
		_w11935_,
		_w11938_,
		_w21185_
	);
	LUT4 #(
		.INIT('h0001)
	) name10673 (
		_w21182_,
		_w21183_,
		_w21184_,
		_w21185_,
		_w21186_
	);
	LUT3 #(
		.INIT('h80)
	) name10674 (
		\wishbone_bd_ram_mem1_reg[204][8]/P0001 ,
		_w11945_,
		_w11954_,
		_w21187_
	);
	LUT3 #(
		.INIT('h80)
	) name10675 (
		\wishbone_bd_ram_mem1_reg[160][8]/P0001 ,
		_w11930_,
		_w11941_,
		_w21188_
	);
	LUT3 #(
		.INIT('h80)
	) name10676 (
		\wishbone_bd_ram_mem1_reg[97][8]/P0001 ,
		_w11965_,
		_w11977_,
		_w21189_
	);
	LUT3 #(
		.INIT('h80)
	) name10677 (
		\wishbone_bd_ram_mem1_reg[120][8]/P0001 ,
		_w11990_,
		_w12012_,
		_w21190_
	);
	LUT4 #(
		.INIT('h0001)
	) name10678 (
		_w21187_,
		_w21188_,
		_w21189_,
		_w21190_,
		_w21191_
	);
	LUT3 #(
		.INIT('h80)
	) name10679 (
		\wishbone_bd_ram_mem1_reg[156][8]/P0001 ,
		_w11954_,
		_w11959_,
		_w21192_
	);
	LUT3 #(
		.INIT('h80)
	) name10680 (
		\wishbone_bd_ram_mem1_reg[31][8]/P0001 ,
		_w11935_,
		_w11973_,
		_w21193_
	);
	LUT3 #(
		.INIT('h80)
	) name10681 (
		\wishbone_bd_ram_mem1_reg[99][8]/P0001 ,
		_w11938_,
		_w11965_,
		_w21194_
	);
	LUT3 #(
		.INIT('h80)
	) name10682 (
		\wishbone_bd_ram_mem1_reg[91][8]/P0001 ,
		_w11936_,
		_w11972_,
		_w21195_
	);
	LUT4 #(
		.INIT('h0001)
	) name10683 (
		_w21192_,
		_w21193_,
		_w21194_,
		_w21195_,
		_w21196_
	);
	LUT3 #(
		.INIT('h80)
	) name10684 (
		\wishbone_bd_ram_mem1_reg[198][8]/P0001 ,
		_w11945_,
		_w11986_,
		_w21197_
	);
	LUT3 #(
		.INIT('h80)
	) name10685 (
		\wishbone_bd_ram_mem1_reg[32][8]/P0001 ,
		_w11941_,
		_w11957_,
		_w21198_
	);
	LUT3 #(
		.INIT('h80)
	) name10686 (
		\wishbone_bd_ram_mem1_reg[49][8]/P0001 ,
		_w11977_,
		_w11979_,
		_w21199_
	);
	LUT3 #(
		.INIT('h80)
	) name10687 (
		\wishbone_bd_ram_mem1_reg[251][8]/P0001 ,
		_w11936_,
		_w11952_,
		_w21200_
	);
	LUT4 #(
		.INIT('h0001)
	) name10688 (
		_w21197_,
		_w21198_,
		_w21199_,
		_w21200_,
		_w21201_
	);
	LUT4 #(
		.INIT('h8000)
	) name10689 (
		_w21186_,
		_w21191_,
		_w21196_,
		_w21201_,
		_w21202_
	);
	LUT3 #(
		.INIT('h80)
	) name10690 (
		\wishbone_bd_ram_mem1_reg[129][8]/P0001 ,
		_w11955_,
		_w11977_,
		_w21203_
	);
	LUT3 #(
		.INIT('h80)
	) name10691 (
		\wishbone_bd_ram_mem1_reg[104][8]/P0001 ,
		_w11965_,
		_w11990_,
		_w21204_
	);
	LUT3 #(
		.INIT('h80)
	) name10692 (
		\wishbone_bd_ram_mem1_reg[107][8]/P0001 ,
		_w11936_,
		_w11965_,
		_w21205_
	);
	LUT3 #(
		.INIT('h80)
	) name10693 (
		\wishbone_bd_ram_mem1_reg[231][8]/P0001 ,
		_w11975_,
		_w11982_,
		_w21206_
	);
	LUT4 #(
		.INIT('h0001)
	) name10694 (
		_w21203_,
		_w21204_,
		_w21205_,
		_w21206_,
		_w21207_
	);
	LUT3 #(
		.INIT('h80)
	) name10695 (
		\wishbone_bd_ram_mem1_reg[181][8]/P0001 ,
		_w11933_,
		_w11942_,
		_w21208_
	);
	LUT3 #(
		.INIT('h80)
	) name10696 (
		\wishbone_bd_ram_mem1_reg[113][8]/P0001 ,
		_w11977_,
		_w12012_,
		_w21209_
	);
	LUT3 #(
		.INIT('h80)
	) name10697 (
		\wishbone_bd_ram_mem1_reg[85][8]/P0001 ,
		_w11933_,
		_w11972_,
		_w21210_
	);
	LUT3 #(
		.INIT('h80)
	) name10698 (
		\wishbone_bd_ram_mem1_reg[30][8]/P0001 ,
		_w11935_,
		_w11948_,
		_w21211_
	);
	LUT4 #(
		.INIT('h0001)
	) name10699 (
		_w21208_,
		_w21209_,
		_w21210_,
		_w21211_,
		_w21212_
	);
	LUT3 #(
		.INIT('h80)
	) name10700 (
		\wishbone_bd_ram_mem1_reg[202][8]/P0001 ,
		_w11944_,
		_w11945_,
		_w21213_
	);
	LUT3 #(
		.INIT('h80)
	) name10701 (
		\wishbone_bd_ram_mem1_reg[86][8]/P0001 ,
		_w11972_,
		_w11986_,
		_w21214_
	);
	LUT3 #(
		.INIT('h80)
	) name10702 (
		\wishbone_bd_ram_mem1_reg[137][8]/P0001 ,
		_w11955_,
		_w11968_,
		_w21215_
	);
	LUT3 #(
		.INIT('h80)
	) name10703 (
		\wishbone_bd_ram_mem1_reg[29][8]/P0001 ,
		_w11935_,
		_w11966_,
		_w21216_
	);
	LUT4 #(
		.INIT('h0001)
	) name10704 (
		_w21213_,
		_w21214_,
		_w21215_,
		_w21216_,
		_w21217_
	);
	LUT3 #(
		.INIT('h80)
	) name10705 (
		\wishbone_bd_ram_mem1_reg[159][8]/P0001 ,
		_w11959_,
		_w11973_,
		_w21218_
	);
	LUT3 #(
		.INIT('h80)
	) name10706 (
		\wishbone_bd_ram_mem1_reg[240][8]/P0001 ,
		_w11941_,
		_w11952_,
		_w21219_
	);
	LUT3 #(
		.INIT('h80)
	) name10707 (
		\wishbone_bd_ram_mem1_reg[16][8]/P0001 ,
		_w11935_,
		_w11941_,
		_w21220_
	);
	LUT3 #(
		.INIT('h80)
	) name10708 (
		\wishbone_bd_ram_mem1_reg[68][8]/P0001 ,
		_w11929_,
		_w11949_,
		_w21221_
	);
	LUT4 #(
		.INIT('h0001)
	) name10709 (
		_w21218_,
		_w21219_,
		_w21220_,
		_w21221_,
		_w21222_
	);
	LUT4 #(
		.INIT('h8000)
	) name10710 (
		_w21207_,
		_w21212_,
		_w21217_,
		_w21222_,
		_w21223_
	);
	LUT4 #(
		.INIT('h8000)
	) name10711 (
		_w21160_,
		_w21181_,
		_w21202_,
		_w21223_,
		_w21224_
	);
	LUT3 #(
		.INIT('h80)
	) name10712 (
		\wishbone_bd_ram_mem1_reg[78][8]/P0001 ,
		_w11948_,
		_w11949_,
		_w21225_
	);
	LUT3 #(
		.INIT('h80)
	) name10713 (
		\wishbone_bd_ram_mem1_reg[228][8]/P0001 ,
		_w11929_,
		_w11982_,
		_w21226_
	);
	LUT3 #(
		.INIT('h80)
	) name10714 (
		\wishbone_bd_ram_mem1_reg[236][8]/P0001 ,
		_w11954_,
		_w11982_,
		_w21227_
	);
	LUT3 #(
		.INIT('h80)
	) name10715 (
		\wishbone_bd_ram_mem1_reg[144][8]/P0001 ,
		_w11941_,
		_w11959_,
		_w21228_
	);
	LUT4 #(
		.INIT('h0001)
	) name10716 (
		_w21225_,
		_w21226_,
		_w21227_,
		_w21228_,
		_w21229_
	);
	LUT3 #(
		.INIT('h80)
	) name10717 (
		\wishbone_bd_ram_mem1_reg[166][8]/P0001 ,
		_w11930_,
		_w11986_,
		_w21230_
	);
	LUT3 #(
		.INIT('h80)
	) name10718 (
		\wishbone_bd_ram_mem1_reg[133][8]/P0001 ,
		_w11933_,
		_w11955_,
		_w21231_
	);
	LUT3 #(
		.INIT('h80)
	) name10719 (
		\wishbone_bd_ram_mem1_reg[170][8]/P0001 ,
		_w11930_,
		_w11944_,
		_w21232_
	);
	LUT3 #(
		.INIT('h80)
	) name10720 (
		\wishbone_bd_ram_mem1_reg[173][8]/P0001 ,
		_w11930_,
		_w11966_,
		_w21233_
	);
	LUT4 #(
		.INIT('h0001)
	) name10721 (
		_w21230_,
		_w21231_,
		_w21232_,
		_w21233_,
		_w21234_
	);
	LUT3 #(
		.INIT('h80)
	) name10722 (
		\wishbone_bd_ram_mem1_reg[237][8]/P0001 ,
		_w11966_,
		_w11982_,
		_w21235_
	);
	LUT3 #(
		.INIT('h80)
	) name10723 (
		\wishbone_bd_ram_mem1_reg[59][8]/P0001 ,
		_w11936_,
		_w11979_,
		_w21236_
	);
	LUT3 #(
		.INIT('h80)
	) name10724 (
		\wishbone_bd_ram_mem1_reg[184][8]/P0001 ,
		_w11942_,
		_w11990_,
		_w21237_
	);
	LUT3 #(
		.INIT('h80)
	) name10725 (
		\wishbone_bd_ram_mem1_reg[95][8]/P0001 ,
		_w11972_,
		_w11973_,
		_w21238_
	);
	LUT4 #(
		.INIT('h0001)
	) name10726 (
		_w21235_,
		_w21236_,
		_w21237_,
		_w21238_,
		_w21239_
	);
	LUT3 #(
		.INIT('h80)
	) name10727 (
		\wishbone_bd_ram_mem1_reg[186][8]/P0001 ,
		_w11942_,
		_w11944_,
		_w21240_
	);
	LUT3 #(
		.INIT('h80)
	) name10728 (
		\wishbone_bd_ram_mem1_reg[131][8]/P0001 ,
		_w11938_,
		_w11955_,
		_w21241_
	);
	LUT3 #(
		.INIT('h80)
	) name10729 (
		\wishbone_bd_ram_mem1_reg[143][8]/P0001 ,
		_w11955_,
		_w11973_,
		_w21242_
	);
	LUT3 #(
		.INIT('h80)
	) name10730 (
		\wishbone_bd_ram_mem1_reg[193][8]/P0001 ,
		_w11945_,
		_w11977_,
		_w21243_
	);
	LUT4 #(
		.INIT('h0001)
	) name10731 (
		_w21240_,
		_w21241_,
		_w21242_,
		_w21243_,
		_w21244_
	);
	LUT4 #(
		.INIT('h8000)
	) name10732 (
		_w21229_,
		_w21234_,
		_w21239_,
		_w21244_,
		_w21245_
	);
	LUT3 #(
		.INIT('h80)
	) name10733 (
		\wishbone_bd_ram_mem1_reg[98][8]/P0001 ,
		_w11963_,
		_w11965_,
		_w21246_
	);
	LUT3 #(
		.INIT('h80)
	) name10734 (
		\wishbone_bd_ram_mem1_reg[84][8]/P0001 ,
		_w11929_,
		_w11972_,
		_w21247_
	);
	LUT3 #(
		.INIT('h80)
	) name10735 (
		\wishbone_bd_ram_mem1_reg[148][8]/P0001 ,
		_w11929_,
		_w11959_,
		_w21248_
	);
	LUT3 #(
		.INIT('h80)
	) name10736 (
		\wishbone_bd_ram_mem1_reg[115][8]/P0001 ,
		_w11938_,
		_w12012_,
		_w21249_
	);
	LUT4 #(
		.INIT('h0001)
	) name10737 (
		_w21246_,
		_w21247_,
		_w21248_,
		_w21249_,
		_w21250_
	);
	LUT3 #(
		.INIT('h80)
	) name10738 (
		\wishbone_bd_ram_mem1_reg[2][8]/P0001 ,
		_w11932_,
		_w11963_,
		_w21251_
	);
	LUT3 #(
		.INIT('h80)
	) name10739 (
		\wishbone_bd_ram_mem1_reg[56][8]/P0001 ,
		_w11979_,
		_w11990_,
		_w21252_
	);
	LUT3 #(
		.INIT('h80)
	) name10740 (
		\wishbone_bd_ram_mem1_reg[27][8]/P0001 ,
		_w11935_,
		_w11936_,
		_w21253_
	);
	LUT3 #(
		.INIT('h80)
	) name10741 (
		\wishbone_bd_ram_mem1_reg[189][8]/P0001 ,
		_w11942_,
		_w11966_,
		_w21254_
	);
	LUT4 #(
		.INIT('h0001)
	) name10742 (
		_w21251_,
		_w21252_,
		_w21253_,
		_w21254_,
		_w21255_
	);
	LUT3 #(
		.INIT('h80)
	) name10743 (
		\wishbone_bd_ram_mem1_reg[50][8]/P0001 ,
		_w11963_,
		_w11979_,
		_w21256_
	);
	LUT3 #(
		.INIT('h80)
	) name10744 (
		\wishbone_bd_ram_mem1_reg[177][8]/P0001 ,
		_w11942_,
		_w11977_,
		_w21257_
	);
	LUT3 #(
		.INIT('h80)
	) name10745 (
		\wishbone_bd_ram_mem1_reg[135][8]/P0001 ,
		_w11955_,
		_w11975_,
		_w21258_
	);
	LUT3 #(
		.INIT('h80)
	) name10746 (
		\wishbone_bd_ram_mem1_reg[51][8]/P0001 ,
		_w11938_,
		_w11979_,
		_w21259_
	);
	LUT4 #(
		.INIT('h0001)
	) name10747 (
		_w21256_,
		_w21257_,
		_w21258_,
		_w21259_,
		_w21260_
	);
	LUT3 #(
		.INIT('h80)
	) name10748 (
		\wishbone_bd_ram_mem1_reg[3][8]/P0001 ,
		_w11932_,
		_w11938_,
		_w21261_
	);
	LUT3 #(
		.INIT('h80)
	) name10749 (
		\wishbone_bd_ram_mem1_reg[253][8]/P0001 ,
		_w11952_,
		_w11966_,
		_w21262_
	);
	LUT3 #(
		.INIT('h80)
	) name10750 (
		\wishbone_bd_ram_mem1_reg[191][8]/P0001 ,
		_w11942_,
		_w11973_,
		_w21263_
	);
	LUT3 #(
		.INIT('h80)
	) name10751 (
		\wishbone_bd_ram_mem1_reg[152][8]/P0001 ,
		_w11959_,
		_w11990_,
		_w21264_
	);
	LUT4 #(
		.INIT('h0001)
	) name10752 (
		_w21261_,
		_w21262_,
		_w21263_,
		_w21264_,
		_w21265_
	);
	LUT4 #(
		.INIT('h8000)
	) name10753 (
		_w21250_,
		_w21255_,
		_w21260_,
		_w21265_,
		_w21266_
	);
	LUT3 #(
		.INIT('h80)
	) name10754 (
		\wishbone_bd_ram_mem1_reg[165][8]/P0001 ,
		_w11930_,
		_w11933_,
		_w21267_
	);
	LUT3 #(
		.INIT('h80)
	) name10755 (
		\wishbone_bd_ram_mem1_reg[10][8]/P0001 ,
		_w11932_,
		_w11944_,
		_w21268_
	);
	LUT3 #(
		.INIT('h80)
	) name10756 (
		\wishbone_bd_ram_mem1_reg[125][8]/P0001 ,
		_w11966_,
		_w12012_,
		_w21269_
	);
	LUT3 #(
		.INIT('h80)
	) name10757 (
		\wishbone_bd_ram_mem1_reg[140][8]/P0001 ,
		_w11954_,
		_w11955_,
		_w21270_
	);
	LUT4 #(
		.INIT('h0001)
	) name10758 (
		_w21267_,
		_w21268_,
		_w21269_,
		_w21270_,
		_w21271_
	);
	LUT3 #(
		.INIT('h80)
	) name10759 (
		\wishbone_bd_ram_mem1_reg[205][8]/P0001 ,
		_w11945_,
		_w11966_,
		_w21272_
	);
	LUT3 #(
		.INIT('h80)
	) name10760 (
		\wishbone_bd_ram_mem1_reg[201][8]/P0001 ,
		_w11945_,
		_w11968_,
		_w21273_
	);
	LUT3 #(
		.INIT('h80)
	) name10761 (
		\wishbone_bd_ram_mem1_reg[1][8]/P0001 ,
		_w11932_,
		_w11977_,
		_w21274_
	);
	LUT3 #(
		.INIT('h80)
	) name10762 (
		\wishbone_bd_ram_mem1_reg[96][8]/P0001 ,
		_w11941_,
		_w11965_,
		_w21275_
	);
	LUT4 #(
		.INIT('h0001)
	) name10763 (
		_w21272_,
		_w21273_,
		_w21274_,
		_w21275_,
		_w21276_
	);
	LUT3 #(
		.INIT('h80)
	) name10764 (
		\wishbone_bd_ram_mem1_reg[213][8]/P0001 ,
		_w11933_,
		_w11984_,
		_w21277_
	);
	LUT3 #(
		.INIT('h80)
	) name10765 (
		\wishbone_bd_ram_mem1_reg[161][8]/P0001 ,
		_w11930_,
		_w11977_,
		_w21278_
	);
	LUT3 #(
		.INIT('h80)
	) name10766 (
		\wishbone_bd_ram_mem1_reg[163][8]/P0001 ,
		_w11930_,
		_w11938_,
		_w21279_
	);
	LUT3 #(
		.INIT('h80)
	) name10767 (
		\wishbone_bd_ram_mem1_reg[185][8]/P0001 ,
		_w11942_,
		_w11968_,
		_w21280_
	);
	LUT4 #(
		.INIT('h0001)
	) name10768 (
		_w21277_,
		_w21278_,
		_w21279_,
		_w21280_,
		_w21281_
	);
	LUT3 #(
		.INIT('h80)
	) name10769 (
		\wishbone_bd_ram_mem1_reg[121][8]/P0001 ,
		_w11968_,
		_w12012_,
		_w21282_
	);
	LUT3 #(
		.INIT('h80)
	) name10770 (
		\wishbone_bd_ram_mem1_reg[254][8]/P0001 ,
		_w11948_,
		_w11952_,
		_w21283_
	);
	LUT3 #(
		.INIT('h80)
	) name10771 (
		\wishbone_bd_ram_mem1_reg[101][8]/P0001 ,
		_w11933_,
		_w11965_,
		_w21284_
	);
	LUT3 #(
		.INIT('h80)
	) name10772 (
		\wishbone_bd_ram_mem1_reg[162][8]/P0001 ,
		_w11930_,
		_w11963_,
		_w21285_
	);
	LUT4 #(
		.INIT('h0001)
	) name10773 (
		_w21282_,
		_w21283_,
		_w21284_,
		_w21285_,
		_w21286_
	);
	LUT4 #(
		.INIT('h8000)
	) name10774 (
		_w21271_,
		_w21276_,
		_w21281_,
		_w21286_,
		_w21287_
	);
	LUT3 #(
		.INIT('h80)
	) name10775 (
		\wishbone_bd_ram_mem1_reg[119][8]/P0001 ,
		_w11975_,
		_w12012_,
		_w21288_
	);
	LUT3 #(
		.INIT('h80)
	) name10776 (
		\wishbone_bd_ram_mem1_reg[138][8]/P0001 ,
		_w11944_,
		_w11955_,
		_w21289_
	);
	LUT3 #(
		.INIT('h80)
	) name10777 (
		\wishbone_bd_ram_mem1_reg[241][8]/P0001 ,
		_w11952_,
		_w11977_,
		_w21290_
	);
	LUT3 #(
		.INIT('h80)
	) name10778 (
		\wishbone_bd_ram_mem1_reg[36][8]/P0001 ,
		_w11929_,
		_w11957_,
		_w21291_
	);
	LUT4 #(
		.INIT('h0001)
	) name10779 (
		_w21288_,
		_w21289_,
		_w21290_,
		_w21291_,
		_w21292_
	);
	LUT3 #(
		.INIT('h80)
	) name10780 (
		\wishbone_bd_ram_mem1_reg[168][8]/P0001 ,
		_w11930_,
		_w11990_,
		_w21293_
	);
	LUT3 #(
		.INIT('h80)
	) name10781 (
		\wishbone_bd_ram_mem1_reg[221][8]/P0001 ,
		_w11966_,
		_w11984_,
		_w21294_
	);
	LUT3 #(
		.INIT('h80)
	) name10782 (
		\wishbone_bd_ram_mem1_reg[25][8]/P0001 ,
		_w11935_,
		_w11968_,
		_w21295_
	);
	LUT3 #(
		.INIT('h80)
	) name10783 (
		\wishbone_bd_ram_mem1_reg[218][8]/P0001 ,
		_w11944_,
		_w11984_,
		_w21296_
	);
	LUT4 #(
		.INIT('h0001)
	) name10784 (
		_w21293_,
		_w21294_,
		_w21295_,
		_w21296_,
		_w21297_
	);
	LUT3 #(
		.INIT('h80)
	) name10785 (
		\wishbone_bd_ram_mem1_reg[58][8]/P0001 ,
		_w11944_,
		_w11979_,
		_w21298_
	);
	LUT3 #(
		.INIT('h80)
	) name10786 (
		\wishbone_bd_ram_mem1_reg[123][8]/P0001 ,
		_w11936_,
		_w12012_,
		_w21299_
	);
	LUT3 #(
		.INIT('h80)
	) name10787 (
		\wishbone_bd_ram_mem1_reg[75][8]/P0001 ,
		_w11936_,
		_w11949_,
		_w21300_
	);
	LUT3 #(
		.INIT('h80)
	) name10788 (
		\wishbone_bd_ram_mem1_reg[215][8]/P0001 ,
		_w11975_,
		_w11984_,
		_w21301_
	);
	LUT4 #(
		.INIT('h0001)
	) name10789 (
		_w21298_,
		_w21299_,
		_w21300_,
		_w21301_,
		_w21302_
	);
	LUT3 #(
		.INIT('h80)
	) name10790 (
		\wishbone_bd_ram_mem1_reg[200][8]/P0001 ,
		_w11945_,
		_w11990_,
		_w21303_
	);
	LUT3 #(
		.INIT('h80)
	) name10791 (
		\wishbone_bd_ram_mem1_reg[249][8]/P0001 ,
		_w11952_,
		_w11968_,
		_w21304_
	);
	LUT3 #(
		.INIT('h80)
	) name10792 (
		\wishbone_bd_ram_mem1_reg[151][8]/P0001 ,
		_w11959_,
		_w11975_,
		_w21305_
	);
	LUT3 #(
		.INIT('h80)
	) name10793 (
		\wishbone_bd_ram_mem1_reg[157][8]/P0001 ,
		_w11959_,
		_w11966_,
		_w21306_
	);
	LUT4 #(
		.INIT('h0001)
	) name10794 (
		_w21303_,
		_w21304_,
		_w21305_,
		_w21306_,
		_w21307_
	);
	LUT4 #(
		.INIT('h8000)
	) name10795 (
		_w21292_,
		_w21297_,
		_w21302_,
		_w21307_,
		_w21308_
	);
	LUT4 #(
		.INIT('h8000)
	) name10796 (
		_w21245_,
		_w21266_,
		_w21287_,
		_w21308_,
		_w21309_
	);
	LUT3 #(
		.INIT('h80)
	) name10797 (
		\wishbone_bd_ram_mem1_reg[21][8]/P0001 ,
		_w11933_,
		_w11935_,
		_w21310_
	);
	LUT3 #(
		.INIT('h80)
	) name10798 (
		\wishbone_bd_ram_mem1_reg[164][8]/P0001 ,
		_w11929_,
		_w11930_,
		_w21311_
	);
	LUT3 #(
		.INIT('h80)
	) name10799 (
		\wishbone_bd_ram_mem1_reg[81][8]/P0001 ,
		_w11972_,
		_w11977_,
		_w21312_
	);
	LUT3 #(
		.INIT('h80)
	) name10800 (
		\wishbone_bd_ram_mem1_reg[187][8]/P0001 ,
		_w11936_,
		_w11942_,
		_w21313_
	);
	LUT4 #(
		.INIT('h0001)
	) name10801 (
		_w21310_,
		_w21311_,
		_w21312_,
		_w21313_,
		_w21314_
	);
	LUT3 #(
		.INIT('h80)
	) name10802 (
		\wishbone_bd_ram_mem1_reg[126][8]/P0001 ,
		_w11948_,
		_w12012_,
		_w21315_
	);
	LUT3 #(
		.INIT('h80)
	) name10803 (
		\wishbone_bd_ram_mem1_reg[209][8]/P0001 ,
		_w11977_,
		_w11984_,
		_w21316_
	);
	LUT3 #(
		.INIT('h80)
	) name10804 (
		\wishbone_bd_ram_mem1_reg[245][8]/P0001 ,
		_w11933_,
		_w11952_,
		_w21317_
	);
	LUT3 #(
		.INIT('h80)
	) name10805 (
		\wishbone_bd_ram_mem1_reg[208][8]/P0001 ,
		_w11941_,
		_w11984_,
		_w21318_
	);
	LUT4 #(
		.INIT('h0001)
	) name10806 (
		_w21315_,
		_w21316_,
		_w21317_,
		_w21318_,
		_w21319_
	);
	LUT3 #(
		.INIT('h80)
	) name10807 (
		\wishbone_bd_ram_mem1_reg[146][8]/P0001 ,
		_w11959_,
		_w11963_,
		_w21320_
	);
	LUT3 #(
		.INIT('h80)
	) name10808 (
		\wishbone_bd_ram_mem1_reg[67][8]/P0001 ,
		_w11938_,
		_w11949_,
		_w21321_
	);
	LUT3 #(
		.INIT('h80)
	) name10809 (
		\wishbone_bd_ram_mem1_reg[183][8]/P0001 ,
		_w11942_,
		_w11975_,
		_w21322_
	);
	LUT3 #(
		.INIT('h80)
	) name10810 (
		\wishbone_bd_ram_mem1_reg[167][8]/P0001 ,
		_w11930_,
		_w11975_,
		_w21323_
	);
	LUT4 #(
		.INIT('h0001)
	) name10811 (
		_w21320_,
		_w21321_,
		_w21322_,
		_w21323_,
		_w21324_
	);
	LUT3 #(
		.INIT('h80)
	) name10812 (
		\wishbone_bd_ram_mem1_reg[38][8]/P0001 ,
		_w11957_,
		_w11986_,
		_w21325_
	);
	LUT3 #(
		.INIT('h80)
	) name10813 (
		\wishbone_bd_ram_mem1_reg[230][8]/P0001 ,
		_w11982_,
		_w11986_,
		_w21326_
	);
	LUT3 #(
		.INIT('h80)
	) name10814 (
		\wishbone_bd_ram_mem1_reg[124][8]/P0001 ,
		_w11954_,
		_w12012_,
		_w21327_
	);
	LUT3 #(
		.INIT('h80)
	) name10815 (
		\wishbone_bd_ram_mem1_reg[73][8]/P0001 ,
		_w11949_,
		_w11968_,
		_w21328_
	);
	LUT4 #(
		.INIT('h0001)
	) name10816 (
		_w21325_,
		_w21326_,
		_w21327_,
		_w21328_,
		_w21329_
	);
	LUT4 #(
		.INIT('h8000)
	) name10817 (
		_w21314_,
		_w21319_,
		_w21324_,
		_w21329_,
		_w21330_
	);
	LUT3 #(
		.INIT('h80)
	) name10818 (
		\wishbone_bd_ram_mem1_reg[246][8]/P0001 ,
		_w11952_,
		_w11986_,
		_w21331_
	);
	LUT3 #(
		.INIT('h80)
	) name10819 (
		\wishbone_bd_ram_mem1_reg[65][8]/P0001 ,
		_w11949_,
		_w11977_,
		_w21332_
	);
	LUT3 #(
		.INIT('h80)
	) name10820 (
		\wishbone_bd_ram_mem1_reg[64][8]/P0001 ,
		_w11941_,
		_w11949_,
		_w21333_
	);
	LUT3 #(
		.INIT('h80)
	) name10821 (
		\wishbone_bd_ram_mem1_reg[103][8]/P0001 ,
		_w11965_,
		_w11975_,
		_w21334_
	);
	LUT4 #(
		.INIT('h0001)
	) name10822 (
		_w21331_,
		_w21332_,
		_w21333_,
		_w21334_,
		_w21335_
	);
	LUT3 #(
		.INIT('h80)
	) name10823 (
		\wishbone_bd_ram_mem1_reg[250][8]/P0001 ,
		_w11944_,
		_w11952_,
		_w21336_
	);
	LUT3 #(
		.INIT('h80)
	) name10824 (
		\wishbone_bd_ram_mem1_reg[110][8]/P0001 ,
		_w11948_,
		_w11965_,
		_w21337_
	);
	LUT3 #(
		.INIT('h80)
	) name10825 (
		\wishbone_bd_ram_mem1_reg[222][8]/P0001 ,
		_w11948_,
		_w11984_,
		_w21338_
	);
	LUT3 #(
		.INIT('h80)
	) name10826 (
		\wishbone_bd_ram_mem1_reg[158][8]/P0001 ,
		_w11948_,
		_w11959_,
		_w21339_
	);
	LUT4 #(
		.INIT('h0001)
	) name10827 (
		_w21336_,
		_w21337_,
		_w21338_,
		_w21339_,
		_w21340_
	);
	LUT3 #(
		.INIT('h80)
	) name10828 (
		\wishbone_bd_ram_mem1_reg[149][8]/P0001 ,
		_w11933_,
		_w11959_,
		_w21341_
	);
	LUT3 #(
		.INIT('h80)
	) name10829 (
		\wishbone_bd_ram_mem1_reg[8][8]/P0001 ,
		_w11932_,
		_w11990_,
		_w21342_
	);
	LUT3 #(
		.INIT('h80)
	) name10830 (
		\wishbone_bd_ram_mem1_reg[11][8]/P0001 ,
		_w11932_,
		_w11936_,
		_w21343_
	);
	LUT3 #(
		.INIT('h80)
	) name10831 (
		\wishbone_bd_ram_mem1_reg[55][8]/P0001 ,
		_w11975_,
		_w11979_,
		_w21344_
	);
	LUT4 #(
		.INIT('h0001)
	) name10832 (
		_w21341_,
		_w21342_,
		_w21343_,
		_w21344_,
		_w21345_
	);
	LUT3 #(
		.INIT('h80)
	) name10833 (
		\wishbone_bd_ram_mem1_reg[109][8]/P0001 ,
		_w11965_,
		_w11966_,
		_w21346_
	);
	LUT3 #(
		.INIT('h80)
	) name10834 (
		\wishbone_bd_ram_mem1_reg[219][8]/P0001 ,
		_w11936_,
		_w11984_,
		_w21347_
	);
	LUT3 #(
		.INIT('h80)
	) name10835 (
		\wishbone_bd_ram_mem1_reg[71][8]/P0001 ,
		_w11949_,
		_w11975_,
		_w21348_
	);
	LUT3 #(
		.INIT('h80)
	) name10836 (
		\wishbone_bd_ram_mem1_reg[54][8]/P0001 ,
		_w11979_,
		_w11986_,
		_w21349_
	);
	LUT4 #(
		.INIT('h0001)
	) name10837 (
		_w21346_,
		_w21347_,
		_w21348_,
		_w21349_,
		_w21350_
	);
	LUT4 #(
		.INIT('h8000)
	) name10838 (
		_w21335_,
		_w21340_,
		_w21345_,
		_w21350_,
		_w21351_
	);
	LUT3 #(
		.INIT('h80)
	) name10839 (
		\wishbone_bd_ram_mem1_reg[225][8]/P0001 ,
		_w11977_,
		_w11982_,
		_w21352_
	);
	LUT3 #(
		.INIT('h80)
	) name10840 (
		\wishbone_bd_ram_mem1_reg[7][8]/P0001 ,
		_w11932_,
		_w11975_,
		_w21353_
	);
	LUT3 #(
		.INIT('h80)
	) name10841 (
		\wishbone_bd_ram_mem1_reg[9][8]/P0001 ,
		_w11932_,
		_w11968_,
		_w21354_
	);
	LUT3 #(
		.INIT('h80)
	) name10842 (
		\wishbone_bd_ram_mem1_reg[242][8]/P0001 ,
		_w11952_,
		_w11963_,
		_w21355_
	);
	LUT4 #(
		.INIT('h0001)
	) name10843 (
		_w21352_,
		_w21353_,
		_w21354_,
		_w21355_,
		_w21356_
	);
	LUT3 #(
		.INIT('h80)
	) name10844 (
		\wishbone_bd_ram_mem1_reg[207][8]/P0001 ,
		_w11945_,
		_w11973_,
		_w21357_
	);
	LUT3 #(
		.INIT('h80)
	) name10845 (
		\wishbone_bd_ram_mem1_reg[90][8]/P0001 ,
		_w11944_,
		_w11972_,
		_w21358_
	);
	LUT3 #(
		.INIT('h80)
	) name10846 (
		\wishbone_bd_ram_mem1_reg[150][8]/P0001 ,
		_w11959_,
		_w11986_,
		_w21359_
	);
	LUT3 #(
		.INIT('h80)
	) name10847 (
		\wishbone_bd_ram_mem1_reg[147][8]/P0001 ,
		_w11938_,
		_w11959_,
		_w21360_
	);
	LUT4 #(
		.INIT('h0001)
	) name10848 (
		_w21357_,
		_w21358_,
		_w21359_,
		_w21360_,
		_w21361_
	);
	LUT3 #(
		.INIT('h80)
	) name10849 (
		\wishbone_bd_ram_mem1_reg[52][8]/P0001 ,
		_w11929_,
		_w11979_,
		_w21362_
	);
	LUT3 #(
		.INIT('h80)
	) name10850 (
		\wishbone_bd_ram_mem1_reg[105][8]/P0001 ,
		_w11965_,
		_w11968_,
		_w21363_
	);
	LUT3 #(
		.INIT('h80)
	) name10851 (
		\wishbone_bd_ram_mem1_reg[79][8]/P0001 ,
		_w11949_,
		_w11973_,
		_w21364_
	);
	LUT3 #(
		.INIT('h80)
	) name10852 (
		\wishbone_bd_ram_mem1_reg[224][8]/P0001 ,
		_w11941_,
		_w11982_,
		_w21365_
	);
	LUT4 #(
		.INIT('h0001)
	) name10853 (
		_w21362_,
		_w21363_,
		_w21364_,
		_w21365_,
		_w21366_
	);
	LUT3 #(
		.INIT('h80)
	) name10854 (
		\wishbone_bd_ram_mem1_reg[61][8]/P0001 ,
		_w11966_,
		_w11979_,
		_w21367_
	);
	LUT3 #(
		.INIT('h80)
	) name10855 (
		\wishbone_bd_ram_mem1_reg[93][8]/P0001 ,
		_w11966_,
		_w11972_,
		_w21368_
	);
	LUT3 #(
		.INIT('h80)
	) name10856 (
		\wishbone_bd_ram_mem1_reg[83][8]/P0001 ,
		_w11938_,
		_w11972_,
		_w21369_
	);
	LUT3 #(
		.INIT('h80)
	) name10857 (
		\wishbone_bd_ram_mem1_reg[41][8]/P0001 ,
		_w11957_,
		_w11968_,
		_w21370_
	);
	LUT4 #(
		.INIT('h0001)
	) name10858 (
		_w21367_,
		_w21368_,
		_w21369_,
		_w21370_,
		_w21371_
	);
	LUT4 #(
		.INIT('h8000)
	) name10859 (
		_w21356_,
		_w21361_,
		_w21366_,
		_w21371_,
		_w21372_
	);
	LUT3 #(
		.INIT('h80)
	) name10860 (
		\wishbone_bd_ram_mem1_reg[197][8]/P0001 ,
		_w11933_,
		_w11945_,
		_w21373_
	);
	LUT3 #(
		.INIT('h80)
	) name10861 (
		\wishbone_bd_ram_mem1_reg[203][8]/P0001 ,
		_w11936_,
		_w11945_,
		_w21374_
	);
	LUT3 #(
		.INIT('h80)
	) name10862 (
		\wishbone_bd_ram_mem1_reg[116][8]/P0001 ,
		_w11929_,
		_w12012_,
		_w21375_
	);
	LUT3 #(
		.INIT('h80)
	) name10863 (
		\wishbone_bd_ram_mem1_reg[6][8]/P0001 ,
		_w11932_,
		_w11986_,
		_w21376_
	);
	LUT4 #(
		.INIT('h0001)
	) name10864 (
		_w21373_,
		_w21374_,
		_w21375_,
		_w21376_,
		_w21377_
	);
	LUT3 #(
		.INIT('h80)
	) name10865 (
		\wishbone_bd_ram_mem1_reg[130][8]/P0001 ,
		_w11955_,
		_w11963_,
		_w21378_
	);
	LUT3 #(
		.INIT('h80)
	) name10866 (
		\wishbone_bd_ram_mem1_reg[243][8]/P0001 ,
		_w11938_,
		_w11952_,
		_w21379_
	);
	LUT3 #(
		.INIT('h80)
	) name10867 (
		\wishbone_bd_ram_mem1_reg[227][8]/P0001 ,
		_w11938_,
		_w11982_,
		_w21380_
	);
	LUT3 #(
		.INIT('h80)
	) name10868 (
		\wishbone_bd_ram_mem1_reg[235][8]/P0001 ,
		_w11936_,
		_w11982_,
		_w21381_
	);
	LUT4 #(
		.INIT('h0001)
	) name10869 (
		_w21378_,
		_w21379_,
		_w21380_,
		_w21381_,
		_w21382_
	);
	LUT3 #(
		.INIT('h80)
	) name10870 (
		\wishbone_bd_ram_mem1_reg[238][8]/P0001 ,
		_w11948_,
		_w11982_,
		_w21383_
	);
	LUT3 #(
		.INIT('h80)
	) name10871 (
		\wishbone_bd_ram_mem1_reg[128][8]/P0001 ,
		_w11941_,
		_w11955_,
		_w21384_
	);
	LUT3 #(
		.INIT('h80)
	) name10872 (
		\wishbone_bd_ram_mem1_reg[214][8]/P0001 ,
		_w11984_,
		_w11986_,
		_w21385_
	);
	LUT3 #(
		.INIT('h80)
	) name10873 (
		\wishbone_bd_ram_mem1_reg[172][8]/P0001 ,
		_w11930_,
		_w11954_,
		_w21386_
	);
	LUT4 #(
		.INIT('h0001)
	) name10874 (
		_w21383_,
		_w21384_,
		_w21385_,
		_w21386_,
		_w21387_
	);
	LUT3 #(
		.INIT('h80)
	) name10875 (
		\wishbone_bd_ram_mem1_reg[15][8]/P0001 ,
		_w11932_,
		_w11973_,
		_w21388_
	);
	LUT3 #(
		.INIT('h80)
	) name10876 (
		\wishbone_bd_ram_mem1_reg[47][8]/P0001 ,
		_w11957_,
		_w11973_,
		_w21389_
	);
	LUT3 #(
		.INIT('h80)
	) name10877 (
		\wishbone_bd_ram_mem1_reg[114][8]/P0001 ,
		_w11963_,
		_w12012_,
		_w21390_
	);
	LUT3 #(
		.INIT('h80)
	) name10878 (
		\wishbone_bd_ram_mem1_reg[106][8]/P0001 ,
		_w11944_,
		_w11965_,
		_w21391_
	);
	LUT4 #(
		.INIT('h0001)
	) name10879 (
		_w21388_,
		_w21389_,
		_w21390_,
		_w21391_,
		_w21392_
	);
	LUT4 #(
		.INIT('h8000)
	) name10880 (
		_w21377_,
		_w21382_,
		_w21387_,
		_w21392_,
		_w21393_
	);
	LUT4 #(
		.INIT('h8000)
	) name10881 (
		_w21330_,
		_w21351_,
		_w21372_,
		_w21393_,
		_w21394_
	);
	LUT3 #(
		.INIT('h80)
	) name10882 (
		\wishbone_bd_ram_mem1_reg[34][8]/P0001 ,
		_w11957_,
		_w11963_,
		_w21395_
	);
	LUT3 #(
		.INIT('h80)
	) name10883 (
		\wishbone_bd_ram_mem1_reg[139][8]/P0001 ,
		_w11936_,
		_w11955_,
		_w21396_
	);
	LUT3 #(
		.INIT('h80)
	) name10884 (
		\wishbone_bd_ram_mem1_reg[45][8]/P0001 ,
		_w11957_,
		_w11966_,
		_w21397_
	);
	LUT3 #(
		.INIT('h80)
	) name10885 (
		\wishbone_bd_ram_mem1_reg[100][8]/P0001 ,
		_w11929_,
		_w11965_,
		_w21398_
	);
	LUT4 #(
		.INIT('h0001)
	) name10886 (
		_w21395_,
		_w21396_,
		_w21397_,
		_w21398_,
		_w21399_
	);
	LUT3 #(
		.INIT('h80)
	) name10887 (
		\wishbone_bd_ram_mem1_reg[102][8]/P0001 ,
		_w11965_,
		_w11986_,
		_w21400_
	);
	LUT3 #(
		.INIT('h80)
	) name10888 (
		\wishbone_bd_ram_mem1_reg[53][8]/P0001 ,
		_w11933_,
		_w11979_,
		_w21401_
	);
	LUT3 #(
		.INIT('h80)
	) name10889 (
		\wishbone_bd_ram_mem1_reg[80][8]/P0001 ,
		_w11941_,
		_w11972_,
		_w21402_
	);
	LUT3 #(
		.INIT('h80)
	) name10890 (
		\wishbone_bd_ram_mem1_reg[70][8]/P0001 ,
		_w11949_,
		_w11986_,
		_w21403_
	);
	LUT4 #(
		.INIT('h0001)
	) name10891 (
		_w21400_,
		_w21401_,
		_w21402_,
		_w21403_,
		_w21404_
	);
	LUT3 #(
		.INIT('h80)
	) name10892 (
		\wishbone_bd_ram_mem1_reg[142][8]/P0001 ,
		_w11948_,
		_w11955_,
		_w21405_
	);
	LUT3 #(
		.INIT('h80)
	) name10893 (
		\wishbone_bd_ram_mem1_reg[169][8]/P0001 ,
		_w11930_,
		_w11968_,
		_w21406_
	);
	LUT3 #(
		.INIT('h80)
	) name10894 (
		\wishbone_bd_ram_mem1_reg[74][8]/P0001 ,
		_w11944_,
		_w11949_,
		_w21407_
	);
	LUT3 #(
		.INIT('h80)
	) name10895 (
		\wishbone_bd_ram_mem1_reg[212][8]/P0001 ,
		_w11929_,
		_w11984_,
		_w21408_
	);
	LUT4 #(
		.INIT('h0001)
	) name10896 (
		_w21405_,
		_w21406_,
		_w21407_,
		_w21408_,
		_w21409_
	);
	LUT3 #(
		.INIT('h80)
	) name10897 (
		\wishbone_bd_ram_mem1_reg[14][8]/P0001 ,
		_w11932_,
		_w11948_,
		_w21410_
	);
	LUT3 #(
		.INIT('h80)
	) name10898 (
		\wishbone_bd_ram_mem1_reg[13][8]/P0001 ,
		_w11932_,
		_w11966_,
		_w21411_
	);
	LUT3 #(
		.INIT('h80)
	) name10899 (
		\wishbone_bd_ram_mem1_reg[216][8]/P0001 ,
		_w11984_,
		_w11990_,
		_w21412_
	);
	LUT3 #(
		.INIT('h80)
	) name10900 (
		\wishbone_bd_ram_mem1_reg[26][8]/P0001 ,
		_w11935_,
		_w11944_,
		_w21413_
	);
	LUT4 #(
		.INIT('h0001)
	) name10901 (
		_w21410_,
		_w21411_,
		_w21412_,
		_w21413_,
		_w21414_
	);
	LUT4 #(
		.INIT('h8000)
	) name10902 (
		_w21399_,
		_w21404_,
		_w21409_,
		_w21414_,
		_w21415_
	);
	LUT3 #(
		.INIT('h80)
	) name10903 (
		\wishbone_bd_ram_mem1_reg[77][8]/P0001 ,
		_w11949_,
		_w11966_,
		_w21416_
	);
	LUT3 #(
		.INIT('h80)
	) name10904 (
		\wishbone_bd_ram_mem1_reg[217][8]/P0001 ,
		_w11968_,
		_w11984_,
		_w21417_
	);
	LUT3 #(
		.INIT('h80)
	) name10905 (
		\wishbone_bd_ram_mem1_reg[20][8]/P0001 ,
		_w11929_,
		_w11935_,
		_w21418_
	);
	LUT3 #(
		.INIT('h80)
	) name10906 (
		\wishbone_bd_ram_mem1_reg[88][8]/P0001 ,
		_w11972_,
		_w11990_,
		_w21419_
	);
	LUT4 #(
		.INIT('h0001)
	) name10907 (
		_w21416_,
		_w21417_,
		_w21418_,
		_w21419_,
		_w21420_
	);
	LUT3 #(
		.INIT('h80)
	) name10908 (
		\wishbone_bd_ram_mem1_reg[39][8]/P0001 ,
		_w11957_,
		_w11975_,
		_w21421_
	);
	LUT3 #(
		.INIT('h80)
	) name10909 (
		\wishbone_bd_ram_mem1_reg[82][8]/P0001 ,
		_w11963_,
		_w11972_,
		_w21422_
	);
	LUT3 #(
		.INIT('h80)
	) name10910 (
		\wishbone_bd_ram_mem1_reg[22][8]/P0001 ,
		_w11935_,
		_w11986_,
		_w21423_
	);
	LUT3 #(
		.INIT('h80)
	) name10911 (
		\wishbone_bd_ram_mem1_reg[28][8]/P0001 ,
		_w11935_,
		_w11954_,
		_w21424_
	);
	LUT4 #(
		.INIT('h0001)
	) name10912 (
		_w21421_,
		_w21422_,
		_w21423_,
		_w21424_,
		_w21425_
	);
	LUT3 #(
		.INIT('h80)
	) name10913 (
		\wishbone_bd_ram_mem1_reg[199][8]/P0001 ,
		_w11945_,
		_w11975_,
		_w21426_
	);
	LUT3 #(
		.INIT('h80)
	) name10914 (
		\wishbone_bd_ram_mem1_reg[234][8]/P0001 ,
		_w11944_,
		_w11982_,
		_w21427_
	);
	LUT3 #(
		.INIT('h80)
	) name10915 (
		\wishbone_bd_ram_mem1_reg[154][8]/P0001 ,
		_w11944_,
		_w11959_,
		_w21428_
	);
	LUT3 #(
		.INIT('h80)
	) name10916 (
		\wishbone_bd_ram_mem1_reg[141][8]/P0001 ,
		_w11955_,
		_w11966_,
		_w21429_
	);
	LUT4 #(
		.INIT('h0001)
	) name10917 (
		_w21426_,
		_w21427_,
		_w21428_,
		_w21429_,
		_w21430_
	);
	LUT3 #(
		.INIT('h80)
	) name10918 (
		\wishbone_bd_ram_mem1_reg[69][8]/P0001 ,
		_w11933_,
		_w11949_,
		_w21431_
	);
	LUT3 #(
		.INIT('h80)
	) name10919 (
		\wishbone_bd_ram_mem1_reg[60][8]/P0001 ,
		_w11954_,
		_w11979_,
		_w21432_
	);
	LUT3 #(
		.INIT('h80)
	) name10920 (
		\wishbone_bd_ram_mem1_reg[233][8]/P0001 ,
		_w11968_,
		_w11982_,
		_w21433_
	);
	LUT3 #(
		.INIT('h80)
	) name10921 (
		\wishbone_bd_ram_mem1_reg[122][8]/P0001 ,
		_w11944_,
		_w12012_,
		_w21434_
	);
	LUT4 #(
		.INIT('h0001)
	) name10922 (
		_w21431_,
		_w21432_,
		_w21433_,
		_w21434_,
		_w21435_
	);
	LUT4 #(
		.INIT('h8000)
	) name10923 (
		_w21420_,
		_w21425_,
		_w21430_,
		_w21435_,
		_w21436_
	);
	LUT3 #(
		.INIT('h80)
	) name10924 (
		\wishbone_bd_ram_mem1_reg[179][8]/P0001 ,
		_w11938_,
		_w11942_,
		_w21437_
	);
	LUT3 #(
		.INIT('h80)
	) name10925 (
		\wishbone_bd_ram_mem1_reg[40][8]/P0001 ,
		_w11957_,
		_w11990_,
		_w21438_
	);
	LUT3 #(
		.INIT('h80)
	) name10926 (
		\wishbone_bd_ram_mem1_reg[244][8]/P0001 ,
		_w11929_,
		_w11952_,
		_w21439_
	);
	LUT3 #(
		.INIT('h80)
	) name10927 (
		\wishbone_bd_ram_mem1_reg[63][8]/P0001 ,
		_w11973_,
		_w11979_,
		_w21440_
	);
	LUT4 #(
		.INIT('h0001)
	) name10928 (
		_w21437_,
		_w21438_,
		_w21439_,
		_w21440_,
		_w21441_
	);
	LUT3 #(
		.INIT('h80)
	) name10929 (
		\wishbone_bd_ram_mem1_reg[192][8]/P0001 ,
		_w11941_,
		_w11945_,
		_w21442_
	);
	LUT3 #(
		.INIT('h80)
	) name10930 (
		\wishbone_bd_ram_mem1_reg[94][8]/P0001 ,
		_w11948_,
		_w11972_,
		_w21443_
	);
	LUT3 #(
		.INIT('h80)
	) name10931 (
		\wishbone_bd_ram_mem1_reg[248][8]/P0001 ,
		_w11952_,
		_w11990_,
		_w21444_
	);
	LUT3 #(
		.INIT('h80)
	) name10932 (
		\wishbone_bd_ram_mem1_reg[175][8]/P0001 ,
		_w11930_,
		_w11973_,
		_w21445_
	);
	LUT4 #(
		.INIT('h0001)
	) name10933 (
		_w21442_,
		_w21443_,
		_w21444_,
		_w21445_,
		_w21446_
	);
	LUT3 #(
		.INIT('h80)
	) name10934 (
		\wishbone_bd_ram_mem1_reg[0][8]/P0001 ,
		_w11932_,
		_w11941_,
		_w21447_
	);
	LUT3 #(
		.INIT('h80)
	) name10935 (
		\wishbone_bd_ram_mem1_reg[23][8]/P0001 ,
		_w11935_,
		_w11975_,
		_w21448_
	);
	LUT3 #(
		.INIT('h80)
	) name10936 (
		\wishbone_bd_ram_mem1_reg[37][8]/P0001 ,
		_w11933_,
		_w11957_,
		_w21449_
	);
	LUT3 #(
		.INIT('h80)
	) name10937 (
		\wishbone_bd_ram_mem1_reg[112][8]/P0001 ,
		_w11941_,
		_w12012_,
		_w21450_
	);
	LUT4 #(
		.INIT('h0001)
	) name10938 (
		_w21447_,
		_w21448_,
		_w21449_,
		_w21450_,
		_w21451_
	);
	LUT3 #(
		.INIT('h80)
	) name10939 (
		\wishbone_bd_ram_mem1_reg[194][8]/P0001 ,
		_w11945_,
		_w11963_,
		_w21452_
	);
	LUT3 #(
		.INIT('h80)
	) name10940 (
		\wishbone_bd_ram_mem1_reg[153][8]/P0001 ,
		_w11959_,
		_w11968_,
		_w21453_
	);
	LUT3 #(
		.INIT('h80)
	) name10941 (
		\wishbone_bd_ram_mem1_reg[206][8]/P0001 ,
		_w11945_,
		_w11948_,
		_w21454_
	);
	LUT3 #(
		.INIT('h80)
	) name10942 (
		\wishbone_bd_ram_mem1_reg[17][8]/P0001 ,
		_w11935_,
		_w11977_,
		_w21455_
	);
	LUT4 #(
		.INIT('h0001)
	) name10943 (
		_w21452_,
		_w21453_,
		_w21454_,
		_w21455_,
		_w21456_
	);
	LUT4 #(
		.INIT('h8000)
	) name10944 (
		_w21441_,
		_w21446_,
		_w21451_,
		_w21456_,
		_w21457_
	);
	LUT3 #(
		.INIT('h80)
	) name10945 (
		\wishbone_bd_ram_mem1_reg[182][8]/P0001 ,
		_w11942_,
		_w11986_,
		_w21458_
	);
	LUT3 #(
		.INIT('h80)
	) name10946 (
		\wishbone_bd_ram_mem1_reg[136][8]/P0001 ,
		_w11955_,
		_w11990_,
		_w21459_
	);
	LUT3 #(
		.INIT('h80)
	) name10947 (
		\wishbone_bd_ram_mem1_reg[195][8]/P0001 ,
		_w11938_,
		_w11945_,
		_w21460_
	);
	LUT3 #(
		.INIT('h80)
	) name10948 (
		\wishbone_bd_ram_mem1_reg[108][8]/P0001 ,
		_w11954_,
		_w11965_,
		_w21461_
	);
	LUT4 #(
		.INIT('h0001)
	) name10949 (
		_w21458_,
		_w21459_,
		_w21460_,
		_w21461_,
		_w21462_
	);
	LUT3 #(
		.INIT('h80)
	) name10950 (
		\wishbone_bd_ram_mem1_reg[12][8]/P0001 ,
		_w11932_,
		_w11954_,
		_w21463_
	);
	LUT3 #(
		.INIT('h80)
	) name10951 (
		\wishbone_bd_ram_mem1_reg[62][8]/P0001 ,
		_w11948_,
		_w11979_,
		_w21464_
	);
	LUT3 #(
		.INIT('h80)
	) name10952 (
		\wishbone_bd_ram_mem1_reg[155][8]/P0001 ,
		_w11936_,
		_w11959_,
		_w21465_
	);
	LUT3 #(
		.INIT('h80)
	) name10953 (
		\wishbone_bd_ram_mem1_reg[247][8]/P0001 ,
		_w11952_,
		_w11975_,
		_w21466_
	);
	LUT4 #(
		.INIT('h0001)
	) name10954 (
		_w21463_,
		_w21464_,
		_w21465_,
		_w21466_,
		_w21467_
	);
	LUT3 #(
		.INIT('h80)
	) name10955 (
		\wishbone_bd_ram_mem1_reg[76][8]/P0001 ,
		_w11949_,
		_w11954_,
		_w21468_
	);
	LUT3 #(
		.INIT('h80)
	) name10956 (
		\wishbone_bd_ram_mem1_reg[87][8]/P0001 ,
		_w11972_,
		_w11975_,
		_w21469_
	);
	LUT3 #(
		.INIT('h80)
	) name10957 (
		\wishbone_bd_ram_mem1_reg[132][8]/P0001 ,
		_w11929_,
		_w11955_,
		_w21470_
	);
	LUT3 #(
		.INIT('h80)
	) name10958 (
		\wishbone_bd_ram_mem1_reg[196][8]/P0001 ,
		_w11929_,
		_w11945_,
		_w21471_
	);
	LUT4 #(
		.INIT('h0001)
	) name10959 (
		_w21468_,
		_w21469_,
		_w21470_,
		_w21471_,
		_w21472_
	);
	LUT3 #(
		.INIT('h80)
	) name10960 (
		\wishbone_bd_ram_mem1_reg[134][8]/P0001 ,
		_w11955_,
		_w11986_,
		_w21473_
	);
	LUT3 #(
		.INIT('h80)
	) name10961 (
		\wishbone_bd_ram_mem1_reg[176][8]/P0001 ,
		_w11941_,
		_w11942_,
		_w21474_
	);
	LUT3 #(
		.INIT('h80)
	) name10962 (
		\wishbone_bd_ram_mem1_reg[24][8]/P0001 ,
		_w11935_,
		_w11990_,
		_w21475_
	);
	LUT3 #(
		.INIT('h80)
	) name10963 (
		\wishbone_bd_ram_mem1_reg[220][8]/P0001 ,
		_w11954_,
		_w11984_,
		_w21476_
	);
	LUT4 #(
		.INIT('h0001)
	) name10964 (
		_w21473_,
		_w21474_,
		_w21475_,
		_w21476_,
		_w21477_
	);
	LUT4 #(
		.INIT('h8000)
	) name10965 (
		_w21462_,
		_w21467_,
		_w21472_,
		_w21477_,
		_w21478_
	);
	LUT4 #(
		.INIT('h8000)
	) name10966 (
		_w21415_,
		_w21436_,
		_w21457_,
		_w21478_,
		_w21479_
	);
	LUT4 #(
		.INIT('h8000)
	) name10967 (
		_w21224_,
		_w21309_,
		_w21394_,
		_w21479_,
		_w21480_
	);
	LUT4 #(
		.INIT('h1555)
	) name10968 (
		wb_rst_i_pad,
		_w21126_,
		_w21130_,
		_w21138_,
		_w21481_
	);
	LUT3 #(
		.INIT('hba)
	) name10969 (
		_w21139_,
		_w21480_,
		_w21481_,
		_w21482_
	);
	LUT4 #(
		.INIT('h0002)
	) name10970 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21483_
	);
	LUT3 #(
		.INIT('h80)
	) name10971 (
		_w18757_,
		_w18762_,
		_w21483_,
		_w21484_
	);
	LUT3 #(
		.INIT('h80)
	) name10972 (
		\ethreg1_MIIRX_DATA_DataOut_reg[9]/NET0131 ,
		_w18785_,
		_w18786_,
		_w21485_
	);
	LUT4 #(
		.INIT('h0008)
	) name10973 (
		\ethreg1_RXHASH0_1_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21486_
	);
	LUT3 #(
		.INIT('h80)
	) name10974 (
		_w18757_,
		_w18758_,
		_w21486_,
		_w21487_
	);
	LUT4 #(
		.INIT('h0008)
	) name10975 (
		\ethreg1_RXHASH1_1_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21488_
	);
	LUT3 #(
		.INIT('h80)
	) name10976 (
		_w18757_,
		_w18762_,
		_w21488_,
		_w21489_
	);
	LUT4 #(
		.INIT('h0001)
	) name10977 (
		_w21484_,
		_w21485_,
		_w21487_,
		_w21489_,
		_w21490_
	);
	LUT4 #(
		.INIT('h0002)
	) name10978 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21491_
	);
	LUT4 #(
		.INIT('h0020)
	) name10979 (
		\ethreg1_TXCTRL_1_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21492_
	);
	LUT4 #(
		.INIT('h777f)
	) name10980 (
		_w18757_,
		_w18758_,
		_w21491_,
		_w21492_,
		_w21493_
	);
	LUT2 #(
		.INIT('h8)
	) name10981 (
		_w18752_,
		_w21493_,
		_w21494_
	);
	LUT3 #(
		.INIT('h80)
	) name10982 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[1]/NET0131 ,
		_w18785_,
		_w18798_,
		_w21495_
	);
	LUT3 #(
		.INIT('h80)
	) name10983 (
		\ethreg1_MODER_1_DataOut_reg[1]/NET0131 ,
		_w18800_,
		_w18801_,
		_w21496_
	);
	LUT3 #(
		.INIT('h80)
	) name10984 (
		\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 ,
		_w18753_,
		_w18754_,
		_w21497_
	);
	LUT3 #(
		.INIT('h80)
	) name10985 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[1]/NET0131 ,
		_w18798_,
		_w18805_,
		_w21498_
	);
	LUT4 #(
		.INIT('h0001)
	) name10986 (
		_w21495_,
		_w21496_,
		_w21497_,
		_w21498_,
		_w21499_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10987 (
		_w18752_,
		_w21490_,
		_w21493_,
		_w21499_,
		_w21500_
	);
	LUT3 #(
		.INIT('h80)
	) name10988 (
		\wishbone_bd_ram_mem1_reg[39][9]/P0001 ,
		_w11957_,
		_w11975_,
		_w21501_
	);
	LUT3 #(
		.INIT('h80)
	) name10989 (
		\wishbone_bd_ram_mem1_reg[109][9]/P0001 ,
		_w11965_,
		_w11966_,
		_w21502_
	);
	LUT3 #(
		.INIT('h80)
	) name10990 (
		\wishbone_bd_ram_mem1_reg[82][9]/P0001 ,
		_w11963_,
		_w11972_,
		_w21503_
	);
	LUT3 #(
		.INIT('h80)
	) name10991 (
		\wishbone_bd_ram_mem1_reg[32][9]/P0001 ,
		_w11941_,
		_w11957_,
		_w21504_
	);
	LUT4 #(
		.INIT('h0001)
	) name10992 (
		_w21501_,
		_w21502_,
		_w21503_,
		_w21504_,
		_w21505_
	);
	LUT3 #(
		.INIT('h80)
	) name10993 (
		\wishbone_bd_ram_mem1_reg[48][9]/P0001 ,
		_w11941_,
		_w11979_,
		_w21506_
	);
	LUT3 #(
		.INIT('h80)
	) name10994 (
		\wishbone_bd_ram_mem1_reg[241][9]/P0001 ,
		_w11952_,
		_w11977_,
		_w21507_
	);
	LUT3 #(
		.INIT('h80)
	) name10995 (
		\wishbone_bd_ram_mem1_reg[57][9]/P0001 ,
		_w11968_,
		_w11979_,
		_w21508_
	);
	LUT3 #(
		.INIT('h80)
	) name10996 (
		\wishbone_bd_ram_mem1_reg[209][9]/P0001 ,
		_w11977_,
		_w11984_,
		_w21509_
	);
	LUT4 #(
		.INIT('h0001)
	) name10997 (
		_w21506_,
		_w21507_,
		_w21508_,
		_w21509_,
		_w21510_
	);
	LUT3 #(
		.INIT('h80)
	) name10998 (
		\wishbone_bd_ram_mem1_reg[178][9]/P0001 ,
		_w11942_,
		_w11963_,
		_w21511_
	);
	LUT3 #(
		.INIT('h80)
	) name10999 (
		\wishbone_bd_ram_mem1_reg[244][9]/P0001 ,
		_w11929_,
		_w11952_,
		_w21512_
	);
	LUT3 #(
		.INIT('h80)
	) name11000 (
		\wishbone_bd_ram_mem1_reg[160][9]/P0001 ,
		_w11930_,
		_w11941_,
		_w21513_
	);
	LUT3 #(
		.INIT('h80)
	) name11001 (
		\wishbone_bd_ram_mem1_reg[133][9]/P0001 ,
		_w11933_,
		_w11955_,
		_w21514_
	);
	LUT4 #(
		.INIT('h0001)
	) name11002 (
		_w21511_,
		_w21512_,
		_w21513_,
		_w21514_,
		_w21515_
	);
	LUT3 #(
		.INIT('h80)
	) name11003 (
		\wishbone_bd_ram_mem1_reg[7][9]/P0001 ,
		_w11932_,
		_w11975_,
		_w21516_
	);
	LUT3 #(
		.INIT('h80)
	) name11004 (
		\wishbone_bd_ram_mem1_reg[238][9]/P0001 ,
		_w11948_,
		_w11982_,
		_w21517_
	);
	LUT3 #(
		.INIT('h80)
	) name11005 (
		\wishbone_bd_ram_mem1_reg[36][9]/P0001 ,
		_w11929_,
		_w11957_,
		_w21518_
	);
	LUT3 #(
		.INIT('h80)
	) name11006 (
		\wishbone_bd_ram_mem1_reg[251][9]/P0001 ,
		_w11936_,
		_w11952_,
		_w21519_
	);
	LUT4 #(
		.INIT('h0001)
	) name11007 (
		_w21516_,
		_w21517_,
		_w21518_,
		_w21519_,
		_w21520_
	);
	LUT4 #(
		.INIT('h8000)
	) name11008 (
		_w21505_,
		_w21510_,
		_w21515_,
		_w21520_,
		_w21521_
	);
	LUT3 #(
		.INIT('h80)
	) name11009 (
		\wishbone_bd_ram_mem1_reg[107][9]/P0001 ,
		_w11936_,
		_w11965_,
		_w21522_
	);
	LUT3 #(
		.INIT('h80)
	) name11010 (
		\wishbone_bd_ram_mem1_reg[174][9]/P0001 ,
		_w11930_,
		_w11948_,
		_w21523_
	);
	LUT3 #(
		.INIT('h80)
	) name11011 (
		\wishbone_bd_ram_mem1_reg[1][9]/P0001 ,
		_w11932_,
		_w11977_,
		_w21524_
	);
	LUT3 #(
		.INIT('h80)
	) name11012 (
		\wishbone_bd_ram_mem1_reg[142][9]/P0001 ,
		_w11948_,
		_w11955_,
		_w21525_
	);
	LUT4 #(
		.INIT('h0001)
	) name11013 (
		_w21522_,
		_w21523_,
		_w21524_,
		_w21525_,
		_w21526_
	);
	LUT3 #(
		.INIT('h80)
	) name11014 (
		\wishbone_bd_ram_mem1_reg[194][9]/P0001 ,
		_w11945_,
		_w11963_,
		_w21527_
	);
	LUT3 #(
		.INIT('h80)
	) name11015 (
		\wishbone_bd_ram_mem1_reg[224][9]/P0001 ,
		_w11941_,
		_w11982_,
		_w21528_
	);
	LUT3 #(
		.INIT('h80)
	) name11016 (
		\wishbone_bd_ram_mem1_reg[185][9]/P0001 ,
		_w11942_,
		_w11968_,
		_w21529_
	);
	LUT3 #(
		.INIT('h80)
	) name11017 (
		\wishbone_bd_ram_mem1_reg[27][9]/P0001 ,
		_w11935_,
		_w11936_,
		_w21530_
	);
	LUT4 #(
		.INIT('h0001)
	) name11018 (
		_w21527_,
		_w21528_,
		_w21529_,
		_w21530_,
		_w21531_
	);
	LUT3 #(
		.INIT('h80)
	) name11019 (
		\wishbone_bd_ram_mem1_reg[95][9]/P0001 ,
		_w11972_,
		_w11973_,
		_w21532_
	);
	LUT3 #(
		.INIT('h80)
	) name11020 (
		\wishbone_bd_ram_mem1_reg[249][9]/P0001 ,
		_w11952_,
		_w11968_,
		_w21533_
	);
	LUT3 #(
		.INIT('h80)
	) name11021 (
		\wishbone_bd_ram_mem1_reg[201][9]/P0001 ,
		_w11945_,
		_w11968_,
		_w21534_
	);
	LUT3 #(
		.INIT('h80)
	) name11022 (
		\wishbone_bd_ram_mem1_reg[40][9]/P0001 ,
		_w11957_,
		_w11990_,
		_w21535_
	);
	LUT4 #(
		.INIT('h0001)
	) name11023 (
		_w21532_,
		_w21533_,
		_w21534_,
		_w21535_,
		_w21536_
	);
	LUT3 #(
		.INIT('h80)
	) name11024 (
		\wishbone_bd_ram_mem1_reg[52][9]/P0001 ,
		_w11929_,
		_w11979_,
		_w21537_
	);
	LUT3 #(
		.INIT('h80)
	) name11025 (
		\wishbone_bd_ram_mem1_reg[126][9]/P0001 ,
		_w11948_,
		_w12012_,
		_w21538_
	);
	LUT3 #(
		.INIT('h80)
	) name11026 (
		\wishbone_bd_ram_mem1_reg[171][9]/P0001 ,
		_w11930_,
		_w11936_,
		_w21539_
	);
	LUT3 #(
		.INIT('h80)
	) name11027 (
		\wishbone_bd_ram_mem1_reg[250][9]/P0001 ,
		_w11944_,
		_w11952_,
		_w21540_
	);
	LUT4 #(
		.INIT('h0001)
	) name11028 (
		_w21537_,
		_w21538_,
		_w21539_,
		_w21540_,
		_w21541_
	);
	LUT4 #(
		.INIT('h8000)
	) name11029 (
		_w21526_,
		_w21531_,
		_w21536_,
		_w21541_,
		_w21542_
	);
	LUT3 #(
		.INIT('h80)
	) name11030 (
		\wishbone_bd_ram_mem1_reg[223][9]/P0001 ,
		_w11973_,
		_w11984_,
		_w21543_
	);
	LUT3 #(
		.INIT('h80)
	) name11031 (
		\wishbone_bd_ram_mem1_reg[87][9]/P0001 ,
		_w11972_,
		_w11975_,
		_w21544_
	);
	LUT3 #(
		.INIT('h80)
	) name11032 (
		\wishbone_bd_ram_mem1_reg[97][9]/P0001 ,
		_w11965_,
		_w11977_,
		_w21545_
	);
	LUT3 #(
		.INIT('h80)
	) name11033 (
		\wishbone_bd_ram_mem1_reg[4][9]/P0001 ,
		_w11929_,
		_w11932_,
		_w21546_
	);
	LUT4 #(
		.INIT('h0001)
	) name11034 (
		_w21543_,
		_w21544_,
		_w21545_,
		_w21546_,
		_w21547_
	);
	LUT3 #(
		.INIT('h80)
	) name11035 (
		\wishbone_bd_ram_mem1_reg[197][9]/P0001 ,
		_w11933_,
		_w11945_,
		_w21548_
	);
	LUT3 #(
		.INIT('h80)
	) name11036 (
		\wishbone_bd_ram_mem1_reg[64][9]/P0001 ,
		_w11941_,
		_w11949_,
		_w21549_
	);
	LUT3 #(
		.INIT('h80)
	) name11037 (
		\wishbone_bd_ram_mem1_reg[206][9]/P0001 ,
		_w11945_,
		_w11948_,
		_w21550_
	);
	LUT3 #(
		.INIT('h80)
	) name11038 (
		\wishbone_bd_ram_mem1_reg[102][9]/P0001 ,
		_w11965_,
		_w11986_,
		_w21551_
	);
	LUT4 #(
		.INIT('h0001)
	) name11039 (
		_w21548_,
		_w21549_,
		_w21550_,
		_w21551_,
		_w21552_
	);
	LUT3 #(
		.INIT('h80)
	) name11040 (
		\wishbone_bd_ram_mem1_reg[189][9]/P0001 ,
		_w11942_,
		_w11966_,
		_w21553_
	);
	LUT3 #(
		.INIT('h80)
	) name11041 (
		\wishbone_bd_ram_mem1_reg[181][9]/P0001 ,
		_w11933_,
		_w11942_,
		_w21554_
	);
	LUT3 #(
		.INIT('h80)
	) name11042 (
		\wishbone_bd_ram_mem1_reg[129][9]/P0001 ,
		_w11955_,
		_w11977_,
		_w21555_
	);
	LUT3 #(
		.INIT('h80)
	) name11043 (
		\wishbone_bd_ram_mem1_reg[235][9]/P0001 ,
		_w11936_,
		_w11982_,
		_w21556_
	);
	LUT4 #(
		.INIT('h0001)
	) name11044 (
		_w21553_,
		_w21554_,
		_w21555_,
		_w21556_,
		_w21557_
	);
	LUT3 #(
		.INIT('h80)
	) name11045 (
		\wishbone_bd_ram_mem1_reg[202][9]/P0001 ,
		_w11944_,
		_w11945_,
		_w21558_
	);
	LUT3 #(
		.INIT('h80)
	) name11046 (
		\wishbone_bd_ram_mem1_reg[217][9]/P0001 ,
		_w11968_,
		_w11984_,
		_w21559_
	);
	LUT3 #(
		.INIT('h80)
	) name11047 (
		\wishbone_bd_ram_mem1_reg[157][9]/P0001 ,
		_w11959_,
		_w11966_,
		_w21560_
	);
	LUT3 #(
		.INIT('h80)
	) name11048 (
		\wishbone_bd_ram_mem1_reg[215][9]/P0001 ,
		_w11975_,
		_w11984_,
		_w21561_
	);
	LUT4 #(
		.INIT('h0001)
	) name11049 (
		_w21558_,
		_w21559_,
		_w21560_,
		_w21561_,
		_w21562_
	);
	LUT4 #(
		.INIT('h8000)
	) name11050 (
		_w21547_,
		_w21552_,
		_w21557_,
		_w21562_,
		_w21563_
	);
	LUT3 #(
		.INIT('h80)
	) name11051 (
		\wishbone_bd_ram_mem1_reg[134][9]/P0001 ,
		_w11955_,
		_w11986_,
		_w21564_
	);
	LUT3 #(
		.INIT('h80)
	) name11052 (
		\wishbone_bd_ram_mem1_reg[170][9]/P0001 ,
		_w11930_,
		_w11944_,
		_w21565_
	);
	LUT3 #(
		.INIT('h80)
	) name11053 (
		\wishbone_bd_ram_mem1_reg[45][9]/P0001 ,
		_w11957_,
		_w11966_,
		_w21566_
	);
	LUT3 #(
		.INIT('h80)
	) name11054 (
		\wishbone_bd_ram_mem1_reg[120][9]/P0001 ,
		_w11990_,
		_w12012_,
		_w21567_
	);
	LUT4 #(
		.INIT('h0001)
	) name11055 (
		_w21564_,
		_w21565_,
		_w21566_,
		_w21567_,
		_w21568_
	);
	LUT3 #(
		.INIT('h80)
	) name11056 (
		\wishbone_bd_ram_mem1_reg[42][9]/P0001 ,
		_w11944_,
		_w11957_,
		_w21569_
	);
	LUT3 #(
		.INIT('h80)
	) name11057 (
		\wishbone_bd_ram_mem1_reg[208][9]/P0001 ,
		_w11941_,
		_w11984_,
		_w21570_
	);
	LUT3 #(
		.INIT('h80)
	) name11058 (
		\wishbone_bd_ram_mem1_reg[85][9]/P0001 ,
		_w11933_,
		_w11972_,
		_w21571_
	);
	LUT3 #(
		.INIT('h80)
	) name11059 (
		\wishbone_bd_ram_mem1_reg[17][9]/P0001 ,
		_w11935_,
		_w11977_,
		_w21572_
	);
	LUT4 #(
		.INIT('h0001)
	) name11060 (
		_w21569_,
		_w21570_,
		_w21571_,
		_w21572_,
		_w21573_
	);
	LUT3 #(
		.INIT('h80)
	) name11061 (
		\wishbone_bd_ram_mem1_reg[132][9]/P0001 ,
		_w11929_,
		_w11955_,
		_w21574_
	);
	LUT3 #(
		.INIT('h80)
	) name11062 (
		\wishbone_bd_ram_mem1_reg[86][9]/P0001 ,
		_w11972_,
		_w11986_,
		_w21575_
	);
	LUT3 #(
		.INIT('h80)
	) name11063 (
		\wishbone_bd_ram_mem1_reg[117][9]/P0001 ,
		_w11933_,
		_w12012_,
		_w21576_
	);
	LUT3 #(
		.INIT('h80)
	) name11064 (
		\wishbone_bd_ram_mem1_reg[56][9]/P0001 ,
		_w11979_,
		_w11990_,
		_w21577_
	);
	LUT4 #(
		.INIT('h0001)
	) name11065 (
		_w21574_,
		_w21575_,
		_w21576_,
		_w21577_,
		_w21578_
	);
	LUT3 #(
		.INIT('h80)
	) name11066 (
		\wishbone_bd_ram_mem1_reg[10][9]/P0001 ,
		_w11932_,
		_w11944_,
		_w21579_
	);
	LUT3 #(
		.INIT('h80)
	) name11067 (
		\wishbone_bd_ram_mem1_reg[83][9]/P0001 ,
		_w11938_,
		_w11972_,
		_w21580_
	);
	LUT3 #(
		.INIT('h80)
	) name11068 (
		\wishbone_bd_ram_mem1_reg[21][9]/P0001 ,
		_w11933_,
		_w11935_,
		_w21581_
	);
	LUT3 #(
		.INIT('h80)
	) name11069 (
		\wishbone_bd_ram_mem1_reg[156][9]/P0001 ,
		_w11954_,
		_w11959_,
		_w21582_
	);
	LUT4 #(
		.INIT('h0001)
	) name11070 (
		_w21579_,
		_w21580_,
		_w21581_,
		_w21582_,
		_w21583_
	);
	LUT4 #(
		.INIT('h8000)
	) name11071 (
		_w21568_,
		_w21573_,
		_w21578_,
		_w21583_,
		_w21584_
	);
	LUT4 #(
		.INIT('h8000)
	) name11072 (
		_w21521_,
		_w21542_,
		_w21563_,
		_w21584_,
		_w21585_
	);
	LUT3 #(
		.INIT('h80)
	) name11073 (
		\wishbone_bd_ram_mem1_reg[73][9]/P0001 ,
		_w11949_,
		_w11968_,
		_w21586_
	);
	LUT3 #(
		.INIT('h80)
	) name11074 (
		\wishbone_bd_ram_mem1_reg[186][9]/P0001 ,
		_w11942_,
		_w11944_,
		_w21587_
	);
	LUT3 #(
		.INIT('h80)
	) name11075 (
		\wishbone_bd_ram_mem1_reg[236][9]/P0001 ,
		_w11954_,
		_w11982_,
		_w21588_
	);
	LUT3 #(
		.INIT('h80)
	) name11076 (
		\wishbone_bd_ram_mem1_reg[130][9]/P0001 ,
		_w11955_,
		_w11963_,
		_w21589_
	);
	LUT4 #(
		.INIT('h0001)
	) name11077 (
		_w21586_,
		_w21587_,
		_w21588_,
		_w21589_,
		_w21590_
	);
	LUT3 #(
		.INIT('h80)
	) name11078 (
		\wishbone_bd_ram_mem1_reg[68][9]/P0001 ,
		_w11929_,
		_w11949_,
		_w21591_
	);
	LUT3 #(
		.INIT('h80)
	) name11079 (
		\wishbone_bd_ram_mem1_reg[195][9]/P0001 ,
		_w11938_,
		_w11945_,
		_w21592_
	);
	LUT3 #(
		.INIT('h80)
	) name11080 (
		\wishbone_bd_ram_mem1_reg[166][9]/P0001 ,
		_w11930_,
		_w11986_,
		_w21593_
	);
	LUT3 #(
		.INIT('h80)
	) name11081 (
		\wishbone_bd_ram_mem1_reg[106][9]/P0001 ,
		_w11944_,
		_w11965_,
		_w21594_
	);
	LUT4 #(
		.INIT('h0001)
	) name11082 (
		_w21591_,
		_w21592_,
		_w21593_,
		_w21594_,
		_w21595_
	);
	LUT3 #(
		.INIT('h80)
	) name11083 (
		\wishbone_bd_ram_mem1_reg[139][9]/P0001 ,
		_w11936_,
		_w11955_,
		_w21596_
	);
	LUT3 #(
		.INIT('h80)
	) name11084 (
		\wishbone_bd_ram_mem1_reg[123][9]/P0001 ,
		_w11936_,
		_w12012_,
		_w21597_
	);
	LUT3 #(
		.INIT('h80)
	) name11085 (
		\wishbone_bd_ram_mem1_reg[196][9]/P0001 ,
		_w11929_,
		_w11945_,
		_w21598_
	);
	LUT3 #(
		.INIT('h80)
	) name11086 (
		\wishbone_bd_ram_mem1_reg[204][9]/P0001 ,
		_w11945_,
		_w11954_,
		_w21599_
	);
	LUT4 #(
		.INIT('h0001)
	) name11087 (
		_w21596_,
		_w21597_,
		_w21598_,
		_w21599_,
		_w21600_
	);
	LUT3 #(
		.INIT('h80)
	) name11088 (
		\wishbone_bd_ram_mem1_reg[193][9]/P0001 ,
		_w11945_,
		_w11977_,
		_w21601_
	);
	LUT3 #(
		.INIT('h80)
	) name11089 (
		\wishbone_bd_ram_mem1_reg[149][9]/P0001 ,
		_w11933_,
		_w11959_,
		_w21602_
	);
	LUT3 #(
		.INIT('h80)
	) name11090 (
		\wishbone_bd_ram_mem1_reg[151][9]/P0001 ,
		_w11959_,
		_w11975_,
		_w21603_
	);
	LUT3 #(
		.INIT('h80)
	) name11091 (
		\wishbone_bd_ram_mem1_reg[154][9]/P0001 ,
		_w11944_,
		_w11959_,
		_w21604_
	);
	LUT4 #(
		.INIT('h0001)
	) name11092 (
		_w21601_,
		_w21602_,
		_w21603_,
		_w21604_,
		_w21605_
	);
	LUT4 #(
		.INIT('h8000)
	) name11093 (
		_w21590_,
		_w21595_,
		_w21600_,
		_w21605_,
		_w21606_
	);
	LUT3 #(
		.INIT('h80)
	) name11094 (
		\wishbone_bd_ram_mem1_reg[84][9]/P0001 ,
		_w11929_,
		_w11972_,
		_w21607_
	);
	LUT3 #(
		.INIT('h80)
	) name11095 (
		\wishbone_bd_ram_mem1_reg[173][9]/P0001 ,
		_w11930_,
		_w11966_,
		_w21608_
	);
	LUT3 #(
		.INIT('h80)
	) name11096 (
		\wishbone_bd_ram_mem1_reg[119][9]/P0001 ,
		_w11975_,
		_w12012_,
		_w21609_
	);
	LUT3 #(
		.INIT('h80)
	) name11097 (
		\wishbone_bd_ram_mem1_reg[25][9]/P0001 ,
		_w11935_,
		_w11968_,
		_w21610_
	);
	LUT4 #(
		.INIT('h0001)
	) name11098 (
		_w21607_,
		_w21608_,
		_w21609_,
		_w21610_,
		_w21611_
	);
	LUT3 #(
		.INIT('h80)
	) name11099 (
		\wishbone_bd_ram_mem1_reg[9][9]/P0001 ,
		_w11932_,
		_w11968_,
		_w21612_
	);
	LUT3 #(
		.INIT('h80)
	) name11100 (
		\wishbone_bd_ram_mem1_reg[20][9]/P0001 ,
		_w11929_,
		_w11935_,
		_w21613_
	);
	LUT3 #(
		.INIT('h80)
	) name11101 (
		\wishbone_bd_ram_mem1_reg[30][9]/P0001 ,
		_w11935_,
		_w11948_,
		_w21614_
	);
	LUT3 #(
		.INIT('h80)
	) name11102 (
		\wishbone_bd_ram_mem1_reg[144][9]/P0001 ,
		_w11941_,
		_w11959_,
		_w21615_
	);
	LUT4 #(
		.INIT('h0001)
	) name11103 (
		_w21612_,
		_w21613_,
		_w21614_,
		_w21615_,
		_w21616_
	);
	LUT3 #(
		.INIT('h80)
	) name11104 (
		\wishbone_bd_ram_mem1_reg[13][9]/P0001 ,
		_w11932_,
		_w11966_,
		_w21617_
	);
	LUT3 #(
		.INIT('h80)
	) name11105 (
		\wishbone_bd_ram_mem1_reg[111][9]/P0001 ,
		_w11965_,
		_w11973_,
		_w21618_
	);
	LUT3 #(
		.INIT('h80)
	) name11106 (
		\wishbone_bd_ram_mem1_reg[118][9]/P0001 ,
		_w11986_,
		_w12012_,
		_w21619_
	);
	LUT3 #(
		.INIT('h80)
	) name11107 (
		\wishbone_bd_ram_mem1_reg[22][9]/P0001 ,
		_w11935_,
		_w11986_,
		_w21620_
	);
	LUT4 #(
		.INIT('h0001)
	) name11108 (
		_w21617_,
		_w21618_,
		_w21619_,
		_w21620_,
		_w21621_
	);
	LUT3 #(
		.INIT('h80)
	) name11109 (
		\wishbone_bd_ram_mem1_reg[231][9]/P0001 ,
		_w11975_,
		_w11982_,
		_w21622_
	);
	LUT3 #(
		.INIT('h80)
	) name11110 (
		\wishbone_bd_ram_mem1_reg[254][9]/P0001 ,
		_w11948_,
		_w11952_,
		_w21623_
	);
	LUT3 #(
		.INIT('h80)
	) name11111 (
		\wishbone_bd_ram_mem1_reg[205][9]/P0001 ,
		_w11945_,
		_w11966_,
		_w21624_
	);
	LUT3 #(
		.INIT('h80)
	) name11112 (
		\wishbone_bd_ram_mem1_reg[138][9]/P0001 ,
		_w11944_,
		_w11955_,
		_w21625_
	);
	LUT4 #(
		.INIT('h0001)
	) name11113 (
		_w21622_,
		_w21623_,
		_w21624_,
		_w21625_,
		_w21626_
	);
	LUT4 #(
		.INIT('h8000)
	) name11114 (
		_w21611_,
		_w21616_,
		_w21621_,
		_w21626_,
		_w21627_
	);
	LUT3 #(
		.INIT('h80)
	) name11115 (
		\wishbone_bd_ram_mem1_reg[165][9]/P0001 ,
		_w11930_,
		_w11933_,
		_w21628_
	);
	LUT3 #(
		.INIT('h80)
	) name11116 (
		\wishbone_bd_ram_mem1_reg[237][9]/P0001 ,
		_w11966_,
		_w11982_,
		_w21629_
	);
	LUT3 #(
		.INIT('h80)
	) name11117 (
		\wishbone_bd_ram_mem1_reg[146][9]/P0001 ,
		_w11959_,
		_w11963_,
		_w21630_
	);
	LUT3 #(
		.INIT('h80)
	) name11118 (
		\wishbone_bd_ram_mem1_reg[127][9]/P0001 ,
		_w11973_,
		_w12012_,
		_w21631_
	);
	LUT4 #(
		.INIT('h0001)
	) name11119 (
		_w21628_,
		_w21629_,
		_w21630_,
		_w21631_,
		_w21632_
	);
	LUT3 #(
		.INIT('h80)
	) name11120 (
		\wishbone_bd_ram_mem1_reg[220][9]/P0001 ,
		_w11954_,
		_w11984_,
		_w21633_
	);
	LUT3 #(
		.INIT('h80)
	) name11121 (
		\wishbone_bd_ram_mem1_reg[246][9]/P0001 ,
		_w11952_,
		_w11986_,
		_w21634_
	);
	LUT3 #(
		.INIT('h80)
	) name11122 (
		\wishbone_bd_ram_mem1_reg[2][9]/P0001 ,
		_w11932_,
		_w11963_,
		_w21635_
	);
	LUT3 #(
		.INIT('h80)
	) name11123 (
		\wishbone_bd_ram_mem1_reg[77][9]/P0001 ,
		_w11949_,
		_w11966_,
		_w21636_
	);
	LUT4 #(
		.INIT('h0001)
	) name11124 (
		_w21633_,
		_w21634_,
		_w21635_,
		_w21636_,
		_w21637_
	);
	LUT3 #(
		.INIT('h80)
	) name11125 (
		\wishbone_bd_ram_mem1_reg[213][9]/P0001 ,
		_w11933_,
		_w11984_,
		_w21638_
	);
	LUT3 #(
		.INIT('h80)
	) name11126 (
		\wishbone_bd_ram_mem1_reg[34][9]/P0001 ,
		_w11957_,
		_w11963_,
		_w21639_
	);
	LUT3 #(
		.INIT('h80)
	) name11127 (
		\wishbone_bd_ram_mem1_reg[184][9]/P0001 ,
		_w11942_,
		_w11990_,
		_w21640_
	);
	LUT3 #(
		.INIT('h80)
	) name11128 (
		\wishbone_bd_ram_mem1_reg[54][9]/P0001 ,
		_w11979_,
		_w11986_,
		_w21641_
	);
	LUT4 #(
		.INIT('h0001)
	) name11129 (
		_w21638_,
		_w21639_,
		_w21640_,
		_w21641_,
		_w21642_
	);
	LUT3 #(
		.INIT('h80)
	) name11130 (
		\wishbone_bd_ram_mem1_reg[180][9]/P0001 ,
		_w11929_,
		_w11942_,
		_w21643_
	);
	LUT3 #(
		.INIT('h80)
	) name11131 (
		\wishbone_bd_ram_mem1_reg[252][9]/P0001 ,
		_w11952_,
		_w11954_,
		_w21644_
	);
	LUT3 #(
		.INIT('h80)
	) name11132 (
		\wishbone_bd_ram_mem1_reg[167][9]/P0001 ,
		_w11930_,
		_w11975_,
		_w21645_
	);
	LUT3 #(
		.INIT('h80)
	) name11133 (
		\wishbone_bd_ram_mem1_reg[92][9]/P0001 ,
		_w11954_,
		_w11972_,
		_w21646_
	);
	LUT4 #(
		.INIT('h0001)
	) name11134 (
		_w21643_,
		_w21644_,
		_w21645_,
		_w21646_,
		_w21647_
	);
	LUT4 #(
		.INIT('h8000)
	) name11135 (
		_w21632_,
		_w21637_,
		_w21642_,
		_w21647_,
		_w21648_
	);
	LUT3 #(
		.INIT('h80)
	) name11136 (
		\wishbone_bd_ram_mem1_reg[61][9]/P0001 ,
		_w11966_,
		_w11979_,
		_w21649_
	);
	LUT3 #(
		.INIT('h80)
	) name11137 (
		\wishbone_bd_ram_mem1_reg[99][9]/P0001 ,
		_w11938_,
		_w11965_,
		_w21650_
	);
	LUT3 #(
		.INIT('h80)
	) name11138 (
		\wishbone_bd_ram_mem1_reg[228][9]/P0001 ,
		_w11929_,
		_w11982_,
		_w21651_
	);
	LUT3 #(
		.INIT('h80)
	) name11139 (
		\wishbone_bd_ram_mem1_reg[115][9]/P0001 ,
		_w11938_,
		_w12012_,
		_w21652_
	);
	LUT4 #(
		.INIT('h0001)
	) name11140 (
		_w21649_,
		_w21650_,
		_w21651_,
		_w21652_,
		_w21653_
	);
	LUT3 #(
		.INIT('h80)
	) name11141 (
		\wishbone_bd_ram_mem1_reg[168][9]/P0001 ,
		_w11930_,
		_w11990_,
		_w21654_
	);
	LUT3 #(
		.INIT('h80)
	) name11142 (
		\wishbone_bd_ram_mem1_reg[227][9]/P0001 ,
		_w11938_,
		_w11982_,
		_w21655_
	);
	LUT3 #(
		.INIT('h80)
	) name11143 (
		\wishbone_bd_ram_mem1_reg[55][9]/P0001 ,
		_w11975_,
		_w11979_,
		_w21656_
	);
	LUT3 #(
		.INIT('h80)
	) name11144 (
		\wishbone_bd_ram_mem1_reg[116][9]/P0001 ,
		_w11929_,
		_w12012_,
		_w21657_
	);
	LUT4 #(
		.INIT('h0001)
	) name11145 (
		_w21654_,
		_w21655_,
		_w21656_,
		_w21657_,
		_w21658_
	);
	LUT3 #(
		.INIT('h80)
	) name11146 (
		\wishbone_bd_ram_mem1_reg[49][9]/P0001 ,
		_w11977_,
		_w11979_,
		_w21659_
	);
	LUT3 #(
		.INIT('h80)
	) name11147 (
		\wishbone_bd_ram_mem1_reg[100][9]/P0001 ,
		_w11929_,
		_w11965_,
		_w21660_
	);
	LUT3 #(
		.INIT('h80)
	) name11148 (
		\wishbone_bd_ram_mem1_reg[80][9]/P0001 ,
		_w11941_,
		_w11972_,
		_w21661_
	);
	LUT3 #(
		.INIT('h80)
	) name11149 (
		\wishbone_bd_ram_mem1_reg[90][9]/P0001 ,
		_w11944_,
		_w11972_,
		_w21662_
	);
	LUT4 #(
		.INIT('h0001)
	) name11150 (
		_w21659_,
		_w21660_,
		_w21661_,
		_w21662_,
		_w21663_
	);
	LUT3 #(
		.INIT('h80)
	) name11151 (
		\wishbone_bd_ram_mem1_reg[255][9]/P0001 ,
		_w11952_,
		_w11973_,
		_w21664_
	);
	LUT3 #(
		.INIT('h80)
	) name11152 (
		\wishbone_bd_ram_mem1_reg[207][9]/P0001 ,
		_w11945_,
		_w11973_,
		_w21665_
	);
	LUT3 #(
		.INIT('h80)
	) name11153 (
		\wishbone_bd_ram_mem1_reg[121][9]/P0001 ,
		_w11968_,
		_w12012_,
		_w21666_
	);
	LUT3 #(
		.INIT('h80)
	) name11154 (
		\wishbone_bd_ram_mem1_reg[29][9]/P0001 ,
		_w11935_,
		_w11966_,
		_w21667_
	);
	LUT4 #(
		.INIT('h0001)
	) name11155 (
		_w21664_,
		_w21665_,
		_w21666_,
		_w21667_,
		_w21668_
	);
	LUT4 #(
		.INIT('h8000)
	) name11156 (
		_w21653_,
		_w21658_,
		_w21663_,
		_w21668_,
		_w21669_
	);
	LUT4 #(
		.INIT('h8000)
	) name11157 (
		_w21606_,
		_w21627_,
		_w21648_,
		_w21669_,
		_w21670_
	);
	LUT3 #(
		.INIT('h80)
	) name11158 (
		\wishbone_bd_ram_mem1_reg[0][9]/P0001 ,
		_w11932_,
		_w11941_,
		_w21671_
	);
	LUT3 #(
		.INIT('h80)
	) name11159 (
		\wishbone_bd_ram_mem1_reg[164][9]/P0001 ,
		_w11929_,
		_w11930_,
		_w21672_
	);
	LUT3 #(
		.INIT('h80)
	) name11160 (
		\wishbone_bd_ram_mem1_reg[65][9]/P0001 ,
		_w11949_,
		_w11977_,
		_w21673_
	);
	LUT3 #(
		.INIT('h80)
	) name11161 (
		\wishbone_bd_ram_mem1_reg[47][9]/P0001 ,
		_w11957_,
		_w11973_,
		_w21674_
	);
	LUT4 #(
		.INIT('h0001)
	) name11162 (
		_w21671_,
		_w21672_,
		_w21673_,
		_w21674_,
		_w21675_
	);
	LUT3 #(
		.INIT('h80)
	) name11163 (
		\wishbone_bd_ram_mem1_reg[148][9]/P0001 ,
		_w11929_,
		_w11959_,
		_w21676_
	);
	LUT3 #(
		.INIT('h80)
	) name11164 (
		\wishbone_bd_ram_mem1_reg[58][9]/P0001 ,
		_w11944_,
		_w11979_,
		_w21677_
	);
	LUT3 #(
		.INIT('h80)
	) name11165 (
		\wishbone_bd_ram_mem1_reg[245][9]/P0001 ,
		_w11933_,
		_w11952_,
		_w21678_
	);
	LUT3 #(
		.INIT('h80)
	) name11166 (
		\wishbone_bd_ram_mem1_reg[137][9]/P0001 ,
		_w11955_,
		_w11968_,
		_w21679_
	);
	LUT4 #(
		.INIT('h0001)
	) name11167 (
		_w21676_,
		_w21677_,
		_w21678_,
		_w21679_,
		_w21680_
	);
	LUT3 #(
		.INIT('h80)
	) name11168 (
		\wishbone_bd_ram_mem1_reg[182][9]/P0001 ,
		_w11942_,
		_w11986_,
		_w21681_
	);
	LUT3 #(
		.INIT('h80)
	) name11169 (
		\wishbone_bd_ram_mem1_reg[67][9]/P0001 ,
		_w11938_,
		_w11949_,
		_w21682_
	);
	LUT3 #(
		.INIT('h80)
	) name11170 (
		\wishbone_bd_ram_mem1_reg[24][9]/P0001 ,
		_w11935_,
		_w11990_,
		_w21683_
	);
	LUT3 #(
		.INIT('h80)
	) name11171 (
		\wishbone_bd_ram_mem1_reg[71][9]/P0001 ,
		_w11949_,
		_w11975_,
		_w21684_
	);
	LUT4 #(
		.INIT('h0001)
	) name11172 (
		_w21681_,
		_w21682_,
		_w21683_,
		_w21684_,
		_w21685_
	);
	LUT3 #(
		.INIT('h80)
	) name11173 (
		\wishbone_bd_ram_mem1_reg[113][9]/P0001 ,
		_w11977_,
		_w12012_,
		_w21686_
	);
	LUT3 #(
		.INIT('h80)
	) name11174 (
		\wishbone_bd_ram_mem1_reg[192][9]/P0001 ,
		_w11941_,
		_w11945_,
		_w21687_
	);
	LUT3 #(
		.INIT('h80)
	) name11175 (
		\wishbone_bd_ram_mem1_reg[222][9]/P0001 ,
		_w11948_,
		_w11984_,
		_w21688_
	);
	LUT3 #(
		.INIT('h80)
	) name11176 (
		\wishbone_bd_ram_mem1_reg[75][9]/P0001 ,
		_w11936_,
		_w11949_,
		_w21689_
	);
	LUT4 #(
		.INIT('h0001)
	) name11177 (
		_w21686_,
		_w21687_,
		_w21688_,
		_w21689_,
		_w21690_
	);
	LUT4 #(
		.INIT('h8000)
	) name11178 (
		_w21675_,
		_w21680_,
		_w21685_,
		_w21690_,
		_w21691_
	);
	LUT3 #(
		.INIT('h80)
	) name11179 (
		\wishbone_bd_ram_mem1_reg[221][9]/P0001 ,
		_w11966_,
		_w11984_,
		_w21692_
	);
	LUT3 #(
		.INIT('h80)
	) name11180 (
		\wishbone_bd_ram_mem1_reg[72][9]/P0001 ,
		_w11949_,
		_w11990_,
		_w21693_
	);
	LUT3 #(
		.INIT('h80)
	) name11181 (
		\wishbone_bd_ram_mem1_reg[37][9]/P0001 ,
		_w11933_,
		_w11957_,
		_w21694_
	);
	LUT3 #(
		.INIT('h80)
	) name11182 (
		\wishbone_bd_ram_mem1_reg[161][9]/P0001 ,
		_w11930_,
		_w11977_,
		_w21695_
	);
	LUT4 #(
		.INIT('h0001)
	) name11183 (
		_w21692_,
		_w21693_,
		_w21694_,
		_w21695_,
		_w21696_
	);
	LUT3 #(
		.INIT('h80)
	) name11184 (
		\wishbone_bd_ram_mem1_reg[190][9]/P0001 ,
		_w11942_,
		_w11948_,
		_w21697_
	);
	LUT3 #(
		.INIT('h80)
	) name11185 (
		\wishbone_bd_ram_mem1_reg[253][9]/P0001 ,
		_w11952_,
		_w11966_,
		_w21698_
	);
	LUT3 #(
		.INIT('h80)
	) name11186 (
		\wishbone_bd_ram_mem1_reg[158][9]/P0001 ,
		_w11948_,
		_w11959_,
		_w21699_
	);
	LUT3 #(
		.INIT('h80)
	) name11187 (
		\wishbone_bd_ram_mem1_reg[38][9]/P0001 ,
		_w11957_,
		_w11986_,
		_w21700_
	);
	LUT4 #(
		.INIT('h0001)
	) name11188 (
		_w21697_,
		_w21698_,
		_w21699_,
		_w21700_,
		_w21701_
	);
	LUT3 #(
		.INIT('h80)
	) name11189 (
		\wishbone_bd_ram_mem1_reg[135][9]/P0001 ,
		_w11955_,
		_w11975_,
		_w21702_
	);
	LUT3 #(
		.INIT('h80)
	) name11190 (
		\wishbone_bd_ram_mem1_reg[5][9]/P0001 ,
		_w11932_,
		_w11933_,
		_w21703_
	);
	LUT3 #(
		.INIT('h80)
	) name11191 (
		\wishbone_bd_ram_mem1_reg[28][9]/P0001 ,
		_w11935_,
		_w11954_,
		_w21704_
	);
	LUT3 #(
		.INIT('h80)
	) name11192 (
		\wishbone_bd_ram_mem1_reg[159][9]/P0001 ,
		_w11959_,
		_w11973_,
		_w21705_
	);
	LUT4 #(
		.INIT('h0001)
	) name11193 (
		_w21702_,
		_w21703_,
		_w21704_,
		_w21705_,
		_w21706_
	);
	LUT3 #(
		.INIT('h80)
	) name11194 (
		\wishbone_bd_ram_mem1_reg[6][9]/P0001 ,
		_w11932_,
		_w11986_,
		_w21707_
	);
	LUT3 #(
		.INIT('h80)
	) name11195 (
		\wishbone_bd_ram_mem1_reg[51][9]/P0001 ,
		_w11938_,
		_w11979_,
		_w21708_
	);
	LUT3 #(
		.INIT('h80)
	) name11196 (
		\wishbone_bd_ram_mem1_reg[147][9]/P0001 ,
		_w11938_,
		_w11959_,
		_w21709_
	);
	LUT3 #(
		.INIT('h80)
	) name11197 (
		\wishbone_bd_ram_mem1_reg[230][9]/P0001 ,
		_w11982_,
		_w11986_,
		_w21710_
	);
	LUT4 #(
		.INIT('h0001)
	) name11198 (
		_w21707_,
		_w21708_,
		_w21709_,
		_w21710_,
		_w21711_
	);
	LUT4 #(
		.INIT('h8000)
	) name11199 (
		_w21696_,
		_w21701_,
		_w21706_,
		_w21711_,
		_w21712_
	);
	LUT3 #(
		.INIT('h80)
	) name11200 (
		\wishbone_bd_ram_mem1_reg[239][9]/P0001 ,
		_w11973_,
		_w11982_,
		_w21713_
	);
	LUT3 #(
		.INIT('h80)
	) name11201 (
		\wishbone_bd_ram_mem1_reg[19][9]/P0001 ,
		_w11935_,
		_w11938_,
		_w21714_
	);
	LUT3 #(
		.INIT('h80)
	) name11202 (
		\wishbone_bd_ram_mem1_reg[44][9]/P0001 ,
		_w11954_,
		_w11957_,
		_w21715_
	);
	LUT3 #(
		.INIT('h80)
	) name11203 (
		\wishbone_bd_ram_mem1_reg[191][9]/P0001 ,
		_w11942_,
		_w11973_,
		_w21716_
	);
	LUT4 #(
		.INIT('h0001)
	) name11204 (
		_w21713_,
		_w21714_,
		_w21715_,
		_w21716_,
		_w21717_
	);
	LUT3 #(
		.INIT('h80)
	) name11205 (
		\wishbone_bd_ram_mem1_reg[31][9]/P0001 ,
		_w11935_,
		_w11973_,
		_w21718_
	);
	LUT3 #(
		.INIT('h80)
	) name11206 (
		\wishbone_bd_ram_mem1_reg[89][9]/P0001 ,
		_w11968_,
		_w11972_,
		_w21719_
	);
	LUT3 #(
		.INIT('h80)
	) name11207 (
		\wishbone_bd_ram_mem1_reg[136][9]/P0001 ,
		_w11955_,
		_w11990_,
		_w21720_
	);
	LUT3 #(
		.INIT('h80)
	) name11208 (
		\wishbone_bd_ram_mem1_reg[23][9]/P0001 ,
		_w11935_,
		_w11975_,
		_w21721_
	);
	LUT4 #(
		.INIT('h0001)
	) name11209 (
		_w21718_,
		_w21719_,
		_w21720_,
		_w21721_,
		_w21722_
	);
	LUT3 #(
		.INIT('h80)
	) name11210 (
		\wishbone_bd_ram_mem1_reg[3][9]/P0001 ,
		_w11932_,
		_w11938_,
		_w21723_
	);
	LUT3 #(
		.INIT('h80)
	) name11211 (
		\wishbone_bd_ram_mem1_reg[216][9]/P0001 ,
		_w11984_,
		_w11990_,
		_w21724_
	);
	LUT3 #(
		.INIT('h80)
	) name11212 (
		\wishbone_bd_ram_mem1_reg[104][9]/P0001 ,
		_w11965_,
		_w11990_,
		_w21725_
	);
	LUT3 #(
		.INIT('h80)
	) name11213 (
		\wishbone_bd_ram_mem1_reg[183][9]/P0001 ,
		_w11942_,
		_w11975_,
		_w21726_
	);
	LUT4 #(
		.INIT('h0001)
	) name11214 (
		_w21723_,
		_w21724_,
		_w21725_,
		_w21726_,
		_w21727_
	);
	LUT3 #(
		.INIT('h80)
	) name11215 (
		\wishbone_bd_ram_mem1_reg[128][9]/P0001 ,
		_w11941_,
		_w11955_,
		_w21728_
	);
	LUT3 #(
		.INIT('h80)
	) name11216 (
		\wishbone_bd_ram_mem1_reg[93][9]/P0001 ,
		_w11966_,
		_w11972_,
		_w21729_
	);
	LUT3 #(
		.INIT('h80)
	) name11217 (
		\wishbone_bd_ram_mem1_reg[105][9]/P0001 ,
		_w11965_,
		_w11968_,
		_w21730_
	);
	LUT3 #(
		.INIT('h80)
	) name11218 (
		\wishbone_bd_ram_mem1_reg[243][9]/P0001 ,
		_w11938_,
		_w11952_,
		_w21731_
	);
	LUT4 #(
		.INIT('h0001)
	) name11219 (
		_w21728_,
		_w21729_,
		_w21730_,
		_w21731_,
		_w21732_
	);
	LUT4 #(
		.INIT('h8000)
	) name11220 (
		_w21717_,
		_w21722_,
		_w21727_,
		_w21732_,
		_w21733_
	);
	LUT3 #(
		.INIT('h80)
	) name11221 (
		\wishbone_bd_ram_mem1_reg[200][9]/P0001 ,
		_w11945_,
		_w11990_,
		_w21734_
	);
	LUT3 #(
		.INIT('h80)
	) name11222 (
		\wishbone_bd_ram_mem1_reg[179][9]/P0001 ,
		_w11938_,
		_w11942_,
		_w21735_
	);
	LUT3 #(
		.INIT('h80)
	) name11223 (
		\wishbone_bd_ram_mem1_reg[59][9]/P0001 ,
		_w11936_,
		_w11979_,
		_w21736_
	);
	LUT3 #(
		.INIT('h80)
	) name11224 (
		\wishbone_bd_ram_mem1_reg[11][9]/P0001 ,
		_w11932_,
		_w11936_,
		_w21737_
	);
	LUT4 #(
		.INIT('h0001)
	) name11225 (
		_w21734_,
		_w21735_,
		_w21736_,
		_w21737_,
		_w21738_
	);
	LUT3 #(
		.INIT('h80)
	) name11226 (
		\wishbone_bd_ram_mem1_reg[177][9]/P0001 ,
		_w11942_,
		_w11977_,
		_w21739_
	);
	LUT3 #(
		.INIT('h80)
	) name11227 (
		\wishbone_bd_ram_mem1_reg[247][9]/P0001 ,
		_w11952_,
		_w11975_,
		_w21740_
	);
	LUT3 #(
		.INIT('h80)
	) name11228 (
		\wishbone_bd_ram_mem1_reg[229][9]/P0001 ,
		_w11933_,
		_w11982_,
		_w21741_
	);
	LUT3 #(
		.INIT('h80)
	) name11229 (
		\wishbone_bd_ram_mem1_reg[175][9]/P0001 ,
		_w11930_,
		_w11973_,
		_w21742_
	);
	LUT4 #(
		.INIT('h0001)
	) name11230 (
		_w21739_,
		_w21740_,
		_w21741_,
		_w21742_,
		_w21743_
	);
	LUT3 #(
		.INIT('h80)
	) name11231 (
		\wishbone_bd_ram_mem1_reg[225][9]/P0001 ,
		_w11977_,
		_w11982_,
		_w21744_
	);
	LUT3 #(
		.INIT('h80)
	) name11232 (
		\wishbone_bd_ram_mem1_reg[62][9]/P0001 ,
		_w11948_,
		_w11979_,
		_w21745_
	);
	LUT3 #(
		.INIT('h80)
	) name11233 (
		\wishbone_bd_ram_mem1_reg[219][9]/P0001 ,
		_w11936_,
		_w11984_,
		_w21746_
	);
	LUT3 #(
		.INIT('h80)
	) name11234 (
		\wishbone_bd_ram_mem1_reg[172][9]/P0001 ,
		_w11930_,
		_w11954_,
		_w21747_
	);
	LUT4 #(
		.INIT('h0001)
	) name11235 (
		_w21744_,
		_w21745_,
		_w21746_,
		_w21747_,
		_w21748_
	);
	LUT3 #(
		.INIT('h80)
	) name11236 (
		\wishbone_bd_ram_mem1_reg[46][9]/P0001 ,
		_w11948_,
		_w11957_,
		_w21749_
	);
	LUT3 #(
		.INIT('h80)
	) name11237 (
		\wishbone_bd_ram_mem1_reg[232][9]/P0001 ,
		_w11982_,
		_w11990_,
		_w21750_
	);
	LUT3 #(
		.INIT('h80)
	) name11238 (
		\wishbone_bd_ram_mem1_reg[79][9]/P0001 ,
		_w11949_,
		_w11973_,
		_w21751_
	);
	LUT3 #(
		.INIT('h80)
	) name11239 (
		\wishbone_bd_ram_mem1_reg[50][9]/P0001 ,
		_w11963_,
		_w11979_,
		_w21752_
	);
	LUT4 #(
		.INIT('h0001)
	) name11240 (
		_w21749_,
		_w21750_,
		_w21751_,
		_w21752_,
		_w21753_
	);
	LUT4 #(
		.INIT('h8000)
	) name11241 (
		_w21738_,
		_w21743_,
		_w21748_,
		_w21753_,
		_w21754_
	);
	LUT4 #(
		.INIT('h8000)
	) name11242 (
		_w21691_,
		_w21712_,
		_w21733_,
		_w21754_,
		_w21755_
	);
	LUT3 #(
		.INIT('h80)
	) name11243 (
		\wishbone_bd_ram_mem1_reg[26][9]/P0001 ,
		_w11935_,
		_w11944_,
		_w21756_
	);
	LUT3 #(
		.INIT('h80)
	) name11244 (
		\wishbone_bd_ram_mem1_reg[124][9]/P0001 ,
		_w11954_,
		_w12012_,
		_w21757_
	);
	LUT3 #(
		.INIT('h80)
	) name11245 (
		\wishbone_bd_ram_mem1_reg[33][9]/P0001 ,
		_w11957_,
		_w11977_,
		_w21758_
	);
	LUT3 #(
		.INIT('h80)
	) name11246 (
		\wishbone_bd_ram_mem1_reg[112][9]/P0001 ,
		_w11941_,
		_w12012_,
		_w21759_
	);
	LUT4 #(
		.INIT('h0001)
	) name11247 (
		_w21756_,
		_w21757_,
		_w21758_,
		_w21759_,
		_w21760_
	);
	LUT3 #(
		.INIT('h80)
	) name11248 (
		\wishbone_bd_ram_mem1_reg[145][9]/P0001 ,
		_w11959_,
		_w11977_,
		_w21761_
	);
	LUT3 #(
		.INIT('h80)
	) name11249 (
		\wishbone_bd_ram_mem1_reg[218][9]/P0001 ,
		_w11944_,
		_w11984_,
		_w21762_
	);
	LUT3 #(
		.INIT('h80)
	) name11250 (
		\wishbone_bd_ram_mem1_reg[78][9]/P0001 ,
		_w11948_,
		_w11949_,
		_w21763_
	);
	LUT3 #(
		.INIT('h80)
	) name11251 (
		\wishbone_bd_ram_mem1_reg[53][9]/P0001 ,
		_w11933_,
		_w11979_,
		_w21764_
	);
	LUT4 #(
		.INIT('h0001)
	) name11252 (
		_w21761_,
		_w21762_,
		_w21763_,
		_w21764_,
		_w21765_
	);
	LUT3 #(
		.INIT('h80)
	) name11253 (
		\wishbone_bd_ram_mem1_reg[155][9]/P0001 ,
		_w11936_,
		_w11959_,
		_w21766_
	);
	LUT3 #(
		.INIT('h80)
	) name11254 (
		\wishbone_bd_ram_mem1_reg[163][9]/P0001 ,
		_w11930_,
		_w11938_,
		_w21767_
	);
	LUT3 #(
		.INIT('h80)
	) name11255 (
		\wishbone_bd_ram_mem1_reg[74][9]/P0001 ,
		_w11944_,
		_w11949_,
		_w21768_
	);
	LUT3 #(
		.INIT('h80)
	) name11256 (
		\wishbone_bd_ram_mem1_reg[212][9]/P0001 ,
		_w11929_,
		_w11984_,
		_w21769_
	);
	LUT4 #(
		.INIT('h0001)
	) name11257 (
		_w21766_,
		_w21767_,
		_w21768_,
		_w21769_,
		_w21770_
	);
	LUT3 #(
		.INIT('h80)
	) name11258 (
		\wishbone_bd_ram_mem1_reg[15][9]/P0001 ,
		_w11932_,
		_w11973_,
		_w21771_
	);
	LUT3 #(
		.INIT('h80)
	) name11259 (
		\wishbone_bd_ram_mem1_reg[8][9]/P0001 ,
		_w11932_,
		_w11990_,
		_w21772_
	);
	LUT3 #(
		.INIT('h80)
	) name11260 (
		\wishbone_bd_ram_mem1_reg[169][9]/P0001 ,
		_w11930_,
		_w11968_,
		_w21773_
	);
	LUT3 #(
		.INIT('h80)
	) name11261 (
		\wishbone_bd_ram_mem1_reg[141][9]/P0001 ,
		_w11955_,
		_w11966_,
		_w21774_
	);
	LUT4 #(
		.INIT('h0001)
	) name11262 (
		_w21771_,
		_w21772_,
		_w21773_,
		_w21774_,
		_w21775_
	);
	LUT4 #(
		.INIT('h8000)
	) name11263 (
		_w21760_,
		_w21765_,
		_w21770_,
		_w21775_,
		_w21776_
	);
	LUT3 #(
		.INIT('h80)
	) name11264 (
		\wishbone_bd_ram_mem1_reg[43][9]/P0001 ,
		_w11936_,
		_w11957_,
		_w21777_
	);
	LUT3 #(
		.INIT('h80)
	) name11265 (
		\wishbone_bd_ram_mem1_reg[70][9]/P0001 ,
		_w11949_,
		_w11986_,
		_w21778_
	);
	LUT3 #(
		.INIT('h80)
	) name11266 (
		\wishbone_bd_ram_mem1_reg[60][9]/P0001 ,
		_w11954_,
		_w11979_,
		_w21779_
	);
	LUT3 #(
		.INIT('h80)
	) name11267 (
		\wishbone_bd_ram_mem1_reg[88][9]/P0001 ,
		_w11972_,
		_w11990_,
		_w21780_
	);
	LUT4 #(
		.INIT('h0001)
	) name11268 (
		_w21777_,
		_w21778_,
		_w21779_,
		_w21780_,
		_w21781_
	);
	LUT3 #(
		.INIT('h80)
	) name11269 (
		\wishbone_bd_ram_mem1_reg[96][9]/P0001 ,
		_w11941_,
		_w11965_,
		_w21782_
	);
	LUT3 #(
		.INIT('h80)
	) name11270 (
		\wishbone_bd_ram_mem1_reg[81][9]/P0001 ,
		_w11972_,
		_w11977_,
		_w21783_
	);
	LUT3 #(
		.INIT('h80)
	) name11271 (
		\wishbone_bd_ram_mem1_reg[14][9]/P0001 ,
		_w11932_,
		_w11948_,
		_w21784_
	);
	LUT3 #(
		.INIT('h80)
	) name11272 (
		\wishbone_bd_ram_mem1_reg[66][9]/P0001 ,
		_w11949_,
		_w11963_,
		_w21785_
	);
	LUT4 #(
		.INIT('h0001)
	) name11273 (
		_w21782_,
		_w21783_,
		_w21784_,
		_w21785_,
		_w21786_
	);
	LUT3 #(
		.INIT('h80)
	) name11274 (
		\wishbone_bd_ram_mem1_reg[203][9]/P0001 ,
		_w11936_,
		_w11945_,
		_w21787_
	);
	LUT3 #(
		.INIT('h80)
	) name11275 (
		\wishbone_bd_ram_mem1_reg[234][9]/P0001 ,
		_w11944_,
		_w11982_,
		_w21788_
	);
	LUT3 #(
		.INIT('h80)
	) name11276 (
		\wishbone_bd_ram_mem1_reg[198][9]/P0001 ,
		_w11945_,
		_w11986_,
		_w21789_
	);
	LUT3 #(
		.INIT('h80)
	) name11277 (
		\wishbone_bd_ram_mem1_reg[131][9]/P0001 ,
		_w11938_,
		_w11955_,
		_w21790_
	);
	LUT4 #(
		.INIT('h0001)
	) name11278 (
		_w21787_,
		_w21788_,
		_w21789_,
		_w21790_,
		_w21791_
	);
	LUT3 #(
		.INIT('h80)
	) name11279 (
		\wishbone_bd_ram_mem1_reg[69][9]/P0001 ,
		_w11933_,
		_w11949_,
		_w21792_
	);
	LUT3 #(
		.INIT('h80)
	) name11280 (
		\wishbone_bd_ram_mem1_reg[108][9]/P0001 ,
		_w11954_,
		_w11965_,
		_w21793_
	);
	LUT3 #(
		.INIT('h80)
	) name11281 (
		\wishbone_bd_ram_mem1_reg[248][9]/P0001 ,
		_w11952_,
		_w11990_,
		_w21794_
	);
	LUT3 #(
		.INIT('h80)
	) name11282 (
		\wishbone_bd_ram_mem1_reg[101][9]/P0001 ,
		_w11933_,
		_w11965_,
		_w21795_
	);
	LUT4 #(
		.INIT('h0001)
	) name11283 (
		_w21792_,
		_w21793_,
		_w21794_,
		_w21795_,
		_w21796_
	);
	LUT4 #(
		.INIT('h8000)
	) name11284 (
		_w21781_,
		_w21786_,
		_w21791_,
		_w21796_,
		_w21797_
	);
	LUT3 #(
		.INIT('h80)
	) name11285 (
		\wishbone_bd_ram_mem1_reg[211][9]/P0001 ,
		_w11938_,
		_w11984_,
		_w21798_
	);
	LUT3 #(
		.INIT('h80)
	) name11286 (
		\wishbone_bd_ram_mem1_reg[187][9]/P0001 ,
		_w11936_,
		_w11942_,
		_w21799_
	);
	LUT3 #(
		.INIT('h80)
	) name11287 (
		\wishbone_bd_ram_mem1_reg[140][9]/P0001 ,
		_w11954_,
		_w11955_,
		_w21800_
	);
	LUT3 #(
		.INIT('h80)
	) name11288 (
		\wishbone_bd_ram_mem1_reg[162][9]/P0001 ,
		_w11930_,
		_w11963_,
		_w21801_
	);
	LUT4 #(
		.INIT('h0001)
	) name11289 (
		_w21798_,
		_w21799_,
		_w21800_,
		_w21801_,
		_w21802_
	);
	LUT3 #(
		.INIT('h80)
	) name11290 (
		\wishbone_bd_ram_mem1_reg[125][9]/P0001 ,
		_w11966_,
		_w12012_,
		_w21803_
	);
	LUT3 #(
		.INIT('h80)
	) name11291 (
		\wishbone_bd_ram_mem1_reg[91][9]/P0001 ,
		_w11936_,
		_w11972_,
		_w21804_
	);
	LUT3 #(
		.INIT('h80)
	) name11292 (
		\wishbone_bd_ram_mem1_reg[152][9]/P0001 ,
		_w11959_,
		_w11990_,
		_w21805_
	);
	LUT3 #(
		.INIT('h80)
	) name11293 (
		\wishbone_bd_ram_mem1_reg[94][9]/P0001 ,
		_w11948_,
		_w11972_,
		_w21806_
	);
	LUT4 #(
		.INIT('h0001)
	) name11294 (
		_w21803_,
		_w21804_,
		_w21805_,
		_w21806_,
		_w21807_
	);
	LUT3 #(
		.INIT('h80)
	) name11295 (
		\wishbone_bd_ram_mem1_reg[12][9]/P0001 ,
		_w11932_,
		_w11954_,
		_w21808_
	);
	LUT3 #(
		.INIT('h80)
	) name11296 (
		\wishbone_bd_ram_mem1_reg[35][9]/P0001 ,
		_w11938_,
		_w11957_,
		_w21809_
	);
	LUT3 #(
		.INIT('h80)
	) name11297 (
		\wishbone_bd_ram_mem1_reg[16][9]/P0001 ,
		_w11935_,
		_w11941_,
		_w21810_
	);
	LUT3 #(
		.INIT('h80)
	) name11298 (
		\wishbone_bd_ram_mem1_reg[103][9]/P0001 ,
		_w11965_,
		_w11975_,
		_w21811_
	);
	LUT4 #(
		.INIT('h0001)
	) name11299 (
		_w21808_,
		_w21809_,
		_w21810_,
		_w21811_,
		_w21812_
	);
	LUT3 #(
		.INIT('h80)
	) name11300 (
		\wishbone_bd_ram_mem1_reg[233][9]/P0001 ,
		_w11968_,
		_w11982_,
		_w21813_
	);
	LUT3 #(
		.INIT('h80)
	) name11301 (
		\wishbone_bd_ram_mem1_reg[143][9]/P0001 ,
		_w11955_,
		_w11973_,
		_w21814_
	);
	LUT3 #(
		.INIT('h80)
	) name11302 (
		\wishbone_bd_ram_mem1_reg[226][9]/P0001 ,
		_w11963_,
		_w11982_,
		_w21815_
	);
	LUT3 #(
		.INIT('h80)
	) name11303 (
		\wishbone_bd_ram_mem1_reg[18][9]/P0001 ,
		_w11935_,
		_w11963_,
		_w21816_
	);
	LUT4 #(
		.INIT('h0001)
	) name11304 (
		_w21813_,
		_w21814_,
		_w21815_,
		_w21816_,
		_w21817_
	);
	LUT4 #(
		.INIT('h8000)
	) name11305 (
		_w21802_,
		_w21807_,
		_w21812_,
		_w21817_,
		_w21818_
	);
	LUT3 #(
		.INIT('h80)
	) name11306 (
		\wishbone_bd_ram_mem1_reg[153][9]/P0001 ,
		_w11959_,
		_w11968_,
		_w21819_
	);
	LUT3 #(
		.INIT('h80)
	) name11307 (
		\wishbone_bd_ram_mem1_reg[122][9]/P0001 ,
		_w11944_,
		_w12012_,
		_w21820_
	);
	LUT3 #(
		.INIT('h80)
	) name11308 (
		\wishbone_bd_ram_mem1_reg[98][9]/P0001 ,
		_w11963_,
		_w11965_,
		_w21821_
	);
	LUT3 #(
		.INIT('h80)
	) name11309 (
		\wishbone_bd_ram_mem1_reg[110][9]/P0001 ,
		_w11948_,
		_w11965_,
		_w21822_
	);
	LUT4 #(
		.INIT('h0001)
	) name11310 (
		_w21819_,
		_w21820_,
		_w21821_,
		_w21822_,
		_w21823_
	);
	LUT3 #(
		.INIT('h80)
	) name11311 (
		\wishbone_bd_ram_mem1_reg[240][9]/P0001 ,
		_w11941_,
		_w11952_,
		_w21824_
	);
	LUT3 #(
		.INIT('h80)
	) name11312 (
		\wishbone_bd_ram_mem1_reg[114][9]/P0001 ,
		_w11963_,
		_w12012_,
		_w21825_
	);
	LUT3 #(
		.INIT('h80)
	) name11313 (
		\wishbone_bd_ram_mem1_reg[150][9]/P0001 ,
		_w11959_,
		_w11986_,
		_w21826_
	);
	LUT3 #(
		.INIT('h80)
	) name11314 (
		\wishbone_bd_ram_mem1_reg[242][9]/P0001 ,
		_w11952_,
		_w11963_,
		_w21827_
	);
	LUT4 #(
		.INIT('h0001)
	) name11315 (
		_w21824_,
		_w21825_,
		_w21826_,
		_w21827_,
		_w21828_
	);
	LUT3 #(
		.INIT('h80)
	) name11316 (
		\wishbone_bd_ram_mem1_reg[76][9]/P0001 ,
		_w11949_,
		_w11954_,
		_w21829_
	);
	LUT3 #(
		.INIT('h80)
	) name11317 (
		\wishbone_bd_ram_mem1_reg[214][9]/P0001 ,
		_w11984_,
		_w11986_,
		_w21830_
	);
	LUT3 #(
		.INIT('h80)
	) name11318 (
		\wishbone_bd_ram_mem1_reg[210][9]/P0001 ,
		_w11963_,
		_w11984_,
		_w21831_
	);
	LUT3 #(
		.INIT('h80)
	) name11319 (
		\wishbone_bd_ram_mem1_reg[188][9]/P0001 ,
		_w11942_,
		_w11954_,
		_w21832_
	);
	LUT4 #(
		.INIT('h0001)
	) name11320 (
		_w21829_,
		_w21830_,
		_w21831_,
		_w21832_,
		_w21833_
	);
	LUT3 #(
		.INIT('h80)
	) name11321 (
		\wishbone_bd_ram_mem1_reg[63][9]/P0001 ,
		_w11973_,
		_w11979_,
		_w21834_
	);
	LUT3 #(
		.INIT('h80)
	) name11322 (
		\wishbone_bd_ram_mem1_reg[176][9]/P0001 ,
		_w11941_,
		_w11942_,
		_w21835_
	);
	LUT3 #(
		.INIT('h80)
	) name11323 (
		\wishbone_bd_ram_mem1_reg[41][9]/P0001 ,
		_w11957_,
		_w11968_,
		_w21836_
	);
	LUT3 #(
		.INIT('h80)
	) name11324 (
		\wishbone_bd_ram_mem1_reg[199][9]/P0001 ,
		_w11945_,
		_w11975_,
		_w21837_
	);
	LUT4 #(
		.INIT('h0001)
	) name11325 (
		_w21834_,
		_w21835_,
		_w21836_,
		_w21837_,
		_w21838_
	);
	LUT4 #(
		.INIT('h8000)
	) name11326 (
		_w21823_,
		_w21828_,
		_w21833_,
		_w21838_,
		_w21839_
	);
	LUT4 #(
		.INIT('h8000)
	) name11327 (
		_w21776_,
		_w21797_,
		_w21818_,
		_w21839_,
		_w21840_
	);
	LUT4 #(
		.INIT('h8000)
	) name11328 (
		_w21585_,
		_w21670_,
		_w21755_,
		_w21840_,
		_w21841_
	);
	LUT4 #(
		.INIT('h1555)
	) name11329 (
		wb_rst_i_pad,
		_w21490_,
		_w21494_,
		_w21499_,
		_w21842_
	);
	LUT3 #(
		.INIT('hba)
	) name11330 (
		_w21500_,
		_w21841_,
		_w21842_,
		_w21843_
	);
	LUT3 #(
		.INIT('h80)
	) name11331 (
		\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 ,
		_w18753_,
		_w18754_,
		_w21844_
	);
	LUT4 #(
		.INIT('h0008)
	) name11332 (
		\ethreg1_RXHASH0_2_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21845_
	);
	LUT3 #(
		.INIT('h80)
	) name11333 (
		_w18757_,
		_w18758_,
		_w21845_,
		_w21846_
	);
	LUT4 #(
		.INIT('h0008)
	) name11334 (
		\ethreg1_RXHASH1_2_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21847_
	);
	LUT3 #(
		.INIT('h80)
	) name11335 (
		_w18757_,
		_w18762_,
		_w21847_,
		_w21848_
	);
	LUT4 #(
		.INIT('h0002)
	) name11336 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21849_
	);
	LUT3 #(
		.INIT('h80)
	) name11337 (
		_w18757_,
		_w18758_,
		_w21849_,
		_w21850_
	);
	LUT4 #(
		.INIT('h0002)
	) name11338 (
		_w18752_,
		_w21846_,
		_w21848_,
		_w21850_,
		_w21851_
	);
	LUT3 #(
		.INIT('h8a)
	) name11339 (
		_w18752_,
		_w21844_,
		_w21851_,
		_w21852_
	);
	LUT3 #(
		.INIT('h45)
	) name11340 (
		wb_rst_i_pad,
		_w21844_,
		_w21851_,
		_w21853_
	);
	LUT3 #(
		.INIT('hdc)
	) name11341 (
		_w14512_,
		_w21852_,
		_w21853_,
		_w21854_
	);
	LUT4 #(
		.INIT('h0002)
	) name11342 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21855_
	);
	LUT3 #(
		.INIT('h80)
	) name11343 (
		_w18757_,
		_w18762_,
		_w21855_,
		_w21856_
	);
	LUT3 #(
		.INIT('h80)
	) name11344 (
		\ethreg1_MIIRX_DATA_DataOut_reg[11]/NET0131 ,
		_w18785_,
		_w18786_,
		_w21857_
	);
	LUT4 #(
		.INIT('h0008)
	) name11345 (
		\ethreg1_RXHASH0_1_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21858_
	);
	LUT3 #(
		.INIT('h80)
	) name11346 (
		_w18757_,
		_w18758_,
		_w21858_,
		_w21859_
	);
	LUT4 #(
		.INIT('h0008)
	) name11347 (
		\ethreg1_RXHASH1_1_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21860_
	);
	LUT3 #(
		.INIT('h80)
	) name11348 (
		_w18757_,
		_w18762_,
		_w21860_,
		_w21861_
	);
	LUT4 #(
		.INIT('h0001)
	) name11349 (
		_w21856_,
		_w21857_,
		_w21859_,
		_w21861_,
		_w21862_
	);
	LUT4 #(
		.INIT('h0002)
	) name11350 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21863_
	);
	LUT4 #(
		.INIT('h0020)
	) name11351 (
		\ethreg1_TXCTRL_1_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w21864_
	);
	LUT4 #(
		.INIT('h777f)
	) name11352 (
		_w18757_,
		_w18758_,
		_w21863_,
		_w21864_,
		_w21865_
	);
	LUT2 #(
		.INIT('h8)
	) name11353 (
		_w18752_,
		_w21865_,
		_w21866_
	);
	LUT3 #(
		.INIT('h80)
	) name11354 (
		\ethreg1_MODER_1_DataOut_reg[3]/NET0131 ,
		_w18800_,
		_w18801_,
		_w21867_
	);
	LUT3 #(
		.INIT('h80)
	) name11355 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[3]/NET0131 ,
		_w18785_,
		_w18798_,
		_w21868_
	);
	LUT3 #(
		.INIT('h80)
	) name11356 (
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		_w18753_,
		_w18754_,
		_w21869_
	);
	LUT3 #(
		.INIT('h80)
	) name11357 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[3]/NET0131 ,
		_w18798_,
		_w18805_,
		_w21870_
	);
	LUT4 #(
		.INIT('h0001)
	) name11358 (
		_w21867_,
		_w21868_,
		_w21869_,
		_w21870_,
		_w21871_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name11359 (
		_w18752_,
		_w21862_,
		_w21865_,
		_w21871_,
		_w21872_
	);
	LUT3 #(
		.INIT('h80)
	) name11360 (
		\wishbone_bd_ram_mem1_reg[16][11]/P0001 ,
		_w11935_,
		_w11941_,
		_w21873_
	);
	LUT3 #(
		.INIT('h80)
	) name11361 (
		\wishbone_bd_ram_mem1_reg[84][11]/P0001 ,
		_w11929_,
		_w11972_,
		_w21874_
	);
	LUT3 #(
		.INIT('h80)
	) name11362 (
		\wishbone_bd_ram_mem1_reg[18][11]/P0001 ,
		_w11935_,
		_w11963_,
		_w21875_
	);
	LUT3 #(
		.INIT('h80)
	) name11363 (
		\wishbone_bd_ram_mem1_reg[138][11]/P0001 ,
		_w11944_,
		_w11955_,
		_w21876_
	);
	LUT4 #(
		.INIT('h0001)
	) name11364 (
		_w21873_,
		_w21874_,
		_w21875_,
		_w21876_,
		_w21877_
	);
	LUT3 #(
		.INIT('h80)
	) name11365 (
		\wishbone_bd_ram_mem1_reg[31][11]/P0001 ,
		_w11935_,
		_w11973_,
		_w21878_
	);
	LUT3 #(
		.INIT('h80)
	) name11366 (
		\wishbone_bd_ram_mem1_reg[142][11]/P0001 ,
		_w11948_,
		_w11955_,
		_w21879_
	);
	LUT3 #(
		.INIT('h80)
	) name11367 (
		\wishbone_bd_ram_mem1_reg[58][11]/P0001 ,
		_w11944_,
		_w11979_,
		_w21880_
	);
	LUT3 #(
		.INIT('h80)
	) name11368 (
		\wishbone_bd_ram_mem1_reg[4][11]/P0001 ,
		_w11929_,
		_w11932_,
		_w21881_
	);
	LUT4 #(
		.INIT('h0001)
	) name11369 (
		_w21878_,
		_w21879_,
		_w21880_,
		_w21881_,
		_w21882_
	);
	LUT3 #(
		.INIT('h80)
	) name11370 (
		\wishbone_bd_ram_mem1_reg[210][11]/P0001 ,
		_w11963_,
		_w11984_,
		_w21883_
	);
	LUT3 #(
		.INIT('h80)
	) name11371 (
		\wishbone_bd_ram_mem1_reg[151][11]/P0001 ,
		_w11959_,
		_w11975_,
		_w21884_
	);
	LUT3 #(
		.INIT('h80)
	) name11372 (
		\wishbone_bd_ram_mem1_reg[80][11]/P0001 ,
		_w11941_,
		_w11972_,
		_w21885_
	);
	LUT3 #(
		.INIT('h80)
	) name11373 (
		\wishbone_bd_ram_mem1_reg[83][11]/P0001 ,
		_w11938_,
		_w11972_,
		_w21886_
	);
	LUT4 #(
		.INIT('h0001)
	) name11374 (
		_w21883_,
		_w21884_,
		_w21885_,
		_w21886_,
		_w21887_
	);
	LUT3 #(
		.INIT('h80)
	) name11375 (
		\wishbone_bd_ram_mem1_reg[110][11]/P0001 ,
		_w11948_,
		_w11965_,
		_w21888_
	);
	LUT3 #(
		.INIT('h80)
	) name11376 (
		\wishbone_bd_ram_mem1_reg[239][11]/P0001 ,
		_w11973_,
		_w11982_,
		_w21889_
	);
	LUT3 #(
		.INIT('h80)
	) name11377 (
		\wishbone_bd_ram_mem1_reg[178][11]/P0001 ,
		_w11942_,
		_w11963_,
		_w21890_
	);
	LUT3 #(
		.INIT('h80)
	) name11378 (
		\wishbone_bd_ram_mem1_reg[179][11]/P0001 ,
		_w11938_,
		_w11942_,
		_w21891_
	);
	LUT4 #(
		.INIT('h0001)
	) name11379 (
		_w21888_,
		_w21889_,
		_w21890_,
		_w21891_,
		_w21892_
	);
	LUT4 #(
		.INIT('h8000)
	) name11380 (
		_w21877_,
		_w21882_,
		_w21887_,
		_w21892_,
		_w21893_
	);
	LUT3 #(
		.INIT('h80)
	) name11381 (
		\wishbone_bd_ram_mem1_reg[161][11]/P0001 ,
		_w11930_,
		_w11977_,
		_w21894_
	);
	LUT3 #(
		.INIT('h80)
	) name11382 (
		\wishbone_bd_ram_mem1_reg[224][11]/P0001 ,
		_w11941_,
		_w11982_,
		_w21895_
	);
	LUT3 #(
		.INIT('h80)
	) name11383 (
		\wishbone_bd_ram_mem1_reg[146][11]/P0001 ,
		_w11959_,
		_w11963_,
		_w21896_
	);
	LUT3 #(
		.INIT('h80)
	) name11384 (
		\wishbone_bd_ram_mem1_reg[168][11]/P0001 ,
		_w11930_,
		_w11990_,
		_w21897_
	);
	LUT4 #(
		.INIT('h0001)
	) name11385 (
		_w21894_,
		_w21895_,
		_w21896_,
		_w21897_,
		_w21898_
	);
	LUT3 #(
		.INIT('h80)
	) name11386 (
		\wishbone_bd_ram_mem1_reg[48][11]/P0001 ,
		_w11941_,
		_w11979_,
		_w21899_
	);
	LUT3 #(
		.INIT('h80)
	) name11387 (
		\wishbone_bd_ram_mem1_reg[231][11]/P0001 ,
		_w11975_,
		_w11982_,
		_w21900_
	);
	LUT3 #(
		.INIT('h80)
	) name11388 (
		\wishbone_bd_ram_mem1_reg[136][11]/P0001 ,
		_w11955_,
		_w11990_,
		_w21901_
	);
	LUT3 #(
		.INIT('h80)
	) name11389 (
		\wishbone_bd_ram_mem1_reg[127][11]/P0001 ,
		_w11973_,
		_w12012_,
		_w21902_
	);
	LUT4 #(
		.INIT('h0001)
	) name11390 (
		_w21899_,
		_w21900_,
		_w21901_,
		_w21902_,
		_w21903_
	);
	LUT3 #(
		.INIT('h80)
	) name11391 (
		\wishbone_bd_ram_mem1_reg[189][11]/P0001 ,
		_w11942_,
		_w11966_,
		_w21904_
	);
	LUT3 #(
		.INIT('h80)
	) name11392 (
		\wishbone_bd_ram_mem1_reg[237][11]/P0001 ,
		_w11966_,
		_w11982_,
		_w21905_
	);
	LUT3 #(
		.INIT('h80)
	) name11393 (
		\wishbone_bd_ram_mem1_reg[213][11]/P0001 ,
		_w11933_,
		_w11984_,
		_w21906_
	);
	LUT3 #(
		.INIT('h80)
	) name11394 (
		\wishbone_bd_ram_mem1_reg[42][11]/P0001 ,
		_w11944_,
		_w11957_,
		_w21907_
	);
	LUT4 #(
		.INIT('h0001)
	) name11395 (
		_w21904_,
		_w21905_,
		_w21906_,
		_w21907_,
		_w21908_
	);
	LUT3 #(
		.INIT('h80)
	) name11396 (
		\wishbone_bd_ram_mem1_reg[65][11]/P0001 ,
		_w11949_,
		_w11977_,
		_w21909_
	);
	LUT3 #(
		.INIT('h80)
	) name11397 (
		\wishbone_bd_ram_mem1_reg[197][11]/P0001 ,
		_w11933_,
		_w11945_,
		_w21910_
	);
	LUT3 #(
		.INIT('h80)
	) name11398 (
		\wishbone_bd_ram_mem1_reg[125][11]/P0001 ,
		_w11966_,
		_w12012_,
		_w21911_
	);
	LUT3 #(
		.INIT('h80)
	) name11399 (
		\wishbone_bd_ram_mem1_reg[202][11]/P0001 ,
		_w11944_,
		_w11945_,
		_w21912_
	);
	LUT4 #(
		.INIT('h0001)
	) name11400 (
		_w21909_,
		_w21910_,
		_w21911_,
		_w21912_,
		_w21913_
	);
	LUT4 #(
		.INIT('h8000)
	) name11401 (
		_w21898_,
		_w21903_,
		_w21908_,
		_w21913_,
		_w21914_
	);
	LUT3 #(
		.INIT('h80)
	) name11402 (
		\wishbone_bd_ram_mem1_reg[175][11]/P0001 ,
		_w11930_,
		_w11973_,
		_w21915_
	);
	LUT3 #(
		.INIT('h80)
	) name11403 (
		\wishbone_bd_ram_mem1_reg[71][11]/P0001 ,
		_w11949_,
		_w11975_,
		_w21916_
	);
	LUT3 #(
		.INIT('h80)
	) name11404 (
		\wishbone_bd_ram_mem1_reg[196][11]/P0001 ,
		_w11929_,
		_w11945_,
		_w21917_
	);
	LUT3 #(
		.INIT('h80)
	) name11405 (
		\wishbone_bd_ram_mem1_reg[119][11]/P0001 ,
		_w11975_,
		_w12012_,
		_w21918_
	);
	LUT4 #(
		.INIT('h0001)
	) name11406 (
		_w21915_,
		_w21916_,
		_w21917_,
		_w21918_,
		_w21919_
	);
	LUT3 #(
		.INIT('h80)
	) name11407 (
		\wishbone_bd_ram_mem1_reg[164][11]/P0001 ,
		_w11929_,
		_w11930_,
		_w21920_
	);
	LUT3 #(
		.INIT('h80)
	) name11408 (
		\wishbone_bd_ram_mem1_reg[78][11]/P0001 ,
		_w11948_,
		_w11949_,
		_w21921_
	);
	LUT3 #(
		.INIT('h80)
	) name11409 (
		\wishbone_bd_ram_mem1_reg[35][11]/P0001 ,
		_w11938_,
		_w11957_,
		_w21922_
	);
	LUT3 #(
		.INIT('h80)
	) name11410 (
		\wishbone_bd_ram_mem1_reg[160][11]/P0001 ,
		_w11930_,
		_w11941_,
		_w21923_
	);
	LUT4 #(
		.INIT('h0001)
	) name11411 (
		_w21920_,
		_w21921_,
		_w21922_,
		_w21923_,
		_w21924_
	);
	LUT3 #(
		.INIT('h80)
	) name11412 (
		\wishbone_bd_ram_mem1_reg[96][11]/P0001 ,
		_w11941_,
		_w11965_,
		_w21925_
	);
	LUT3 #(
		.INIT('h80)
	) name11413 (
		\wishbone_bd_ram_mem1_reg[6][11]/P0001 ,
		_w11932_,
		_w11986_,
		_w21926_
	);
	LUT3 #(
		.INIT('h80)
	) name11414 (
		\wishbone_bd_ram_mem1_reg[54][11]/P0001 ,
		_w11979_,
		_w11986_,
		_w21927_
	);
	LUT3 #(
		.INIT('h80)
	) name11415 (
		\wishbone_bd_ram_mem1_reg[194][11]/P0001 ,
		_w11945_,
		_w11963_,
		_w21928_
	);
	LUT4 #(
		.INIT('h0001)
	) name11416 (
		_w21925_,
		_w21926_,
		_w21927_,
		_w21928_,
		_w21929_
	);
	LUT3 #(
		.INIT('h80)
	) name11417 (
		\wishbone_bd_ram_mem1_reg[207][11]/P0001 ,
		_w11945_,
		_w11973_,
		_w21930_
	);
	LUT3 #(
		.INIT('h80)
	) name11418 (
		\wishbone_bd_ram_mem1_reg[32][11]/P0001 ,
		_w11941_,
		_w11957_,
		_w21931_
	);
	LUT3 #(
		.INIT('h80)
	) name11419 (
		\wishbone_bd_ram_mem1_reg[203][11]/P0001 ,
		_w11936_,
		_w11945_,
		_w21932_
	);
	LUT3 #(
		.INIT('h80)
	) name11420 (
		\wishbone_bd_ram_mem1_reg[7][11]/P0001 ,
		_w11932_,
		_w11975_,
		_w21933_
	);
	LUT4 #(
		.INIT('h0001)
	) name11421 (
		_w21930_,
		_w21931_,
		_w21932_,
		_w21933_,
		_w21934_
	);
	LUT4 #(
		.INIT('h8000)
	) name11422 (
		_w21919_,
		_w21924_,
		_w21929_,
		_w21934_,
		_w21935_
	);
	LUT3 #(
		.INIT('h80)
	) name11423 (
		\wishbone_bd_ram_mem1_reg[91][11]/P0001 ,
		_w11936_,
		_w11972_,
		_w21936_
	);
	LUT3 #(
		.INIT('h80)
	) name11424 (
		\wishbone_bd_ram_mem1_reg[44][11]/P0001 ,
		_w11954_,
		_w11957_,
		_w21937_
	);
	LUT3 #(
		.INIT('h80)
	) name11425 (
		\wishbone_bd_ram_mem1_reg[30][11]/P0001 ,
		_w11935_,
		_w11948_,
		_w21938_
	);
	LUT3 #(
		.INIT('h80)
	) name11426 (
		\wishbone_bd_ram_mem1_reg[220][11]/P0001 ,
		_w11954_,
		_w11984_,
		_w21939_
	);
	LUT4 #(
		.INIT('h0001)
	) name11427 (
		_w21936_,
		_w21937_,
		_w21938_,
		_w21939_,
		_w21940_
	);
	LUT3 #(
		.INIT('h80)
	) name11428 (
		\wishbone_bd_ram_mem1_reg[214][11]/P0001 ,
		_w11984_,
		_w11986_,
		_w21941_
	);
	LUT3 #(
		.INIT('h80)
	) name11429 (
		\wishbone_bd_ram_mem1_reg[173][11]/P0001 ,
		_w11930_,
		_w11966_,
		_w21942_
	);
	LUT3 #(
		.INIT('h80)
	) name11430 (
		\wishbone_bd_ram_mem1_reg[20][11]/P0001 ,
		_w11929_,
		_w11935_,
		_w21943_
	);
	LUT3 #(
		.INIT('h80)
	) name11431 (
		\wishbone_bd_ram_mem1_reg[40][11]/P0001 ,
		_w11957_,
		_w11990_,
		_w21944_
	);
	LUT4 #(
		.INIT('h0001)
	) name11432 (
		_w21941_,
		_w21942_,
		_w21943_,
		_w21944_,
		_w21945_
	);
	LUT3 #(
		.INIT('h80)
	) name11433 (
		\wishbone_bd_ram_mem1_reg[181][11]/P0001 ,
		_w11933_,
		_w11942_,
		_w21946_
	);
	LUT3 #(
		.INIT('h80)
	) name11434 (
		\wishbone_bd_ram_mem1_reg[26][11]/P0001 ,
		_w11935_,
		_w11944_,
		_w21947_
	);
	LUT3 #(
		.INIT('h80)
	) name11435 (
		\wishbone_bd_ram_mem1_reg[147][11]/P0001 ,
		_w11938_,
		_w11959_,
		_w21948_
	);
	LUT3 #(
		.INIT('h80)
	) name11436 (
		\wishbone_bd_ram_mem1_reg[211][11]/P0001 ,
		_w11938_,
		_w11984_,
		_w21949_
	);
	LUT4 #(
		.INIT('h0001)
	) name11437 (
		_w21946_,
		_w21947_,
		_w21948_,
		_w21949_,
		_w21950_
	);
	LUT3 #(
		.INIT('h80)
	) name11438 (
		\wishbone_bd_ram_mem1_reg[75][11]/P0001 ,
		_w11936_,
		_w11949_,
		_w21951_
	);
	LUT3 #(
		.INIT('h80)
	) name11439 (
		\wishbone_bd_ram_mem1_reg[10][11]/P0001 ,
		_w11932_,
		_w11944_,
		_w21952_
	);
	LUT3 #(
		.INIT('h80)
	) name11440 (
		\wishbone_bd_ram_mem1_reg[12][11]/P0001 ,
		_w11932_,
		_w11954_,
		_w21953_
	);
	LUT3 #(
		.INIT('h80)
	) name11441 (
		\wishbone_bd_ram_mem1_reg[61][11]/P0001 ,
		_w11966_,
		_w11979_,
		_w21954_
	);
	LUT4 #(
		.INIT('h0001)
	) name11442 (
		_w21951_,
		_w21952_,
		_w21953_,
		_w21954_,
		_w21955_
	);
	LUT4 #(
		.INIT('h8000)
	) name11443 (
		_w21940_,
		_w21945_,
		_w21950_,
		_w21955_,
		_w21956_
	);
	LUT4 #(
		.INIT('h8000)
	) name11444 (
		_w21893_,
		_w21914_,
		_w21935_,
		_w21956_,
		_w21957_
	);
	LUT3 #(
		.INIT('h80)
	) name11445 (
		\wishbone_bd_ram_mem1_reg[121][11]/P0001 ,
		_w11968_,
		_w12012_,
		_w21958_
	);
	LUT3 #(
		.INIT('h80)
	) name11446 (
		\wishbone_bd_ram_mem1_reg[176][11]/P0001 ,
		_w11941_,
		_w11942_,
		_w21959_
	);
	LUT3 #(
		.INIT('h80)
	) name11447 (
		\wishbone_bd_ram_mem1_reg[242][11]/P0001 ,
		_w11952_,
		_w11963_,
		_w21960_
	);
	LUT3 #(
		.INIT('h80)
	) name11448 (
		\wishbone_bd_ram_mem1_reg[79][11]/P0001 ,
		_w11949_,
		_w11973_,
		_w21961_
	);
	LUT4 #(
		.INIT('h0001)
	) name11449 (
		_w21958_,
		_w21959_,
		_w21960_,
		_w21961_,
		_w21962_
	);
	LUT3 #(
		.INIT('h80)
	) name11450 (
		\wishbone_bd_ram_mem1_reg[182][11]/P0001 ,
		_w11942_,
		_w11986_,
		_w21963_
	);
	LUT3 #(
		.INIT('h80)
	) name11451 (
		\wishbone_bd_ram_mem1_reg[74][11]/P0001 ,
		_w11944_,
		_w11949_,
		_w21964_
	);
	LUT3 #(
		.INIT('h80)
	) name11452 (
		\wishbone_bd_ram_mem1_reg[131][11]/P0001 ,
		_w11938_,
		_w11955_,
		_w21965_
	);
	LUT3 #(
		.INIT('h80)
	) name11453 (
		\wishbone_bd_ram_mem1_reg[38][11]/P0001 ,
		_w11957_,
		_w11986_,
		_w21966_
	);
	LUT4 #(
		.INIT('h0001)
	) name11454 (
		_w21963_,
		_w21964_,
		_w21965_,
		_w21966_,
		_w21967_
	);
	LUT3 #(
		.INIT('h80)
	) name11455 (
		\wishbone_bd_ram_mem1_reg[221][11]/P0001 ,
		_w11966_,
		_w11984_,
		_w21968_
	);
	LUT3 #(
		.INIT('h80)
	) name11456 (
		\wishbone_bd_ram_mem1_reg[218][11]/P0001 ,
		_w11944_,
		_w11984_,
		_w21969_
	);
	LUT3 #(
		.INIT('h80)
	) name11457 (
		\wishbone_bd_ram_mem1_reg[162][11]/P0001 ,
		_w11930_,
		_w11963_,
		_w21970_
	);
	LUT3 #(
		.INIT('h80)
	) name11458 (
		\wishbone_bd_ram_mem1_reg[21][11]/P0001 ,
		_w11933_,
		_w11935_,
		_w21971_
	);
	LUT4 #(
		.INIT('h0001)
	) name11459 (
		_w21968_,
		_w21969_,
		_w21970_,
		_w21971_,
		_w21972_
	);
	LUT3 #(
		.INIT('h80)
	) name11460 (
		\wishbone_bd_ram_mem1_reg[245][11]/P0001 ,
		_w11933_,
		_w11952_,
		_w21973_
	);
	LUT3 #(
		.INIT('h80)
	) name11461 (
		\wishbone_bd_ram_mem1_reg[56][11]/P0001 ,
		_w11979_,
		_w11990_,
		_w21974_
	);
	LUT3 #(
		.INIT('h80)
	) name11462 (
		\wishbone_bd_ram_mem1_reg[183][11]/P0001 ,
		_w11942_,
		_w11975_,
		_w21975_
	);
	LUT3 #(
		.INIT('h80)
	) name11463 (
		\wishbone_bd_ram_mem1_reg[124][11]/P0001 ,
		_w11954_,
		_w12012_,
		_w21976_
	);
	LUT4 #(
		.INIT('h0001)
	) name11464 (
		_w21973_,
		_w21974_,
		_w21975_,
		_w21976_,
		_w21977_
	);
	LUT4 #(
		.INIT('h8000)
	) name11465 (
		_w21962_,
		_w21967_,
		_w21972_,
		_w21977_,
		_w21978_
	);
	LUT3 #(
		.INIT('h80)
	) name11466 (
		\wishbone_bd_ram_mem1_reg[64][11]/P0001 ,
		_w11941_,
		_w11949_,
		_w21979_
	);
	LUT3 #(
		.INIT('h80)
	) name11467 (
		\wishbone_bd_ram_mem1_reg[95][11]/P0001 ,
		_w11972_,
		_w11973_,
		_w21980_
	);
	LUT3 #(
		.INIT('h80)
	) name11468 (
		\wishbone_bd_ram_mem1_reg[68][11]/P0001 ,
		_w11929_,
		_w11949_,
		_w21981_
	);
	LUT3 #(
		.INIT('h80)
	) name11469 (
		\wishbone_bd_ram_mem1_reg[46][11]/P0001 ,
		_w11948_,
		_w11957_,
		_w21982_
	);
	LUT4 #(
		.INIT('h0001)
	) name11470 (
		_w21979_,
		_w21980_,
		_w21981_,
		_w21982_,
		_w21983_
	);
	LUT3 #(
		.INIT('h80)
	) name11471 (
		\wishbone_bd_ram_mem1_reg[69][11]/P0001 ,
		_w11933_,
		_w11949_,
		_w21984_
	);
	LUT3 #(
		.INIT('h80)
	) name11472 (
		\wishbone_bd_ram_mem1_reg[157][11]/P0001 ,
		_w11959_,
		_w11966_,
		_w21985_
	);
	LUT3 #(
		.INIT('h80)
	) name11473 (
		\wishbone_bd_ram_mem1_reg[106][11]/P0001 ,
		_w11944_,
		_w11965_,
		_w21986_
	);
	LUT3 #(
		.INIT('h80)
	) name11474 (
		\wishbone_bd_ram_mem1_reg[177][11]/P0001 ,
		_w11942_,
		_w11977_,
		_w21987_
	);
	LUT4 #(
		.INIT('h0001)
	) name11475 (
		_w21984_,
		_w21985_,
		_w21986_,
		_w21987_,
		_w21988_
	);
	LUT3 #(
		.INIT('h80)
	) name11476 (
		\wishbone_bd_ram_mem1_reg[27][11]/P0001 ,
		_w11935_,
		_w11936_,
		_w21989_
	);
	LUT3 #(
		.INIT('h80)
	) name11477 (
		\wishbone_bd_ram_mem1_reg[190][11]/P0001 ,
		_w11942_,
		_w11948_,
		_w21990_
	);
	LUT3 #(
		.INIT('h80)
	) name11478 (
		\wishbone_bd_ram_mem1_reg[107][11]/P0001 ,
		_w11936_,
		_w11965_,
		_w21991_
	);
	LUT3 #(
		.INIT('h80)
	) name11479 (
		\wishbone_bd_ram_mem1_reg[36][11]/P0001 ,
		_w11929_,
		_w11957_,
		_w21992_
	);
	LUT4 #(
		.INIT('h0001)
	) name11480 (
		_w21989_,
		_w21990_,
		_w21991_,
		_w21992_,
		_w21993_
	);
	LUT3 #(
		.INIT('h80)
	) name11481 (
		\wishbone_bd_ram_mem1_reg[118][11]/P0001 ,
		_w11986_,
		_w12012_,
		_w21994_
	);
	LUT3 #(
		.INIT('h80)
	) name11482 (
		\wishbone_bd_ram_mem1_reg[28][11]/P0001 ,
		_w11935_,
		_w11954_,
		_w21995_
	);
	LUT3 #(
		.INIT('h80)
	) name11483 (
		\wishbone_bd_ram_mem1_reg[171][11]/P0001 ,
		_w11930_,
		_w11936_,
		_w21996_
	);
	LUT3 #(
		.INIT('h80)
	) name11484 (
		\wishbone_bd_ram_mem1_reg[163][11]/P0001 ,
		_w11930_,
		_w11938_,
		_w21997_
	);
	LUT4 #(
		.INIT('h0001)
	) name11485 (
		_w21994_,
		_w21995_,
		_w21996_,
		_w21997_,
		_w21998_
	);
	LUT4 #(
		.INIT('h8000)
	) name11486 (
		_w21983_,
		_w21988_,
		_w21993_,
		_w21998_,
		_w21999_
	);
	LUT3 #(
		.INIT('h80)
	) name11487 (
		\wishbone_bd_ram_mem1_reg[246][11]/P0001 ,
		_w11952_,
		_w11986_,
		_w22000_
	);
	LUT3 #(
		.INIT('h80)
	) name11488 (
		\wishbone_bd_ram_mem1_reg[122][11]/P0001 ,
		_w11944_,
		_w12012_,
		_w22001_
	);
	LUT3 #(
		.INIT('h80)
	) name11489 (
		\wishbone_bd_ram_mem1_reg[174][11]/P0001 ,
		_w11930_,
		_w11948_,
		_w22002_
	);
	LUT3 #(
		.INIT('h80)
	) name11490 (
		\wishbone_bd_ram_mem1_reg[180][11]/P0001 ,
		_w11929_,
		_w11942_,
		_w22003_
	);
	LUT4 #(
		.INIT('h0001)
	) name11491 (
		_w22000_,
		_w22001_,
		_w22002_,
		_w22003_,
		_w22004_
	);
	LUT3 #(
		.INIT('h80)
	) name11492 (
		\wishbone_bd_ram_mem1_reg[8][11]/P0001 ,
		_w11932_,
		_w11990_,
		_w22005_
	);
	LUT3 #(
		.INIT('h80)
	) name11493 (
		\wishbone_bd_ram_mem1_reg[234][11]/P0001 ,
		_w11944_,
		_w11982_,
		_w22006_
	);
	LUT3 #(
		.INIT('h80)
	) name11494 (
		\wishbone_bd_ram_mem1_reg[148][11]/P0001 ,
		_w11929_,
		_w11959_,
		_w22007_
	);
	LUT3 #(
		.INIT('h80)
	) name11495 (
		\wishbone_bd_ram_mem1_reg[98][11]/P0001 ,
		_w11963_,
		_w11965_,
		_w22008_
	);
	LUT4 #(
		.INIT('h0001)
	) name11496 (
		_w22005_,
		_w22006_,
		_w22007_,
		_w22008_,
		_w22009_
	);
	LUT3 #(
		.INIT('h80)
	) name11497 (
		\wishbone_bd_ram_mem1_reg[222][11]/P0001 ,
		_w11948_,
		_w11984_,
		_w22010_
	);
	LUT3 #(
		.INIT('h80)
	) name11498 (
		\wishbone_bd_ram_mem1_reg[191][11]/P0001 ,
		_w11942_,
		_w11973_,
		_w22011_
	);
	LUT3 #(
		.INIT('h80)
	) name11499 (
		\wishbone_bd_ram_mem1_reg[99][11]/P0001 ,
		_w11938_,
		_w11965_,
		_w22012_
	);
	LUT3 #(
		.INIT('h80)
	) name11500 (
		\wishbone_bd_ram_mem1_reg[192][11]/P0001 ,
		_w11941_,
		_w11945_,
		_w22013_
	);
	LUT4 #(
		.INIT('h0001)
	) name11501 (
		_w22010_,
		_w22011_,
		_w22012_,
		_w22013_,
		_w22014_
	);
	LUT3 #(
		.INIT('h80)
	) name11502 (
		\wishbone_bd_ram_mem1_reg[90][11]/P0001 ,
		_w11944_,
		_w11972_,
		_w22015_
	);
	LUT3 #(
		.INIT('h80)
	) name11503 (
		\wishbone_bd_ram_mem1_reg[206][11]/P0001 ,
		_w11945_,
		_w11948_,
		_w22016_
	);
	LUT3 #(
		.INIT('h80)
	) name11504 (
		\wishbone_bd_ram_mem1_reg[82][11]/P0001 ,
		_w11963_,
		_w11972_,
		_w22017_
	);
	LUT3 #(
		.INIT('h80)
	) name11505 (
		\wishbone_bd_ram_mem1_reg[111][11]/P0001 ,
		_w11965_,
		_w11973_,
		_w22018_
	);
	LUT4 #(
		.INIT('h0001)
	) name11506 (
		_w22015_,
		_w22016_,
		_w22017_,
		_w22018_,
		_w22019_
	);
	LUT4 #(
		.INIT('h8000)
	) name11507 (
		_w22004_,
		_w22009_,
		_w22014_,
		_w22019_,
		_w22020_
	);
	LUT3 #(
		.INIT('h80)
	) name11508 (
		\wishbone_bd_ram_mem1_reg[62][11]/P0001 ,
		_w11948_,
		_w11979_,
		_w22021_
	);
	LUT3 #(
		.INIT('h80)
	) name11509 (
		\wishbone_bd_ram_mem1_reg[134][11]/P0001 ,
		_w11955_,
		_w11986_,
		_w22022_
	);
	LUT3 #(
		.INIT('h80)
	) name11510 (
		\wishbone_bd_ram_mem1_reg[184][11]/P0001 ,
		_w11942_,
		_w11990_,
		_w22023_
	);
	LUT3 #(
		.INIT('h80)
	) name11511 (
		\wishbone_bd_ram_mem1_reg[219][11]/P0001 ,
		_w11936_,
		_w11984_,
		_w22024_
	);
	LUT4 #(
		.INIT('h0001)
	) name11512 (
		_w22021_,
		_w22022_,
		_w22023_,
		_w22024_,
		_w22025_
	);
	LUT3 #(
		.INIT('h80)
	) name11513 (
		\wishbone_bd_ram_mem1_reg[123][11]/P0001 ,
		_w11936_,
		_w12012_,
		_w22026_
	);
	LUT3 #(
		.INIT('h80)
	) name11514 (
		\wishbone_bd_ram_mem1_reg[217][11]/P0001 ,
		_w11968_,
		_w11984_,
		_w22027_
	);
	LUT3 #(
		.INIT('h80)
	) name11515 (
		\wishbone_bd_ram_mem1_reg[250][11]/P0001 ,
		_w11944_,
		_w11952_,
		_w22028_
	);
	LUT3 #(
		.INIT('h80)
	) name11516 (
		\wishbone_bd_ram_mem1_reg[154][11]/P0001 ,
		_w11944_,
		_w11959_,
		_w22029_
	);
	LUT4 #(
		.INIT('h0001)
	) name11517 (
		_w22026_,
		_w22027_,
		_w22028_,
		_w22029_,
		_w22030_
	);
	LUT3 #(
		.INIT('h80)
	) name11518 (
		\wishbone_bd_ram_mem1_reg[185][11]/P0001 ,
		_w11942_,
		_w11968_,
		_w22031_
	);
	LUT3 #(
		.INIT('h80)
	) name11519 (
		\wishbone_bd_ram_mem1_reg[232][11]/P0001 ,
		_w11982_,
		_w11990_,
		_w22032_
	);
	LUT3 #(
		.INIT('h80)
	) name11520 (
		\wishbone_bd_ram_mem1_reg[55][11]/P0001 ,
		_w11975_,
		_w11979_,
		_w22033_
	);
	LUT3 #(
		.INIT('h80)
	) name11521 (
		\wishbone_bd_ram_mem1_reg[101][11]/P0001 ,
		_w11933_,
		_w11965_,
		_w22034_
	);
	LUT4 #(
		.INIT('h0001)
	) name11522 (
		_w22031_,
		_w22032_,
		_w22033_,
		_w22034_,
		_w22035_
	);
	LUT3 #(
		.INIT('h80)
	) name11523 (
		\wishbone_bd_ram_mem1_reg[33][11]/P0001 ,
		_w11957_,
		_w11977_,
		_w22036_
	);
	LUT3 #(
		.INIT('h80)
	) name11524 (
		\wishbone_bd_ram_mem1_reg[253][11]/P0001 ,
		_w11952_,
		_w11966_,
		_w22037_
	);
	LUT3 #(
		.INIT('h80)
	) name11525 (
		\wishbone_bd_ram_mem1_reg[113][11]/P0001 ,
		_w11977_,
		_w12012_,
		_w22038_
	);
	LUT3 #(
		.INIT('h80)
	) name11526 (
		\wishbone_bd_ram_mem1_reg[153][11]/P0001 ,
		_w11959_,
		_w11968_,
		_w22039_
	);
	LUT4 #(
		.INIT('h0001)
	) name11527 (
		_w22036_,
		_w22037_,
		_w22038_,
		_w22039_,
		_w22040_
	);
	LUT4 #(
		.INIT('h8000)
	) name11528 (
		_w22025_,
		_w22030_,
		_w22035_,
		_w22040_,
		_w22041_
	);
	LUT4 #(
		.INIT('h8000)
	) name11529 (
		_w21978_,
		_w21999_,
		_w22020_,
		_w22041_,
		_w22042_
	);
	LUT3 #(
		.INIT('h80)
	) name11530 (
		\wishbone_bd_ram_mem1_reg[103][11]/P0001 ,
		_w11965_,
		_w11975_,
		_w22043_
	);
	LUT3 #(
		.INIT('h80)
	) name11531 (
		\wishbone_bd_ram_mem1_reg[205][11]/P0001 ,
		_w11945_,
		_w11966_,
		_w22044_
	);
	LUT3 #(
		.INIT('h80)
	) name11532 (
		\wishbone_bd_ram_mem1_reg[132][11]/P0001 ,
		_w11929_,
		_w11955_,
		_w22045_
	);
	LUT3 #(
		.INIT('h80)
	) name11533 (
		\wishbone_bd_ram_mem1_reg[247][11]/P0001 ,
		_w11952_,
		_w11975_,
		_w22046_
	);
	LUT4 #(
		.INIT('h0001)
	) name11534 (
		_w22043_,
		_w22044_,
		_w22045_,
		_w22046_,
		_w22047_
	);
	LUT3 #(
		.INIT('h80)
	) name11535 (
		\wishbone_bd_ram_mem1_reg[200][11]/P0001 ,
		_w11945_,
		_w11990_,
		_w22048_
	);
	LUT3 #(
		.INIT('h80)
	) name11536 (
		\wishbone_bd_ram_mem1_reg[114][11]/P0001 ,
		_w11963_,
		_w12012_,
		_w22049_
	);
	LUT3 #(
		.INIT('h80)
	) name11537 (
		\wishbone_bd_ram_mem1_reg[252][11]/P0001 ,
		_w11952_,
		_w11954_,
		_w22050_
	);
	LUT3 #(
		.INIT('h80)
	) name11538 (
		\wishbone_bd_ram_mem1_reg[201][11]/P0001 ,
		_w11945_,
		_w11968_,
		_w22051_
	);
	LUT4 #(
		.INIT('h0001)
	) name11539 (
		_w22048_,
		_w22049_,
		_w22050_,
		_w22051_,
		_w22052_
	);
	LUT3 #(
		.INIT('h80)
	) name11540 (
		\wishbone_bd_ram_mem1_reg[236][11]/P0001 ,
		_w11954_,
		_w11982_,
		_w22053_
	);
	LUT3 #(
		.INIT('h80)
	) name11541 (
		\wishbone_bd_ram_mem1_reg[2][11]/P0001 ,
		_w11932_,
		_w11963_,
		_w22054_
	);
	LUT3 #(
		.INIT('h80)
	) name11542 (
		\wishbone_bd_ram_mem1_reg[199][11]/P0001 ,
		_w11945_,
		_w11975_,
		_w22055_
	);
	LUT3 #(
		.INIT('h80)
	) name11543 (
		\wishbone_bd_ram_mem1_reg[81][11]/P0001 ,
		_w11972_,
		_w11977_,
		_w22056_
	);
	LUT4 #(
		.INIT('h0001)
	) name11544 (
		_w22053_,
		_w22054_,
		_w22055_,
		_w22056_,
		_w22057_
	);
	LUT3 #(
		.INIT('h80)
	) name11545 (
		\wishbone_bd_ram_mem1_reg[241][11]/P0001 ,
		_w11952_,
		_w11977_,
		_w22058_
	);
	LUT3 #(
		.INIT('h80)
	) name11546 (
		\wishbone_bd_ram_mem1_reg[141][11]/P0001 ,
		_w11955_,
		_w11966_,
		_w22059_
	);
	LUT3 #(
		.INIT('h80)
	) name11547 (
		\wishbone_bd_ram_mem1_reg[51][11]/P0001 ,
		_w11938_,
		_w11979_,
		_w22060_
	);
	LUT3 #(
		.INIT('h80)
	) name11548 (
		\wishbone_bd_ram_mem1_reg[129][11]/P0001 ,
		_w11955_,
		_w11977_,
		_w22061_
	);
	LUT4 #(
		.INIT('h0001)
	) name11549 (
		_w22058_,
		_w22059_,
		_w22060_,
		_w22061_,
		_w22062_
	);
	LUT4 #(
		.INIT('h8000)
	) name11550 (
		_w22047_,
		_w22052_,
		_w22057_,
		_w22062_,
		_w22063_
	);
	LUT3 #(
		.INIT('h80)
	) name11551 (
		\wishbone_bd_ram_mem1_reg[14][11]/P0001 ,
		_w11932_,
		_w11948_,
		_w22064_
	);
	LUT3 #(
		.INIT('h80)
	) name11552 (
		\wishbone_bd_ram_mem1_reg[128][11]/P0001 ,
		_w11941_,
		_w11955_,
		_w22065_
	);
	LUT3 #(
		.INIT('h80)
	) name11553 (
		\wishbone_bd_ram_mem1_reg[144][11]/P0001 ,
		_w11941_,
		_w11959_,
		_w22066_
	);
	LUT3 #(
		.INIT('h80)
	) name11554 (
		\wishbone_bd_ram_mem1_reg[170][11]/P0001 ,
		_w11930_,
		_w11944_,
		_w22067_
	);
	LUT4 #(
		.INIT('h0001)
	) name11555 (
		_w22064_,
		_w22065_,
		_w22066_,
		_w22067_,
		_w22068_
	);
	LUT3 #(
		.INIT('h80)
	) name11556 (
		\wishbone_bd_ram_mem1_reg[150][11]/P0001 ,
		_w11959_,
		_w11986_,
		_w22069_
	);
	LUT3 #(
		.INIT('h80)
	) name11557 (
		\wishbone_bd_ram_mem1_reg[216][11]/P0001 ,
		_w11984_,
		_w11990_,
		_w22070_
	);
	LUT3 #(
		.INIT('h80)
	) name11558 (
		\wishbone_bd_ram_mem1_reg[208][11]/P0001 ,
		_w11941_,
		_w11984_,
		_w22071_
	);
	LUT3 #(
		.INIT('h80)
	) name11559 (
		\wishbone_bd_ram_mem1_reg[115][11]/P0001 ,
		_w11938_,
		_w12012_,
		_w22072_
	);
	LUT4 #(
		.INIT('h0001)
	) name11560 (
		_w22069_,
		_w22070_,
		_w22071_,
		_w22072_,
		_w22073_
	);
	LUT3 #(
		.INIT('h80)
	) name11561 (
		\wishbone_bd_ram_mem1_reg[49][11]/P0001 ,
		_w11977_,
		_w11979_,
		_w22074_
	);
	LUT3 #(
		.INIT('h80)
	) name11562 (
		\wishbone_bd_ram_mem1_reg[104][11]/P0001 ,
		_w11965_,
		_w11990_,
		_w22075_
	);
	LUT3 #(
		.INIT('h80)
	) name11563 (
		\wishbone_bd_ram_mem1_reg[76][11]/P0001 ,
		_w11949_,
		_w11954_,
		_w22076_
	);
	LUT3 #(
		.INIT('h80)
	) name11564 (
		\wishbone_bd_ram_mem1_reg[73][11]/P0001 ,
		_w11949_,
		_w11968_,
		_w22077_
	);
	LUT4 #(
		.INIT('h0001)
	) name11565 (
		_w22074_,
		_w22075_,
		_w22076_,
		_w22077_,
		_w22078_
	);
	LUT3 #(
		.INIT('h80)
	) name11566 (
		\wishbone_bd_ram_mem1_reg[186][11]/P0001 ,
		_w11942_,
		_w11944_,
		_w22079_
	);
	LUT3 #(
		.INIT('h80)
	) name11567 (
		\wishbone_bd_ram_mem1_reg[25][11]/P0001 ,
		_w11935_,
		_w11968_,
		_w22080_
	);
	LUT3 #(
		.INIT('h80)
	) name11568 (
		\wishbone_bd_ram_mem1_reg[188][11]/P0001 ,
		_w11942_,
		_w11954_,
		_w22081_
	);
	LUT3 #(
		.INIT('h80)
	) name11569 (
		\wishbone_bd_ram_mem1_reg[172][11]/P0001 ,
		_w11930_,
		_w11954_,
		_w22082_
	);
	LUT4 #(
		.INIT('h0001)
	) name11570 (
		_w22079_,
		_w22080_,
		_w22081_,
		_w22082_,
		_w22083_
	);
	LUT4 #(
		.INIT('h8000)
	) name11571 (
		_w22068_,
		_w22073_,
		_w22078_,
		_w22083_,
		_w22084_
	);
	LUT3 #(
		.INIT('h80)
	) name11572 (
		\wishbone_bd_ram_mem1_reg[215][11]/P0001 ,
		_w11975_,
		_w11984_,
		_w22085_
	);
	LUT3 #(
		.INIT('h80)
	) name11573 (
		\wishbone_bd_ram_mem1_reg[93][11]/P0001 ,
		_w11966_,
		_w11972_,
		_w22086_
	);
	LUT3 #(
		.INIT('h80)
	) name11574 (
		\wishbone_bd_ram_mem1_reg[120][11]/P0001 ,
		_w11990_,
		_w12012_,
		_w22087_
	);
	LUT3 #(
		.INIT('h80)
	) name11575 (
		\wishbone_bd_ram_mem1_reg[212][11]/P0001 ,
		_w11929_,
		_w11984_,
		_w22088_
	);
	LUT4 #(
		.INIT('h0001)
	) name11576 (
		_w22085_,
		_w22086_,
		_w22087_,
		_w22088_,
		_w22089_
	);
	LUT3 #(
		.INIT('h80)
	) name11577 (
		\wishbone_bd_ram_mem1_reg[227][11]/P0001 ,
		_w11938_,
		_w11982_,
		_w22090_
	);
	LUT3 #(
		.INIT('h80)
	) name11578 (
		\wishbone_bd_ram_mem1_reg[255][11]/P0001 ,
		_w11952_,
		_w11973_,
		_w22091_
	);
	LUT3 #(
		.INIT('h80)
	) name11579 (
		\wishbone_bd_ram_mem1_reg[53][11]/P0001 ,
		_w11933_,
		_w11979_,
		_w22092_
	);
	LUT3 #(
		.INIT('h80)
	) name11580 (
		\wishbone_bd_ram_mem1_reg[169][11]/P0001 ,
		_w11930_,
		_w11968_,
		_w22093_
	);
	LUT4 #(
		.INIT('h0001)
	) name11581 (
		_w22090_,
		_w22091_,
		_w22092_,
		_w22093_,
		_w22094_
	);
	LUT3 #(
		.INIT('h80)
	) name11582 (
		\wishbone_bd_ram_mem1_reg[72][11]/P0001 ,
		_w11949_,
		_w11990_,
		_w22095_
	);
	LUT3 #(
		.INIT('h80)
	) name11583 (
		\wishbone_bd_ram_mem1_reg[66][11]/P0001 ,
		_w11949_,
		_w11963_,
		_w22096_
	);
	LUT3 #(
		.INIT('h80)
	) name11584 (
		\wishbone_bd_ram_mem1_reg[108][11]/P0001 ,
		_w11954_,
		_w11965_,
		_w22097_
	);
	LUT3 #(
		.INIT('h80)
	) name11585 (
		\wishbone_bd_ram_mem1_reg[243][11]/P0001 ,
		_w11938_,
		_w11952_,
		_w22098_
	);
	LUT4 #(
		.INIT('h0001)
	) name11586 (
		_w22095_,
		_w22096_,
		_w22097_,
		_w22098_,
		_w22099_
	);
	LUT3 #(
		.INIT('h80)
	) name11587 (
		\wishbone_bd_ram_mem1_reg[47][11]/P0001 ,
		_w11957_,
		_w11973_,
		_w22100_
	);
	LUT3 #(
		.INIT('h80)
	) name11588 (
		\wishbone_bd_ram_mem1_reg[117][11]/P0001 ,
		_w11933_,
		_w12012_,
		_w22101_
	);
	LUT3 #(
		.INIT('h80)
	) name11589 (
		\wishbone_bd_ram_mem1_reg[112][11]/P0001 ,
		_w11941_,
		_w12012_,
		_w22102_
	);
	LUT3 #(
		.INIT('h80)
	) name11590 (
		\wishbone_bd_ram_mem1_reg[87][11]/P0001 ,
		_w11972_,
		_w11975_,
		_w22103_
	);
	LUT4 #(
		.INIT('h0001)
	) name11591 (
		_w22100_,
		_w22101_,
		_w22102_,
		_w22103_,
		_w22104_
	);
	LUT4 #(
		.INIT('h8000)
	) name11592 (
		_w22089_,
		_w22094_,
		_w22099_,
		_w22104_,
		_w22105_
	);
	LUT3 #(
		.INIT('h80)
	) name11593 (
		\wishbone_bd_ram_mem1_reg[223][11]/P0001 ,
		_w11973_,
		_w11984_,
		_w22106_
	);
	LUT3 #(
		.INIT('h80)
	) name11594 (
		\wishbone_bd_ram_mem1_reg[43][11]/P0001 ,
		_w11936_,
		_w11957_,
		_w22107_
	);
	LUT3 #(
		.INIT('h80)
	) name11595 (
		\wishbone_bd_ram_mem1_reg[233][11]/P0001 ,
		_w11968_,
		_w11982_,
		_w22108_
	);
	LUT3 #(
		.INIT('h80)
	) name11596 (
		\wishbone_bd_ram_mem1_reg[152][11]/P0001 ,
		_w11959_,
		_w11990_,
		_w22109_
	);
	LUT4 #(
		.INIT('h0001)
	) name11597 (
		_w22106_,
		_w22107_,
		_w22108_,
		_w22109_,
		_w22110_
	);
	LUT3 #(
		.INIT('h80)
	) name11598 (
		\wishbone_bd_ram_mem1_reg[67][11]/P0001 ,
		_w11938_,
		_w11949_,
		_w22111_
	);
	LUT3 #(
		.INIT('h80)
	) name11599 (
		\wishbone_bd_ram_mem1_reg[9][11]/P0001 ,
		_w11932_,
		_w11968_,
		_w22112_
	);
	LUT3 #(
		.INIT('h80)
	) name11600 (
		\wishbone_bd_ram_mem1_reg[100][11]/P0001 ,
		_w11929_,
		_w11965_,
		_w22113_
	);
	LUT3 #(
		.INIT('h80)
	) name11601 (
		\wishbone_bd_ram_mem1_reg[0][11]/P0001 ,
		_w11932_,
		_w11941_,
		_w22114_
	);
	LUT4 #(
		.INIT('h0001)
	) name11602 (
		_w22111_,
		_w22112_,
		_w22113_,
		_w22114_,
		_w22115_
	);
	LUT3 #(
		.INIT('h80)
	) name11603 (
		\wishbone_bd_ram_mem1_reg[41][11]/P0001 ,
		_w11957_,
		_w11968_,
		_w22116_
	);
	LUT3 #(
		.INIT('h80)
	) name11604 (
		\wishbone_bd_ram_mem1_reg[89][11]/P0001 ,
		_w11968_,
		_w11972_,
		_w22117_
	);
	LUT3 #(
		.INIT('h80)
	) name11605 (
		\wishbone_bd_ram_mem1_reg[45][11]/P0001 ,
		_w11957_,
		_w11966_,
		_w22118_
	);
	LUT3 #(
		.INIT('h80)
	) name11606 (
		\wishbone_bd_ram_mem1_reg[248][11]/P0001 ,
		_w11952_,
		_w11990_,
		_w22119_
	);
	LUT4 #(
		.INIT('h0001)
	) name11607 (
		_w22116_,
		_w22117_,
		_w22118_,
		_w22119_,
		_w22120_
	);
	LUT3 #(
		.INIT('h80)
	) name11608 (
		\wishbone_bd_ram_mem1_reg[109][11]/P0001 ,
		_w11965_,
		_w11966_,
		_w22121_
	);
	LUT3 #(
		.INIT('h80)
	) name11609 (
		\wishbone_bd_ram_mem1_reg[88][11]/P0001 ,
		_w11972_,
		_w11990_,
		_w22122_
	);
	LUT3 #(
		.INIT('h80)
	) name11610 (
		\wishbone_bd_ram_mem1_reg[3][11]/P0001 ,
		_w11932_,
		_w11938_,
		_w22123_
	);
	LUT3 #(
		.INIT('h80)
	) name11611 (
		\wishbone_bd_ram_mem1_reg[17][11]/P0001 ,
		_w11935_,
		_w11977_,
		_w22124_
	);
	LUT4 #(
		.INIT('h0001)
	) name11612 (
		_w22121_,
		_w22122_,
		_w22123_,
		_w22124_,
		_w22125_
	);
	LUT4 #(
		.INIT('h8000)
	) name11613 (
		_w22110_,
		_w22115_,
		_w22120_,
		_w22125_,
		_w22126_
	);
	LUT4 #(
		.INIT('h8000)
	) name11614 (
		_w22063_,
		_w22084_,
		_w22105_,
		_w22126_,
		_w22127_
	);
	LUT3 #(
		.INIT('h80)
	) name11615 (
		\wishbone_bd_ram_mem1_reg[37][11]/P0001 ,
		_w11933_,
		_w11957_,
		_w22128_
	);
	LUT3 #(
		.INIT('h80)
	) name11616 (
		\wishbone_bd_ram_mem1_reg[167][11]/P0001 ,
		_w11930_,
		_w11975_,
		_w22129_
	);
	LUT3 #(
		.INIT('h80)
	) name11617 (
		\wishbone_bd_ram_mem1_reg[254][11]/P0001 ,
		_w11948_,
		_w11952_,
		_w22130_
	);
	LUT3 #(
		.INIT('h80)
	) name11618 (
		\wishbone_bd_ram_mem1_reg[198][11]/P0001 ,
		_w11945_,
		_w11986_,
		_w22131_
	);
	LUT4 #(
		.INIT('h0001)
	) name11619 (
		_w22128_,
		_w22129_,
		_w22130_,
		_w22131_,
		_w22132_
	);
	LUT3 #(
		.INIT('h80)
	) name11620 (
		\wishbone_bd_ram_mem1_reg[50][11]/P0001 ,
		_w11963_,
		_w11979_,
		_w22133_
	);
	LUT3 #(
		.INIT('h80)
	) name11621 (
		\wishbone_bd_ram_mem1_reg[229][11]/P0001 ,
		_w11933_,
		_w11982_,
		_w22134_
	);
	LUT3 #(
		.INIT('h80)
	) name11622 (
		\wishbone_bd_ram_mem1_reg[130][11]/P0001 ,
		_w11955_,
		_w11963_,
		_w22135_
	);
	LUT3 #(
		.INIT('h80)
	) name11623 (
		\wishbone_bd_ram_mem1_reg[187][11]/P0001 ,
		_w11936_,
		_w11942_,
		_w22136_
	);
	LUT4 #(
		.INIT('h0001)
	) name11624 (
		_w22133_,
		_w22134_,
		_w22135_,
		_w22136_,
		_w22137_
	);
	LUT3 #(
		.INIT('h80)
	) name11625 (
		\wishbone_bd_ram_mem1_reg[22][11]/P0001 ,
		_w11935_,
		_w11986_,
		_w22138_
	);
	LUT3 #(
		.INIT('h80)
	) name11626 (
		\wishbone_bd_ram_mem1_reg[193][11]/P0001 ,
		_w11945_,
		_w11977_,
		_w22139_
	);
	LUT3 #(
		.INIT('h80)
	) name11627 (
		\wishbone_bd_ram_mem1_reg[11][11]/P0001 ,
		_w11932_,
		_w11936_,
		_w22140_
	);
	LUT3 #(
		.INIT('h80)
	) name11628 (
		\wishbone_bd_ram_mem1_reg[145][11]/P0001 ,
		_w11959_,
		_w11977_,
		_w22141_
	);
	LUT4 #(
		.INIT('h0001)
	) name11629 (
		_w22138_,
		_w22139_,
		_w22140_,
		_w22141_,
		_w22142_
	);
	LUT3 #(
		.INIT('h80)
	) name11630 (
		\wishbone_bd_ram_mem1_reg[105][11]/P0001 ,
		_w11965_,
		_w11968_,
		_w22143_
	);
	LUT3 #(
		.INIT('h80)
	) name11631 (
		\wishbone_bd_ram_mem1_reg[52][11]/P0001 ,
		_w11929_,
		_w11979_,
		_w22144_
	);
	LUT3 #(
		.INIT('h80)
	) name11632 (
		\wishbone_bd_ram_mem1_reg[155][11]/P0001 ,
		_w11936_,
		_w11959_,
		_w22145_
	);
	LUT3 #(
		.INIT('h80)
	) name11633 (
		\wishbone_bd_ram_mem1_reg[85][11]/P0001 ,
		_w11933_,
		_w11972_,
		_w22146_
	);
	LUT4 #(
		.INIT('h0001)
	) name11634 (
		_w22143_,
		_w22144_,
		_w22145_,
		_w22146_,
		_w22147_
	);
	LUT4 #(
		.INIT('h8000)
	) name11635 (
		_w22132_,
		_w22137_,
		_w22142_,
		_w22147_,
		_w22148_
	);
	LUT3 #(
		.INIT('h80)
	) name11636 (
		\wishbone_bd_ram_mem1_reg[24][11]/P0001 ,
		_w11935_,
		_w11990_,
		_w22149_
	);
	LUT3 #(
		.INIT('h80)
	) name11637 (
		\wishbone_bd_ram_mem1_reg[240][11]/P0001 ,
		_w11941_,
		_w11952_,
		_w22150_
	);
	LUT3 #(
		.INIT('h80)
	) name11638 (
		\wishbone_bd_ram_mem1_reg[230][11]/P0001 ,
		_w11982_,
		_w11986_,
		_w22151_
	);
	LUT3 #(
		.INIT('h80)
	) name11639 (
		\wishbone_bd_ram_mem1_reg[126][11]/P0001 ,
		_w11948_,
		_w12012_,
		_w22152_
	);
	LUT4 #(
		.INIT('h0001)
	) name11640 (
		_w22149_,
		_w22150_,
		_w22151_,
		_w22152_,
		_w22153_
	);
	LUT3 #(
		.INIT('h80)
	) name11641 (
		\wishbone_bd_ram_mem1_reg[39][11]/P0001 ,
		_w11957_,
		_w11975_,
		_w22154_
	);
	LUT3 #(
		.INIT('h80)
	) name11642 (
		\wishbone_bd_ram_mem1_reg[133][11]/P0001 ,
		_w11933_,
		_w11955_,
		_w22155_
	);
	LUT3 #(
		.INIT('h80)
	) name11643 (
		\wishbone_bd_ram_mem1_reg[159][11]/P0001 ,
		_w11959_,
		_w11973_,
		_w22156_
	);
	LUT3 #(
		.INIT('h80)
	) name11644 (
		\wishbone_bd_ram_mem1_reg[139][11]/P0001 ,
		_w11936_,
		_w11955_,
		_w22157_
	);
	LUT4 #(
		.INIT('h0001)
	) name11645 (
		_w22154_,
		_w22155_,
		_w22156_,
		_w22157_,
		_w22158_
	);
	LUT3 #(
		.INIT('h80)
	) name11646 (
		\wishbone_bd_ram_mem1_reg[60][11]/P0001 ,
		_w11954_,
		_w11979_,
		_w22159_
	);
	LUT3 #(
		.INIT('h80)
	) name11647 (
		\wishbone_bd_ram_mem1_reg[228][11]/P0001 ,
		_w11929_,
		_w11982_,
		_w22160_
	);
	LUT3 #(
		.INIT('h80)
	) name11648 (
		\wishbone_bd_ram_mem1_reg[92][11]/P0001 ,
		_w11954_,
		_w11972_,
		_w22161_
	);
	LUT3 #(
		.INIT('h80)
	) name11649 (
		\wishbone_bd_ram_mem1_reg[13][11]/P0001 ,
		_w11932_,
		_w11966_,
		_w22162_
	);
	LUT4 #(
		.INIT('h0001)
	) name11650 (
		_w22159_,
		_w22160_,
		_w22161_,
		_w22162_,
		_w22163_
	);
	LUT3 #(
		.INIT('h80)
	) name11651 (
		\wishbone_bd_ram_mem1_reg[5][11]/P0001 ,
		_w11932_,
		_w11933_,
		_w22164_
	);
	LUT3 #(
		.INIT('h80)
	) name11652 (
		\wishbone_bd_ram_mem1_reg[143][11]/P0001 ,
		_w11955_,
		_w11973_,
		_w22165_
	);
	LUT3 #(
		.INIT('h80)
	) name11653 (
		\wishbone_bd_ram_mem1_reg[226][11]/P0001 ,
		_w11963_,
		_w11982_,
		_w22166_
	);
	LUT3 #(
		.INIT('h80)
	) name11654 (
		\wishbone_bd_ram_mem1_reg[70][11]/P0001 ,
		_w11949_,
		_w11986_,
		_w22167_
	);
	LUT4 #(
		.INIT('h0001)
	) name11655 (
		_w22164_,
		_w22165_,
		_w22166_,
		_w22167_,
		_w22168_
	);
	LUT4 #(
		.INIT('h8000)
	) name11656 (
		_w22153_,
		_w22158_,
		_w22163_,
		_w22168_,
		_w22169_
	);
	LUT3 #(
		.INIT('h80)
	) name11657 (
		\wishbone_bd_ram_mem1_reg[235][11]/P0001 ,
		_w11936_,
		_w11982_,
		_w22170_
	);
	LUT3 #(
		.INIT('h80)
	) name11658 (
		\wishbone_bd_ram_mem1_reg[135][11]/P0001 ,
		_w11955_,
		_w11975_,
		_w22171_
	);
	LUT3 #(
		.INIT('h80)
	) name11659 (
		\wishbone_bd_ram_mem1_reg[149][11]/P0001 ,
		_w11933_,
		_w11959_,
		_w22172_
	);
	LUT3 #(
		.INIT('h80)
	) name11660 (
		\wishbone_bd_ram_mem1_reg[63][11]/P0001 ,
		_w11973_,
		_w11979_,
		_w22173_
	);
	LUT4 #(
		.INIT('h0001)
	) name11661 (
		_w22170_,
		_w22171_,
		_w22172_,
		_w22173_,
		_w22174_
	);
	LUT3 #(
		.INIT('h80)
	) name11662 (
		\wishbone_bd_ram_mem1_reg[156][11]/P0001 ,
		_w11954_,
		_w11959_,
		_w22175_
	);
	LUT3 #(
		.INIT('h80)
	) name11663 (
		\wishbone_bd_ram_mem1_reg[225][11]/P0001 ,
		_w11977_,
		_w11982_,
		_w22176_
	);
	LUT3 #(
		.INIT('h80)
	) name11664 (
		\wishbone_bd_ram_mem1_reg[238][11]/P0001 ,
		_w11948_,
		_w11982_,
		_w22177_
	);
	LUT3 #(
		.INIT('h80)
	) name11665 (
		\wishbone_bd_ram_mem1_reg[57][11]/P0001 ,
		_w11968_,
		_w11979_,
		_w22178_
	);
	LUT4 #(
		.INIT('h0001)
	) name11666 (
		_w22175_,
		_w22176_,
		_w22177_,
		_w22178_,
		_w22179_
	);
	LUT3 #(
		.INIT('h80)
	) name11667 (
		\wishbone_bd_ram_mem1_reg[86][11]/P0001 ,
		_w11972_,
		_w11986_,
		_w22180_
	);
	LUT3 #(
		.INIT('h80)
	) name11668 (
		\wishbone_bd_ram_mem1_reg[19][11]/P0001 ,
		_w11935_,
		_w11938_,
		_w22181_
	);
	LUT3 #(
		.INIT('h80)
	) name11669 (
		\wishbone_bd_ram_mem1_reg[166][11]/P0001 ,
		_w11930_,
		_w11986_,
		_w22182_
	);
	LUT3 #(
		.INIT('h80)
	) name11670 (
		\wishbone_bd_ram_mem1_reg[34][11]/P0001 ,
		_w11957_,
		_w11963_,
		_w22183_
	);
	LUT4 #(
		.INIT('h0001)
	) name11671 (
		_w22180_,
		_w22181_,
		_w22182_,
		_w22183_,
		_w22184_
	);
	LUT3 #(
		.INIT('h80)
	) name11672 (
		\wishbone_bd_ram_mem1_reg[251][11]/P0001 ,
		_w11936_,
		_w11952_,
		_w22185_
	);
	LUT3 #(
		.INIT('h80)
	) name11673 (
		\wishbone_bd_ram_mem1_reg[77][11]/P0001 ,
		_w11949_,
		_w11966_,
		_w22186_
	);
	LUT3 #(
		.INIT('h80)
	) name11674 (
		\wishbone_bd_ram_mem1_reg[165][11]/P0001 ,
		_w11930_,
		_w11933_,
		_w22187_
	);
	LUT3 #(
		.INIT('h80)
	) name11675 (
		\wishbone_bd_ram_mem1_reg[244][11]/P0001 ,
		_w11929_,
		_w11952_,
		_w22188_
	);
	LUT4 #(
		.INIT('h0001)
	) name11676 (
		_w22185_,
		_w22186_,
		_w22187_,
		_w22188_,
		_w22189_
	);
	LUT4 #(
		.INIT('h8000)
	) name11677 (
		_w22174_,
		_w22179_,
		_w22184_,
		_w22189_,
		_w22190_
	);
	LUT3 #(
		.INIT('h80)
	) name11678 (
		\wishbone_bd_ram_mem1_reg[102][11]/P0001 ,
		_w11965_,
		_w11986_,
		_w22191_
	);
	LUT3 #(
		.INIT('h80)
	) name11679 (
		\wishbone_bd_ram_mem1_reg[158][11]/P0001 ,
		_w11948_,
		_w11959_,
		_w22192_
	);
	LUT3 #(
		.INIT('h80)
	) name11680 (
		\wishbone_bd_ram_mem1_reg[140][11]/P0001 ,
		_w11954_,
		_w11955_,
		_w22193_
	);
	LUT3 #(
		.INIT('h80)
	) name11681 (
		\wishbone_bd_ram_mem1_reg[137][11]/P0001 ,
		_w11955_,
		_w11968_,
		_w22194_
	);
	LUT4 #(
		.INIT('h0001)
	) name11682 (
		_w22191_,
		_w22192_,
		_w22193_,
		_w22194_,
		_w22195_
	);
	LUT3 #(
		.INIT('h80)
	) name11683 (
		\wishbone_bd_ram_mem1_reg[116][11]/P0001 ,
		_w11929_,
		_w12012_,
		_w22196_
	);
	LUT3 #(
		.INIT('h80)
	) name11684 (
		\wishbone_bd_ram_mem1_reg[29][11]/P0001 ,
		_w11935_,
		_w11966_,
		_w22197_
	);
	LUT3 #(
		.INIT('h80)
	) name11685 (
		\wishbone_bd_ram_mem1_reg[59][11]/P0001 ,
		_w11936_,
		_w11979_,
		_w22198_
	);
	LUT3 #(
		.INIT('h80)
	) name11686 (
		\wishbone_bd_ram_mem1_reg[204][11]/P0001 ,
		_w11945_,
		_w11954_,
		_w22199_
	);
	LUT4 #(
		.INIT('h0001)
	) name11687 (
		_w22196_,
		_w22197_,
		_w22198_,
		_w22199_,
		_w22200_
	);
	LUT3 #(
		.INIT('h80)
	) name11688 (
		\wishbone_bd_ram_mem1_reg[15][11]/P0001 ,
		_w11932_,
		_w11973_,
		_w22201_
	);
	LUT3 #(
		.INIT('h80)
	) name11689 (
		\wishbone_bd_ram_mem1_reg[97][11]/P0001 ,
		_w11965_,
		_w11977_,
		_w22202_
	);
	LUT3 #(
		.INIT('h80)
	) name11690 (
		\wishbone_bd_ram_mem1_reg[94][11]/P0001 ,
		_w11948_,
		_w11972_,
		_w22203_
	);
	LUT3 #(
		.INIT('h80)
	) name11691 (
		\wishbone_bd_ram_mem1_reg[195][11]/P0001 ,
		_w11938_,
		_w11945_,
		_w22204_
	);
	LUT4 #(
		.INIT('h0001)
	) name11692 (
		_w22201_,
		_w22202_,
		_w22203_,
		_w22204_,
		_w22205_
	);
	LUT3 #(
		.INIT('h80)
	) name11693 (
		\wishbone_bd_ram_mem1_reg[23][11]/P0001 ,
		_w11935_,
		_w11975_,
		_w22206_
	);
	LUT3 #(
		.INIT('h80)
	) name11694 (
		\wishbone_bd_ram_mem1_reg[249][11]/P0001 ,
		_w11952_,
		_w11968_,
		_w22207_
	);
	LUT3 #(
		.INIT('h80)
	) name11695 (
		\wishbone_bd_ram_mem1_reg[1][11]/P0001 ,
		_w11932_,
		_w11977_,
		_w22208_
	);
	LUT3 #(
		.INIT('h80)
	) name11696 (
		\wishbone_bd_ram_mem1_reg[209][11]/P0001 ,
		_w11977_,
		_w11984_,
		_w22209_
	);
	LUT4 #(
		.INIT('h0001)
	) name11697 (
		_w22206_,
		_w22207_,
		_w22208_,
		_w22209_,
		_w22210_
	);
	LUT4 #(
		.INIT('h8000)
	) name11698 (
		_w22195_,
		_w22200_,
		_w22205_,
		_w22210_,
		_w22211_
	);
	LUT4 #(
		.INIT('h8000)
	) name11699 (
		_w22148_,
		_w22169_,
		_w22190_,
		_w22211_,
		_w22212_
	);
	LUT4 #(
		.INIT('h8000)
	) name11700 (
		_w21957_,
		_w22042_,
		_w22127_,
		_w22212_,
		_w22213_
	);
	LUT4 #(
		.INIT('h1555)
	) name11701 (
		wb_rst_i_pad,
		_w21862_,
		_w21866_,
		_w21871_,
		_w22214_
	);
	LUT3 #(
		.INIT('hba)
	) name11702 (
		_w21872_,
		_w22213_,
		_w22214_,
		_w22215_
	);
	LUT4 #(
		.INIT('h0001)
	) name11703 (
		\wishbone_TxLength_reg[10]/NET0131 ,
		\wishbone_TxLength_reg[7]/NET0131 ,
		\wishbone_TxLength_reg[8]/NET0131 ,
		\wishbone_TxLength_reg[9]/NET0131 ,
		_w22216_
	);
	LUT3 #(
		.INIT('h80)
	) name11704 (
		_w12309_,
		_w12310_,
		_w22216_,
		_w22217_
	);
	LUT2 #(
		.INIT('h4)
	) name11705 (
		_w14878_,
		_w22217_,
		_w22218_
	);
	LUT3 #(
		.INIT('h48)
	) name11706 (
		\wishbone_TxLength_reg[11]/NET0131 ,
		_w15777_,
		_w22218_,
		_w22219_
	);
	LUT3 #(
		.INIT('hf2)
	) name11707 (
		_w12303_,
		_w17356_,
		_w22219_,
		_w22220_
	);
	LUT3 #(
		.INIT('h80)
	) name11708 (
		\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 ,
		_w18753_,
		_w18754_,
		_w22221_
	);
	LUT4 #(
		.INIT('h0008)
	) name11709 (
		\ethreg1_RXHASH1_0_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22222_
	);
	LUT3 #(
		.INIT('h80)
	) name11710 (
		_w18757_,
		_w18762_,
		_w22222_,
		_w22223_
	);
	LUT3 #(
		.INIT('h80)
	) name11711 (
		\ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131 ,
		_w18786_,
		_w18801_,
		_w22224_
	);
	LUT4 #(
		.INIT('h0008)
	) name11712 (
		\ethreg1_RXHASH0_0_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22225_
	);
	LUT3 #(
		.INIT('h80)
	) name11713 (
		_w18757_,
		_w18758_,
		_w22225_,
		_w22226_
	);
	LUT3 #(
		.INIT('h80)
	) name11714 (
		\ethreg1_IPGT_0_DataOut_reg[2]/NET0131 ,
		_w19646_,
		_w19655_,
		_w22227_
	);
	LUT4 #(
		.INIT('h0001)
	) name11715 (
		_w22223_,
		_w22224_,
		_w22226_,
		_w22227_,
		_w22228_
	);
	LUT3 #(
		.INIT('h80)
	) name11716 (
		\ethreg1_INT_MASK_0_DataOut_reg[2]/NET0131 ,
		_w18801_,
		_w19655_,
		_w22229_
	);
	LUT4 #(
		.INIT('h0002)
	) name11717 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22230_
	);
	LUT3 #(
		.INIT('h80)
	) name11718 (
		_w18757_,
		_w18762_,
		_w22230_,
		_w22231_
	);
	LUT3 #(
		.INIT('h80)
	) name11719 (
		\ethreg1_MIIRX_DATA_DataOut_reg[2]/NET0131 ,
		_w18785_,
		_w18786_,
		_w22232_
	);
	LUT3 #(
		.INIT('h80)
	) name11720 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[2]/NET0131 ,
		_w18798_,
		_w18801_,
		_w22233_
	);
	LUT4 #(
		.INIT('h0001)
	) name11721 (
		_w22229_,
		_w22231_,
		_w22232_,
		_w22233_,
		_w22234_
	);
	LUT3 #(
		.INIT('h40)
	) name11722 (
		_w22221_,
		_w22228_,
		_w22234_,
		_w22235_
	);
	LUT4 #(
		.INIT('h0002)
	) name11723 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22236_
	);
	LUT4 #(
		.INIT('h0020)
	) name11724 (
		\ethreg1_TXCTRL_0_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22237_
	);
	LUT4 #(
		.INIT('h777f)
	) name11725 (
		_w18757_,
		_w18758_,
		_w22236_,
		_w22237_,
		_w22238_
	);
	LUT3 #(
		.INIT('h80)
	) name11726 (
		\ethreg1_IPGR1_0_DataOut_reg[2]/NET0131 ,
		_w18785_,
		_w18800_,
		_w22239_
	);
	LUT3 #(
		.INIT('h80)
	) name11727 (
		\ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131 ,
		_w18798_,
		_w19646_,
		_w22240_
	);
	LUT4 #(
		.INIT('h0008)
	) name11728 (
		_w18752_,
		_w22238_,
		_w22239_,
		_w22240_,
		_w22241_
	);
	LUT3 #(
		.INIT('h80)
	) name11729 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[2]/NET0131 ,
		_w18785_,
		_w18798_,
		_w22242_
	);
	LUT3 #(
		.INIT('h80)
	) name11730 (
		\miim1_Nvalid_reg/NET0131 ,
		_w18786_,
		_w18805_,
		_w22243_
	);
	LUT3 #(
		.INIT('h80)
	) name11731 (
		\ethreg1_MIICOMMAND2_DataOut_reg[0]/NET0131 ,
		_w18786_,
		_w19646_,
		_w22244_
	);
	LUT3 #(
		.INIT('h80)
	) name11732 (
		\ethreg1_irq_rxb_reg/NET0131 ,
		_w18800_,
		_w19646_,
		_w22245_
	);
	LUT4 #(
		.INIT('h0001)
	) name11733 (
		_w22242_,
		_w22243_,
		_w22244_,
		_w22245_,
		_w22246_
	);
	LUT3 #(
		.INIT('h80)
	) name11734 (
		\ethreg1_MODER_0_DataOut_reg[2]/NET0131 ,
		_w18800_,
		_w18801_,
		_w22247_
	);
	LUT3 #(
		.INIT('h80)
	) name11735 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[2]/NET0131 ,
		_w18798_,
		_w18805_,
		_w22248_
	);
	LUT3 #(
		.INIT('h80)
	) name11736 (
		\ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131 ,
		_w18805_,
		_w19655_,
		_w22249_
	);
	LUT3 #(
		.INIT('h80)
	) name11737 (
		\ethreg1_IPGR2_0_DataOut_reg[2]/NET0131 ,
		_w18800_,
		_w18805_,
		_w22250_
	);
	LUT4 #(
		.INIT('h0001)
	) name11738 (
		_w22247_,
		_w22248_,
		_w22249_,
		_w22250_,
		_w22251_
	);
	LUT3 #(
		.INIT('h80)
	) name11739 (
		_w22241_,
		_w22246_,
		_w22251_,
		_w22252_
	);
	LUT3 #(
		.INIT('h2a)
	) name11740 (
		_w18752_,
		_w22235_,
		_w22252_,
		_w22253_
	);
	LUT3 #(
		.INIT('h80)
	) name11741 (
		\wishbone_bd_ram_mem0_reg[43][2]/P0001 ,
		_w11936_,
		_w11957_,
		_w22254_
	);
	LUT3 #(
		.INIT('h80)
	) name11742 (
		\wishbone_bd_ram_mem0_reg[13][2]/P0001 ,
		_w11932_,
		_w11966_,
		_w22255_
	);
	LUT3 #(
		.INIT('h80)
	) name11743 (
		\wishbone_bd_ram_mem0_reg[50][2]/P0001 ,
		_w11963_,
		_w11979_,
		_w22256_
	);
	LUT3 #(
		.INIT('h80)
	) name11744 (
		\wishbone_bd_ram_mem0_reg[87][2]/P0001 ,
		_w11972_,
		_w11975_,
		_w22257_
	);
	LUT4 #(
		.INIT('h0001)
	) name11745 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22257_,
		_w22258_
	);
	LUT3 #(
		.INIT('h80)
	) name11746 (
		\wishbone_bd_ram_mem0_reg[91][2]/P0001 ,
		_w11936_,
		_w11972_,
		_w22259_
	);
	LUT3 #(
		.INIT('h80)
	) name11747 (
		\wishbone_bd_ram_mem0_reg[193][2]/P0001 ,
		_w11945_,
		_w11977_,
		_w22260_
	);
	LUT3 #(
		.INIT('h80)
	) name11748 (
		\wishbone_bd_ram_mem0_reg[160][2]/P0001 ,
		_w11930_,
		_w11941_,
		_w22261_
	);
	LUT3 #(
		.INIT('h80)
	) name11749 (
		\wishbone_bd_ram_mem0_reg[236][2]/P0001 ,
		_w11954_,
		_w11982_,
		_w22262_
	);
	LUT4 #(
		.INIT('h0001)
	) name11750 (
		_w22259_,
		_w22260_,
		_w22261_,
		_w22262_,
		_w22263_
	);
	LUT3 #(
		.INIT('h80)
	) name11751 (
		\wishbone_bd_ram_mem0_reg[240][2]/P0001 ,
		_w11941_,
		_w11952_,
		_w22264_
	);
	LUT3 #(
		.INIT('h80)
	) name11752 (
		\wishbone_bd_ram_mem0_reg[179][2]/P0001 ,
		_w11938_,
		_w11942_,
		_w22265_
	);
	LUT3 #(
		.INIT('h80)
	) name11753 (
		\wishbone_bd_ram_mem0_reg[34][2]/P0001 ,
		_w11957_,
		_w11963_,
		_w22266_
	);
	LUT3 #(
		.INIT('h80)
	) name11754 (
		\wishbone_bd_ram_mem0_reg[186][2]/P0001 ,
		_w11942_,
		_w11944_,
		_w22267_
	);
	LUT4 #(
		.INIT('h0001)
	) name11755 (
		_w22264_,
		_w22265_,
		_w22266_,
		_w22267_,
		_w22268_
	);
	LUT3 #(
		.INIT('h80)
	) name11756 (
		\wishbone_bd_ram_mem0_reg[28][2]/P0001 ,
		_w11935_,
		_w11954_,
		_w22269_
	);
	LUT3 #(
		.INIT('h80)
	) name11757 (
		\wishbone_bd_ram_mem0_reg[248][2]/P0001 ,
		_w11952_,
		_w11990_,
		_w22270_
	);
	LUT3 #(
		.INIT('h80)
	) name11758 (
		\wishbone_bd_ram_mem0_reg[11][2]/P0001 ,
		_w11932_,
		_w11936_,
		_w22271_
	);
	LUT3 #(
		.INIT('h80)
	) name11759 (
		\wishbone_bd_ram_mem0_reg[231][2]/P0001 ,
		_w11975_,
		_w11982_,
		_w22272_
	);
	LUT4 #(
		.INIT('h0001)
	) name11760 (
		_w22269_,
		_w22270_,
		_w22271_,
		_w22272_,
		_w22273_
	);
	LUT4 #(
		.INIT('h8000)
	) name11761 (
		_w22258_,
		_w22263_,
		_w22268_,
		_w22273_,
		_w22274_
	);
	LUT3 #(
		.INIT('h80)
	) name11762 (
		\wishbone_bd_ram_mem0_reg[104][2]/P0001 ,
		_w11965_,
		_w11990_,
		_w22275_
	);
	LUT3 #(
		.INIT('h80)
	) name11763 (
		\wishbone_bd_ram_mem0_reg[153][2]/P0001 ,
		_w11959_,
		_w11968_,
		_w22276_
	);
	LUT3 #(
		.INIT('h80)
	) name11764 (
		\wishbone_bd_ram_mem0_reg[44][2]/P0001 ,
		_w11954_,
		_w11957_,
		_w22277_
	);
	LUT3 #(
		.INIT('h80)
	) name11765 (
		\wishbone_bd_ram_mem0_reg[59][2]/P0001 ,
		_w11936_,
		_w11979_,
		_w22278_
	);
	LUT4 #(
		.INIT('h0001)
	) name11766 (
		_w22275_,
		_w22276_,
		_w22277_,
		_w22278_,
		_w22279_
	);
	LUT3 #(
		.INIT('h80)
	) name11767 (
		\wishbone_bd_ram_mem0_reg[233][2]/P0001 ,
		_w11968_,
		_w11982_,
		_w22280_
	);
	LUT3 #(
		.INIT('h80)
	) name11768 (
		\wishbone_bd_ram_mem0_reg[183][2]/P0001 ,
		_w11942_,
		_w11975_,
		_w22281_
	);
	LUT3 #(
		.INIT('h80)
	) name11769 (
		\wishbone_bd_ram_mem0_reg[70][2]/P0001 ,
		_w11949_,
		_w11986_,
		_w22282_
	);
	LUT3 #(
		.INIT('h80)
	) name11770 (
		\wishbone_bd_ram_mem0_reg[2][2]/P0001 ,
		_w11932_,
		_w11963_,
		_w22283_
	);
	LUT4 #(
		.INIT('h0001)
	) name11771 (
		_w22280_,
		_w22281_,
		_w22282_,
		_w22283_,
		_w22284_
	);
	LUT3 #(
		.INIT('h80)
	) name11772 (
		\wishbone_bd_ram_mem0_reg[166][2]/P0001 ,
		_w11930_,
		_w11986_,
		_w22285_
	);
	LUT3 #(
		.INIT('h80)
	) name11773 (
		\wishbone_bd_ram_mem0_reg[207][2]/P0001 ,
		_w11945_,
		_w11973_,
		_w22286_
	);
	LUT3 #(
		.INIT('h80)
	) name11774 (
		\wishbone_bd_ram_mem0_reg[178][2]/P0001 ,
		_w11942_,
		_w11963_,
		_w22287_
	);
	LUT3 #(
		.INIT('h80)
	) name11775 (
		\wishbone_bd_ram_mem0_reg[118][2]/P0001 ,
		_w11986_,
		_w12012_,
		_w22288_
	);
	LUT4 #(
		.INIT('h0001)
	) name11776 (
		_w22285_,
		_w22286_,
		_w22287_,
		_w22288_,
		_w22289_
	);
	LUT3 #(
		.INIT('h80)
	) name11777 (
		\wishbone_bd_ram_mem0_reg[1][2]/P0001 ,
		_w11932_,
		_w11977_,
		_w22290_
	);
	LUT3 #(
		.INIT('h80)
	) name11778 (
		\wishbone_bd_ram_mem0_reg[170][2]/P0001 ,
		_w11930_,
		_w11944_,
		_w22291_
	);
	LUT3 #(
		.INIT('h80)
	) name11779 (
		\wishbone_bd_ram_mem0_reg[103][2]/P0001 ,
		_w11965_,
		_w11975_,
		_w22292_
	);
	LUT3 #(
		.INIT('h80)
	) name11780 (
		\wishbone_bd_ram_mem0_reg[194][2]/P0001 ,
		_w11945_,
		_w11963_,
		_w22293_
	);
	LUT4 #(
		.INIT('h0001)
	) name11781 (
		_w22290_,
		_w22291_,
		_w22292_,
		_w22293_,
		_w22294_
	);
	LUT4 #(
		.INIT('h8000)
	) name11782 (
		_w22279_,
		_w22284_,
		_w22289_,
		_w22294_,
		_w22295_
	);
	LUT3 #(
		.INIT('h80)
	) name11783 (
		\wishbone_bd_ram_mem0_reg[88][2]/P0001 ,
		_w11972_,
		_w11990_,
		_w22296_
	);
	LUT3 #(
		.INIT('h80)
	) name11784 (
		\wishbone_bd_ram_mem0_reg[82][2]/P0001 ,
		_w11963_,
		_w11972_,
		_w22297_
	);
	LUT3 #(
		.INIT('h80)
	) name11785 (
		\wishbone_bd_ram_mem0_reg[169][2]/P0001 ,
		_w11930_,
		_w11968_,
		_w22298_
	);
	LUT3 #(
		.INIT('h80)
	) name11786 (
		\wishbone_bd_ram_mem0_reg[84][2]/P0001 ,
		_w11929_,
		_w11972_,
		_w22299_
	);
	LUT4 #(
		.INIT('h0001)
	) name11787 (
		_w22296_,
		_w22297_,
		_w22298_,
		_w22299_,
		_w22300_
	);
	LUT3 #(
		.INIT('h80)
	) name11788 (
		\wishbone_bd_ram_mem0_reg[199][2]/P0001 ,
		_w11945_,
		_w11975_,
		_w22301_
	);
	LUT3 #(
		.INIT('h80)
	) name11789 (
		\wishbone_bd_ram_mem0_reg[164][2]/P0001 ,
		_w11929_,
		_w11930_,
		_w22302_
	);
	LUT3 #(
		.INIT('h80)
	) name11790 (
		\wishbone_bd_ram_mem0_reg[249][2]/P0001 ,
		_w11952_,
		_w11968_,
		_w22303_
	);
	LUT3 #(
		.INIT('h80)
	) name11791 (
		\wishbone_bd_ram_mem0_reg[98][2]/P0001 ,
		_w11963_,
		_w11965_,
		_w22304_
	);
	LUT4 #(
		.INIT('h0001)
	) name11792 (
		_w22301_,
		_w22302_,
		_w22303_,
		_w22304_,
		_w22305_
	);
	LUT3 #(
		.INIT('h80)
	) name11793 (
		\wishbone_bd_ram_mem0_reg[143][2]/P0001 ,
		_w11955_,
		_w11973_,
		_w22306_
	);
	LUT3 #(
		.INIT('h80)
	) name11794 (
		\wishbone_bd_ram_mem0_reg[7][2]/P0001 ,
		_w11932_,
		_w11975_,
		_w22307_
	);
	LUT3 #(
		.INIT('h80)
	) name11795 (
		\wishbone_bd_ram_mem0_reg[142][2]/P0001 ,
		_w11948_,
		_w11955_,
		_w22308_
	);
	LUT3 #(
		.INIT('h80)
	) name11796 (
		\wishbone_bd_ram_mem0_reg[237][2]/P0001 ,
		_w11966_,
		_w11982_,
		_w22309_
	);
	LUT4 #(
		.INIT('h0001)
	) name11797 (
		_w22306_,
		_w22307_,
		_w22308_,
		_w22309_,
		_w22310_
	);
	LUT3 #(
		.INIT('h80)
	) name11798 (
		\wishbone_bd_ram_mem0_reg[112][2]/P0001 ,
		_w11941_,
		_w12012_,
		_w22311_
	);
	LUT3 #(
		.INIT('h80)
	) name11799 (
		\wishbone_bd_ram_mem0_reg[245][2]/P0001 ,
		_w11933_,
		_w11952_,
		_w22312_
	);
	LUT3 #(
		.INIT('h80)
	) name11800 (
		\wishbone_bd_ram_mem0_reg[57][2]/P0001 ,
		_w11968_,
		_w11979_,
		_w22313_
	);
	LUT3 #(
		.INIT('h80)
	) name11801 (
		\wishbone_bd_ram_mem0_reg[206][2]/P0001 ,
		_w11945_,
		_w11948_,
		_w22314_
	);
	LUT4 #(
		.INIT('h0001)
	) name11802 (
		_w22311_,
		_w22312_,
		_w22313_,
		_w22314_,
		_w22315_
	);
	LUT4 #(
		.INIT('h8000)
	) name11803 (
		_w22300_,
		_w22305_,
		_w22310_,
		_w22315_,
		_w22316_
	);
	LUT3 #(
		.INIT('h80)
	) name11804 (
		\wishbone_bd_ram_mem0_reg[214][2]/P0001 ,
		_w11984_,
		_w11986_,
		_w22317_
	);
	LUT3 #(
		.INIT('h80)
	) name11805 (
		\wishbone_bd_ram_mem0_reg[174][2]/P0001 ,
		_w11930_,
		_w11948_,
		_w22318_
	);
	LUT3 #(
		.INIT('h80)
	) name11806 (
		\wishbone_bd_ram_mem0_reg[96][2]/P0001 ,
		_w11941_,
		_w11965_,
		_w22319_
	);
	LUT3 #(
		.INIT('h80)
	) name11807 (
		\wishbone_bd_ram_mem0_reg[189][2]/P0001 ,
		_w11942_,
		_w11966_,
		_w22320_
	);
	LUT4 #(
		.INIT('h0001)
	) name11808 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22321_
	);
	LUT3 #(
		.INIT('h80)
	) name11809 (
		\wishbone_bd_ram_mem0_reg[190][2]/P0001 ,
		_w11942_,
		_w11948_,
		_w22322_
	);
	LUT3 #(
		.INIT('h80)
	) name11810 (
		\wishbone_bd_ram_mem0_reg[140][2]/P0001 ,
		_w11954_,
		_w11955_,
		_w22323_
	);
	LUT3 #(
		.INIT('h80)
	) name11811 (
		\wishbone_bd_ram_mem0_reg[149][2]/P0001 ,
		_w11933_,
		_w11959_,
		_w22324_
	);
	LUT3 #(
		.INIT('h80)
	) name11812 (
		\wishbone_bd_ram_mem0_reg[24][2]/P0001 ,
		_w11935_,
		_w11990_,
		_w22325_
	);
	LUT4 #(
		.INIT('h0001)
	) name11813 (
		_w22322_,
		_w22323_,
		_w22324_,
		_w22325_,
		_w22326_
	);
	LUT3 #(
		.INIT('h80)
	) name11814 (
		\wishbone_bd_ram_mem0_reg[210][2]/P0001 ,
		_w11963_,
		_w11984_,
		_w22327_
	);
	LUT3 #(
		.INIT('h80)
	) name11815 (
		\wishbone_bd_ram_mem0_reg[47][2]/P0001 ,
		_w11957_,
		_w11973_,
		_w22328_
	);
	LUT3 #(
		.INIT('h80)
	) name11816 (
		\wishbone_bd_ram_mem0_reg[195][2]/P0001 ,
		_w11938_,
		_w11945_,
		_w22329_
	);
	LUT3 #(
		.INIT('h80)
	) name11817 (
		\wishbone_bd_ram_mem0_reg[39][2]/P0001 ,
		_w11957_,
		_w11975_,
		_w22330_
	);
	LUT4 #(
		.INIT('h0001)
	) name11818 (
		_w22327_,
		_w22328_,
		_w22329_,
		_w22330_,
		_w22331_
	);
	LUT3 #(
		.INIT('h80)
	) name11819 (
		\wishbone_bd_ram_mem0_reg[163][2]/P0001 ,
		_w11930_,
		_w11938_,
		_w22332_
	);
	LUT3 #(
		.INIT('h80)
	) name11820 (
		\wishbone_bd_ram_mem0_reg[73][2]/P0001 ,
		_w11949_,
		_w11968_,
		_w22333_
	);
	LUT3 #(
		.INIT('h80)
	) name11821 (
		\wishbone_bd_ram_mem0_reg[64][2]/P0001 ,
		_w11941_,
		_w11949_,
		_w22334_
	);
	LUT3 #(
		.INIT('h80)
	) name11822 (
		\wishbone_bd_ram_mem0_reg[145][2]/P0001 ,
		_w11959_,
		_w11977_,
		_w22335_
	);
	LUT4 #(
		.INIT('h0001)
	) name11823 (
		_w22332_,
		_w22333_,
		_w22334_,
		_w22335_,
		_w22336_
	);
	LUT4 #(
		.INIT('h8000)
	) name11824 (
		_w22321_,
		_w22326_,
		_w22331_,
		_w22336_,
		_w22337_
	);
	LUT4 #(
		.INIT('h8000)
	) name11825 (
		_w22274_,
		_w22295_,
		_w22316_,
		_w22337_,
		_w22338_
	);
	LUT3 #(
		.INIT('h80)
	) name11826 (
		\wishbone_bd_ram_mem0_reg[157][2]/P0001 ,
		_w11959_,
		_w11966_,
		_w22339_
	);
	LUT3 #(
		.INIT('h80)
	) name11827 (
		\wishbone_bd_ram_mem0_reg[124][2]/P0001 ,
		_w11954_,
		_w12012_,
		_w22340_
	);
	LUT3 #(
		.INIT('h80)
	) name11828 (
		\wishbone_bd_ram_mem0_reg[113][2]/P0001 ,
		_w11977_,
		_w12012_,
		_w22341_
	);
	LUT3 #(
		.INIT('h80)
	) name11829 (
		\wishbone_bd_ram_mem0_reg[146][2]/P0001 ,
		_w11959_,
		_w11963_,
		_w22342_
	);
	LUT4 #(
		.INIT('h0001)
	) name11830 (
		_w22339_,
		_w22340_,
		_w22341_,
		_w22342_,
		_w22343_
	);
	LUT3 #(
		.INIT('h80)
	) name11831 (
		\wishbone_bd_ram_mem0_reg[212][2]/P0001 ,
		_w11929_,
		_w11984_,
		_w22344_
	);
	LUT3 #(
		.INIT('h80)
	) name11832 (
		\wishbone_bd_ram_mem0_reg[25][2]/P0001 ,
		_w11935_,
		_w11968_,
		_w22345_
	);
	LUT3 #(
		.INIT('h80)
	) name11833 (
		\wishbone_bd_ram_mem0_reg[85][2]/P0001 ,
		_w11933_,
		_w11972_,
		_w22346_
	);
	LUT3 #(
		.INIT('h80)
	) name11834 (
		\wishbone_bd_ram_mem0_reg[72][2]/P0001 ,
		_w11949_,
		_w11990_,
		_w22347_
	);
	LUT4 #(
		.INIT('h0001)
	) name11835 (
		_w22344_,
		_w22345_,
		_w22346_,
		_w22347_,
		_w22348_
	);
	LUT3 #(
		.INIT('h80)
	) name11836 (
		\wishbone_bd_ram_mem0_reg[196][2]/P0001 ,
		_w11929_,
		_w11945_,
		_w22349_
	);
	LUT3 #(
		.INIT('h80)
	) name11837 (
		\wishbone_bd_ram_mem0_reg[100][2]/P0001 ,
		_w11929_,
		_w11965_,
		_w22350_
	);
	LUT3 #(
		.INIT('h80)
	) name11838 (
		\wishbone_bd_ram_mem0_reg[198][2]/P0001 ,
		_w11945_,
		_w11986_,
		_w22351_
	);
	LUT3 #(
		.INIT('h80)
	) name11839 (
		\wishbone_bd_ram_mem0_reg[224][2]/P0001 ,
		_w11941_,
		_w11982_,
		_w22352_
	);
	LUT4 #(
		.INIT('h0001)
	) name11840 (
		_w22349_,
		_w22350_,
		_w22351_,
		_w22352_,
		_w22353_
	);
	LUT3 #(
		.INIT('h80)
	) name11841 (
		\wishbone_bd_ram_mem0_reg[188][2]/P0001 ,
		_w11942_,
		_w11954_,
		_w22354_
	);
	LUT3 #(
		.INIT('h80)
	) name11842 (
		\wishbone_bd_ram_mem0_reg[26][2]/P0001 ,
		_w11935_,
		_w11944_,
		_w22355_
	);
	LUT3 #(
		.INIT('h80)
	) name11843 (
		\wishbone_bd_ram_mem0_reg[108][2]/P0001 ,
		_w11954_,
		_w11965_,
		_w22356_
	);
	LUT3 #(
		.INIT('h80)
	) name11844 (
		\wishbone_bd_ram_mem0_reg[228][2]/P0001 ,
		_w11929_,
		_w11982_,
		_w22357_
	);
	LUT4 #(
		.INIT('h0001)
	) name11845 (
		_w22354_,
		_w22355_,
		_w22356_,
		_w22357_,
		_w22358_
	);
	LUT4 #(
		.INIT('h8000)
	) name11846 (
		_w22343_,
		_w22348_,
		_w22353_,
		_w22358_,
		_w22359_
	);
	LUT3 #(
		.INIT('h80)
	) name11847 (
		\wishbone_bd_ram_mem0_reg[80][2]/P0001 ,
		_w11941_,
		_w11972_,
		_w22360_
	);
	LUT3 #(
		.INIT('h80)
	) name11848 (
		\wishbone_bd_ram_mem0_reg[235][2]/P0001 ,
		_w11936_,
		_w11982_,
		_w22361_
	);
	LUT3 #(
		.INIT('h80)
	) name11849 (
		\wishbone_bd_ram_mem0_reg[135][2]/P0001 ,
		_w11955_,
		_w11975_,
		_w22362_
	);
	LUT3 #(
		.INIT('h80)
	) name11850 (
		\wishbone_bd_ram_mem0_reg[31][2]/P0001 ,
		_w11935_,
		_w11973_,
		_w22363_
	);
	LUT4 #(
		.INIT('h0001)
	) name11851 (
		_w22360_,
		_w22361_,
		_w22362_,
		_w22363_,
		_w22364_
	);
	LUT3 #(
		.INIT('h80)
	) name11852 (
		\wishbone_bd_ram_mem0_reg[8][2]/P0001 ,
		_w11932_,
		_w11990_,
		_w22365_
	);
	LUT3 #(
		.INIT('h80)
	) name11853 (
		\wishbone_bd_ram_mem0_reg[60][2]/P0001 ,
		_w11954_,
		_w11979_,
		_w22366_
	);
	LUT3 #(
		.INIT('h80)
	) name11854 (
		\wishbone_bd_ram_mem0_reg[42][2]/P0001 ,
		_w11944_,
		_w11957_,
		_w22367_
	);
	LUT3 #(
		.INIT('h80)
	) name11855 (
		\wishbone_bd_ram_mem0_reg[95][2]/P0001 ,
		_w11972_,
		_w11973_,
		_w22368_
	);
	LUT4 #(
		.INIT('h0001)
	) name11856 (
		_w22365_,
		_w22366_,
		_w22367_,
		_w22368_,
		_w22369_
	);
	LUT3 #(
		.INIT('h80)
	) name11857 (
		\wishbone_bd_ram_mem0_reg[16][2]/P0001 ,
		_w11935_,
		_w11941_,
		_w22370_
	);
	LUT3 #(
		.INIT('h80)
	) name11858 (
		\wishbone_bd_ram_mem0_reg[219][2]/P0001 ,
		_w11936_,
		_w11984_,
		_w22371_
	);
	LUT3 #(
		.INIT('h80)
	) name11859 (
		\wishbone_bd_ram_mem0_reg[38][2]/P0001 ,
		_w11957_,
		_w11986_,
		_w22372_
	);
	LUT3 #(
		.INIT('h80)
	) name11860 (
		\wishbone_bd_ram_mem0_reg[23][2]/P0001 ,
		_w11935_,
		_w11975_,
		_w22373_
	);
	LUT4 #(
		.INIT('h0001)
	) name11861 (
		_w22370_,
		_w22371_,
		_w22372_,
		_w22373_,
		_w22374_
	);
	LUT3 #(
		.INIT('h80)
	) name11862 (
		\wishbone_bd_ram_mem0_reg[121][2]/P0001 ,
		_w11968_,
		_w12012_,
		_w22375_
	);
	LUT3 #(
		.INIT('h80)
	) name11863 (
		\wishbone_bd_ram_mem0_reg[246][2]/P0001 ,
		_w11952_,
		_w11986_,
		_w22376_
	);
	LUT3 #(
		.INIT('h80)
	) name11864 (
		\wishbone_bd_ram_mem0_reg[200][2]/P0001 ,
		_w11945_,
		_w11990_,
		_w22377_
	);
	LUT3 #(
		.INIT('h80)
	) name11865 (
		\wishbone_bd_ram_mem0_reg[136][2]/P0001 ,
		_w11955_,
		_w11990_,
		_w22378_
	);
	LUT4 #(
		.INIT('h0001)
	) name11866 (
		_w22375_,
		_w22376_,
		_w22377_,
		_w22378_,
		_w22379_
	);
	LUT4 #(
		.INIT('h8000)
	) name11867 (
		_w22364_,
		_w22369_,
		_w22374_,
		_w22379_,
		_w22380_
	);
	LUT3 #(
		.INIT('h80)
	) name11868 (
		\wishbone_bd_ram_mem0_reg[76][2]/P0001 ,
		_w11949_,
		_w11954_,
		_w22381_
	);
	LUT3 #(
		.INIT('h80)
	) name11869 (
		\wishbone_bd_ram_mem0_reg[132][2]/P0001 ,
		_w11929_,
		_w11955_,
		_w22382_
	);
	LUT3 #(
		.INIT('h80)
	) name11870 (
		\wishbone_bd_ram_mem0_reg[102][2]/P0001 ,
		_w11965_,
		_w11986_,
		_w22383_
	);
	LUT3 #(
		.INIT('h80)
	) name11871 (
		\wishbone_bd_ram_mem0_reg[114][2]/P0001 ,
		_w11963_,
		_w12012_,
		_w22384_
	);
	LUT4 #(
		.INIT('h0001)
	) name11872 (
		_w22381_,
		_w22382_,
		_w22383_,
		_w22384_,
		_w22385_
	);
	LUT3 #(
		.INIT('h80)
	) name11873 (
		\wishbone_bd_ram_mem0_reg[242][2]/P0001 ,
		_w11952_,
		_w11963_,
		_w22386_
	);
	LUT3 #(
		.INIT('h80)
	) name11874 (
		\wishbone_bd_ram_mem0_reg[238][2]/P0001 ,
		_w11948_,
		_w11982_,
		_w22387_
	);
	LUT3 #(
		.INIT('h80)
	) name11875 (
		\wishbone_bd_ram_mem0_reg[223][2]/P0001 ,
		_w11973_,
		_w11984_,
		_w22388_
	);
	LUT3 #(
		.INIT('h80)
	) name11876 (
		\wishbone_bd_ram_mem0_reg[86][2]/P0001 ,
		_w11972_,
		_w11986_,
		_w22389_
	);
	LUT4 #(
		.INIT('h0001)
	) name11877 (
		_w22386_,
		_w22387_,
		_w22388_,
		_w22389_,
		_w22390_
	);
	LUT3 #(
		.INIT('h80)
	) name11878 (
		\wishbone_bd_ram_mem0_reg[221][2]/P0001 ,
		_w11966_,
		_w11984_,
		_w22391_
	);
	LUT3 #(
		.INIT('h80)
	) name11879 (
		\wishbone_bd_ram_mem0_reg[131][2]/P0001 ,
		_w11938_,
		_w11955_,
		_w22392_
	);
	LUT3 #(
		.INIT('h80)
	) name11880 (
		\wishbone_bd_ram_mem0_reg[222][2]/P0001 ,
		_w11948_,
		_w11984_,
		_w22393_
	);
	LUT3 #(
		.INIT('h80)
	) name11881 (
		\wishbone_bd_ram_mem0_reg[255][2]/P0001 ,
		_w11952_,
		_w11973_,
		_w22394_
	);
	LUT4 #(
		.INIT('h0001)
	) name11882 (
		_w22391_,
		_w22392_,
		_w22393_,
		_w22394_,
		_w22395_
	);
	LUT3 #(
		.INIT('h80)
	) name11883 (
		\wishbone_bd_ram_mem0_reg[192][2]/P0001 ,
		_w11941_,
		_w11945_,
		_w22396_
	);
	LUT3 #(
		.INIT('h80)
	) name11884 (
		\wishbone_bd_ram_mem0_reg[62][2]/P0001 ,
		_w11948_,
		_w11979_,
		_w22397_
	);
	LUT3 #(
		.INIT('h80)
	) name11885 (
		\wishbone_bd_ram_mem0_reg[137][2]/P0001 ,
		_w11955_,
		_w11968_,
		_w22398_
	);
	LUT3 #(
		.INIT('h80)
	) name11886 (
		\wishbone_bd_ram_mem0_reg[93][2]/P0001 ,
		_w11966_,
		_w11972_,
		_w22399_
	);
	LUT4 #(
		.INIT('h0001)
	) name11887 (
		_w22396_,
		_w22397_,
		_w22398_,
		_w22399_,
		_w22400_
	);
	LUT4 #(
		.INIT('h8000)
	) name11888 (
		_w22385_,
		_w22390_,
		_w22395_,
		_w22400_,
		_w22401_
	);
	LUT3 #(
		.INIT('h80)
	) name11889 (
		\wishbone_bd_ram_mem0_reg[3][2]/P0001 ,
		_w11932_,
		_w11938_,
		_w22402_
	);
	LUT3 #(
		.INIT('h80)
	) name11890 (
		\wishbone_bd_ram_mem0_reg[10][2]/P0001 ,
		_w11932_,
		_w11944_,
		_w22403_
	);
	LUT3 #(
		.INIT('h80)
	) name11891 (
		\wishbone_bd_ram_mem0_reg[12][2]/P0001 ,
		_w11932_,
		_w11954_,
		_w22404_
	);
	LUT3 #(
		.INIT('h80)
	) name11892 (
		\wishbone_bd_ram_mem0_reg[109][2]/P0001 ,
		_w11965_,
		_w11966_,
		_w22405_
	);
	LUT4 #(
		.INIT('h0001)
	) name11893 (
		_w22402_,
		_w22403_,
		_w22404_,
		_w22405_,
		_w22406_
	);
	LUT3 #(
		.INIT('h80)
	) name11894 (
		\wishbone_bd_ram_mem0_reg[150][2]/P0001 ,
		_w11959_,
		_w11986_,
		_w22407_
	);
	LUT3 #(
		.INIT('h80)
	) name11895 (
		\wishbone_bd_ram_mem0_reg[253][2]/P0001 ,
		_w11952_,
		_w11966_,
		_w22408_
	);
	LUT3 #(
		.INIT('h80)
	) name11896 (
		\wishbone_bd_ram_mem0_reg[159][2]/P0001 ,
		_w11959_,
		_w11973_,
		_w22409_
	);
	LUT3 #(
		.INIT('h80)
	) name11897 (
		\wishbone_bd_ram_mem0_reg[138][2]/P0001 ,
		_w11944_,
		_w11955_,
		_w22410_
	);
	LUT4 #(
		.INIT('h0001)
	) name11898 (
		_w22407_,
		_w22408_,
		_w22409_,
		_w22410_,
		_w22411_
	);
	LUT3 #(
		.INIT('h80)
	) name11899 (
		\wishbone_bd_ram_mem0_reg[175][2]/P0001 ,
		_w11930_,
		_w11973_,
		_w22412_
	);
	LUT3 #(
		.INIT('h80)
	) name11900 (
		\wishbone_bd_ram_mem0_reg[229][2]/P0001 ,
		_w11933_,
		_w11982_,
		_w22413_
	);
	LUT3 #(
		.INIT('h80)
	) name11901 (
		\wishbone_bd_ram_mem0_reg[51][2]/P0001 ,
		_w11938_,
		_w11979_,
		_w22414_
	);
	LUT3 #(
		.INIT('h80)
	) name11902 (
		\wishbone_bd_ram_mem0_reg[250][2]/P0001 ,
		_w11944_,
		_w11952_,
		_w22415_
	);
	LUT4 #(
		.INIT('h0001)
	) name11903 (
		_w22412_,
		_w22413_,
		_w22414_,
		_w22415_,
		_w22416_
	);
	LUT3 #(
		.INIT('h80)
	) name11904 (
		\wishbone_bd_ram_mem0_reg[191][2]/P0001 ,
		_w11942_,
		_w11973_,
		_w22417_
	);
	LUT3 #(
		.INIT('h80)
	) name11905 (
		\wishbone_bd_ram_mem0_reg[202][2]/P0001 ,
		_w11944_,
		_w11945_,
		_w22418_
	);
	LUT3 #(
		.INIT('h80)
	) name11906 (
		\wishbone_bd_ram_mem0_reg[180][2]/P0001 ,
		_w11929_,
		_w11942_,
		_w22419_
	);
	LUT3 #(
		.INIT('h80)
	) name11907 (
		\wishbone_bd_ram_mem0_reg[119][2]/P0001 ,
		_w11975_,
		_w12012_,
		_w22420_
	);
	LUT4 #(
		.INIT('h0001)
	) name11908 (
		_w22417_,
		_w22418_,
		_w22419_,
		_w22420_,
		_w22421_
	);
	LUT4 #(
		.INIT('h8000)
	) name11909 (
		_w22406_,
		_w22411_,
		_w22416_,
		_w22421_,
		_w22422_
	);
	LUT4 #(
		.INIT('h8000)
	) name11910 (
		_w22359_,
		_w22380_,
		_w22401_,
		_w22422_,
		_w22423_
	);
	LUT3 #(
		.INIT('h80)
	) name11911 (
		\wishbone_bd_ram_mem0_reg[9][2]/P0001 ,
		_w11932_,
		_w11968_,
		_w22424_
	);
	LUT3 #(
		.INIT('h80)
	) name11912 (
		\wishbone_bd_ram_mem0_reg[69][2]/P0001 ,
		_w11933_,
		_w11949_,
		_w22425_
	);
	LUT3 #(
		.INIT('h80)
	) name11913 (
		\wishbone_bd_ram_mem0_reg[218][2]/P0001 ,
		_w11944_,
		_w11984_,
		_w22426_
	);
	LUT3 #(
		.INIT('h80)
	) name11914 (
		\wishbone_bd_ram_mem0_reg[225][2]/P0001 ,
		_w11977_,
		_w11982_,
		_w22427_
	);
	LUT4 #(
		.INIT('h0001)
	) name11915 (
		_w22424_,
		_w22425_,
		_w22426_,
		_w22427_,
		_w22428_
	);
	LUT3 #(
		.INIT('h80)
	) name11916 (
		\wishbone_bd_ram_mem0_reg[20][2]/P0001 ,
		_w11929_,
		_w11935_,
		_w22429_
	);
	LUT3 #(
		.INIT('h80)
	) name11917 (
		\wishbone_bd_ram_mem0_reg[67][2]/P0001 ,
		_w11938_,
		_w11949_,
		_w22430_
	);
	LUT3 #(
		.INIT('h80)
	) name11918 (
		\wishbone_bd_ram_mem0_reg[181][2]/P0001 ,
		_w11933_,
		_w11942_,
		_w22431_
	);
	LUT3 #(
		.INIT('h80)
	) name11919 (
		\wishbone_bd_ram_mem0_reg[155][2]/P0001 ,
		_w11936_,
		_w11959_,
		_w22432_
	);
	LUT4 #(
		.INIT('h0001)
	) name11920 (
		_w22429_,
		_w22430_,
		_w22431_,
		_w22432_,
		_w22433_
	);
	LUT3 #(
		.INIT('h80)
	) name11921 (
		\wishbone_bd_ram_mem0_reg[144][2]/P0001 ,
		_w11941_,
		_w11959_,
		_w22434_
	);
	LUT3 #(
		.INIT('h80)
	) name11922 (
		\wishbone_bd_ram_mem0_reg[33][2]/P0001 ,
		_w11957_,
		_w11977_,
		_w22435_
	);
	LUT3 #(
		.INIT('h80)
	) name11923 (
		\wishbone_bd_ram_mem0_reg[209][2]/P0001 ,
		_w11977_,
		_w11984_,
		_w22436_
	);
	LUT3 #(
		.INIT('h80)
	) name11924 (
		\wishbone_bd_ram_mem0_reg[165][2]/P0001 ,
		_w11930_,
		_w11933_,
		_w22437_
	);
	LUT4 #(
		.INIT('h0001)
	) name11925 (
		_w22434_,
		_w22435_,
		_w22436_,
		_w22437_,
		_w22438_
	);
	LUT3 #(
		.INIT('h80)
	) name11926 (
		\wishbone_bd_ram_mem0_reg[128][2]/P0001 ,
		_w11941_,
		_w11955_,
		_w22439_
	);
	LUT3 #(
		.INIT('h80)
	) name11927 (
		\wishbone_bd_ram_mem0_reg[182][2]/P0001 ,
		_w11942_,
		_w11986_,
		_w22440_
	);
	LUT3 #(
		.INIT('h80)
	) name11928 (
		\wishbone_bd_ram_mem0_reg[158][2]/P0001 ,
		_w11948_,
		_w11959_,
		_w22441_
	);
	LUT3 #(
		.INIT('h80)
	) name11929 (
		\wishbone_bd_ram_mem0_reg[148][2]/P0001 ,
		_w11929_,
		_w11959_,
		_w22442_
	);
	LUT4 #(
		.INIT('h0001)
	) name11930 (
		_w22439_,
		_w22440_,
		_w22441_,
		_w22442_,
		_w22443_
	);
	LUT4 #(
		.INIT('h8000)
	) name11931 (
		_w22428_,
		_w22433_,
		_w22438_,
		_w22443_,
		_w22444_
	);
	LUT3 #(
		.INIT('h80)
	) name11932 (
		\wishbone_bd_ram_mem0_reg[252][2]/P0001 ,
		_w11952_,
		_w11954_,
		_w22445_
	);
	LUT3 #(
		.INIT('h80)
	) name11933 (
		\wishbone_bd_ram_mem0_reg[152][2]/P0001 ,
		_w11959_,
		_w11990_,
		_w22446_
	);
	LUT3 #(
		.INIT('h80)
	) name11934 (
		\wishbone_bd_ram_mem0_reg[5][2]/P0001 ,
		_w11932_,
		_w11933_,
		_w22447_
	);
	LUT3 #(
		.INIT('h80)
	) name11935 (
		\wishbone_bd_ram_mem0_reg[120][2]/P0001 ,
		_w11990_,
		_w12012_,
		_w22448_
	);
	LUT4 #(
		.INIT('h0001)
	) name11936 (
		_w22445_,
		_w22446_,
		_w22447_,
		_w22448_,
		_w22449_
	);
	LUT3 #(
		.INIT('h80)
	) name11937 (
		\wishbone_bd_ram_mem0_reg[226][2]/P0001 ,
		_w11963_,
		_w11982_,
		_w22450_
	);
	LUT3 #(
		.INIT('h80)
	) name11938 (
		\wishbone_bd_ram_mem0_reg[139][2]/P0001 ,
		_w11936_,
		_w11955_,
		_w22451_
	);
	LUT3 #(
		.INIT('h80)
	) name11939 (
		\wishbone_bd_ram_mem0_reg[105][2]/P0001 ,
		_w11965_,
		_w11968_,
		_w22452_
	);
	LUT3 #(
		.INIT('h80)
	) name11940 (
		\wishbone_bd_ram_mem0_reg[162][2]/P0001 ,
		_w11930_,
		_w11963_,
		_w22453_
	);
	LUT4 #(
		.INIT('h0001)
	) name11941 (
		_w22450_,
		_w22451_,
		_w22452_,
		_w22453_,
		_w22454_
	);
	LUT3 #(
		.INIT('h80)
	) name11942 (
		\wishbone_bd_ram_mem0_reg[161][2]/P0001 ,
		_w11930_,
		_w11977_,
		_w22455_
	);
	LUT3 #(
		.INIT('h80)
	) name11943 (
		\wishbone_bd_ram_mem0_reg[40][2]/P0001 ,
		_w11957_,
		_w11990_,
		_w22456_
	);
	LUT3 #(
		.INIT('h80)
	) name11944 (
		\wishbone_bd_ram_mem0_reg[14][2]/P0001 ,
		_w11932_,
		_w11948_,
		_w22457_
	);
	LUT3 #(
		.INIT('h80)
	) name11945 (
		\wishbone_bd_ram_mem0_reg[6][2]/P0001 ,
		_w11932_,
		_w11986_,
		_w22458_
	);
	LUT4 #(
		.INIT('h0001)
	) name11946 (
		_w22455_,
		_w22456_,
		_w22457_,
		_w22458_,
		_w22459_
	);
	LUT3 #(
		.INIT('h80)
	) name11947 (
		\wishbone_bd_ram_mem0_reg[66][2]/P0001 ,
		_w11949_,
		_w11963_,
		_w22460_
	);
	LUT3 #(
		.INIT('h80)
	) name11948 (
		\wishbone_bd_ram_mem0_reg[55][2]/P0001 ,
		_w11975_,
		_w11979_,
		_w22461_
	);
	LUT3 #(
		.INIT('h80)
	) name11949 (
		\wishbone_bd_ram_mem0_reg[15][2]/P0001 ,
		_w11932_,
		_w11973_,
		_w22462_
	);
	LUT3 #(
		.INIT('h80)
	) name11950 (
		\wishbone_bd_ram_mem0_reg[116][2]/P0001 ,
		_w11929_,
		_w12012_,
		_w22463_
	);
	LUT4 #(
		.INIT('h0001)
	) name11951 (
		_w22460_,
		_w22461_,
		_w22462_,
		_w22463_,
		_w22464_
	);
	LUT4 #(
		.INIT('h8000)
	) name11952 (
		_w22449_,
		_w22454_,
		_w22459_,
		_w22464_,
		_w22465_
	);
	LUT3 #(
		.INIT('h80)
	) name11953 (
		\wishbone_bd_ram_mem0_reg[172][2]/P0001 ,
		_w11930_,
		_w11954_,
		_w22466_
	);
	LUT3 #(
		.INIT('h80)
	) name11954 (
		\wishbone_bd_ram_mem0_reg[83][2]/P0001 ,
		_w11938_,
		_w11972_,
		_w22467_
	);
	LUT3 #(
		.INIT('h80)
	) name11955 (
		\wishbone_bd_ram_mem0_reg[21][2]/P0001 ,
		_w11933_,
		_w11935_,
		_w22468_
	);
	LUT3 #(
		.INIT('h80)
	) name11956 (
		\wishbone_bd_ram_mem0_reg[127][2]/P0001 ,
		_w11973_,
		_w12012_,
		_w22469_
	);
	LUT4 #(
		.INIT('h0001)
	) name11957 (
		_w22466_,
		_w22467_,
		_w22468_,
		_w22469_,
		_w22470_
	);
	LUT3 #(
		.INIT('h80)
	) name11958 (
		\wishbone_bd_ram_mem0_reg[217][2]/P0001 ,
		_w11968_,
		_w11984_,
		_w22471_
	);
	LUT3 #(
		.INIT('h80)
	) name11959 (
		\wishbone_bd_ram_mem0_reg[147][2]/P0001 ,
		_w11938_,
		_w11959_,
		_w22472_
	);
	LUT3 #(
		.INIT('h80)
	) name11960 (
		\wishbone_bd_ram_mem0_reg[208][2]/P0001 ,
		_w11941_,
		_w11984_,
		_w22473_
	);
	LUT3 #(
		.INIT('h80)
	) name11961 (
		\wishbone_bd_ram_mem0_reg[115][2]/P0001 ,
		_w11938_,
		_w12012_,
		_w22474_
	);
	LUT4 #(
		.INIT('h0001)
	) name11962 (
		_w22471_,
		_w22472_,
		_w22473_,
		_w22474_,
		_w22475_
	);
	LUT3 #(
		.INIT('h80)
	) name11963 (
		\wishbone_bd_ram_mem0_reg[68][2]/P0001 ,
		_w11929_,
		_w11949_,
		_w22476_
	);
	LUT3 #(
		.INIT('h80)
	) name11964 (
		\wishbone_bd_ram_mem0_reg[176][2]/P0001 ,
		_w11941_,
		_w11942_,
		_w22477_
	);
	LUT3 #(
		.INIT('h80)
	) name11965 (
		\wishbone_bd_ram_mem0_reg[78][2]/P0001 ,
		_w11948_,
		_w11949_,
		_w22478_
	);
	LUT3 #(
		.INIT('h80)
	) name11966 (
		\wishbone_bd_ram_mem0_reg[151][2]/P0001 ,
		_w11959_,
		_w11975_,
		_w22479_
	);
	LUT4 #(
		.INIT('h0001)
	) name11967 (
		_w22476_,
		_w22477_,
		_w22478_,
		_w22479_,
		_w22480_
	);
	LUT3 #(
		.INIT('h80)
	) name11968 (
		\wishbone_bd_ram_mem0_reg[141][2]/P0001 ,
		_w11955_,
		_w11966_,
		_w22481_
	);
	LUT3 #(
		.INIT('h80)
	) name11969 (
		\wishbone_bd_ram_mem0_reg[54][2]/P0001 ,
		_w11979_,
		_w11986_,
		_w22482_
	);
	LUT3 #(
		.INIT('h80)
	) name11970 (
		\wishbone_bd_ram_mem0_reg[81][2]/P0001 ,
		_w11972_,
		_w11977_,
		_w22483_
	);
	LUT3 #(
		.INIT('h80)
	) name11971 (
		\wishbone_bd_ram_mem0_reg[22][2]/P0001 ,
		_w11935_,
		_w11986_,
		_w22484_
	);
	LUT4 #(
		.INIT('h0001)
	) name11972 (
		_w22481_,
		_w22482_,
		_w22483_,
		_w22484_,
		_w22485_
	);
	LUT4 #(
		.INIT('h8000)
	) name11973 (
		_w22470_,
		_w22475_,
		_w22480_,
		_w22485_,
		_w22486_
	);
	LUT3 #(
		.INIT('h80)
	) name11974 (
		\wishbone_bd_ram_mem0_reg[126][2]/P0001 ,
		_w11948_,
		_w12012_,
		_w22487_
	);
	LUT3 #(
		.INIT('h80)
	) name11975 (
		\wishbone_bd_ram_mem0_reg[211][2]/P0001 ,
		_w11938_,
		_w11984_,
		_w22488_
	);
	LUT3 #(
		.INIT('h80)
	) name11976 (
		\wishbone_bd_ram_mem0_reg[63][2]/P0001 ,
		_w11973_,
		_w11979_,
		_w22489_
	);
	LUT3 #(
		.INIT('h80)
	) name11977 (
		\wishbone_bd_ram_mem0_reg[239][2]/P0001 ,
		_w11973_,
		_w11982_,
		_w22490_
	);
	LUT4 #(
		.INIT('h0001)
	) name11978 (
		_w22487_,
		_w22488_,
		_w22489_,
		_w22490_,
		_w22491_
	);
	LUT3 #(
		.INIT('h80)
	) name11979 (
		\wishbone_bd_ram_mem0_reg[17][2]/P0001 ,
		_w11935_,
		_w11977_,
		_w22492_
	);
	LUT3 #(
		.INIT('h80)
	) name11980 (
		\wishbone_bd_ram_mem0_reg[205][2]/P0001 ,
		_w11945_,
		_w11966_,
		_w22493_
	);
	LUT3 #(
		.INIT('h80)
	) name11981 (
		\wishbone_bd_ram_mem0_reg[187][2]/P0001 ,
		_w11936_,
		_w11942_,
		_w22494_
	);
	LUT3 #(
		.INIT('h80)
	) name11982 (
		\wishbone_bd_ram_mem0_reg[204][2]/P0001 ,
		_w11945_,
		_w11954_,
		_w22495_
	);
	LUT4 #(
		.INIT('h0001)
	) name11983 (
		_w22492_,
		_w22493_,
		_w22494_,
		_w22495_,
		_w22496_
	);
	LUT3 #(
		.INIT('h80)
	) name11984 (
		\wishbone_bd_ram_mem0_reg[201][2]/P0001 ,
		_w11945_,
		_w11968_,
		_w22497_
	);
	LUT3 #(
		.INIT('h80)
	) name11985 (
		\wishbone_bd_ram_mem0_reg[173][2]/P0001 ,
		_w11930_,
		_w11966_,
		_w22498_
	);
	LUT3 #(
		.INIT('h80)
	) name11986 (
		\wishbone_bd_ram_mem0_reg[75][2]/P0001 ,
		_w11936_,
		_w11949_,
		_w22499_
	);
	LUT3 #(
		.INIT('h80)
	) name11987 (
		\wishbone_bd_ram_mem0_reg[94][2]/P0001 ,
		_w11948_,
		_w11972_,
		_w22500_
	);
	LUT4 #(
		.INIT('h0001)
	) name11988 (
		_w22497_,
		_w22498_,
		_w22499_,
		_w22500_,
		_w22501_
	);
	LUT3 #(
		.INIT('h80)
	) name11989 (
		\wishbone_bd_ram_mem0_reg[122][2]/P0001 ,
		_w11944_,
		_w12012_,
		_w22502_
	);
	LUT3 #(
		.INIT('h80)
	) name11990 (
		\wishbone_bd_ram_mem0_reg[29][2]/P0001 ,
		_w11935_,
		_w11966_,
		_w22503_
	);
	LUT3 #(
		.INIT('h80)
	) name11991 (
		\wishbone_bd_ram_mem0_reg[65][2]/P0001 ,
		_w11949_,
		_w11977_,
		_w22504_
	);
	LUT3 #(
		.INIT('h80)
	) name11992 (
		\wishbone_bd_ram_mem0_reg[18][2]/P0001 ,
		_w11935_,
		_w11963_,
		_w22505_
	);
	LUT4 #(
		.INIT('h0001)
	) name11993 (
		_w22502_,
		_w22503_,
		_w22504_,
		_w22505_,
		_w22506_
	);
	LUT4 #(
		.INIT('h8000)
	) name11994 (
		_w22491_,
		_w22496_,
		_w22501_,
		_w22506_,
		_w22507_
	);
	LUT4 #(
		.INIT('h8000)
	) name11995 (
		_w22444_,
		_w22465_,
		_w22486_,
		_w22507_,
		_w22508_
	);
	LUT3 #(
		.INIT('h80)
	) name11996 (
		\wishbone_bd_ram_mem0_reg[134][2]/P0001 ,
		_w11955_,
		_w11986_,
		_w22509_
	);
	LUT3 #(
		.INIT('h80)
	) name11997 (
		\wishbone_bd_ram_mem0_reg[111][2]/P0001 ,
		_w11965_,
		_w11973_,
		_w22510_
	);
	LUT3 #(
		.INIT('h80)
	) name11998 (
		\wishbone_bd_ram_mem0_reg[129][2]/P0001 ,
		_w11955_,
		_w11977_,
		_w22511_
	);
	LUT3 #(
		.INIT('h80)
	) name11999 (
		\wishbone_bd_ram_mem0_reg[92][2]/P0001 ,
		_w11954_,
		_w11972_,
		_w22512_
	);
	LUT4 #(
		.INIT('h0001)
	) name12000 (
		_w22509_,
		_w22510_,
		_w22511_,
		_w22512_,
		_w22513_
	);
	LUT3 #(
		.INIT('h80)
	) name12001 (
		\wishbone_bd_ram_mem0_reg[107][2]/P0001 ,
		_w11936_,
		_w11965_,
		_w22514_
	);
	LUT3 #(
		.INIT('h80)
	) name12002 (
		\wishbone_bd_ram_mem0_reg[101][2]/P0001 ,
		_w11933_,
		_w11965_,
		_w22515_
	);
	LUT3 #(
		.INIT('h80)
	) name12003 (
		\wishbone_bd_ram_mem0_reg[184][2]/P0001 ,
		_w11942_,
		_w11990_,
		_w22516_
	);
	LUT3 #(
		.INIT('h80)
	) name12004 (
		\wishbone_bd_ram_mem0_reg[215][2]/P0001 ,
		_w11975_,
		_w11984_,
		_w22517_
	);
	LUT4 #(
		.INIT('h0001)
	) name12005 (
		_w22514_,
		_w22515_,
		_w22516_,
		_w22517_,
		_w22518_
	);
	LUT3 #(
		.INIT('h80)
	) name12006 (
		\wishbone_bd_ram_mem0_reg[99][2]/P0001 ,
		_w11938_,
		_w11965_,
		_w22519_
	);
	LUT3 #(
		.INIT('h80)
	) name12007 (
		\wishbone_bd_ram_mem0_reg[213][2]/P0001 ,
		_w11933_,
		_w11984_,
		_w22520_
	);
	LUT3 #(
		.INIT('h80)
	) name12008 (
		\wishbone_bd_ram_mem0_reg[41][2]/P0001 ,
		_w11957_,
		_w11968_,
		_w22521_
	);
	LUT3 #(
		.INIT('h80)
	) name12009 (
		\wishbone_bd_ram_mem0_reg[220][2]/P0001 ,
		_w11954_,
		_w11984_,
		_w22522_
	);
	LUT4 #(
		.INIT('h0001)
	) name12010 (
		_w22519_,
		_w22520_,
		_w22521_,
		_w22522_,
		_w22523_
	);
	LUT3 #(
		.INIT('h80)
	) name12011 (
		\wishbone_bd_ram_mem0_reg[46][2]/P0001 ,
		_w11948_,
		_w11957_,
		_w22524_
	);
	LUT3 #(
		.INIT('h80)
	) name12012 (
		\wishbone_bd_ram_mem0_reg[4][2]/P0001 ,
		_w11929_,
		_w11932_,
		_w22525_
	);
	LUT3 #(
		.INIT('h80)
	) name12013 (
		\wishbone_bd_ram_mem0_reg[168][2]/P0001 ,
		_w11930_,
		_w11990_,
		_w22526_
	);
	LUT3 #(
		.INIT('h80)
	) name12014 (
		\wishbone_bd_ram_mem0_reg[56][2]/P0001 ,
		_w11979_,
		_w11990_,
		_w22527_
	);
	LUT4 #(
		.INIT('h0001)
	) name12015 (
		_w22524_,
		_w22525_,
		_w22526_,
		_w22527_,
		_w22528_
	);
	LUT4 #(
		.INIT('h8000)
	) name12016 (
		_w22513_,
		_w22518_,
		_w22523_,
		_w22528_,
		_w22529_
	);
	LUT3 #(
		.INIT('h80)
	) name12017 (
		\wishbone_bd_ram_mem0_reg[89][2]/P0001 ,
		_w11968_,
		_w11972_,
		_w22530_
	);
	LUT3 #(
		.INIT('h80)
	) name12018 (
		\wishbone_bd_ram_mem0_reg[74][2]/P0001 ,
		_w11944_,
		_w11949_,
		_w22531_
	);
	LUT3 #(
		.INIT('h80)
	) name12019 (
		\wishbone_bd_ram_mem0_reg[203][2]/P0001 ,
		_w11936_,
		_w11945_,
		_w22532_
	);
	LUT3 #(
		.INIT('h80)
	) name12020 (
		\wishbone_bd_ram_mem0_reg[90][2]/P0001 ,
		_w11944_,
		_w11972_,
		_w22533_
	);
	LUT4 #(
		.INIT('h0001)
	) name12021 (
		_w22530_,
		_w22531_,
		_w22532_,
		_w22533_,
		_w22534_
	);
	LUT3 #(
		.INIT('h80)
	) name12022 (
		\wishbone_bd_ram_mem0_reg[171][2]/P0001 ,
		_w11930_,
		_w11936_,
		_w22535_
	);
	LUT3 #(
		.INIT('h80)
	) name12023 (
		\wishbone_bd_ram_mem0_reg[156][2]/P0001 ,
		_w11954_,
		_w11959_,
		_w22536_
	);
	LUT3 #(
		.INIT('h80)
	) name12024 (
		\wishbone_bd_ram_mem0_reg[32][2]/P0001 ,
		_w11941_,
		_w11957_,
		_w22537_
	);
	LUT3 #(
		.INIT('h80)
	) name12025 (
		\wishbone_bd_ram_mem0_reg[35][2]/P0001 ,
		_w11938_,
		_w11957_,
		_w22538_
	);
	LUT4 #(
		.INIT('h0001)
	) name12026 (
		_w22535_,
		_w22536_,
		_w22537_,
		_w22538_,
		_w22539_
	);
	LUT3 #(
		.INIT('h80)
	) name12027 (
		\wishbone_bd_ram_mem0_reg[185][2]/P0001 ,
		_w11942_,
		_w11968_,
		_w22540_
	);
	LUT3 #(
		.INIT('h80)
	) name12028 (
		\wishbone_bd_ram_mem0_reg[110][2]/P0001 ,
		_w11948_,
		_w11965_,
		_w22541_
	);
	LUT3 #(
		.INIT('h80)
	) name12029 (
		\wishbone_bd_ram_mem0_reg[232][2]/P0001 ,
		_w11982_,
		_w11990_,
		_w22542_
	);
	LUT3 #(
		.INIT('h80)
	) name12030 (
		\wishbone_bd_ram_mem0_reg[61][2]/P0001 ,
		_w11966_,
		_w11979_,
		_w22543_
	);
	LUT4 #(
		.INIT('h0001)
	) name12031 (
		_w22540_,
		_w22541_,
		_w22542_,
		_w22543_,
		_w22544_
	);
	LUT3 #(
		.INIT('h80)
	) name12032 (
		\wishbone_bd_ram_mem0_reg[27][2]/P0001 ,
		_w11935_,
		_w11936_,
		_w22545_
	);
	LUT3 #(
		.INIT('h80)
	) name12033 (
		\wishbone_bd_ram_mem0_reg[77][2]/P0001 ,
		_w11949_,
		_w11966_,
		_w22546_
	);
	LUT3 #(
		.INIT('h80)
	) name12034 (
		\wishbone_bd_ram_mem0_reg[216][2]/P0001 ,
		_w11984_,
		_w11990_,
		_w22547_
	);
	LUT3 #(
		.INIT('h80)
	) name12035 (
		\wishbone_bd_ram_mem0_reg[167][2]/P0001 ,
		_w11930_,
		_w11975_,
		_w22548_
	);
	LUT4 #(
		.INIT('h0001)
	) name12036 (
		_w22545_,
		_w22546_,
		_w22547_,
		_w22548_,
		_w22549_
	);
	LUT4 #(
		.INIT('h8000)
	) name12037 (
		_w22534_,
		_w22539_,
		_w22544_,
		_w22549_,
		_w22550_
	);
	LUT3 #(
		.INIT('h80)
	) name12038 (
		\wishbone_bd_ram_mem0_reg[247][2]/P0001 ,
		_w11952_,
		_w11975_,
		_w22551_
	);
	LUT3 #(
		.INIT('h80)
	) name12039 (
		\wishbone_bd_ram_mem0_reg[58][2]/P0001 ,
		_w11944_,
		_w11979_,
		_w22552_
	);
	LUT3 #(
		.INIT('h80)
	) name12040 (
		\wishbone_bd_ram_mem0_reg[197][2]/P0001 ,
		_w11933_,
		_w11945_,
		_w22553_
	);
	LUT3 #(
		.INIT('h80)
	) name12041 (
		\wishbone_bd_ram_mem0_reg[234][2]/P0001 ,
		_w11944_,
		_w11982_,
		_w22554_
	);
	LUT4 #(
		.INIT('h0001)
	) name12042 (
		_w22551_,
		_w22552_,
		_w22553_,
		_w22554_,
		_w22555_
	);
	LUT3 #(
		.INIT('h80)
	) name12043 (
		\wishbone_bd_ram_mem0_reg[19][2]/P0001 ,
		_w11935_,
		_w11938_,
		_w22556_
	);
	LUT3 #(
		.INIT('h80)
	) name12044 (
		\wishbone_bd_ram_mem0_reg[37][2]/P0001 ,
		_w11933_,
		_w11957_,
		_w22557_
	);
	LUT3 #(
		.INIT('h80)
	) name12045 (
		\wishbone_bd_ram_mem0_reg[123][2]/P0001 ,
		_w11936_,
		_w12012_,
		_w22558_
	);
	LUT3 #(
		.INIT('h80)
	) name12046 (
		\wishbone_bd_ram_mem0_reg[244][2]/P0001 ,
		_w11929_,
		_w11952_,
		_w22559_
	);
	LUT4 #(
		.INIT('h0001)
	) name12047 (
		_w22556_,
		_w22557_,
		_w22558_,
		_w22559_,
		_w22560_
	);
	LUT3 #(
		.INIT('h80)
	) name12048 (
		\wishbone_bd_ram_mem0_reg[79][2]/P0001 ,
		_w11949_,
		_w11973_,
		_w22561_
	);
	LUT3 #(
		.INIT('h80)
	) name12049 (
		\wishbone_bd_ram_mem0_reg[71][2]/P0001 ,
		_w11949_,
		_w11975_,
		_w22562_
	);
	LUT3 #(
		.INIT('h80)
	) name12050 (
		\wishbone_bd_ram_mem0_reg[30][2]/P0001 ,
		_w11935_,
		_w11948_,
		_w22563_
	);
	LUT3 #(
		.INIT('h80)
	) name12051 (
		\wishbone_bd_ram_mem0_reg[133][2]/P0001 ,
		_w11933_,
		_w11955_,
		_w22564_
	);
	LUT4 #(
		.INIT('h0001)
	) name12052 (
		_w22561_,
		_w22562_,
		_w22563_,
		_w22564_,
		_w22565_
	);
	LUT3 #(
		.INIT('h80)
	) name12053 (
		\wishbone_bd_ram_mem0_reg[254][2]/P0001 ,
		_w11948_,
		_w11952_,
		_w22566_
	);
	LUT3 #(
		.INIT('h80)
	) name12054 (
		\wishbone_bd_ram_mem0_reg[230][2]/P0001 ,
		_w11982_,
		_w11986_,
		_w22567_
	);
	LUT3 #(
		.INIT('h80)
	) name12055 (
		\wishbone_bd_ram_mem0_reg[227][2]/P0001 ,
		_w11938_,
		_w11982_,
		_w22568_
	);
	LUT3 #(
		.INIT('h80)
	) name12056 (
		\wishbone_bd_ram_mem0_reg[52][2]/P0001 ,
		_w11929_,
		_w11979_,
		_w22569_
	);
	LUT4 #(
		.INIT('h0001)
	) name12057 (
		_w22566_,
		_w22567_,
		_w22568_,
		_w22569_,
		_w22570_
	);
	LUT4 #(
		.INIT('h8000)
	) name12058 (
		_w22555_,
		_w22560_,
		_w22565_,
		_w22570_,
		_w22571_
	);
	LUT3 #(
		.INIT('h80)
	) name12059 (
		\wishbone_bd_ram_mem0_reg[125][2]/P0001 ,
		_w11966_,
		_w12012_,
		_w22572_
	);
	LUT3 #(
		.INIT('h80)
	) name12060 (
		\wishbone_bd_ram_mem0_reg[45][2]/P0001 ,
		_w11957_,
		_w11966_,
		_w22573_
	);
	LUT3 #(
		.INIT('h80)
	) name12061 (
		\wishbone_bd_ram_mem0_reg[106][2]/P0001 ,
		_w11944_,
		_w11965_,
		_w22574_
	);
	LUT3 #(
		.INIT('h80)
	) name12062 (
		\wishbone_bd_ram_mem0_reg[130][2]/P0001 ,
		_w11955_,
		_w11963_,
		_w22575_
	);
	LUT4 #(
		.INIT('h0001)
	) name12063 (
		_w22572_,
		_w22573_,
		_w22574_,
		_w22575_,
		_w22576_
	);
	LUT3 #(
		.INIT('h80)
	) name12064 (
		\wishbone_bd_ram_mem0_reg[53][2]/P0001 ,
		_w11933_,
		_w11979_,
		_w22577_
	);
	LUT3 #(
		.INIT('h80)
	) name12065 (
		\wishbone_bd_ram_mem0_reg[49][2]/P0001 ,
		_w11977_,
		_w11979_,
		_w22578_
	);
	LUT3 #(
		.INIT('h80)
	) name12066 (
		\wishbone_bd_ram_mem0_reg[117][2]/P0001 ,
		_w11933_,
		_w12012_,
		_w22579_
	);
	LUT3 #(
		.INIT('h80)
	) name12067 (
		\wishbone_bd_ram_mem0_reg[177][2]/P0001 ,
		_w11942_,
		_w11977_,
		_w22580_
	);
	LUT4 #(
		.INIT('h0001)
	) name12068 (
		_w22577_,
		_w22578_,
		_w22579_,
		_w22580_,
		_w22581_
	);
	LUT3 #(
		.INIT('h80)
	) name12069 (
		\wishbone_bd_ram_mem0_reg[36][2]/P0001 ,
		_w11929_,
		_w11957_,
		_w22582_
	);
	LUT3 #(
		.INIT('h80)
	) name12070 (
		\wishbone_bd_ram_mem0_reg[251][2]/P0001 ,
		_w11936_,
		_w11952_,
		_w22583_
	);
	LUT3 #(
		.INIT('h80)
	) name12071 (
		\wishbone_bd_ram_mem0_reg[241][2]/P0001 ,
		_w11952_,
		_w11977_,
		_w22584_
	);
	LUT3 #(
		.INIT('h80)
	) name12072 (
		\wishbone_bd_ram_mem0_reg[97][2]/P0001 ,
		_w11965_,
		_w11977_,
		_w22585_
	);
	LUT4 #(
		.INIT('h0001)
	) name12073 (
		_w22582_,
		_w22583_,
		_w22584_,
		_w22585_,
		_w22586_
	);
	LUT3 #(
		.INIT('h80)
	) name12074 (
		\wishbone_bd_ram_mem0_reg[48][2]/P0001 ,
		_w11941_,
		_w11979_,
		_w22587_
	);
	LUT3 #(
		.INIT('h80)
	) name12075 (
		\wishbone_bd_ram_mem0_reg[154][2]/P0001 ,
		_w11944_,
		_w11959_,
		_w22588_
	);
	LUT3 #(
		.INIT('h80)
	) name12076 (
		\wishbone_bd_ram_mem0_reg[0][2]/P0001 ,
		_w11932_,
		_w11941_,
		_w22589_
	);
	LUT3 #(
		.INIT('h80)
	) name12077 (
		\wishbone_bd_ram_mem0_reg[243][2]/P0001 ,
		_w11938_,
		_w11952_,
		_w22590_
	);
	LUT4 #(
		.INIT('h0001)
	) name12078 (
		_w22587_,
		_w22588_,
		_w22589_,
		_w22590_,
		_w22591_
	);
	LUT4 #(
		.INIT('h8000)
	) name12079 (
		_w22576_,
		_w22581_,
		_w22586_,
		_w22591_,
		_w22592_
	);
	LUT4 #(
		.INIT('h8000)
	) name12080 (
		_w22529_,
		_w22550_,
		_w22571_,
		_w22592_,
		_w22593_
	);
	LUT4 #(
		.INIT('h8000)
	) name12081 (
		_w22338_,
		_w22423_,
		_w22508_,
		_w22593_,
		_w22594_
	);
	LUT3 #(
		.INIT('h15)
	) name12082 (
		wb_rst_i_pad,
		_w22235_,
		_w22252_,
		_w22595_
	);
	LUT3 #(
		.INIT('hba)
	) name12083 (
		_w22253_,
		_w22594_,
		_w22595_,
		_w22596_
	);
	LUT3 #(
		.INIT('h80)
	) name12084 (
		\ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131 ,
		_w18753_,
		_w18754_,
		_w22597_
	);
	LUT3 #(
		.INIT('h80)
	) name12085 (
		\ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131 ,
		_w18805_,
		_w19655_,
		_w22598_
	);
	LUT3 #(
		.INIT('h80)
	) name12086 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[0]/NET0131 ,
		_w18798_,
		_w18801_,
		_w22599_
	);
	LUT3 #(
		.INIT('h80)
	) name12087 (
		\ethreg1_MIIMODER_0_DataOut_reg[0]/NET0131 ,
		_w18786_,
		_w18801_,
		_w22600_
	);
	LUT3 #(
		.INIT('h80)
	) name12088 (
		\ethreg1_INT_MASK_0_DataOut_reg[0]/NET0131 ,
		_w18801_,
		_w19655_,
		_w22601_
	);
	LUT4 #(
		.INIT('h0001)
	) name12089 (
		_w22598_,
		_w22599_,
		_w22600_,
		_w22601_,
		_w22602_
	);
	LUT3 #(
		.INIT('h80)
	) name12090 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[0]/NET0131 ,
		_w18785_,
		_w18798_,
		_w22603_
	);
	LUT4 #(
		.INIT('h0002)
	) name12091 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22604_
	);
	LUT3 #(
		.INIT('h80)
	) name12092 (
		_w18757_,
		_w18762_,
		_w22604_,
		_w22605_
	);
	LUT3 #(
		.INIT('h80)
	) name12093 (
		\miim1_shftrg_LinkFail_reg/NET0131 ,
		_w18786_,
		_w18805_,
		_w22606_
	);
	LUT3 #(
		.INIT('h80)
	) name12094 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[0]/NET0131 ,
		_w18798_,
		_w18805_,
		_w22607_
	);
	LUT4 #(
		.INIT('h0001)
	) name12095 (
		_w22603_,
		_w22605_,
		_w22606_,
		_w22607_,
		_w22608_
	);
	LUT3 #(
		.INIT('h40)
	) name12096 (
		_w22597_,
		_w22602_,
		_w22608_,
		_w22609_
	);
	LUT3 #(
		.INIT('h80)
	) name12097 (
		\ethreg1_IPGT_0_DataOut_reg[0]/NET0131 ,
		_w19646_,
		_w19655_,
		_w22610_
	);
	LUT4 #(
		.INIT('h0002)
	) name12098 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22611_
	);
	LUT3 #(
		.INIT('h80)
	) name12099 (
		_w18757_,
		_w18758_,
		_w22611_,
		_w22612_
	);
	LUT3 #(
		.INIT('h80)
	) name12100 (
		\ethreg1_IPGR1_0_DataOut_reg[0]/NET0131 ,
		_w18785_,
		_w18800_,
		_w22613_
	);
	LUT3 #(
		.INIT('h80)
	) name12101 (
		\ethreg1_MIIRX_DATA_DataOut_reg[0]/NET0131 ,
		_w18785_,
		_w18786_,
		_w22614_
	);
	LUT4 #(
		.INIT('h0001)
	) name12102 (
		_w22610_,
		_w22612_,
		_w22613_,
		_w22614_,
		_w22615_
	);
	LUT4 #(
		.INIT('h0008)
	) name12103 (
		\ethreg1_RXHASH1_0_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22616_
	);
	LUT3 #(
		.INIT('h80)
	) name12104 (
		_w18757_,
		_w18762_,
		_w22616_,
		_w22617_
	);
	LUT3 #(
		.INIT('h80)
	) name12105 (
		\ethreg1_MODER_0_DataOut_reg[0]/NET0131 ,
		_w18800_,
		_w18801_,
		_w22618_
	);
	LUT4 #(
		.INIT('h0008)
	) name12106 (
		\ethreg1_RXHASH0_0_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22619_
	);
	LUT3 #(
		.INIT('h80)
	) name12107 (
		_w18757_,
		_w18758_,
		_w22619_,
		_w22620_
	);
	LUT3 #(
		.INIT('h80)
	) name12108 (
		\ethreg1_IPGR2_0_DataOut_reg[0]/NET0131 ,
		_w18800_,
		_w18805_,
		_w22621_
	);
	LUT4 #(
		.INIT('h0001)
	) name12109 (
		_w22617_,
		_w22618_,
		_w22620_,
		_w22621_,
		_w22622_
	);
	LUT4 #(
		.INIT('h0020)
	) name12110 (
		\ethreg1_TXCTRL_0_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22623_
	);
	LUT3 #(
		.INIT('h80)
	) name12111 (
		_w18757_,
		_w18758_,
		_w22623_,
		_w22624_
	);
	LUT3 #(
		.INIT('h80)
	) name12112 (
		\ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131 ,
		_w18798_,
		_w19646_,
		_w22625_
	);
	LUT3 #(
		.INIT('h80)
	) name12113 (
		\ethreg1_irq_txb_reg/NET0131 ,
		_w18800_,
		_w19646_,
		_w22626_
	);
	LUT3 #(
		.INIT('h80)
	) name12114 (
		\ethreg1_MIICOMMAND0_DataOut_reg[0]/NET0131 ,
		_w18786_,
		_w19646_,
		_w22627_
	);
	LUT4 #(
		.INIT('h0001)
	) name12115 (
		_w22624_,
		_w22625_,
		_w22626_,
		_w22627_,
		_w22628_
	);
	LUT4 #(
		.INIT('h8000)
	) name12116 (
		_w18752_,
		_w22615_,
		_w22622_,
		_w22628_,
		_w22629_
	);
	LUT3 #(
		.INIT('h2a)
	) name12117 (
		_w18752_,
		_w22609_,
		_w22629_,
		_w22630_
	);
	LUT3 #(
		.INIT('h15)
	) name12118 (
		wb_rst_i_pad,
		_w22609_,
		_w22629_,
		_w22631_
	);
	LUT3 #(
		.INIT('hdc)
	) name12119 (
		_w19524_,
		_w22630_,
		_w22631_,
		_w22632_
	);
	LUT3 #(
		.INIT('h80)
	) name12120 (
		\ethreg1_irq_txe_reg/NET0131 ,
		_w18800_,
		_w19646_,
		_w22633_
	);
	LUT3 #(
		.INIT('h80)
	) name12121 (
		\ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131 ,
		_w18798_,
		_w19646_,
		_w22634_
	);
	LUT4 #(
		.INIT('h0001)
	) name12122 (
		\miim1_InProgress_reg/NET0131 ,
		\miim1_Nvalid_reg/NET0131 ,
		\miim1_RStatStart_reg/NET0131 ,
		\miim1_SyncStatMdcEn_reg/NET0131 ,
		_w22635_
	);
	LUT4 #(
		.INIT('h0001)
	) name12123 (
		\ethreg1_MIICOMMAND2_DataOut_reg[0]/NET0131 ,
		\miim1_EndBusy_reg/NET0131 ,
		\miim1_InProgress_q3_reg/NET0131 ,
		\miim1_WCtrlDataStart_reg/NET0131 ,
		_w22636_
	);
	LUT4 #(
		.INIT('h0888)
	) name12124 (
		_w18786_,
		_w18805_,
		_w22635_,
		_w22636_,
		_w22637_
	);
	LUT3 #(
		.INIT('h80)
	) name12125 (
		\ethreg1_MODER_0_DataOut_reg[1]/NET0131 ,
		_w18800_,
		_w18801_,
		_w22638_
	);
	LUT4 #(
		.INIT('h0001)
	) name12126 (
		_w22633_,
		_w22634_,
		_w22637_,
		_w22638_,
		_w22639_
	);
	LUT3 #(
		.INIT('h80)
	) name12127 (
		\ethreg1_IPGR1_0_DataOut_reg[1]/NET0131 ,
		_w18785_,
		_w18800_,
		_w22640_
	);
	LUT3 #(
		.INIT('h80)
	) name12128 (
		\ethreg1_INT_MASK_0_DataOut_reg[1]/NET0131 ,
		_w18801_,
		_w19655_,
		_w22641_
	);
	LUT3 #(
		.INIT('h80)
	) name12129 (
		\ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131 ,
		_w18753_,
		_w18754_,
		_w22642_
	);
	LUT3 #(
		.INIT('h80)
	) name12130 (
		\ethreg1_IPGT_0_DataOut_reg[1]/NET0131 ,
		_w19646_,
		_w19655_,
		_w22643_
	);
	LUT4 #(
		.INIT('h0001)
	) name12131 (
		_w22640_,
		_w22641_,
		_w22642_,
		_w22643_,
		_w22644_
	);
	LUT2 #(
		.INIT('h8)
	) name12132 (
		_w22639_,
		_w22644_,
		_w22645_
	);
	LUT3 #(
		.INIT('h80)
	) name12133 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[1]/NET0131 ,
		_w18798_,
		_w18801_,
		_w22646_
	);
	LUT4 #(
		.INIT('h0002)
	) name12134 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22647_
	);
	LUT3 #(
		.INIT('h80)
	) name12135 (
		_w18757_,
		_w18758_,
		_w22647_,
		_w22648_
	);
	LUT3 #(
		.INIT('h80)
	) name12136 (
		\ethreg1_IPGR2_0_DataOut_reg[1]/NET0131 ,
		_w18800_,
		_w18805_,
		_w22649_
	);
	LUT4 #(
		.INIT('h0008)
	) name12137 (
		\ethreg1_RXHASH0_0_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22650_
	);
	LUT3 #(
		.INIT('h80)
	) name12138 (
		_w18757_,
		_w18758_,
		_w22650_,
		_w22651_
	);
	LUT4 #(
		.INIT('h0001)
	) name12139 (
		_w22646_,
		_w22648_,
		_w22649_,
		_w22651_,
		_w22652_
	);
	LUT3 #(
		.INIT('h02)
	) name12140 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[6]_pad ,
		\wb_adr_i[8]_pad ,
		_w22653_
	);
	LUT3 #(
		.INIT('h80)
	) name12141 (
		\ethreg1_MIICOMMAND1_DataOut_reg[0]/NET0131 ,
		_w18786_,
		_w22653_,
		_w22654_
	);
	LUT2 #(
		.INIT('h2)
	) name12142 (
		_w18752_,
		_w22654_,
		_w22655_
	);
	LUT3 #(
		.INIT('h80)
	) name12143 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[1]/NET0131 ,
		_w18785_,
		_w18798_,
		_w22656_
	);
	LUT4 #(
		.INIT('h0002)
	) name12144 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22657_
	);
	LUT3 #(
		.INIT('h80)
	) name12145 (
		_w18757_,
		_w18762_,
		_w22657_,
		_w22658_
	);
	LUT3 #(
		.INIT('h80)
	) name12146 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[1]/NET0131 ,
		_w18798_,
		_w18805_,
		_w22659_
	);
	LUT3 #(
		.INIT('h80)
	) name12147 (
		\ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131 ,
		_w18805_,
		_w19655_,
		_w22660_
	);
	LUT4 #(
		.INIT('h0001)
	) name12148 (
		_w22656_,
		_w22658_,
		_w22659_,
		_w22660_,
		_w22661_
	);
	LUT4 #(
		.INIT('h0008)
	) name12149 (
		\ethreg1_RXHASH1_0_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22662_
	);
	LUT3 #(
		.INIT('h80)
	) name12150 (
		_w18757_,
		_w18762_,
		_w22662_,
		_w22663_
	);
	LUT4 #(
		.INIT('h0020)
	) name12151 (
		\ethreg1_TXCTRL_0_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22664_
	);
	LUT3 #(
		.INIT('h80)
	) name12152 (
		_w18757_,
		_w18758_,
		_w22664_,
		_w22665_
	);
	LUT3 #(
		.INIT('h80)
	) name12153 (
		\ethreg1_MIIRX_DATA_DataOut_reg[1]/NET0131 ,
		_w18785_,
		_w18786_,
		_w22666_
	);
	LUT3 #(
		.INIT('h80)
	) name12154 (
		\ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131 ,
		_w18786_,
		_w18801_,
		_w22667_
	);
	LUT4 #(
		.INIT('h0001)
	) name12155 (
		_w22663_,
		_w22665_,
		_w22666_,
		_w22667_,
		_w22668_
	);
	LUT4 #(
		.INIT('h8000)
	) name12156 (
		_w22652_,
		_w22655_,
		_w22661_,
		_w22668_,
		_w22669_
	);
	LUT3 #(
		.INIT('h2a)
	) name12157 (
		_w18752_,
		_w22645_,
		_w22669_,
		_w22670_
	);
	LUT3 #(
		.INIT('h15)
	) name12158 (
		wb_rst_i_pad,
		_w22645_,
		_w22669_,
		_w22671_
	);
	LUT3 #(
		.INIT('hdc)
	) name12159 (
		_w14151_,
		_w22670_,
		_w22671_,
		_w22672_
	);
	LUT4 #(
		.INIT('h050d)
	) name12160 (
		\wishbone_TxLength_reg[7]/NET0131 ,
		_w12311_,
		_w13399_,
		_w14878_,
		_w22673_
	);
	LUT2 #(
		.INIT('h2)
	) name12161 (
		_w15777_,
		_w22673_,
		_w22674_
	);
	LUT3 #(
		.INIT('hf2)
	) name12162 (
		_w12303_,
		_w18401_,
		_w22674_,
		_w22675_
	);
	LUT3 #(
		.INIT('h70)
	) name12163 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_TxLength_reg[5]/NET0131 ,
		_w22676_
	);
	LUT2 #(
		.INIT('h4)
	) name12164 (
		_w12302_,
		_w22676_,
		_w22677_
	);
	LUT4 #(
		.INIT('h01fe)
	) name12165 (
		\wishbone_TxLength_reg[2]/NET0131 ,
		\wishbone_TxLength_reg[3]/NET0131 ,
		\wishbone_TxLength_reg[4]/NET0131 ,
		\wishbone_TxLength_reg[5]/NET0131 ,
		_w22678_
	);
	LUT4 #(
		.INIT('h0800)
	) name12166 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		\wishbone_TxLength_reg[5]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		_w22679_
	);
	LUT3 #(
		.INIT('h01)
	) name12167 (
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w22678_,
		_w22679_,
		_w22680_
	);
	LUT3 #(
		.INIT('h08)
	) name12168 (
		\wishbone_TxLength_reg[5]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w22681_
	);
	LUT2 #(
		.INIT('h8)
	) name12169 (
		_w14516_,
		_w22681_,
		_w22682_
	);
	LUT2 #(
		.INIT('h1)
	) name12170 (
		_w22680_,
		_w22682_,
		_w22683_
	);
	LUT3 #(
		.INIT('h80)
	) name12171 (
		_w14519_,
		_w14520_,
		_w19165_,
		_w22684_
	);
	LUT3 #(
		.INIT('h80)
	) name12172 (
		\wishbone_TxLength_reg[5]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w22685_
	);
	LUT3 #(
		.INIT('h70)
	) name12173 (
		_w12309_,
		_w14520_,
		_w22685_,
		_w22686_
	);
	LUT3 #(
		.INIT('hb7)
	) name12174 (
		\wishbone_TxLength_reg[5]/NET0131 ,
		_w14526_,
		_w14527_,
		_w22687_
	);
	LUT3 #(
		.INIT('h10)
	) name12175 (
		_w22684_,
		_w22686_,
		_w22687_,
		_w22688_
	);
	LUT4 #(
		.INIT('h0444)
	) name12176 (
		_w12302_,
		_w12304_,
		_w12312_,
		_w12317_,
		_w22689_
	);
	LUT4 #(
		.INIT('h4055)
	) name12177 (
		_w22677_,
		_w22683_,
		_w22688_,
		_w22689_,
		_w22690_
	);
	LUT3 #(
		.INIT('h2f)
	) name12178 (
		_w12303_,
		_w18058_,
		_w22690_,
		_w22691_
	);
	LUT4 #(
		.INIT('h0020)
	) name12179 (
		\ethreg1_TXCTRL_2_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22692_
	);
	LUT3 #(
		.INIT('h80)
	) name12180 (
		_w18757_,
		_w18758_,
		_w22692_,
		_w22693_
	);
	LUT3 #(
		.INIT('h80)
	) name12181 (
		\ethreg1_MODER_2_DataOut_reg[0]/NET0131 ,
		_w18800_,
		_w18801_,
		_w22694_
	);
	LUT4 #(
		.INIT('h0008)
	) name12182 (
		\ethreg1_RXHASH0_2_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22695_
	);
	LUT3 #(
		.INIT('h80)
	) name12183 (
		_w18757_,
		_w18758_,
		_w22695_,
		_w22696_
	);
	LUT3 #(
		.INIT('h01)
	) name12184 (
		_w22693_,
		_w22694_,
		_w22696_,
		_w22697_
	);
	LUT4 #(
		.INIT('h0008)
	) name12185 (
		\ethreg1_RXHASH1_2_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22698_
	);
	LUT3 #(
		.INIT('h80)
	) name12186 (
		_w18757_,
		_w18762_,
		_w22698_,
		_w22699_
	);
	LUT4 #(
		.INIT('h0002)
	) name12187 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22700_
	);
	LUT3 #(
		.INIT('h80)
	) name12188 (
		_w18757_,
		_w18758_,
		_w22700_,
		_w22701_
	);
	LUT3 #(
		.INIT('h80)
	) name12189 (
		\ethreg1_COLLCONF_2_DataOut_reg[0]/NET0131 ,
		_w18753_,
		_w19641_,
		_w22702_
	);
	LUT3 #(
		.INIT('h80)
	) name12190 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		_w18753_,
		_w18754_,
		_w22703_
	);
	LUT4 #(
		.INIT('h0001)
	) name12191 (
		_w22699_,
		_w22701_,
		_w22702_,
		_w22703_,
		_w22704_
	);
	LUT3 #(
		.INIT('h2a)
	) name12192 (
		_w18752_,
		_w22697_,
		_w22704_,
		_w22705_
	);
	LUT4 #(
		.INIT('h5455)
	) name12193 (
		wb_rst_i_pad,
		wb_we_i_pad,
		_w18750_,
		_w18751_,
		_w22706_
	);
	LUT3 #(
		.INIT('hdc)
	) name12194 (
		_w16122_,
		_w22705_,
		_w22706_,
		_w22707_
	);
	LUT3 #(
		.INIT('h80)
	) name12195 (
		\ethreg1_IPGT_0_DataOut_reg[6]/NET0131 ,
		_w19646_,
		_w19655_,
		_w22708_
	);
	LUT4 #(
		.INIT('h0008)
	) name12196 (
		\ethreg1_RXHASH1_0_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22709_
	);
	LUT3 #(
		.INIT('h80)
	) name12197 (
		_w18757_,
		_w18762_,
		_w22709_,
		_w22710_
	);
	LUT3 #(
		.INIT('h80)
	) name12198 (
		\ethreg1_IPGR2_0_DataOut_reg[6]/NET0131 ,
		_w18800_,
		_w18805_,
		_w22711_
	);
	LUT3 #(
		.INIT('h80)
	) name12199 (
		\ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131 ,
		_w18786_,
		_w18801_,
		_w22712_
	);
	LUT4 #(
		.INIT('h0001)
	) name12200 (
		_w22708_,
		_w22710_,
		_w22711_,
		_w22712_,
		_w22713_
	);
	LUT2 #(
		.INIT('h8)
	) name12201 (
		_w18752_,
		_w22713_,
		_w22714_
	);
	LUT3 #(
		.INIT('h80)
	) name12202 (
		\ethreg1_IPGR1_0_DataOut_reg[6]/NET0131 ,
		_w18785_,
		_w18800_,
		_w22715_
	);
	LUT3 #(
		.INIT('h80)
	) name12203 (
		\ethreg1_MODER_0_DataOut_reg[6]/NET0131 ,
		_w18800_,
		_w18801_,
		_w22716_
	);
	LUT3 #(
		.INIT('h80)
	) name12204 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[6]/NET0131 ,
		_w18798_,
		_w18801_,
		_w22717_
	);
	LUT4 #(
		.INIT('h0002)
	) name12205 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22718_
	);
	LUT3 #(
		.INIT('h80)
	) name12206 (
		_w18757_,
		_w18762_,
		_w22718_,
		_w22719_
	);
	LUT4 #(
		.INIT('h0001)
	) name12207 (
		_w22715_,
		_w22716_,
		_w22717_,
		_w22719_,
		_w22720_
	);
	LUT4 #(
		.INIT('h0008)
	) name12208 (
		\ethreg1_RXHASH0_0_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22721_
	);
	LUT3 #(
		.INIT('h80)
	) name12209 (
		_w18757_,
		_w18758_,
		_w22721_,
		_w22722_
	);
	LUT3 #(
		.INIT('h80)
	) name12210 (
		\ethreg1_INT_MASK_0_DataOut_reg[6]/NET0131 ,
		_w18801_,
		_w19655_,
		_w22723_
	);
	LUT4 #(
		.INIT('h0002)
	) name12211 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22724_
	);
	LUT4 #(
		.INIT('h0020)
	) name12212 (
		\ethreg1_TXCTRL_0_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22725_
	);
	LUT4 #(
		.INIT('h777f)
	) name12213 (
		_w18757_,
		_w18758_,
		_w22724_,
		_w22725_,
		_w22726_
	);
	LUT3 #(
		.INIT('h10)
	) name12214 (
		_w22722_,
		_w22723_,
		_w22726_,
		_w22727_
	);
	LUT3 #(
		.INIT('h80)
	) name12215 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[6]/NET0131 ,
		_w18798_,
		_w18805_,
		_w22728_
	);
	LUT3 #(
		.INIT('h80)
	) name12216 (
		\ethreg1_irq_rxc_reg/NET0131 ,
		_w18800_,
		_w19646_,
		_w22729_
	);
	LUT3 #(
		.INIT('h80)
	) name12217 (
		\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 ,
		_w18753_,
		_w18754_,
		_w22730_
	);
	LUT3 #(
		.INIT('h80)
	) name12218 (
		\ethreg1_MIIRX_DATA_DataOut_reg[6]/NET0131 ,
		_w18785_,
		_w18786_,
		_w22731_
	);
	LUT4 #(
		.INIT('h0001)
	) name12219 (
		_w22728_,
		_w22729_,
		_w22730_,
		_w22731_,
		_w22732_
	);
	LUT3 #(
		.INIT('h80)
	) name12220 (
		_w22720_,
		_w22727_,
		_w22732_,
		_w22733_
	);
	LUT3 #(
		.INIT('h2a)
	) name12221 (
		_w18752_,
		_w22713_,
		_w22733_,
		_w22734_
	);
	LUT3 #(
		.INIT('h80)
	) name12222 (
		\wishbone_bd_ram_mem0_reg[80][6]/P0001 ,
		_w11941_,
		_w11972_,
		_w22735_
	);
	LUT3 #(
		.INIT('h80)
	) name12223 (
		\wishbone_bd_ram_mem0_reg[33][6]/P0001 ,
		_w11957_,
		_w11977_,
		_w22736_
	);
	LUT3 #(
		.INIT('h80)
	) name12224 (
		\wishbone_bd_ram_mem0_reg[21][6]/P0001 ,
		_w11933_,
		_w11935_,
		_w22737_
	);
	LUT3 #(
		.INIT('h80)
	) name12225 (
		\wishbone_bd_ram_mem0_reg[73][6]/P0001 ,
		_w11949_,
		_w11968_,
		_w22738_
	);
	LUT4 #(
		.INIT('h0001)
	) name12226 (
		_w22735_,
		_w22736_,
		_w22737_,
		_w22738_,
		_w22739_
	);
	LUT3 #(
		.INIT('h80)
	) name12227 (
		\wishbone_bd_ram_mem0_reg[210][6]/P0001 ,
		_w11963_,
		_w11984_,
		_w22740_
	);
	LUT3 #(
		.INIT('h80)
	) name12228 (
		\wishbone_bd_ram_mem0_reg[121][6]/P0001 ,
		_w11968_,
		_w12012_,
		_w22741_
	);
	LUT3 #(
		.INIT('h80)
	) name12229 (
		\wishbone_bd_ram_mem0_reg[149][6]/P0001 ,
		_w11933_,
		_w11959_,
		_w22742_
	);
	LUT3 #(
		.INIT('h80)
	) name12230 (
		\wishbone_bd_ram_mem0_reg[183][6]/P0001 ,
		_w11942_,
		_w11975_,
		_w22743_
	);
	LUT4 #(
		.INIT('h0001)
	) name12231 (
		_w22740_,
		_w22741_,
		_w22742_,
		_w22743_,
		_w22744_
	);
	LUT3 #(
		.INIT('h80)
	) name12232 (
		\wishbone_bd_ram_mem0_reg[249][6]/P0001 ,
		_w11952_,
		_w11968_,
		_w22745_
	);
	LUT3 #(
		.INIT('h80)
	) name12233 (
		\wishbone_bd_ram_mem0_reg[255][6]/P0001 ,
		_w11952_,
		_w11973_,
		_w22746_
	);
	LUT3 #(
		.INIT('h80)
	) name12234 (
		\wishbone_bd_ram_mem0_reg[84][6]/P0001 ,
		_w11929_,
		_w11972_,
		_w22747_
	);
	LUT3 #(
		.INIT('h80)
	) name12235 (
		\wishbone_bd_ram_mem0_reg[237][6]/P0001 ,
		_w11966_,
		_w11982_,
		_w22748_
	);
	LUT4 #(
		.INIT('h0001)
	) name12236 (
		_w22745_,
		_w22746_,
		_w22747_,
		_w22748_,
		_w22749_
	);
	LUT3 #(
		.INIT('h80)
	) name12237 (
		\wishbone_bd_ram_mem0_reg[51][6]/P0001 ,
		_w11938_,
		_w11979_,
		_w22750_
	);
	LUT3 #(
		.INIT('h80)
	) name12238 (
		\wishbone_bd_ram_mem0_reg[252][6]/P0001 ,
		_w11952_,
		_w11954_,
		_w22751_
	);
	LUT3 #(
		.INIT('h80)
	) name12239 (
		\wishbone_bd_ram_mem0_reg[32][6]/P0001 ,
		_w11941_,
		_w11957_,
		_w22752_
	);
	LUT3 #(
		.INIT('h80)
	) name12240 (
		\wishbone_bd_ram_mem0_reg[144][6]/P0001 ,
		_w11941_,
		_w11959_,
		_w22753_
	);
	LUT4 #(
		.INIT('h0001)
	) name12241 (
		_w22750_,
		_w22751_,
		_w22752_,
		_w22753_,
		_w22754_
	);
	LUT4 #(
		.INIT('h8000)
	) name12242 (
		_w22739_,
		_w22744_,
		_w22749_,
		_w22754_,
		_w22755_
	);
	LUT3 #(
		.INIT('h80)
	) name12243 (
		\wishbone_bd_ram_mem0_reg[89][6]/P0001 ,
		_w11968_,
		_w11972_,
		_w22756_
	);
	LUT3 #(
		.INIT('h80)
	) name12244 (
		\wishbone_bd_ram_mem0_reg[104][6]/P0001 ,
		_w11965_,
		_w11990_,
		_w22757_
	);
	LUT3 #(
		.INIT('h80)
	) name12245 (
		\wishbone_bd_ram_mem0_reg[194][6]/P0001 ,
		_w11945_,
		_w11963_,
		_w22758_
	);
	LUT3 #(
		.INIT('h80)
	) name12246 (
		\wishbone_bd_ram_mem0_reg[92][6]/P0001 ,
		_w11954_,
		_w11972_,
		_w22759_
	);
	LUT4 #(
		.INIT('h0001)
	) name12247 (
		_w22756_,
		_w22757_,
		_w22758_,
		_w22759_,
		_w22760_
	);
	LUT3 #(
		.INIT('h80)
	) name12248 (
		\wishbone_bd_ram_mem0_reg[221][6]/P0001 ,
		_w11966_,
		_w11984_,
		_w22761_
	);
	LUT3 #(
		.INIT('h80)
	) name12249 (
		\wishbone_bd_ram_mem0_reg[127][6]/P0001 ,
		_w11973_,
		_w12012_,
		_w22762_
	);
	LUT3 #(
		.INIT('h80)
	) name12250 (
		\wishbone_bd_ram_mem0_reg[74][6]/P0001 ,
		_w11944_,
		_w11949_,
		_w22763_
	);
	LUT3 #(
		.INIT('h80)
	) name12251 (
		\wishbone_bd_ram_mem0_reg[4][6]/P0001 ,
		_w11929_,
		_w11932_,
		_w22764_
	);
	LUT4 #(
		.INIT('h0001)
	) name12252 (
		_w22761_,
		_w22762_,
		_w22763_,
		_w22764_,
		_w22765_
	);
	LUT3 #(
		.INIT('h80)
	) name12253 (
		\wishbone_bd_ram_mem0_reg[174][6]/P0001 ,
		_w11930_,
		_w11948_,
		_w22766_
	);
	LUT3 #(
		.INIT('h80)
	) name12254 (
		\wishbone_bd_ram_mem0_reg[178][6]/P0001 ,
		_w11942_,
		_w11963_,
		_w22767_
	);
	LUT3 #(
		.INIT('h80)
	) name12255 (
		\wishbone_bd_ram_mem0_reg[217][6]/P0001 ,
		_w11968_,
		_w11984_,
		_w22768_
	);
	LUT3 #(
		.INIT('h80)
	) name12256 (
		\wishbone_bd_ram_mem0_reg[72][6]/P0001 ,
		_w11949_,
		_w11990_,
		_w22769_
	);
	LUT4 #(
		.INIT('h0001)
	) name12257 (
		_w22766_,
		_w22767_,
		_w22768_,
		_w22769_,
		_w22770_
	);
	LUT3 #(
		.INIT('h80)
	) name12258 (
		\wishbone_bd_ram_mem0_reg[79][6]/P0001 ,
		_w11949_,
		_w11973_,
		_w22771_
	);
	LUT3 #(
		.INIT('h80)
	) name12259 (
		\wishbone_bd_ram_mem0_reg[212][6]/P0001 ,
		_w11929_,
		_w11984_,
		_w22772_
	);
	LUT3 #(
		.INIT('h80)
	) name12260 (
		\wishbone_bd_ram_mem0_reg[151][6]/P0001 ,
		_w11959_,
		_w11975_,
		_w22773_
	);
	LUT3 #(
		.INIT('h80)
	) name12261 (
		\wishbone_bd_ram_mem0_reg[225][6]/P0001 ,
		_w11977_,
		_w11982_,
		_w22774_
	);
	LUT4 #(
		.INIT('h0001)
	) name12262 (
		_w22771_,
		_w22772_,
		_w22773_,
		_w22774_,
		_w22775_
	);
	LUT4 #(
		.INIT('h8000)
	) name12263 (
		_w22760_,
		_w22765_,
		_w22770_,
		_w22775_,
		_w22776_
	);
	LUT3 #(
		.INIT('h80)
	) name12264 (
		\wishbone_bd_ram_mem0_reg[197][6]/P0001 ,
		_w11933_,
		_w11945_,
		_w22777_
	);
	LUT3 #(
		.INIT('h80)
	) name12265 (
		\wishbone_bd_ram_mem0_reg[208][6]/P0001 ,
		_w11941_,
		_w11984_,
		_w22778_
	);
	LUT3 #(
		.INIT('h80)
	) name12266 (
		\wishbone_bd_ram_mem0_reg[176][6]/P0001 ,
		_w11941_,
		_w11942_,
		_w22779_
	);
	LUT3 #(
		.INIT('h80)
	) name12267 (
		\wishbone_bd_ram_mem0_reg[65][6]/P0001 ,
		_w11949_,
		_w11977_,
		_w22780_
	);
	LUT4 #(
		.INIT('h0001)
	) name12268 (
		_w22777_,
		_w22778_,
		_w22779_,
		_w22780_,
		_w22781_
	);
	LUT3 #(
		.INIT('h80)
	) name12269 (
		\wishbone_bd_ram_mem0_reg[3][6]/P0001 ,
		_w11932_,
		_w11938_,
		_w22782_
	);
	LUT3 #(
		.INIT('h80)
	) name12270 (
		\wishbone_bd_ram_mem0_reg[85][6]/P0001 ,
		_w11933_,
		_w11972_,
		_w22783_
	);
	LUT3 #(
		.INIT('h80)
	) name12271 (
		\wishbone_bd_ram_mem0_reg[9][6]/P0001 ,
		_w11932_,
		_w11968_,
		_w22784_
	);
	LUT3 #(
		.INIT('h80)
	) name12272 (
		\wishbone_bd_ram_mem0_reg[145][6]/P0001 ,
		_w11959_,
		_w11977_,
		_w22785_
	);
	LUT4 #(
		.INIT('h0001)
	) name12273 (
		_w22782_,
		_w22783_,
		_w22784_,
		_w22785_,
		_w22786_
	);
	LUT3 #(
		.INIT('h80)
	) name12274 (
		\wishbone_bd_ram_mem0_reg[64][6]/P0001 ,
		_w11941_,
		_w11949_,
		_w22787_
	);
	LUT3 #(
		.INIT('h80)
	) name12275 (
		\wishbone_bd_ram_mem0_reg[147][6]/P0001 ,
		_w11938_,
		_w11959_,
		_w22788_
	);
	LUT3 #(
		.INIT('h80)
	) name12276 (
		\wishbone_bd_ram_mem0_reg[218][6]/P0001 ,
		_w11944_,
		_w11984_,
		_w22789_
	);
	LUT3 #(
		.INIT('h80)
	) name12277 (
		\wishbone_bd_ram_mem0_reg[188][6]/P0001 ,
		_w11942_,
		_w11954_,
		_w22790_
	);
	LUT4 #(
		.INIT('h0001)
	) name12278 (
		_w22787_,
		_w22788_,
		_w22789_,
		_w22790_,
		_w22791_
	);
	LUT3 #(
		.INIT('h80)
	) name12279 (
		\wishbone_bd_ram_mem0_reg[139][6]/P0001 ,
		_w11936_,
		_w11955_,
		_w22792_
	);
	LUT3 #(
		.INIT('h80)
	) name12280 (
		\wishbone_bd_ram_mem0_reg[207][6]/P0001 ,
		_w11945_,
		_w11973_,
		_w22793_
	);
	LUT3 #(
		.INIT('h80)
	) name12281 (
		\wishbone_bd_ram_mem0_reg[128][6]/P0001 ,
		_w11941_,
		_w11955_,
		_w22794_
	);
	LUT3 #(
		.INIT('h80)
	) name12282 (
		\wishbone_bd_ram_mem0_reg[216][6]/P0001 ,
		_w11984_,
		_w11990_,
		_w22795_
	);
	LUT4 #(
		.INIT('h0001)
	) name12283 (
		_w22792_,
		_w22793_,
		_w22794_,
		_w22795_,
		_w22796_
	);
	LUT4 #(
		.INIT('h8000)
	) name12284 (
		_w22781_,
		_w22786_,
		_w22791_,
		_w22796_,
		_w22797_
	);
	LUT3 #(
		.INIT('h80)
	) name12285 (
		\wishbone_bd_ram_mem0_reg[138][6]/P0001 ,
		_w11944_,
		_w11955_,
		_w22798_
	);
	LUT3 #(
		.INIT('h80)
	) name12286 (
		\wishbone_bd_ram_mem0_reg[177][6]/P0001 ,
		_w11942_,
		_w11977_,
		_w22799_
	);
	LUT3 #(
		.INIT('h80)
	) name12287 (
		\wishbone_bd_ram_mem0_reg[171][6]/P0001 ,
		_w11930_,
		_w11936_,
		_w22800_
	);
	LUT3 #(
		.INIT('h80)
	) name12288 (
		\wishbone_bd_ram_mem0_reg[182][6]/P0001 ,
		_w11942_,
		_w11986_,
		_w22801_
	);
	LUT4 #(
		.INIT('h0001)
	) name12289 (
		_w22798_,
		_w22799_,
		_w22800_,
		_w22801_,
		_w22802_
	);
	LUT3 #(
		.INIT('h80)
	) name12290 (
		\wishbone_bd_ram_mem0_reg[181][6]/P0001 ,
		_w11933_,
		_w11942_,
		_w22803_
	);
	LUT3 #(
		.INIT('h80)
	) name12291 (
		\wishbone_bd_ram_mem0_reg[113][6]/P0001 ,
		_w11977_,
		_w12012_,
		_w22804_
	);
	LUT3 #(
		.INIT('h80)
	) name12292 (
		\wishbone_bd_ram_mem0_reg[49][6]/P0001 ,
		_w11977_,
		_w11979_,
		_w22805_
	);
	LUT3 #(
		.INIT('h80)
	) name12293 (
		\wishbone_bd_ram_mem0_reg[13][6]/P0001 ,
		_w11932_,
		_w11966_,
		_w22806_
	);
	LUT4 #(
		.INIT('h0001)
	) name12294 (
		_w22803_,
		_w22804_,
		_w22805_,
		_w22806_,
		_w22807_
	);
	LUT3 #(
		.INIT('h80)
	) name12295 (
		\wishbone_bd_ram_mem0_reg[154][6]/P0001 ,
		_w11944_,
		_w11959_,
		_w22808_
	);
	LUT3 #(
		.INIT('h80)
	) name12296 (
		\wishbone_bd_ram_mem0_reg[118][6]/P0001 ,
		_w11986_,
		_w12012_,
		_w22809_
	);
	LUT3 #(
		.INIT('h80)
	) name12297 (
		\wishbone_bd_ram_mem0_reg[137][6]/P0001 ,
		_w11955_,
		_w11968_,
		_w22810_
	);
	LUT3 #(
		.INIT('h80)
	) name12298 (
		\wishbone_bd_ram_mem0_reg[20][6]/P0001 ,
		_w11929_,
		_w11935_,
		_w22811_
	);
	LUT4 #(
		.INIT('h0001)
	) name12299 (
		_w22808_,
		_w22809_,
		_w22810_,
		_w22811_,
		_w22812_
	);
	LUT3 #(
		.INIT('h80)
	) name12300 (
		\wishbone_bd_ram_mem0_reg[76][6]/P0001 ,
		_w11949_,
		_w11954_,
		_w22813_
	);
	LUT3 #(
		.INIT('h80)
	) name12301 (
		\wishbone_bd_ram_mem0_reg[109][6]/P0001 ,
		_w11965_,
		_w11966_,
		_w22814_
	);
	LUT3 #(
		.INIT('h80)
	) name12302 (
		\wishbone_bd_ram_mem0_reg[2][6]/P0001 ,
		_w11932_,
		_w11963_,
		_w22815_
	);
	LUT3 #(
		.INIT('h80)
	) name12303 (
		\wishbone_bd_ram_mem0_reg[186][6]/P0001 ,
		_w11942_,
		_w11944_,
		_w22816_
	);
	LUT4 #(
		.INIT('h0001)
	) name12304 (
		_w22813_,
		_w22814_,
		_w22815_,
		_w22816_,
		_w22817_
	);
	LUT4 #(
		.INIT('h8000)
	) name12305 (
		_w22802_,
		_w22807_,
		_w22812_,
		_w22817_,
		_w22818_
	);
	LUT4 #(
		.INIT('h8000)
	) name12306 (
		_w22755_,
		_w22776_,
		_w22797_,
		_w22818_,
		_w22819_
	);
	LUT3 #(
		.INIT('h80)
	) name12307 (
		\wishbone_bd_ram_mem0_reg[61][6]/P0001 ,
		_w11966_,
		_w11979_,
		_w22820_
	);
	LUT3 #(
		.INIT('h80)
	) name12308 (
		\wishbone_bd_ram_mem0_reg[162][6]/P0001 ,
		_w11930_,
		_w11963_,
		_w22821_
	);
	LUT3 #(
		.INIT('h80)
	) name12309 (
		\wishbone_bd_ram_mem0_reg[203][6]/P0001 ,
		_w11936_,
		_w11945_,
		_w22822_
	);
	LUT3 #(
		.INIT('h80)
	) name12310 (
		\wishbone_bd_ram_mem0_reg[231][6]/P0001 ,
		_w11975_,
		_w11982_,
		_w22823_
	);
	LUT4 #(
		.INIT('h0001)
	) name12311 (
		_w22820_,
		_w22821_,
		_w22822_,
		_w22823_,
		_w22824_
	);
	LUT3 #(
		.INIT('h80)
	) name12312 (
		\wishbone_bd_ram_mem0_reg[223][6]/P0001 ,
		_w11973_,
		_w11984_,
		_w22825_
	);
	LUT3 #(
		.INIT('h80)
	) name12313 (
		\wishbone_bd_ram_mem0_reg[196][6]/P0001 ,
		_w11929_,
		_w11945_,
		_w22826_
	);
	LUT3 #(
		.INIT('h80)
	) name12314 (
		\wishbone_bd_ram_mem0_reg[62][6]/P0001 ,
		_w11948_,
		_w11979_,
		_w22827_
	);
	LUT3 #(
		.INIT('h80)
	) name12315 (
		\wishbone_bd_ram_mem0_reg[52][6]/P0001 ,
		_w11929_,
		_w11979_,
		_w22828_
	);
	LUT4 #(
		.INIT('h0001)
	) name12316 (
		_w22825_,
		_w22826_,
		_w22827_,
		_w22828_,
		_w22829_
	);
	LUT3 #(
		.INIT('h80)
	) name12317 (
		\wishbone_bd_ram_mem0_reg[193][6]/P0001 ,
		_w11945_,
		_w11977_,
		_w22830_
	);
	LUT3 #(
		.INIT('h80)
	) name12318 (
		\wishbone_bd_ram_mem0_reg[59][6]/P0001 ,
		_w11936_,
		_w11979_,
		_w22831_
	);
	LUT3 #(
		.INIT('h80)
	) name12319 (
		\wishbone_bd_ram_mem0_reg[71][6]/P0001 ,
		_w11949_,
		_w11975_,
		_w22832_
	);
	LUT3 #(
		.INIT('h80)
	) name12320 (
		\wishbone_bd_ram_mem0_reg[191][6]/P0001 ,
		_w11942_,
		_w11973_,
		_w22833_
	);
	LUT4 #(
		.INIT('h0001)
	) name12321 (
		_w22830_,
		_w22831_,
		_w22832_,
		_w22833_,
		_w22834_
	);
	LUT3 #(
		.INIT('h80)
	) name12322 (
		\wishbone_bd_ram_mem0_reg[198][6]/P0001 ,
		_w11945_,
		_w11986_,
		_w22835_
	);
	LUT3 #(
		.INIT('h80)
	) name12323 (
		\wishbone_bd_ram_mem0_reg[98][6]/P0001 ,
		_w11963_,
		_w11965_,
		_w22836_
	);
	LUT3 #(
		.INIT('h80)
	) name12324 (
		\wishbone_bd_ram_mem0_reg[120][6]/P0001 ,
		_w11990_,
		_w12012_,
		_w22837_
	);
	LUT3 #(
		.INIT('h80)
	) name12325 (
		\wishbone_bd_ram_mem0_reg[63][6]/P0001 ,
		_w11973_,
		_w11979_,
		_w22838_
	);
	LUT4 #(
		.INIT('h0001)
	) name12326 (
		_w22835_,
		_w22836_,
		_w22837_,
		_w22838_,
		_w22839_
	);
	LUT4 #(
		.INIT('h8000)
	) name12327 (
		_w22824_,
		_w22829_,
		_w22834_,
		_w22839_,
		_w22840_
	);
	LUT3 #(
		.INIT('h80)
	) name12328 (
		\wishbone_bd_ram_mem0_reg[161][6]/P0001 ,
		_w11930_,
		_w11977_,
		_w22841_
	);
	LUT3 #(
		.INIT('h80)
	) name12329 (
		\wishbone_bd_ram_mem0_reg[243][6]/P0001 ,
		_w11938_,
		_w11952_,
		_w22842_
	);
	LUT3 #(
		.INIT('h80)
	) name12330 (
		\wishbone_bd_ram_mem0_reg[38][6]/P0001 ,
		_w11957_,
		_w11986_,
		_w22843_
	);
	LUT3 #(
		.INIT('h80)
	) name12331 (
		\wishbone_bd_ram_mem0_reg[22][6]/P0001 ,
		_w11935_,
		_w11986_,
		_w22844_
	);
	LUT4 #(
		.INIT('h0001)
	) name12332 (
		_w22841_,
		_w22842_,
		_w22843_,
		_w22844_,
		_w22845_
	);
	LUT3 #(
		.INIT('h80)
	) name12333 (
		\wishbone_bd_ram_mem0_reg[58][6]/P0001 ,
		_w11944_,
		_w11979_,
		_w22846_
	);
	LUT3 #(
		.INIT('h80)
	) name12334 (
		\wishbone_bd_ram_mem0_reg[56][6]/P0001 ,
		_w11979_,
		_w11990_,
		_w22847_
	);
	LUT3 #(
		.INIT('h80)
	) name12335 (
		\wishbone_bd_ram_mem0_reg[126][6]/P0001 ,
		_w11948_,
		_w12012_,
		_w22848_
	);
	LUT3 #(
		.INIT('h80)
	) name12336 (
		\wishbone_bd_ram_mem0_reg[125][6]/P0001 ,
		_w11966_,
		_w12012_,
		_w22849_
	);
	LUT4 #(
		.INIT('h0001)
	) name12337 (
		_w22846_,
		_w22847_,
		_w22848_,
		_w22849_,
		_w22850_
	);
	LUT3 #(
		.INIT('h80)
	) name12338 (
		\wishbone_bd_ram_mem0_reg[44][6]/P0001 ,
		_w11954_,
		_w11957_,
		_w22851_
	);
	LUT3 #(
		.INIT('h80)
	) name12339 (
		\wishbone_bd_ram_mem0_reg[94][6]/P0001 ,
		_w11948_,
		_w11972_,
		_w22852_
	);
	LUT3 #(
		.INIT('h80)
	) name12340 (
		\wishbone_bd_ram_mem0_reg[29][6]/P0001 ,
		_w11935_,
		_w11966_,
		_w22853_
	);
	LUT3 #(
		.INIT('h80)
	) name12341 (
		\wishbone_bd_ram_mem0_reg[66][6]/P0001 ,
		_w11949_,
		_w11963_,
		_w22854_
	);
	LUT4 #(
		.INIT('h0001)
	) name12342 (
		_w22851_,
		_w22852_,
		_w22853_,
		_w22854_,
		_w22855_
	);
	LUT3 #(
		.INIT('h80)
	) name12343 (
		\wishbone_bd_ram_mem0_reg[130][6]/P0001 ,
		_w11955_,
		_w11963_,
		_w22856_
	);
	LUT3 #(
		.INIT('h80)
	) name12344 (
		\wishbone_bd_ram_mem0_reg[18][6]/P0001 ,
		_w11935_,
		_w11963_,
		_w22857_
	);
	LUT3 #(
		.INIT('h80)
	) name12345 (
		\wishbone_bd_ram_mem0_reg[199][6]/P0001 ,
		_w11945_,
		_w11975_,
		_w22858_
	);
	LUT3 #(
		.INIT('h80)
	) name12346 (
		\wishbone_bd_ram_mem0_reg[45][6]/P0001 ,
		_w11957_,
		_w11966_,
		_w22859_
	);
	LUT4 #(
		.INIT('h0001)
	) name12347 (
		_w22856_,
		_w22857_,
		_w22858_,
		_w22859_,
		_w22860_
	);
	LUT4 #(
		.INIT('h8000)
	) name12348 (
		_w22845_,
		_w22850_,
		_w22855_,
		_w22860_,
		_w22861_
	);
	LUT3 #(
		.INIT('h80)
	) name12349 (
		\wishbone_bd_ram_mem0_reg[19][6]/P0001 ,
		_w11935_,
		_w11938_,
		_w22862_
	);
	LUT3 #(
		.INIT('h80)
	) name12350 (
		\wishbone_bd_ram_mem0_reg[133][6]/P0001 ,
		_w11933_,
		_w11955_,
		_w22863_
	);
	LUT3 #(
		.INIT('h80)
	) name12351 (
		\wishbone_bd_ram_mem0_reg[96][6]/P0001 ,
		_w11941_,
		_w11965_,
		_w22864_
	);
	LUT3 #(
		.INIT('h80)
	) name12352 (
		\wishbone_bd_ram_mem0_reg[224][6]/P0001 ,
		_w11941_,
		_w11982_,
		_w22865_
	);
	LUT4 #(
		.INIT('h0001)
	) name12353 (
		_w22862_,
		_w22863_,
		_w22864_,
		_w22865_,
		_w22866_
	);
	LUT3 #(
		.INIT('h80)
	) name12354 (
		\wishbone_bd_ram_mem0_reg[114][6]/P0001 ,
		_w11963_,
		_w12012_,
		_w22867_
	);
	LUT3 #(
		.INIT('h80)
	) name12355 (
		\wishbone_bd_ram_mem0_reg[227][6]/P0001 ,
		_w11938_,
		_w11982_,
		_w22868_
	);
	LUT3 #(
		.INIT('h80)
	) name12356 (
		\wishbone_bd_ram_mem0_reg[1][6]/P0001 ,
		_w11932_,
		_w11977_,
		_w22869_
	);
	LUT3 #(
		.INIT('h80)
	) name12357 (
		\wishbone_bd_ram_mem0_reg[60][6]/P0001 ,
		_w11954_,
		_w11979_,
		_w22870_
	);
	LUT4 #(
		.INIT('h0001)
	) name12358 (
		_w22867_,
		_w22868_,
		_w22869_,
		_w22870_,
		_w22871_
	);
	LUT3 #(
		.INIT('h80)
	) name12359 (
		\wishbone_bd_ram_mem0_reg[219][6]/P0001 ,
		_w11936_,
		_w11984_,
		_w22872_
	);
	LUT3 #(
		.INIT('h80)
	) name12360 (
		\wishbone_bd_ram_mem0_reg[179][6]/P0001 ,
		_w11938_,
		_w11942_,
		_w22873_
	);
	LUT3 #(
		.INIT('h80)
	) name12361 (
		\wishbone_bd_ram_mem0_reg[146][6]/P0001 ,
		_w11959_,
		_w11963_,
		_w22874_
	);
	LUT3 #(
		.INIT('h80)
	) name12362 (
		\wishbone_bd_ram_mem0_reg[204][6]/P0001 ,
		_w11945_,
		_w11954_,
		_w22875_
	);
	LUT4 #(
		.INIT('h0001)
	) name12363 (
		_w22872_,
		_w22873_,
		_w22874_,
		_w22875_,
		_w22876_
	);
	LUT3 #(
		.INIT('h80)
	) name12364 (
		\wishbone_bd_ram_mem0_reg[88][6]/P0001 ,
		_w11972_,
		_w11990_,
		_w22877_
	);
	LUT3 #(
		.INIT('h80)
	) name12365 (
		\wishbone_bd_ram_mem0_reg[254][6]/P0001 ,
		_w11948_,
		_w11952_,
		_w22878_
	);
	LUT3 #(
		.INIT('h80)
	) name12366 (
		\wishbone_bd_ram_mem0_reg[87][6]/P0001 ,
		_w11972_,
		_w11975_,
		_w22879_
	);
	LUT3 #(
		.INIT('h80)
	) name12367 (
		\wishbone_bd_ram_mem0_reg[100][6]/P0001 ,
		_w11929_,
		_w11965_,
		_w22880_
	);
	LUT4 #(
		.INIT('h0001)
	) name12368 (
		_w22877_,
		_w22878_,
		_w22879_,
		_w22880_,
		_w22881_
	);
	LUT4 #(
		.INIT('h8000)
	) name12369 (
		_w22866_,
		_w22871_,
		_w22876_,
		_w22881_,
		_w22882_
	);
	LUT3 #(
		.INIT('h80)
	) name12370 (
		\wishbone_bd_ram_mem0_reg[26][6]/P0001 ,
		_w11935_,
		_w11944_,
		_w22883_
	);
	LUT3 #(
		.INIT('h80)
	) name12371 (
		\wishbone_bd_ram_mem0_reg[117][6]/P0001 ,
		_w11933_,
		_w12012_,
		_w22884_
	);
	LUT3 #(
		.INIT('h80)
	) name12372 (
		\wishbone_bd_ram_mem0_reg[241][6]/P0001 ,
		_w11952_,
		_w11977_,
		_w22885_
	);
	LUT3 #(
		.INIT('h80)
	) name12373 (
		\wishbone_bd_ram_mem0_reg[248][6]/P0001 ,
		_w11952_,
		_w11990_,
		_w22886_
	);
	LUT4 #(
		.INIT('h0001)
	) name12374 (
		_w22883_,
		_w22884_,
		_w22885_,
		_w22886_,
		_w22887_
	);
	LUT3 #(
		.INIT('h80)
	) name12375 (
		\wishbone_bd_ram_mem0_reg[53][6]/P0001 ,
		_w11933_,
		_w11979_,
		_w22888_
	);
	LUT3 #(
		.INIT('h80)
	) name12376 (
		\wishbone_bd_ram_mem0_reg[187][6]/P0001 ,
		_w11936_,
		_w11942_,
		_w22889_
	);
	LUT3 #(
		.INIT('h80)
	) name12377 (
		\wishbone_bd_ram_mem0_reg[36][6]/P0001 ,
		_w11929_,
		_w11957_,
		_w22890_
	);
	LUT3 #(
		.INIT('h80)
	) name12378 (
		\wishbone_bd_ram_mem0_reg[155][6]/P0001 ,
		_w11936_,
		_w11959_,
		_w22891_
	);
	LUT4 #(
		.INIT('h0001)
	) name12379 (
		_w22888_,
		_w22889_,
		_w22890_,
		_w22891_,
		_w22892_
	);
	LUT3 #(
		.INIT('h80)
	) name12380 (
		\wishbone_bd_ram_mem0_reg[211][6]/P0001 ,
		_w11938_,
		_w11984_,
		_w22893_
	);
	LUT3 #(
		.INIT('h80)
	) name12381 (
		\wishbone_bd_ram_mem0_reg[81][6]/P0001 ,
		_w11972_,
		_w11977_,
		_w22894_
	);
	LUT3 #(
		.INIT('h80)
	) name12382 (
		\wishbone_bd_ram_mem0_reg[35][6]/P0001 ,
		_w11938_,
		_w11957_,
		_w22895_
	);
	LUT3 #(
		.INIT('h80)
	) name12383 (
		\wishbone_bd_ram_mem0_reg[238][6]/P0001 ,
		_w11948_,
		_w11982_,
		_w22896_
	);
	LUT4 #(
		.INIT('h0001)
	) name12384 (
		_w22893_,
		_w22894_,
		_w22895_,
		_w22896_,
		_w22897_
	);
	LUT3 #(
		.INIT('h80)
	) name12385 (
		\wishbone_bd_ram_mem0_reg[244][6]/P0001 ,
		_w11929_,
		_w11952_,
		_w22898_
	);
	LUT3 #(
		.INIT('h80)
	) name12386 (
		\wishbone_bd_ram_mem0_reg[215][6]/P0001 ,
		_w11975_,
		_w11984_,
		_w22899_
	);
	LUT3 #(
		.INIT('h80)
	) name12387 (
		\wishbone_bd_ram_mem0_reg[153][6]/P0001 ,
		_w11959_,
		_w11968_,
		_w22900_
	);
	LUT3 #(
		.INIT('h80)
	) name12388 (
		\wishbone_bd_ram_mem0_reg[131][6]/P0001 ,
		_w11938_,
		_w11955_,
		_w22901_
	);
	LUT4 #(
		.INIT('h0001)
	) name12389 (
		_w22898_,
		_w22899_,
		_w22900_,
		_w22901_,
		_w22902_
	);
	LUT4 #(
		.INIT('h8000)
	) name12390 (
		_w22887_,
		_w22892_,
		_w22897_,
		_w22902_,
		_w22903_
	);
	LUT4 #(
		.INIT('h8000)
	) name12391 (
		_w22840_,
		_w22861_,
		_w22882_,
		_w22903_,
		_w22904_
	);
	LUT3 #(
		.INIT('h80)
	) name12392 (
		\wishbone_bd_ram_mem0_reg[50][6]/P0001 ,
		_w11963_,
		_w11979_,
		_w22905_
	);
	LUT3 #(
		.INIT('h80)
	) name12393 (
		\wishbone_bd_ram_mem0_reg[12][6]/P0001 ,
		_w11932_,
		_w11954_,
		_w22906_
	);
	LUT3 #(
		.INIT('h80)
	) name12394 (
		\wishbone_bd_ram_mem0_reg[99][6]/P0001 ,
		_w11938_,
		_w11965_,
		_w22907_
	);
	LUT3 #(
		.INIT('h80)
	) name12395 (
		\wishbone_bd_ram_mem0_reg[206][6]/P0001 ,
		_w11945_,
		_w11948_,
		_w22908_
	);
	LUT4 #(
		.INIT('h0001)
	) name12396 (
		_w22905_,
		_w22906_,
		_w22907_,
		_w22908_,
		_w22909_
	);
	LUT3 #(
		.INIT('h80)
	) name12397 (
		\wishbone_bd_ram_mem0_reg[141][6]/P0001 ,
		_w11955_,
		_w11966_,
		_w22910_
	);
	LUT3 #(
		.INIT('h80)
	) name12398 (
		\wishbone_bd_ram_mem0_reg[40][6]/P0001 ,
		_w11957_,
		_w11990_,
		_w22911_
	);
	LUT3 #(
		.INIT('h80)
	) name12399 (
		\wishbone_bd_ram_mem0_reg[229][6]/P0001 ,
		_w11933_,
		_w11982_,
		_w22912_
	);
	LUT3 #(
		.INIT('h80)
	) name12400 (
		\wishbone_bd_ram_mem0_reg[57][6]/P0001 ,
		_w11968_,
		_w11979_,
		_w22913_
	);
	LUT4 #(
		.INIT('h0001)
	) name12401 (
		_w22910_,
		_w22911_,
		_w22912_,
		_w22913_,
		_w22914_
	);
	LUT3 #(
		.INIT('h80)
	) name12402 (
		\wishbone_bd_ram_mem0_reg[143][6]/P0001 ,
		_w11955_,
		_w11973_,
		_w22915_
	);
	LUT3 #(
		.INIT('h80)
	) name12403 (
		\wishbone_bd_ram_mem0_reg[17][6]/P0001 ,
		_w11935_,
		_w11977_,
		_w22916_
	);
	LUT3 #(
		.INIT('h80)
	) name12404 (
		\wishbone_bd_ram_mem0_reg[236][6]/P0001 ,
		_w11954_,
		_w11982_,
		_w22917_
	);
	LUT3 #(
		.INIT('h80)
	) name12405 (
		\wishbone_bd_ram_mem0_reg[168][6]/P0001 ,
		_w11930_,
		_w11990_,
		_w22918_
	);
	LUT4 #(
		.INIT('h0001)
	) name12406 (
		_w22915_,
		_w22916_,
		_w22917_,
		_w22918_,
		_w22919_
	);
	LUT3 #(
		.INIT('h80)
	) name12407 (
		\wishbone_bd_ram_mem0_reg[148][6]/P0001 ,
		_w11929_,
		_w11959_,
		_w22920_
	);
	LUT3 #(
		.INIT('h80)
	) name12408 (
		\wishbone_bd_ram_mem0_reg[132][6]/P0001 ,
		_w11929_,
		_w11955_,
		_w22921_
	);
	LUT3 #(
		.INIT('h80)
	) name12409 (
		\wishbone_bd_ram_mem0_reg[124][6]/P0001 ,
		_w11954_,
		_w12012_,
		_w22922_
	);
	LUT3 #(
		.INIT('h80)
	) name12410 (
		\wishbone_bd_ram_mem0_reg[163][6]/P0001 ,
		_w11930_,
		_w11938_,
		_w22923_
	);
	LUT4 #(
		.INIT('h0001)
	) name12411 (
		_w22920_,
		_w22921_,
		_w22922_,
		_w22923_,
		_w22924_
	);
	LUT4 #(
		.INIT('h8000)
	) name12412 (
		_w22909_,
		_w22914_,
		_w22919_,
		_w22924_,
		_w22925_
	);
	LUT3 #(
		.INIT('h80)
	) name12413 (
		\wishbone_bd_ram_mem0_reg[240][6]/P0001 ,
		_w11941_,
		_w11952_,
		_w22926_
	);
	LUT3 #(
		.INIT('h80)
	) name12414 (
		\wishbone_bd_ram_mem0_reg[68][6]/P0001 ,
		_w11929_,
		_w11949_,
		_w22927_
	);
	LUT3 #(
		.INIT('h80)
	) name12415 (
		\wishbone_bd_ram_mem0_reg[28][6]/P0001 ,
		_w11935_,
		_w11954_,
		_w22928_
	);
	LUT3 #(
		.INIT('h80)
	) name12416 (
		\wishbone_bd_ram_mem0_reg[103][6]/P0001 ,
		_w11965_,
		_w11975_,
		_w22929_
	);
	LUT4 #(
		.INIT('h0001)
	) name12417 (
		_w22926_,
		_w22927_,
		_w22928_,
		_w22929_,
		_w22930_
	);
	LUT3 #(
		.INIT('h80)
	) name12418 (
		\wishbone_bd_ram_mem0_reg[246][6]/P0001 ,
		_w11952_,
		_w11986_,
		_w22931_
	);
	LUT3 #(
		.INIT('h80)
	) name12419 (
		\wishbone_bd_ram_mem0_reg[110][6]/P0001 ,
		_w11948_,
		_w11965_,
		_w22932_
	);
	LUT3 #(
		.INIT('h80)
	) name12420 (
		\wishbone_bd_ram_mem0_reg[91][6]/P0001 ,
		_w11936_,
		_w11972_,
		_w22933_
	);
	LUT3 #(
		.INIT('h80)
	) name12421 (
		\wishbone_bd_ram_mem0_reg[234][6]/P0001 ,
		_w11944_,
		_w11982_,
		_w22934_
	);
	LUT4 #(
		.INIT('h0001)
	) name12422 (
		_w22931_,
		_w22932_,
		_w22933_,
		_w22934_,
		_w22935_
	);
	LUT3 #(
		.INIT('h80)
	) name12423 (
		\wishbone_bd_ram_mem0_reg[95][6]/P0001 ,
		_w11972_,
		_w11973_,
		_w22936_
	);
	LUT3 #(
		.INIT('h80)
	) name12424 (
		\wishbone_bd_ram_mem0_reg[8][6]/P0001 ,
		_w11932_,
		_w11990_,
		_w22937_
	);
	LUT3 #(
		.INIT('h80)
	) name12425 (
		\wishbone_bd_ram_mem0_reg[70][6]/P0001 ,
		_w11949_,
		_w11986_,
		_w22938_
	);
	LUT3 #(
		.INIT('h80)
	) name12426 (
		\wishbone_bd_ram_mem0_reg[83][6]/P0001 ,
		_w11938_,
		_w11972_,
		_w22939_
	);
	LUT4 #(
		.INIT('h0001)
	) name12427 (
		_w22936_,
		_w22937_,
		_w22938_,
		_w22939_,
		_w22940_
	);
	LUT3 #(
		.INIT('h80)
	) name12428 (
		\wishbone_bd_ram_mem0_reg[101][6]/P0001 ,
		_w11933_,
		_w11965_,
		_w22941_
	);
	LUT3 #(
		.INIT('h80)
	) name12429 (
		\wishbone_bd_ram_mem0_reg[7][6]/P0001 ,
		_w11932_,
		_w11975_,
		_w22942_
	);
	LUT3 #(
		.INIT('h80)
	) name12430 (
		\wishbone_bd_ram_mem0_reg[142][6]/P0001 ,
		_w11948_,
		_w11955_,
		_w22943_
	);
	LUT3 #(
		.INIT('h80)
	) name12431 (
		\wishbone_bd_ram_mem0_reg[54][6]/P0001 ,
		_w11979_,
		_w11986_,
		_w22944_
	);
	LUT4 #(
		.INIT('h0001)
	) name12432 (
		_w22941_,
		_w22942_,
		_w22943_,
		_w22944_,
		_w22945_
	);
	LUT4 #(
		.INIT('h8000)
	) name12433 (
		_w22930_,
		_w22935_,
		_w22940_,
		_w22945_,
		_w22946_
	);
	LUT3 #(
		.INIT('h80)
	) name12434 (
		\wishbone_bd_ram_mem0_reg[226][6]/P0001 ,
		_w11963_,
		_w11982_,
		_w22947_
	);
	LUT3 #(
		.INIT('h80)
	) name12435 (
		\wishbone_bd_ram_mem0_reg[23][6]/P0001 ,
		_w11935_,
		_w11975_,
		_w22948_
	);
	LUT3 #(
		.INIT('h80)
	) name12436 (
		\wishbone_bd_ram_mem0_reg[30][6]/P0001 ,
		_w11935_,
		_w11948_,
		_w22949_
	);
	LUT3 #(
		.INIT('h80)
	) name12437 (
		\wishbone_bd_ram_mem0_reg[209][6]/P0001 ,
		_w11977_,
		_w11984_,
		_w22950_
	);
	LUT4 #(
		.INIT('h0001)
	) name12438 (
		_w22947_,
		_w22948_,
		_w22949_,
		_w22950_,
		_w22951_
	);
	LUT3 #(
		.INIT('h80)
	) name12439 (
		\wishbone_bd_ram_mem0_reg[245][6]/P0001 ,
		_w11933_,
		_w11952_,
		_w22952_
	);
	LUT3 #(
		.INIT('h80)
	) name12440 (
		\wishbone_bd_ram_mem0_reg[166][6]/P0001 ,
		_w11930_,
		_w11986_,
		_w22953_
	);
	LUT3 #(
		.INIT('h80)
	) name12441 (
		\wishbone_bd_ram_mem0_reg[97][6]/P0001 ,
		_w11965_,
		_w11977_,
		_w22954_
	);
	LUT3 #(
		.INIT('h80)
	) name12442 (
		\wishbone_bd_ram_mem0_reg[31][6]/P0001 ,
		_w11935_,
		_w11973_,
		_w22955_
	);
	LUT4 #(
		.INIT('h0001)
	) name12443 (
		_w22952_,
		_w22953_,
		_w22954_,
		_w22955_,
		_w22956_
	);
	LUT3 #(
		.INIT('h80)
	) name12444 (
		\wishbone_bd_ram_mem0_reg[69][6]/P0001 ,
		_w11933_,
		_w11949_,
		_w22957_
	);
	LUT3 #(
		.INIT('h80)
	) name12445 (
		\wishbone_bd_ram_mem0_reg[195][6]/P0001 ,
		_w11938_,
		_w11945_,
		_w22958_
	);
	LUT3 #(
		.INIT('h80)
	) name12446 (
		\wishbone_bd_ram_mem0_reg[160][6]/P0001 ,
		_w11930_,
		_w11941_,
		_w22959_
	);
	LUT3 #(
		.INIT('h80)
	) name12447 (
		\wishbone_bd_ram_mem0_reg[175][6]/P0001 ,
		_w11930_,
		_w11973_,
		_w22960_
	);
	LUT4 #(
		.INIT('h0001)
	) name12448 (
		_w22957_,
		_w22958_,
		_w22959_,
		_w22960_,
		_w22961_
	);
	LUT3 #(
		.INIT('h80)
	) name12449 (
		\wishbone_bd_ram_mem0_reg[157][6]/P0001 ,
		_w11959_,
		_w11966_,
		_w22962_
	);
	LUT3 #(
		.INIT('h80)
	) name12450 (
		\wishbone_bd_ram_mem0_reg[122][6]/P0001 ,
		_w11944_,
		_w12012_,
		_w22963_
	);
	LUT3 #(
		.INIT('h80)
	) name12451 (
		\wishbone_bd_ram_mem0_reg[167][6]/P0001 ,
		_w11930_,
		_w11975_,
		_w22964_
	);
	LUT3 #(
		.INIT('h80)
	) name12452 (
		\wishbone_bd_ram_mem0_reg[41][6]/P0001 ,
		_w11957_,
		_w11968_,
		_w22965_
	);
	LUT4 #(
		.INIT('h0001)
	) name12453 (
		_w22962_,
		_w22963_,
		_w22964_,
		_w22965_,
		_w22966_
	);
	LUT4 #(
		.INIT('h8000)
	) name12454 (
		_w22951_,
		_w22956_,
		_w22961_,
		_w22966_,
		_w22967_
	);
	LUT3 #(
		.INIT('h80)
	) name12455 (
		\wishbone_bd_ram_mem0_reg[242][6]/P0001 ,
		_w11952_,
		_w11963_,
		_w22968_
	);
	LUT3 #(
		.INIT('h80)
	) name12456 (
		\wishbone_bd_ram_mem0_reg[220][6]/P0001 ,
		_w11954_,
		_w11984_,
		_w22969_
	);
	LUT3 #(
		.INIT('h80)
	) name12457 (
		\wishbone_bd_ram_mem0_reg[123][6]/P0001 ,
		_w11936_,
		_w12012_,
		_w22970_
	);
	LUT3 #(
		.INIT('h80)
	) name12458 (
		\wishbone_bd_ram_mem0_reg[6][6]/P0001 ,
		_w11932_,
		_w11986_,
		_w22971_
	);
	LUT4 #(
		.INIT('h0001)
	) name12459 (
		_w22968_,
		_w22969_,
		_w22970_,
		_w22971_,
		_w22972_
	);
	LUT3 #(
		.INIT('h80)
	) name12460 (
		\wishbone_bd_ram_mem0_reg[189][6]/P0001 ,
		_w11942_,
		_w11966_,
		_w22973_
	);
	LUT3 #(
		.INIT('h80)
	) name12461 (
		\wishbone_bd_ram_mem0_reg[55][6]/P0001 ,
		_w11975_,
		_w11979_,
		_w22974_
	);
	LUT3 #(
		.INIT('h80)
	) name12462 (
		\wishbone_bd_ram_mem0_reg[190][6]/P0001 ,
		_w11942_,
		_w11948_,
		_w22975_
	);
	LUT3 #(
		.INIT('h80)
	) name12463 (
		\wishbone_bd_ram_mem0_reg[170][6]/P0001 ,
		_w11930_,
		_w11944_,
		_w22976_
	);
	LUT4 #(
		.INIT('h0001)
	) name12464 (
		_w22973_,
		_w22974_,
		_w22975_,
		_w22976_,
		_w22977_
	);
	LUT3 #(
		.INIT('h80)
	) name12465 (
		\wishbone_bd_ram_mem0_reg[250][6]/P0001 ,
		_w11944_,
		_w11952_,
		_w22978_
	);
	LUT3 #(
		.INIT('h80)
	) name12466 (
		\wishbone_bd_ram_mem0_reg[119][6]/P0001 ,
		_w11975_,
		_w12012_,
		_w22979_
	);
	LUT3 #(
		.INIT('h80)
	) name12467 (
		\wishbone_bd_ram_mem0_reg[159][6]/P0001 ,
		_w11959_,
		_w11973_,
		_w22980_
	);
	LUT3 #(
		.INIT('h80)
	) name12468 (
		\wishbone_bd_ram_mem0_reg[232][6]/P0001 ,
		_w11982_,
		_w11990_,
		_w22981_
	);
	LUT4 #(
		.INIT('h0001)
	) name12469 (
		_w22978_,
		_w22979_,
		_w22980_,
		_w22981_,
		_w22982_
	);
	LUT3 #(
		.INIT('h80)
	) name12470 (
		\wishbone_bd_ram_mem0_reg[75][6]/P0001 ,
		_w11936_,
		_w11949_,
		_w22983_
	);
	LUT3 #(
		.INIT('h80)
	) name12471 (
		\wishbone_bd_ram_mem0_reg[47][6]/P0001 ,
		_w11957_,
		_w11973_,
		_w22984_
	);
	LUT3 #(
		.INIT('h80)
	) name12472 (
		\wishbone_bd_ram_mem0_reg[42][6]/P0001 ,
		_w11944_,
		_w11957_,
		_w22985_
	);
	LUT3 #(
		.INIT('h80)
	) name12473 (
		\wishbone_bd_ram_mem0_reg[0][6]/P0001 ,
		_w11932_,
		_w11941_,
		_w22986_
	);
	LUT4 #(
		.INIT('h0001)
	) name12474 (
		_w22983_,
		_w22984_,
		_w22985_,
		_w22986_,
		_w22987_
	);
	LUT4 #(
		.INIT('h8000)
	) name12475 (
		_w22972_,
		_w22977_,
		_w22982_,
		_w22987_,
		_w22988_
	);
	LUT4 #(
		.INIT('h8000)
	) name12476 (
		_w22925_,
		_w22946_,
		_w22967_,
		_w22988_,
		_w22989_
	);
	LUT3 #(
		.INIT('h80)
	) name12477 (
		\wishbone_bd_ram_mem0_reg[34][6]/P0001 ,
		_w11957_,
		_w11963_,
		_w22990_
	);
	LUT3 #(
		.INIT('h80)
	) name12478 (
		\wishbone_bd_ram_mem0_reg[222][6]/P0001 ,
		_w11948_,
		_w11984_,
		_w22991_
	);
	LUT3 #(
		.INIT('h80)
	) name12479 (
		\wishbone_bd_ram_mem0_reg[152][6]/P0001 ,
		_w11959_,
		_w11990_,
		_w22992_
	);
	LUT3 #(
		.INIT('h80)
	) name12480 (
		\wishbone_bd_ram_mem0_reg[93][6]/P0001 ,
		_w11966_,
		_w11972_,
		_w22993_
	);
	LUT4 #(
		.INIT('h0001)
	) name12481 (
		_w22990_,
		_w22991_,
		_w22992_,
		_w22993_,
		_w22994_
	);
	LUT3 #(
		.INIT('h80)
	) name12482 (
		\wishbone_bd_ram_mem0_reg[102][6]/P0001 ,
		_w11965_,
		_w11986_,
		_w22995_
	);
	LUT3 #(
		.INIT('h80)
	) name12483 (
		\wishbone_bd_ram_mem0_reg[129][6]/P0001 ,
		_w11955_,
		_w11977_,
		_w22996_
	);
	LUT3 #(
		.INIT('h80)
	) name12484 (
		\wishbone_bd_ram_mem0_reg[164][6]/P0001 ,
		_w11929_,
		_w11930_,
		_w22997_
	);
	LUT3 #(
		.INIT('h80)
	) name12485 (
		\wishbone_bd_ram_mem0_reg[233][6]/P0001 ,
		_w11968_,
		_w11982_,
		_w22998_
	);
	LUT4 #(
		.INIT('h0001)
	) name12486 (
		_w22995_,
		_w22996_,
		_w22997_,
		_w22998_,
		_w22999_
	);
	LUT3 #(
		.INIT('h80)
	) name12487 (
		\wishbone_bd_ram_mem0_reg[136][6]/P0001 ,
		_w11955_,
		_w11990_,
		_w23000_
	);
	LUT3 #(
		.INIT('h80)
	) name12488 (
		\wishbone_bd_ram_mem0_reg[239][6]/P0001 ,
		_w11973_,
		_w11982_,
		_w23001_
	);
	LUT3 #(
		.INIT('h80)
	) name12489 (
		\wishbone_bd_ram_mem0_reg[25][6]/P0001 ,
		_w11935_,
		_w11968_,
		_w23002_
	);
	LUT3 #(
		.INIT('h80)
	) name12490 (
		\wishbone_bd_ram_mem0_reg[106][6]/P0001 ,
		_w11944_,
		_w11965_,
		_w23003_
	);
	LUT4 #(
		.INIT('h0001)
	) name12491 (
		_w23000_,
		_w23001_,
		_w23002_,
		_w23003_,
		_w23004_
	);
	LUT3 #(
		.INIT('h80)
	) name12492 (
		\wishbone_bd_ram_mem0_reg[14][6]/P0001 ,
		_w11932_,
		_w11948_,
		_w23005_
	);
	LUT3 #(
		.INIT('h80)
	) name12493 (
		\wishbone_bd_ram_mem0_reg[5][6]/P0001 ,
		_w11932_,
		_w11933_,
		_w23006_
	);
	LUT3 #(
		.INIT('h80)
	) name12494 (
		\wishbone_bd_ram_mem0_reg[134][6]/P0001 ,
		_w11955_,
		_w11986_,
		_w23007_
	);
	LUT3 #(
		.INIT('h80)
	) name12495 (
		\wishbone_bd_ram_mem0_reg[77][6]/P0001 ,
		_w11949_,
		_w11966_,
		_w23008_
	);
	LUT4 #(
		.INIT('h0001)
	) name12496 (
		_w23005_,
		_w23006_,
		_w23007_,
		_w23008_,
		_w23009_
	);
	LUT4 #(
		.INIT('h8000)
	) name12497 (
		_w22994_,
		_w22999_,
		_w23004_,
		_w23009_,
		_w23010_
	);
	LUT3 #(
		.INIT('h80)
	) name12498 (
		\wishbone_bd_ram_mem0_reg[180][6]/P0001 ,
		_w11929_,
		_w11942_,
		_w23011_
	);
	LUT3 #(
		.INIT('h80)
	) name12499 (
		\wishbone_bd_ram_mem0_reg[46][6]/P0001 ,
		_w11948_,
		_w11957_,
		_w23012_
	);
	LUT3 #(
		.INIT('h80)
	) name12500 (
		\wishbone_bd_ram_mem0_reg[78][6]/P0001 ,
		_w11948_,
		_w11949_,
		_w23013_
	);
	LUT3 #(
		.INIT('h80)
	) name12501 (
		\wishbone_bd_ram_mem0_reg[230][6]/P0001 ,
		_w11982_,
		_w11986_,
		_w23014_
	);
	LUT4 #(
		.INIT('h0001)
	) name12502 (
		_w23011_,
		_w23012_,
		_w23013_,
		_w23014_,
		_w23015_
	);
	LUT3 #(
		.INIT('h80)
	) name12503 (
		\wishbone_bd_ram_mem0_reg[107][6]/P0001 ,
		_w11936_,
		_w11965_,
		_w23016_
	);
	LUT3 #(
		.INIT('h80)
	) name12504 (
		\wishbone_bd_ram_mem0_reg[165][6]/P0001 ,
		_w11930_,
		_w11933_,
		_w23017_
	);
	LUT3 #(
		.INIT('h80)
	) name12505 (
		\wishbone_bd_ram_mem0_reg[15][6]/P0001 ,
		_w11932_,
		_w11973_,
		_w23018_
	);
	LUT3 #(
		.INIT('h80)
	) name12506 (
		\wishbone_bd_ram_mem0_reg[115][6]/P0001 ,
		_w11938_,
		_w12012_,
		_w23019_
	);
	LUT4 #(
		.INIT('h0001)
	) name12507 (
		_w23016_,
		_w23017_,
		_w23018_,
		_w23019_,
		_w23020_
	);
	LUT3 #(
		.INIT('h80)
	) name12508 (
		\wishbone_bd_ram_mem0_reg[140][6]/P0001 ,
		_w11954_,
		_w11955_,
		_w23021_
	);
	LUT3 #(
		.INIT('h80)
	) name12509 (
		\wishbone_bd_ram_mem0_reg[202][6]/P0001 ,
		_w11944_,
		_w11945_,
		_w23022_
	);
	LUT3 #(
		.INIT('h80)
	) name12510 (
		\wishbone_bd_ram_mem0_reg[112][6]/P0001 ,
		_w11941_,
		_w12012_,
		_w23023_
	);
	LUT3 #(
		.INIT('h80)
	) name12511 (
		\wishbone_bd_ram_mem0_reg[135][6]/P0001 ,
		_w11955_,
		_w11975_,
		_w23024_
	);
	LUT4 #(
		.INIT('h0001)
	) name12512 (
		_w23021_,
		_w23022_,
		_w23023_,
		_w23024_,
		_w23025_
	);
	LUT3 #(
		.INIT('h80)
	) name12513 (
		\wishbone_bd_ram_mem0_reg[43][6]/P0001 ,
		_w11936_,
		_w11957_,
		_w23026_
	);
	LUT3 #(
		.INIT('h80)
	) name12514 (
		\wishbone_bd_ram_mem0_reg[86][6]/P0001 ,
		_w11972_,
		_w11986_,
		_w23027_
	);
	LUT3 #(
		.INIT('h80)
	) name12515 (
		\wishbone_bd_ram_mem0_reg[213][6]/P0001 ,
		_w11933_,
		_w11984_,
		_w23028_
	);
	LUT3 #(
		.INIT('h80)
	) name12516 (
		\wishbone_bd_ram_mem0_reg[150][6]/P0001 ,
		_w11959_,
		_w11986_,
		_w23029_
	);
	LUT4 #(
		.INIT('h0001)
	) name12517 (
		_w23026_,
		_w23027_,
		_w23028_,
		_w23029_,
		_w23030_
	);
	LUT4 #(
		.INIT('h8000)
	) name12518 (
		_w23015_,
		_w23020_,
		_w23025_,
		_w23030_,
		_w23031_
	);
	LUT3 #(
		.INIT('h80)
	) name12519 (
		\wishbone_bd_ram_mem0_reg[173][6]/P0001 ,
		_w11930_,
		_w11966_,
		_w23032_
	);
	LUT3 #(
		.INIT('h80)
	) name12520 (
		\wishbone_bd_ram_mem0_reg[67][6]/P0001 ,
		_w11938_,
		_w11949_,
		_w23033_
	);
	LUT3 #(
		.INIT('h80)
	) name12521 (
		\wishbone_bd_ram_mem0_reg[205][6]/P0001 ,
		_w11945_,
		_w11966_,
		_w23034_
	);
	LUT3 #(
		.INIT('h80)
	) name12522 (
		\wishbone_bd_ram_mem0_reg[158][6]/P0001 ,
		_w11948_,
		_w11959_,
		_w23035_
	);
	LUT4 #(
		.INIT('h0001)
	) name12523 (
		_w23032_,
		_w23033_,
		_w23034_,
		_w23035_,
		_w23036_
	);
	LUT3 #(
		.INIT('h80)
	) name12524 (
		\wishbone_bd_ram_mem0_reg[192][6]/P0001 ,
		_w11941_,
		_w11945_,
		_w23037_
	);
	LUT3 #(
		.INIT('h80)
	) name12525 (
		\wishbone_bd_ram_mem0_reg[169][6]/P0001 ,
		_w11930_,
		_w11968_,
		_w23038_
	);
	LUT3 #(
		.INIT('h80)
	) name12526 (
		\wishbone_bd_ram_mem0_reg[201][6]/P0001 ,
		_w11945_,
		_w11968_,
		_w23039_
	);
	LUT3 #(
		.INIT('h80)
	) name12527 (
		\wishbone_bd_ram_mem0_reg[200][6]/P0001 ,
		_w11945_,
		_w11990_,
		_w23040_
	);
	LUT4 #(
		.INIT('h0001)
	) name12528 (
		_w23037_,
		_w23038_,
		_w23039_,
		_w23040_,
		_w23041_
	);
	LUT3 #(
		.INIT('h80)
	) name12529 (
		\wishbone_bd_ram_mem0_reg[16][6]/P0001 ,
		_w11935_,
		_w11941_,
		_w23042_
	);
	LUT3 #(
		.INIT('h80)
	) name12530 (
		\wishbone_bd_ram_mem0_reg[11][6]/P0001 ,
		_w11932_,
		_w11936_,
		_w23043_
	);
	LUT3 #(
		.INIT('h80)
	) name12531 (
		\wishbone_bd_ram_mem0_reg[24][6]/P0001 ,
		_w11935_,
		_w11990_,
		_w23044_
	);
	LUT3 #(
		.INIT('h80)
	) name12532 (
		\wishbone_bd_ram_mem0_reg[184][6]/P0001 ,
		_w11942_,
		_w11990_,
		_w23045_
	);
	LUT4 #(
		.INIT('h0001)
	) name12533 (
		_w23042_,
		_w23043_,
		_w23044_,
		_w23045_,
		_w23046_
	);
	LUT3 #(
		.INIT('h80)
	) name12534 (
		\wishbone_bd_ram_mem0_reg[214][6]/P0001 ,
		_w11984_,
		_w11986_,
		_w23047_
	);
	LUT3 #(
		.INIT('h80)
	) name12535 (
		\wishbone_bd_ram_mem0_reg[108][6]/P0001 ,
		_w11954_,
		_w11965_,
		_w23048_
	);
	LUT3 #(
		.INIT('h80)
	) name12536 (
		\wishbone_bd_ram_mem0_reg[10][6]/P0001 ,
		_w11932_,
		_w11944_,
		_w23049_
	);
	LUT3 #(
		.INIT('h80)
	) name12537 (
		\wishbone_bd_ram_mem0_reg[27][6]/P0001 ,
		_w11935_,
		_w11936_,
		_w23050_
	);
	LUT4 #(
		.INIT('h0001)
	) name12538 (
		_w23047_,
		_w23048_,
		_w23049_,
		_w23050_,
		_w23051_
	);
	LUT4 #(
		.INIT('h8000)
	) name12539 (
		_w23036_,
		_w23041_,
		_w23046_,
		_w23051_,
		_w23052_
	);
	LUT3 #(
		.INIT('h80)
	) name12540 (
		\wishbone_bd_ram_mem0_reg[39][6]/P0001 ,
		_w11957_,
		_w11975_,
		_w23053_
	);
	LUT3 #(
		.INIT('h80)
	) name12541 (
		\wishbone_bd_ram_mem0_reg[116][6]/P0001 ,
		_w11929_,
		_w12012_,
		_w23054_
	);
	LUT3 #(
		.INIT('h80)
	) name12542 (
		\wishbone_bd_ram_mem0_reg[90][6]/P0001 ,
		_w11944_,
		_w11972_,
		_w23055_
	);
	LUT3 #(
		.INIT('h80)
	) name12543 (
		\wishbone_bd_ram_mem0_reg[156][6]/P0001 ,
		_w11954_,
		_w11959_,
		_w23056_
	);
	LUT4 #(
		.INIT('h0001)
	) name12544 (
		_w23053_,
		_w23054_,
		_w23055_,
		_w23056_,
		_w23057_
	);
	LUT3 #(
		.INIT('h80)
	) name12545 (
		\wishbone_bd_ram_mem0_reg[251][6]/P0001 ,
		_w11936_,
		_w11952_,
		_w23058_
	);
	LUT3 #(
		.INIT('h80)
	) name12546 (
		\wishbone_bd_ram_mem0_reg[235][6]/P0001 ,
		_w11936_,
		_w11982_,
		_w23059_
	);
	LUT3 #(
		.INIT('h80)
	) name12547 (
		\wishbone_bd_ram_mem0_reg[111][6]/P0001 ,
		_w11965_,
		_w11973_,
		_w23060_
	);
	LUT3 #(
		.INIT('h80)
	) name12548 (
		\wishbone_bd_ram_mem0_reg[247][6]/P0001 ,
		_w11952_,
		_w11975_,
		_w23061_
	);
	LUT4 #(
		.INIT('h0001)
	) name12549 (
		_w23058_,
		_w23059_,
		_w23060_,
		_w23061_,
		_w23062_
	);
	LUT3 #(
		.INIT('h80)
	) name12550 (
		\wishbone_bd_ram_mem0_reg[48][6]/P0001 ,
		_w11941_,
		_w11979_,
		_w23063_
	);
	LUT3 #(
		.INIT('h80)
	) name12551 (
		\wishbone_bd_ram_mem0_reg[253][6]/P0001 ,
		_w11952_,
		_w11966_,
		_w23064_
	);
	LUT3 #(
		.INIT('h80)
	) name12552 (
		\wishbone_bd_ram_mem0_reg[172][6]/P0001 ,
		_w11930_,
		_w11954_,
		_w23065_
	);
	LUT3 #(
		.INIT('h80)
	) name12553 (
		\wishbone_bd_ram_mem0_reg[228][6]/P0001 ,
		_w11929_,
		_w11982_,
		_w23066_
	);
	LUT4 #(
		.INIT('h0001)
	) name12554 (
		_w23063_,
		_w23064_,
		_w23065_,
		_w23066_,
		_w23067_
	);
	LUT3 #(
		.INIT('h80)
	) name12555 (
		\wishbone_bd_ram_mem0_reg[82][6]/P0001 ,
		_w11963_,
		_w11972_,
		_w23068_
	);
	LUT3 #(
		.INIT('h80)
	) name12556 (
		\wishbone_bd_ram_mem0_reg[105][6]/P0001 ,
		_w11965_,
		_w11968_,
		_w23069_
	);
	LUT3 #(
		.INIT('h80)
	) name12557 (
		\wishbone_bd_ram_mem0_reg[37][6]/P0001 ,
		_w11933_,
		_w11957_,
		_w23070_
	);
	LUT3 #(
		.INIT('h80)
	) name12558 (
		\wishbone_bd_ram_mem0_reg[185][6]/P0001 ,
		_w11942_,
		_w11968_,
		_w23071_
	);
	LUT4 #(
		.INIT('h0001)
	) name12559 (
		_w23068_,
		_w23069_,
		_w23070_,
		_w23071_,
		_w23072_
	);
	LUT4 #(
		.INIT('h8000)
	) name12560 (
		_w23057_,
		_w23062_,
		_w23067_,
		_w23072_,
		_w23073_
	);
	LUT4 #(
		.INIT('h8000)
	) name12561 (
		_w23010_,
		_w23031_,
		_w23052_,
		_w23073_,
		_w23074_
	);
	LUT4 #(
		.INIT('h8000)
	) name12562 (
		_w22819_,
		_w22904_,
		_w22989_,
		_w23074_,
		_w23075_
	);
	LUT3 #(
		.INIT('h15)
	) name12563 (
		wb_rst_i_pad,
		_w22714_,
		_w22733_,
		_w23076_
	);
	LUT3 #(
		.INIT('hba)
	) name12564 (
		_w22734_,
		_w23075_,
		_w23076_,
		_w23077_
	);
	LUT4 #(
		.INIT('h0008)
	) name12565 (
		\ethreg1_RXHASH1_2_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23078_
	);
	LUT3 #(
		.INIT('h80)
	) name12566 (
		_w18757_,
		_w18762_,
		_w23078_,
		_w23079_
	);
	LUT4 #(
		.INIT('h0002)
	) name12567 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23080_
	);
	LUT3 #(
		.INIT('h80)
	) name12568 (
		_w18757_,
		_w18758_,
		_w23080_,
		_w23081_
	);
	LUT4 #(
		.INIT('h0008)
	) name12569 (
		\ethreg1_RXHASH0_2_DataOut_reg[1]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23082_
	);
	LUT3 #(
		.INIT('h80)
	) name12570 (
		_w18757_,
		_w18758_,
		_w23082_,
		_w23083_
	);
	LUT4 #(
		.INIT('h0002)
	) name12571 (
		_w18752_,
		_w23079_,
		_w23081_,
		_w23083_,
		_w23084_
	);
	LUT3 #(
		.INIT('h80)
	) name12572 (
		\ethreg1_COLLCONF_2_DataOut_reg[1]/NET0131 ,
		_w18753_,
		_w19641_,
		_w23085_
	);
	LUT3 #(
		.INIT('h80)
	) name12573 (
		\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 ,
		_w18753_,
		_w18754_,
		_w23086_
	);
	LUT2 #(
		.INIT('h1)
	) name12574 (
		_w23085_,
		_w23086_,
		_w23087_
	);
	LUT3 #(
		.INIT('h2a)
	) name12575 (
		_w18752_,
		_w23084_,
		_w23087_,
		_w23088_
	);
	LUT3 #(
		.INIT('h15)
	) name12576 (
		wb_rst_i_pad,
		_w23084_,
		_w23087_,
		_w23089_
	);
	LUT3 #(
		.INIT('hdc)
	) name12577 (
		_w16814_,
		_w23088_,
		_w23089_,
		_w23090_
	);
	LUT4 #(
		.INIT('h0008)
	) name12578 (
		\ethreg1_RXHASH1_2_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23091_
	);
	LUT3 #(
		.INIT('h80)
	) name12579 (
		_w18757_,
		_w18762_,
		_w23091_,
		_w23092_
	);
	LUT4 #(
		.INIT('h0002)
	) name12580 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23093_
	);
	LUT3 #(
		.INIT('h80)
	) name12581 (
		_w18757_,
		_w18758_,
		_w23093_,
		_w23094_
	);
	LUT4 #(
		.INIT('h0008)
	) name12582 (
		\ethreg1_RXHASH0_2_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23095_
	);
	LUT3 #(
		.INIT('h80)
	) name12583 (
		_w18757_,
		_w18758_,
		_w23095_,
		_w23096_
	);
	LUT4 #(
		.INIT('h0002)
	) name12584 (
		_w18752_,
		_w23092_,
		_w23094_,
		_w23096_,
		_w23097_
	);
	LUT3 #(
		.INIT('h80)
	) name12585 (
		\ethreg1_COLLCONF_2_DataOut_reg[2]/NET0131 ,
		_w18753_,
		_w19641_,
		_w23098_
	);
	LUT3 #(
		.INIT('h80)
	) name12586 (
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		_w18753_,
		_w18754_,
		_w23099_
	);
	LUT2 #(
		.INIT('h1)
	) name12587 (
		_w23098_,
		_w23099_,
		_w23100_
	);
	LUT3 #(
		.INIT('h2a)
	) name12588 (
		_w18752_,
		_w23097_,
		_w23100_,
		_w23101_
	);
	LUT3 #(
		.INIT('h15)
	) name12589 (
		wb_rst_i_pad,
		_w23097_,
		_w23100_,
		_w23102_
	);
	LUT3 #(
		.INIT('hdc)
	) name12590 (
		_w15775_,
		_w23101_,
		_w23102_,
		_w23103_
	);
	LUT4 #(
		.INIT('h0008)
	) name12591 (
		\ethreg1_RXHASH1_2_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23104_
	);
	LUT3 #(
		.INIT('h80)
	) name12592 (
		_w18757_,
		_w18762_,
		_w23104_,
		_w23105_
	);
	LUT4 #(
		.INIT('h0002)
	) name12593 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23106_
	);
	LUT3 #(
		.INIT('h80)
	) name12594 (
		_w18757_,
		_w18758_,
		_w23106_,
		_w23107_
	);
	LUT4 #(
		.INIT('h0008)
	) name12595 (
		\ethreg1_RXHASH0_2_DataOut_reg[3]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23108_
	);
	LUT3 #(
		.INIT('h80)
	) name12596 (
		_w18757_,
		_w18758_,
		_w23108_,
		_w23109_
	);
	LUT4 #(
		.INIT('h0002)
	) name12597 (
		_w18752_,
		_w23105_,
		_w23107_,
		_w23109_,
		_w23110_
	);
	LUT3 #(
		.INIT('h80)
	) name12598 (
		\ethreg1_COLLCONF_2_DataOut_reg[3]/NET0131 ,
		_w18753_,
		_w19641_,
		_w23111_
	);
	LUT3 #(
		.INIT('h80)
	) name12599 (
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		_w18753_,
		_w18754_,
		_w23112_
	);
	LUT2 #(
		.INIT('h1)
	) name12600 (
		_w23111_,
		_w23112_,
		_w23113_
	);
	LUT3 #(
		.INIT('h2a)
	) name12601 (
		_w18752_,
		_w23110_,
		_w23113_,
		_w23114_
	);
	LUT3 #(
		.INIT('h15)
	) name12602 (
		wb_rst_i_pad,
		_w23110_,
		_w23113_,
		_w23115_
	);
	LUT3 #(
		.INIT('hdc)
	) name12603 (
		_w17713_,
		_w23114_,
		_w23115_,
		_w23116_
	);
	LUT3 #(
		.INIT('h80)
	) name12604 (
		\wishbone_RxPointerMSB_reg[15]/NET0131 ,
		\wishbone_RxPointerMSB_reg[16]/NET0131 ,
		\wishbone_RxPointerMSB_reg[17]/NET0131 ,
		_w23117_
	);
	LUT4 #(
		.INIT('h1333)
	) name12605 (
		\wishbone_RxPointerMSB_reg[18]/NET0131 ,
		\wishbone_RxPointerMSB_reg[19]/NET0131 ,
		_w15288_,
		_w23117_,
		_w23118_
	);
	LUT2 #(
		.INIT('h8)
	) name12606 (
		\wishbone_RxPointerMSB_reg[15]/NET0131 ,
		_w15289_,
		_w23119_
	);
	LUT3 #(
		.INIT('h15)
	) name12607 (
		_w13807_,
		_w15288_,
		_w23119_,
		_w23120_
	);
	LUT2 #(
		.INIT('h4)
	) name12608 (
		_w23118_,
		_w23120_,
		_w23121_
	);
	LUT3 #(
		.INIT('hf2)
	) name12609 (
		_w15282_,
		_w17713_,
		_w23121_,
		_w23122_
	);
	LUT3 #(
		.INIT('h15)
	) name12610 (
		\wishbone_RxPointerMSB_reg[20]/NET0131 ,
		_w15288_,
		_w23119_,
		_w23123_
	);
	LUT3 #(
		.INIT('h15)
	) name12611 (
		_w13807_,
		_w15288_,
		_w15291_,
		_w23124_
	);
	LUT2 #(
		.INIT('h4)
	) name12612 (
		_w23123_,
		_w23124_,
		_w23125_
	);
	LUT3 #(
		.INIT('hf4)
	) name12613 (
		_w14512_,
		_w15282_,
		_w23125_,
		_w23126_
	);
	LUT4 #(
		.INIT('heddd)
	) name12614 (
		\wishbone_RxPointerMSB_reg[21]/NET0131 ,
		_w13807_,
		_w15288_,
		_w15291_,
		_w23127_
	);
	LUT3 #(
		.INIT('h2f)
	) name12615 (
		_w15282_,
		_w18058_,
		_w23127_,
		_w23128_
	);
	LUT4 #(
		.INIT('h1333)
	) name12616 (
		\wishbone_RxPointerMSB_reg[21]/NET0131 ,
		\wishbone_RxPointerMSB_reg[22]/NET0131 ,
		_w15288_,
		_w15291_,
		_w23129_
	);
	LUT4 #(
		.INIT('h1555)
	) name12617 (
		_w13807_,
		_w15288_,
		_w15291_,
		_w15292_,
		_w23130_
	);
	LUT2 #(
		.INIT('h4)
	) name12618 (
		_w23129_,
		_w23130_,
		_w23131_
	);
	LUT3 #(
		.INIT('hf2)
	) name12619 (
		_w15282_,
		_w18746_,
		_w23131_,
		_w23132_
	);
	LUT4 #(
		.INIT('h1555)
	) name12620 (
		\wishbone_RxPointerMSB_reg[23]/NET0131 ,
		_w15288_,
		_w15291_,
		_w15292_,
		_w23133_
	);
	LUT3 #(
		.INIT('h80)
	) name12621 (
		\wishbone_RxPointerMSB_reg[21]/NET0131 ,
		\wishbone_RxPointerMSB_reg[22]/NET0131 ,
		\wishbone_RxPointerMSB_reg[23]/NET0131 ,
		_w23134_
	);
	LUT4 #(
		.INIT('h1555)
	) name12622 (
		_w13807_,
		_w15288_,
		_w15291_,
		_w23134_,
		_w23135_
	);
	LUT2 #(
		.INIT('h4)
	) name12623 (
		_w23133_,
		_w23135_,
		_w23136_
	);
	LUT3 #(
		.INIT('hf2)
	) name12624 (
		_w15282_,
		_w18401_,
		_w23136_,
		_w23137_
	);
	LUT4 #(
		.INIT('h1555)
	) name12625 (
		\wishbone_RxPointerMSB_reg[24]/NET0131 ,
		_w15288_,
		_w15291_,
		_w23134_,
		_w23138_
	);
	LUT4 #(
		.INIT('h1555)
	) name12626 (
		_w13807_,
		_w15288_,
		_w15291_,
		_w15293_,
		_w23139_
	);
	LUT2 #(
		.INIT('h4)
	) name12627 (
		_w23138_,
		_w23139_,
		_w23140_
	);
	LUT3 #(
		.INIT('hf4)
	) name12628 (
		_w13397_,
		_w15282_,
		_w23140_,
		_w23141_
	);
	LUT4 #(
		.INIT('h70f0)
	) name12629 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxPointerMSB_reg[25]/NET0131 ,
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w23142_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12630 (
		_w15288_,
		_w15291_,
		_w15293_,
		_w23142_,
		_w23143_
	);
	LUT4 #(
		.INIT('h070f)
	) name12631 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxPointerMSB_reg[25]/NET0131 ,
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w23144_
	);
	LUT4 #(
		.INIT('h8000)
	) name12632 (
		_w15288_,
		_w15291_,
		_w15293_,
		_w23144_,
		_w23145_
	);
	LUT2 #(
		.INIT('h1)
	) name12633 (
		_w23143_,
		_w23145_,
		_w23146_
	);
	LUT3 #(
		.INIT('h4f)
	) name12634 (
		_w15222_,
		_w15282_,
		_w23146_,
		_w23147_
	);
	LUT2 #(
		.INIT('h8)
	) name12635 (
		\wishbone_RxPointerMSB_reg[25]/NET0131 ,
		\wishbone_RxPointerMSB_reg[26]/NET0131 ,
		_w23148_
	);
	LUT4 #(
		.INIT('h8000)
	) name12636 (
		_w15288_,
		_w15291_,
		_w15293_,
		_w23148_,
		_w23149_
	);
	LUT4 #(
		.INIT('h8000)
	) name12637 (
		_w15288_,
		_w15291_,
		_w15293_,
		_w23142_,
		_w23150_
	);
	LUT4 #(
		.INIT('h70f0)
	) name12638 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxPointerMSB_reg[26]/NET0131 ,
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w23151_
	);
	LUT3 #(
		.INIT('h54)
	) name12639 (
		_w23149_,
		_w23150_,
		_w23151_,
		_w23152_
	);
	LUT3 #(
		.INIT('hf4)
	) name12640 (
		_w14872_,
		_w15282_,
		_w23152_,
		_w23153_
	);
	LUT3 #(
		.INIT('h80)
	) name12641 (
		\wishbone_RxPointerMSB_reg[25]/NET0131 ,
		\wishbone_RxPointerMSB_reg[26]/NET0131 ,
		\wishbone_RxPointerMSB_reg[27]/NET0131 ,
		_w23154_
	);
	LUT4 #(
		.INIT('h8000)
	) name12642 (
		_w15288_,
		_w15291_,
		_w15293_,
		_w23154_,
		_w23155_
	);
	LUT4 #(
		.INIT('h0032)
	) name12643 (
		\wishbone_RxPointerMSB_reg[27]/NET0131 ,
		_w13807_,
		_w23149_,
		_w23155_,
		_w23156_
	);
	LUT3 #(
		.INIT('hf2)
	) name12644 (
		_w15282_,
		_w17356_,
		_w23156_,
		_w23157_
	);
	LUT4 #(
		.INIT('h8000)
	) name12645 (
		\wishbone_RxPointerMSB_reg[25]/NET0131 ,
		\wishbone_RxPointerMSB_reg[26]/NET0131 ,
		\wishbone_RxPointerMSB_reg[27]/NET0131 ,
		\wishbone_RxPointerMSB_reg[28]/NET0131 ,
		_w23158_
	);
	LUT4 #(
		.INIT('h8000)
	) name12646 (
		_w15288_,
		_w15291_,
		_w15293_,
		_w23158_,
		_w23159_
	);
	LUT4 #(
		.INIT('h0032)
	) name12647 (
		\wishbone_RxPointerMSB_reg[28]/NET0131 ,
		_w13807_,
		_w23155_,
		_w23159_,
		_w23160_
	);
	LUT3 #(
		.INIT('hf4)
	) name12648 (
		_w12301_,
		_w15282_,
		_w23160_,
		_w23161_
	);
	LUT4 #(
		.INIT('h0302)
	) name12649 (
		\wishbone_RxPointerMSB_reg[29]/NET0131 ,
		_w13807_,
		_w15297_,
		_w23159_,
		_w23162_
	);
	LUT3 #(
		.INIT('hf4)
	) name12650 (
		_w12668_,
		_w15282_,
		_w23162_,
		_w23163_
	);
	LUT3 #(
		.INIT('h12)
	) name12651 (
		\wishbone_RxPointerMSB_reg[31]/NET0131 ,
		_w13807_,
		_w15300_,
		_w23164_
	);
	LUT4 #(
		.INIT('h5154)
	) name12652 (
		wb_rst_i_pad,
		\wishbone_RxPointerMSB_reg[31]/NET0131 ,
		_w13807_,
		_w15300_,
		_w23165_
	);
	LUT3 #(
		.INIT('hdc)
	) name12653 (
		_w16469_,
		_w23164_,
		_w23165_,
		_w23166_
	);
	LUT2 #(
		.INIT('h8)
	) name12654 (
		\wishbone_RxPointerMSB_reg[7]/NET0131 ,
		\wishbone_RxPointerMSB_reg[8]/NET0131 ,
		_w23167_
	);
	LUT4 #(
		.INIT('h1555)
	) name12655 (
		\wishbone_RxPointerMSB_reg[9]/NET0131 ,
		_w15283_,
		_w15284_,
		_w23167_,
		_w23168_
	);
	LUT3 #(
		.INIT('h80)
	) name12656 (
		\wishbone_RxPointerMSB_reg[7]/NET0131 ,
		\wishbone_RxPointerMSB_reg[8]/NET0131 ,
		\wishbone_RxPointerMSB_reg[9]/NET0131 ,
		_w23169_
	);
	LUT4 #(
		.INIT('h1555)
	) name12657 (
		_w13807_,
		_w15283_,
		_w15284_,
		_w23169_,
		_w23170_
	);
	LUT2 #(
		.INIT('h4)
	) name12658 (
		_w23168_,
		_w23170_,
		_w23171_
	);
	LUT3 #(
		.INIT('hf2)
	) name12659 (
		_w15282_,
		_w21841_,
		_w23171_,
		_w23172_
	);
	LUT2 #(
		.INIT('h8)
	) name12660 (
		\wishbone_TxPointerMSB_reg[18]/NET0131 ,
		\wishbone_TxPointerMSB_reg[19]/NET0131 ,
		_w23173_
	);
	LUT3 #(
		.INIT('h80)
	) name12661 (
		_w15310_,
		_w15314_,
		_w23173_,
		_w23174_
	);
	LUT4 #(
		.INIT('h70f0)
	) name12662 (
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		\wishbone_TxPointerMSB_reg[19]/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w23175_
	);
	LUT4 #(
		.INIT('h70f0)
	) name12663 (
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		\wishbone_TxPointerMSB_reg[18]/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w23176_
	);
	LUT4 #(
		.INIT('h070f)
	) name12664 (
		_w15310_,
		_w15314_,
		_w23175_,
		_w23176_,
		_w23177_
	);
	LUT2 #(
		.INIT('h1)
	) name12665 (
		_w23174_,
		_w23177_,
		_w23178_
	);
	LUT3 #(
		.INIT('hf4)
	) name12666 (
		_w17713_,
		_w19180_,
		_w23178_,
		_w23179_
	);
	LUT4 #(
		.INIT('h1555)
	) name12667 (
		\wishbone_TxPointerMSB_reg[20]/NET0131 ,
		_w15310_,
		_w15314_,
		_w23173_,
		_w23180_
	);
	LUT4 #(
		.INIT('h1555)
	) name12668 (
		_w15303_,
		_w15310_,
		_w15314_,
		_w15315_,
		_w23181_
	);
	LUT2 #(
		.INIT('h4)
	) name12669 (
		_w23180_,
		_w23181_,
		_w23182_
	);
	LUT3 #(
		.INIT('hf4)
	) name12670 (
		_w14512_,
		_w19180_,
		_w23182_,
		_w23183_
	);
	LUT4 #(
		.INIT('h1555)
	) name12671 (
		\wishbone_TxPointerMSB_reg[21]/NET0131 ,
		_w15310_,
		_w15314_,
		_w15315_,
		_w23184_
	);
	LUT4 #(
		.INIT('h8000)
	) name12672 (
		\wishbone_TxPointerMSB_reg[18]/NET0131 ,
		\wishbone_TxPointerMSB_reg[19]/NET0131 ,
		\wishbone_TxPointerMSB_reg[20]/NET0131 ,
		\wishbone_TxPointerMSB_reg[21]/NET0131 ,
		_w23185_
	);
	LUT4 #(
		.INIT('h1555)
	) name12673 (
		_w15303_,
		_w15310_,
		_w15314_,
		_w23185_,
		_w23186_
	);
	LUT2 #(
		.INIT('h4)
	) name12674 (
		_w23184_,
		_w23186_,
		_w23187_
	);
	LUT3 #(
		.INIT('hf4)
	) name12675 (
		_w18058_,
		_w19180_,
		_w23187_,
		_w23188_
	);
	LUT4 #(
		.INIT('h1555)
	) name12676 (
		\wishbone_TxPointerMSB_reg[22]/NET0131 ,
		_w15310_,
		_w15314_,
		_w23185_,
		_w23189_
	);
	LUT4 #(
		.INIT('h1555)
	) name12677 (
		_w15303_,
		_w15310_,
		_w15314_,
		_w15317_,
		_w23190_
	);
	LUT2 #(
		.INIT('h4)
	) name12678 (
		_w23189_,
		_w23190_,
		_w23191_
	);
	LUT3 #(
		.INIT('hf4)
	) name12679 (
		_w18746_,
		_w19180_,
		_w23191_,
		_w23192_
	);
	LUT4 #(
		.INIT('h70f0)
	) name12680 (
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		\wishbone_TxPointerMSB_reg[23]/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w23193_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12681 (
		_w15310_,
		_w15314_,
		_w15317_,
		_w23193_,
		_w23194_
	);
	LUT4 #(
		.INIT('h070f)
	) name12682 (
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		\wishbone_TxPointerMSB_reg[23]/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w23195_
	);
	LUT4 #(
		.INIT('h8000)
	) name12683 (
		_w15310_,
		_w15314_,
		_w15317_,
		_w23195_,
		_w23196_
	);
	LUT2 #(
		.INIT('h1)
	) name12684 (
		_w23194_,
		_w23196_,
		_w23197_
	);
	LUT3 #(
		.INIT('h4f)
	) name12685 (
		_w18401_,
		_w19180_,
		_w23197_,
		_w23198_
	);
	LUT4 #(
		.INIT('h060c)
	) name12686 (
		\wishbone_TxPointerMSB_reg[23]/NET0131 ,
		\wishbone_TxPointerMSB_reg[24]/NET0131 ,
		_w15303_,
		_w15318_,
		_w23199_
	);
	LUT3 #(
		.INIT('hf4)
	) name12687 (
		_w13397_,
		_w19180_,
		_w23199_,
		_w23200_
	);
	LUT3 #(
		.INIT('h80)
	) name12688 (
		\wishbone_TxPointerMSB_reg[23]/NET0131 ,
		\wishbone_TxPointerMSB_reg[24]/NET0131 ,
		\wishbone_TxPointerMSB_reg[25]/NET0131 ,
		_w23201_
	);
	LUT4 #(
		.INIT('h8000)
	) name12689 (
		_w15310_,
		_w15314_,
		_w15317_,
		_w23201_,
		_w23202_
	);
	LUT4 #(
		.INIT('h70f0)
	) name12690 (
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		\wishbone_TxPointerMSB_reg[25]/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w23203_
	);
	LUT2 #(
		.INIT('h4)
	) name12691 (
		_w15303_,
		_w15320_,
		_w23204_
	);
	LUT4 #(
		.INIT('h8000)
	) name12692 (
		_w15310_,
		_w15314_,
		_w15317_,
		_w23204_,
		_w23205_
	);
	LUT3 #(
		.INIT('h54)
	) name12693 (
		_w23202_,
		_w23203_,
		_w23205_,
		_w23206_
	);
	LUT3 #(
		.INIT('hf4)
	) name12694 (
		_w15222_,
		_w19180_,
		_w23206_,
		_w23207_
	);
	LUT4 #(
		.INIT('h8000)
	) name12695 (
		\wishbone_TxPointerMSB_reg[23]/NET0131 ,
		\wishbone_TxPointerMSB_reg[24]/NET0131 ,
		\wishbone_TxPointerMSB_reg[25]/NET0131 ,
		\wishbone_TxPointerMSB_reg[26]/NET0131 ,
		_w23208_
	);
	LUT4 #(
		.INIT('h8000)
	) name12696 (
		_w15310_,
		_w15314_,
		_w15317_,
		_w23208_,
		_w23209_
	);
	LUT4 #(
		.INIT('h0032)
	) name12697 (
		\wishbone_TxPointerMSB_reg[26]/NET0131 ,
		_w15303_,
		_w23202_,
		_w23209_,
		_w23210_
	);
	LUT3 #(
		.INIT('hf4)
	) name12698 (
		_w14872_,
		_w19180_,
		_w23210_,
		_w23211_
	);
	LUT3 #(
		.INIT('h80)
	) name12699 (
		\wishbone_TxPointerMSB_reg[23]/NET0131 ,
		\wishbone_TxPointerMSB_reg[24]/NET0131 ,
		\wishbone_TxPointerMSB_reg[27]/NET0131 ,
		_w23212_
	);
	LUT2 #(
		.INIT('h8)
	) name12700 (
		_w15319_,
		_w23212_,
		_w23213_
	);
	LUT4 #(
		.INIT('h8000)
	) name12701 (
		_w15310_,
		_w15314_,
		_w15317_,
		_w23213_,
		_w23214_
	);
	LUT4 #(
		.INIT('h0032)
	) name12702 (
		\wishbone_TxPointerMSB_reg[27]/NET0131 ,
		_w15303_,
		_w23209_,
		_w23214_,
		_w23215_
	);
	LUT3 #(
		.INIT('hf4)
	) name12703 (
		_w17356_,
		_w19180_,
		_w23215_,
		_w23216_
	);
	LUT3 #(
		.INIT('hed)
	) name12704 (
		\wishbone_TxPointerMSB_reg[29]/NET0131 ,
		_w15303_,
		_w15323_,
		_w23217_
	);
	LUT3 #(
		.INIT('h4f)
	) name12705 (
		_w12668_,
		_w19180_,
		_w23217_,
		_w23218_
	);
	LUT4 #(
		.INIT('h0302)
	) name12706 (
		\wishbone_TxPointerMSB_reg[28]/NET0131 ,
		_w15303_,
		_w15323_,
		_w23214_,
		_w23219_
	);
	LUT3 #(
		.INIT('hf4)
	) name12707 (
		_w12301_,
		_w19180_,
		_w23219_,
		_w23220_
	);
	LUT4 #(
		.INIT('h8000)
	) name12708 (
		\wishbone_TxPointerMSB_reg[27]/NET0131 ,
		\wishbone_TxPointerMSB_reg[28]/NET0131 ,
		\wishbone_TxPointerMSB_reg[29]/NET0131 ,
		\wishbone_TxPointerMSB_reg[30]/NET0131 ,
		_w23221_
	);
	LUT2 #(
		.INIT('h8)
	) name12709 (
		_w23208_,
		_w23221_,
		_w23222_
	);
	LUT4 #(
		.INIT('h8000)
	) name12710 (
		_w15310_,
		_w15314_,
		_w15317_,
		_w23222_,
		_w23223_
	);
	LUT3 #(
		.INIT('hed)
	) name12711 (
		\wishbone_TxPointerMSB_reg[31]/NET0131 ,
		_w15303_,
		_w23223_,
		_w23224_
	);
	LUT3 #(
		.INIT('h4f)
	) name12712 (
		_w16469_,
		_w19180_,
		_w23224_,
		_w23225_
	);
	LUT2 #(
		.INIT('h8)
	) name12713 (
		\wishbone_TxPointerMSB_reg[7]/NET0131 ,
		\wishbone_TxPointerMSB_reg[8]/NET0131 ,
		_w23226_
	);
	LUT4 #(
		.INIT('h1555)
	) name12714 (
		\wishbone_TxPointerMSB_reg[9]/NET0131 ,
		_w15305_,
		_w15306_,
		_w23226_,
		_w23227_
	);
	LUT4 #(
		.INIT('h1555)
	) name12715 (
		_w15303_,
		_w15305_,
		_w15306_,
		_w15307_,
		_w23228_
	);
	LUT2 #(
		.INIT('h4)
	) name12716 (
		_w23227_,
		_w23228_,
		_w23229_
	);
	LUT3 #(
		.INIT('hf2)
	) name12717 (
		_w19180_,
		_w21841_,
		_w23229_,
		_w23230_
	);
	LUT3 #(
		.INIT('h80)
	) name12718 (
		\ethreg1_MODER_1_DataOut_reg[5]/NET0131 ,
		_w18800_,
		_w18801_,
		_w23231_
	);
	LUT4 #(
		.INIT('h0020)
	) name12719 (
		\ethreg1_TXCTRL_1_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23232_
	);
	LUT3 #(
		.INIT('h80)
	) name12720 (
		_w18757_,
		_w18758_,
		_w23232_,
		_w23233_
	);
	LUT4 #(
		.INIT('h0008)
	) name12721 (
		\ethreg1_RXHASH0_1_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23234_
	);
	LUT3 #(
		.INIT('h80)
	) name12722 (
		_w18757_,
		_w18758_,
		_w23234_,
		_w23235_
	);
	LUT4 #(
		.INIT('h0008)
	) name12723 (
		\ethreg1_RXHASH1_1_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23236_
	);
	LUT3 #(
		.INIT('h80)
	) name12724 (
		_w18757_,
		_w18762_,
		_w23236_,
		_w23237_
	);
	LUT4 #(
		.INIT('h0001)
	) name12725 (
		_w23231_,
		_w23233_,
		_w23235_,
		_w23237_,
		_w23238_
	);
	LUT3 #(
		.INIT('h80)
	) name12726 (
		\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 ,
		_w18753_,
		_w18754_,
		_w23239_
	);
	LUT3 #(
		.INIT('h80)
	) name12727 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[5]/NET0131 ,
		_w18798_,
		_w18805_,
		_w23240_
	);
	LUT4 #(
		.INIT('h0002)
	) name12728 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23241_
	);
	LUT3 #(
		.INIT('h80)
	) name12729 (
		_w18757_,
		_w18758_,
		_w23241_,
		_w23242_
	);
	LUT4 #(
		.INIT('h0002)
	) name12730 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23243_
	);
	LUT3 #(
		.INIT('h80)
	) name12731 (
		_w18757_,
		_w18762_,
		_w23243_,
		_w23244_
	);
	LUT3 #(
		.INIT('h80)
	) name12732 (
		\ethreg1_MIIRX_DATA_DataOut_reg[13]/NET0131 ,
		_w18785_,
		_w18786_,
		_w23245_
	);
	LUT4 #(
		.INIT('h0001)
	) name12733 (
		_w23240_,
		_w23242_,
		_w23244_,
		_w23245_,
		_w23246_
	);
	LUT4 #(
		.INIT('h0800)
	) name12734 (
		_w18752_,
		_w23238_,
		_w23239_,
		_w23246_,
		_w23247_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name12735 (
		_w18752_,
		_w23238_,
		_w23239_,
		_w23246_,
		_w23248_
	);
	LUT3 #(
		.INIT('h80)
	) name12736 (
		\wishbone_bd_ram_mem1_reg[65][13]/P0001 ,
		_w11949_,
		_w11977_,
		_w23249_
	);
	LUT3 #(
		.INIT('h80)
	) name12737 (
		\wishbone_bd_ram_mem1_reg[126][13]/P0001 ,
		_w11948_,
		_w12012_,
		_w23250_
	);
	LUT3 #(
		.INIT('h80)
	) name12738 (
		\wishbone_bd_ram_mem1_reg[57][13]/P0001 ,
		_w11968_,
		_w11979_,
		_w23251_
	);
	LUT3 #(
		.INIT('h80)
	) name12739 (
		\wishbone_bd_ram_mem1_reg[82][13]/P0001 ,
		_w11963_,
		_w11972_,
		_w23252_
	);
	LUT4 #(
		.INIT('h0001)
	) name12740 (
		_w23249_,
		_w23250_,
		_w23251_,
		_w23252_,
		_w23253_
	);
	LUT3 #(
		.INIT('h80)
	) name12741 (
		\wishbone_bd_ram_mem1_reg[188][13]/P0001 ,
		_w11942_,
		_w11954_,
		_w23254_
	);
	LUT3 #(
		.INIT('h80)
	) name12742 (
		\wishbone_bd_ram_mem1_reg[134][13]/P0001 ,
		_w11955_,
		_w11986_,
		_w23255_
	);
	LUT3 #(
		.INIT('h80)
	) name12743 (
		\wishbone_bd_ram_mem1_reg[37][13]/P0001 ,
		_w11933_,
		_w11957_,
		_w23256_
	);
	LUT3 #(
		.INIT('h80)
	) name12744 (
		\wishbone_bd_ram_mem1_reg[203][13]/P0001 ,
		_w11936_,
		_w11945_,
		_w23257_
	);
	LUT4 #(
		.INIT('h0001)
	) name12745 (
		_w23254_,
		_w23255_,
		_w23256_,
		_w23257_,
		_w23258_
	);
	LUT3 #(
		.INIT('h80)
	) name12746 (
		\wishbone_bd_ram_mem1_reg[201][13]/P0001 ,
		_w11945_,
		_w11968_,
		_w23259_
	);
	LUT3 #(
		.INIT('h80)
	) name12747 (
		\wishbone_bd_ram_mem1_reg[209][13]/P0001 ,
		_w11977_,
		_w11984_,
		_w23260_
	);
	LUT3 #(
		.INIT('h80)
	) name12748 (
		\wishbone_bd_ram_mem1_reg[29][13]/P0001 ,
		_w11935_,
		_w11966_,
		_w23261_
	);
	LUT3 #(
		.INIT('h80)
	) name12749 (
		\wishbone_bd_ram_mem1_reg[36][13]/P0001 ,
		_w11929_,
		_w11957_,
		_w23262_
	);
	LUT4 #(
		.INIT('h0001)
	) name12750 (
		_w23259_,
		_w23260_,
		_w23261_,
		_w23262_,
		_w23263_
	);
	LUT3 #(
		.INIT('h80)
	) name12751 (
		\wishbone_bd_ram_mem1_reg[154][13]/P0001 ,
		_w11944_,
		_w11959_,
		_w23264_
	);
	LUT3 #(
		.INIT('h80)
	) name12752 (
		\wishbone_bd_ram_mem1_reg[233][13]/P0001 ,
		_w11968_,
		_w11982_,
		_w23265_
	);
	LUT3 #(
		.INIT('h80)
	) name12753 (
		\wishbone_bd_ram_mem1_reg[87][13]/P0001 ,
		_w11972_,
		_w11975_,
		_w23266_
	);
	LUT3 #(
		.INIT('h80)
	) name12754 (
		\wishbone_bd_ram_mem1_reg[179][13]/P0001 ,
		_w11938_,
		_w11942_,
		_w23267_
	);
	LUT4 #(
		.INIT('h0001)
	) name12755 (
		_w23264_,
		_w23265_,
		_w23266_,
		_w23267_,
		_w23268_
	);
	LUT4 #(
		.INIT('h8000)
	) name12756 (
		_w23253_,
		_w23258_,
		_w23263_,
		_w23268_,
		_w23269_
	);
	LUT3 #(
		.INIT('h80)
	) name12757 (
		\wishbone_bd_ram_mem1_reg[90][13]/P0001 ,
		_w11944_,
		_w11972_,
		_w23270_
	);
	LUT3 #(
		.INIT('h80)
	) name12758 (
		\wishbone_bd_ram_mem1_reg[255][13]/P0001 ,
		_w11952_,
		_w11973_,
		_w23271_
	);
	LUT3 #(
		.INIT('h80)
	) name12759 (
		\wishbone_bd_ram_mem1_reg[177][13]/P0001 ,
		_w11942_,
		_w11977_,
		_w23272_
	);
	LUT3 #(
		.INIT('h80)
	) name12760 (
		\wishbone_bd_ram_mem1_reg[213][13]/P0001 ,
		_w11933_,
		_w11984_,
		_w23273_
	);
	LUT4 #(
		.INIT('h0001)
	) name12761 (
		_w23270_,
		_w23271_,
		_w23272_,
		_w23273_,
		_w23274_
	);
	LUT3 #(
		.INIT('h80)
	) name12762 (
		\wishbone_bd_ram_mem1_reg[184][13]/P0001 ,
		_w11942_,
		_w11990_,
		_w23275_
	);
	LUT3 #(
		.INIT('h80)
	) name12763 (
		\wishbone_bd_ram_mem1_reg[47][13]/P0001 ,
		_w11957_,
		_w11973_,
		_w23276_
	);
	LUT3 #(
		.INIT('h80)
	) name12764 (
		\wishbone_bd_ram_mem1_reg[74][13]/P0001 ,
		_w11944_,
		_w11949_,
		_w23277_
	);
	LUT3 #(
		.INIT('h80)
	) name12765 (
		\wishbone_bd_ram_mem1_reg[84][13]/P0001 ,
		_w11929_,
		_w11972_,
		_w23278_
	);
	LUT4 #(
		.INIT('h0001)
	) name12766 (
		_w23275_,
		_w23276_,
		_w23277_,
		_w23278_,
		_w23279_
	);
	LUT3 #(
		.INIT('h80)
	) name12767 (
		\wishbone_bd_ram_mem1_reg[30][13]/P0001 ,
		_w11935_,
		_w11948_,
		_w23280_
	);
	LUT3 #(
		.INIT('h80)
	) name12768 (
		\wishbone_bd_ram_mem1_reg[54][13]/P0001 ,
		_w11979_,
		_w11986_,
		_w23281_
	);
	LUT3 #(
		.INIT('h80)
	) name12769 (
		\wishbone_bd_ram_mem1_reg[176][13]/P0001 ,
		_w11941_,
		_w11942_,
		_w23282_
	);
	LUT3 #(
		.INIT('h80)
	) name12770 (
		\wishbone_bd_ram_mem1_reg[175][13]/P0001 ,
		_w11930_,
		_w11973_,
		_w23283_
	);
	LUT4 #(
		.INIT('h0001)
	) name12771 (
		_w23280_,
		_w23281_,
		_w23282_,
		_w23283_,
		_w23284_
	);
	LUT3 #(
		.INIT('h80)
	) name12772 (
		\wishbone_bd_ram_mem1_reg[13][13]/P0001 ,
		_w11932_,
		_w11966_,
		_w23285_
	);
	LUT3 #(
		.INIT('h80)
	) name12773 (
		\wishbone_bd_ram_mem1_reg[143][13]/P0001 ,
		_w11955_,
		_w11973_,
		_w23286_
	);
	LUT3 #(
		.INIT('h80)
	) name12774 (
		\wishbone_bd_ram_mem1_reg[5][13]/P0001 ,
		_w11932_,
		_w11933_,
		_w23287_
	);
	LUT3 #(
		.INIT('h80)
	) name12775 (
		\wishbone_bd_ram_mem1_reg[217][13]/P0001 ,
		_w11968_,
		_w11984_,
		_w23288_
	);
	LUT4 #(
		.INIT('h0001)
	) name12776 (
		_w23285_,
		_w23286_,
		_w23287_,
		_w23288_,
		_w23289_
	);
	LUT4 #(
		.INIT('h8000)
	) name12777 (
		_w23274_,
		_w23279_,
		_w23284_,
		_w23289_,
		_w23290_
	);
	LUT3 #(
		.INIT('h80)
	) name12778 (
		\wishbone_bd_ram_mem1_reg[78][13]/P0001 ,
		_w11948_,
		_w11949_,
		_w23291_
	);
	LUT3 #(
		.INIT('h80)
	) name12779 (
		\wishbone_bd_ram_mem1_reg[137][13]/P0001 ,
		_w11955_,
		_w11968_,
		_w23292_
	);
	LUT3 #(
		.INIT('h80)
	) name12780 (
		\wishbone_bd_ram_mem1_reg[115][13]/P0001 ,
		_w11938_,
		_w12012_,
		_w23293_
	);
	LUT3 #(
		.INIT('h80)
	) name12781 (
		\wishbone_bd_ram_mem1_reg[80][13]/P0001 ,
		_w11941_,
		_w11972_,
		_w23294_
	);
	LUT4 #(
		.INIT('h0001)
	) name12782 (
		_w23291_,
		_w23292_,
		_w23293_,
		_w23294_,
		_w23295_
	);
	LUT3 #(
		.INIT('h80)
	) name12783 (
		\wishbone_bd_ram_mem1_reg[182][13]/P0001 ,
		_w11942_,
		_w11986_,
		_w23296_
	);
	LUT3 #(
		.INIT('h80)
	) name12784 (
		\wishbone_bd_ram_mem1_reg[199][13]/P0001 ,
		_w11945_,
		_w11975_,
		_w23297_
	);
	LUT3 #(
		.INIT('h80)
	) name12785 (
		\wishbone_bd_ram_mem1_reg[216][13]/P0001 ,
		_w11984_,
		_w11990_,
		_w23298_
	);
	LUT3 #(
		.INIT('h80)
	) name12786 (
		\wishbone_bd_ram_mem1_reg[146][13]/P0001 ,
		_w11959_,
		_w11963_,
		_w23299_
	);
	LUT4 #(
		.INIT('h0001)
	) name12787 (
		_w23296_,
		_w23297_,
		_w23298_,
		_w23299_,
		_w23300_
	);
	LUT3 #(
		.INIT('h80)
	) name12788 (
		\wishbone_bd_ram_mem1_reg[44][13]/P0001 ,
		_w11954_,
		_w11957_,
		_w23301_
	);
	LUT3 #(
		.INIT('h80)
	) name12789 (
		\wishbone_bd_ram_mem1_reg[219][13]/P0001 ,
		_w11936_,
		_w11984_,
		_w23302_
	);
	LUT3 #(
		.INIT('h80)
	) name12790 (
		\wishbone_bd_ram_mem1_reg[150][13]/P0001 ,
		_w11959_,
		_w11986_,
		_w23303_
	);
	LUT3 #(
		.INIT('h80)
	) name12791 (
		\wishbone_bd_ram_mem1_reg[194][13]/P0001 ,
		_w11945_,
		_w11963_,
		_w23304_
	);
	LUT4 #(
		.INIT('h0001)
	) name12792 (
		_w23301_,
		_w23302_,
		_w23303_,
		_w23304_,
		_w23305_
	);
	LUT3 #(
		.INIT('h80)
	) name12793 (
		\wishbone_bd_ram_mem1_reg[100][13]/P0001 ,
		_w11929_,
		_w11965_,
		_w23306_
	);
	LUT3 #(
		.INIT('h80)
	) name12794 (
		\wishbone_bd_ram_mem1_reg[229][13]/P0001 ,
		_w11933_,
		_w11982_,
		_w23307_
	);
	LUT3 #(
		.INIT('h80)
	) name12795 (
		\wishbone_bd_ram_mem1_reg[96][13]/P0001 ,
		_w11941_,
		_w11965_,
		_w23308_
	);
	LUT3 #(
		.INIT('h80)
	) name12796 (
		\wishbone_bd_ram_mem1_reg[252][13]/P0001 ,
		_w11952_,
		_w11954_,
		_w23309_
	);
	LUT4 #(
		.INIT('h0001)
	) name12797 (
		_w23306_,
		_w23307_,
		_w23308_,
		_w23309_,
		_w23310_
	);
	LUT4 #(
		.INIT('h8000)
	) name12798 (
		_w23295_,
		_w23300_,
		_w23305_,
		_w23310_,
		_w23311_
	);
	LUT3 #(
		.INIT('h80)
	) name12799 (
		\wishbone_bd_ram_mem1_reg[232][13]/P0001 ,
		_w11982_,
		_w11990_,
		_w23312_
	);
	LUT3 #(
		.INIT('h80)
	) name12800 (
		\wishbone_bd_ram_mem1_reg[56][13]/P0001 ,
		_w11979_,
		_w11990_,
		_w23313_
	);
	LUT3 #(
		.INIT('h80)
	) name12801 (
		\wishbone_bd_ram_mem1_reg[171][13]/P0001 ,
		_w11930_,
		_w11936_,
		_w23314_
	);
	LUT3 #(
		.INIT('h80)
	) name12802 (
		\wishbone_bd_ram_mem1_reg[38][13]/P0001 ,
		_w11957_,
		_w11986_,
		_w23315_
	);
	LUT4 #(
		.INIT('h0001)
	) name12803 (
		_w23312_,
		_w23313_,
		_w23314_,
		_w23315_,
		_w23316_
	);
	LUT3 #(
		.INIT('h80)
	) name12804 (
		\wishbone_bd_ram_mem1_reg[97][13]/P0001 ,
		_w11965_,
		_w11977_,
		_w23317_
	);
	LUT3 #(
		.INIT('h80)
	) name12805 (
		\wishbone_bd_ram_mem1_reg[95][13]/P0001 ,
		_w11972_,
		_w11973_,
		_w23318_
	);
	LUT3 #(
		.INIT('h80)
	) name12806 (
		\wishbone_bd_ram_mem1_reg[130][13]/P0001 ,
		_w11955_,
		_w11963_,
		_w23319_
	);
	LUT3 #(
		.INIT('h80)
	) name12807 (
		\wishbone_bd_ram_mem1_reg[107][13]/P0001 ,
		_w11936_,
		_w11965_,
		_w23320_
	);
	LUT4 #(
		.INIT('h0001)
	) name12808 (
		_w23317_,
		_w23318_,
		_w23319_,
		_w23320_,
		_w23321_
	);
	LUT3 #(
		.INIT('h80)
	) name12809 (
		\wishbone_bd_ram_mem1_reg[152][13]/P0001 ,
		_w11959_,
		_w11990_,
		_w23322_
	);
	LUT3 #(
		.INIT('h80)
	) name12810 (
		\wishbone_bd_ram_mem1_reg[145][13]/P0001 ,
		_w11959_,
		_w11977_,
		_w23323_
	);
	LUT3 #(
		.INIT('h80)
	) name12811 (
		\wishbone_bd_ram_mem1_reg[218][13]/P0001 ,
		_w11944_,
		_w11984_,
		_w23324_
	);
	LUT3 #(
		.INIT('h80)
	) name12812 (
		\wishbone_bd_ram_mem1_reg[141][13]/P0001 ,
		_w11955_,
		_w11966_,
		_w23325_
	);
	LUT4 #(
		.INIT('h0001)
	) name12813 (
		_w23322_,
		_w23323_,
		_w23324_,
		_w23325_,
		_w23326_
	);
	LUT3 #(
		.INIT('h80)
	) name12814 (
		\wishbone_bd_ram_mem1_reg[136][13]/P0001 ,
		_w11955_,
		_w11990_,
		_w23327_
	);
	LUT3 #(
		.INIT('h80)
	) name12815 (
		\wishbone_bd_ram_mem1_reg[6][13]/P0001 ,
		_w11932_,
		_w11986_,
		_w23328_
	);
	LUT3 #(
		.INIT('h80)
	) name12816 (
		\wishbone_bd_ram_mem1_reg[180][13]/P0001 ,
		_w11929_,
		_w11942_,
		_w23329_
	);
	LUT3 #(
		.INIT('h80)
	) name12817 (
		\wishbone_bd_ram_mem1_reg[166][13]/P0001 ,
		_w11930_,
		_w11986_,
		_w23330_
	);
	LUT4 #(
		.INIT('h0001)
	) name12818 (
		_w23327_,
		_w23328_,
		_w23329_,
		_w23330_,
		_w23331_
	);
	LUT4 #(
		.INIT('h8000)
	) name12819 (
		_w23316_,
		_w23321_,
		_w23326_,
		_w23331_,
		_w23332_
	);
	LUT4 #(
		.INIT('h8000)
	) name12820 (
		_w23269_,
		_w23290_,
		_w23311_,
		_w23332_,
		_w23333_
	);
	LUT3 #(
		.INIT('h80)
	) name12821 (
		\wishbone_bd_ram_mem1_reg[18][13]/P0001 ,
		_w11935_,
		_w11963_,
		_w23334_
	);
	LUT3 #(
		.INIT('h80)
	) name12822 (
		\wishbone_bd_ram_mem1_reg[76][13]/P0001 ,
		_w11949_,
		_w11954_,
		_w23335_
	);
	LUT3 #(
		.INIT('h80)
	) name12823 (
		\wishbone_bd_ram_mem1_reg[224][13]/P0001 ,
		_w11941_,
		_w11982_,
		_w23336_
	);
	LUT3 #(
		.INIT('h80)
	) name12824 (
		\wishbone_bd_ram_mem1_reg[27][13]/P0001 ,
		_w11935_,
		_w11936_,
		_w23337_
	);
	LUT4 #(
		.INIT('h0001)
	) name12825 (
		_w23334_,
		_w23335_,
		_w23336_,
		_w23337_,
		_w23338_
	);
	LUT3 #(
		.INIT('h80)
	) name12826 (
		\wishbone_bd_ram_mem1_reg[102][13]/P0001 ,
		_w11965_,
		_w11986_,
		_w23339_
	);
	LUT3 #(
		.INIT('h80)
	) name12827 (
		\wishbone_bd_ram_mem1_reg[75][13]/P0001 ,
		_w11936_,
		_w11949_,
		_w23340_
	);
	LUT3 #(
		.INIT('h80)
	) name12828 (
		\wishbone_bd_ram_mem1_reg[8][13]/P0001 ,
		_w11932_,
		_w11990_,
		_w23341_
	);
	LUT3 #(
		.INIT('h80)
	) name12829 (
		\wishbone_bd_ram_mem1_reg[21][13]/P0001 ,
		_w11933_,
		_w11935_,
		_w23342_
	);
	LUT4 #(
		.INIT('h0001)
	) name12830 (
		_w23339_,
		_w23340_,
		_w23341_,
		_w23342_,
		_w23343_
	);
	LUT3 #(
		.INIT('h80)
	) name12831 (
		\wishbone_bd_ram_mem1_reg[45][13]/P0001 ,
		_w11957_,
		_w11966_,
		_w23344_
	);
	LUT3 #(
		.INIT('h80)
	) name12832 (
		\wishbone_bd_ram_mem1_reg[110][13]/P0001 ,
		_w11948_,
		_w11965_,
		_w23345_
	);
	LUT3 #(
		.INIT('h80)
	) name12833 (
		\wishbone_bd_ram_mem1_reg[66][13]/P0001 ,
		_w11949_,
		_w11963_,
		_w23346_
	);
	LUT3 #(
		.INIT('h80)
	) name12834 (
		\wishbone_bd_ram_mem1_reg[170][13]/P0001 ,
		_w11930_,
		_w11944_,
		_w23347_
	);
	LUT4 #(
		.INIT('h0001)
	) name12835 (
		_w23344_,
		_w23345_,
		_w23346_,
		_w23347_,
		_w23348_
	);
	LUT3 #(
		.INIT('h80)
	) name12836 (
		\wishbone_bd_ram_mem1_reg[208][13]/P0001 ,
		_w11941_,
		_w11984_,
		_w23349_
	);
	LUT3 #(
		.INIT('h80)
	) name12837 (
		\wishbone_bd_ram_mem1_reg[79][13]/P0001 ,
		_w11949_,
		_w11973_,
		_w23350_
	);
	LUT3 #(
		.INIT('h80)
	) name12838 (
		\wishbone_bd_ram_mem1_reg[60][13]/P0001 ,
		_w11954_,
		_w11979_,
		_w23351_
	);
	LUT3 #(
		.INIT('h80)
	) name12839 (
		\wishbone_bd_ram_mem1_reg[214][13]/P0001 ,
		_w11984_,
		_w11986_,
		_w23352_
	);
	LUT4 #(
		.INIT('h0001)
	) name12840 (
		_w23349_,
		_w23350_,
		_w23351_,
		_w23352_,
		_w23353_
	);
	LUT4 #(
		.INIT('h8000)
	) name12841 (
		_w23338_,
		_w23343_,
		_w23348_,
		_w23353_,
		_w23354_
	);
	LUT3 #(
		.INIT('h80)
	) name12842 (
		\wishbone_bd_ram_mem1_reg[34][13]/P0001 ,
		_w11957_,
		_w11963_,
		_w23355_
	);
	LUT3 #(
		.INIT('h80)
	) name12843 (
		\wishbone_bd_ram_mem1_reg[247][13]/P0001 ,
		_w11952_,
		_w11975_,
		_w23356_
	);
	LUT3 #(
		.INIT('h80)
	) name12844 (
		\wishbone_bd_ram_mem1_reg[131][13]/P0001 ,
		_w11938_,
		_w11955_,
		_w23357_
	);
	LUT3 #(
		.INIT('h80)
	) name12845 (
		\wishbone_bd_ram_mem1_reg[158][13]/P0001 ,
		_w11948_,
		_w11959_,
		_w23358_
	);
	LUT4 #(
		.INIT('h0001)
	) name12846 (
		_w23355_,
		_w23356_,
		_w23357_,
		_w23358_,
		_w23359_
	);
	LUT3 #(
		.INIT('h80)
	) name12847 (
		\wishbone_bd_ram_mem1_reg[85][13]/P0001 ,
		_w11933_,
		_w11972_,
		_w23360_
	);
	LUT3 #(
		.INIT('h80)
	) name12848 (
		\wishbone_bd_ram_mem1_reg[103][13]/P0001 ,
		_w11965_,
		_w11975_,
		_w23361_
	);
	LUT3 #(
		.INIT('h80)
	) name12849 (
		\wishbone_bd_ram_mem1_reg[114][13]/P0001 ,
		_w11963_,
		_w12012_,
		_w23362_
	);
	LUT3 #(
		.INIT('h80)
	) name12850 (
		\wishbone_bd_ram_mem1_reg[52][13]/P0001 ,
		_w11929_,
		_w11979_,
		_w23363_
	);
	LUT4 #(
		.INIT('h0001)
	) name12851 (
		_w23360_,
		_w23361_,
		_w23362_,
		_w23363_,
		_w23364_
	);
	LUT3 #(
		.INIT('h80)
	) name12852 (
		\wishbone_bd_ram_mem1_reg[24][13]/P0001 ,
		_w11935_,
		_w11990_,
		_w23365_
	);
	LUT3 #(
		.INIT('h80)
	) name12853 (
		\wishbone_bd_ram_mem1_reg[138][13]/P0001 ,
		_w11944_,
		_w11955_,
		_w23366_
	);
	LUT3 #(
		.INIT('h80)
	) name12854 (
		\wishbone_bd_ram_mem1_reg[40][13]/P0001 ,
		_w11957_,
		_w11990_,
		_w23367_
	);
	LUT3 #(
		.INIT('h80)
	) name12855 (
		\wishbone_bd_ram_mem1_reg[31][13]/P0001 ,
		_w11935_,
		_w11973_,
		_w23368_
	);
	LUT4 #(
		.INIT('h0001)
	) name12856 (
		_w23365_,
		_w23366_,
		_w23367_,
		_w23368_,
		_w23369_
	);
	LUT3 #(
		.INIT('h80)
	) name12857 (
		\wishbone_bd_ram_mem1_reg[77][13]/P0001 ,
		_w11949_,
		_w11966_,
		_w23370_
	);
	LUT3 #(
		.INIT('h80)
	) name12858 (
		\wishbone_bd_ram_mem1_reg[239][13]/P0001 ,
		_w11973_,
		_w11982_,
		_w23371_
	);
	LUT3 #(
		.INIT('h80)
	) name12859 (
		\wishbone_bd_ram_mem1_reg[42][13]/P0001 ,
		_w11944_,
		_w11957_,
		_w23372_
	);
	LUT3 #(
		.INIT('h80)
	) name12860 (
		\wishbone_bd_ram_mem1_reg[155][13]/P0001 ,
		_w11936_,
		_w11959_,
		_w23373_
	);
	LUT4 #(
		.INIT('h0001)
	) name12861 (
		_w23370_,
		_w23371_,
		_w23372_,
		_w23373_,
		_w23374_
	);
	LUT4 #(
		.INIT('h8000)
	) name12862 (
		_w23359_,
		_w23364_,
		_w23369_,
		_w23374_,
		_w23375_
	);
	LUT3 #(
		.INIT('h80)
	) name12863 (
		\wishbone_bd_ram_mem1_reg[178][13]/P0001 ,
		_w11942_,
		_w11963_,
		_w23376_
	);
	LUT3 #(
		.INIT('h80)
	) name12864 (
		\wishbone_bd_ram_mem1_reg[92][13]/P0001 ,
		_w11954_,
		_w11972_,
		_w23377_
	);
	LUT3 #(
		.INIT('h80)
	) name12865 (
		\wishbone_bd_ram_mem1_reg[69][13]/P0001 ,
		_w11933_,
		_w11949_,
		_w23378_
	);
	LUT3 #(
		.INIT('h80)
	) name12866 (
		\wishbone_bd_ram_mem1_reg[191][13]/P0001 ,
		_w11942_,
		_w11973_,
		_w23379_
	);
	LUT4 #(
		.INIT('h0001)
	) name12867 (
		_w23376_,
		_w23377_,
		_w23378_,
		_w23379_,
		_w23380_
	);
	LUT3 #(
		.INIT('h80)
	) name12868 (
		\wishbone_bd_ram_mem1_reg[88][13]/P0001 ,
		_w11972_,
		_w11990_,
		_w23381_
	);
	LUT3 #(
		.INIT('h80)
	) name12869 (
		\wishbone_bd_ram_mem1_reg[109][13]/P0001 ,
		_w11965_,
		_w11966_,
		_w23382_
	);
	LUT3 #(
		.INIT('h80)
	) name12870 (
		\wishbone_bd_ram_mem1_reg[50][13]/P0001 ,
		_w11963_,
		_w11979_,
		_w23383_
	);
	LUT3 #(
		.INIT('h80)
	) name12871 (
		\wishbone_bd_ram_mem1_reg[118][13]/P0001 ,
		_w11986_,
		_w12012_,
		_w23384_
	);
	LUT4 #(
		.INIT('h0001)
	) name12872 (
		_w23381_,
		_w23382_,
		_w23383_,
		_w23384_,
		_w23385_
	);
	LUT3 #(
		.INIT('h80)
	) name12873 (
		\wishbone_bd_ram_mem1_reg[7][13]/P0001 ,
		_w11932_,
		_w11975_,
		_w23386_
	);
	LUT3 #(
		.INIT('h80)
	) name12874 (
		\wishbone_bd_ram_mem1_reg[12][13]/P0001 ,
		_w11932_,
		_w11954_,
		_w23387_
	);
	LUT3 #(
		.INIT('h80)
	) name12875 (
		\wishbone_bd_ram_mem1_reg[169][13]/P0001 ,
		_w11930_,
		_w11968_,
		_w23388_
	);
	LUT3 #(
		.INIT('h80)
	) name12876 (
		\wishbone_bd_ram_mem1_reg[49][13]/P0001 ,
		_w11977_,
		_w11979_,
		_w23389_
	);
	LUT4 #(
		.INIT('h0001)
	) name12877 (
		_w23386_,
		_w23387_,
		_w23388_,
		_w23389_,
		_w23390_
	);
	LUT3 #(
		.INIT('h80)
	) name12878 (
		\wishbone_bd_ram_mem1_reg[120][13]/P0001 ,
		_w11990_,
		_w12012_,
		_w23391_
	);
	LUT3 #(
		.INIT('h80)
	) name12879 (
		\wishbone_bd_ram_mem1_reg[237][13]/P0001 ,
		_w11966_,
		_w11982_,
		_w23392_
	);
	LUT3 #(
		.INIT('h80)
	) name12880 (
		\wishbone_bd_ram_mem1_reg[116][13]/P0001 ,
		_w11929_,
		_w12012_,
		_w23393_
	);
	LUT3 #(
		.INIT('h80)
	) name12881 (
		\wishbone_bd_ram_mem1_reg[122][13]/P0001 ,
		_w11944_,
		_w12012_,
		_w23394_
	);
	LUT4 #(
		.INIT('h0001)
	) name12882 (
		_w23391_,
		_w23392_,
		_w23393_,
		_w23394_,
		_w23395_
	);
	LUT4 #(
		.INIT('h8000)
	) name12883 (
		_w23380_,
		_w23385_,
		_w23390_,
		_w23395_,
		_w23396_
	);
	LUT3 #(
		.INIT('h80)
	) name12884 (
		\wishbone_bd_ram_mem1_reg[160][13]/P0001 ,
		_w11930_,
		_w11941_,
		_w23397_
	);
	LUT3 #(
		.INIT('h80)
	) name12885 (
		\wishbone_bd_ram_mem1_reg[167][13]/P0001 ,
		_w11930_,
		_w11975_,
		_w23398_
	);
	LUT3 #(
		.INIT('h80)
	) name12886 (
		\wishbone_bd_ram_mem1_reg[250][13]/P0001 ,
		_w11944_,
		_w11952_,
		_w23399_
	);
	LUT3 #(
		.INIT('h80)
	) name12887 (
		\wishbone_bd_ram_mem1_reg[240][13]/P0001 ,
		_w11941_,
		_w11952_,
		_w23400_
	);
	LUT4 #(
		.INIT('h0001)
	) name12888 (
		_w23397_,
		_w23398_,
		_w23399_,
		_w23400_,
		_w23401_
	);
	LUT3 #(
		.INIT('h80)
	) name12889 (
		\wishbone_bd_ram_mem1_reg[133][13]/P0001 ,
		_w11933_,
		_w11955_,
		_w23402_
	);
	LUT3 #(
		.INIT('h80)
	) name12890 (
		\wishbone_bd_ram_mem1_reg[111][13]/P0001 ,
		_w11965_,
		_w11973_,
		_w23403_
	);
	LUT3 #(
		.INIT('h80)
	) name12891 (
		\wishbone_bd_ram_mem1_reg[206][13]/P0001 ,
		_w11945_,
		_w11948_,
		_w23404_
	);
	LUT3 #(
		.INIT('h80)
	) name12892 (
		\wishbone_bd_ram_mem1_reg[112][13]/P0001 ,
		_w11941_,
		_w12012_,
		_w23405_
	);
	LUT4 #(
		.INIT('h0001)
	) name12893 (
		_w23402_,
		_w23403_,
		_w23404_,
		_w23405_,
		_w23406_
	);
	LUT3 #(
		.INIT('h80)
	) name12894 (
		\wishbone_bd_ram_mem1_reg[200][13]/P0001 ,
		_w11945_,
		_w11990_,
		_w23407_
	);
	LUT3 #(
		.INIT('h80)
	) name12895 (
		\wishbone_bd_ram_mem1_reg[91][13]/P0001 ,
		_w11936_,
		_w11972_,
		_w23408_
	);
	LUT3 #(
		.INIT('h80)
	) name12896 (
		\wishbone_bd_ram_mem1_reg[101][13]/P0001 ,
		_w11933_,
		_w11965_,
		_w23409_
	);
	LUT3 #(
		.INIT('h80)
	) name12897 (
		\wishbone_bd_ram_mem1_reg[132][13]/P0001 ,
		_w11929_,
		_w11955_,
		_w23410_
	);
	LUT4 #(
		.INIT('h0001)
	) name12898 (
		_w23407_,
		_w23408_,
		_w23409_,
		_w23410_,
		_w23411_
	);
	LUT3 #(
		.INIT('h80)
	) name12899 (
		\wishbone_bd_ram_mem1_reg[220][13]/P0001 ,
		_w11954_,
		_w11984_,
		_w23412_
	);
	LUT3 #(
		.INIT('h80)
	) name12900 (
		\wishbone_bd_ram_mem1_reg[251][13]/P0001 ,
		_w11936_,
		_w11952_,
		_w23413_
	);
	LUT3 #(
		.INIT('h80)
	) name12901 (
		\wishbone_bd_ram_mem1_reg[148][13]/P0001 ,
		_w11929_,
		_w11959_,
		_w23414_
	);
	LUT3 #(
		.INIT('h80)
	) name12902 (
		\wishbone_bd_ram_mem1_reg[108][13]/P0001 ,
		_w11954_,
		_w11965_,
		_w23415_
	);
	LUT4 #(
		.INIT('h0001)
	) name12903 (
		_w23412_,
		_w23413_,
		_w23414_,
		_w23415_,
		_w23416_
	);
	LUT4 #(
		.INIT('h8000)
	) name12904 (
		_w23401_,
		_w23406_,
		_w23411_,
		_w23416_,
		_w23417_
	);
	LUT4 #(
		.INIT('h8000)
	) name12905 (
		_w23354_,
		_w23375_,
		_w23396_,
		_w23417_,
		_w23418_
	);
	LUT3 #(
		.INIT('h80)
	) name12906 (
		\wishbone_bd_ram_mem1_reg[153][13]/P0001 ,
		_w11959_,
		_w11968_,
		_w23419_
	);
	LUT3 #(
		.INIT('h80)
	) name12907 (
		\wishbone_bd_ram_mem1_reg[127][13]/P0001 ,
		_w11973_,
		_w12012_,
		_w23420_
	);
	LUT3 #(
		.INIT('h80)
	) name12908 (
		\wishbone_bd_ram_mem1_reg[55][13]/P0001 ,
		_w11975_,
		_w11979_,
		_w23421_
	);
	LUT3 #(
		.INIT('h80)
	) name12909 (
		\wishbone_bd_ram_mem1_reg[53][13]/P0001 ,
		_w11933_,
		_w11979_,
		_w23422_
	);
	LUT4 #(
		.INIT('h0001)
	) name12910 (
		_w23419_,
		_w23420_,
		_w23421_,
		_w23422_,
		_w23423_
	);
	LUT3 #(
		.INIT('h80)
	) name12911 (
		\wishbone_bd_ram_mem1_reg[68][13]/P0001 ,
		_w11929_,
		_w11949_,
		_w23424_
	);
	LUT3 #(
		.INIT('h80)
	) name12912 (
		\wishbone_bd_ram_mem1_reg[17][13]/P0001 ,
		_w11935_,
		_w11977_,
		_w23425_
	);
	LUT3 #(
		.INIT('h80)
	) name12913 (
		\wishbone_bd_ram_mem1_reg[249][13]/P0001 ,
		_w11952_,
		_w11968_,
		_w23426_
	);
	LUT3 #(
		.INIT('h80)
	) name12914 (
		\wishbone_bd_ram_mem1_reg[19][13]/P0001 ,
		_w11935_,
		_w11938_,
		_w23427_
	);
	LUT4 #(
		.INIT('h0001)
	) name12915 (
		_w23424_,
		_w23425_,
		_w23426_,
		_w23427_,
		_w23428_
	);
	LUT3 #(
		.INIT('h80)
	) name12916 (
		\wishbone_bd_ram_mem1_reg[161][13]/P0001 ,
		_w11930_,
		_w11977_,
		_w23429_
	);
	LUT3 #(
		.INIT('h80)
	) name12917 (
		\wishbone_bd_ram_mem1_reg[20][13]/P0001 ,
		_w11929_,
		_w11935_,
		_w23430_
	);
	LUT3 #(
		.INIT('h80)
	) name12918 (
		\wishbone_bd_ram_mem1_reg[86][13]/P0001 ,
		_w11972_,
		_w11986_,
		_w23431_
	);
	LUT3 #(
		.INIT('h80)
	) name12919 (
		\wishbone_bd_ram_mem1_reg[227][13]/P0001 ,
		_w11938_,
		_w11982_,
		_w23432_
	);
	LUT4 #(
		.INIT('h0001)
	) name12920 (
		_w23429_,
		_w23430_,
		_w23431_,
		_w23432_,
		_w23433_
	);
	LUT3 #(
		.INIT('h80)
	) name12921 (
		\wishbone_bd_ram_mem1_reg[104][13]/P0001 ,
		_w11965_,
		_w11990_,
		_w23434_
	);
	LUT3 #(
		.INIT('h80)
	) name12922 (
		\wishbone_bd_ram_mem1_reg[62][13]/P0001 ,
		_w11948_,
		_w11979_,
		_w23435_
	);
	LUT3 #(
		.INIT('h80)
	) name12923 (
		\wishbone_bd_ram_mem1_reg[41][13]/P0001 ,
		_w11957_,
		_w11968_,
		_w23436_
	);
	LUT3 #(
		.INIT('h80)
	) name12924 (
		\wishbone_bd_ram_mem1_reg[117][13]/P0001 ,
		_w11933_,
		_w12012_,
		_w23437_
	);
	LUT4 #(
		.INIT('h0001)
	) name12925 (
		_w23434_,
		_w23435_,
		_w23436_,
		_w23437_,
		_w23438_
	);
	LUT4 #(
		.INIT('h8000)
	) name12926 (
		_w23423_,
		_w23428_,
		_w23433_,
		_w23438_,
		_w23439_
	);
	LUT3 #(
		.INIT('h80)
	) name12927 (
		\wishbone_bd_ram_mem1_reg[172][13]/P0001 ,
		_w11930_,
		_w11954_,
		_w23440_
	);
	LUT3 #(
		.INIT('h80)
	) name12928 (
		\wishbone_bd_ram_mem1_reg[26][13]/P0001 ,
		_w11935_,
		_w11944_,
		_w23441_
	);
	LUT3 #(
		.INIT('h80)
	) name12929 (
		\wishbone_bd_ram_mem1_reg[164][13]/P0001 ,
		_w11929_,
		_w11930_,
		_w23442_
	);
	LUT3 #(
		.INIT('h80)
	) name12930 (
		\wishbone_bd_ram_mem1_reg[3][13]/P0001 ,
		_w11932_,
		_w11938_,
		_w23443_
	);
	LUT4 #(
		.INIT('h0001)
	) name12931 (
		_w23440_,
		_w23441_,
		_w23442_,
		_w23443_,
		_w23444_
	);
	LUT3 #(
		.INIT('h80)
	) name12932 (
		\wishbone_bd_ram_mem1_reg[187][13]/P0001 ,
		_w11936_,
		_w11942_,
		_w23445_
	);
	LUT3 #(
		.INIT('h80)
	) name12933 (
		\wishbone_bd_ram_mem1_reg[10][13]/P0001 ,
		_w11932_,
		_w11944_,
		_w23446_
	);
	LUT3 #(
		.INIT('h80)
	) name12934 (
		\wishbone_bd_ram_mem1_reg[94][13]/P0001 ,
		_w11948_,
		_w11972_,
		_w23447_
	);
	LUT3 #(
		.INIT('h80)
	) name12935 (
		\wishbone_bd_ram_mem1_reg[234][13]/P0001 ,
		_w11944_,
		_w11982_,
		_w23448_
	);
	LUT4 #(
		.INIT('h0001)
	) name12936 (
		_w23445_,
		_w23446_,
		_w23447_,
		_w23448_,
		_w23449_
	);
	LUT3 #(
		.INIT('h80)
	) name12937 (
		\wishbone_bd_ram_mem1_reg[39][13]/P0001 ,
		_w11957_,
		_w11975_,
		_w23450_
	);
	LUT3 #(
		.INIT('h80)
	) name12938 (
		\wishbone_bd_ram_mem1_reg[113][13]/P0001 ,
		_w11977_,
		_w12012_,
		_w23451_
	);
	LUT3 #(
		.INIT('h80)
	) name12939 (
		\wishbone_bd_ram_mem1_reg[168][13]/P0001 ,
		_w11930_,
		_w11990_,
		_w23452_
	);
	LUT3 #(
		.INIT('h80)
	) name12940 (
		\wishbone_bd_ram_mem1_reg[22][13]/P0001 ,
		_w11935_,
		_w11986_,
		_w23453_
	);
	LUT4 #(
		.INIT('h0001)
	) name12941 (
		_w23450_,
		_w23451_,
		_w23452_,
		_w23453_,
		_w23454_
	);
	LUT3 #(
		.INIT('h80)
	) name12942 (
		\wishbone_bd_ram_mem1_reg[195][13]/P0001 ,
		_w11938_,
		_w11945_,
		_w23455_
	);
	LUT3 #(
		.INIT('h80)
	) name12943 (
		\wishbone_bd_ram_mem1_reg[70][13]/P0001 ,
		_w11949_,
		_w11986_,
		_w23456_
	);
	LUT3 #(
		.INIT('h80)
	) name12944 (
		\wishbone_bd_ram_mem1_reg[165][13]/P0001 ,
		_w11930_,
		_w11933_,
		_w23457_
	);
	LUT3 #(
		.INIT('h80)
	) name12945 (
		\wishbone_bd_ram_mem1_reg[71][13]/P0001 ,
		_w11949_,
		_w11975_,
		_w23458_
	);
	LUT4 #(
		.INIT('h0001)
	) name12946 (
		_w23455_,
		_w23456_,
		_w23457_,
		_w23458_,
		_w23459_
	);
	LUT4 #(
		.INIT('h8000)
	) name12947 (
		_w23444_,
		_w23449_,
		_w23454_,
		_w23459_,
		_w23460_
	);
	LUT3 #(
		.INIT('h80)
	) name12948 (
		\wishbone_bd_ram_mem1_reg[81][13]/P0001 ,
		_w11972_,
		_w11977_,
		_w23461_
	);
	LUT3 #(
		.INIT('h80)
	) name12949 (
		\wishbone_bd_ram_mem1_reg[253][13]/P0001 ,
		_w11952_,
		_w11966_,
		_w23462_
	);
	LUT3 #(
		.INIT('h80)
	) name12950 (
		\wishbone_bd_ram_mem1_reg[197][13]/P0001 ,
		_w11933_,
		_w11945_,
		_w23463_
	);
	LUT3 #(
		.INIT('h80)
	) name12951 (
		\wishbone_bd_ram_mem1_reg[174][13]/P0001 ,
		_w11930_,
		_w11948_,
		_w23464_
	);
	LUT4 #(
		.INIT('h0001)
	) name12952 (
		_w23461_,
		_w23462_,
		_w23463_,
		_w23464_,
		_w23465_
	);
	LUT3 #(
		.INIT('h80)
	) name12953 (
		\wishbone_bd_ram_mem1_reg[93][13]/P0001 ,
		_w11966_,
		_w11972_,
		_w23466_
	);
	LUT3 #(
		.INIT('h80)
	) name12954 (
		\wishbone_bd_ram_mem1_reg[125][13]/P0001 ,
		_w11966_,
		_w12012_,
		_w23467_
	);
	LUT3 #(
		.INIT('h80)
	) name12955 (
		\wishbone_bd_ram_mem1_reg[63][13]/P0001 ,
		_w11973_,
		_w11979_,
		_w23468_
	);
	LUT3 #(
		.INIT('h80)
	) name12956 (
		\wishbone_bd_ram_mem1_reg[246][13]/P0001 ,
		_w11952_,
		_w11986_,
		_w23469_
	);
	LUT4 #(
		.INIT('h0001)
	) name12957 (
		_w23466_,
		_w23467_,
		_w23468_,
		_w23469_,
		_w23470_
	);
	LUT3 #(
		.INIT('h80)
	) name12958 (
		\wishbone_bd_ram_mem1_reg[135][13]/P0001 ,
		_w11955_,
		_w11975_,
		_w23471_
	);
	LUT3 #(
		.INIT('h80)
	) name12959 (
		\wishbone_bd_ram_mem1_reg[59][13]/P0001 ,
		_w11936_,
		_w11979_,
		_w23472_
	);
	LUT3 #(
		.INIT('h80)
	) name12960 (
		\wishbone_bd_ram_mem1_reg[61][13]/P0001 ,
		_w11966_,
		_w11979_,
		_w23473_
	);
	LUT3 #(
		.INIT('h80)
	) name12961 (
		\wishbone_bd_ram_mem1_reg[235][13]/P0001 ,
		_w11936_,
		_w11982_,
		_w23474_
	);
	LUT4 #(
		.INIT('h0001)
	) name12962 (
		_w23471_,
		_w23472_,
		_w23473_,
		_w23474_,
		_w23475_
	);
	LUT3 #(
		.INIT('h80)
	) name12963 (
		\wishbone_bd_ram_mem1_reg[149][13]/P0001 ,
		_w11933_,
		_w11959_,
		_w23476_
	);
	LUT3 #(
		.INIT('h80)
	) name12964 (
		\wishbone_bd_ram_mem1_reg[222][13]/P0001 ,
		_w11948_,
		_w11984_,
		_w23477_
	);
	LUT3 #(
		.INIT('h80)
	) name12965 (
		\wishbone_bd_ram_mem1_reg[99][13]/P0001 ,
		_w11938_,
		_w11965_,
		_w23478_
	);
	LUT3 #(
		.INIT('h80)
	) name12966 (
		\wishbone_bd_ram_mem1_reg[248][13]/P0001 ,
		_w11952_,
		_w11990_,
		_w23479_
	);
	LUT4 #(
		.INIT('h0001)
	) name12967 (
		_w23476_,
		_w23477_,
		_w23478_,
		_w23479_,
		_w23480_
	);
	LUT4 #(
		.INIT('h8000)
	) name12968 (
		_w23465_,
		_w23470_,
		_w23475_,
		_w23480_,
		_w23481_
	);
	LUT3 #(
		.INIT('h80)
	) name12969 (
		\wishbone_bd_ram_mem1_reg[211][13]/P0001 ,
		_w11938_,
		_w11984_,
		_w23482_
	);
	LUT3 #(
		.INIT('h80)
	) name12970 (
		\wishbone_bd_ram_mem1_reg[156][13]/P0001 ,
		_w11954_,
		_w11959_,
		_w23483_
	);
	LUT3 #(
		.INIT('h80)
	) name12971 (
		\wishbone_bd_ram_mem1_reg[142][13]/P0001 ,
		_w11948_,
		_w11955_,
		_w23484_
	);
	LUT3 #(
		.INIT('h80)
	) name12972 (
		\wishbone_bd_ram_mem1_reg[51][13]/P0001 ,
		_w11938_,
		_w11979_,
		_w23485_
	);
	LUT4 #(
		.INIT('h0001)
	) name12973 (
		_w23482_,
		_w23483_,
		_w23484_,
		_w23485_,
		_w23486_
	);
	LUT3 #(
		.INIT('h80)
	) name12974 (
		\wishbone_bd_ram_mem1_reg[72][13]/P0001 ,
		_w11949_,
		_w11990_,
		_w23487_
	);
	LUT3 #(
		.INIT('h80)
	) name12975 (
		\wishbone_bd_ram_mem1_reg[223][13]/P0001 ,
		_w11973_,
		_w11984_,
		_w23488_
	);
	LUT3 #(
		.INIT('h80)
	) name12976 (
		\wishbone_bd_ram_mem1_reg[207][13]/P0001 ,
		_w11945_,
		_w11973_,
		_w23489_
	);
	LUT3 #(
		.INIT('h80)
	) name12977 (
		\wishbone_bd_ram_mem1_reg[242][13]/P0001 ,
		_w11952_,
		_w11963_,
		_w23490_
	);
	LUT4 #(
		.INIT('h0001)
	) name12978 (
		_w23487_,
		_w23488_,
		_w23489_,
		_w23490_,
		_w23491_
	);
	LUT3 #(
		.INIT('h80)
	) name12979 (
		\wishbone_bd_ram_mem1_reg[221][13]/P0001 ,
		_w11966_,
		_w11984_,
		_w23492_
	);
	LUT3 #(
		.INIT('h80)
	) name12980 (
		\wishbone_bd_ram_mem1_reg[230][13]/P0001 ,
		_w11982_,
		_w11986_,
		_w23493_
	);
	LUT3 #(
		.INIT('h80)
	) name12981 (
		\wishbone_bd_ram_mem1_reg[35][13]/P0001 ,
		_w11938_,
		_w11957_,
		_w23494_
	);
	LUT3 #(
		.INIT('h80)
	) name12982 (
		\wishbone_bd_ram_mem1_reg[241][13]/P0001 ,
		_w11952_,
		_w11977_,
		_w23495_
	);
	LUT4 #(
		.INIT('h0001)
	) name12983 (
		_w23492_,
		_w23493_,
		_w23494_,
		_w23495_,
		_w23496_
	);
	LUT3 #(
		.INIT('h80)
	) name12984 (
		\wishbone_bd_ram_mem1_reg[215][13]/P0001 ,
		_w11975_,
		_w11984_,
		_w23497_
	);
	LUT3 #(
		.INIT('h80)
	) name12985 (
		\wishbone_bd_ram_mem1_reg[64][13]/P0001 ,
		_w11941_,
		_w11949_,
		_w23498_
	);
	LUT3 #(
		.INIT('h80)
	) name12986 (
		\wishbone_bd_ram_mem1_reg[1][13]/P0001 ,
		_w11932_,
		_w11977_,
		_w23499_
	);
	LUT3 #(
		.INIT('h80)
	) name12987 (
		\wishbone_bd_ram_mem1_reg[58][13]/P0001 ,
		_w11944_,
		_w11979_,
		_w23500_
	);
	LUT4 #(
		.INIT('h0001)
	) name12988 (
		_w23497_,
		_w23498_,
		_w23499_,
		_w23500_,
		_w23501_
	);
	LUT4 #(
		.INIT('h8000)
	) name12989 (
		_w23486_,
		_w23491_,
		_w23496_,
		_w23501_,
		_w23502_
	);
	LUT4 #(
		.INIT('h8000)
	) name12990 (
		_w23439_,
		_w23460_,
		_w23481_,
		_w23502_,
		_w23503_
	);
	LUT3 #(
		.INIT('h80)
	) name12991 (
		\wishbone_bd_ram_mem1_reg[157][13]/P0001 ,
		_w11959_,
		_w11966_,
		_w23504_
	);
	LUT3 #(
		.INIT('h80)
	) name12992 (
		\wishbone_bd_ram_mem1_reg[186][13]/P0001 ,
		_w11942_,
		_w11944_,
		_w23505_
	);
	LUT3 #(
		.INIT('h80)
	) name12993 (
		\wishbone_bd_ram_mem1_reg[105][13]/P0001 ,
		_w11965_,
		_w11968_,
		_w23506_
	);
	LUT3 #(
		.INIT('h80)
	) name12994 (
		\wishbone_bd_ram_mem1_reg[245][13]/P0001 ,
		_w11933_,
		_w11952_,
		_w23507_
	);
	LUT4 #(
		.INIT('h0001)
	) name12995 (
		_w23504_,
		_w23505_,
		_w23506_,
		_w23507_,
		_w23508_
	);
	LUT3 #(
		.INIT('h80)
	) name12996 (
		\wishbone_bd_ram_mem1_reg[33][13]/P0001 ,
		_w11957_,
		_w11977_,
		_w23509_
	);
	LUT3 #(
		.INIT('h80)
	) name12997 (
		\wishbone_bd_ram_mem1_reg[162][13]/P0001 ,
		_w11930_,
		_w11963_,
		_w23510_
	);
	LUT3 #(
		.INIT('h80)
	) name12998 (
		\wishbone_bd_ram_mem1_reg[2][13]/P0001 ,
		_w11932_,
		_w11963_,
		_w23511_
	);
	LUT3 #(
		.INIT('h80)
	) name12999 (
		\wishbone_bd_ram_mem1_reg[238][13]/P0001 ,
		_w11948_,
		_w11982_,
		_w23512_
	);
	LUT4 #(
		.INIT('h0001)
	) name13000 (
		_w23509_,
		_w23510_,
		_w23511_,
		_w23512_,
		_w23513_
	);
	LUT3 #(
		.INIT('h80)
	) name13001 (
		\wishbone_bd_ram_mem1_reg[23][13]/P0001 ,
		_w11935_,
		_w11975_,
		_w23514_
	);
	LUT3 #(
		.INIT('h80)
	) name13002 (
		\wishbone_bd_ram_mem1_reg[124][13]/P0001 ,
		_w11954_,
		_w12012_,
		_w23515_
	);
	LUT3 #(
		.INIT('h80)
	) name13003 (
		\wishbone_bd_ram_mem1_reg[123][13]/P0001 ,
		_w11936_,
		_w12012_,
		_w23516_
	);
	LUT3 #(
		.INIT('h80)
	) name13004 (
		\wishbone_bd_ram_mem1_reg[0][13]/P0001 ,
		_w11932_,
		_w11941_,
		_w23517_
	);
	LUT4 #(
		.INIT('h0001)
	) name13005 (
		_w23514_,
		_w23515_,
		_w23516_,
		_w23517_,
		_w23518_
	);
	LUT3 #(
		.INIT('h80)
	) name13006 (
		\wishbone_bd_ram_mem1_reg[181][13]/P0001 ,
		_w11933_,
		_w11942_,
		_w23519_
	);
	LUT3 #(
		.INIT('h80)
	) name13007 (
		\wishbone_bd_ram_mem1_reg[9][13]/P0001 ,
		_w11932_,
		_w11968_,
		_w23520_
	);
	LUT3 #(
		.INIT('h80)
	) name13008 (
		\wishbone_bd_ram_mem1_reg[14][13]/P0001 ,
		_w11932_,
		_w11948_,
		_w23521_
	);
	LUT3 #(
		.INIT('h80)
	) name13009 (
		\wishbone_bd_ram_mem1_reg[212][13]/P0001 ,
		_w11929_,
		_w11984_,
		_w23522_
	);
	LUT4 #(
		.INIT('h0001)
	) name13010 (
		_w23519_,
		_w23520_,
		_w23521_,
		_w23522_,
		_w23523_
	);
	LUT4 #(
		.INIT('h8000)
	) name13011 (
		_w23508_,
		_w23513_,
		_w23518_,
		_w23523_,
		_w23524_
	);
	LUT3 #(
		.INIT('h80)
	) name13012 (
		\wishbone_bd_ram_mem1_reg[144][13]/P0001 ,
		_w11941_,
		_w11959_,
		_w23525_
	);
	LUT3 #(
		.INIT('h80)
	) name13013 (
		\wishbone_bd_ram_mem1_reg[25][13]/P0001 ,
		_w11935_,
		_w11968_,
		_w23526_
	);
	LUT3 #(
		.INIT('h80)
	) name13014 (
		\wishbone_bd_ram_mem1_reg[89][13]/P0001 ,
		_w11968_,
		_w11972_,
		_w23527_
	);
	LUT3 #(
		.INIT('h80)
	) name13015 (
		\wishbone_bd_ram_mem1_reg[192][13]/P0001 ,
		_w11941_,
		_w11945_,
		_w23528_
	);
	LUT4 #(
		.INIT('h0001)
	) name13016 (
		_w23525_,
		_w23526_,
		_w23527_,
		_w23528_,
		_w23529_
	);
	LUT3 #(
		.INIT('h80)
	) name13017 (
		\wishbone_bd_ram_mem1_reg[151][13]/P0001 ,
		_w11959_,
		_w11975_,
		_w23530_
	);
	LUT3 #(
		.INIT('h80)
	) name13018 (
		\wishbone_bd_ram_mem1_reg[11][13]/P0001 ,
		_w11932_,
		_w11936_,
		_w23531_
	);
	LUT3 #(
		.INIT('h80)
	) name13019 (
		\wishbone_bd_ram_mem1_reg[28][13]/P0001 ,
		_w11935_,
		_w11954_,
		_w23532_
	);
	LUT3 #(
		.INIT('h80)
	) name13020 (
		\wishbone_bd_ram_mem1_reg[226][13]/P0001 ,
		_w11963_,
		_w11982_,
		_w23533_
	);
	LUT4 #(
		.INIT('h0001)
	) name13021 (
		_w23530_,
		_w23531_,
		_w23532_,
		_w23533_,
		_w23534_
	);
	LUT3 #(
		.INIT('h80)
	) name13022 (
		\wishbone_bd_ram_mem1_reg[183][13]/P0001 ,
		_w11942_,
		_w11975_,
		_w23535_
	);
	LUT3 #(
		.INIT('h80)
	) name13023 (
		\wishbone_bd_ram_mem1_reg[15][13]/P0001 ,
		_w11932_,
		_w11973_,
		_w23536_
	);
	LUT3 #(
		.INIT('h80)
	) name13024 (
		\wishbone_bd_ram_mem1_reg[32][13]/P0001 ,
		_w11941_,
		_w11957_,
		_w23537_
	);
	LUT3 #(
		.INIT('h80)
	) name13025 (
		\wishbone_bd_ram_mem1_reg[16][13]/P0001 ,
		_w11935_,
		_w11941_,
		_w23538_
	);
	LUT4 #(
		.INIT('h0001)
	) name13026 (
		_w23535_,
		_w23536_,
		_w23537_,
		_w23538_,
		_w23539_
	);
	LUT3 #(
		.INIT('h80)
	) name13027 (
		\wishbone_bd_ram_mem1_reg[128][13]/P0001 ,
		_w11941_,
		_w11955_,
		_w23540_
	);
	LUT3 #(
		.INIT('h80)
	) name13028 (
		\wishbone_bd_ram_mem1_reg[236][13]/P0001 ,
		_w11954_,
		_w11982_,
		_w23541_
	);
	LUT3 #(
		.INIT('h80)
	) name13029 (
		\wishbone_bd_ram_mem1_reg[198][13]/P0001 ,
		_w11945_,
		_w11986_,
		_w23542_
	);
	LUT3 #(
		.INIT('h80)
	) name13030 (
		\wishbone_bd_ram_mem1_reg[147][13]/P0001 ,
		_w11938_,
		_w11959_,
		_w23543_
	);
	LUT4 #(
		.INIT('h0001)
	) name13031 (
		_w23540_,
		_w23541_,
		_w23542_,
		_w23543_,
		_w23544_
	);
	LUT4 #(
		.INIT('h8000)
	) name13032 (
		_w23529_,
		_w23534_,
		_w23539_,
		_w23544_,
		_w23545_
	);
	LUT3 #(
		.INIT('h80)
	) name13033 (
		\wishbone_bd_ram_mem1_reg[140][13]/P0001 ,
		_w11954_,
		_w11955_,
		_w23546_
	);
	LUT3 #(
		.INIT('h80)
	) name13034 (
		\wishbone_bd_ram_mem1_reg[67][13]/P0001 ,
		_w11938_,
		_w11949_,
		_w23547_
	);
	LUT3 #(
		.INIT('h80)
	) name13035 (
		\wishbone_bd_ram_mem1_reg[185][13]/P0001 ,
		_w11942_,
		_w11968_,
		_w23548_
	);
	LUT3 #(
		.INIT('h80)
	) name13036 (
		\wishbone_bd_ram_mem1_reg[202][13]/P0001 ,
		_w11944_,
		_w11945_,
		_w23549_
	);
	LUT4 #(
		.INIT('h0001)
	) name13037 (
		_w23546_,
		_w23547_,
		_w23548_,
		_w23549_,
		_w23550_
	);
	LUT3 #(
		.INIT('h80)
	) name13038 (
		\wishbone_bd_ram_mem1_reg[244][13]/P0001 ,
		_w11929_,
		_w11952_,
		_w23551_
	);
	LUT3 #(
		.INIT('h80)
	) name13039 (
		\wishbone_bd_ram_mem1_reg[228][13]/P0001 ,
		_w11929_,
		_w11982_,
		_w23552_
	);
	LUT3 #(
		.INIT('h80)
	) name13040 (
		\wishbone_bd_ram_mem1_reg[163][13]/P0001 ,
		_w11930_,
		_w11938_,
		_w23553_
	);
	LUT3 #(
		.INIT('h80)
	) name13041 (
		\wishbone_bd_ram_mem1_reg[121][13]/P0001 ,
		_w11968_,
		_w12012_,
		_w23554_
	);
	LUT4 #(
		.INIT('h0001)
	) name13042 (
		_w23551_,
		_w23552_,
		_w23553_,
		_w23554_,
		_w23555_
	);
	LUT3 #(
		.INIT('h80)
	) name13043 (
		\wishbone_bd_ram_mem1_reg[243][13]/P0001 ,
		_w11938_,
		_w11952_,
		_w23556_
	);
	LUT3 #(
		.INIT('h80)
	) name13044 (
		\wishbone_bd_ram_mem1_reg[210][13]/P0001 ,
		_w11963_,
		_w11984_,
		_w23557_
	);
	LUT3 #(
		.INIT('h80)
	) name13045 (
		\wishbone_bd_ram_mem1_reg[205][13]/P0001 ,
		_w11945_,
		_w11966_,
		_w23558_
	);
	LUT3 #(
		.INIT('h80)
	) name13046 (
		\wishbone_bd_ram_mem1_reg[48][13]/P0001 ,
		_w11941_,
		_w11979_,
		_w23559_
	);
	LUT4 #(
		.INIT('h0001)
	) name13047 (
		_w23556_,
		_w23557_,
		_w23558_,
		_w23559_,
		_w23560_
	);
	LUT3 #(
		.INIT('h80)
	) name13048 (
		\wishbone_bd_ram_mem1_reg[190][13]/P0001 ,
		_w11942_,
		_w11948_,
		_w23561_
	);
	LUT3 #(
		.INIT('h80)
	) name13049 (
		\wishbone_bd_ram_mem1_reg[4][13]/P0001 ,
		_w11929_,
		_w11932_,
		_w23562_
	);
	LUT3 #(
		.INIT('h80)
	) name13050 (
		\wishbone_bd_ram_mem1_reg[193][13]/P0001 ,
		_w11945_,
		_w11977_,
		_w23563_
	);
	LUT3 #(
		.INIT('h80)
	) name13051 (
		\wishbone_bd_ram_mem1_reg[204][13]/P0001 ,
		_w11945_,
		_w11954_,
		_w23564_
	);
	LUT4 #(
		.INIT('h0001)
	) name13052 (
		_w23561_,
		_w23562_,
		_w23563_,
		_w23564_,
		_w23565_
	);
	LUT4 #(
		.INIT('h8000)
	) name13053 (
		_w23550_,
		_w23555_,
		_w23560_,
		_w23565_,
		_w23566_
	);
	LUT3 #(
		.INIT('h80)
	) name13054 (
		\wishbone_bd_ram_mem1_reg[173][13]/P0001 ,
		_w11930_,
		_w11966_,
		_w23567_
	);
	LUT3 #(
		.INIT('h80)
	) name13055 (
		\wishbone_bd_ram_mem1_reg[46][13]/P0001 ,
		_w11948_,
		_w11957_,
		_w23568_
	);
	LUT3 #(
		.INIT('h80)
	) name13056 (
		\wishbone_bd_ram_mem1_reg[119][13]/P0001 ,
		_w11975_,
		_w12012_,
		_w23569_
	);
	LUT3 #(
		.INIT('h80)
	) name13057 (
		\wishbone_bd_ram_mem1_reg[43][13]/P0001 ,
		_w11936_,
		_w11957_,
		_w23570_
	);
	LUT4 #(
		.INIT('h0001)
	) name13058 (
		_w23567_,
		_w23568_,
		_w23569_,
		_w23570_,
		_w23571_
	);
	LUT3 #(
		.INIT('h80)
	) name13059 (
		\wishbone_bd_ram_mem1_reg[196][13]/P0001 ,
		_w11929_,
		_w11945_,
		_w23572_
	);
	LUT3 #(
		.INIT('h80)
	) name13060 (
		\wishbone_bd_ram_mem1_reg[189][13]/P0001 ,
		_w11942_,
		_w11966_,
		_w23573_
	);
	LUT3 #(
		.INIT('h80)
	) name13061 (
		\wishbone_bd_ram_mem1_reg[83][13]/P0001 ,
		_w11938_,
		_w11972_,
		_w23574_
	);
	LUT3 #(
		.INIT('h80)
	) name13062 (
		\wishbone_bd_ram_mem1_reg[231][13]/P0001 ,
		_w11975_,
		_w11982_,
		_w23575_
	);
	LUT4 #(
		.INIT('h0001)
	) name13063 (
		_w23572_,
		_w23573_,
		_w23574_,
		_w23575_,
		_w23576_
	);
	LUT3 #(
		.INIT('h80)
	) name13064 (
		\wishbone_bd_ram_mem1_reg[129][13]/P0001 ,
		_w11955_,
		_w11977_,
		_w23577_
	);
	LUT3 #(
		.INIT('h80)
	) name13065 (
		\wishbone_bd_ram_mem1_reg[254][13]/P0001 ,
		_w11948_,
		_w11952_,
		_w23578_
	);
	LUT3 #(
		.INIT('h80)
	) name13066 (
		\wishbone_bd_ram_mem1_reg[139][13]/P0001 ,
		_w11936_,
		_w11955_,
		_w23579_
	);
	LUT3 #(
		.INIT('h80)
	) name13067 (
		\wishbone_bd_ram_mem1_reg[159][13]/P0001 ,
		_w11959_,
		_w11973_,
		_w23580_
	);
	LUT4 #(
		.INIT('h0001)
	) name13068 (
		_w23577_,
		_w23578_,
		_w23579_,
		_w23580_,
		_w23581_
	);
	LUT3 #(
		.INIT('h80)
	) name13069 (
		\wishbone_bd_ram_mem1_reg[73][13]/P0001 ,
		_w11949_,
		_w11968_,
		_w23582_
	);
	LUT3 #(
		.INIT('h80)
	) name13070 (
		\wishbone_bd_ram_mem1_reg[225][13]/P0001 ,
		_w11977_,
		_w11982_,
		_w23583_
	);
	LUT3 #(
		.INIT('h80)
	) name13071 (
		\wishbone_bd_ram_mem1_reg[106][13]/P0001 ,
		_w11944_,
		_w11965_,
		_w23584_
	);
	LUT3 #(
		.INIT('h80)
	) name13072 (
		\wishbone_bd_ram_mem1_reg[98][13]/P0001 ,
		_w11963_,
		_w11965_,
		_w23585_
	);
	LUT4 #(
		.INIT('h0001)
	) name13073 (
		_w23582_,
		_w23583_,
		_w23584_,
		_w23585_,
		_w23586_
	);
	LUT4 #(
		.INIT('h8000)
	) name13074 (
		_w23571_,
		_w23576_,
		_w23581_,
		_w23586_,
		_w23587_
	);
	LUT4 #(
		.INIT('h8000)
	) name13075 (
		_w23524_,
		_w23545_,
		_w23566_,
		_w23587_,
		_w23588_
	);
	LUT4 #(
		.INIT('h8000)
	) name13076 (
		_w23333_,
		_w23418_,
		_w23503_,
		_w23588_,
		_w23589_
	);
	LUT2 #(
		.INIT('h1)
	) name13077 (
		wb_rst_i_pad,
		_w23247_,
		_w23590_
	);
	LUT3 #(
		.INIT('hba)
	) name13078 (
		_w23248_,
		_w23589_,
		_w23590_,
		_w23591_
	);
	LUT3 #(
		.INIT('h80)
	) name13079 (
		\ethreg1_MODER_1_DataOut_reg[6]/NET0131 ,
		_w18800_,
		_w18801_,
		_w23592_
	);
	LUT4 #(
		.INIT('h0020)
	) name13080 (
		\ethreg1_TXCTRL_1_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23593_
	);
	LUT3 #(
		.INIT('h80)
	) name13081 (
		_w18757_,
		_w18758_,
		_w23593_,
		_w23594_
	);
	LUT4 #(
		.INIT('h0008)
	) name13082 (
		\ethreg1_RXHASH0_1_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23595_
	);
	LUT3 #(
		.INIT('h80)
	) name13083 (
		_w18757_,
		_w18758_,
		_w23595_,
		_w23596_
	);
	LUT4 #(
		.INIT('h0008)
	) name13084 (
		\ethreg1_RXHASH1_1_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23597_
	);
	LUT3 #(
		.INIT('h80)
	) name13085 (
		_w18757_,
		_w18762_,
		_w23597_,
		_w23598_
	);
	LUT4 #(
		.INIT('h0001)
	) name13086 (
		_w23592_,
		_w23594_,
		_w23596_,
		_w23598_,
		_w23599_
	);
	LUT3 #(
		.INIT('h80)
	) name13087 (
		\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 ,
		_w18753_,
		_w18754_,
		_w23600_
	);
	LUT3 #(
		.INIT('h80)
	) name13088 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[6]/NET0131 ,
		_w18798_,
		_w18805_,
		_w23601_
	);
	LUT4 #(
		.INIT('h0002)
	) name13089 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23602_
	);
	LUT3 #(
		.INIT('h80)
	) name13090 (
		_w18757_,
		_w18758_,
		_w23602_,
		_w23603_
	);
	LUT4 #(
		.INIT('h0002)
	) name13091 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23604_
	);
	LUT3 #(
		.INIT('h80)
	) name13092 (
		_w18757_,
		_w18762_,
		_w23604_,
		_w23605_
	);
	LUT3 #(
		.INIT('h80)
	) name13093 (
		\ethreg1_MIIRX_DATA_DataOut_reg[14]/NET0131 ,
		_w18785_,
		_w18786_,
		_w23606_
	);
	LUT4 #(
		.INIT('h0001)
	) name13094 (
		_w23601_,
		_w23603_,
		_w23605_,
		_w23606_,
		_w23607_
	);
	LUT4 #(
		.INIT('h0800)
	) name13095 (
		_w18752_,
		_w23599_,
		_w23600_,
		_w23607_,
		_w23608_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name13096 (
		_w18752_,
		_w23599_,
		_w23600_,
		_w23607_,
		_w23609_
	);
	LUT3 #(
		.INIT('h80)
	) name13097 (
		\wishbone_bd_ram_mem1_reg[107][14]/P0001 ,
		_w11936_,
		_w11965_,
		_w23610_
	);
	LUT3 #(
		.INIT('h80)
	) name13098 (
		\wishbone_bd_ram_mem1_reg[95][14]/P0001 ,
		_w11972_,
		_w11973_,
		_w23611_
	);
	LUT3 #(
		.INIT('h80)
	) name13099 (
		\wishbone_bd_ram_mem1_reg[164][14]/P0001 ,
		_w11929_,
		_w11930_,
		_w23612_
	);
	LUT3 #(
		.INIT('h80)
	) name13100 (
		\wishbone_bd_ram_mem1_reg[207][14]/P0001 ,
		_w11945_,
		_w11973_,
		_w23613_
	);
	LUT4 #(
		.INIT('h0001)
	) name13101 (
		_w23610_,
		_w23611_,
		_w23612_,
		_w23613_,
		_w23614_
	);
	LUT3 #(
		.INIT('h80)
	) name13102 (
		\wishbone_bd_ram_mem1_reg[198][14]/P0001 ,
		_w11945_,
		_w11986_,
		_w23615_
	);
	LUT3 #(
		.INIT('h80)
	) name13103 (
		\wishbone_bd_ram_mem1_reg[137][14]/P0001 ,
		_w11955_,
		_w11968_,
		_w23616_
	);
	LUT3 #(
		.INIT('h80)
	) name13104 (
		\wishbone_bd_ram_mem1_reg[4][14]/P0001 ,
		_w11929_,
		_w11932_,
		_w23617_
	);
	LUT3 #(
		.INIT('h80)
	) name13105 (
		\wishbone_bd_ram_mem1_reg[220][14]/P0001 ,
		_w11954_,
		_w11984_,
		_w23618_
	);
	LUT4 #(
		.INIT('h0001)
	) name13106 (
		_w23615_,
		_w23616_,
		_w23617_,
		_w23618_,
		_w23619_
	);
	LUT3 #(
		.INIT('h80)
	) name13107 (
		\wishbone_bd_ram_mem1_reg[206][14]/P0001 ,
		_w11945_,
		_w11948_,
		_w23620_
	);
	LUT3 #(
		.INIT('h80)
	) name13108 (
		\wishbone_bd_ram_mem1_reg[140][14]/P0001 ,
		_w11954_,
		_w11955_,
		_w23621_
	);
	LUT3 #(
		.INIT('h80)
	) name13109 (
		\wishbone_bd_ram_mem1_reg[2][14]/P0001 ,
		_w11932_,
		_w11963_,
		_w23622_
	);
	LUT3 #(
		.INIT('h80)
	) name13110 (
		\wishbone_bd_ram_mem1_reg[112][14]/P0001 ,
		_w11941_,
		_w12012_,
		_w23623_
	);
	LUT4 #(
		.INIT('h0001)
	) name13111 (
		_w23620_,
		_w23621_,
		_w23622_,
		_w23623_,
		_w23624_
	);
	LUT3 #(
		.INIT('h80)
	) name13112 (
		\wishbone_bd_ram_mem1_reg[45][14]/P0001 ,
		_w11957_,
		_w11966_,
		_w23625_
	);
	LUT3 #(
		.INIT('h80)
	) name13113 (
		\wishbone_bd_ram_mem1_reg[202][14]/P0001 ,
		_w11944_,
		_w11945_,
		_w23626_
	);
	LUT3 #(
		.INIT('h80)
	) name13114 (
		\wishbone_bd_ram_mem1_reg[76][14]/P0001 ,
		_w11949_,
		_w11954_,
		_w23627_
	);
	LUT3 #(
		.INIT('h80)
	) name13115 (
		\wishbone_bd_ram_mem1_reg[170][14]/P0001 ,
		_w11930_,
		_w11944_,
		_w23628_
	);
	LUT4 #(
		.INIT('h0001)
	) name13116 (
		_w23625_,
		_w23626_,
		_w23627_,
		_w23628_,
		_w23629_
	);
	LUT4 #(
		.INIT('h8000)
	) name13117 (
		_w23614_,
		_w23619_,
		_w23624_,
		_w23629_,
		_w23630_
	);
	LUT3 #(
		.INIT('h80)
	) name13118 (
		\wishbone_bd_ram_mem1_reg[0][14]/P0001 ,
		_w11932_,
		_w11941_,
		_w23631_
	);
	LUT3 #(
		.INIT('h80)
	) name13119 (
		\wishbone_bd_ram_mem1_reg[56][14]/P0001 ,
		_w11979_,
		_w11990_,
		_w23632_
	);
	LUT3 #(
		.INIT('h80)
	) name13120 (
		\wishbone_bd_ram_mem1_reg[247][14]/P0001 ,
		_w11952_,
		_w11975_,
		_w23633_
	);
	LUT3 #(
		.INIT('h80)
	) name13121 (
		\wishbone_bd_ram_mem1_reg[101][14]/P0001 ,
		_w11933_,
		_w11965_,
		_w23634_
	);
	LUT4 #(
		.INIT('h0001)
	) name13122 (
		_w23631_,
		_w23632_,
		_w23633_,
		_w23634_,
		_w23635_
	);
	LUT3 #(
		.INIT('h80)
	) name13123 (
		\wishbone_bd_ram_mem1_reg[114][14]/P0001 ,
		_w11963_,
		_w12012_,
		_w23636_
	);
	LUT3 #(
		.INIT('h80)
	) name13124 (
		\wishbone_bd_ram_mem1_reg[209][14]/P0001 ,
		_w11977_,
		_w11984_,
		_w23637_
	);
	LUT3 #(
		.INIT('h80)
	) name13125 (
		\wishbone_bd_ram_mem1_reg[28][14]/P0001 ,
		_w11935_,
		_w11954_,
		_w23638_
	);
	LUT3 #(
		.INIT('h80)
	) name13126 (
		\wishbone_bd_ram_mem1_reg[69][14]/P0001 ,
		_w11933_,
		_w11949_,
		_w23639_
	);
	LUT4 #(
		.INIT('h0001)
	) name13127 (
		_w23636_,
		_w23637_,
		_w23638_,
		_w23639_,
		_w23640_
	);
	LUT3 #(
		.INIT('h80)
	) name13128 (
		\wishbone_bd_ram_mem1_reg[177][14]/P0001 ,
		_w11942_,
		_w11977_,
		_w23641_
	);
	LUT3 #(
		.INIT('h80)
	) name13129 (
		\wishbone_bd_ram_mem1_reg[217][14]/P0001 ,
		_w11968_,
		_w11984_,
		_w23642_
	);
	LUT3 #(
		.INIT('h80)
	) name13130 (
		\wishbone_bd_ram_mem1_reg[194][14]/P0001 ,
		_w11945_,
		_w11963_,
		_w23643_
	);
	LUT3 #(
		.INIT('h80)
	) name13131 (
		\wishbone_bd_ram_mem1_reg[255][14]/P0001 ,
		_w11952_,
		_w11973_,
		_w23644_
	);
	LUT4 #(
		.INIT('h0001)
	) name13132 (
		_w23641_,
		_w23642_,
		_w23643_,
		_w23644_,
		_w23645_
	);
	LUT3 #(
		.INIT('h80)
	) name13133 (
		\wishbone_bd_ram_mem1_reg[242][14]/P0001 ,
		_w11952_,
		_w11963_,
		_w23646_
	);
	LUT3 #(
		.INIT('h80)
	) name13134 (
		\wishbone_bd_ram_mem1_reg[223][14]/P0001 ,
		_w11973_,
		_w11984_,
		_w23647_
	);
	LUT3 #(
		.INIT('h80)
	) name13135 (
		\wishbone_bd_ram_mem1_reg[214][14]/P0001 ,
		_w11984_,
		_w11986_,
		_w23648_
	);
	LUT3 #(
		.INIT('h80)
	) name13136 (
		\wishbone_bd_ram_mem1_reg[190][14]/P0001 ,
		_w11942_,
		_w11948_,
		_w23649_
	);
	LUT4 #(
		.INIT('h0001)
	) name13137 (
		_w23646_,
		_w23647_,
		_w23648_,
		_w23649_,
		_w23650_
	);
	LUT4 #(
		.INIT('h8000)
	) name13138 (
		_w23635_,
		_w23640_,
		_w23645_,
		_w23650_,
		_w23651_
	);
	LUT3 #(
		.INIT('h80)
	) name13139 (
		\wishbone_bd_ram_mem1_reg[224][14]/P0001 ,
		_w11941_,
		_w11982_,
		_w23652_
	);
	LUT3 #(
		.INIT('h80)
	) name13140 (
		\wishbone_bd_ram_mem1_reg[41][14]/P0001 ,
		_w11957_,
		_w11968_,
		_w23653_
	);
	LUT3 #(
		.INIT('h80)
	) name13141 (
		\wishbone_bd_ram_mem1_reg[195][14]/P0001 ,
		_w11938_,
		_w11945_,
		_w23654_
	);
	LUT3 #(
		.INIT('h80)
	) name13142 (
		\wishbone_bd_ram_mem1_reg[183][14]/P0001 ,
		_w11942_,
		_w11975_,
		_w23655_
	);
	LUT4 #(
		.INIT('h0001)
	) name13143 (
		_w23652_,
		_w23653_,
		_w23654_,
		_w23655_,
		_w23656_
	);
	LUT3 #(
		.INIT('h80)
	) name13144 (
		\wishbone_bd_ram_mem1_reg[205][14]/P0001 ,
		_w11945_,
		_w11966_,
		_w23657_
	);
	LUT3 #(
		.INIT('h80)
	) name13145 (
		\wishbone_bd_ram_mem1_reg[12][14]/P0001 ,
		_w11932_,
		_w11954_,
		_w23658_
	);
	LUT3 #(
		.INIT('h80)
	) name13146 (
		\wishbone_bd_ram_mem1_reg[253][14]/P0001 ,
		_w11952_,
		_w11966_,
		_w23659_
	);
	LUT3 #(
		.INIT('h80)
	) name13147 (
		\wishbone_bd_ram_mem1_reg[156][14]/P0001 ,
		_w11954_,
		_w11959_,
		_w23660_
	);
	LUT4 #(
		.INIT('h0001)
	) name13148 (
		_w23657_,
		_w23658_,
		_w23659_,
		_w23660_,
		_w23661_
	);
	LUT3 #(
		.INIT('h80)
	) name13149 (
		\wishbone_bd_ram_mem1_reg[131][14]/P0001 ,
		_w11938_,
		_w11955_,
		_w23662_
	);
	LUT3 #(
		.INIT('h80)
	) name13150 (
		\wishbone_bd_ram_mem1_reg[73][14]/P0001 ,
		_w11949_,
		_w11968_,
		_w23663_
	);
	LUT3 #(
		.INIT('h80)
	) name13151 (
		\wishbone_bd_ram_mem1_reg[31][14]/P0001 ,
		_w11935_,
		_w11973_,
		_w23664_
	);
	LUT3 #(
		.INIT('h80)
	) name13152 (
		\wishbone_bd_ram_mem1_reg[216][14]/P0001 ,
		_w11984_,
		_w11990_,
		_w23665_
	);
	LUT4 #(
		.INIT('h0001)
	) name13153 (
		_w23662_,
		_w23663_,
		_w23664_,
		_w23665_,
		_w23666_
	);
	LUT3 #(
		.INIT('h80)
	) name13154 (
		\wishbone_bd_ram_mem1_reg[231][14]/P0001 ,
		_w11975_,
		_w11982_,
		_w23667_
	);
	LUT3 #(
		.INIT('h80)
	) name13155 (
		\wishbone_bd_ram_mem1_reg[221][14]/P0001 ,
		_w11966_,
		_w11984_,
		_w23668_
	);
	LUT3 #(
		.INIT('h80)
	) name13156 (
		\wishbone_bd_ram_mem1_reg[13][14]/P0001 ,
		_w11932_,
		_w11966_,
		_w23669_
	);
	LUT3 #(
		.INIT('h80)
	) name13157 (
		\wishbone_bd_ram_mem1_reg[238][14]/P0001 ,
		_w11948_,
		_w11982_,
		_w23670_
	);
	LUT4 #(
		.INIT('h0001)
	) name13158 (
		_w23667_,
		_w23668_,
		_w23669_,
		_w23670_,
		_w23671_
	);
	LUT4 #(
		.INIT('h8000)
	) name13159 (
		_w23656_,
		_w23661_,
		_w23666_,
		_w23671_,
		_w23672_
	);
	LUT3 #(
		.INIT('h80)
	) name13160 (
		\wishbone_bd_ram_mem1_reg[123][14]/P0001 ,
		_w11936_,
		_w12012_,
		_w23673_
	);
	LUT3 #(
		.INIT('h80)
	) name13161 (
		\wishbone_bd_ram_mem1_reg[189][14]/P0001 ,
		_w11942_,
		_w11966_,
		_w23674_
	);
	LUT3 #(
		.INIT('h80)
	) name13162 (
		\wishbone_bd_ram_mem1_reg[146][14]/P0001 ,
		_w11959_,
		_w11963_,
		_w23675_
	);
	LUT3 #(
		.INIT('h80)
	) name13163 (
		\wishbone_bd_ram_mem1_reg[72][14]/P0001 ,
		_w11949_,
		_w11990_,
		_w23676_
	);
	LUT4 #(
		.INIT('h0001)
	) name13164 (
		_w23673_,
		_w23674_,
		_w23675_,
		_w23676_,
		_w23677_
	);
	LUT3 #(
		.INIT('h80)
	) name13165 (
		\wishbone_bd_ram_mem1_reg[248][14]/P0001 ,
		_w11952_,
		_w11990_,
		_w23678_
	);
	LUT3 #(
		.INIT('h80)
	) name13166 (
		\wishbone_bd_ram_mem1_reg[126][14]/P0001 ,
		_w11948_,
		_w12012_,
		_w23679_
	);
	LUT3 #(
		.INIT('h80)
	) name13167 (
		\wishbone_bd_ram_mem1_reg[8][14]/P0001 ,
		_w11932_,
		_w11990_,
		_w23680_
	);
	LUT3 #(
		.INIT('h80)
	) name13168 (
		\wishbone_bd_ram_mem1_reg[218][14]/P0001 ,
		_w11944_,
		_w11984_,
		_w23681_
	);
	LUT4 #(
		.INIT('h0001)
	) name13169 (
		_w23678_,
		_w23679_,
		_w23680_,
		_w23681_,
		_w23682_
	);
	LUT3 #(
		.INIT('h80)
	) name13170 (
		\wishbone_bd_ram_mem1_reg[98][14]/P0001 ,
		_w11963_,
		_w11965_,
		_w23683_
	);
	LUT3 #(
		.INIT('h80)
	) name13171 (
		\wishbone_bd_ram_mem1_reg[172][14]/P0001 ,
		_w11930_,
		_w11954_,
		_w23684_
	);
	LUT3 #(
		.INIT('h80)
	) name13172 (
		\wishbone_bd_ram_mem1_reg[53][14]/P0001 ,
		_w11933_,
		_w11979_,
		_w23685_
	);
	LUT3 #(
		.INIT('h80)
	) name13173 (
		\wishbone_bd_ram_mem1_reg[148][14]/P0001 ,
		_w11929_,
		_w11959_,
		_w23686_
	);
	LUT4 #(
		.INIT('h0001)
	) name13174 (
		_w23683_,
		_w23684_,
		_w23685_,
		_w23686_,
		_w23687_
	);
	LUT3 #(
		.INIT('h80)
	) name13175 (
		\wishbone_bd_ram_mem1_reg[134][14]/P0001 ,
		_w11955_,
		_w11986_,
		_w23688_
	);
	LUT3 #(
		.INIT('h80)
	) name13176 (
		\wishbone_bd_ram_mem1_reg[54][14]/P0001 ,
		_w11979_,
		_w11986_,
		_w23689_
	);
	LUT3 #(
		.INIT('h80)
	) name13177 (
		\wishbone_bd_ram_mem1_reg[203][14]/P0001 ,
		_w11936_,
		_w11945_,
		_w23690_
	);
	LUT3 #(
		.INIT('h80)
	) name13178 (
		\wishbone_bd_ram_mem1_reg[230][14]/P0001 ,
		_w11982_,
		_w11986_,
		_w23691_
	);
	LUT4 #(
		.INIT('h0001)
	) name13179 (
		_w23688_,
		_w23689_,
		_w23690_,
		_w23691_,
		_w23692_
	);
	LUT4 #(
		.INIT('h8000)
	) name13180 (
		_w23677_,
		_w23682_,
		_w23687_,
		_w23692_,
		_w23693_
	);
	LUT4 #(
		.INIT('h8000)
	) name13181 (
		_w23630_,
		_w23651_,
		_w23672_,
		_w23693_,
		_w23694_
	);
	LUT3 #(
		.INIT('h80)
	) name13182 (
		\wishbone_bd_ram_mem1_reg[68][14]/P0001 ,
		_w11929_,
		_w11949_,
		_w23695_
	);
	LUT3 #(
		.INIT('h80)
	) name13183 (
		\wishbone_bd_ram_mem1_reg[132][14]/P0001 ,
		_w11929_,
		_w11955_,
		_w23696_
	);
	LUT3 #(
		.INIT('h80)
	) name13184 (
		\wishbone_bd_ram_mem1_reg[87][14]/P0001 ,
		_w11972_,
		_w11975_,
		_w23697_
	);
	LUT3 #(
		.INIT('h80)
	) name13185 (
		\wishbone_bd_ram_mem1_reg[108][14]/P0001 ,
		_w11954_,
		_w11965_,
		_w23698_
	);
	LUT4 #(
		.INIT('h0001)
	) name13186 (
		_w23695_,
		_w23696_,
		_w23697_,
		_w23698_,
		_w23699_
	);
	LUT3 #(
		.INIT('h80)
	) name13187 (
		\wishbone_bd_ram_mem1_reg[197][14]/P0001 ,
		_w11933_,
		_w11945_,
		_w23700_
	);
	LUT3 #(
		.INIT('h80)
	) name13188 (
		\wishbone_bd_ram_mem1_reg[222][14]/P0001 ,
		_w11948_,
		_w11984_,
		_w23701_
	);
	LUT3 #(
		.INIT('h80)
	) name13189 (
		\wishbone_bd_ram_mem1_reg[16][14]/P0001 ,
		_w11935_,
		_w11941_,
		_w23702_
	);
	LUT3 #(
		.INIT('h80)
	) name13190 (
		\wishbone_bd_ram_mem1_reg[135][14]/P0001 ,
		_w11955_,
		_w11975_,
		_w23703_
	);
	LUT4 #(
		.INIT('h0001)
	) name13191 (
		_w23700_,
		_w23701_,
		_w23702_,
		_w23703_,
		_w23704_
	);
	LUT3 #(
		.INIT('h80)
	) name13192 (
		\wishbone_bd_ram_mem1_reg[75][14]/P0001 ,
		_w11936_,
		_w11949_,
		_w23705_
	);
	LUT3 #(
		.INIT('h80)
	) name13193 (
		\wishbone_bd_ram_mem1_reg[70][14]/P0001 ,
		_w11949_,
		_w11986_,
		_w23706_
	);
	LUT3 #(
		.INIT('h80)
	) name13194 (
		\wishbone_bd_ram_mem1_reg[155][14]/P0001 ,
		_w11936_,
		_w11959_,
		_w23707_
	);
	LUT3 #(
		.INIT('h80)
	) name13195 (
		\wishbone_bd_ram_mem1_reg[243][14]/P0001 ,
		_w11938_,
		_w11952_,
		_w23708_
	);
	LUT4 #(
		.INIT('h0001)
	) name13196 (
		_w23705_,
		_w23706_,
		_w23707_,
		_w23708_,
		_w23709_
	);
	LUT3 #(
		.INIT('h80)
	) name13197 (
		\wishbone_bd_ram_mem1_reg[210][14]/P0001 ,
		_w11963_,
		_w11984_,
		_w23710_
	);
	LUT3 #(
		.INIT('h80)
	) name13198 (
		\wishbone_bd_ram_mem1_reg[85][14]/P0001 ,
		_w11933_,
		_w11972_,
		_w23711_
	);
	LUT3 #(
		.INIT('h80)
	) name13199 (
		\wishbone_bd_ram_mem1_reg[50][14]/P0001 ,
		_w11963_,
		_w11979_,
		_w23712_
	);
	LUT3 #(
		.INIT('h80)
	) name13200 (
		\wishbone_bd_ram_mem1_reg[176][14]/P0001 ,
		_w11941_,
		_w11942_,
		_w23713_
	);
	LUT4 #(
		.INIT('h0001)
	) name13201 (
		_w23710_,
		_w23711_,
		_w23712_,
		_w23713_,
		_w23714_
	);
	LUT4 #(
		.INIT('h8000)
	) name13202 (
		_w23699_,
		_w23704_,
		_w23709_,
		_w23714_,
		_w23715_
	);
	LUT3 #(
		.INIT('h80)
	) name13203 (
		\wishbone_bd_ram_mem1_reg[33][14]/P0001 ,
		_w11957_,
		_w11977_,
		_w23716_
	);
	LUT3 #(
		.INIT('h80)
	) name13204 (
		\wishbone_bd_ram_mem1_reg[113][14]/P0001 ,
		_w11977_,
		_w12012_,
		_w23717_
	);
	LUT3 #(
		.INIT('h80)
	) name13205 (
		\wishbone_bd_ram_mem1_reg[44][14]/P0001 ,
		_w11954_,
		_w11957_,
		_w23718_
	);
	LUT3 #(
		.INIT('h80)
	) name13206 (
		\wishbone_bd_ram_mem1_reg[237][14]/P0001 ,
		_w11966_,
		_w11982_,
		_w23719_
	);
	LUT4 #(
		.INIT('h0001)
	) name13207 (
		_w23716_,
		_w23717_,
		_w23718_,
		_w23719_,
		_w23720_
	);
	LUT3 #(
		.INIT('h80)
	) name13208 (
		\wishbone_bd_ram_mem1_reg[18][14]/P0001 ,
		_w11935_,
		_w11963_,
		_w23721_
	);
	LUT3 #(
		.INIT('h80)
	) name13209 (
		\wishbone_bd_ram_mem1_reg[58][14]/P0001 ,
		_w11944_,
		_w11979_,
		_w23722_
	);
	LUT3 #(
		.INIT('h80)
	) name13210 (
		\wishbone_bd_ram_mem1_reg[171][14]/P0001 ,
		_w11930_,
		_w11936_,
		_w23723_
	);
	LUT3 #(
		.INIT('h80)
	) name13211 (
		\wishbone_bd_ram_mem1_reg[118][14]/P0001 ,
		_w11986_,
		_w12012_,
		_w23724_
	);
	LUT4 #(
		.INIT('h0001)
	) name13212 (
		_w23721_,
		_w23722_,
		_w23723_,
		_w23724_,
		_w23725_
	);
	LUT3 #(
		.INIT('h80)
	) name13213 (
		\wishbone_bd_ram_mem1_reg[78][14]/P0001 ,
		_w11948_,
		_w11949_,
		_w23726_
	);
	LUT3 #(
		.INIT('h80)
	) name13214 (
		\wishbone_bd_ram_mem1_reg[46][14]/P0001 ,
		_w11948_,
		_w11957_,
		_w23727_
	);
	LUT3 #(
		.INIT('h80)
	) name13215 (
		\wishbone_bd_ram_mem1_reg[157][14]/P0001 ,
		_w11959_,
		_w11966_,
		_w23728_
	);
	LUT3 #(
		.INIT('h80)
	) name13216 (
		\wishbone_bd_ram_mem1_reg[81][14]/P0001 ,
		_w11972_,
		_w11977_,
		_w23729_
	);
	LUT4 #(
		.INIT('h0001)
	) name13217 (
		_w23726_,
		_w23727_,
		_w23728_,
		_w23729_,
		_w23730_
	);
	LUT3 #(
		.INIT('h80)
	) name13218 (
		\wishbone_bd_ram_mem1_reg[29][14]/P0001 ,
		_w11935_,
		_w11966_,
		_w23731_
	);
	LUT3 #(
		.INIT('h80)
	) name13219 (
		\wishbone_bd_ram_mem1_reg[241][14]/P0001 ,
		_w11952_,
		_w11977_,
		_w23732_
	);
	LUT3 #(
		.INIT('h80)
	) name13220 (
		\wishbone_bd_ram_mem1_reg[211][14]/P0001 ,
		_w11938_,
		_w11984_,
		_w23733_
	);
	LUT3 #(
		.INIT('h80)
	) name13221 (
		\wishbone_bd_ram_mem1_reg[66][14]/P0001 ,
		_w11949_,
		_w11963_,
		_w23734_
	);
	LUT4 #(
		.INIT('h0001)
	) name13222 (
		_w23731_,
		_w23732_,
		_w23733_,
		_w23734_,
		_w23735_
	);
	LUT4 #(
		.INIT('h8000)
	) name13223 (
		_w23720_,
		_w23725_,
		_w23730_,
		_w23735_,
		_w23736_
	);
	LUT3 #(
		.INIT('h80)
	) name13224 (
		\wishbone_bd_ram_mem1_reg[138][14]/P0001 ,
		_w11944_,
		_w11955_,
		_w23737_
	);
	LUT3 #(
		.INIT('h80)
	) name13225 (
		\wishbone_bd_ram_mem1_reg[116][14]/P0001 ,
		_w11929_,
		_w12012_,
		_w23738_
	);
	LUT3 #(
		.INIT('h80)
	) name13226 (
		\wishbone_bd_ram_mem1_reg[121][14]/P0001 ,
		_w11968_,
		_w12012_,
		_w23739_
	);
	LUT3 #(
		.INIT('h80)
	) name13227 (
		\wishbone_bd_ram_mem1_reg[204][14]/P0001 ,
		_w11945_,
		_w11954_,
		_w23740_
	);
	LUT4 #(
		.INIT('h0001)
	) name13228 (
		_w23737_,
		_w23738_,
		_w23739_,
		_w23740_,
		_w23741_
	);
	LUT3 #(
		.INIT('h80)
	) name13229 (
		\wishbone_bd_ram_mem1_reg[212][14]/P0001 ,
		_w11929_,
		_w11984_,
		_w23742_
	);
	LUT3 #(
		.INIT('h80)
	) name13230 (
		\wishbone_bd_ram_mem1_reg[233][14]/P0001 ,
		_w11968_,
		_w11982_,
		_w23743_
	);
	LUT3 #(
		.INIT('h80)
	) name13231 (
		\wishbone_bd_ram_mem1_reg[43][14]/P0001 ,
		_w11936_,
		_w11957_,
		_w23744_
	);
	LUT3 #(
		.INIT('h80)
	) name13232 (
		\wishbone_bd_ram_mem1_reg[27][14]/P0001 ,
		_w11935_,
		_w11936_,
		_w23745_
	);
	LUT4 #(
		.INIT('h0001)
	) name13233 (
		_w23742_,
		_w23743_,
		_w23744_,
		_w23745_,
		_w23746_
	);
	LUT3 #(
		.INIT('h80)
	) name13234 (
		\wishbone_bd_ram_mem1_reg[178][14]/P0001 ,
		_w11942_,
		_w11963_,
		_w23747_
	);
	LUT3 #(
		.INIT('h80)
	) name13235 (
		\wishbone_bd_ram_mem1_reg[1][14]/P0001 ,
		_w11932_,
		_w11977_,
		_w23748_
	);
	LUT3 #(
		.INIT('h80)
	) name13236 (
		\wishbone_bd_ram_mem1_reg[232][14]/P0001 ,
		_w11982_,
		_w11990_,
		_w23749_
	);
	LUT3 #(
		.INIT('h80)
	) name13237 (
		\wishbone_bd_ram_mem1_reg[235][14]/P0001 ,
		_w11936_,
		_w11982_,
		_w23750_
	);
	LUT4 #(
		.INIT('h0001)
	) name13238 (
		_w23747_,
		_w23748_,
		_w23749_,
		_w23750_,
		_w23751_
	);
	LUT3 #(
		.INIT('h80)
	) name13239 (
		\wishbone_bd_ram_mem1_reg[125][14]/P0001 ,
		_w11966_,
		_w12012_,
		_w23752_
	);
	LUT3 #(
		.INIT('h80)
	) name13240 (
		\wishbone_bd_ram_mem1_reg[219][14]/P0001 ,
		_w11936_,
		_w11984_,
		_w23753_
	);
	LUT3 #(
		.INIT('h80)
	) name13241 (
		\wishbone_bd_ram_mem1_reg[11][14]/P0001 ,
		_w11932_,
		_w11936_,
		_w23754_
	);
	LUT3 #(
		.INIT('h80)
	) name13242 (
		\wishbone_bd_ram_mem1_reg[36][14]/P0001 ,
		_w11929_,
		_w11957_,
		_w23755_
	);
	LUT4 #(
		.INIT('h0001)
	) name13243 (
		_w23752_,
		_w23753_,
		_w23754_,
		_w23755_,
		_w23756_
	);
	LUT4 #(
		.INIT('h8000)
	) name13244 (
		_w23741_,
		_w23746_,
		_w23751_,
		_w23756_,
		_w23757_
	);
	LUT3 #(
		.INIT('h80)
	) name13245 (
		\wishbone_bd_ram_mem1_reg[17][14]/P0001 ,
		_w11935_,
		_w11977_,
		_w23758_
	);
	LUT3 #(
		.INIT('h80)
	) name13246 (
		\wishbone_bd_ram_mem1_reg[25][14]/P0001 ,
		_w11935_,
		_w11968_,
		_w23759_
	);
	LUT3 #(
		.INIT('h80)
	) name13247 (
		\wishbone_bd_ram_mem1_reg[105][14]/P0001 ,
		_w11965_,
		_w11968_,
		_w23760_
	);
	LUT3 #(
		.INIT('h80)
	) name13248 (
		\wishbone_bd_ram_mem1_reg[234][14]/P0001 ,
		_w11944_,
		_w11982_,
		_w23761_
	);
	LUT4 #(
		.INIT('h0001)
	) name13249 (
		_w23758_,
		_w23759_,
		_w23760_,
		_w23761_,
		_w23762_
	);
	LUT3 #(
		.INIT('h80)
	) name13250 (
		\wishbone_bd_ram_mem1_reg[14][14]/P0001 ,
		_w11932_,
		_w11948_,
		_w23763_
	);
	LUT3 #(
		.INIT('h80)
	) name13251 (
		\wishbone_bd_ram_mem1_reg[93][14]/P0001 ,
		_w11966_,
		_w11972_,
		_w23764_
	);
	LUT3 #(
		.INIT('h80)
	) name13252 (
		\wishbone_bd_ram_mem1_reg[32][14]/P0001 ,
		_w11941_,
		_w11957_,
		_w23765_
	);
	LUT3 #(
		.INIT('h80)
	) name13253 (
		\wishbone_bd_ram_mem1_reg[215][14]/P0001 ,
		_w11975_,
		_w11984_,
		_w23766_
	);
	LUT4 #(
		.INIT('h0001)
	) name13254 (
		_w23763_,
		_w23764_,
		_w23765_,
		_w23766_,
		_w23767_
	);
	LUT3 #(
		.INIT('h80)
	) name13255 (
		\wishbone_bd_ram_mem1_reg[199][14]/P0001 ,
		_w11945_,
		_w11975_,
		_w23768_
	);
	LUT3 #(
		.INIT('h80)
	) name13256 (
		\wishbone_bd_ram_mem1_reg[133][14]/P0001 ,
		_w11933_,
		_w11955_,
		_w23769_
	);
	LUT3 #(
		.INIT('h80)
	) name13257 (
		\wishbone_bd_ram_mem1_reg[165][14]/P0001 ,
		_w11930_,
		_w11933_,
		_w23770_
	);
	LUT3 #(
		.INIT('h80)
	) name13258 (
		\wishbone_bd_ram_mem1_reg[169][14]/P0001 ,
		_w11930_,
		_w11968_,
		_w23771_
	);
	LUT4 #(
		.INIT('h0001)
	) name13259 (
		_w23768_,
		_w23769_,
		_w23770_,
		_w23771_,
		_w23772_
	);
	LUT3 #(
		.INIT('h80)
	) name13260 (
		\wishbone_bd_ram_mem1_reg[185][14]/P0001 ,
		_w11942_,
		_w11968_,
		_w23773_
	);
	LUT3 #(
		.INIT('h80)
	) name13261 (
		\wishbone_bd_ram_mem1_reg[129][14]/P0001 ,
		_w11955_,
		_w11977_,
		_w23774_
	);
	LUT3 #(
		.INIT('h80)
	) name13262 (
		\wishbone_bd_ram_mem1_reg[240][14]/P0001 ,
		_w11941_,
		_w11952_,
		_w23775_
	);
	LUT3 #(
		.INIT('h80)
	) name13263 (
		\wishbone_bd_ram_mem1_reg[175][14]/P0001 ,
		_w11930_,
		_w11973_,
		_w23776_
	);
	LUT4 #(
		.INIT('h0001)
	) name13264 (
		_w23773_,
		_w23774_,
		_w23775_,
		_w23776_,
		_w23777_
	);
	LUT4 #(
		.INIT('h8000)
	) name13265 (
		_w23762_,
		_w23767_,
		_w23772_,
		_w23777_,
		_w23778_
	);
	LUT4 #(
		.INIT('h8000)
	) name13266 (
		_w23715_,
		_w23736_,
		_w23757_,
		_w23778_,
		_w23779_
	);
	LUT3 #(
		.INIT('h80)
	) name13267 (
		\wishbone_bd_ram_mem1_reg[38][14]/P0001 ,
		_w11957_,
		_w11986_,
		_w23780_
	);
	LUT3 #(
		.INIT('h80)
	) name13268 (
		\wishbone_bd_ram_mem1_reg[119][14]/P0001 ,
		_w11975_,
		_w12012_,
		_w23781_
	);
	LUT3 #(
		.INIT('h80)
	) name13269 (
		\wishbone_bd_ram_mem1_reg[163][14]/P0001 ,
		_w11930_,
		_w11938_,
		_w23782_
	);
	LUT3 #(
		.INIT('h80)
	) name13270 (
		\wishbone_bd_ram_mem1_reg[251][14]/P0001 ,
		_w11936_,
		_w11952_,
		_w23783_
	);
	LUT4 #(
		.INIT('h0001)
	) name13271 (
		_w23780_,
		_w23781_,
		_w23782_,
		_w23783_,
		_w23784_
	);
	LUT3 #(
		.INIT('h80)
	) name13272 (
		\wishbone_bd_ram_mem1_reg[161][14]/P0001 ,
		_w11930_,
		_w11977_,
		_w23785_
	);
	LUT3 #(
		.INIT('h80)
	) name13273 (
		\wishbone_bd_ram_mem1_reg[153][14]/P0001 ,
		_w11959_,
		_w11968_,
		_w23786_
	);
	LUT3 #(
		.INIT('h80)
	) name13274 (
		\wishbone_bd_ram_mem1_reg[84][14]/P0001 ,
		_w11929_,
		_w11972_,
		_w23787_
	);
	LUT3 #(
		.INIT('h80)
	) name13275 (
		\wishbone_bd_ram_mem1_reg[6][14]/P0001 ,
		_w11932_,
		_w11986_,
		_w23788_
	);
	LUT4 #(
		.INIT('h0001)
	) name13276 (
		_w23785_,
		_w23786_,
		_w23787_,
		_w23788_,
		_w23789_
	);
	LUT3 #(
		.INIT('h80)
	) name13277 (
		\wishbone_bd_ram_mem1_reg[180][14]/P0001 ,
		_w11929_,
		_w11942_,
		_w23790_
	);
	LUT3 #(
		.INIT('h80)
	) name13278 (
		\wishbone_bd_ram_mem1_reg[173][14]/P0001 ,
		_w11930_,
		_w11966_,
		_w23791_
	);
	LUT3 #(
		.INIT('h80)
	) name13279 (
		\wishbone_bd_ram_mem1_reg[191][14]/P0001 ,
		_w11942_,
		_w11973_,
		_w23792_
	);
	LUT3 #(
		.INIT('h80)
	) name13280 (
		\wishbone_bd_ram_mem1_reg[19][14]/P0001 ,
		_w11935_,
		_w11938_,
		_w23793_
	);
	LUT4 #(
		.INIT('h0001)
	) name13281 (
		_w23790_,
		_w23791_,
		_w23792_,
		_w23793_,
		_w23794_
	);
	LUT3 #(
		.INIT('h80)
	) name13282 (
		\wishbone_bd_ram_mem1_reg[80][14]/P0001 ,
		_w11941_,
		_w11972_,
		_w23795_
	);
	LUT3 #(
		.INIT('h80)
	) name13283 (
		\wishbone_bd_ram_mem1_reg[34][14]/P0001 ,
		_w11957_,
		_w11963_,
		_w23796_
	);
	LUT3 #(
		.INIT('h80)
	) name13284 (
		\wishbone_bd_ram_mem1_reg[92][14]/P0001 ,
		_w11954_,
		_w11972_,
		_w23797_
	);
	LUT3 #(
		.INIT('h80)
	) name13285 (
		\wishbone_bd_ram_mem1_reg[188][14]/P0001 ,
		_w11942_,
		_w11954_,
		_w23798_
	);
	LUT4 #(
		.INIT('h0001)
	) name13286 (
		_w23795_,
		_w23796_,
		_w23797_,
		_w23798_,
		_w23799_
	);
	LUT4 #(
		.INIT('h8000)
	) name13287 (
		_w23784_,
		_w23789_,
		_w23794_,
		_w23799_,
		_w23800_
	);
	LUT3 #(
		.INIT('h80)
	) name13288 (
		\wishbone_bd_ram_mem1_reg[213][14]/P0001 ,
		_w11933_,
		_w11984_,
		_w23801_
	);
	LUT3 #(
		.INIT('h80)
	) name13289 (
		\wishbone_bd_ram_mem1_reg[144][14]/P0001 ,
		_w11941_,
		_w11959_,
		_w23802_
	);
	LUT3 #(
		.INIT('h80)
	) name13290 (
		\wishbone_bd_ram_mem1_reg[42][14]/P0001 ,
		_w11944_,
		_w11957_,
		_w23803_
	);
	LUT3 #(
		.INIT('h80)
	) name13291 (
		\wishbone_bd_ram_mem1_reg[64][14]/P0001 ,
		_w11941_,
		_w11949_,
		_w23804_
	);
	LUT4 #(
		.INIT('h0001)
	) name13292 (
		_w23801_,
		_w23802_,
		_w23803_,
		_w23804_,
		_w23805_
	);
	LUT3 #(
		.INIT('h80)
	) name13293 (
		\wishbone_bd_ram_mem1_reg[91][14]/P0001 ,
		_w11936_,
		_w11972_,
		_w23806_
	);
	LUT3 #(
		.INIT('h80)
	) name13294 (
		\wishbone_bd_ram_mem1_reg[71][14]/P0001 ,
		_w11949_,
		_w11975_,
		_w23807_
	);
	LUT3 #(
		.INIT('h80)
	) name13295 (
		\wishbone_bd_ram_mem1_reg[7][14]/P0001 ,
		_w11932_,
		_w11975_,
		_w23808_
	);
	LUT3 #(
		.INIT('h80)
	) name13296 (
		\wishbone_bd_ram_mem1_reg[186][14]/P0001 ,
		_w11942_,
		_w11944_,
		_w23809_
	);
	LUT4 #(
		.INIT('h0001)
	) name13297 (
		_w23806_,
		_w23807_,
		_w23808_,
		_w23809_,
		_w23810_
	);
	LUT3 #(
		.INIT('h80)
	) name13298 (
		\wishbone_bd_ram_mem1_reg[236][14]/P0001 ,
		_w11954_,
		_w11982_,
		_w23811_
	);
	LUT3 #(
		.INIT('h80)
	) name13299 (
		\wishbone_bd_ram_mem1_reg[96][14]/P0001 ,
		_w11941_,
		_w11965_,
		_w23812_
	);
	LUT3 #(
		.INIT('h80)
	) name13300 (
		\wishbone_bd_ram_mem1_reg[55][14]/P0001 ,
		_w11975_,
		_w11979_,
		_w23813_
	);
	LUT3 #(
		.INIT('h80)
	) name13301 (
		\wishbone_bd_ram_mem1_reg[252][14]/P0001 ,
		_w11952_,
		_w11954_,
		_w23814_
	);
	LUT4 #(
		.INIT('h0001)
	) name13302 (
		_w23811_,
		_w23812_,
		_w23813_,
		_w23814_,
		_w23815_
	);
	LUT3 #(
		.INIT('h80)
	) name13303 (
		\wishbone_bd_ram_mem1_reg[254][14]/P0001 ,
		_w11948_,
		_w11952_,
		_w23816_
	);
	LUT3 #(
		.INIT('h80)
	) name13304 (
		\wishbone_bd_ram_mem1_reg[139][14]/P0001 ,
		_w11936_,
		_w11955_,
		_w23817_
	);
	LUT3 #(
		.INIT('h80)
	) name13305 (
		\wishbone_bd_ram_mem1_reg[109][14]/P0001 ,
		_w11965_,
		_w11966_,
		_w23818_
	);
	LUT3 #(
		.INIT('h80)
	) name13306 (
		\wishbone_bd_ram_mem1_reg[10][14]/P0001 ,
		_w11932_,
		_w11944_,
		_w23819_
	);
	LUT4 #(
		.INIT('h0001)
	) name13307 (
		_w23816_,
		_w23817_,
		_w23818_,
		_w23819_,
		_w23820_
	);
	LUT4 #(
		.INIT('h8000)
	) name13308 (
		_w23805_,
		_w23810_,
		_w23815_,
		_w23820_,
		_w23821_
	);
	LUT3 #(
		.INIT('h80)
	) name13309 (
		\wishbone_bd_ram_mem1_reg[249][14]/P0001 ,
		_w11952_,
		_w11968_,
		_w23822_
	);
	LUT3 #(
		.INIT('h80)
	) name13310 (
		\wishbone_bd_ram_mem1_reg[15][14]/P0001 ,
		_w11932_,
		_w11973_,
		_w23823_
	);
	LUT3 #(
		.INIT('h80)
	) name13311 (
		\wishbone_bd_ram_mem1_reg[52][14]/P0001 ,
		_w11929_,
		_w11979_,
		_w23824_
	);
	LUT3 #(
		.INIT('h80)
	) name13312 (
		\wishbone_bd_ram_mem1_reg[179][14]/P0001 ,
		_w11938_,
		_w11942_,
		_w23825_
	);
	LUT4 #(
		.INIT('h0001)
	) name13313 (
		_w23822_,
		_w23823_,
		_w23824_,
		_w23825_,
		_w23826_
	);
	LUT3 #(
		.INIT('h80)
	) name13314 (
		\wishbone_bd_ram_mem1_reg[201][14]/P0001 ,
		_w11945_,
		_w11968_,
		_w23827_
	);
	LUT3 #(
		.INIT('h80)
	) name13315 (
		\wishbone_bd_ram_mem1_reg[61][14]/P0001 ,
		_w11966_,
		_w11979_,
		_w23828_
	);
	LUT3 #(
		.INIT('h80)
	) name13316 (
		\wishbone_bd_ram_mem1_reg[245][14]/P0001 ,
		_w11933_,
		_w11952_,
		_w23829_
	);
	LUT3 #(
		.INIT('h80)
	) name13317 (
		\wishbone_bd_ram_mem1_reg[193][14]/P0001 ,
		_w11945_,
		_w11977_,
		_w23830_
	);
	LUT4 #(
		.INIT('h0001)
	) name13318 (
		_w23827_,
		_w23828_,
		_w23829_,
		_w23830_,
		_w23831_
	);
	LUT3 #(
		.INIT('h80)
	) name13319 (
		\wishbone_bd_ram_mem1_reg[62][14]/P0001 ,
		_w11948_,
		_w11979_,
		_w23832_
	);
	LUT3 #(
		.INIT('h80)
	) name13320 (
		\wishbone_bd_ram_mem1_reg[196][14]/P0001 ,
		_w11929_,
		_w11945_,
		_w23833_
	);
	LUT3 #(
		.INIT('h80)
	) name13321 (
		\wishbone_bd_ram_mem1_reg[30][14]/P0001 ,
		_w11935_,
		_w11948_,
		_w23834_
	);
	LUT3 #(
		.INIT('h80)
	) name13322 (
		\wishbone_bd_ram_mem1_reg[128][14]/P0001 ,
		_w11941_,
		_w11955_,
		_w23835_
	);
	LUT4 #(
		.INIT('h0001)
	) name13323 (
		_w23832_,
		_w23833_,
		_w23834_,
		_w23835_,
		_w23836_
	);
	LUT3 #(
		.INIT('h80)
	) name13324 (
		\wishbone_bd_ram_mem1_reg[24][14]/P0001 ,
		_w11935_,
		_w11990_,
		_w23837_
	);
	LUT3 #(
		.INIT('h80)
	) name13325 (
		\wishbone_bd_ram_mem1_reg[88][14]/P0001 ,
		_w11972_,
		_w11990_,
		_w23838_
	);
	LUT3 #(
		.INIT('h80)
	) name13326 (
		\wishbone_bd_ram_mem1_reg[115][14]/P0001 ,
		_w11938_,
		_w12012_,
		_w23839_
	);
	LUT3 #(
		.INIT('h80)
	) name13327 (
		\wishbone_bd_ram_mem1_reg[97][14]/P0001 ,
		_w11965_,
		_w11977_,
		_w23840_
	);
	LUT4 #(
		.INIT('h0001)
	) name13328 (
		_w23837_,
		_w23838_,
		_w23839_,
		_w23840_,
		_w23841_
	);
	LUT4 #(
		.INIT('h8000)
	) name13329 (
		_w23826_,
		_w23831_,
		_w23836_,
		_w23841_,
		_w23842_
	);
	LUT3 #(
		.INIT('h80)
	) name13330 (
		\wishbone_bd_ram_mem1_reg[151][14]/P0001 ,
		_w11959_,
		_w11975_,
		_w23843_
	);
	LUT3 #(
		.INIT('h80)
	) name13331 (
		\wishbone_bd_ram_mem1_reg[39][14]/P0001 ,
		_w11957_,
		_w11975_,
		_w23844_
	);
	LUT3 #(
		.INIT('h80)
	) name13332 (
		\wishbone_bd_ram_mem1_reg[152][14]/P0001 ,
		_w11959_,
		_w11990_,
		_w23845_
	);
	LUT3 #(
		.INIT('h80)
	) name13333 (
		\wishbone_bd_ram_mem1_reg[48][14]/P0001 ,
		_w11941_,
		_w11979_,
		_w23846_
	);
	LUT4 #(
		.INIT('h0001)
	) name13334 (
		_w23843_,
		_w23844_,
		_w23845_,
		_w23846_,
		_w23847_
	);
	LUT3 #(
		.INIT('h80)
	) name13335 (
		\wishbone_bd_ram_mem1_reg[145][14]/P0001 ,
		_w11959_,
		_w11977_,
		_w23848_
	);
	LUT3 #(
		.INIT('h80)
	) name13336 (
		\wishbone_bd_ram_mem1_reg[192][14]/P0001 ,
		_w11941_,
		_w11945_,
		_w23849_
	);
	LUT3 #(
		.INIT('h80)
	) name13337 (
		\wishbone_bd_ram_mem1_reg[51][14]/P0001 ,
		_w11938_,
		_w11979_,
		_w23850_
	);
	LUT3 #(
		.INIT('h80)
	) name13338 (
		\wishbone_bd_ram_mem1_reg[200][14]/P0001 ,
		_w11945_,
		_w11990_,
		_w23851_
	);
	LUT4 #(
		.INIT('h0001)
	) name13339 (
		_w23848_,
		_w23849_,
		_w23850_,
		_w23851_,
		_w23852_
	);
	LUT3 #(
		.INIT('h80)
	) name13340 (
		\wishbone_bd_ram_mem1_reg[187][14]/P0001 ,
		_w11936_,
		_w11942_,
		_w23853_
	);
	LUT3 #(
		.INIT('h80)
	) name13341 (
		\wishbone_bd_ram_mem1_reg[20][14]/P0001 ,
		_w11929_,
		_w11935_,
		_w23854_
	);
	LUT3 #(
		.INIT('h80)
	) name13342 (
		\wishbone_bd_ram_mem1_reg[136][14]/P0001 ,
		_w11955_,
		_w11990_,
		_w23855_
	);
	LUT3 #(
		.INIT('h80)
	) name13343 (
		\wishbone_bd_ram_mem1_reg[110][14]/P0001 ,
		_w11948_,
		_w11965_,
		_w23856_
	);
	LUT4 #(
		.INIT('h0001)
	) name13344 (
		_w23853_,
		_w23854_,
		_w23855_,
		_w23856_,
		_w23857_
	);
	LUT3 #(
		.INIT('h80)
	) name13345 (
		\wishbone_bd_ram_mem1_reg[225][14]/P0001 ,
		_w11977_,
		_w11982_,
		_w23858_
	);
	LUT3 #(
		.INIT('h80)
	) name13346 (
		\wishbone_bd_ram_mem1_reg[3][14]/P0001 ,
		_w11932_,
		_w11938_,
		_w23859_
	);
	LUT3 #(
		.INIT('h80)
	) name13347 (
		\wishbone_bd_ram_mem1_reg[47][14]/P0001 ,
		_w11957_,
		_w11973_,
		_w23860_
	);
	LUT3 #(
		.INIT('h80)
	) name13348 (
		\wishbone_bd_ram_mem1_reg[120][14]/P0001 ,
		_w11990_,
		_w12012_,
		_w23861_
	);
	LUT4 #(
		.INIT('h0001)
	) name13349 (
		_w23858_,
		_w23859_,
		_w23860_,
		_w23861_,
		_w23862_
	);
	LUT4 #(
		.INIT('h8000)
	) name13350 (
		_w23847_,
		_w23852_,
		_w23857_,
		_w23862_,
		_w23863_
	);
	LUT4 #(
		.INIT('h8000)
	) name13351 (
		_w23800_,
		_w23821_,
		_w23842_,
		_w23863_,
		_w23864_
	);
	LUT3 #(
		.INIT('h80)
	) name13352 (
		\wishbone_bd_ram_mem1_reg[49][14]/P0001 ,
		_w11977_,
		_w11979_,
		_w23865_
	);
	LUT3 #(
		.INIT('h80)
	) name13353 (
		\wishbone_bd_ram_mem1_reg[184][14]/P0001 ,
		_w11942_,
		_w11990_,
		_w23866_
	);
	LUT3 #(
		.INIT('h80)
	) name13354 (
		\wishbone_bd_ram_mem1_reg[82][14]/P0001 ,
		_w11963_,
		_w11972_,
		_w23867_
	);
	LUT3 #(
		.INIT('h80)
	) name13355 (
		\wishbone_bd_ram_mem1_reg[142][14]/P0001 ,
		_w11948_,
		_w11955_,
		_w23868_
	);
	LUT4 #(
		.INIT('h0001)
	) name13356 (
		_w23865_,
		_w23866_,
		_w23867_,
		_w23868_,
		_w23869_
	);
	LUT3 #(
		.INIT('h80)
	) name13357 (
		\wishbone_bd_ram_mem1_reg[77][14]/P0001 ,
		_w11949_,
		_w11966_,
		_w23870_
	);
	LUT3 #(
		.INIT('h80)
	) name13358 (
		\wishbone_bd_ram_mem1_reg[22][14]/P0001 ,
		_w11935_,
		_w11986_,
		_w23871_
	);
	LUT3 #(
		.INIT('h80)
	) name13359 (
		\wishbone_bd_ram_mem1_reg[21][14]/P0001 ,
		_w11933_,
		_w11935_,
		_w23872_
	);
	LUT3 #(
		.INIT('h80)
	) name13360 (
		\wishbone_bd_ram_mem1_reg[227][14]/P0001 ,
		_w11938_,
		_w11982_,
		_w23873_
	);
	LUT4 #(
		.INIT('h0001)
	) name13361 (
		_w23870_,
		_w23871_,
		_w23872_,
		_w23873_,
		_w23874_
	);
	LUT3 #(
		.INIT('h80)
	) name13362 (
		\wishbone_bd_ram_mem1_reg[167][14]/P0001 ,
		_w11930_,
		_w11975_,
		_w23875_
	);
	LUT3 #(
		.INIT('h80)
	) name13363 (
		\wishbone_bd_ram_mem1_reg[226][14]/P0001 ,
		_w11963_,
		_w11982_,
		_w23876_
	);
	LUT3 #(
		.INIT('h80)
	) name13364 (
		\wishbone_bd_ram_mem1_reg[83][14]/P0001 ,
		_w11938_,
		_w11972_,
		_w23877_
	);
	LUT3 #(
		.INIT('h80)
	) name13365 (
		\wishbone_bd_ram_mem1_reg[127][14]/P0001 ,
		_w11973_,
		_w12012_,
		_w23878_
	);
	LUT4 #(
		.INIT('h0001)
	) name13366 (
		_w23875_,
		_w23876_,
		_w23877_,
		_w23878_,
		_w23879_
	);
	LUT3 #(
		.INIT('h80)
	) name13367 (
		\wishbone_bd_ram_mem1_reg[162][14]/P0001 ,
		_w11930_,
		_w11963_,
		_w23880_
	);
	LUT3 #(
		.INIT('h80)
	) name13368 (
		\wishbone_bd_ram_mem1_reg[37][14]/P0001 ,
		_w11933_,
		_w11957_,
		_w23881_
	);
	LUT3 #(
		.INIT('h80)
	) name13369 (
		\wishbone_bd_ram_mem1_reg[23][14]/P0001 ,
		_w11935_,
		_w11975_,
		_w23882_
	);
	LUT3 #(
		.INIT('h80)
	) name13370 (
		\wishbone_bd_ram_mem1_reg[57][14]/P0001 ,
		_w11968_,
		_w11979_,
		_w23883_
	);
	LUT4 #(
		.INIT('h0001)
	) name13371 (
		_w23880_,
		_w23881_,
		_w23882_,
		_w23883_,
		_w23884_
	);
	LUT4 #(
		.INIT('h8000)
	) name13372 (
		_w23869_,
		_w23874_,
		_w23879_,
		_w23884_,
		_w23885_
	);
	LUT3 #(
		.INIT('h80)
	) name13373 (
		\wishbone_bd_ram_mem1_reg[143][14]/P0001 ,
		_w11955_,
		_w11973_,
		_w23886_
	);
	LUT3 #(
		.INIT('h80)
	) name13374 (
		\wishbone_bd_ram_mem1_reg[154][14]/P0001 ,
		_w11944_,
		_w11959_,
		_w23887_
	);
	LUT3 #(
		.INIT('h80)
	) name13375 (
		\wishbone_bd_ram_mem1_reg[130][14]/P0001 ,
		_w11955_,
		_w11963_,
		_w23888_
	);
	LUT3 #(
		.INIT('h80)
	) name13376 (
		\wishbone_bd_ram_mem1_reg[103][14]/P0001 ,
		_w11965_,
		_w11975_,
		_w23889_
	);
	LUT4 #(
		.INIT('h0001)
	) name13377 (
		_w23886_,
		_w23887_,
		_w23888_,
		_w23889_,
		_w23890_
	);
	LUT3 #(
		.INIT('h80)
	) name13378 (
		\wishbone_bd_ram_mem1_reg[149][14]/P0001 ,
		_w11933_,
		_w11959_,
		_w23891_
	);
	LUT3 #(
		.INIT('h80)
	) name13379 (
		\wishbone_bd_ram_mem1_reg[35][14]/P0001 ,
		_w11938_,
		_w11957_,
		_w23892_
	);
	LUT3 #(
		.INIT('h80)
	) name13380 (
		\wishbone_bd_ram_mem1_reg[147][14]/P0001 ,
		_w11938_,
		_w11959_,
		_w23893_
	);
	LUT3 #(
		.INIT('h80)
	) name13381 (
		\wishbone_bd_ram_mem1_reg[159][14]/P0001 ,
		_w11959_,
		_w11973_,
		_w23894_
	);
	LUT4 #(
		.INIT('h0001)
	) name13382 (
		_w23891_,
		_w23892_,
		_w23893_,
		_w23894_,
		_w23895_
	);
	LUT3 #(
		.INIT('h80)
	) name13383 (
		\wishbone_bd_ram_mem1_reg[250][14]/P0001 ,
		_w11944_,
		_w11952_,
		_w23896_
	);
	LUT3 #(
		.INIT('h80)
	) name13384 (
		\wishbone_bd_ram_mem1_reg[79][14]/P0001 ,
		_w11949_,
		_w11973_,
		_w23897_
	);
	LUT3 #(
		.INIT('h80)
	) name13385 (
		\wishbone_bd_ram_mem1_reg[74][14]/P0001 ,
		_w11944_,
		_w11949_,
		_w23898_
	);
	LUT3 #(
		.INIT('h80)
	) name13386 (
		\wishbone_bd_ram_mem1_reg[160][14]/P0001 ,
		_w11930_,
		_w11941_,
		_w23899_
	);
	LUT4 #(
		.INIT('h0001)
	) name13387 (
		_w23896_,
		_w23897_,
		_w23898_,
		_w23899_,
		_w23900_
	);
	LUT3 #(
		.INIT('h80)
	) name13388 (
		\wishbone_bd_ram_mem1_reg[102][14]/P0001 ,
		_w11965_,
		_w11986_,
		_w23901_
	);
	LUT3 #(
		.INIT('h80)
	) name13389 (
		\wishbone_bd_ram_mem1_reg[141][14]/P0001 ,
		_w11955_,
		_w11966_,
		_w23902_
	);
	LUT3 #(
		.INIT('h80)
	) name13390 (
		\wishbone_bd_ram_mem1_reg[239][14]/P0001 ,
		_w11973_,
		_w11982_,
		_w23903_
	);
	LUT3 #(
		.INIT('h80)
	) name13391 (
		\wishbone_bd_ram_mem1_reg[63][14]/P0001 ,
		_w11973_,
		_w11979_,
		_w23904_
	);
	LUT4 #(
		.INIT('h0001)
	) name13392 (
		_w23901_,
		_w23902_,
		_w23903_,
		_w23904_,
		_w23905_
	);
	LUT4 #(
		.INIT('h8000)
	) name13393 (
		_w23890_,
		_w23895_,
		_w23900_,
		_w23905_,
		_w23906_
	);
	LUT3 #(
		.INIT('h80)
	) name13394 (
		\wishbone_bd_ram_mem1_reg[26][14]/P0001 ,
		_w11935_,
		_w11944_,
		_w23907_
	);
	LUT3 #(
		.INIT('h80)
	) name13395 (
		\wishbone_bd_ram_mem1_reg[9][14]/P0001 ,
		_w11932_,
		_w11968_,
		_w23908_
	);
	LUT3 #(
		.INIT('h80)
	) name13396 (
		\wishbone_bd_ram_mem1_reg[89][14]/P0001 ,
		_w11968_,
		_w11972_,
		_w23909_
	);
	LUT3 #(
		.INIT('h80)
	) name13397 (
		\wishbone_bd_ram_mem1_reg[150][14]/P0001 ,
		_w11959_,
		_w11986_,
		_w23910_
	);
	LUT4 #(
		.INIT('h0001)
	) name13398 (
		_w23907_,
		_w23908_,
		_w23909_,
		_w23910_,
		_w23911_
	);
	LUT3 #(
		.INIT('h80)
	) name13399 (
		\wishbone_bd_ram_mem1_reg[104][14]/P0001 ,
		_w11965_,
		_w11990_,
		_w23912_
	);
	LUT3 #(
		.INIT('h80)
	) name13400 (
		\wishbone_bd_ram_mem1_reg[99][14]/P0001 ,
		_w11938_,
		_w11965_,
		_w23913_
	);
	LUT3 #(
		.INIT('h80)
	) name13401 (
		\wishbone_bd_ram_mem1_reg[208][14]/P0001 ,
		_w11941_,
		_w11984_,
		_w23914_
	);
	LUT3 #(
		.INIT('h80)
	) name13402 (
		\wishbone_bd_ram_mem1_reg[166][14]/P0001 ,
		_w11930_,
		_w11986_,
		_w23915_
	);
	LUT4 #(
		.INIT('h0001)
	) name13403 (
		_w23912_,
		_w23913_,
		_w23914_,
		_w23915_,
		_w23916_
	);
	LUT3 #(
		.INIT('h80)
	) name13404 (
		\wishbone_bd_ram_mem1_reg[5][14]/P0001 ,
		_w11932_,
		_w11933_,
		_w23917_
	);
	LUT3 #(
		.INIT('h80)
	) name13405 (
		\wishbone_bd_ram_mem1_reg[229][14]/P0001 ,
		_w11933_,
		_w11982_,
		_w23918_
	);
	LUT3 #(
		.INIT('h80)
	) name13406 (
		\wishbone_bd_ram_mem1_reg[182][14]/P0001 ,
		_w11942_,
		_w11986_,
		_w23919_
	);
	LUT3 #(
		.INIT('h80)
	) name13407 (
		\wishbone_bd_ram_mem1_reg[94][14]/P0001 ,
		_w11948_,
		_w11972_,
		_w23920_
	);
	LUT4 #(
		.INIT('h0001)
	) name13408 (
		_w23917_,
		_w23918_,
		_w23919_,
		_w23920_,
		_w23921_
	);
	LUT3 #(
		.INIT('h80)
	) name13409 (
		\wishbone_bd_ram_mem1_reg[117][14]/P0001 ,
		_w11933_,
		_w12012_,
		_w23922_
	);
	LUT3 #(
		.INIT('h80)
	) name13410 (
		\wishbone_bd_ram_mem1_reg[67][14]/P0001 ,
		_w11938_,
		_w11949_,
		_w23923_
	);
	LUT3 #(
		.INIT('h80)
	) name13411 (
		\wishbone_bd_ram_mem1_reg[246][14]/P0001 ,
		_w11952_,
		_w11986_,
		_w23924_
	);
	LUT3 #(
		.INIT('h80)
	) name13412 (
		\wishbone_bd_ram_mem1_reg[111][14]/P0001 ,
		_w11965_,
		_w11973_,
		_w23925_
	);
	LUT4 #(
		.INIT('h0001)
	) name13413 (
		_w23922_,
		_w23923_,
		_w23924_,
		_w23925_,
		_w23926_
	);
	LUT4 #(
		.INIT('h8000)
	) name13414 (
		_w23911_,
		_w23916_,
		_w23921_,
		_w23926_,
		_w23927_
	);
	LUT3 #(
		.INIT('h80)
	) name13415 (
		\wishbone_bd_ram_mem1_reg[174][14]/P0001 ,
		_w11930_,
		_w11948_,
		_w23928_
	);
	LUT3 #(
		.INIT('h80)
	) name13416 (
		\wishbone_bd_ram_mem1_reg[244][14]/P0001 ,
		_w11929_,
		_w11952_,
		_w23929_
	);
	LUT3 #(
		.INIT('h80)
	) name13417 (
		\wishbone_bd_ram_mem1_reg[40][14]/P0001 ,
		_w11957_,
		_w11990_,
		_w23930_
	);
	LUT3 #(
		.INIT('h80)
	) name13418 (
		\wishbone_bd_ram_mem1_reg[90][14]/P0001 ,
		_w11944_,
		_w11972_,
		_w23931_
	);
	LUT4 #(
		.INIT('h0001)
	) name13419 (
		_w23928_,
		_w23929_,
		_w23930_,
		_w23931_,
		_w23932_
	);
	LUT3 #(
		.INIT('h80)
	) name13420 (
		\wishbone_bd_ram_mem1_reg[100][14]/P0001 ,
		_w11929_,
		_w11965_,
		_w23933_
	);
	LUT3 #(
		.INIT('h80)
	) name13421 (
		\wishbone_bd_ram_mem1_reg[60][14]/P0001 ,
		_w11954_,
		_w11979_,
		_w23934_
	);
	LUT3 #(
		.INIT('h80)
	) name13422 (
		\wishbone_bd_ram_mem1_reg[168][14]/P0001 ,
		_w11930_,
		_w11990_,
		_w23935_
	);
	LUT3 #(
		.INIT('h80)
	) name13423 (
		\wishbone_bd_ram_mem1_reg[106][14]/P0001 ,
		_w11944_,
		_w11965_,
		_w23936_
	);
	LUT4 #(
		.INIT('h0001)
	) name13424 (
		_w23933_,
		_w23934_,
		_w23935_,
		_w23936_,
		_w23937_
	);
	LUT3 #(
		.INIT('h80)
	) name13425 (
		\wishbone_bd_ram_mem1_reg[124][14]/P0001 ,
		_w11954_,
		_w12012_,
		_w23938_
	);
	LUT3 #(
		.INIT('h80)
	) name13426 (
		\wishbone_bd_ram_mem1_reg[181][14]/P0001 ,
		_w11933_,
		_w11942_,
		_w23939_
	);
	LUT3 #(
		.INIT('h80)
	) name13427 (
		\wishbone_bd_ram_mem1_reg[228][14]/P0001 ,
		_w11929_,
		_w11982_,
		_w23940_
	);
	LUT3 #(
		.INIT('h80)
	) name13428 (
		\wishbone_bd_ram_mem1_reg[122][14]/P0001 ,
		_w11944_,
		_w12012_,
		_w23941_
	);
	LUT4 #(
		.INIT('h0001)
	) name13429 (
		_w23938_,
		_w23939_,
		_w23940_,
		_w23941_,
		_w23942_
	);
	LUT3 #(
		.INIT('h80)
	) name13430 (
		\wishbone_bd_ram_mem1_reg[158][14]/P0001 ,
		_w11948_,
		_w11959_,
		_w23943_
	);
	LUT3 #(
		.INIT('h80)
	) name13431 (
		\wishbone_bd_ram_mem1_reg[59][14]/P0001 ,
		_w11936_,
		_w11979_,
		_w23944_
	);
	LUT3 #(
		.INIT('h80)
	) name13432 (
		\wishbone_bd_ram_mem1_reg[65][14]/P0001 ,
		_w11949_,
		_w11977_,
		_w23945_
	);
	LUT3 #(
		.INIT('h80)
	) name13433 (
		\wishbone_bd_ram_mem1_reg[86][14]/P0001 ,
		_w11972_,
		_w11986_,
		_w23946_
	);
	LUT4 #(
		.INIT('h0001)
	) name13434 (
		_w23943_,
		_w23944_,
		_w23945_,
		_w23946_,
		_w23947_
	);
	LUT4 #(
		.INIT('h8000)
	) name13435 (
		_w23932_,
		_w23937_,
		_w23942_,
		_w23947_,
		_w23948_
	);
	LUT4 #(
		.INIT('h8000)
	) name13436 (
		_w23885_,
		_w23906_,
		_w23927_,
		_w23948_,
		_w23949_
	);
	LUT4 #(
		.INIT('h8000)
	) name13437 (
		_w23694_,
		_w23779_,
		_w23864_,
		_w23949_,
		_w23950_
	);
	LUT2 #(
		.INIT('h1)
	) name13438 (
		wb_rst_i_pad,
		_w23608_,
		_w23951_
	);
	LUT3 #(
		.INIT('hba)
	) name13439 (
		_w23609_,
		_w23950_,
		_w23951_,
		_w23952_
	);
	LUT3 #(
		.INIT('h80)
	) name13440 (
		\ethreg1_MODER_1_DataOut_reg[7]/NET0131 ,
		_w18800_,
		_w18801_,
		_w23953_
	);
	LUT4 #(
		.INIT('h0020)
	) name13441 (
		\ethreg1_TXCTRL_1_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23954_
	);
	LUT3 #(
		.INIT('h80)
	) name13442 (
		_w18757_,
		_w18758_,
		_w23954_,
		_w23955_
	);
	LUT4 #(
		.INIT('h0008)
	) name13443 (
		\ethreg1_RXHASH0_1_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23956_
	);
	LUT3 #(
		.INIT('h80)
	) name13444 (
		_w18757_,
		_w18758_,
		_w23956_,
		_w23957_
	);
	LUT4 #(
		.INIT('h0008)
	) name13445 (
		\ethreg1_RXHASH1_1_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23958_
	);
	LUT3 #(
		.INIT('h80)
	) name13446 (
		_w18757_,
		_w18762_,
		_w23958_,
		_w23959_
	);
	LUT4 #(
		.INIT('h0001)
	) name13447 (
		_w23953_,
		_w23955_,
		_w23957_,
		_w23959_,
		_w23960_
	);
	LUT3 #(
		.INIT('h80)
	) name13448 (
		\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131 ,
		_w18753_,
		_w18754_,
		_w23961_
	);
	LUT3 #(
		.INIT('h80)
	) name13449 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[7]/NET0131 ,
		_w18798_,
		_w18805_,
		_w23962_
	);
	LUT4 #(
		.INIT('h0002)
	) name13450 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23963_
	);
	LUT3 #(
		.INIT('h80)
	) name13451 (
		_w18757_,
		_w18758_,
		_w23963_,
		_w23964_
	);
	LUT4 #(
		.INIT('h0002)
	) name13452 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w23965_
	);
	LUT3 #(
		.INIT('h80)
	) name13453 (
		_w18757_,
		_w18762_,
		_w23965_,
		_w23966_
	);
	LUT3 #(
		.INIT('h80)
	) name13454 (
		\ethreg1_MIIRX_DATA_DataOut_reg[15]/NET0131 ,
		_w18785_,
		_w18786_,
		_w23967_
	);
	LUT4 #(
		.INIT('h0001)
	) name13455 (
		_w23962_,
		_w23964_,
		_w23966_,
		_w23967_,
		_w23968_
	);
	LUT4 #(
		.INIT('h0800)
	) name13456 (
		_w18752_,
		_w23960_,
		_w23961_,
		_w23968_,
		_w23969_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name13457 (
		_w18752_,
		_w23960_,
		_w23961_,
		_w23968_,
		_w23970_
	);
	LUT2 #(
		.INIT('h1)
	) name13458 (
		wb_rst_i_pad,
		_w23969_,
		_w23971_
	);
	LUT3 #(
		.INIT('hdc)
	) name13459 (
		_w13800_,
		_w23970_,
		_w23971_,
		_w23972_
	);
	LUT2 #(
		.INIT('h8)
	) name13460 (
		\wishbone_RxPointerMSB_reg[11]/NET0131 ,
		\wishbone_RxPointerMSB_reg[12]/NET0131 ,
		_w23973_
	);
	LUT4 #(
		.INIT('h8000)
	) name13461 (
		_w15283_,
		_w15284_,
		_w15285_,
		_w23973_,
		_w23974_
	);
	LUT4 #(
		.INIT('h060c)
	) name13462 (
		\wishbone_RxPointerMSB_reg[11]/NET0131 ,
		\wishbone_RxPointerMSB_reg[12]/NET0131 ,
		_w13807_,
		_w15286_,
		_w23975_
	);
	LUT3 #(
		.INIT('hf2)
	) name13463 (
		_w15282_,
		_w19149_,
		_w23975_,
		_w23976_
	);
	LUT3 #(
		.INIT('h80)
	) name13464 (
		\wishbone_RxPointerMSB_reg[11]/NET0131 ,
		\wishbone_RxPointerMSB_reg[12]/NET0131 ,
		\wishbone_RxPointerMSB_reg[13]/NET0131 ,
		_w23977_
	);
	LUT4 #(
		.INIT('h8000)
	) name13465 (
		_w15283_,
		_w15284_,
		_w15285_,
		_w23977_,
		_w23978_
	);
	LUT4 #(
		.INIT('h0302)
	) name13466 (
		\wishbone_RxPointerMSB_reg[14]/NET0131 ,
		_w13807_,
		_w15288_,
		_w23978_,
		_w23979_
	);
	LUT3 #(
		.INIT('hf2)
	) name13467 (
		_w15282_,
		_w23950_,
		_w23979_,
		_w23980_
	);
	LUT3 #(
		.INIT('h12)
	) name13468 (
		\wishbone_RxPointerMSB_reg[4]/NET0131 ,
		_w13807_,
		_w15283_,
		_w23981_
	);
	LUT3 #(
		.INIT('hf2)
	) name13469 (
		_w15282_,
		_w20382_,
		_w23981_,
		_w23982_
	);
	LUT2 #(
		.INIT('h8)
	) name13470 (
		\wishbone_RxPointerMSB_reg[4]/NET0131 ,
		\wishbone_RxPointerMSB_reg[5]/NET0131 ,
		_w23983_
	);
	LUT4 #(
		.INIT('h060c)
	) name13471 (
		\wishbone_RxPointerMSB_reg[4]/NET0131 ,
		\wishbone_RxPointerMSB_reg[5]/NET0131 ,
		_w13807_,
		_w15283_,
		_w23984_
	);
	LUT3 #(
		.INIT('hf2)
	) name13472 (
		_w15282_,
		_w20754_,
		_w23984_,
		_w23985_
	);
	LUT4 #(
		.INIT('heddd)
	) name13473 (
		\wishbone_RxPointerMSB_reg[7]/NET0131 ,
		_w13807_,
		_w15283_,
		_w15284_,
		_w23986_
	);
	LUT3 #(
		.INIT('h2f)
	) name13474 (
		_w15282_,
		_w21117_,
		_w23986_,
		_w23987_
	);
	LUT3 #(
		.INIT('h15)
	) name13475 (
		\wishbone_RxPointerMSB_reg[6]/NET0131 ,
		_w15283_,
		_w23983_,
		_w23988_
	);
	LUT3 #(
		.INIT('h15)
	) name13476 (
		_w13807_,
		_w15283_,
		_w15284_,
		_w23989_
	);
	LUT2 #(
		.INIT('h4)
	) name13477 (
		_w23988_,
		_w23989_,
		_w23990_
	);
	LUT3 #(
		.INIT('hf2)
	) name13478 (
		_w15282_,
		_w23075_,
		_w23990_,
		_w23991_
	);
	LUT2 #(
		.INIT('h8)
	) name13479 (
		\wishbone_TxPointerMSB_reg[10]/NET0131 ,
		\wishbone_TxPointerMSB_reg[11]/NET0131 ,
		_w23992_
	);
	LUT4 #(
		.INIT('h8000)
	) name13480 (
		_w15305_,
		_w15306_,
		_w15307_,
		_w23992_,
		_w23993_
	);
	LUT4 #(
		.INIT('h0302)
	) name13481 (
		\wishbone_TxPointerMSB_reg[12]/NET0131 ,
		_w15303_,
		_w15310_,
		_w23993_,
		_w23994_
	);
	LUT3 #(
		.INIT('hf4)
	) name13482 (
		_w19149_,
		_w19180_,
		_w23994_,
		_w23995_
	);
	LUT4 #(
		.INIT('h060c)
	) name13483 (
		\wishbone_TxPointerMSB_reg[13]/NET0131 ,
		\wishbone_TxPointerMSB_reg[14]/NET0131 ,
		_w15303_,
		_w15310_,
		_w23996_
	);
	LUT3 #(
		.INIT('hf2)
	) name13484 (
		_w19180_,
		_w23950_,
		_w23996_,
		_w23997_
	);
	LUT3 #(
		.INIT('h12)
	) name13485 (
		\wishbone_TxPointerMSB_reg[4]/NET0131 ,
		_w15303_,
		_w15305_,
		_w23998_
	);
	LUT3 #(
		.INIT('hf2)
	) name13486 (
		_w19180_,
		_w20382_,
		_w23998_,
		_w23999_
	);
	LUT2 #(
		.INIT('h8)
	) name13487 (
		\wishbone_TxPointerMSB_reg[4]/NET0131 ,
		\wishbone_TxPointerMSB_reg[5]/NET0131 ,
		_w24000_
	);
	LUT4 #(
		.INIT('h060c)
	) name13488 (
		\wishbone_TxPointerMSB_reg[4]/NET0131 ,
		\wishbone_TxPointerMSB_reg[5]/NET0131 ,
		_w15303_,
		_w15305_,
		_w24001_
	);
	LUT3 #(
		.INIT('hf2)
	) name13489 (
		_w19180_,
		_w20754_,
		_w24001_,
		_w24002_
	);
	LUT3 #(
		.INIT('h15)
	) name13490 (
		\wishbone_TxPointerMSB_reg[6]/NET0131 ,
		_w15305_,
		_w24000_,
		_w24003_
	);
	LUT3 #(
		.INIT('h15)
	) name13491 (
		_w15303_,
		_w15305_,
		_w15306_,
		_w24004_
	);
	LUT2 #(
		.INIT('h4)
	) name13492 (
		_w24003_,
		_w24004_,
		_w24005_
	);
	LUT3 #(
		.INIT('hf2)
	) name13493 (
		_w19180_,
		_w23075_,
		_w24005_,
		_w24006_
	);
	LUT4 #(
		.INIT('heddd)
	) name13494 (
		\wishbone_TxPointerMSB_reg[7]/NET0131 ,
		_w15303_,
		_w15305_,
		_w15306_,
		_w24007_
	);
	LUT3 #(
		.INIT('h2f)
	) name13495 (
		_w19180_,
		_w21117_,
		_w24007_,
		_w24008_
	);
	LUT4 #(
		.INIT('h70f0)
	) name13496 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxPointerMSB_reg[11]/NET0131 ,
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w24009_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13497 (
		_w15283_,
		_w15284_,
		_w15285_,
		_w24009_,
		_w24010_
	);
	LUT4 #(
		.INIT('h070f)
	) name13498 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxPointerMSB_reg[11]/NET0131 ,
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w24011_
	);
	LUT4 #(
		.INIT('h8000)
	) name13499 (
		_w15283_,
		_w15284_,
		_w15285_,
		_w24011_,
		_w24012_
	);
	LUT2 #(
		.INIT('h1)
	) name13500 (
		_w24010_,
		_w24012_,
		_w24013_
	);
	LUT3 #(
		.INIT('h2f)
	) name13501 (
		_w15282_,
		_w22213_,
		_w24013_,
		_w24014_
	);
	LUT4 #(
		.INIT('h0032)
	) name13502 (
		\wishbone_RxPointerMSB_reg[13]/NET0131 ,
		_w13807_,
		_w23974_,
		_w23978_,
		_w24015_
	);
	LUT3 #(
		.INIT('hf2)
	) name13503 (
		_w15282_,
		_w23589_,
		_w24015_,
		_w24016_
	);
	LUT3 #(
		.INIT('hed)
	) name13504 (
		\wishbone_RxPointerMSB_reg[15]/NET0131 ,
		_w13807_,
		_w15288_,
		_w24017_
	);
	LUT3 #(
		.INIT('h4f)
	) name13505 (
		_w13800_,
		_w15282_,
		_w24017_,
		_w24018_
	);
	LUT2 #(
		.INIT('h8)
	) name13506 (
		\wishbone_RxPointerMSB_reg[15]/NET0131 ,
		\wishbone_RxPointerMSB_reg[16]/NET0131 ,
		_w24019_
	);
	LUT4 #(
		.INIT('h060c)
	) name13507 (
		\wishbone_RxPointerMSB_reg[15]/NET0131 ,
		\wishbone_RxPointerMSB_reg[16]/NET0131 ,
		_w13807_,
		_w15288_,
		_w24020_
	);
	LUT3 #(
		.INIT('hf2)
	) name13508 (
		_w15282_,
		_w16122_,
		_w24020_,
		_w24021_
	);
	LUT3 #(
		.INIT('h15)
	) name13509 (
		\wishbone_RxPointerMSB_reg[17]/NET0131 ,
		_w15288_,
		_w24019_,
		_w24022_
	);
	LUT3 #(
		.INIT('h15)
	) name13510 (
		_w13807_,
		_w15288_,
		_w23117_,
		_w24023_
	);
	LUT2 #(
		.INIT('h4)
	) name13511 (
		_w24022_,
		_w24023_,
		_w24024_
	);
	LUT3 #(
		.INIT('hf2)
	) name13512 (
		_w15282_,
		_w16814_,
		_w24024_,
		_w24025_
	);
	LUT4 #(
		.INIT('heddd)
	) name13513 (
		\wishbone_RxPointerMSB_reg[18]/NET0131 ,
		_w13807_,
		_w15288_,
		_w23117_,
		_w24026_
	);
	LUT3 #(
		.INIT('h2f)
	) name13514 (
		_w15282_,
		_w15775_,
		_w24026_,
		_w24027_
	);
	LUT3 #(
		.INIT('h12)
	) name13515 (
		\wishbone_RxPointerMSB_reg[2]/NET0131 ,
		_w13807_,
		_w13809_,
		_w24028_
	);
	LUT3 #(
		.INIT('hf2)
	) name13516 (
		_w15282_,
		_w22594_,
		_w24028_,
		_w24029_
	);
	LUT4 #(
		.INIT('h007f)
	) name13517 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_RxPointerMSB_reg[2]/NET0131 ,
		\wishbone_RxPointerMSB_reg[3]/NET0131 ,
		_w24030_
	);
	LUT3 #(
		.INIT('h01)
	) name13518 (
		_w13807_,
		_w15283_,
		_w24030_,
		_w24031_
	);
	LUT3 #(
		.INIT('hf2)
	) name13519 (
		_w15282_,
		_w20008_,
		_w24031_,
		_w24032_
	);
	LUT4 #(
		.INIT('h1333)
	) name13520 (
		\wishbone_RxPointerMSB_reg[7]/NET0131 ,
		\wishbone_RxPointerMSB_reg[8]/NET0131 ,
		_w15283_,
		_w15284_,
		_w24033_
	);
	LUT4 #(
		.INIT('h1555)
	) name13521 (
		_w13807_,
		_w15283_,
		_w15284_,
		_w23167_,
		_w24034_
	);
	LUT2 #(
		.INIT('h4)
	) name13522 (
		_w24033_,
		_w24034_,
		_w24035_
	);
	LUT3 #(
		.INIT('hf2)
	) name13523 (
		_w15282_,
		_w21480_,
		_w24035_,
		_w24036_
	);
	LUT4 #(
		.INIT('h70f0)
	) name13524 (
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		\wishbone_TxPointerMSB_reg[10]/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w24037_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13525 (
		_w15305_,
		_w15306_,
		_w15307_,
		_w24037_,
		_w24038_
	);
	LUT4 #(
		.INIT('h070f)
	) name13526 (
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		\wishbone_TxPointerMSB_reg[10]/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w24039_
	);
	LUT4 #(
		.INIT('h8000)
	) name13527 (
		_w15305_,
		_w15306_,
		_w15307_,
		_w24039_,
		_w24040_
	);
	LUT2 #(
		.INIT('h1)
	) name13528 (
		_w24038_,
		_w24040_,
		_w24041_
	);
	LUT3 #(
		.INIT('h80)
	) name13529 (
		\wishbone_bd_ram_mem1_reg[20][10]/P0001 ,
		_w11929_,
		_w11935_,
		_w24042_
	);
	LUT3 #(
		.INIT('h80)
	) name13530 (
		\wishbone_bd_ram_mem1_reg[88][10]/P0001 ,
		_w11972_,
		_w11990_,
		_w24043_
	);
	LUT3 #(
		.INIT('h80)
	) name13531 (
		\wishbone_bd_ram_mem1_reg[33][10]/P0001 ,
		_w11957_,
		_w11977_,
		_w24044_
	);
	LUT3 #(
		.INIT('h80)
	) name13532 (
		\wishbone_bd_ram_mem1_reg[222][10]/P0001 ,
		_w11948_,
		_w11984_,
		_w24045_
	);
	LUT4 #(
		.INIT('h0001)
	) name13533 (
		_w24042_,
		_w24043_,
		_w24044_,
		_w24045_,
		_w24046_
	);
	LUT3 #(
		.INIT('h80)
	) name13534 (
		\wishbone_bd_ram_mem1_reg[134][10]/P0001 ,
		_w11955_,
		_w11986_,
		_w24047_
	);
	LUT3 #(
		.INIT('h80)
	) name13535 (
		\wishbone_bd_ram_mem1_reg[199][10]/P0001 ,
		_w11945_,
		_w11975_,
		_w24048_
	);
	LUT3 #(
		.INIT('h80)
	) name13536 (
		\wishbone_bd_ram_mem1_reg[112][10]/P0001 ,
		_w11941_,
		_w12012_,
		_w24049_
	);
	LUT3 #(
		.INIT('h80)
	) name13537 (
		\wishbone_bd_ram_mem1_reg[78][10]/P0001 ,
		_w11948_,
		_w11949_,
		_w24050_
	);
	LUT4 #(
		.INIT('h0001)
	) name13538 (
		_w24047_,
		_w24048_,
		_w24049_,
		_w24050_,
		_w24051_
	);
	LUT3 #(
		.INIT('h80)
	) name13539 (
		\wishbone_bd_ram_mem1_reg[208][10]/P0001 ,
		_w11941_,
		_w11984_,
		_w24052_
	);
	LUT3 #(
		.INIT('h80)
	) name13540 (
		\wishbone_bd_ram_mem1_reg[107][10]/P0001 ,
		_w11936_,
		_w11965_,
		_w24053_
	);
	LUT3 #(
		.INIT('h80)
	) name13541 (
		\wishbone_bd_ram_mem1_reg[118][10]/P0001 ,
		_w11986_,
		_w12012_,
		_w24054_
	);
	LUT3 #(
		.INIT('h80)
	) name13542 (
		\wishbone_bd_ram_mem1_reg[155][10]/P0001 ,
		_w11936_,
		_w11959_,
		_w24055_
	);
	LUT4 #(
		.INIT('h0001)
	) name13543 (
		_w24052_,
		_w24053_,
		_w24054_,
		_w24055_,
		_w24056_
	);
	LUT3 #(
		.INIT('h80)
	) name13544 (
		\wishbone_bd_ram_mem1_reg[193][10]/P0001 ,
		_w11945_,
		_w11977_,
		_w24057_
	);
	LUT3 #(
		.INIT('h80)
	) name13545 (
		\wishbone_bd_ram_mem1_reg[116][10]/P0001 ,
		_w11929_,
		_w12012_,
		_w24058_
	);
	LUT3 #(
		.INIT('h80)
	) name13546 (
		\wishbone_bd_ram_mem1_reg[251][10]/P0001 ,
		_w11936_,
		_w11952_,
		_w24059_
	);
	LUT3 #(
		.INIT('h80)
	) name13547 (
		\wishbone_bd_ram_mem1_reg[113][10]/P0001 ,
		_w11977_,
		_w12012_,
		_w24060_
	);
	LUT4 #(
		.INIT('h0001)
	) name13548 (
		_w24057_,
		_w24058_,
		_w24059_,
		_w24060_,
		_w24061_
	);
	LUT4 #(
		.INIT('h8000)
	) name13549 (
		_w24046_,
		_w24051_,
		_w24056_,
		_w24061_,
		_w24062_
	);
	LUT3 #(
		.INIT('h80)
	) name13550 (
		\wishbone_bd_ram_mem1_reg[200][10]/P0001 ,
		_w11945_,
		_w11990_,
		_w24063_
	);
	LUT3 #(
		.INIT('h80)
	) name13551 (
		\wishbone_bd_ram_mem1_reg[148][10]/P0001 ,
		_w11929_,
		_w11959_,
		_w24064_
	);
	LUT3 #(
		.INIT('h80)
	) name13552 (
		\wishbone_bd_ram_mem1_reg[230][10]/P0001 ,
		_w11982_,
		_w11986_,
		_w24065_
	);
	LUT3 #(
		.INIT('h80)
	) name13553 (
		\wishbone_bd_ram_mem1_reg[14][10]/P0001 ,
		_w11932_,
		_w11948_,
		_w24066_
	);
	LUT4 #(
		.INIT('h0001)
	) name13554 (
		_w24063_,
		_w24064_,
		_w24065_,
		_w24066_,
		_w24067_
	);
	LUT3 #(
		.INIT('h80)
	) name13555 (
		\wishbone_bd_ram_mem1_reg[38][10]/P0001 ,
		_w11957_,
		_w11986_,
		_w24068_
	);
	LUT3 #(
		.INIT('h80)
	) name13556 (
		\wishbone_bd_ram_mem1_reg[64][10]/P0001 ,
		_w11941_,
		_w11949_,
		_w24069_
	);
	LUT3 #(
		.INIT('h80)
	) name13557 (
		\wishbone_bd_ram_mem1_reg[132][10]/P0001 ,
		_w11929_,
		_w11955_,
		_w24070_
	);
	LUT3 #(
		.INIT('h80)
	) name13558 (
		\wishbone_bd_ram_mem1_reg[235][10]/P0001 ,
		_w11936_,
		_w11982_,
		_w24071_
	);
	LUT4 #(
		.INIT('h0001)
	) name13559 (
		_w24068_,
		_w24069_,
		_w24070_,
		_w24071_,
		_w24072_
	);
	LUT3 #(
		.INIT('h80)
	) name13560 (
		\wishbone_bd_ram_mem1_reg[255][10]/P0001 ,
		_w11952_,
		_w11973_,
		_w24073_
	);
	LUT3 #(
		.INIT('h80)
	) name13561 (
		\wishbone_bd_ram_mem1_reg[71][10]/P0001 ,
		_w11949_,
		_w11975_,
		_w24074_
	);
	LUT3 #(
		.INIT('h80)
	) name13562 (
		\wishbone_bd_ram_mem1_reg[127][10]/P0001 ,
		_w11973_,
		_w12012_,
		_w24075_
	);
	LUT3 #(
		.INIT('h80)
	) name13563 (
		\wishbone_bd_ram_mem1_reg[21][10]/P0001 ,
		_w11933_,
		_w11935_,
		_w24076_
	);
	LUT4 #(
		.INIT('h0001)
	) name13564 (
		_w24073_,
		_w24074_,
		_w24075_,
		_w24076_,
		_w24077_
	);
	LUT3 #(
		.INIT('h80)
	) name13565 (
		\wishbone_bd_ram_mem1_reg[17][10]/P0001 ,
		_w11935_,
		_w11977_,
		_w24078_
	);
	LUT3 #(
		.INIT('h80)
	) name13566 (
		\wishbone_bd_ram_mem1_reg[0][10]/P0001 ,
		_w11932_,
		_w11941_,
		_w24079_
	);
	LUT3 #(
		.INIT('h80)
	) name13567 (
		\wishbone_bd_ram_mem1_reg[27][10]/P0001 ,
		_w11935_,
		_w11936_,
		_w24080_
	);
	LUT3 #(
		.INIT('h80)
	) name13568 (
		\wishbone_bd_ram_mem1_reg[158][10]/P0001 ,
		_w11948_,
		_w11959_,
		_w24081_
	);
	LUT4 #(
		.INIT('h0001)
	) name13569 (
		_w24078_,
		_w24079_,
		_w24080_,
		_w24081_,
		_w24082_
	);
	LUT4 #(
		.INIT('h8000)
	) name13570 (
		_w24067_,
		_w24072_,
		_w24077_,
		_w24082_,
		_w24083_
	);
	LUT3 #(
		.INIT('h80)
	) name13571 (
		\wishbone_bd_ram_mem1_reg[247][10]/P0001 ,
		_w11952_,
		_w11975_,
		_w24084_
	);
	LUT3 #(
		.INIT('h80)
	) name13572 (
		\wishbone_bd_ram_mem1_reg[180][10]/P0001 ,
		_w11929_,
		_w11942_,
		_w24085_
	);
	LUT3 #(
		.INIT('h80)
	) name13573 (
		\wishbone_bd_ram_mem1_reg[225][10]/P0001 ,
		_w11977_,
		_w11982_,
		_w24086_
	);
	LUT3 #(
		.INIT('h80)
	) name13574 (
		\wishbone_bd_ram_mem1_reg[145][10]/P0001 ,
		_w11959_,
		_w11977_,
		_w24087_
	);
	LUT4 #(
		.INIT('h0001)
	) name13575 (
		_w24084_,
		_w24085_,
		_w24086_,
		_w24087_,
		_w24088_
	);
	LUT3 #(
		.INIT('h80)
	) name13576 (
		\wishbone_bd_ram_mem1_reg[49][10]/P0001 ,
		_w11977_,
		_w11979_,
		_w24089_
	);
	LUT3 #(
		.INIT('h80)
	) name13577 (
		\wishbone_bd_ram_mem1_reg[128][10]/P0001 ,
		_w11941_,
		_w11955_,
		_w24090_
	);
	LUT3 #(
		.INIT('h80)
	) name13578 (
		\wishbone_bd_ram_mem1_reg[245][10]/P0001 ,
		_w11933_,
		_w11952_,
		_w24091_
	);
	LUT3 #(
		.INIT('h80)
	) name13579 (
		\wishbone_bd_ram_mem1_reg[120][10]/P0001 ,
		_w11990_,
		_w12012_,
		_w24092_
	);
	LUT4 #(
		.INIT('h0001)
	) name13580 (
		_w24089_,
		_w24090_,
		_w24091_,
		_w24092_,
		_w24093_
	);
	LUT3 #(
		.INIT('h80)
	) name13581 (
		\wishbone_bd_ram_mem1_reg[106][10]/P0001 ,
		_w11944_,
		_w11965_,
		_w24094_
	);
	LUT3 #(
		.INIT('h80)
	) name13582 (
		\wishbone_bd_ram_mem1_reg[212][10]/P0001 ,
		_w11929_,
		_w11984_,
		_w24095_
	);
	LUT3 #(
		.INIT('h80)
	) name13583 (
		\wishbone_bd_ram_mem1_reg[246][10]/P0001 ,
		_w11952_,
		_w11986_,
		_w24096_
	);
	LUT3 #(
		.INIT('h80)
	) name13584 (
		\wishbone_bd_ram_mem1_reg[181][10]/P0001 ,
		_w11933_,
		_w11942_,
		_w24097_
	);
	LUT4 #(
		.INIT('h0001)
	) name13585 (
		_w24094_,
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_
	);
	LUT3 #(
		.INIT('h80)
	) name13586 (
		\wishbone_bd_ram_mem1_reg[196][10]/P0001 ,
		_w11929_,
		_w11945_,
		_w24099_
	);
	LUT3 #(
		.INIT('h80)
	) name13587 (
		\wishbone_bd_ram_mem1_reg[81][10]/P0001 ,
		_w11972_,
		_w11977_,
		_w24100_
	);
	LUT3 #(
		.INIT('h80)
	) name13588 (
		\wishbone_bd_ram_mem1_reg[183][10]/P0001 ,
		_w11942_,
		_w11975_,
		_w24101_
	);
	LUT3 #(
		.INIT('h80)
	) name13589 (
		\wishbone_bd_ram_mem1_reg[250][10]/P0001 ,
		_w11944_,
		_w11952_,
		_w24102_
	);
	LUT4 #(
		.INIT('h0001)
	) name13590 (
		_w24099_,
		_w24100_,
		_w24101_,
		_w24102_,
		_w24103_
	);
	LUT4 #(
		.INIT('h8000)
	) name13591 (
		_w24088_,
		_w24093_,
		_w24098_,
		_w24103_,
		_w24104_
	);
	LUT3 #(
		.INIT('h80)
	) name13592 (
		\wishbone_bd_ram_mem1_reg[241][10]/P0001 ,
		_w11952_,
		_w11977_,
		_w24105_
	);
	LUT3 #(
		.INIT('h80)
	) name13593 (
		\wishbone_bd_ram_mem1_reg[146][10]/P0001 ,
		_w11959_,
		_w11963_,
		_w24106_
	);
	LUT3 #(
		.INIT('h80)
	) name13594 (
		\wishbone_bd_ram_mem1_reg[18][10]/P0001 ,
		_w11935_,
		_w11963_,
		_w24107_
	);
	LUT3 #(
		.INIT('h80)
	) name13595 (
		\wishbone_bd_ram_mem1_reg[58][10]/P0001 ,
		_w11944_,
		_w11979_,
		_w24108_
	);
	LUT4 #(
		.INIT('h0001)
	) name13596 (
		_w24105_,
		_w24106_,
		_w24107_,
		_w24108_,
		_w24109_
	);
	LUT3 #(
		.INIT('h80)
	) name13597 (
		\wishbone_bd_ram_mem1_reg[83][10]/P0001 ,
		_w11938_,
		_w11972_,
		_w24110_
	);
	LUT3 #(
		.INIT('h80)
	) name13598 (
		\wishbone_bd_ram_mem1_reg[79][10]/P0001 ,
		_w11949_,
		_w11973_,
		_w24111_
	);
	LUT3 #(
		.INIT('h80)
	) name13599 (
		\wishbone_bd_ram_mem1_reg[204][10]/P0001 ,
		_w11945_,
		_w11954_,
		_w24112_
	);
	LUT3 #(
		.INIT('h80)
	) name13600 (
		\wishbone_bd_ram_mem1_reg[243][10]/P0001 ,
		_w11938_,
		_w11952_,
		_w24113_
	);
	LUT4 #(
		.INIT('h0001)
	) name13601 (
		_w24110_,
		_w24111_,
		_w24112_,
		_w24113_,
		_w24114_
	);
	LUT3 #(
		.INIT('h80)
	) name13602 (
		\wishbone_bd_ram_mem1_reg[24][10]/P0001 ,
		_w11935_,
		_w11990_,
		_w24115_
	);
	LUT3 #(
		.INIT('h80)
	) name13603 (
		\wishbone_bd_ram_mem1_reg[149][10]/P0001 ,
		_w11933_,
		_w11959_,
		_w24116_
	);
	LUT3 #(
		.INIT('h80)
	) name13604 (
		\wishbone_bd_ram_mem1_reg[32][10]/P0001 ,
		_w11941_,
		_w11957_,
		_w24117_
	);
	LUT3 #(
		.INIT('h80)
	) name13605 (
		\wishbone_bd_ram_mem1_reg[42][10]/P0001 ,
		_w11944_,
		_w11957_,
		_w24118_
	);
	LUT4 #(
		.INIT('h0001)
	) name13606 (
		_w24115_,
		_w24116_,
		_w24117_,
		_w24118_,
		_w24119_
	);
	LUT3 #(
		.INIT('h80)
	) name13607 (
		\wishbone_bd_ram_mem1_reg[133][10]/P0001 ,
		_w11933_,
		_w11955_,
		_w24120_
	);
	LUT3 #(
		.INIT('h80)
	) name13608 (
		\wishbone_bd_ram_mem1_reg[52][10]/P0001 ,
		_w11929_,
		_w11979_,
		_w24121_
	);
	LUT3 #(
		.INIT('h80)
	) name13609 (
		\wishbone_bd_ram_mem1_reg[136][10]/P0001 ,
		_w11955_,
		_w11990_,
		_w24122_
	);
	LUT3 #(
		.INIT('h80)
	) name13610 (
		\wishbone_bd_ram_mem1_reg[86][10]/P0001 ,
		_w11972_,
		_w11986_,
		_w24123_
	);
	LUT4 #(
		.INIT('h0001)
	) name13611 (
		_w24120_,
		_w24121_,
		_w24122_,
		_w24123_,
		_w24124_
	);
	LUT4 #(
		.INIT('h8000)
	) name13612 (
		_w24109_,
		_w24114_,
		_w24119_,
		_w24124_,
		_w24125_
	);
	LUT4 #(
		.INIT('h8000)
	) name13613 (
		_w24062_,
		_w24083_,
		_w24104_,
		_w24125_,
		_w24126_
	);
	LUT3 #(
		.INIT('h80)
	) name13614 (
		\wishbone_bd_ram_mem1_reg[103][10]/P0001 ,
		_w11965_,
		_w11975_,
		_w24127_
	);
	LUT3 #(
		.INIT('h80)
	) name13615 (
		\wishbone_bd_ram_mem1_reg[56][10]/P0001 ,
		_w11979_,
		_w11990_,
		_w24128_
	);
	LUT3 #(
		.INIT('h80)
	) name13616 (
		\wishbone_bd_ram_mem1_reg[220][10]/P0001 ,
		_w11954_,
		_w11984_,
		_w24129_
	);
	LUT3 #(
		.INIT('h80)
	) name13617 (
		\wishbone_bd_ram_mem1_reg[131][10]/P0001 ,
		_w11938_,
		_w11955_,
		_w24130_
	);
	LUT4 #(
		.INIT('h0001)
	) name13618 (
		_w24127_,
		_w24128_,
		_w24129_,
		_w24130_,
		_w24131_
	);
	LUT3 #(
		.INIT('h80)
	) name13619 (
		\wishbone_bd_ram_mem1_reg[141][10]/P0001 ,
		_w11955_,
		_w11966_,
		_w24132_
	);
	LUT3 #(
		.INIT('h80)
	) name13620 (
		\wishbone_bd_ram_mem1_reg[137][10]/P0001 ,
		_w11955_,
		_w11968_,
		_w24133_
	);
	LUT3 #(
		.INIT('h80)
	) name13621 (
		\wishbone_bd_ram_mem1_reg[191][10]/P0001 ,
		_w11942_,
		_w11973_,
		_w24134_
	);
	LUT3 #(
		.INIT('h80)
	) name13622 (
		\wishbone_bd_ram_mem1_reg[177][10]/P0001 ,
		_w11942_,
		_w11977_,
		_w24135_
	);
	LUT4 #(
		.INIT('h0001)
	) name13623 (
		_w24132_,
		_w24133_,
		_w24134_,
		_w24135_,
		_w24136_
	);
	LUT3 #(
		.INIT('h80)
	) name13624 (
		\wishbone_bd_ram_mem1_reg[70][10]/P0001 ,
		_w11949_,
		_w11986_,
		_w24137_
	);
	LUT3 #(
		.INIT('h80)
	) name13625 (
		\wishbone_bd_ram_mem1_reg[10][10]/P0001 ,
		_w11932_,
		_w11944_,
		_w24138_
	);
	LUT3 #(
		.INIT('h80)
	) name13626 (
		\wishbone_bd_ram_mem1_reg[219][10]/P0001 ,
		_w11936_,
		_w11984_,
		_w24139_
	);
	LUT3 #(
		.INIT('h80)
	) name13627 (
		\wishbone_bd_ram_mem1_reg[236][10]/P0001 ,
		_w11954_,
		_w11982_,
		_w24140_
	);
	LUT4 #(
		.INIT('h0001)
	) name13628 (
		_w24137_,
		_w24138_,
		_w24139_,
		_w24140_,
		_w24141_
	);
	LUT3 #(
		.INIT('h80)
	) name13629 (
		\wishbone_bd_ram_mem1_reg[228][10]/P0001 ,
		_w11929_,
		_w11982_,
		_w24142_
	);
	LUT3 #(
		.INIT('h80)
	) name13630 (
		\wishbone_bd_ram_mem1_reg[65][10]/P0001 ,
		_w11949_,
		_w11977_,
		_w24143_
	);
	LUT3 #(
		.INIT('h80)
	) name13631 (
		\wishbone_bd_ram_mem1_reg[189][10]/P0001 ,
		_w11942_,
		_w11966_,
		_w24144_
	);
	LUT3 #(
		.INIT('h80)
	) name13632 (
		\wishbone_bd_ram_mem1_reg[82][10]/P0001 ,
		_w11963_,
		_w11972_,
		_w24145_
	);
	LUT4 #(
		.INIT('h0001)
	) name13633 (
		_w24142_,
		_w24143_,
		_w24144_,
		_w24145_,
		_w24146_
	);
	LUT4 #(
		.INIT('h8000)
	) name13634 (
		_w24131_,
		_w24136_,
		_w24141_,
		_w24146_,
		_w24147_
	);
	LUT3 #(
		.INIT('h80)
	) name13635 (
		\wishbone_bd_ram_mem1_reg[210][10]/P0001 ,
		_w11963_,
		_w11984_,
		_w24148_
	);
	LUT3 #(
		.INIT('h80)
	) name13636 (
		\wishbone_bd_ram_mem1_reg[159][10]/P0001 ,
		_w11959_,
		_w11973_,
		_w24149_
	);
	LUT3 #(
		.INIT('h80)
	) name13637 (
		\wishbone_bd_ram_mem1_reg[43][10]/P0001 ,
		_w11936_,
		_w11957_,
		_w24150_
	);
	LUT3 #(
		.INIT('h80)
	) name13638 (
		\wishbone_bd_ram_mem1_reg[253][10]/P0001 ,
		_w11952_,
		_w11966_,
		_w24151_
	);
	LUT4 #(
		.INIT('h0001)
	) name13639 (
		_w24148_,
		_w24149_,
		_w24150_,
		_w24151_,
		_w24152_
	);
	LUT3 #(
		.INIT('h80)
	) name13640 (
		\wishbone_bd_ram_mem1_reg[124][10]/P0001 ,
		_w11954_,
		_w12012_,
		_w24153_
	);
	LUT3 #(
		.INIT('h80)
	) name13641 (
		\wishbone_bd_ram_mem1_reg[3][10]/P0001 ,
		_w11932_,
		_w11938_,
		_w24154_
	);
	LUT3 #(
		.INIT('h80)
	) name13642 (
		\wishbone_bd_ram_mem1_reg[164][10]/P0001 ,
		_w11929_,
		_w11930_,
		_w24155_
	);
	LUT3 #(
		.INIT('h80)
	) name13643 (
		\wishbone_bd_ram_mem1_reg[29][10]/P0001 ,
		_w11935_,
		_w11966_,
		_w24156_
	);
	LUT4 #(
		.INIT('h0001)
	) name13644 (
		_w24153_,
		_w24154_,
		_w24155_,
		_w24156_,
		_w24157_
	);
	LUT3 #(
		.INIT('h80)
	) name13645 (
		\wishbone_bd_ram_mem1_reg[77][10]/P0001 ,
		_w11949_,
		_w11966_,
		_w24158_
	);
	LUT3 #(
		.INIT('h80)
	) name13646 (
		\wishbone_bd_ram_mem1_reg[249][10]/P0001 ,
		_w11952_,
		_w11968_,
		_w24159_
	);
	LUT3 #(
		.INIT('h80)
	) name13647 (
		\wishbone_bd_ram_mem1_reg[119][10]/P0001 ,
		_w11975_,
		_w12012_,
		_w24160_
	);
	LUT3 #(
		.INIT('h80)
	) name13648 (
		\wishbone_bd_ram_mem1_reg[92][10]/P0001 ,
		_w11954_,
		_w11972_,
		_w24161_
	);
	LUT4 #(
		.INIT('h0001)
	) name13649 (
		_w24158_,
		_w24159_,
		_w24160_,
		_w24161_,
		_w24162_
	);
	LUT3 #(
		.INIT('h80)
	) name13650 (
		\wishbone_bd_ram_mem1_reg[60][10]/P0001 ,
		_w11954_,
		_w11979_,
		_w24163_
	);
	LUT3 #(
		.INIT('h80)
	) name13651 (
		\wishbone_bd_ram_mem1_reg[30][10]/P0001 ,
		_w11935_,
		_w11948_,
		_w24164_
	);
	LUT3 #(
		.INIT('h80)
	) name13652 (
		\wishbone_bd_ram_mem1_reg[242][10]/P0001 ,
		_w11952_,
		_w11963_,
		_w24165_
	);
	LUT3 #(
		.INIT('h80)
	) name13653 (
		\wishbone_bd_ram_mem1_reg[48][10]/P0001 ,
		_w11941_,
		_w11979_,
		_w24166_
	);
	LUT4 #(
		.INIT('h0001)
	) name13654 (
		_w24163_,
		_w24164_,
		_w24165_,
		_w24166_,
		_w24167_
	);
	LUT4 #(
		.INIT('h8000)
	) name13655 (
		_w24152_,
		_w24157_,
		_w24162_,
		_w24167_,
		_w24168_
	);
	LUT3 #(
		.INIT('h80)
	) name13656 (
		\wishbone_bd_ram_mem1_reg[28][10]/P0001 ,
		_w11935_,
		_w11954_,
		_w24169_
	);
	LUT3 #(
		.INIT('h80)
	) name13657 (
		\wishbone_bd_ram_mem1_reg[100][10]/P0001 ,
		_w11929_,
		_w11965_,
		_w24170_
	);
	LUT3 #(
		.INIT('h80)
	) name13658 (
		\wishbone_bd_ram_mem1_reg[102][10]/P0001 ,
		_w11965_,
		_w11986_,
		_w24171_
	);
	LUT3 #(
		.INIT('h80)
	) name13659 (
		\wishbone_bd_ram_mem1_reg[161][10]/P0001 ,
		_w11930_,
		_w11977_,
		_w24172_
	);
	LUT4 #(
		.INIT('h0001)
	) name13660 (
		_w24169_,
		_w24170_,
		_w24171_,
		_w24172_,
		_w24173_
	);
	LUT3 #(
		.INIT('h80)
	) name13661 (
		\wishbone_bd_ram_mem1_reg[90][10]/P0001 ,
		_w11944_,
		_w11972_,
		_w24174_
	);
	LUT3 #(
		.INIT('h80)
	) name13662 (
		\wishbone_bd_ram_mem1_reg[252][10]/P0001 ,
		_w11952_,
		_w11954_,
		_w24175_
	);
	LUT3 #(
		.INIT('h80)
	) name13663 (
		\wishbone_bd_ram_mem1_reg[39][10]/P0001 ,
		_w11957_,
		_w11975_,
		_w24176_
	);
	LUT3 #(
		.INIT('h80)
	) name13664 (
		\wishbone_bd_ram_mem1_reg[175][10]/P0001 ,
		_w11930_,
		_w11973_,
		_w24177_
	);
	LUT4 #(
		.INIT('h0001)
	) name13665 (
		_w24174_,
		_w24175_,
		_w24176_,
		_w24177_,
		_w24178_
	);
	LUT3 #(
		.INIT('h80)
	) name13666 (
		\wishbone_bd_ram_mem1_reg[184][10]/P0001 ,
		_w11942_,
		_w11990_,
		_w24179_
	);
	LUT3 #(
		.INIT('h80)
	) name13667 (
		\wishbone_bd_ram_mem1_reg[139][10]/P0001 ,
		_w11936_,
		_w11955_,
		_w24180_
	);
	LUT3 #(
		.INIT('h80)
	) name13668 (
		\wishbone_bd_ram_mem1_reg[93][10]/P0001 ,
		_w11966_,
		_w11972_,
		_w24181_
	);
	LUT3 #(
		.INIT('h80)
	) name13669 (
		\wishbone_bd_ram_mem1_reg[76][10]/P0001 ,
		_w11949_,
		_w11954_,
		_w24182_
	);
	LUT4 #(
		.INIT('h0001)
	) name13670 (
		_w24179_,
		_w24180_,
		_w24181_,
		_w24182_,
		_w24183_
	);
	LUT3 #(
		.INIT('h80)
	) name13671 (
		\wishbone_bd_ram_mem1_reg[151][10]/P0001 ,
		_w11959_,
		_w11975_,
		_w24184_
	);
	LUT3 #(
		.INIT('h80)
	) name13672 (
		\wishbone_bd_ram_mem1_reg[240][10]/P0001 ,
		_w11941_,
		_w11952_,
		_w24185_
	);
	LUT3 #(
		.INIT('h80)
	) name13673 (
		\wishbone_bd_ram_mem1_reg[122][10]/P0001 ,
		_w11944_,
		_w12012_,
		_w24186_
	);
	LUT3 #(
		.INIT('h80)
	) name13674 (
		\wishbone_bd_ram_mem1_reg[215][10]/P0001 ,
		_w11975_,
		_w11984_,
		_w24187_
	);
	LUT4 #(
		.INIT('h0001)
	) name13675 (
		_w24184_,
		_w24185_,
		_w24186_,
		_w24187_,
		_w24188_
	);
	LUT4 #(
		.INIT('h8000)
	) name13676 (
		_w24173_,
		_w24178_,
		_w24183_,
		_w24188_,
		_w24189_
	);
	LUT3 #(
		.INIT('h80)
	) name13677 (
		\wishbone_bd_ram_mem1_reg[22][10]/P0001 ,
		_w11935_,
		_w11986_,
		_w24190_
	);
	LUT3 #(
		.INIT('h80)
	) name13678 (
		\wishbone_bd_ram_mem1_reg[140][10]/P0001 ,
		_w11954_,
		_w11955_,
		_w24191_
	);
	LUT3 #(
		.INIT('h80)
	) name13679 (
		\wishbone_bd_ram_mem1_reg[111][10]/P0001 ,
		_w11965_,
		_w11973_,
		_w24192_
	);
	LUT3 #(
		.INIT('h80)
	) name13680 (
		\wishbone_bd_ram_mem1_reg[165][10]/P0001 ,
		_w11930_,
		_w11933_,
		_w24193_
	);
	LUT4 #(
		.INIT('h0001)
	) name13681 (
		_w24190_,
		_w24191_,
		_w24192_,
		_w24193_,
		_w24194_
	);
	LUT3 #(
		.INIT('h80)
	) name13682 (
		\wishbone_bd_ram_mem1_reg[206][10]/P0001 ,
		_w11945_,
		_w11948_,
		_w24195_
	);
	LUT3 #(
		.INIT('h80)
	) name13683 (
		\wishbone_bd_ram_mem1_reg[163][10]/P0001 ,
		_w11930_,
		_w11938_,
		_w24196_
	);
	LUT3 #(
		.INIT('h80)
	) name13684 (
		\wishbone_bd_ram_mem1_reg[187][10]/P0001 ,
		_w11936_,
		_w11942_,
		_w24197_
	);
	LUT3 #(
		.INIT('h80)
	) name13685 (
		\wishbone_bd_ram_mem1_reg[162][10]/P0001 ,
		_w11930_,
		_w11963_,
		_w24198_
	);
	LUT4 #(
		.INIT('h0001)
	) name13686 (
		_w24195_,
		_w24196_,
		_w24197_,
		_w24198_,
		_w24199_
	);
	LUT3 #(
		.INIT('h80)
	) name13687 (
		\wishbone_bd_ram_mem1_reg[12][10]/P0001 ,
		_w11932_,
		_w11954_,
		_w24200_
	);
	LUT3 #(
		.INIT('h80)
	) name13688 (
		\wishbone_bd_ram_mem1_reg[99][10]/P0001 ,
		_w11938_,
		_w11965_,
		_w24201_
	);
	LUT3 #(
		.INIT('h80)
	) name13689 (
		\wishbone_bd_ram_mem1_reg[41][10]/P0001 ,
		_w11957_,
		_w11968_,
		_w24202_
	);
	LUT3 #(
		.INIT('h80)
	) name13690 (
		\wishbone_bd_ram_mem1_reg[54][10]/P0001 ,
		_w11979_,
		_w11986_,
		_w24203_
	);
	LUT4 #(
		.INIT('h0001)
	) name13691 (
		_w24200_,
		_w24201_,
		_w24202_,
		_w24203_,
		_w24204_
	);
	LUT3 #(
		.INIT('h80)
	) name13692 (
		\wishbone_bd_ram_mem1_reg[44][10]/P0001 ,
		_w11954_,
		_w11957_,
		_w24205_
	);
	LUT3 #(
		.INIT('h80)
	) name13693 (
		\wishbone_bd_ram_mem1_reg[188][10]/P0001 ,
		_w11942_,
		_w11954_,
		_w24206_
	);
	LUT3 #(
		.INIT('h80)
	) name13694 (
		\wishbone_bd_ram_mem1_reg[31][10]/P0001 ,
		_w11935_,
		_w11973_,
		_w24207_
	);
	LUT3 #(
		.INIT('h80)
	) name13695 (
		\wishbone_bd_ram_mem1_reg[96][10]/P0001 ,
		_w11941_,
		_w11965_,
		_w24208_
	);
	LUT4 #(
		.INIT('h0001)
	) name13696 (
		_w24205_,
		_w24206_,
		_w24207_,
		_w24208_,
		_w24209_
	);
	LUT4 #(
		.INIT('h8000)
	) name13697 (
		_w24194_,
		_w24199_,
		_w24204_,
		_w24209_,
		_w24210_
	);
	LUT4 #(
		.INIT('h8000)
	) name13698 (
		_w24147_,
		_w24168_,
		_w24189_,
		_w24210_,
		_w24211_
	);
	LUT3 #(
		.INIT('h80)
	) name13699 (
		\wishbone_bd_ram_mem1_reg[182][10]/P0001 ,
		_w11942_,
		_w11986_,
		_w24212_
	);
	LUT3 #(
		.INIT('h80)
	) name13700 (
		\wishbone_bd_ram_mem1_reg[9][10]/P0001 ,
		_w11932_,
		_w11968_,
		_w24213_
	);
	LUT3 #(
		.INIT('h80)
	) name13701 (
		\wishbone_bd_ram_mem1_reg[110][10]/P0001 ,
		_w11948_,
		_w11965_,
		_w24214_
	);
	LUT3 #(
		.INIT('h80)
	) name13702 (
		\wishbone_bd_ram_mem1_reg[85][10]/P0001 ,
		_w11933_,
		_w11972_,
		_w24215_
	);
	LUT4 #(
		.INIT('h0001)
	) name13703 (
		_w24212_,
		_w24213_,
		_w24214_,
		_w24215_,
		_w24216_
	);
	LUT3 #(
		.INIT('h80)
	) name13704 (
		\wishbone_bd_ram_mem1_reg[171][10]/P0001 ,
		_w11930_,
		_w11936_,
		_w24217_
	);
	LUT3 #(
		.INIT('h80)
	) name13705 (
		\wishbone_bd_ram_mem1_reg[72][10]/P0001 ,
		_w11949_,
		_w11990_,
		_w24218_
	);
	LUT3 #(
		.INIT('h80)
	) name13706 (
		\wishbone_bd_ram_mem1_reg[221][10]/P0001 ,
		_w11966_,
		_w11984_,
		_w24219_
	);
	LUT3 #(
		.INIT('h80)
	) name13707 (
		\wishbone_bd_ram_mem1_reg[227][10]/P0001 ,
		_w11938_,
		_w11982_,
		_w24220_
	);
	LUT4 #(
		.INIT('h0001)
	) name13708 (
		_w24217_,
		_w24218_,
		_w24219_,
		_w24220_,
		_w24221_
	);
	LUT3 #(
		.INIT('h80)
	) name13709 (
		\wishbone_bd_ram_mem1_reg[125][10]/P0001 ,
		_w11966_,
		_w12012_,
		_w24222_
	);
	LUT3 #(
		.INIT('h80)
	) name13710 (
		\wishbone_bd_ram_mem1_reg[153][10]/P0001 ,
		_w11959_,
		_w11968_,
		_w24223_
	);
	LUT3 #(
		.INIT('h80)
	) name13711 (
		\wishbone_bd_ram_mem1_reg[179][10]/P0001 ,
		_w11938_,
		_w11942_,
		_w24224_
	);
	LUT3 #(
		.INIT('h80)
	) name13712 (
		\wishbone_bd_ram_mem1_reg[129][10]/P0001 ,
		_w11955_,
		_w11977_,
		_w24225_
	);
	LUT4 #(
		.INIT('h0001)
	) name13713 (
		_w24222_,
		_w24223_,
		_w24224_,
		_w24225_,
		_w24226_
	);
	LUT3 #(
		.INIT('h80)
	) name13714 (
		\wishbone_bd_ram_mem1_reg[168][10]/P0001 ,
		_w11930_,
		_w11990_,
		_w24227_
	);
	LUT3 #(
		.INIT('h80)
	) name13715 (
		\wishbone_bd_ram_mem1_reg[143][10]/P0001 ,
		_w11955_,
		_w11973_,
		_w24228_
	);
	LUT3 #(
		.INIT('h80)
	) name13716 (
		\wishbone_bd_ram_mem1_reg[248][10]/P0001 ,
		_w11952_,
		_w11990_,
		_w24229_
	);
	LUT3 #(
		.INIT('h80)
	) name13717 (
		\wishbone_bd_ram_mem1_reg[51][10]/P0001 ,
		_w11938_,
		_w11979_,
		_w24230_
	);
	LUT4 #(
		.INIT('h0001)
	) name13718 (
		_w24227_,
		_w24228_,
		_w24229_,
		_w24230_,
		_w24231_
	);
	LUT4 #(
		.INIT('h8000)
	) name13719 (
		_w24216_,
		_w24221_,
		_w24226_,
		_w24231_,
		_w24232_
	);
	LUT3 #(
		.INIT('h80)
	) name13720 (
		\wishbone_bd_ram_mem1_reg[94][10]/P0001 ,
		_w11948_,
		_w11972_,
		_w24233_
	);
	LUT3 #(
		.INIT('h80)
	) name13721 (
		\wishbone_bd_ram_mem1_reg[50][10]/P0001 ,
		_w11963_,
		_w11979_,
		_w24234_
	);
	LUT3 #(
		.INIT('h80)
	) name13722 (
		\wishbone_bd_ram_mem1_reg[67][10]/P0001 ,
		_w11938_,
		_w11949_,
		_w24235_
	);
	LUT3 #(
		.INIT('h80)
	) name13723 (
		\wishbone_bd_ram_mem1_reg[84][10]/P0001 ,
		_w11929_,
		_w11972_,
		_w24236_
	);
	LUT4 #(
		.INIT('h0001)
	) name13724 (
		_w24233_,
		_w24234_,
		_w24235_,
		_w24236_,
		_w24237_
	);
	LUT3 #(
		.INIT('h80)
	) name13725 (
		\wishbone_bd_ram_mem1_reg[217][10]/P0001 ,
		_w11968_,
		_w11984_,
		_w24238_
	);
	LUT3 #(
		.INIT('h80)
	) name13726 (
		\wishbone_bd_ram_mem1_reg[87][10]/P0001 ,
		_w11972_,
		_w11975_,
		_w24239_
	);
	LUT3 #(
		.INIT('h80)
	) name13727 (
		\wishbone_bd_ram_mem1_reg[238][10]/P0001 ,
		_w11948_,
		_w11982_,
		_w24240_
	);
	LUT3 #(
		.INIT('h80)
	) name13728 (
		\wishbone_bd_ram_mem1_reg[55][10]/P0001 ,
		_w11975_,
		_w11979_,
		_w24241_
	);
	LUT4 #(
		.INIT('h0001)
	) name13729 (
		_w24238_,
		_w24239_,
		_w24240_,
		_w24241_,
		_w24242_
	);
	LUT3 #(
		.INIT('h80)
	) name13730 (
		\wishbone_bd_ram_mem1_reg[166][10]/P0001 ,
		_w11930_,
		_w11986_,
		_w24243_
	);
	LUT3 #(
		.INIT('h80)
	) name13731 (
		\wishbone_bd_ram_mem1_reg[95][10]/P0001 ,
		_w11972_,
		_w11973_,
		_w24244_
	);
	LUT3 #(
		.INIT('h80)
	) name13732 (
		\wishbone_bd_ram_mem1_reg[178][10]/P0001 ,
		_w11942_,
		_w11963_,
		_w24245_
	);
	LUT3 #(
		.INIT('h80)
	) name13733 (
		\wishbone_bd_ram_mem1_reg[25][10]/P0001 ,
		_w11935_,
		_w11968_,
		_w24246_
	);
	LUT4 #(
		.INIT('h0001)
	) name13734 (
		_w24243_,
		_w24244_,
		_w24245_,
		_w24246_,
		_w24247_
	);
	LUT3 #(
		.INIT('h80)
	) name13735 (
		\wishbone_bd_ram_mem1_reg[232][10]/P0001 ,
		_w11982_,
		_w11990_,
		_w24248_
	);
	LUT3 #(
		.INIT('h80)
	) name13736 (
		\wishbone_bd_ram_mem1_reg[46][10]/P0001 ,
		_w11948_,
		_w11957_,
		_w24249_
	);
	LUT3 #(
		.INIT('h80)
	) name13737 (
		\wishbone_bd_ram_mem1_reg[74][10]/P0001 ,
		_w11944_,
		_w11949_,
		_w24250_
	);
	LUT3 #(
		.INIT('h80)
	) name13738 (
		\wishbone_bd_ram_mem1_reg[214][10]/P0001 ,
		_w11984_,
		_w11986_,
		_w24251_
	);
	LUT4 #(
		.INIT('h0001)
	) name13739 (
		_w24248_,
		_w24249_,
		_w24250_,
		_w24251_,
		_w24252_
	);
	LUT4 #(
		.INIT('h8000)
	) name13740 (
		_w24237_,
		_w24242_,
		_w24247_,
		_w24252_,
		_w24253_
	);
	LUT3 #(
		.INIT('h80)
	) name13741 (
		\wishbone_bd_ram_mem1_reg[254][10]/P0001 ,
		_w11948_,
		_w11952_,
		_w24254_
	);
	LUT3 #(
		.INIT('h80)
	) name13742 (
		\wishbone_bd_ram_mem1_reg[6][10]/P0001 ,
		_w11932_,
		_w11986_,
		_w24255_
	);
	LUT3 #(
		.INIT('h80)
	) name13743 (
		\wishbone_bd_ram_mem1_reg[2][10]/P0001 ,
		_w11932_,
		_w11963_,
		_w24256_
	);
	LUT3 #(
		.INIT('h80)
	) name13744 (
		\wishbone_bd_ram_mem1_reg[8][10]/P0001 ,
		_w11932_,
		_w11990_,
		_w24257_
	);
	LUT4 #(
		.INIT('h0001)
	) name13745 (
		_w24254_,
		_w24255_,
		_w24256_,
		_w24257_,
		_w24258_
	);
	LUT3 #(
		.INIT('h80)
	) name13746 (
		\wishbone_bd_ram_mem1_reg[194][10]/P0001 ,
		_w11945_,
		_w11963_,
		_w24259_
	);
	LUT3 #(
		.INIT('h80)
	) name13747 (
		\wishbone_bd_ram_mem1_reg[231][10]/P0001 ,
		_w11975_,
		_w11982_,
		_w24260_
	);
	LUT3 #(
		.INIT('h80)
	) name13748 (
		\wishbone_bd_ram_mem1_reg[169][10]/P0001 ,
		_w11930_,
		_w11968_,
		_w24261_
	);
	LUT3 #(
		.INIT('h80)
	) name13749 (
		\wishbone_bd_ram_mem1_reg[105][10]/P0001 ,
		_w11965_,
		_w11968_,
		_w24262_
	);
	LUT4 #(
		.INIT('h0001)
	) name13750 (
		_w24259_,
		_w24260_,
		_w24261_,
		_w24262_,
		_w24263_
	);
	LUT3 #(
		.INIT('h80)
	) name13751 (
		\wishbone_bd_ram_mem1_reg[130][10]/P0001 ,
		_w11955_,
		_w11963_,
		_w24264_
	);
	LUT3 #(
		.INIT('h80)
	) name13752 (
		\wishbone_bd_ram_mem1_reg[186][10]/P0001 ,
		_w11942_,
		_w11944_,
		_w24265_
	);
	LUT3 #(
		.INIT('h80)
	) name13753 (
		\wishbone_bd_ram_mem1_reg[223][10]/P0001 ,
		_w11973_,
		_w11984_,
		_w24266_
	);
	LUT3 #(
		.INIT('h80)
	) name13754 (
		\wishbone_bd_ram_mem1_reg[144][10]/P0001 ,
		_w11941_,
		_w11959_,
		_w24267_
	);
	LUT4 #(
		.INIT('h0001)
	) name13755 (
		_w24264_,
		_w24265_,
		_w24266_,
		_w24267_,
		_w24268_
	);
	LUT3 #(
		.INIT('h80)
	) name13756 (
		\wishbone_bd_ram_mem1_reg[205][10]/P0001 ,
		_w11945_,
		_w11966_,
		_w24269_
	);
	LUT3 #(
		.INIT('h80)
	) name13757 (
		\wishbone_bd_ram_mem1_reg[150][10]/P0001 ,
		_w11959_,
		_w11986_,
		_w24270_
	);
	LUT3 #(
		.INIT('h80)
	) name13758 (
		\wishbone_bd_ram_mem1_reg[239][10]/P0001 ,
		_w11973_,
		_w11982_,
		_w24271_
	);
	LUT3 #(
		.INIT('h80)
	) name13759 (
		\wishbone_bd_ram_mem1_reg[172][10]/P0001 ,
		_w11930_,
		_w11954_,
		_w24272_
	);
	LUT4 #(
		.INIT('h0001)
	) name13760 (
		_w24269_,
		_w24270_,
		_w24271_,
		_w24272_,
		_w24273_
	);
	LUT4 #(
		.INIT('h8000)
	) name13761 (
		_w24258_,
		_w24263_,
		_w24268_,
		_w24273_,
		_w24274_
	);
	LUT3 #(
		.INIT('h80)
	) name13762 (
		\wishbone_bd_ram_mem1_reg[13][10]/P0001 ,
		_w11932_,
		_w11966_,
		_w24275_
	);
	LUT3 #(
		.INIT('h80)
	) name13763 (
		\wishbone_bd_ram_mem1_reg[45][10]/P0001 ,
		_w11957_,
		_w11966_,
		_w24276_
	);
	LUT3 #(
		.INIT('h80)
	) name13764 (
		\wishbone_bd_ram_mem1_reg[109][10]/P0001 ,
		_w11965_,
		_w11966_,
		_w24277_
	);
	LUT3 #(
		.INIT('h80)
	) name13765 (
		\wishbone_bd_ram_mem1_reg[63][10]/P0001 ,
		_w11973_,
		_w11979_,
		_w24278_
	);
	LUT4 #(
		.INIT('h0001)
	) name13766 (
		_w24275_,
		_w24276_,
		_w24277_,
		_w24278_,
		_w24279_
	);
	LUT3 #(
		.INIT('h80)
	) name13767 (
		\wishbone_bd_ram_mem1_reg[34][10]/P0001 ,
		_w11957_,
		_w11963_,
		_w24280_
	);
	LUT3 #(
		.INIT('h80)
	) name13768 (
		\wishbone_bd_ram_mem1_reg[198][10]/P0001 ,
		_w11945_,
		_w11986_,
		_w24281_
	);
	LUT3 #(
		.INIT('h80)
	) name13769 (
		\wishbone_bd_ram_mem1_reg[226][10]/P0001 ,
		_w11963_,
		_w11982_,
		_w24282_
	);
	LUT3 #(
		.INIT('h80)
	) name13770 (
		\wishbone_bd_ram_mem1_reg[244][10]/P0001 ,
		_w11929_,
		_w11952_,
		_w24283_
	);
	LUT4 #(
		.INIT('h0001)
	) name13771 (
		_w24280_,
		_w24281_,
		_w24282_,
		_w24283_,
		_w24284_
	);
	LUT3 #(
		.INIT('h80)
	) name13772 (
		\wishbone_bd_ram_mem1_reg[66][10]/P0001 ,
		_w11949_,
		_w11963_,
		_w24285_
	);
	LUT3 #(
		.INIT('h80)
	) name13773 (
		\wishbone_bd_ram_mem1_reg[192][10]/P0001 ,
		_w11941_,
		_w11945_,
		_w24286_
	);
	LUT3 #(
		.INIT('h80)
	) name13774 (
		\wishbone_bd_ram_mem1_reg[195][10]/P0001 ,
		_w11938_,
		_w11945_,
		_w24287_
	);
	LUT3 #(
		.INIT('h80)
	) name13775 (
		\wishbone_bd_ram_mem1_reg[160][10]/P0001 ,
		_w11930_,
		_w11941_,
		_w24288_
	);
	LUT4 #(
		.INIT('h0001)
	) name13776 (
		_w24285_,
		_w24286_,
		_w24287_,
		_w24288_,
		_w24289_
	);
	LUT3 #(
		.INIT('h80)
	) name13777 (
		\wishbone_bd_ram_mem1_reg[35][10]/P0001 ,
		_w11938_,
		_w11957_,
		_w24290_
	);
	LUT3 #(
		.INIT('h80)
	) name13778 (
		\wishbone_bd_ram_mem1_reg[173][10]/P0001 ,
		_w11930_,
		_w11966_,
		_w24291_
	);
	LUT3 #(
		.INIT('h80)
	) name13779 (
		\wishbone_bd_ram_mem1_reg[233][10]/P0001 ,
		_w11968_,
		_w11982_,
		_w24292_
	);
	LUT3 #(
		.INIT('h80)
	) name13780 (
		\wishbone_bd_ram_mem1_reg[40][10]/P0001 ,
		_w11957_,
		_w11990_,
		_w24293_
	);
	LUT4 #(
		.INIT('h0001)
	) name13781 (
		_w24290_,
		_w24291_,
		_w24292_,
		_w24293_,
		_w24294_
	);
	LUT4 #(
		.INIT('h8000)
	) name13782 (
		_w24279_,
		_w24284_,
		_w24289_,
		_w24294_,
		_w24295_
	);
	LUT4 #(
		.INIT('h8000)
	) name13783 (
		_w24232_,
		_w24253_,
		_w24274_,
		_w24295_,
		_w24296_
	);
	LUT3 #(
		.INIT('h80)
	) name13784 (
		\wishbone_bd_ram_mem1_reg[4][10]/P0001 ,
		_w11929_,
		_w11932_,
		_w24297_
	);
	LUT3 #(
		.INIT('h80)
	) name13785 (
		\wishbone_bd_ram_mem1_reg[190][10]/P0001 ,
		_w11942_,
		_w11948_,
		_w24298_
	);
	LUT3 #(
		.INIT('h80)
	) name13786 (
		\wishbone_bd_ram_mem1_reg[213][10]/P0001 ,
		_w11933_,
		_w11984_,
		_w24299_
	);
	LUT3 #(
		.INIT('h80)
	) name13787 (
		\wishbone_bd_ram_mem1_reg[101][10]/P0001 ,
		_w11933_,
		_w11965_,
		_w24300_
	);
	LUT4 #(
		.INIT('h0001)
	) name13788 (
		_w24297_,
		_w24298_,
		_w24299_,
		_w24300_,
		_w24301_
	);
	LUT3 #(
		.INIT('h80)
	) name13789 (
		\wishbone_bd_ram_mem1_reg[126][10]/P0001 ,
		_w11948_,
		_w12012_,
		_w24302_
	);
	LUT3 #(
		.INIT('h80)
	) name13790 (
		\wishbone_bd_ram_mem1_reg[207][10]/P0001 ,
		_w11945_,
		_w11973_,
		_w24303_
	);
	LUT3 #(
		.INIT('h80)
	) name13791 (
		\wishbone_bd_ram_mem1_reg[157][10]/P0001 ,
		_w11959_,
		_w11966_,
		_w24304_
	);
	LUT3 #(
		.INIT('h80)
	) name13792 (
		\wishbone_bd_ram_mem1_reg[19][10]/P0001 ,
		_w11935_,
		_w11938_,
		_w24305_
	);
	LUT4 #(
		.INIT('h0001)
	) name13793 (
		_w24302_,
		_w24303_,
		_w24304_,
		_w24305_,
		_w24306_
	);
	LUT3 #(
		.INIT('h80)
	) name13794 (
		\wishbone_bd_ram_mem1_reg[117][10]/P0001 ,
		_w11933_,
		_w12012_,
		_w24307_
	);
	LUT3 #(
		.INIT('h80)
	) name13795 (
		\wishbone_bd_ram_mem1_reg[142][10]/P0001 ,
		_w11948_,
		_w11955_,
		_w24308_
	);
	LUT3 #(
		.INIT('h80)
	) name13796 (
		\wishbone_bd_ram_mem1_reg[154][10]/P0001 ,
		_w11944_,
		_w11959_,
		_w24309_
	);
	LUT3 #(
		.INIT('h80)
	) name13797 (
		\wishbone_bd_ram_mem1_reg[156][10]/P0001 ,
		_w11954_,
		_w11959_,
		_w24310_
	);
	LUT4 #(
		.INIT('h0001)
	) name13798 (
		_w24307_,
		_w24308_,
		_w24309_,
		_w24310_,
		_w24311_
	);
	LUT3 #(
		.INIT('h80)
	) name13799 (
		\wishbone_bd_ram_mem1_reg[97][10]/P0001 ,
		_w11965_,
		_w11977_,
		_w24312_
	);
	LUT3 #(
		.INIT('h80)
	) name13800 (
		\wishbone_bd_ram_mem1_reg[16][10]/P0001 ,
		_w11935_,
		_w11941_,
		_w24313_
	);
	LUT3 #(
		.INIT('h80)
	) name13801 (
		\wishbone_bd_ram_mem1_reg[201][10]/P0001 ,
		_w11945_,
		_w11968_,
		_w24314_
	);
	LUT3 #(
		.INIT('h80)
	) name13802 (
		\wishbone_bd_ram_mem1_reg[59][10]/P0001 ,
		_w11936_,
		_w11979_,
		_w24315_
	);
	LUT4 #(
		.INIT('h0001)
	) name13803 (
		_w24312_,
		_w24313_,
		_w24314_,
		_w24315_,
		_w24316_
	);
	LUT4 #(
		.INIT('h8000)
	) name13804 (
		_w24301_,
		_w24306_,
		_w24311_,
		_w24316_,
		_w24317_
	);
	LUT3 #(
		.INIT('h80)
	) name13805 (
		\wishbone_bd_ram_mem1_reg[62][10]/P0001 ,
		_w11948_,
		_w11979_,
		_w24318_
	);
	LUT3 #(
		.INIT('h80)
	) name13806 (
		\wishbone_bd_ram_mem1_reg[75][10]/P0001 ,
		_w11936_,
		_w11949_,
		_w24319_
	);
	LUT3 #(
		.INIT('h80)
	) name13807 (
		\wishbone_bd_ram_mem1_reg[61][10]/P0001 ,
		_w11966_,
		_w11979_,
		_w24320_
	);
	LUT3 #(
		.INIT('h80)
	) name13808 (
		\wishbone_bd_ram_mem1_reg[211][10]/P0001 ,
		_w11938_,
		_w11984_,
		_w24321_
	);
	LUT4 #(
		.INIT('h0001)
	) name13809 (
		_w24318_,
		_w24319_,
		_w24320_,
		_w24321_,
		_w24322_
	);
	LUT3 #(
		.INIT('h80)
	) name13810 (
		\wishbone_bd_ram_mem1_reg[89][10]/P0001 ,
		_w11968_,
		_w11972_,
		_w24323_
	);
	LUT3 #(
		.INIT('h80)
	) name13811 (
		\wishbone_bd_ram_mem1_reg[218][10]/P0001 ,
		_w11944_,
		_w11984_,
		_w24324_
	);
	LUT3 #(
		.INIT('h80)
	) name13812 (
		\wishbone_bd_ram_mem1_reg[23][10]/P0001 ,
		_w11935_,
		_w11975_,
		_w24325_
	);
	LUT3 #(
		.INIT('h80)
	) name13813 (
		\wishbone_bd_ram_mem1_reg[11][10]/P0001 ,
		_w11932_,
		_w11936_,
		_w24326_
	);
	LUT4 #(
		.INIT('h0001)
	) name13814 (
		_w24323_,
		_w24324_,
		_w24325_,
		_w24326_,
		_w24327_
	);
	LUT3 #(
		.INIT('h80)
	) name13815 (
		\wishbone_bd_ram_mem1_reg[197][10]/P0001 ,
		_w11933_,
		_w11945_,
		_w24328_
	);
	LUT3 #(
		.INIT('h80)
	) name13816 (
		\wishbone_bd_ram_mem1_reg[36][10]/P0001 ,
		_w11929_,
		_w11957_,
		_w24329_
	);
	LUT3 #(
		.INIT('h80)
	) name13817 (
		\wishbone_bd_ram_mem1_reg[216][10]/P0001 ,
		_w11984_,
		_w11990_,
		_w24330_
	);
	LUT3 #(
		.INIT('h80)
	) name13818 (
		\wishbone_bd_ram_mem1_reg[26][10]/P0001 ,
		_w11935_,
		_w11944_,
		_w24331_
	);
	LUT4 #(
		.INIT('h0001)
	) name13819 (
		_w24328_,
		_w24329_,
		_w24330_,
		_w24331_,
		_w24332_
	);
	LUT3 #(
		.INIT('h80)
	) name13820 (
		\wishbone_bd_ram_mem1_reg[37][10]/P0001 ,
		_w11933_,
		_w11957_,
		_w24333_
	);
	LUT3 #(
		.INIT('h80)
	) name13821 (
		\wishbone_bd_ram_mem1_reg[57][10]/P0001 ,
		_w11968_,
		_w11979_,
		_w24334_
	);
	LUT3 #(
		.INIT('h80)
	) name13822 (
		\wishbone_bd_ram_mem1_reg[7][10]/P0001 ,
		_w11932_,
		_w11975_,
		_w24335_
	);
	LUT3 #(
		.INIT('h80)
	) name13823 (
		\wishbone_bd_ram_mem1_reg[108][10]/P0001 ,
		_w11954_,
		_w11965_,
		_w24336_
	);
	LUT4 #(
		.INIT('h0001)
	) name13824 (
		_w24333_,
		_w24334_,
		_w24335_,
		_w24336_,
		_w24337_
	);
	LUT4 #(
		.INIT('h8000)
	) name13825 (
		_w24322_,
		_w24327_,
		_w24332_,
		_w24337_,
		_w24338_
	);
	LUT3 #(
		.INIT('h80)
	) name13826 (
		\wishbone_bd_ram_mem1_reg[203][10]/P0001 ,
		_w11936_,
		_w11945_,
		_w24339_
	);
	LUT3 #(
		.INIT('h80)
	) name13827 (
		\wishbone_bd_ram_mem1_reg[121][10]/P0001 ,
		_w11968_,
		_w12012_,
		_w24340_
	);
	LUT3 #(
		.INIT('h80)
	) name13828 (
		\wishbone_bd_ram_mem1_reg[209][10]/P0001 ,
		_w11977_,
		_w11984_,
		_w24341_
	);
	LUT3 #(
		.INIT('h80)
	) name13829 (
		\wishbone_bd_ram_mem1_reg[91][10]/P0001 ,
		_w11936_,
		_w11972_,
		_w24342_
	);
	LUT4 #(
		.INIT('h0001)
	) name13830 (
		_w24339_,
		_w24340_,
		_w24341_,
		_w24342_,
		_w24343_
	);
	LUT3 #(
		.INIT('h80)
	) name13831 (
		\wishbone_bd_ram_mem1_reg[98][10]/P0001 ,
		_w11963_,
		_w11965_,
		_w24344_
	);
	LUT3 #(
		.INIT('h80)
	) name13832 (
		\wishbone_bd_ram_mem1_reg[237][10]/P0001 ,
		_w11966_,
		_w11982_,
		_w24345_
	);
	LUT3 #(
		.INIT('h80)
	) name13833 (
		\wishbone_bd_ram_mem1_reg[234][10]/P0001 ,
		_w11944_,
		_w11982_,
		_w24346_
	);
	LUT3 #(
		.INIT('h80)
	) name13834 (
		\wishbone_bd_ram_mem1_reg[47][10]/P0001 ,
		_w11957_,
		_w11973_,
		_w24347_
	);
	LUT4 #(
		.INIT('h0001)
	) name13835 (
		_w24344_,
		_w24345_,
		_w24346_,
		_w24347_,
		_w24348_
	);
	LUT3 #(
		.INIT('h80)
	) name13836 (
		\wishbone_bd_ram_mem1_reg[1][10]/P0001 ,
		_w11932_,
		_w11977_,
		_w24349_
	);
	LUT3 #(
		.INIT('h80)
	) name13837 (
		\wishbone_bd_ram_mem1_reg[135][10]/P0001 ,
		_w11955_,
		_w11975_,
		_w24350_
	);
	LUT3 #(
		.INIT('h80)
	) name13838 (
		\wishbone_bd_ram_mem1_reg[104][10]/P0001 ,
		_w11965_,
		_w11990_,
		_w24351_
	);
	LUT3 #(
		.INIT('h80)
	) name13839 (
		\wishbone_bd_ram_mem1_reg[176][10]/P0001 ,
		_w11941_,
		_w11942_,
		_w24352_
	);
	LUT4 #(
		.INIT('h0001)
	) name13840 (
		_w24349_,
		_w24350_,
		_w24351_,
		_w24352_,
		_w24353_
	);
	LUT3 #(
		.INIT('h80)
	) name13841 (
		\wishbone_bd_ram_mem1_reg[229][10]/P0001 ,
		_w11933_,
		_w11982_,
		_w24354_
	);
	LUT3 #(
		.INIT('h80)
	) name13842 (
		\wishbone_bd_ram_mem1_reg[170][10]/P0001 ,
		_w11930_,
		_w11944_,
		_w24355_
	);
	LUT3 #(
		.INIT('h80)
	) name13843 (
		\wishbone_bd_ram_mem1_reg[53][10]/P0001 ,
		_w11933_,
		_w11979_,
		_w24356_
	);
	LUT3 #(
		.INIT('h80)
	) name13844 (
		\wishbone_bd_ram_mem1_reg[185][10]/P0001 ,
		_w11942_,
		_w11968_,
		_w24357_
	);
	LUT4 #(
		.INIT('h0001)
	) name13845 (
		_w24354_,
		_w24355_,
		_w24356_,
		_w24357_,
		_w24358_
	);
	LUT4 #(
		.INIT('h8000)
	) name13846 (
		_w24343_,
		_w24348_,
		_w24353_,
		_w24358_,
		_w24359_
	);
	LUT3 #(
		.INIT('h80)
	) name13847 (
		\wishbone_bd_ram_mem1_reg[80][10]/P0001 ,
		_w11941_,
		_w11972_,
		_w24360_
	);
	LUT3 #(
		.INIT('h80)
	) name13848 (
		\wishbone_bd_ram_mem1_reg[138][10]/P0001 ,
		_w11944_,
		_w11955_,
		_w24361_
	);
	LUT3 #(
		.INIT('h80)
	) name13849 (
		\wishbone_bd_ram_mem1_reg[224][10]/P0001 ,
		_w11941_,
		_w11982_,
		_w24362_
	);
	LUT3 #(
		.INIT('h80)
	) name13850 (
		\wishbone_bd_ram_mem1_reg[174][10]/P0001 ,
		_w11930_,
		_w11948_,
		_w24363_
	);
	LUT4 #(
		.INIT('h0001)
	) name13851 (
		_w24360_,
		_w24361_,
		_w24362_,
		_w24363_,
		_w24364_
	);
	LUT3 #(
		.INIT('h80)
	) name13852 (
		\wishbone_bd_ram_mem1_reg[15][10]/P0001 ,
		_w11932_,
		_w11973_,
		_w24365_
	);
	LUT3 #(
		.INIT('h80)
	) name13853 (
		\wishbone_bd_ram_mem1_reg[5][10]/P0001 ,
		_w11932_,
		_w11933_,
		_w24366_
	);
	LUT3 #(
		.INIT('h80)
	) name13854 (
		\wishbone_bd_ram_mem1_reg[73][10]/P0001 ,
		_w11949_,
		_w11968_,
		_w24367_
	);
	LUT3 #(
		.INIT('h80)
	) name13855 (
		\wishbone_bd_ram_mem1_reg[114][10]/P0001 ,
		_w11963_,
		_w12012_,
		_w24368_
	);
	LUT4 #(
		.INIT('h0001)
	) name13856 (
		_w24365_,
		_w24366_,
		_w24367_,
		_w24368_,
		_w24369_
	);
	LUT3 #(
		.INIT('h80)
	) name13857 (
		\wishbone_bd_ram_mem1_reg[147][10]/P0001 ,
		_w11938_,
		_w11959_,
		_w24370_
	);
	LUT3 #(
		.INIT('h80)
	) name13858 (
		\wishbone_bd_ram_mem1_reg[167][10]/P0001 ,
		_w11930_,
		_w11975_,
		_w24371_
	);
	LUT3 #(
		.INIT('h80)
	) name13859 (
		\wishbone_bd_ram_mem1_reg[202][10]/P0001 ,
		_w11944_,
		_w11945_,
		_w24372_
	);
	LUT3 #(
		.INIT('h80)
	) name13860 (
		\wishbone_bd_ram_mem1_reg[115][10]/P0001 ,
		_w11938_,
		_w12012_,
		_w24373_
	);
	LUT4 #(
		.INIT('h0001)
	) name13861 (
		_w24370_,
		_w24371_,
		_w24372_,
		_w24373_,
		_w24374_
	);
	LUT3 #(
		.INIT('h80)
	) name13862 (
		\wishbone_bd_ram_mem1_reg[123][10]/P0001 ,
		_w11936_,
		_w12012_,
		_w24375_
	);
	LUT3 #(
		.INIT('h80)
	) name13863 (
		\wishbone_bd_ram_mem1_reg[152][10]/P0001 ,
		_w11959_,
		_w11990_,
		_w24376_
	);
	LUT3 #(
		.INIT('h80)
	) name13864 (
		\wishbone_bd_ram_mem1_reg[69][10]/P0001 ,
		_w11933_,
		_w11949_,
		_w24377_
	);
	LUT3 #(
		.INIT('h80)
	) name13865 (
		\wishbone_bd_ram_mem1_reg[68][10]/P0001 ,
		_w11929_,
		_w11949_,
		_w24378_
	);
	LUT4 #(
		.INIT('h0001)
	) name13866 (
		_w24375_,
		_w24376_,
		_w24377_,
		_w24378_,
		_w24379_
	);
	LUT4 #(
		.INIT('h8000)
	) name13867 (
		_w24364_,
		_w24369_,
		_w24374_,
		_w24379_,
		_w24380_
	);
	LUT4 #(
		.INIT('h8000)
	) name13868 (
		_w24317_,
		_w24338_,
		_w24359_,
		_w24380_,
		_w24381_
	);
	LUT4 #(
		.INIT('h8000)
	) name13869 (
		_w24126_,
		_w24211_,
		_w24296_,
		_w24381_,
		_w24382_
	);
	LUT3 #(
		.INIT('h3b)
	) name13870 (
		_w19180_,
		_w24041_,
		_w24382_,
		_w24383_
	);
	LUT4 #(
		.INIT('h060c)
	) name13871 (
		\wishbone_TxPointerMSB_reg[10]/NET0131 ,
		\wishbone_TxPointerMSB_reg[11]/NET0131 ,
		_w15303_,
		_w15308_,
		_w24384_
	);
	LUT3 #(
		.INIT('hf2)
	) name13872 (
		_w19180_,
		_w22213_,
		_w24384_,
		_w24385_
	);
	LUT3 #(
		.INIT('hed)
	) name13873 (
		\wishbone_TxPointerMSB_reg[13]/NET0131 ,
		_w15303_,
		_w15310_,
		_w24386_
	);
	LUT3 #(
		.INIT('h2f)
	) name13874 (
		_w19180_,
		_w23589_,
		_w24386_,
		_w24387_
	);
	LUT3 #(
		.INIT('h80)
	) name13875 (
		\wishbone_TxPointerMSB_reg[13]/NET0131 ,
		\wishbone_TxPointerMSB_reg[14]/NET0131 ,
		\wishbone_TxPointerMSB_reg[15]/NET0131 ,
		_w24388_
	);
	LUT4 #(
		.INIT('h1222)
	) name13876 (
		\wishbone_TxPointerMSB_reg[15]/NET0131 ,
		_w15303_,
		_w15310_,
		_w15312_,
		_w24389_
	);
	LUT3 #(
		.INIT('hf4)
	) name13877 (
		_w13800_,
		_w19180_,
		_w24389_,
		_w24390_
	);
	LUT3 #(
		.INIT('h15)
	) name13878 (
		\wishbone_TxPointerMSB_reg[16]/NET0131 ,
		_w15310_,
		_w24388_,
		_w24391_
	);
	LUT4 #(
		.INIT('h8000)
	) name13879 (
		\wishbone_TxPointerMSB_reg[13]/NET0131 ,
		\wishbone_TxPointerMSB_reg[14]/NET0131 ,
		\wishbone_TxPointerMSB_reg[15]/NET0131 ,
		\wishbone_TxPointerMSB_reg[16]/NET0131 ,
		_w24392_
	);
	LUT3 #(
		.INIT('h15)
	) name13880 (
		_w15303_,
		_w15310_,
		_w24392_,
		_w24393_
	);
	LUT2 #(
		.INIT('h4)
	) name13881 (
		_w24391_,
		_w24393_,
		_w24394_
	);
	LUT3 #(
		.INIT('hf4)
	) name13882 (
		_w16122_,
		_w19180_,
		_w24394_,
		_w24395_
	);
	LUT3 #(
		.INIT('h15)
	) name13883 (
		\wishbone_TxPointerMSB_reg[17]/NET0131 ,
		_w15310_,
		_w24392_,
		_w24396_
	);
	LUT3 #(
		.INIT('h15)
	) name13884 (
		_w15303_,
		_w15310_,
		_w15314_,
		_w24397_
	);
	LUT2 #(
		.INIT('h4)
	) name13885 (
		_w24396_,
		_w24397_,
		_w24398_
	);
	LUT3 #(
		.INIT('hf4)
	) name13886 (
		_w16814_,
		_w19180_,
		_w24398_,
		_w24399_
	);
	LUT4 #(
		.INIT('heddd)
	) name13887 (
		\wishbone_TxPointerMSB_reg[18]/NET0131 ,
		_w15303_,
		_w15310_,
		_w15314_,
		_w24400_
	);
	LUT3 #(
		.INIT('h4f)
	) name13888 (
		_w15775_,
		_w19180_,
		_w24400_,
		_w24401_
	);
	LUT3 #(
		.INIT('h12)
	) name13889 (
		\wishbone_TxPointerMSB_reg[2]/NET0131 ,
		_w15303_,
		_w15304_,
		_w24402_
	);
	LUT3 #(
		.INIT('hf2)
	) name13890 (
		_w19180_,
		_w22594_,
		_w24402_,
		_w24403_
	);
	LUT4 #(
		.INIT('h00bf)
	) name13891 (
		\wishbone_BlockingIncrementTxPointer_reg/NET0131 ,
		\wishbone_IncrTxPointer_reg/NET0131 ,
		\wishbone_TxPointerMSB_reg[2]/NET0131 ,
		\wishbone_TxPointerMSB_reg[3]/NET0131 ,
		_w24404_
	);
	LUT3 #(
		.INIT('h01)
	) name13892 (
		_w15303_,
		_w15305_,
		_w24404_,
		_w24405_
	);
	LUT3 #(
		.INIT('hf2)
	) name13893 (
		_w19180_,
		_w20008_,
		_w24405_,
		_w24406_
	);
	LUT4 #(
		.INIT('h1333)
	) name13894 (
		\wishbone_TxPointerMSB_reg[7]/NET0131 ,
		\wishbone_TxPointerMSB_reg[8]/NET0131 ,
		_w15305_,
		_w15306_,
		_w24407_
	);
	LUT4 #(
		.INIT('h1555)
	) name13895 (
		_w15303_,
		_w15305_,
		_w15306_,
		_w23226_,
		_w24408_
	);
	LUT2 #(
		.INIT('h4)
	) name13896 (
		_w24407_,
		_w24408_,
		_w24409_
	);
	LUT3 #(
		.INIT('hf2)
	) name13897 (
		_w19180_,
		_w21480_,
		_w24409_,
		_w24410_
	);
	LUT4 #(
		.INIT('h0001)
	) name13898 (
		\miim1_clkgen_Counter_reg[0]/NET0131 ,
		\miim1_clkgen_Counter_reg[1]/NET0131 ,
		\miim1_clkgen_Counter_reg[2]/NET0131 ,
		\miim1_clkgen_Counter_reg[3]/NET0131 ,
		_w24411_
	);
	LUT2 #(
		.INIT('h9)
	) name13899 (
		\miim1_clkgen_Counter_reg[4]/NET0131 ,
		_w24411_,
		_w24412_
	);
	LUT2 #(
		.INIT('h1)
	) name13900 (
		\ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131 ,
		_w24413_
	);
	LUT2 #(
		.INIT('h1)
	) name13901 (
		\ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131 ,
		_w24414_
	);
	LUT4 #(
		.INIT('h0001)
	) name13902 (
		\ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131 ,
		_w24415_
	);
	LUT3 #(
		.INIT('h01)
	) name13903 (
		\ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131 ,
		_w24416_
	);
	LUT2 #(
		.INIT('h4)
	) name13904 (
		_w24415_,
		_w24416_,
		_w24417_
	);
	LUT4 #(
		.INIT('h88cc)
	) name13905 (
		\ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131 ,
		_w24414_,
		_w24416_,
		_w24418_
	);
	LUT3 #(
		.INIT('h20)
	) name13906 (
		_w24413_,
		_w24414_,
		_w24416_,
		_w24419_
	);
	LUT3 #(
		.INIT('h01)
	) name13907 (
		\miim1_clkgen_Counter_reg[4]/NET0131 ,
		\miim1_clkgen_Counter_reg[5]/NET0131 ,
		\miim1_clkgen_Counter_reg[6]/NET0131 ,
		_w24420_
	);
	LUT2 #(
		.INIT('h8)
	) name13908 (
		_w24411_,
		_w24420_,
		_w24421_
	);
	LUT4 #(
		.INIT('h5455)
	) name13909 (
		_w24412_,
		_w24418_,
		_w24419_,
		_w24421_,
		_w24422_
	);
	LUT3 #(
		.INIT('h80)
	) name13910 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w24423_
	);
	LUT2 #(
		.INIT('h8)
	) name13911 (
		\wishbone_LastByteIn_reg/NET0131 ,
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		_w24424_
	);
	LUT2 #(
		.INIT('h8)
	) name13912 (
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w24425_
	);
	LUT4 #(
		.INIT('h8000)
	) name13913 (
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		\wishbone_RxEnableWindow_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w24426_
	);
	LUT3 #(
		.INIT('h80)
	) name13914 (
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_RxEnableWindow_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w24427_
	);
	LUT4 #(
		.INIT('h3666)
	) name13915 (
		\wishbone_LastByteIn_reg/NET0131 ,
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		\wishbone_RxEnableWindow_reg/NET0131 ,
		_w24425_,
		_w24428_
	);
	LUT2 #(
		.INIT('h1)
	) name13916 (
		\RxAbort_wb_reg/NET0131 ,
		\wishbone_ShiftEnded_rck_reg/NET0131 ,
		_w24429_
	);
	LUT2 #(
		.INIT('h4)
	) name13917 (
		_w13420_,
		_w24429_,
		_w24430_
	);
	LUT3 #(
		.INIT('he0)
	) name13918 (
		_w24423_,
		_w24428_,
		_w24430_,
		_w24431_
	);
	LUT3 #(
		.INIT('h60)
	) name13919 (
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		_w13032_,
		_w13040_,
		_w24432_
	);
	LUT4 #(
		.INIT('hc400)
	) name13920 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131 ,
		\maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w24433_
	);
	LUT2 #(
		.INIT('h8)
	) name13921 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		_w24434_
	);
	LUT2 #(
		.INIT('h8)
	) name13922 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		_w24435_
	);
	LUT4 #(
		.INIT('h1555)
	) name13923 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131 ,
		_w24433_,
		_w24434_,
		_w24435_,
		_w24436_
	);
	LUT3 #(
		.INIT('h80)
	) name13924 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131 ,
		_w24437_
	);
	LUT4 #(
		.INIT('h1555)
	) name13925 (
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		_w24433_,
		_w24434_,
		_w24437_,
		_w24438_
	);
	LUT2 #(
		.INIT('h4)
	) name13926 (
		_w24436_,
		_w24438_,
		_w24439_
	);
	LUT4 #(
		.INIT('hddde)
	) name13927 (
		\wishbone_RxByteCnt_reg[1]/NET0131 ,
		_w24423_,
		_w24424_,
		_w24426_,
		_w24440_
	);
	LUT2 #(
		.INIT('h9)
	) name13928 (
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w24441_
	);
	LUT3 #(
		.INIT('h4c)
	) name13929 (
		_w24423_,
		_w24429_,
		_w24441_,
		_w24442_
	);
	LUT2 #(
		.INIT('h8)
	) name13930 (
		_w24440_,
		_w24442_,
		_w24443_
	);
	LUT3 #(
		.INIT('h10)
	) name13931 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131 ,
		_w24444_
	);
	LUT4 #(
		.INIT('h4000)
	) name13932 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w24445_
	);
	LUT4 #(
		.INIT('h5111)
	) name13933 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		_w24433_,
		_w24444_,
		_w24445_,
		_w24446_
	);
	LUT3 #(
		.INIT('h13)
	) name13934 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		_w24433_,
		_w24447_
	);
	LUT2 #(
		.INIT('h4)
	) name13935 (
		_w24446_,
		_w24447_,
		_w24448_
	);
	LUT4 #(
		.INIT('h1222)
	) name13936 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		_w24433_,
		_w24434_,
		_w24449_
	);
	LUT4 #(
		.INIT('h1333)
	) name13937 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		_w24433_,
		_w24434_,
		_w24450_
	);
	LUT4 #(
		.INIT('h1555)
	) name13938 (
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		_w24433_,
		_w24434_,
		_w24435_,
		_w24451_
	);
	LUT2 #(
		.INIT('h4)
	) name13939 (
		_w24450_,
		_w24451_,
		_w24452_
	);
	LUT4 #(
		.INIT('h6a00)
	) name13940 (
		\txethmac1_txcounters1_ByteCnt_reg[10]/NET0131 ,
		_w13034_,
		_w13036_,
		_w13040_,
		_w24453_
	);
	LUT4 #(
		.INIT('h1555)
	) name13941 (
		\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 ,
		_w13027_,
		_w13034_,
		_w13036_,
		_w24454_
	);
	LUT3 #(
		.INIT('h80)
	) name13942 (
		\txethmac1_txcounters1_ByteCnt_reg[10]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[11]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 ,
		_w24455_
	);
	LUT4 #(
		.INIT('h70f0)
	) name13943 (
		_w13034_,
		_w13036_,
		_w13040_,
		_w24455_,
		_w24456_
	);
	LUT2 #(
		.INIT('h4)
	) name13944 (
		_w24454_,
		_w24456_,
		_w24457_
	);
	LUT2 #(
		.INIT('h8)
	) name13945 (
		\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 ,
		_w13029_,
		_w24458_
	);
	LUT3 #(
		.INIT('h80)
	) name13946 (
		\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[13]/NET0131 ,
		_w13029_,
		_w24459_
	);
	LUT4 #(
		.INIT('h60a0)
	) name13947 (
		\txethmac1_txcounters1_ByteCnt_reg[13]/NET0131 ,
		_w13032_,
		_w13040_,
		_w24458_,
		_w24460_
	);
	LUT3 #(
		.INIT('h15)
	) name13948 (
		\txethmac1_txcounters1_ByteCnt_reg[14]/NET0131 ,
		_w13032_,
		_w24459_,
		_w24461_
	);
	LUT2 #(
		.INIT('h8)
	) name13949 (
		\txethmac1_txcounters1_ByteCnt_reg[13]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[14]/NET0131 ,
		_w24462_
	);
	LUT3 #(
		.INIT('h80)
	) name13950 (
		\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 ,
		_w13029_,
		_w24462_,
		_w24463_
	);
	LUT3 #(
		.INIT('h4c)
	) name13951 (
		_w13032_,
		_w13040_,
		_w24463_,
		_w24464_
	);
	LUT2 #(
		.INIT('h4)
	) name13952 (
		_w24461_,
		_w24464_,
		_w24465_
	);
	LUT4 #(
		.INIT('h0444)
	) name13953 (
		_w13022_,
		_w13025_,
		_w13029_,
		_w13031_,
		_w24466_
	);
	LUT4 #(
		.INIT('h6c00)
	) name13954 (
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		_w13032_,
		_w13040_,
		_w24467_
	);
	LUT4 #(
		.INIT('h3020)
	) name13955 (
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		_w13034_,
		_w13040_,
		_w24466_,
		_w24468_
	);
	LUT4 #(
		.INIT('h0004)
	) name13956 (
		\txethmac1_PacketFinished_q_reg/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		_w10936_,
		_w10937_,
		_w24469_
	);
	LUT3 #(
		.INIT('h70)
	) name13957 (
		_w10791_,
		_w10967_,
		_w24469_,
		_w24470_
	);
	LUT4 #(
		.INIT('h0001)
	) name13958 (
		\txethmac1_PacketFinished_q_reg/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		_w10936_,
		_w10937_,
		_w24471_
	);
	LUT3 #(
		.INIT('h70)
	) name13959 (
		_w10791_,
		_w10967_,
		_w24471_,
		_w24472_
	);
	LUT3 #(
		.INIT('he4)
	) name13960 (
		_w13034_,
		_w24470_,
		_w24472_,
		_w24473_
	);
	LUT2 #(
		.INIT('h8)
	) name13961 (
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w24474_
	);
	LUT4 #(
		.INIT('h6c00)
	) name13962 (
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w13034_,
		_w13040_,
		_w24475_
	);
	LUT3 #(
		.INIT('h15)
	) name13963 (
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		_w13034_,
		_w24474_,
		_w24476_
	);
	LUT3 #(
		.INIT('h80)
	) name13964 (
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		_w24477_
	);
	LUT3 #(
		.INIT('h4c)
	) name13965 (
		_w13034_,
		_w13040_,
		_w24477_,
		_w24478_
	);
	LUT2 #(
		.INIT('h4)
	) name13966 (
		_w24476_,
		_w24478_,
		_w24479_
	);
	LUT4 #(
		.INIT('h60a0)
	) name13967 (
		\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 ,
		_w13034_,
		_w13040_,
		_w24477_,
		_w24480_
	);
	LUT4 #(
		.INIT('h1333)
	) name13968 (
		\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[7]/NET0131 ,
		_w13034_,
		_w24477_,
		_w24481_
	);
	LUT4 #(
		.INIT('h70f0)
	) name13969 (
		_w13023_,
		_w13034_,
		_w13040_,
		_w24477_,
		_w24482_
	);
	LUT2 #(
		.INIT('h4)
	) name13970 (
		_w24481_,
		_w24482_,
		_w24483_
	);
	LUT4 #(
		.INIT('h1555)
	) name13971 (
		\txethmac1_txcounters1_ByteCnt_reg[8]/NET0131 ,
		_w13023_,
		_w13034_,
		_w24477_,
		_w24484_
	);
	LUT3 #(
		.INIT('h80)
	) name13972 (
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		_w13023_,
		_w13024_,
		_w24485_
	);
	LUT3 #(
		.INIT('h4c)
	) name13973 (
		_w13034_,
		_w13040_,
		_w24485_,
		_w24486_
	);
	LUT2 #(
		.INIT('h4)
	) name13974 (
		_w24484_,
		_w24486_,
		_w24487_
	);
	LUT3 #(
		.INIT('h80)
	) name13975 (
		_w13023_,
		_w13024_,
		_w13026_,
		_w24488_
	);
	LUT4 #(
		.INIT('h1500)
	) name13976 (
		_w13022_,
		_w13029_,
		_w13031_,
		_w24488_,
		_w24489_
	);
	LUT4 #(
		.INIT('h8000)
	) name13977 (
		\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 ,
		_w13023_,
		_w13024_,
		_w13026_,
		_w24490_
	);
	LUT4 #(
		.INIT('h1500)
	) name13978 (
		_w13022_,
		_w13029_,
		_w13031_,
		_w24490_,
		_w24491_
	);
	LUT4 #(
		.INIT('h00c8)
	) name13979 (
		\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 ,
		_w13040_,
		_w24489_,
		_w24491_,
		_w24492_
	);
	LUT4 #(
		.INIT('h1000)
	) name13980 (
		\txethmac1_txcrc_Crc_reg[3]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11776_,
		_w11779_,
		_w24493_
	);
	LUT3 #(
		.INIT('h40)
	) name13981 (
		\txethmac1_txcrc_Crc_reg[3]/NET0131 ,
		_w10913_,
		_w10914_,
		_w24494_
	);
	LUT3 #(
		.INIT('hcd)
	) name13982 (
		_w11782_,
		_w24493_,
		_w24494_,
		_w24495_
	);
	LUT2 #(
		.INIT('h1)
	) name13983 (
		\txethmac1_txcrc_Crc_reg[2]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w24496_
	);
	LUT3 #(
		.INIT('h60)
	) name13984 (
		_w11105_,
		_w11106_,
		_w24496_,
		_w24497_
	);
	LUT3 #(
		.INIT('h40)
	) name13985 (
		\txethmac1_txcrc_Crc_reg[2]/NET0131 ,
		_w10913_,
		_w10914_,
		_w24498_
	);
	LUT4 #(
		.INIT('h090f)
	) name13986 (
		_w11105_,
		_w11106_,
		_w24498_,
		_w11110_,
		_w24499_
	);
	LUT2 #(
		.INIT('he)
	) name13987 (
		_w24497_,
		_w24499_,
		_w24500_
	);
	LUT3 #(
		.INIT('h0e)
	) name13988 (
		m_wb_ack_i_pad,
		m_wb_err_i_pad,
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w24501_
	);
	LUT3 #(
		.INIT('he1)
	) name13989 (
		m_wb_ack_i_pad,
		m_wb_err_i_pad,
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w24502_
	);
	LUT4 #(
		.INIT('h000b)
	) name13990 (
		\wishbone_BlockReadTxDataFromMemory_reg/NET0131 ,
		\wishbone_ReadTxDataFromMemory_reg/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[4]/NET0131 ,
		_w24503_
	);
	LUT2 #(
		.INIT('h8)
	) name13991 (
		_w11866_,
		_w24503_,
		_w24504_
	);
	LUT3 #(
		.INIT('h20)
	) name13992 (
		_w11866_,
		_w24502_,
		_w24503_,
		_w24505_
	);
	LUT2 #(
		.INIT('h1)
	) name13993 (
		_w11893_,
		_w11898_,
		_w24506_
	);
	LUT4 #(
		.INIT('h8000)
	) name13994 (
		_w11866_,
		_w11892_,
		_w11893_,
		_w24503_,
		_w24507_
	);
	LUT2 #(
		.INIT('h4)
	) name13995 (
		_w11892_,
		_w24502_,
		_w24508_
	);
	LUT4 #(
		.INIT('h000b)
	) name13996 (
		_w24505_,
		_w24506_,
		_w24507_,
		_w24508_,
		_w24509_
	);
	LUT2 #(
		.INIT('h8)
	) name13997 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_rx_burst_en_reg/NET0131 ,
		_w24510_
	);
	LUT3 #(
		.INIT('h70)
	) name13998 (
		_w11866_,
		_w11867_,
		_w24510_,
		_w24511_
	);
	LUT4 #(
		.INIT('h1000)
	) name13999 (
		\wishbone_BlockReadTxDataFromMemory_reg/NET0131 ,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_ReadTxDataFromMemory_reg/NET0131 ,
		\wishbone_tx_burst_en_reg/NET0131 ,
		_w24512_
	);
	LUT3 #(
		.INIT('h08)
	) name14000 (
		_w11898_,
		_w24501_,
		_w24512_,
		_w24513_
	);
	LUT3 #(
		.INIT('h10)
	) name14001 (
		_w24504_,
		_w24511_,
		_w24513_,
		_w24514_
	);
	LUT4 #(
		.INIT('h3233)
	) name14002 (
		_w24504_,
		_w24505_,
		_w24511_,
		_w24513_,
		_w24515_
	);
	LUT3 #(
		.INIT('h2a)
	) name14003 (
		\m_wb_sel_o[0]_pad ,
		_w24509_,
		_w24515_,
		_w24516_
	);
	LUT2 #(
		.INIT('hd)
	) name14004 (
		_w11907_,
		_w24516_,
		_w24517_
	);
	LUT2 #(
		.INIT('h2)
	) name14005 (
		\macstatus1_InvalidSymbol_reg/NET0131 ,
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		_w24518_
	);
	LUT4 #(
		.INIT('h13df)
	) name14006 (
		\RxEnSync_reg/NET0131 ,
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		mrxerr_pad_i_pad,
		mtxerr_pad_o_pad,
		_w24519_
	);
	LUT2 #(
		.INIT('h1)
	) name14007 (
		_w10576_,
		_w24519_,
		_w24520_
	);
	LUT4 #(
		.INIT('h0100)
	) name14008 (
		_w10578_,
		_w10588_,
		_w10943_,
		_w11045_,
		_w24521_
	);
	LUT3 #(
		.INIT('hea)
	) name14009 (
		_w24518_,
		_w24520_,
		_w24521_,
		_w24522_
	);
	LUT3 #(
		.INIT('h70)
	) name14010 (
		\wishbone_ShiftEndedSync_c1_reg/NET0131 ,
		\wishbone_ShiftEndedSync_c2_reg/NET0131 ,
		\wishbone_ShiftEnded_rck_reg/NET0131 ,
		_w24523_
	);
	LUT2 #(
		.INIT('h8)
	) name14011 (
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w24524_
	);
	LUT3 #(
		.INIT('h80)
	) name14012 (
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		\wishbone_RxByteCnt_reg[1]/NET0131 ,
		\wishbone_RxEnableWindow_reg/NET0131 ,
		_w24525_
	);
	LUT4 #(
		.INIT('h0111)
	) name14013 (
		\wishbone_LastByteIn_reg/NET0131 ,
		_w24523_,
		_w24524_,
		_w24525_,
		_w24526_
	);
	LUT2 #(
		.INIT('h1)
	) name14014 (
		_w13424_,
		_w24523_,
		_w24527_
	);
	LUT4 #(
		.INIT('h0105)
	) name14015 (
		\RxAbort_wb_reg/NET0131 ,
		_w13423_,
		_w24526_,
		_w24527_,
		_w24528_
	);
	LUT4 #(
		.INIT('h060c)
	) name14016 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		_w24433_,
		_w24529_
	);
	LUT2 #(
		.INIT('h2)
	) name14017 (
		m_wb_stb_o_pad,
		_w24509_,
		_w24530_
	);
	LUT2 #(
		.INIT('hd)
	) name14018 (
		_w11907_,
		_w24530_,
		_w24531_
	);
	LUT3 #(
		.INIT('h08)
	) name14019 (
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w24532_
	);
	LUT4 #(
		.INIT('h008f)
	) name14020 (
		_w11866_,
		_w11867_,
		_w11883_,
		_w24532_,
		_w24533_
	);
	LUT3 #(
		.INIT('h20)
	) name14021 (
		\wishbone_tx_burst_en_reg/NET0131 ,
		_w11882_,
		_w24533_,
		_w24534_
	);
	LUT4 #(
		.INIT('h3233)
	) name14022 (
		_w24504_,
		_w24507_,
		_w24511_,
		_w24513_,
		_w24535_
	);
	LUT3 #(
		.INIT('ha8)
	) name14023 (
		\wishbone_tx_burst_en_reg/NET0131 ,
		_w11882_,
		_w11884_,
		_w24536_
	);
	LUT2 #(
		.INIT('h8)
	) name14024 (
		\wishbone_TxLength_reg[3]/NET0131 ,
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w24537_
	);
	LUT4 #(
		.INIT('he000)
	) name14025 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		\wishbone_TxLength_reg[2]/NET0131 ,
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w24538_
	);
	LUT2 #(
		.INIT('h1)
	) name14026 (
		_w24537_,
		_w24538_,
		_w24539_
	);
	LUT4 #(
		.INIT('h8000)
	) name14027 (
		_w12307_,
		_w12310_,
		_w12314_,
		_w12316_,
		_w24540_
	);
	LUT3 #(
		.INIT('h07)
	) name14028 (
		\wishbone_tx_fifo_cnt_reg[2]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w24541_
	);
	LUT3 #(
		.INIT('h70)
	) name14029 (
		_w24539_,
		_w24540_,
		_w24541_,
		_w24542_
	);
	LUT4 #(
		.INIT('hfbea)
	) name14030 (
		_w24534_,
		_w24535_,
		_w24536_,
		_w24542_,
		_w24543_
	);
	LUT4 #(
		.INIT('hcfef)
	) name14031 (
		\wishbone_IncrTxPointer_reg/NET0131 ,
		_w11890_,
		_w11900_,
		_w24509_,
		_w24544_
	);
	LUT3 #(
		.INIT('h80)
	) name14032 (
		_w11891_,
		_w11897_,
		_w11898_,
		_w24545_
	);
	LUT2 #(
		.INIT('h4)
	) name14033 (
		_w11896_,
		_w24545_,
		_w24546_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name14034 (
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w11866_,
		_w11868_,
		_w24503_,
		_w24547_
	);
	LUT3 #(
		.INIT('h70)
	) name14035 (
		_w11903_,
		_w11904_,
		_w24547_,
		_w24548_
	);
	LUT4 #(
		.INIT('h0100)
	) name14036 (
		_w11890_,
		_w11902_,
		_w24546_,
		_w24548_,
		_w24549_
	);
	LUT2 #(
		.INIT('he)
	) name14037 (
		_w24514_,
		_w24549_,
		_w24550_
	);
	LUT2 #(
		.INIT('h1)
	) name14038 (
		\txethmac1_StatusLatch_reg/NET0131 ,
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		_w24551_
	);
	LUT4 #(
		.INIT('h2033)
	) name14039 (
		_w10834_,
		_w10836_,
		_w10975_,
		_w24551_,
		_w24552_
	);
	LUT4 #(
		.INIT('h0001)
	) name14040 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		\rxethmac1_rxstatem1_StatePreamble_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w24553_
	);
	LUT4 #(
		.INIT('h0405)
	) name14041 (
		_w10576_,
		_w11562_,
		_w24519_,
		_w24553_,
		_w24554_
	);
	LUT2 #(
		.INIT('h4)
	) name14042 (
		\wishbone_WriteRxDataToFifoSync2_reg/NET0131 ,
		\wishbone_WriteRxDataToFifo_reg/NET0131 ,
		_w24555_
	);
	LUT2 #(
		.INIT('h1)
	) name14043 (
		_w13424_,
		_w24555_,
		_w24556_
	);
	LUT3 #(
		.INIT('h15)
	) name14044 (
		\RxAbort_wb_reg/NET0131 ,
		_w13423_,
		_w24556_,
		_w24557_
	);
	LUT4 #(
		.INIT('h01fe)
	) name14045 (
		\miim1_clkgen_Counter_reg[0]/NET0131 ,
		\miim1_clkgen_Counter_reg[1]/NET0131 ,
		\miim1_clkgen_Counter_reg[2]/NET0131 ,
		\miim1_clkgen_Counter_reg[3]/NET0131 ,
		_w24558_
	);
	LUT3 #(
		.INIT('h70)
	) name14046 (
		_w24411_,
		_w24420_,
		_w24558_,
		_w24559_
	);
	LUT4 #(
		.INIT('h006f)
	) name14047 (
		\ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131 ,
		_w24417_,
		_w24421_,
		_w24559_,
		_w24560_
	);
	LUT3 #(
		.INIT('h80)
	) name14048 (
		mdc_pad_o_pad,
		_w24411_,
		_w24420_,
		_w24561_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name14049 (
		mdc_pad_o_pad,
		\miim1_shftrg_ShiftReg_reg[1]/NET0131 ,
		_w24411_,
		_w24420_,
		_w24562_
	);
	LUT4 #(
		.INIT('h1333)
	) name14050 (
		mdc_pad_o_pad,
		\miim1_shftrg_ShiftReg_reg[1]/NET0131 ,
		_w24411_,
		_w24420_,
		_w24563_
	);
	LUT4 #(
		.INIT('h0002)
	) name14051 (
		\ethreg1_MIIMODER_1_DataOut_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[2]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		\miim1_BitCounter_reg[4]/NET0131 ,
		_w24564_
	);
	LUT4 #(
		.INIT('h0001)
	) name14052 (
		\miim1_BitCounter_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[1]/NET0131 ,
		\miim1_BitCounter_reg[5]/NET0131 ,
		\miim1_BitCounter_reg[6]/NET0131 ,
		_w24565_
	);
	LUT2 #(
		.INIT('h8)
	) name14053 (
		_w24564_,
		_w24565_,
		_w24566_
	);
	LUT3 #(
		.INIT('h80)
	) name14054 (
		\miim1_InProgress_reg/NET0131 ,
		_w24564_,
		_w24565_,
		_w24567_
	);
	LUT4 #(
		.INIT('h0100)
	) name14055 (
		\miim1_BitCounter_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[1]/NET0131 ,
		\miim1_BitCounter_reg[2]/NET0131 ,
		\miim1_BitCounter_reg[5]/NET0131 ,
		_w24568_
	);
	LUT3 #(
		.INIT('h10)
	) name14056 (
		\miim1_BitCounter_reg[4]/NET0131 ,
		\miim1_BitCounter_reg[6]/NET0131 ,
		\miim1_InProgress_reg/NET0131 ,
		_w24569_
	);
	LUT2 #(
		.INIT('h1)
	) name14057 (
		\ethreg1_MIIMODER_1_DataOut_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24570_
	);
	LUT3 #(
		.INIT('h80)
	) name14058 (
		_w24568_,
		_w24569_,
		_w24570_,
		_w24571_
	);
	LUT4 #(
		.INIT('h0200)
	) name14059 (
		\miim1_BitCounter_reg[3]/NET0131 ,
		\miim1_BitCounter_reg[4]/NET0131 ,
		\miim1_BitCounter_reg[6]/NET0131 ,
		\miim1_InProgress_reg/NET0131 ,
		_w24572_
	);
	LUT4 #(
		.INIT('h2000)
	) name14060 (
		\miim1_BitCounter_reg[4]/NET0131 ,
		\miim1_BitCounter_reg[6]/NET0131 ,
		\miim1_InProgress_reg/NET0131 ,
		\miim1_WriteOp_reg/NET0131 ,
		_w24573_
	);
	LUT3 #(
		.INIT('hac)
	) name14061 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_MIITX_DATA_1_DataOut_reg[1]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24574_
	);
	LUT4 #(
		.INIT('h5777)
	) name14062 (
		_w24568_,
		_w24572_,
		_w24573_,
		_w24574_,
		_w24575_
	);
	LUT4 #(
		.INIT('h5700)
	) name14063 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[2]/NET0131 ,
		_w24567_,
		_w24571_,
		_w24575_,
		_w24576_
	);
	LUT4 #(
		.INIT('h222a)
	) name14064 (
		\miim1_shftrg_ShiftReg_reg[0]/NET0131 ,
		_w24568_,
		_w24572_,
		_w24573_,
		_w24577_
	);
	LUT4 #(
		.INIT('h5455)
	) name14065 (
		_w24562_,
		_w24567_,
		_w24571_,
		_w24577_,
		_w24578_
	);
	LUT3 #(
		.INIT('h15)
	) name14066 (
		_w24563_,
		_w24576_,
		_w24578_,
		_w24579_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name14067 (
		mdc_pad_o_pad,
		\miim1_shftrg_ShiftReg_reg[2]/NET0131 ,
		_w24411_,
		_w24420_,
		_w24580_
	);
	LUT4 #(
		.INIT('h1333)
	) name14068 (
		mdc_pad_o_pad,
		\miim1_shftrg_ShiftReg_reg[2]/NET0131 ,
		_w24411_,
		_w24420_,
		_w24581_
	);
	LUT3 #(
		.INIT('ha8)
	) name14069 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[3]/NET0131 ,
		_w24567_,
		_w24571_,
		_w24582_
	);
	LUT2 #(
		.INIT('h2)
	) name14070 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[2]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24583_
	);
	LUT3 #(
		.INIT('h80)
	) name14071 (
		_w24568_,
		_w24573_,
		_w24583_,
		_w24584_
	);
	LUT2 #(
		.INIT('h8)
	) name14072 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[2]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24585_
	);
	LUT3 #(
		.INIT('h80)
	) name14073 (
		_w24568_,
		_w24573_,
		_w24585_,
		_w24586_
	);
	LUT3 #(
		.INIT('h80)
	) name14074 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[0]/NET0131 ,
		_w24568_,
		_w24572_,
		_w24587_
	);
	LUT3 #(
		.INIT('h01)
	) name14075 (
		_w24584_,
		_w24586_,
		_w24587_,
		_w24588_
	);
	LUT4 #(
		.INIT('h222a)
	) name14076 (
		\miim1_shftrg_ShiftReg_reg[1]/NET0131 ,
		_w24568_,
		_w24572_,
		_w24573_,
		_w24589_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name14077 (
		_w24567_,
		_w24571_,
		_w24580_,
		_w24589_,
		_w24590_
	);
	LUT4 #(
		.INIT('h4555)
	) name14078 (
		_w24581_,
		_w24582_,
		_w24588_,
		_w24590_,
		_w24591_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name14079 (
		mdc_pad_o_pad,
		\miim1_shftrg_ShiftReg_reg[3]/NET0131 ,
		_w24411_,
		_w24420_,
		_w24592_
	);
	LUT4 #(
		.INIT('h1333)
	) name14080 (
		mdc_pad_o_pad,
		\miim1_shftrg_ShiftReg_reg[3]/NET0131 ,
		_w24411_,
		_w24420_,
		_w24593_
	);
	LUT3 #(
		.INIT('ha8)
	) name14081 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[4]/NET0131 ,
		_w24567_,
		_w24571_,
		_w24594_
	);
	LUT2 #(
		.INIT('h2)
	) name14082 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[3]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24595_
	);
	LUT3 #(
		.INIT('h80)
	) name14083 (
		_w24568_,
		_w24573_,
		_w24595_,
		_w24596_
	);
	LUT2 #(
		.INIT('h8)
	) name14084 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[3]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24597_
	);
	LUT3 #(
		.INIT('h80)
	) name14085 (
		_w24568_,
		_w24573_,
		_w24597_,
		_w24598_
	);
	LUT3 #(
		.INIT('h80)
	) name14086 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[1]/NET0131 ,
		_w24568_,
		_w24572_,
		_w24599_
	);
	LUT3 #(
		.INIT('h01)
	) name14087 (
		_w24596_,
		_w24598_,
		_w24599_,
		_w24600_
	);
	LUT4 #(
		.INIT('h222a)
	) name14088 (
		\miim1_shftrg_ShiftReg_reg[2]/NET0131 ,
		_w24568_,
		_w24572_,
		_w24573_,
		_w24601_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name14089 (
		_w24567_,
		_w24571_,
		_w24592_,
		_w24601_,
		_w24602_
	);
	LUT4 #(
		.INIT('h4555)
	) name14090 (
		_w24593_,
		_w24594_,
		_w24600_,
		_w24602_,
		_w24603_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name14091 (
		mdc_pad_o_pad,
		\miim1_shftrg_ShiftReg_reg[4]/NET0131 ,
		_w24411_,
		_w24420_,
		_w24604_
	);
	LUT4 #(
		.INIT('h1333)
	) name14092 (
		mdc_pad_o_pad,
		\miim1_shftrg_ShiftReg_reg[4]/NET0131 ,
		_w24411_,
		_w24420_,
		_w24605_
	);
	LUT3 #(
		.INIT('ha8)
	) name14093 (
		\miim1_WriteOp_reg/NET0131 ,
		_w24567_,
		_w24571_,
		_w24606_
	);
	LUT2 #(
		.INIT('h2)
	) name14094 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[4]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24607_
	);
	LUT3 #(
		.INIT('h80)
	) name14095 (
		_w24568_,
		_w24573_,
		_w24607_,
		_w24608_
	);
	LUT2 #(
		.INIT('h8)
	) name14096 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[4]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24609_
	);
	LUT3 #(
		.INIT('h80)
	) name14097 (
		_w24568_,
		_w24573_,
		_w24609_,
		_w24610_
	);
	LUT3 #(
		.INIT('h80)
	) name14098 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[2]/NET0131 ,
		_w24568_,
		_w24572_,
		_w24611_
	);
	LUT3 #(
		.INIT('h01)
	) name14099 (
		_w24608_,
		_w24610_,
		_w24611_,
		_w24612_
	);
	LUT4 #(
		.INIT('h222a)
	) name14100 (
		\miim1_shftrg_ShiftReg_reg[3]/NET0131 ,
		_w24568_,
		_w24572_,
		_w24573_,
		_w24613_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name14101 (
		_w24567_,
		_w24571_,
		_w24604_,
		_w24613_,
		_w24614_
	);
	LUT4 #(
		.INIT('h4555)
	) name14102 (
		_w24605_,
		_w24606_,
		_w24612_,
		_w24614_,
		_w24615_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name14103 (
		mdc_pad_o_pad,
		\miim1_shftrg_ShiftReg_reg[5]/NET0131 ,
		_w24411_,
		_w24420_,
		_w24616_
	);
	LUT4 #(
		.INIT('h1333)
	) name14104 (
		mdc_pad_o_pad,
		\miim1_shftrg_ShiftReg_reg[5]/NET0131 ,
		_w24411_,
		_w24420_,
		_w24617_
	);
	LUT3 #(
		.INIT('h54)
	) name14105 (
		\miim1_WriteOp_reg/NET0131 ,
		_w24567_,
		_w24571_,
		_w24618_
	);
	LUT2 #(
		.INIT('h2)
	) name14106 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[5]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24619_
	);
	LUT3 #(
		.INIT('h80)
	) name14107 (
		_w24568_,
		_w24573_,
		_w24619_,
		_w24620_
	);
	LUT2 #(
		.INIT('h8)
	) name14108 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[5]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24621_
	);
	LUT3 #(
		.INIT('h80)
	) name14109 (
		_w24568_,
		_w24573_,
		_w24621_,
		_w24622_
	);
	LUT3 #(
		.INIT('h80)
	) name14110 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[3]/NET0131 ,
		_w24568_,
		_w24572_,
		_w24623_
	);
	LUT3 #(
		.INIT('h01)
	) name14111 (
		_w24620_,
		_w24622_,
		_w24623_,
		_w24624_
	);
	LUT4 #(
		.INIT('h222a)
	) name14112 (
		\miim1_shftrg_ShiftReg_reg[4]/NET0131 ,
		_w24568_,
		_w24572_,
		_w24573_,
		_w24625_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name14113 (
		_w24567_,
		_w24571_,
		_w24616_,
		_w24625_,
		_w24626_
	);
	LUT4 #(
		.INIT('h4555)
	) name14114 (
		_w24617_,
		_w24618_,
		_w24624_,
		_w24626_,
		_w24627_
	);
	LUT3 #(
		.INIT('h80)
	) name14115 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[4]/NET0131 ,
		_w24568_,
		_w24572_,
		_w24628_
	);
	LUT2 #(
		.INIT('h2)
	) name14116 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[6]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24629_
	);
	LUT3 #(
		.INIT('h80)
	) name14117 (
		_w24568_,
		_w24573_,
		_w24629_,
		_w24630_
	);
	LUT4 #(
		.INIT('h0001)
	) name14118 (
		_w24567_,
		_w24571_,
		_w24628_,
		_w24630_,
		_w24631_
	);
	LUT4 #(
		.INIT('h222a)
	) name14119 (
		\miim1_shftrg_ShiftReg_reg[5]/NET0131 ,
		_w24568_,
		_w24572_,
		_w24573_,
		_w24632_
	);
	LUT2 #(
		.INIT('h8)
	) name14120 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[6]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24633_
	);
	LUT3 #(
		.INIT('h80)
	) name14121 (
		_w24568_,
		_w24573_,
		_w24633_,
		_w24634_
	);
	LUT2 #(
		.INIT('h1)
	) name14122 (
		_w24632_,
		_w24634_,
		_w24635_
	);
	LUT4 #(
		.INIT('h2eee)
	) name14123 (
		\miim1_shftrg_ShiftReg_reg[6]/NET0131 ,
		_w24561_,
		_w24631_,
		_w24635_,
		_w24636_
	);
	LUT3 #(
		.INIT('h10)
	) name14124 (
		\txethmac1_TxAbort_reg/NET0131 ,
		_w11065_,
		_w11068_,
		_w24637_
	);
	LUT3 #(
		.INIT('h07)
	) name14125 (
		_w10834_,
		_w10975_,
		_w11075_,
		_w24638_
	);
	LUT3 #(
		.INIT('h07)
	) name14126 (
		_w11062_,
		_w24637_,
		_w24638_,
		_w24639_
	);
	LUT2 #(
		.INIT('h4)
	) name14127 (
		\ethreg1_RXHASH1_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24640_
	);
	LUT4 #(
		.INIT('h0c08)
	) name14128 (
		\ethreg1_RXHASH0_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24641_
	);
	LUT3 #(
		.INIT('h45)
	) name14129 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w24640_,
		_w24641_,
		_w24642_
	);
	LUT2 #(
		.INIT('h4)
	) name14130 (
		\ethreg1_RXHASH1_0_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24643_
	);
	LUT4 #(
		.INIT('h0302)
	) name14131 (
		\ethreg1_RXHASH0_0_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24644_
	);
	LUT2 #(
		.INIT('h4)
	) name14132 (
		_w24643_,
		_w24644_,
		_w24645_
	);
	LUT2 #(
		.INIT('h4)
	) name14133 (
		\ethreg1_RXHASH1_3_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24646_
	);
	LUT4 #(
		.INIT('hc080)
	) name14134 (
		\ethreg1_RXHASH0_3_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24647_
	);
	LUT2 #(
		.INIT('h4)
	) name14135 (
		\ethreg1_RXHASH1_2_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24648_
	);
	LUT4 #(
		.INIT('h3020)
	) name14136 (
		\ethreg1_RXHASH0_2_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24649_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14137 (
		_w24646_,
		_w24647_,
		_w24648_,
		_w24649_,
		_w24650_
	);
	LUT3 #(
		.INIT('h20)
	) name14138 (
		_w24642_,
		_w24645_,
		_w24650_,
		_w24651_
	);
	LUT2 #(
		.INIT('h4)
	) name14139 (
		\ethreg1_RXHASH1_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24652_
	);
	LUT4 #(
		.INIT('h0c08)
	) name14140 (
		\ethreg1_RXHASH0_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24653_
	);
	LUT3 #(
		.INIT('h8a)
	) name14141 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w24652_,
		_w24653_,
		_w24654_
	);
	LUT2 #(
		.INIT('h4)
	) name14142 (
		\ethreg1_RXHASH1_0_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24655_
	);
	LUT4 #(
		.INIT('h0302)
	) name14143 (
		\ethreg1_RXHASH0_0_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24656_
	);
	LUT2 #(
		.INIT('h4)
	) name14144 (
		_w24655_,
		_w24656_,
		_w24657_
	);
	LUT2 #(
		.INIT('h4)
	) name14145 (
		\ethreg1_RXHASH1_2_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24658_
	);
	LUT4 #(
		.INIT('h3020)
	) name14146 (
		\ethreg1_RXHASH0_2_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24659_
	);
	LUT2 #(
		.INIT('h4)
	) name14147 (
		\ethreg1_RXHASH1_3_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24660_
	);
	LUT4 #(
		.INIT('hc080)
	) name14148 (
		\ethreg1_RXHASH0_3_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24661_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14149 (
		_w24658_,
		_w24659_,
		_w24660_,
		_w24661_,
		_w24662_
	);
	LUT3 #(
		.INIT('h20)
	) name14150 (
		_w24654_,
		_w24657_,
		_w24662_,
		_w24663_
	);
	LUT2 #(
		.INIT('h2)
	) name14151 (
		\rxethmac1_CrcHash_reg[1]/P0001 ,
		\rxethmac1_CrcHash_reg[2]/P0001 ,
		_w24664_
	);
	LUT3 #(
		.INIT('h10)
	) name14152 (
		_w24651_,
		_w24663_,
		_w24664_,
		_w24665_
	);
	LUT2 #(
		.INIT('h4)
	) name14153 (
		\ethreg1_RXHASH1_0_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24666_
	);
	LUT4 #(
		.INIT('h0302)
	) name14154 (
		\ethreg1_RXHASH0_0_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24667_
	);
	LUT3 #(
		.INIT('h8a)
	) name14155 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w24666_,
		_w24667_,
		_w24668_
	);
	LUT2 #(
		.INIT('h4)
	) name14156 (
		\ethreg1_RXHASH1_2_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24669_
	);
	LUT4 #(
		.INIT('h3020)
	) name14157 (
		\ethreg1_RXHASH0_2_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24670_
	);
	LUT2 #(
		.INIT('h4)
	) name14158 (
		_w24669_,
		_w24670_,
		_w24671_
	);
	LUT2 #(
		.INIT('h4)
	) name14159 (
		\ethreg1_RXHASH1_1_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24672_
	);
	LUT4 #(
		.INIT('h0c08)
	) name14160 (
		\ethreg1_RXHASH0_1_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24673_
	);
	LUT2 #(
		.INIT('h4)
	) name14161 (
		\ethreg1_RXHASH1_3_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24674_
	);
	LUT4 #(
		.INIT('hc080)
	) name14162 (
		\ethreg1_RXHASH0_3_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24675_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14163 (
		_w24672_,
		_w24673_,
		_w24674_,
		_w24675_,
		_w24676_
	);
	LUT3 #(
		.INIT('h20)
	) name14164 (
		_w24668_,
		_w24671_,
		_w24676_,
		_w24677_
	);
	LUT2 #(
		.INIT('h4)
	) name14165 (
		\ethreg1_RXHASH1_3_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24678_
	);
	LUT4 #(
		.INIT('hc080)
	) name14166 (
		\ethreg1_RXHASH0_3_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24679_
	);
	LUT3 #(
		.INIT('h45)
	) name14167 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w24678_,
		_w24679_,
		_w24680_
	);
	LUT2 #(
		.INIT('h4)
	) name14168 (
		\ethreg1_RXHASH1_0_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24681_
	);
	LUT4 #(
		.INIT('h0302)
	) name14169 (
		\ethreg1_RXHASH0_0_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24682_
	);
	LUT2 #(
		.INIT('h4)
	) name14170 (
		_w24681_,
		_w24682_,
		_w24683_
	);
	LUT2 #(
		.INIT('h4)
	) name14171 (
		\ethreg1_RXHASH1_2_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24684_
	);
	LUT4 #(
		.INIT('h3020)
	) name14172 (
		\ethreg1_RXHASH0_2_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24685_
	);
	LUT2 #(
		.INIT('h4)
	) name14173 (
		\ethreg1_RXHASH1_1_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24686_
	);
	LUT4 #(
		.INIT('h0c08)
	) name14174 (
		\ethreg1_RXHASH0_1_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24687_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14175 (
		_w24684_,
		_w24685_,
		_w24686_,
		_w24687_,
		_w24688_
	);
	LUT3 #(
		.INIT('h20)
	) name14176 (
		_w24680_,
		_w24683_,
		_w24688_,
		_w24689_
	);
	LUT2 #(
		.INIT('h1)
	) name14177 (
		\rxethmac1_CrcHash_reg[1]/P0001 ,
		\rxethmac1_CrcHash_reg[2]/P0001 ,
		_w24690_
	);
	LUT3 #(
		.INIT('h10)
	) name14178 (
		_w24677_,
		_w24689_,
		_w24690_,
		_w24691_
	);
	LUT2 #(
		.INIT('h1)
	) name14179 (
		_w24665_,
		_w24691_,
		_w24692_
	);
	LUT2 #(
		.INIT('h8)
	) name14180 (
		\rxethmac1_CrcHashGood_reg/P0001 ,
		\rxethmac1_Multicast_reg/NET0131 ,
		_w24693_
	);
	LUT2 #(
		.INIT('h4)
	) name14181 (
		\ethreg1_RXHASH1_0_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24694_
	);
	LUT4 #(
		.INIT('h0302)
	) name14182 (
		\ethreg1_RXHASH0_0_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24695_
	);
	LUT3 #(
		.INIT('h45)
	) name14183 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w24694_,
		_w24695_,
		_w24696_
	);
	LUT2 #(
		.INIT('h4)
	) name14184 (
		\ethreg1_RXHASH1_3_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24697_
	);
	LUT4 #(
		.INIT('hc080)
	) name14185 (
		\ethreg1_RXHASH0_3_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24698_
	);
	LUT2 #(
		.INIT('h4)
	) name14186 (
		_w24697_,
		_w24698_,
		_w24699_
	);
	LUT2 #(
		.INIT('h4)
	) name14187 (
		\ethreg1_RXHASH1_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24700_
	);
	LUT4 #(
		.INIT('h0c08)
	) name14188 (
		\ethreg1_RXHASH0_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24701_
	);
	LUT2 #(
		.INIT('h4)
	) name14189 (
		\ethreg1_RXHASH1_2_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24702_
	);
	LUT4 #(
		.INIT('h3020)
	) name14190 (
		\ethreg1_RXHASH0_2_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24703_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14191 (
		_w24700_,
		_w24701_,
		_w24702_,
		_w24703_,
		_w24704_
	);
	LUT3 #(
		.INIT('h20)
	) name14192 (
		_w24696_,
		_w24699_,
		_w24704_,
		_w24705_
	);
	LUT2 #(
		.INIT('h4)
	) name14193 (
		\ethreg1_RXHASH1_0_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24706_
	);
	LUT4 #(
		.INIT('h0302)
	) name14194 (
		\ethreg1_RXHASH0_0_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24707_
	);
	LUT3 #(
		.INIT('h8a)
	) name14195 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w24706_,
		_w24707_,
		_w24708_
	);
	LUT2 #(
		.INIT('h4)
	) name14196 (
		\ethreg1_RXHASH1_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24709_
	);
	LUT4 #(
		.INIT('h0c08)
	) name14197 (
		\ethreg1_RXHASH0_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24710_
	);
	LUT2 #(
		.INIT('h4)
	) name14198 (
		_w24709_,
		_w24710_,
		_w24711_
	);
	LUT2 #(
		.INIT('h4)
	) name14199 (
		\ethreg1_RXHASH1_2_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24712_
	);
	LUT4 #(
		.INIT('h3020)
	) name14200 (
		\ethreg1_RXHASH0_2_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24713_
	);
	LUT2 #(
		.INIT('h4)
	) name14201 (
		\ethreg1_RXHASH1_3_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24714_
	);
	LUT4 #(
		.INIT('hc080)
	) name14202 (
		\ethreg1_RXHASH0_3_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24715_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14203 (
		_w24712_,
		_w24713_,
		_w24714_,
		_w24715_,
		_w24716_
	);
	LUT3 #(
		.INIT('h20)
	) name14204 (
		_w24708_,
		_w24711_,
		_w24716_,
		_w24717_
	);
	LUT2 #(
		.INIT('h8)
	) name14205 (
		\rxethmac1_CrcHash_reg[1]/P0001 ,
		\rxethmac1_CrcHash_reg[2]/P0001 ,
		_w24718_
	);
	LUT3 #(
		.INIT('h10)
	) name14206 (
		_w24705_,
		_w24717_,
		_w24718_,
		_w24719_
	);
	LUT2 #(
		.INIT('h4)
	) name14207 (
		\ethreg1_RXHASH1_3_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24720_
	);
	LUT4 #(
		.INIT('hc080)
	) name14208 (
		\ethreg1_RXHASH0_3_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24721_
	);
	LUT3 #(
		.INIT('h8a)
	) name14209 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w24720_,
		_w24721_,
		_w24722_
	);
	LUT2 #(
		.INIT('h4)
	) name14210 (
		\ethreg1_RXHASH1_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24723_
	);
	LUT4 #(
		.INIT('h0c08)
	) name14211 (
		\ethreg1_RXHASH0_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24724_
	);
	LUT2 #(
		.INIT('h4)
	) name14212 (
		_w24723_,
		_w24724_,
		_w24725_
	);
	LUT2 #(
		.INIT('h4)
	) name14213 (
		\ethreg1_RXHASH1_2_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24726_
	);
	LUT4 #(
		.INIT('h3020)
	) name14214 (
		\ethreg1_RXHASH0_2_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24727_
	);
	LUT2 #(
		.INIT('h4)
	) name14215 (
		\ethreg1_RXHASH1_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24728_
	);
	LUT4 #(
		.INIT('h0302)
	) name14216 (
		\ethreg1_RXHASH0_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24729_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14217 (
		_w24726_,
		_w24727_,
		_w24728_,
		_w24729_,
		_w24730_
	);
	LUT3 #(
		.INIT('h20)
	) name14218 (
		_w24722_,
		_w24725_,
		_w24730_,
		_w24731_
	);
	LUT2 #(
		.INIT('h4)
	) name14219 (
		\ethreg1_RXHASH1_0_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24732_
	);
	LUT4 #(
		.INIT('h0302)
	) name14220 (
		\ethreg1_RXHASH0_0_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24733_
	);
	LUT3 #(
		.INIT('h45)
	) name14221 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w24732_,
		_w24733_,
		_w24734_
	);
	LUT2 #(
		.INIT('h4)
	) name14222 (
		\ethreg1_RXHASH1_3_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24735_
	);
	LUT4 #(
		.INIT('hc080)
	) name14223 (
		\ethreg1_RXHASH0_3_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24736_
	);
	LUT2 #(
		.INIT('h4)
	) name14224 (
		_w24735_,
		_w24736_,
		_w24737_
	);
	LUT2 #(
		.INIT('h4)
	) name14225 (
		\ethreg1_RXHASH1_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24738_
	);
	LUT4 #(
		.INIT('h0c08)
	) name14226 (
		\ethreg1_RXHASH0_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24739_
	);
	LUT2 #(
		.INIT('h4)
	) name14227 (
		\ethreg1_RXHASH1_2_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24740_
	);
	LUT4 #(
		.INIT('h3020)
	) name14228 (
		\ethreg1_RXHASH0_2_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w24741_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14229 (
		_w24738_,
		_w24739_,
		_w24740_,
		_w24741_,
		_w24742_
	);
	LUT3 #(
		.INIT('h20)
	) name14230 (
		_w24734_,
		_w24737_,
		_w24742_,
		_w24743_
	);
	LUT2 #(
		.INIT('h4)
	) name14231 (
		\rxethmac1_CrcHash_reg[1]/P0001 ,
		\rxethmac1_CrcHash_reg[2]/P0001 ,
		_w24744_
	);
	LUT3 #(
		.INIT('h10)
	) name14232 (
		_w24731_,
		_w24743_,
		_w24744_,
		_w24745_
	);
	LUT3 #(
		.INIT('h02)
	) name14233 (
		_w24693_,
		_w24719_,
		_w24745_,
		_w24746_
	);
	LUT3 #(
		.INIT('h07)
	) name14234 (
		\rxethmac1_CrcHashGood_reg/P0001 ,
		\rxethmac1_Multicast_reg/NET0131 ,
		\rxethmac1_rxaddrcheck1_MulticastOK_reg/NET0131 ,
		_w24747_
	);
	LUT2 #(
		.INIT('h2)
	) name14235 (
		_w11795_,
		_w24747_,
		_w24748_
	);
	LUT3 #(
		.INIT('h70)
	) name14236 (
		_w24692_,
		_w24746_,
		_w24748_,
		_w24749_
	);
	LUT4 #(
		.INIT('h4000)
	) name14237 (
		\wb_adr_i[11]_pad ,
		wb_cyc_i_pad,
		\wb_sel_i[0]_pad ,
		wb_stb_i_pad,
		_w24750_
	);
	LUT2 #(
		.INIT('h4)
	) name14238 (
		_w18750_,
		_w24750_,
		_w24751_
	);
	LUT2 #(
		.INIT('h4)
	) name14239 (
		\wb_adr_i[10]_pad ,
		wb_we_i_pad,
		_w24752_
	);
	LUT3 #(
		.INIT('h40)
	) name14240 (
		_w18750_,
		_w24750_,
		_w24752_,
		_w24753_
	);
	LUT2 #(
		.INIT('h4)
	) name14241 (
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w24754_
	);
	LUT4 #(
		.INIT('h0001)
	) name14242 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[6]_pad ,
		\wb_dat_i[10]_pad ,
		_w24755_
	);
	LUT2 #(
		.INIT('h8)
	) name14243 (
		_w24754_,
		_w24755_,
		_w24756_
	);
	LUT4 #(
		.INIT('h0001)
	) name14244 (
		\wb_dat_i[15]_pad ,
		\wb_dat_i[16]_pad ,
		\wb_dat_i[17]_pad ,
		\wb_dat_i[18]_pad ,
		_w24757_
	);
	LUT4 #(
		.INIT('h0001)
	) name14245 (
		\wb_dat_i[11]_pad ,
		\wb_dat_i[12]_pad ,
		\wb_dat_i[13]_pad ,
		\wb_dat_i[14]_pad ,
		_w24758_
	);
	LUT4 #(
		.INIT('h0001)
	) name14246 (
		\wb_dat_i[23]_pad ,
		\wb_dat_i[24]_pad ,
		\wb_dat_i[25]_pad ,
		\wb_dat_i[26]_pad ,
		_w24759_
	);
	LUT4 #(
		.INIT('h0001)
	) name14247 (
		\wb_dat_i[19]_pad ,
		\wb_dat_i[20]_pad ,
		\wb_dat_i[21]_pad ,
		\wb_dat_i[22]_pad ,
		_w24760_
	);
	LUT4 #(
		.INIT('h8000)
	) name14248 (
		_w24757_,
		_w24758_,
		_w24759_,
		_w24760_,
		_w24761_
	);
	LUT3 #(
		.INIT('h01)
	) name14249 (
		\wb_dat_i[4]_pad ,
		\wb_dat_i[5]_pad ,
		\wb_dat_i[6]_pad ,
		_w24762_
	);
	LUT4 #(
		.INIT('h0001)
	) name14250 (
		\wb_dat_i[0]_pad ,
		\wb_dat_i[1]_pad ,
		\wb_dat_i[2]_pad ,
		\wb_dat_i[3]_pad ,
		_w24763_
	);
	LUT3 #(
		.INIT('h2a)
	) name14251 (
		\wb_dat_i[7]_pad ,
		_w24762_,
		_w24763_,
		_w24764_
	);
	LUT3 #(
		.INIT('h01)
	) name14252 (
		\wb_adr_i[7]_pad ,
		\wb_adr_i[8]_pad ,
		\wb_adr_i[9]_pad ,
		_w24765_
	);
	LUT3 #(
		.INIT('h01)
	) name14253 (
		\wb_dat_i[31]_pad ,
		\wb_dat_i[8]_pad ,
		\wb_dat_i[9]_pad ,
		_w24766_
	);
	LUT4 #(
		.INIT('h0001)
	) name14254 (
		\wb_dat_i[27]_pad ,
		\wb_dat_i[28]_pad ,
		\wb_dat_i[29]_pad ,
		\wb_dat_i[30]_pad ,
		_w24767_
	);
	LUT3 #(
		.INIT('h80)
	) name14255 (
		_w24765_,
		_w24766_,
		_w24767_,
		_w24768_
	);
	LUT4 #(
		.INIT('h0800)
	) name14256 (
		_w24756_,
		_w24761_,
		_w24764_,
		_w24768_,
		_w24769_
	);
	LUT2 #(
		.INIT('h8)
	) name14257 (
		_w24753_,
		_w24769_,
		_w24770_
	);
	LUT2 #(
		.INIT('h1)
	) name14258 (
		\rxethmac1_crcrx_Crc_reg[17]/NET0131 ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w24771_
	);
	LUT4 #(
		.INIT('h02ff)
	) name14259 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		_w10542_,
		_w10543_,
		_w24771_,
		_w24772_
	);
	LUT3 #(
		.INIT('h14)
	) name14260 (
		\rxethmac1_crcrx_Crc_reg[2]/NET0131 ,
		_w10580_,
		_w10590_,
		_w24773_
	);
	LUT4 #(
		.INIT('h7000)
	) name14261 (
		_w10554_,
		_w10573_,
		_w10577_,
		_w24773_,
		_w24774_
	);
	LUT2 #(
		.INIT('h4)
	) name14262 (
		\rxethmac1_crcrx_Crc_reg[2]/NET0131 ,
		_w10582_,
		_w24775_
	);
	LUT3 #(
		.INIT('hab)
	) name14263 (
		_w24774_,
		_w24775_,
		_w10958_,
		_w24776_
	);
	LUT2 #(
		.INIT('h2)
	) name14264 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24777_
	);
	LUT4 #(
		.INIT('h1000)
	) name14265 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_OpCodeOK_reg/NET0131 ,
		\maccontrol1_receivecontrol1_TypeLengthOK_reg/NET0131 ,
		_w24778_
	);
	LUT2 #(
		.INIT('h2)
	) name14266 (
		\maccontrol1_receivecontrol1_AddressOK_reg/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24779_
	);
	LUT4 #(
		.INIT('heccc)
	) name14267 (
		_w11921_,
		_w24777_,
		_w24778_,
		_w24779_,
		_w24780_
	);
	LUT4 #(
		.INIT('h1000)
	) name14268 (
		\txethmac1_txcrc_Crc_reg[0]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11776_,
		_w11779_,
		_w24781_
	);
	LUT3 #(
		.INIT('h40)
	) name14269 (
		\txethmac1_txcrc_Crc_reg[0]/NET0131 ,
		_w10913_,
		_w10914_,
		_w24782_
	);
	LUT3 #(
		.INIT('hcd)
	) name14270 (
		_w11782_,
		_w24781_,
		_w24782_,
		_w24783_
	);
	LUT4 #(
		.INIT('h2000)
	) name14271 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w24784_
	);
	LUT2 #(
		.INIT('h2)
	) name14272 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[0]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24785_
	);
	LUT2 #(
		.INIT('h2)
	) name14273 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24786_
	);
	LUT4 #(
		.INIT('hf870)
	) name14274 (
		_w24444_,
		_w24784_,
		_w24785_,
		_w24786_,
		_w24787_
	);
	LUT4 #(
		.INIT('h1000)
	) name14275 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w24788_
	);
	LUT2 #(
		.INIT('h2)
	) name14276 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[10]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24789_
	);
	LUT2 #(
		.INIT('h2)
	) name14277 (
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24790_
	);
	LUT4 #(
		.INIT('hf870)
	) name14278 (
		_w24444_,
		_w24788_,
		_w24789_,
		_w24790_,
		_w24791_
	);
	LUT2 #(
		.INIT('h2)
	) name14279 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[11]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24792_
	);
	LUT2 #(
		.INIT('h2)
	) name14280 (
		\rxethmac1_RxData_reg[3]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24793_
	);
	LUT4 #(
		.INIT('hf870)
	) name14281 (
		_w24444_,
		_w24788_,
		_w24792_,
		_w24793_,
		_w24794_
	);
	LUT2 #(
		.INIT('h2)
	) name14282 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[12]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24795_
	);
	LUT2 #(
		.INIT('h2)
	) name14283 (
		\rxethmac1_RxData_reg[4]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24796_
	);
	LUT4 #(
		.INIT('hf870)
	) name14284 (
		_w24444_,
		_w24788_,
		_w24795_,
		_w24796_,
		_w24797_
	);
	LUT2 #(
		.INIT('h2)
	) name14285 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[13]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24798_
	);
	LUT2 #(
		.INIT('h2)
	) name14286 (
		\rxethmac1_RxData_reg[5]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24799_
	);
	LUT4 #(
		.INIT('hf870)
	) name14287 (
		_w24444_,
		_w24788_,
		_w24798_,
		_w24799_,
		_w24800_
	);
	LUT2 #(
		.INIT('h2)
	) name14288 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[14]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24801_
	);
	LUT2 #(
		.INIT('h2)
	) name14289 (
		\rxethmac1_RxData_reg[6]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24802_
	);
	LUT4 #(
		.INIT('hf870)
	) name14290 (
		_w24444_,
		_w24788_,
		_w24801_,
		_w24802_,
		_w24803_
	);
	LUT2 #(
		.INIT('h2)
	) name14291 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[15]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24804_
	);
	LUT2 #(
		.INIT('h2)
	) name14292 (
		\rxethmac1_RxData_reg[7]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24805_
	);
	LUT4 #(
		.INIT('hf870)
	) name14293 (
		_w24444_,
		_w24788_,
		_w24804_,
		_w24805_,
		_w24806_
	);
	LUT2 #(
		.INIT('h2)
	) name14294 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[1]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24807_
	);
	LUT2 #(
		.INIT('h2)
	) name14295 (
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24808_
	);
	LUT4 #(
		.INIT('hf870)
	) name14296 (
		_w24444_,
		_w24784_,
		_w24807_,
		_w24808_,
		_w24809_
	);
	LUT2 #(
		.INIT('h2)
	) name14297 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[2]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24810_
	);
	LUT4 #(
		.INIT('hf780)
	) name14298 (
		_w24444_,
		_w24784_,
		_w24790_,
		_w24810_,
		_w24811_
	);
	LUT2 #(
		.INIT('h2)
	) name14299 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[3]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24812_
	);
	LUT4 #(
		.INIT('hf780)
	) name14300 (
		_w24444_,
		_w24784_,
		_w24793_,
		_w24812_,
		_w24813_
	);
	LUT2 #(
		.INIT('h2)
	) name14301 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[4]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24814_
	);
	LUT4 #(
		.INIT('hf780)
	) name14302 (
		_w24444_,
		_w24784_,
		_w24796_,
		_w24814_,
		_w24815_
	);
	LUT2 #(
		.INIT('h2)
	) name14303 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[5]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24816_
	);
	LUT4 #(
		.INIT('hf780)
	) name14304 (
		_w24444_,
		_w24784_,
		_w24799_,
		_w24816_,
		_w24817_
	);
	LUT2 #(
		.INIT('h2)
	) name14305 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[6]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24818_
	);
	LUT4 #(
		.INIT('hf780)
	) name14306 (
		_w24444_,
		_w24784_,
		_w24802_,
		_w24818_,
		_w24819_
	);
	LUT2 #(
		.INIT('h2)
	) name14307 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[7]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24820_
	);
	LUT4 #(
		.INIT('hf780)
	) name14308 (
		_w24444_,
		_w24784_,
		_w24805_,
		_w24820_,
		_w24821_
	);
	LUT2 #(
		.INIT('h2)
	) name14309 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[8]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24822_
	);
	LUT4 #(
		.INIT('hdf80)
	) name14310 (
		_w24444_,
		_w24786_,
		_w24788_,
		_w24822_,
		_w24823_
	);
	LUT2 #(
		.INIT('h2)
	) name14311 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[9]/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w24824_
	);
	LUT4 #(
		.INIT('hf780)
	) name14312 (
		_w24444_,
		_w24788_,
		_w24808_,
		_w24824_,
		_w24825_
	);
	LUT3 #(
		.INIT('h2a)
	) name14313 (
		\m_wb_sel_o[1]_pad ,
		_w24509_,
		_w24515_,
		_w24826_
	);
	LUT2 #(
		.INIT('h8)
	) name14314 (
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w24827_
	);
	LUT3 #(
		.INIT('h40)
	) name14315 (
		_w11890_,
		_w11900_,
		_w24827_,
		_w24828_
	);
	LUT3 #(
		.INIT('hab)
	) name14316 (
		_w24826_,
		_w11907_,
		_w24828_,
		_w24829_
	);
	LUT3 #(
		.INIT('h54)
	) name14317 (
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w11902_,
		_w11905_,
		_w24830_
	);
	LUT3 #(
		.INIT('h2a)
	) name14318 (
		\m_wb_sel_o[2]_pad ,
		_w24509_,
		_w24515_,
		_w24831_
	);
	LUT3 #(
		.INIT('hfd)
	) name14319 (
		_w11901_,
		_w24830_,
		_w24831_,
		_w24832_
	);
	LUT3 #(
		.INIT('h2a)
	) name14320 (
		\m_wb_sel_o[3]_pad ,
		_w24509_,
		_w24515_,
		_w24833_
	);
	LUT2 #(
		.INIT('h1)
	) name14321 (
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w24834_
	);
	LUT3 #(
		.INIT('he0)
	) name14322 (
		_w11902_,
		_w11905_,
		_w24834_,
		_w24835_
	);
	LUT3 #(
		.INIT('hfd)
	) name14323 (
		_w11901_,
		_w24833_,
		_w24835_,
		_w24836_
	);
	LUT3 #(
		.INIT('h0b)
	) name14324 (
		_w24505_,
		_w24506_,
		_w24508_,
		_w24837_
	);
	LUT3 #(
		.INIT('h8a)
	) name14325 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		_w24514_,
		_w24837_,
		_w24838_
	);
	LUT2 #(
		.INIT('hd)
	) name14326 (
		_w11906_,
		_w24838_,
		_w24839_
	);
	LUT3 #(
		.INIT('h8a)
	) name14327 (
		\wishbone_MasterWbTX_reg/NET0131 ,
		_w24514_,
		_w24837_,
		_w24840_
	);
	LUT2 #(
		.INIT('hd)
	) name14328 (
		_w11901_,
		_w24840_,
		_w24841_
	);
	LUT2 #(
		.INIT('h1)
	) name14329 (
		\macstatus1_RxColWindow_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		_w24842_
	);
	LUT4 #(
		.INIT('h956a)
	) name14330 (
		\ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w24843_
	);
	LUT3 #(
		.INIT('h96)
	) name14331 (
		\ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		_w24844_
	);
	LUT2 #(
		.INIT('h6)
	) name14332 (
		\ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		_w24845_
	);
	LUT4 #(
		.INIT('h2100)
	) name14333 (
		\ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131 ,
		mcoll_pad_i_pad,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		_w24846_
	);
	LUT4 #(
		.INIT('h0100)
	) name14334 (
		_w24843_,
		_w24844_,
		_w24845_,
		_w24846_,
		_w24847_
	);
	LUT3 #(
		.INIT('h96)
	) name14335 (
		\ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w11135_,
		_w24848_
	);
	LUT4 #(
		.INIT('h69a5)
	) name14336 (
		\ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		_w11134_,
		_w24849_
	);
	LUT4 #(
		.INIT('h5155)
	) name14337 (
		_w24842_,
		_w24847_,
		_w24848_,
		_w24849_,
		_w24850_
	);
	LUT4 #(
		.INIT('h0007)
	) name14338 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131 ,
		_w24851_
	);
	LUT2 #(
		.INIT('h8)
	) name14339 (
		_w10514_,
		_w24851_,
		_w24852_
	);
	LUT3 #(
		.INIT('h2a)
	) name14340 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10519_,
		_w24852_,
		_w24853_
	);
	LUT2 #(
		.INIT('h8)
	) name14341 (
		\rxethmac1_DelayData_reg/NET0131 ,
		\rxethmac1_RxData_d_reg[0]/NET0131 ,
		_w24854_
	);
	LUT4 #(
		.INIT('hd500)
	) name14342 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10519_,
		_w24852_,
		_w24854_,
		_w24855_
	);
	LUT2 #(
		.INIT('h8)
	) name14343 (
		\rxethmac1_LatchedByte_reg[0]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w24856_
	);
	LUT3 #(
		.INIT('h70)
	) name14344 (
		_w10519_,
		_w24852_,
		_w24856_,
		_w24857_
	);
	LUT2 #(
		.INIT('he)
	) name14345 (
		_w24855_,
		_w24857_,
		_w24858_
	);
	LUT2 #(
		.INIT('h2)
	) name14346 (
		\txethmac1_StopExcessiveDeferOccured_reg/NET0131 ,
		_w10836_,
		_w24859_
	);
	LUT3 #(
		.INIT('hf8)
	) name14347 (
		_w10834_,
		_w10844_,
		_w24859_,
		_w24860_
	);
	LUT2 #(
		.INIT('h8)
	) name14348 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24861_
	);
	LUT3 #(
		.INIT('h80)
	) name14349 (
		_w24444_,
		_w24445_,
		_w24861_,
		_w24862_
	);
	LUT2 #(
		.INIT('h2)
	) name14350 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[0]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24863_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14351 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24863_,
		_w24864_
	);
	LUT2 #(
		.INIT('he)
	) name14352 (
		_w24862_,
		_w24864_,
		_w24865_
	);
	LUT2 #(
		.INIT('h8)
	) name14353 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[10]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24866_
	);
	LUT3 #(
		.INIT('h80)
	) name14354 (
		_w24444_,
		_w24445_,
		_w24866_,
		_w24867_
	);
	LUT2 #(
		.INIT('h2)
	) name14355 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[10]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24868_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14356 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24868_,
		_w24869_
	);
	LUT2 #(
		.INIT('he)
	) name14357 (
		_w24867_,
		_w24869_,
		_w24870_
	);
	LUT2 #(
		.INIT('h8)
	) name14358 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[11]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24871_
	);
	LUT3 #(
		.INIT('h80)
	) name14359 (
		_w24444_,
		_w24445_,
		_w24871_,
		_w24872_
	);
	LUT2 #(
		.INIT('h2)
	) name14360 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[11]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24873_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14361 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24873_,
		_w24874_
	);
	LUT2 #(
		.INIT('he)
	) name14362 (
		_w24872_,
		_w24874_,
		_w24875_
	);
	LUT2 #(
		.INIT('h8)
	) name14363 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[12]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24876_
	);
	LUT3 #(
		.INIT('h80)
	) name14364 (
		_w24444_,
		_w24445_,
		_w24876_,
		_w24877_
	);
	LUT2 #(
		.INIT('h2)
	) name14365 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[12]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24878_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14366 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24878_,
		_w24879_
	);
	LUT2 #(
		.INIT('he)
	) name14367 (
		_w24877_,
		_w24879_,
		_w24880_
	);
	LUT2 #(
		.INIT('h8)
	) name14368 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[13]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24881_
	);
	LUT3 #(
		.INIT('h80)
	) name14369 (
		_w24444_,
		_w24445_,
		_w24881_,
		_w24882_
	);
	LUT2 #(
		.INIT('h2)
	) name14370 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[13]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24883_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14371 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24883_,
		_w24884_
	);
	LUT2 #(
		.INIT('he)
	) name14372 (
		_w24882_,
		_w24884_,
		_w24885_
	);
	LUT2 #(
		.INIT('h8)
	) name14373 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[15]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24886_
	);
	LUT3 #(
		.INIT('h80)
	) name14374 (
		_w24444_,
		_w24445_,
		_w24886_,
		_w24887_
	);
	LUT2 #(
		.INIT('h2)
	) name14375 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[15]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24888_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14376 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24888_,
		_w24889_
	);
	LUT2 #(
		.INIT('he)
	) name14377 (
		_w24887_,
		_w24889_,
		_w24890_
	);
	LUT2 #(
		.INIT('h8)
	) name14378 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[14]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24891_
	);
	LUT3 #(
		.INIT('h80)
	) name14379 (
		_w24444_,
		_w24445_,
		_w24891_,
		_w24892_
	);
	LUT2 #(
		.INIT('h2)
	) name14380 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[14]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24893_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14381 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24893_,
		_w24894_
	);
	LUT2 #(
		.INIT('he)
	) name14382 (
		_w24892_,
		_w24894_,
		_w24895_
	);
	LUT2 #(
		.INIT('h8)
	) name14383 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24896_
	);
	LUT3 #(
		.INIT('h80)
	) name14384 (
		_w24444_,
		_w24445_,
		_w24896_,
		_w24897_
	);
	LUT2 #(
		.INIT('h2)
	) name14385 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[1]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24898_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14386 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24898_,
		_w24899_
	);
	LUT2 #(
		.INIT('he)
	) name14387 (
		_w24897_,
		_w24899_,
		_w24900_
	);
	LUT2 #(
		.INIT('h8)
	) name14388 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24901_
	);
	LUT3 #(
		.INIT('h80)
	) name14389 (
		_w24444_,
		_w24445_,
		_w24901_,
		_w24902_
	);
	LUT2 #(
		.INIT('h2)
	) name14390 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[2]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24903_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14391 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24903_,
		_w24904_
	);
	LUT2 #(
		.INIT('he)
	) name14392 (
		_w24902_,
		_w24904_,
		_w24905_
	);
	LUT2 #(
		.INIT('h8)
	) name14393 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[3]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24906_
	);
	LUT3 #(
		.INIT('h80)
	) name14394 (
		_w24444_,
		_w24445_,
		_w24906_,
		_w24907_
	);
	LUT2 #(
		.INIT('h2)
	) name14395 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[3]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24908_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14396 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24908_,
		_w24909_
	);
	LUT2 #(
		.INIT('he)
	) name14397 (
		_w24907_,
		_w24909_,
		_w24910_
	);
	LUT2 #(
		.INIT('h8)
	) name14398 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[4]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24911_
	);
	LUT3 #(
		.INIT('h80)
	) name14399 (
		_w24444_,
		_w24445_,
		_w24911_,
		_w24912_
	);
	LUT2 #(
		.INIT('h2)
	) name14400 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[4]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24913_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14401 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24913_,
		_w24914_
	);
	LUT2 #(
		.INIT('he)
	) name14402 (
		_w24912_,
		_w24914_,
		_w24915_
	);
	LUT2 #(
		.INIT('h8)
	) name14403 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[5]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24916_
	);
	LUT3 #(
		.INIT('h80)
	) name14404 (
		_w24444_,
		_w24445_,
		_w24916_,
		_w24917_
	);
	LUT2 #(
		.INIT('h2)
	) name14405 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[5]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24918_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14406 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24918_,
		_w24919_
	);
	LUT2 #(
		.INIT('he)
	) name14407 (
		_w24917_,
		_w24919_,
		_w24920_
	);
	LUT2 #(
		.INIT('h8)
	) name14408 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[6]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24921_
	);
	LUT3 #(
		.INIT('h80)
	) name14409 (
		_w24444_,
		_w24445_,
		_w24921_,
		_w24922_
	);
	LUT2 #(
		.INIT('h2)
	) name14410 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[6]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24923_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14411 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24923_,
		_w24924_
	);
	LUT2 #(
		.INIT('he)
	) name14412 (
		_w24922_,
		_w24924_,
		_w24925_
	);
	LUT2 #(
		.INIT('h8)
	) name14413 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[7]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24926_
	);
	LUT3 #(
		.INIT('h80)
	) name14414 (
		_w24444_,
		_w24445_,
		_w24926_,
		_w24927_
	);
	LUT2 #(
		.INIT('h2)
	) name14415 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[7]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24928_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14416 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24928_,
		_w24929_
	);
	LUT2 #(
		.INIT('he)
	) name14417 (
		_w24927_,
		_w24929_,
		_w24930_
	);
	LUT2 #(
		.INIT('h8)
	) name14418 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[8]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24931_
	);
	LUT3 #(
		.INIT('h80)
	) name14419 (
		_w24444_,
		_w24445_,
		_w24931_,
		_w24932_
	);
	LUT2 #(
		.INIT('h2)
	) name14420 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[8]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24933_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14421 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24933_,
		_w24934_
	);
	LUT2 #(
		.INIT('he)
	) name14422 (
		_w24932_,
		_w24934_,
		_w24935_
	);
	LUT2 #(
		.INIT('h8)
	) name14423 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[9]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24936_
	);
	LUT3 #(
		.INIT('h80)
	) name14424 (
		_w24444_,
		_w24445_,
		_w24936_,
		_w24937_
	);
	LUT2 #(
		.INIT('h2)
	) name14425 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[9]/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w24938_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14426 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w24444_,
		_w24445_,
		_w24938_,
		_w24939_
	);
	LUT2 #(
		.INIT('he)
	) name14427 (
		_w24937_,
		_w24939_,
		_w24940_
	);
	LUT4 #(
		.INIT('h0400)
	) name14428 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_LastByteIn_reg/NET0131 ,
		\wishbone_RxEnableWindow_reg/NET0131 ,
		_w24941_
	);
	LUT4 #(
		.INIT('h535c)
	) name14429 (
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		_w13419_,
		_w24941_,
		_w24942_
	);
	LUT4 #(
		.INIT('h060c)
	) name14430 (
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		_w13419_,
		_w24941_,
		_w24943_
	);
	LUT4 #(
		.INIT('h0880)
	) name14431 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w24944_
	);
	LUT2 #(
		.INIT('he)
	) name14432 (
		_w24943_,
		_w24944_,
		_w24945_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name14433 (
		mdc_pad_o_pad,
		\miim1_shftrg_ShiftReg_reg[0]/NET0131 ,
		_w24411_,
		_w24420_,
		_w24946_
	);
	LUT4 #(
		.INIT('h1333)
	) name14434 (
		mdc_pad_o_pad,
		\miim1_shftrg_ShiftReg_reg[0]/NET0131 ,
		_w24411_,
		_w24420_,
		_w24947_
	);
	LUT2 #(
		.INIT('h2)
	) name14435 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24948_
	);
	LUT2 #(
		.INIT('h8)
	) name14436 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24949_
	);
	LUT4 #(
		.INIT('h777f)
	) name14437 (
		_w24568_,
		_w24573_,
		_w24948_,
		_w24949_,
		_w24950_
	);
	LUT4 #(
		.INIT('h5700)
	) name14438 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[1]/NET0131 ,
		_w24567_,
		_w24571_,
		_w24950_,
		_w24951_
	);
	LUT4 #(
		.INIT('h222a)
	) name14439 (
		md_pad_i_pad,
		_w24568_,
		_w24572_,
		_w24573_,
		_w24952_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name14440 (
		_w24567_,
		_w24571_,
		_w24946_,
		_w24952_,
		_w24953_
	);
	LUT3 #(
		.INIT('h15)
	) name14441 (
		_w24947_,
		_w24951_,
		_w24953_,
		_w24954_
	);
	LUT4 #(
		.INIT('h222a)
	) name14442 (
		\miim1_shftrg_ShiftReg_reg[6]/NET0131 ,
		_w24568_,
		_w24572_,
		_w24573_,
		_w24955_
	);
	LUT3 #(
		.INIT('h10)
	) name14443 (
		_w24567_,
		_w24571_,
		_w24955_,
		_w24956_
	);
	LUT2 #(
		.INIT('h2)
	) name14444 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[7]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24957_
	);
	LUT3 #(
		.INIT('h80)
	) name14445 (
		_w24568_,
		_w24573_,
		_w24957_,
		_w24958_
	);
	LUT2 #(
		.INIT('h8)
	) name14446 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[7]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24959_
	);
	LUT3 #(
		.INIT('h80)
	) name14447 (
		_w24568_,
		_w24573_,
		_w24959_,
		_w24960_
	);
	LUT3 #(
		.INIT('h80)
	) name14448 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[0]/NET0131 ,
		_w24568_,
		_w24572_,
		_w24961_
	);
	LUT3 #(
		.INIT('h01)
	) name14449 (
		_w24958_,
		_w24960_,
		_w24961_,
		_w24962_
	);
	LUT4 #(
		.INIT('he2ee)
	) name14450 (
		\miim1_shftrg_ShiftReg_reg[7]/NET0131 ,
		_w24561_,
		_w24956_,
		_w24962_,
		_w24963_
	);
	LUT3 #(
		.INIT('h64)
	) name14451 (
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		_w11890_,
		_w24535_,
		_w24964_
	);
	LUT3 #(
		.INIT('h87)
	) name14452 (
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w24965_
	);
	LUT4 #(
		.INIT('h008f)
	) name14453 (
		_w11866_,
		_w11867_,
		_w11883_,
		_w24965_,
		_w24966_
	);
	LUT2 #(
		.INIT('h4)
	) name14454 (
		_w11882_,
		_w24966_,
		_w24967_
	);
	LUT3 #(
		.INIT('ha8)
	) name14455 (
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w11882_,
		_w11884_,
		_w24968_
	);
	LUT3 #(
		.INIT('hec)
	) name14456 (
		_w24535_,
		_w24967_,
		_w24968_,
		_w24969_
	);
	LUT2 #(
		.INIT('h4)
	) name14457 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		_w24970_
	);
	LUT4 #(
		.INIT('h0001)
	) name14458 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24971_
	);
	LUT3 #(
		.INIT('ha8)
	) name14459 (
		\wishbone_rx_fifo_fifo_reg[0][0]/P0001 ,
		_w24970_,
		_w24971_,
		_w24972_
	);
	LUT4 #(
		.INIT('h8000)
	) name14460 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24973_
	);
	LUT4 #(
		.INIT('h0200)
	) name14461 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24974_
	);
	LUT4 #(
		.INIT('h135f)
	) name14462 (
		\wishbone_rx_fifo_fifo_reg[15][0]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][0]/P0001 ,
		_w24973_,
		_w24974_,
		_w24975_
	);
	LUT4 #(
		.INIT('h0100)
	) name14463 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24976_
	);
	LUT4 #(
		.INIT('h0002)
	) name14464 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24977_
	);
	LUT4 #(
		.INIT('h153f)
	) name14465 (
		\wishbone_rx_fifo_fifo_reg[1][0]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][0]/P0001 ,
		_w24976_,
		_w24977_,
		_w24978_
	);
	LUT4 #(
		.INIT('h0040)
	) name14466 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24979_
	);
	LUT4 #(
		.INIT('h0400)
	) name14467 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24980_
	);
	LUT4 #(
		.INIT('h153f)
	) name14468 (
		\wishbone_rx_fifo_fifo_reg[10][0]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][0]/P0001 ,
		_w24979_,
		_w24980_,
		_w24981_
	);
	LUT4 #(
		.INIT('h0080)
	) name14469 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24982_
	);
	LUT4 #(
		.INIT('h0010)
	) name14470 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24983_
	);
	LUT4 #(
		.INIT('h153f)
	) name14471 (
		\wishbone_rx_fifo_fifo_reg[4][0]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][0]/P0001 ,
		_w24982_,
		_w24983_,
		_w24984_
	);
	LUT4 #(
		.INIT('h8000)
	) name14472 (
		_w24975_,
		_w24978_,
		_w24981_,
		_w24984_,
		_w24985_
	);
	LUT4 #(
		.INIT('h0008)
	) name14473 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24986_
	);
	LUT2 #(
		.INIT('h8)
	) name14474 (
		\wishbone_rx_fifo_fifo_reg[3][0]/P0001 ,
		_w24986_,
		_w24987_
	);
	LUT4 #(
		.INIT('h2000)
	) name14475 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24988_
	);
	LUT4 #(
		.INIT('h0800)
	) name14476 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24989_
	);
	LUT4 #(
		.INIT('h153f)
	) name14477 (
		\wishbone_rx_fifo_fifo_reg[11][0]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[13][0]/P0001 ,
		_w24988_,
		_w24989_,
		_w24990_
	);
	LUT4 #(
		.INIT('h0004)
	) name14478 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24991_
	);
	LUT4 #(
		.INIT('h0020)
	) name14479 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24992_
	);
	LUT4 #(
		.INIT('h135f)
	) name14480 (
		\wishbone_rx_fifo_fifo_reg[2][0]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][0]/P0001 ,
		_w24991_,
		_w24992_,
		_w24993_
	);
	LUT4 #(
		.INIT('h4000)
	) name14481 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24994_
	);
	LUT4 #(
		.INIT('h1000)
	) name14482 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24995_
	);
	LUT4 #(
		.INIT('h153f)
	) name14483 (
		\wishbone_rx_fifo_fifo_reg[12][0]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[14][0]/P0001 ,
		_w24994_,
		_w24995_,
		_w24996_
	);
	LUT4 #(
		.INIT('h4000)
	) name14484 (
		_w24987_,
		_w24990_,
		_w24993_,
		_w24996_,
		_w24997_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14485 (
		_w24970_,
		_w24972_,
		_w24985_,
		_w24997_,
		_w24998_
	);
	LUT4 #(
		.INIT('h153f)
	) name14486 (
		\wishbone_rx_fifo_fifo_reg[11][10]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[3][10]/P0001 ,
		_w24986_,
		_w24989_,
		_w24999_
	);
	LUT4 #(
		.INIT('h135f)
	) name14487 (
		\wishbone_rx_fifo_fifo_reg[15][10]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][10]/P0001 ,
		_w24973_,
		_w24979_,
		_w25000_
	);
	LUT3 #(
		.INIT('h13)
	) name14488 (
		\wishbone_rx_fifo_fifo_reg[5][10]/P0001 ,
		_w24970_,
		_w24992_,
		_w25001_
	);
	LUT4 #(
		.INIT('h135f)
	) name14489 (
		\wishbone_rx_fifo_fifo_reg[1][10]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][10]/P0001 ,
		_w24977_,
		_w24982_,
		_w25002_
	);
	LUT4 #(
		.INIT('h8000)
	) name14490 (
		_w24999_,
		_w25000_,
		_w25001_,
		_w25002_,
		_w25003_
	);
	LUT4 #(
		.INIT('h135f)
	) name14491 (
		\wishbone_rx_fifo_fifo_reg[10][10]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[12][10]/P0001 ,
		_w24980_,
		_w24995_,
		_w25004_
	);
	LUT4 #(
		.INIT('h153f)
	) name14492 (
		\wishbone_rx_fifo_fifo_reg[13][10]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][10]/P0001 ,
		_w24974_,
		_w24988_,
		_w25005_
	);
	LUT4 #(
		.INIT('h153f)
	) name14493 (
		\wishbone_rx_fifo_fifo_reg[14][10]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][10]/P0001 ,
		_w24991_,
		_w24994_,
		_w25006_
	);
	LUT4 #(
		.INIT('h153f)
	) name14494 (
		\wishbone_rx_fifo_fifo_reg[4][10]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][10]/P0001 ,
		_w24976_,
		_w24983_,
		_w25007_
	);
	LUT4 #(
		.INIT('h8000)
	) name14495 (
		_w25004_,
		_w25005_,
		_w25006_,
		_w25007_,
		_w25008_
	);
	LUT3 #(
		.INIT('h04)
	) name14496 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[0][10]/P0001 ,
		_w25009_
	);
	LUT2 #(
		.INIT('h8)
	) name14497 (
		\wishbone_rx_fifo_fifo_reg[0][10]/P0001 ,
		_w24971_,
		_w25010_
	);
	LUT4 #(
		.INIT('hff07)
	) name14498 (
		_w25003_,
		_w25008_,
		_w25009_,
		_w25010_,
		_w25011_
	);
	LUT3 #(
		.INIT('ha8)
	) name14499 (
		\wishbone_rx_fifo_fifo_reg[0][11]/P0001 ,
		_w24970_,
		_w24971_,
		_w25012_
	);
	LUT4 #(
		.INIT('h153f)
	) name14500 (
		\wishbone_rx_fifo_fifo_reg[5][11]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][11]/P0001 ,
		_w24974_,
		_w24992_,
		_w25013_
	);
	LUT4 #(
		.INIT('h135f)
	) name14501 (
		\wishbone_rx_fifo_fifo_reg[10][11]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[13][11]/P0001 ,
		_w24980_,
		_w24988_,
		_w25014_
	);
	LUT4 #(
		.INIT('h153f)
	) name14502 (
		\wishbone_rx_fifo_fifo_reg[12][11]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][11]/P0001 ,
		_w24979_,
		_w24995_,
		_w25015_
	);
	LUT4 #(
		.INIT('h153f)
	) name14503 (
		\wishbone_rx_fifo_fifo_reg[11][11]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][11]/P0001 ,
		_w24976_,
		_w24989_,
		_w25016_
	);
	LUT4 #(
		.INIT('h8000)
	) name14504 (
		_w25013_,
		_w25014_,
		_w25015_,
		_w25016_,
		_w25017_
	);
	LUT2 #(
		.INIT('h8)
	) name14505 (
		\wishbone_rx_fifo_fifo_reg[2][11]/P0001 ,
		_w24991_,
		_w25018_
	);
	LUT4 #(
		.INIT('h153f)
	) name14506 (
		\wishbone_rx_fifo_fifo_reg[14][11]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][11]/P0001 ,
		_w24982_,
		_w24994_,
		_w25019_
	);
	LUT4 #(
		.INIT('h135f)
	) name14507 (
		\wishbone_rx_fifo_fifo_reg[15][11]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][11]/P0001 ,
		_w24973_,
		_w24977_,
		_w25020_
	);
	LUT4 #(
		.INIT('h153f)
	) name14508 (
		\wishbone_rx_fifo_fifo_reg[3][11]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][11]/P0001 ,
		_w24983_,
		_w24986_,
		_w25021_
	);
	LUT4 #(
		.INIT('h4000)
	) name14509 (
		_w25018_,
		_w25019_,
		_w25020_,
		_w25021_,
		_w25022_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14510 (
		_w24970_,
		_w25012_,
		_w25017_,
		_w25022_,
		_w25023_
	);
	LUT4 #(
		.INIT('h135f)
	) name14511 (
		\wishbone_rx_fifo_fifo_reg[11][12]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][12]/P0001 ,
		_w24989_,
		_w24992_,
		_w25024_
	);
	LUT4 #(
		.INIT('h153f)
	) name14512 (
		\wishbone_rx_fifo_fifo_reg[10][12]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][12]/P0001 ,
		_w24977_,
		_w24980_,
		_w25025_
	);
	LUT3 #(
		.INIT('h13)
	) name14513 (
		\wishbone_rx_fifo_fifo_reg[3][12]/P0001 ,
		_w24970_,
		_w24986_,
		_w25026_
	);
	LUT4 #(
		.INIT('h153f)
	) name14514 (
		\wishbone_rx_fifo_fifo_reg[14][12]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][12]/P0001 ,
		_w24991_,
		_w24994_,
		_w25027_
	);
	LUT4 #(
		.INIT('h8000)
	) name14515 (
		_w25024_,
		_w25025_,
		_w25026_,
		_w25027_,
		_w25028_
	);
	LUT4 #(
		.INIT('h153f)
	) name14516 (
		\wishbone_rx_fifo_fifo_reg[12][12]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][12]/P0001 ,
		_w24974_,
		_w24995_,
		_w25029_
	);
	LUT4 #(
		.INIT('h153f)
	) name14517 (
		\wishbone_rx_fifo_fifo_reg[13][12]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][12]/P0001 ,
		_w24979_,
		_w24988_,
		_w25030_
	);
	LUT4 #(
		.INIT('h153f)
	) name14518 (
		\wishbone_rx_fifo_fifo_reg[4][12]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][12]/P0001 ,
		_w24976_,
		_w24983_,
		_w25031_
	);
	LUT4 #(
		.INIT('h135f)
	) name14519 (
		\wishbone_rx_fifo_fifo_reg[15][12]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][12]/P0001 ,
		_w24973_,
		_w24982_,
		_w25032_
	);
	LUT4 #(
		.INIT('h8000)
	) name14520 (
		_w25029_,
		_w25030_,
		_w25031_,
		_w25032_,
		_w25033_
	);
	LUT3 #(
		.INIT('h04)
	) name14521 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[0][12]/P0001 ,
		_w25034_
	);
	LUT2 #(
		.INIT('h8)
	) name14522 (
		\wishbone_rx_fifo_fifo_reg[0][12]/P0001 ,
		_w24971_,
		_w25035_
	);
	LUT4 #(
		.INIT('hff07)
	) name14523 (
		_w25028_,
		_w25033_,
		_w25034_,
		_w25035_,
		_w25036_
	);
	LUT3 #(
		.INIT('ha8)
	) name14524 (
		\wishbone_rx_fifo_fifo_reg[0][13]/P0001 ,
		_w24970_,
		_w24971_,
		_w25037_
	);
	LUT4 #(
		.INIT('h135f)
	) name14525 (
		\wishbone_rx_fifo_fifo_reg[10][13]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][13]/P0001 ,
		_w24980_,
		_w24992_,
		_w25038_
	);
	LUT4 #(
		.INIT('h153f)
	) name14526 (
		\wishbone_rx_fifo_fifo_reg[14][13]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][13]/P0001 ,
		_w24983_,
		_w24994_,
		_w25039_
	);
	LUT4 #(
		.INIT('h153f)
	) name14527 (
		\wishbone_rx_fifo_fifo_reg[3][13]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][13]/P0001 ,
		_w24974_,
		_w24986_,
		_w25040_
	);
	LUT4 #(
		.INIT('h153f)
	) name14528 (
		\wishbone_rx_fifo_fifo_reg[7][13]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][13]/P0001 ,
		_w24976_,
		_w24982_,
		_w25041_
	);
	LUT4 #(
		.INIT('h8000)
	) name14529 (
		_w25038_,
		_w25039_,
		_w25040_,
		_w25041_,
		_w25042_
	);
	LUT2 #(
		.INIT('h8)
	) name14530 (
		\wishbone_rx_fifo_fifo_reg[6][13]/P0001 ,
		_w24979_,
		_w25043_
	);
	LUT4 #(
		.INIT('h153f)
	) name14531 (
		\wishbone_rx_fifo_fifo_reg[11][13]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[15][13]/P0001 ,
		_w24973_,
		_w24989_,
		_w25044_
	);
	LUT4 #(
		.INIT('h153f)
	) name14532 (
		\wishbone_rx_fifo_fifo_reg[13][13]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][13]/P0001 ,
		_w24977_,
		_w24988_,
		_w25045_
	);
	LUT4 #(
		.INIT('h153f)
	) name14533 (
		\wishbone_rx_fifo_fifo_reg[12][13]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][13]/P0001 ,
		_w24991_,
		_w24995_,
		_w25046_
	);
	LUT4 #(
		.INIT('h4000)
	) name14534 (
		_w25043_,
		_w25044_,
		_w25045_,
		_w25046_,
		_w25047_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14535 (
		_w24970_,
		_w25037_,
		_w25042_,
		_w25047_,
		_w25048_
	);
	LUT4 #(
		.INIT('h153f)
	) name14536 (
		\wishbone_rx_fifo_fifo_reg[11][14]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[3][14]/P0001 ,
		_w24986_,
		_w24989_,
		_w25049_
	);
	LUT4 #(
		.INIT('h153f)
	) name14537 (
		\wishbone_rx_fifo_fifo_reg[6][14]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][14]/P0001 ,
		_w24976_,
		_w24979_,
		_w25050_
	);
	LUT3 #(
		.INIT('h13)
	) name14538 (
		\wishbone_rx_fifo_fifo_reg[12][14]/P0001 ,
		_w24970_,
		_w24995_,
		_w25051_
	);
	LUT4 #(
		.INIT('h135f)
	) name14539 (
		\wishbone_rx_fifo_fifo_reg[2][14]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][14]/P0001 ,
		_w24991_,
		_w24992_,
		_w25052_
	);
	LUT4 #(
		.INIT('h8000)
	) name14540 (
		_w25049_,
		_w25050_,
		_w25051_,
		_w25052_,
		_w25053_
	);
	LUT4 #(
		.INIT('h153f)
	) name14541 (
		\wishbone_rx_fifo_fifo_reg[10][14]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][14]/P0001 ,
		_w24977_,
		_w24980_,
		_w25054_
	);
	LUT4 #(
		.INIT('h153f)
	) name14542 (
		\wishbone_rx_fifo_fifo_reg[4][14]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][14]/P0001 ,
		_w24974_,
		_w24983_,
		_w25055_
	);
	LUT4 #(
		.INIT('h153f)
	) name14543 (
		\wishbone_rx_fifo_fifo_reg[13][14]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[15][14]/P0001 ,
		_w24973_,
		_w24988_,
		_w25056_
	);
	LUT4 #(
		.INIT('h153f)
	) name14544 (
		\wishbone_rx_fifo_fifo_reg[14][14]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][14]/P0001 ,
		_w24982_,
		_w24994_,
		_w25057_
	);
	LUT4 #(
		.INIT('h8000)
	) name14545 (
		_w25054_,
		_w25055_,
		_w25056_,
		_w25057_,
		_w25058_
	);
	LUT3 #(
		.INIT('h04)
	) name14546 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[0][14]/P0001 ,
		_w25059_
	);
	LUT2 #(
		.INIT('h8)
	) name14547 (
		\wishbone_rx_fifo_fifo_reg[0][14]/P0001 ,
		_w24971_,
		_w25060_
	);
	LUT4 #(
		.INIT('hff07)
	) name14548 (
		_w25053_,
		_w25058_,
		_w25059_,
		_w25060_,
		_w25061_
	);
	LUT3 #(
		.INIT('ha8)
	) name14549 (
		\wishbone_rx_fifo_fifo_reg[0][15]/P0001 ,
		_w24970_,
		_w24971_,
		_w25062_
	);
	LUT4 #(
		.INIT('h153f)
	) name14550 (
		\wishbone_rx_fifo_fifo_reg[14][15]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][15]/P0001 ,
		_w24979_,
		_w24994_,
		_w25063_
	);
	LUT4 #(
		.INIT('h153f)
	) name14551 (
		\wishbone_rx_fifo_fifo_reg[10][15]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][15]/P0001 ,
		_w24977_,
		_w24980_,
		_w25064_
	);
	LUT4 #(
		.INIT('h153f)
	) name14552 (
		\wishbone_rx_fifo_fifo_reg[12][15]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][15]/P0001 ,
		_w24992_,
		_w24995_,
		_w25065_
	);
	LUT4 #(
		.INIT('h153f)
	) name14553 (
		\wishbone_rx_fifo_fifo_reg[4][15]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][15]/P0001 ,
		_w24976_,
		_w24983_,
		_w25066_
	);
	LUT4 #(
		.INIT('h8000)
	) name14554 (
		_w25063_,
		_w25064_,
		_w25065_,
		_w25066_,
		_w25067_
	);
	LUT2 #(
		.INIT('h8)
	) name14555 (
		\wishbone_rx_fifo_fifo_reg[11][15]/P0001 ,
		_w24989_,
		_w25068_
	);
	LUT4 #(
		.INIT('h135f)
	) name14556 (
		\wishbone_rx_fifo_fifo_reg[15][15]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[3][15]/P0001 ,
		_w24973_,
		_w24986_,
		_w25069_
	);
	LUT4 #(
		.INIT('h153f)
	) name14557 (
		\wishbone_rx_fifo_fifo_reg[2][15]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][15]/P0001 ,
		_w24982_,
		_w24991_,
		_w25070_
	);
	LUT4 #(
		.INIT('h153f)
	) name14558 (
		\wishbone_rx_fifo_fifo_reg[13][15]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][15]/P0001 ,
		_w24974_,
		_w24988_,
		_w25071_
	);
	LUT4 #(
		.INIT('h4000)
	) name14559 (
		_w25068_,
		_w25069_,
		_w25070_,
		_w25071_,
		_w25072_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14560 (
		_w24970_,
		_w25062_,
		_w25067_,
		_w25072_,
		_w25073_
	);
	LUT4 #(
		.INIT('h153f)
	) name14561 (
		\wishbone_rx_fifo_fifo_reg[11][16]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][16]/P0001 ,
		_w24974_,
		_w24989_,
		_w25074_
	);
	LUT4 #(
		.INIT('h135f)
	) name14562 (
		\wishbone_rx_fifo_fifo_reg[15][16]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][16]/P0001 ,
		_w24973_,
		_w24979_,
		_w25075_
	);
	LUT3 #(
		.INIT('h13)
	) name14563 (
		\wishbone_rx_fifo_fifo_reg[12][16]/P0001 ,
		_w24970_,
		_w24995_,
		_w25076_
	);
	LUT4 #(
		.INIT('h135f)
	) name14564 (
		\wishbone_rx_fifo_fifo_reg[1][16]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[3][16]/P0001 ,
		_w24977_,
		_w24986_,
		_w25077_
	);
	LUT4 #(
		.INIT('h8000)
	) name14565 (
		_w25074_,
		_w25075_,
		_w25076_,
		_w25077_,
		_w25078_
	);
	LUT4 #(
		.INIT('h135f)
	) name14566 (
		\wishbone_rx_fifo_fifo_reg[10][16]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][16]/P0001 ,
		_w24980_,
		_w24992_,
		_w25079_
	);
	LUT4 #(
		.INIT('h153f)
	) name14567 (
		\wishbone_rx_fifo_fifo_reg[2][16]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][16]/P0001 ,
		_w24983_,
		_w24991_,
		_w25080_
	);
	LUT4 #(
		.INIT('h153f)
	) name14568 (
		\wishbone_rx_fifo_fifo_reg[7][16]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][16]/P0001 ,
		_w24976_,
		_w24982_,
		_w25081_
	);
	LUT4 #(
		.INIT('h135f)
	) name14569 (
		\wishbone_rx_fifo_fifo_reg[13][16]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[14][16]/P0001 ,
		_w24988_,
		_w24994_,
		_w25082_
	);
	LUT4 #(
		.INIT('h8000)
	) name14570 (
		_w25079_,
		_w25080_,
		_w25081_,
		_w25082_,
		_w25083_
	);
	LUT3 #(
		.INIT('h04)
	) name14571 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[0][16]/P0001 ,
		_w25084_
	);
	LUT2 #(
		.INIT('h8)
	) name14572 (
		\wishbone_rx_fifo_fifo_reg[0][16]/P0001 ,
		_w24971_,
		_w25085_
	);
	LUT4 #(
		.INIT('hff07)
	) name14573 (
		_w25078_,
		_w25083_,
		_w25084_,
		_w25085_,
		_w25086_
	);
	LUT3 #(
		.INIT('ha8)
	) name14574 (
		\wishbone_rx_fifo_fifo_reg[0][17]/P0001 ,
		_w24970_,
		_w24971_,
		_w25087_
	);
	LUT4 #(
		.INIT('h153f)
	) name14575 (
		\wishbone_rx_fifo_fifo_reg[14][17]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][17]/P0001 ,
		_w24974_,
		_w24994_,
		_w25088_
	);
	LUT4 #(
		.INIT('h153f)
	) name14576 (
		\wishbone_rx_fifo_fifo_reg[10][17]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][17]/P0001 ,
		_w24977_,
		_w24980_,
		_w25089_
	);
	LUT4 #(
		.INIT('h153f)
	) name14577 (
		\wishbone_rx_fifo_fifo_reg[12][17]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][17]/P0001 ,
		_w24992_,
		_w24995_,
		_w25090_
	);
	LUT4 #(
		.INIT('h153f)
	) name14578 (
		\wishbone_rx_fifo_fifo_reg[4][17]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][17]/P0001 ,
		_w24976_,
		_w24983_,
		_w25091_
	);
	LUT4 #(
		.INIT('h8000)
	) name14579 (
		_w25088_,
		_w25089_,
		_w25090_,
		_w25091_,
		_w25092_
	);
	LUT2 #(
		.INIT('h8)
	) name14580 (
		\wishbone_rx_fifo_fifo_reg[11][17]/P0001 ,
		_w24989_,
		_w25093_
	);
	LUT4 #(
		.INIT('h135f)
	) name14581 (
		\wishbone_rx_fifo_fifo_reg[15][17]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[3][17]/P0001 ,
		_w24973_,
		_w24986_,
		_w25094_
	);
	LUT4 #(
		.INIT('h153f)
	) name14582 (
		\wishbone_rx_fifo_fifo_reg[2][17]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][17]/P0001 ,
		_w24982_,
		_w24991_,
		_w25095_
	);
	LUT4 #(
		.INIT('h153f)
	) name14583 (
		\wishbone_rx_fifo_fifo_reg[13][17]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][17]/P0001 ,
		_w24979_,
		_w24988_,
		_w25096_
	);
	LUT4 #(
		.INIT('h4000)
	) name14584 (
		_w25093_,
		_w25094_,
		_w25095_,
		_w25096_,
		_w25097_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14585 (
		_w24970_,
		_w25087_,
		_w25092_,
		_w25097_,
		_w25098_
	);
	LUT3 #(
		.INIT('ha8)
	) name14586 (
		\wishbone_rx_fifo_fifo_reg[0][18]/P0001 ,
		_w24970_,
		_w24971_,
		_w25099_
	);
	LUT4 #(
		.INIT('h153f)
	) name14587 (
		\wishbone_rx_fifo_fifo_reg[10][18]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][18]/P0001 ,
		_w24979_,
		_w24980_,
		_w25100_
	);
	LUT4 #(
		.INIT('h153f)
	) name14588 (
		\wishbone_rx_fifo_fifo_reg[12][18]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][18]/P0001 ,
		_w24983_,
		_w24995_,
		_w25101_
	);
	LUT4 #(
		.INIT('h153f)
	) name14589 (
		\wishbone_rx_fifo_fifo_reg[3][18]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][18]/P0001 ,
		_w24974_,
		_w24986_,
		_w25102_
	);
	LUT4 #(
		.INIT('h153f)
	) name14590 (
		\wishbone_rx_fifo_fifo_reg[5][18]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][18]/P0001 ,
		_w24982_,
		_w24992_,
		_w25103_
	);
	LUT4 #(
		.INIT('h8000)
	) name14591 (
		_w25100_,
		_w25101_,
		_w25102_,
		_w25103_,
		_w25104_
	);
	LUT2 #(
		.INIT('h8)
	) name14592 (
		\wishbone_rx_fifo_fifo_reg[15][18]/P0001 ,
		_w24973_,
		_w25105_
	);
	LUT4 #(
		.INIT('h153f)
	) name14593 (
		\wishbone_rx_fifo_fifo_reg[11][18]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][18]/P0001 ,
		_w24976_,
		_w24989_,
		_w25106_
	);
	LUT4 #(
		.INIT('h153f)
	) name14594 (
		\wishbone_rx_fifo_fifo_reg[13][18]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][18]/P0001 ,
		_w24977_,
		_w24988_,
		_w25107_
	);
	LUT4 #(
		.INIT('h153f)
	) name14595 (
		\wishbone_rx_fifo_fifo_reg[14][18]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][18]/P0001 ,
		_w24991_,
		_w24994_,
		_w25108_
	);
	LUT4 #(
		.INIT('h4000)
	) name14596 (
		_w25105_,
		_w25106_,
		_w25107_,
		_w25108_,
		_w25109_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14597 (
		_w24970_,
		_w25099_,
		_w25104_,
		_w25109_,
		_w25110_
	);
	LUT3 #(
		.INIT('ha8)
	) name14598 (
		\wishbone_rx_fifo_fifo_reg[0][19]/P0001 ,
		_w24970_,
		_w24971_,
		_w25111_
	);
	LUT4 #(
		.INIT('h153f)
	) name14599 (
		\wishbone_rx_fifo_fifo_reg[2][19]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[3][19]/P0001 ,
		_w24986_,
		_w24991_,
		_w25112_
	);
	LUT4 #(
		.INIT('h135f)
	) name14600 (
		\wishbone_rx_fifo_fifo_reg[4][19]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][19]/P0001 ,
		_w24983_,
		_w24992_,
		_w25113_
	);
	LUT4 #(
		.INIT('h153f)
	) name14601 (
		\wishbone_rx_fifo_fifo_reg[8][19]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][19]/P0001 ,
		_w24974_,
		_w24976_,
		_w25114_
	);
	LUT4 #(
		.INIT('h153f)
	) name14602 (
		\wishbone_rx_fifo_fifo_reg[12][19]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[13][19]/P0001 ,
		_w24988_,
		_w24995_,
		_w25115_
	);
	LUT4 #(
		.INIT('h8000)
	) name14603 (
		_w25112_,
		_w25113_,
		_w25114_,
		_w25115_,
		_w25116_
	);
	LUT2 #(
		.INIT('h8)
	) name14604 (
		\wishbone_rx_fifo_fifo_reg[14][19]/P0001 ,
		_w24994_,
		_w25117_
	);
	LUT4 #(
		.INIT('h135f)
	) name14605 (
		\wishbone_rx_fifo_fifo_reg[15][19]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][19]/P0001 ,
		_w24973_,
		_w24979_,
		_w25118_
	);
	LUT4 #(
		.INIT('h135f)
	) name14606 (
		\wishbone_rx_fifo_fifo_reg[10][19]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][19]/P0001 ,
		_w24980_,
		_w24982_,
		_w25119_
	);
	LUT4 #(
		.INIT('h153f)
	) name14607 (
		\wishbone_rx_fifo_fifo_reg[11][19]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][19]/P0001 ,
		_w24977_,
		_w24989_,
		_w25120_
	);
	LUT4 #(
		.INIT('h4000)
	) name14608 (
		_w25117_,
		_w25118_,
		_w25119_,
		_w25120_,
		_w25121_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14609 (
		_w24970_,
		_w25111_,
		_w25116_,
		_w25121_,
		_w25122_
	);
	LUT4 #(
		.INIT('h153f)
	) name14610 (
		\wishbone_rx_fifo_fifo_reg[11][1]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][1]/P0001 ,
		_w24974_,
		_w24989_,
		_w25123_
	);
	LUT4 #(
		.INIT('h135f)
	) name14611 (
		\wishbone_rx_fifo_fifo_reg[15][1]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][1]/P0001 ,
		_w24973_,
		_w24979_,
		_w25124_
	);
	LUT3 #(
		.INIT('h13)
	) name14612 (
		\wishbone_rx_fifo_fifo_reg[5][1]/P0001 ,
		_w24970_,
		_w24992_,
		_w25125_
	);
	LUT4 #(
		.INIT('h135f)
	) name14613 (
		\wishbone_rx_fifo_fifo_reg[1][1]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[3][1]/P0001 ,
		_w24977_,
		_w24986_,
		_w25126_
	);
	LUT4 #(
		.INIT('h8000)
	) name14614 (
		_w25123_,
		_w25124_,
		_w25125_,
		_w25126_,
		_w25127_
	);
	LUT4 #(
		.INIT('h135f)
	) name14615 (
		\wishbone_rx_fifo_fifo_reg[10][1]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[14][1]/P0001 ,
		_w24980_,
		_w24994_,
		_w25128_
	);
	LUT4 #(
		.INIT('h153f)
	) name14616 (
		\wishbone_rx_fifo_fifo_reg[2][1]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][1]/P0001 ,
		_w24983_,
		_w24991_,
		_w25129_
	);
	LUT4 #(
		.INIT('h153f)
	) name14617 (
		\wishbone_rx_fifo_fifo_reg[7][1]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][1]/P0001 ,
		_w24976_,
		_w24982_,
		_w25130_
	);
	LUT4 #(
		.INIT('h153f)
	) name14618 (
		\wishbone_rx_fifo_fifo_reg[12][1]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[13][1]/P0001 ,
		_w24988_,
		_w24995_,
		_w25131_
	);
	LUT4 #(
		.INIT('h8000)
	) name14619 (
		_w25128_,
		_w25129_,
		_w25130_,
		_w25131_,
		_w25132_
	);
	LUT3 #(
		.INIT('h04)
	) name14620 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[0][1]/P0001 ,
		_w25133_
	);
	LUT2 #(
		.INIT('h8)
	) name14621 (
		\wishbone_rx_fifo_fifo_reg[0][1]/P0001 ,
		_w24971_,
		_w25134_
	);
	LUT4 #(
		.INIT('hff07)
	) name14622 (
		_w25127_,
		_w25132_,
		_w25133_,
		_w25134_,
		_w25135_
	);
	LUT4 #(
		.INIT('h153f)
	) name14623 (
		\wishbone_rx_fifo_fifo_reg[14][20]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][20]/P0001 ,
		_w24977_,
		_w24994_,
		_w25136_
	);
	LUT4 #(
		.INIT('h153f)
	) name14624 (
		\wishbone_rx_fifo_fifo_reg[2][20]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][20]/P0001 ,
		_w24979_,
		_w24991_,
		_w25137_
	);
	LUT3 #(
		.INIT('h13)
	) name14625 (
		\wishbone_rx_fifo_fifo_reg[10][20]/P0001 ,
		_w24970_,
		_w24980_,
		_w25138_
	);
	LUT4 #(
		.INIT('h153f)
	) name14626 (
		\wishbone_rx_fifo_fifo_reg[11][20]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[13][20]/P0001 ,
		_w24988_,
		_w24989_,
		_w25139_
	);
	LUT4 #(
		.INIT('h8000)
	) name14627 (
		_w25136_,
		_w25137_,
		_w25138_,
		_w25139_,
		_w25140_
	);
	LUT4 #(
		.INIT('h135f)
	) name14628 (
		\wishbone_rx_fifo_fifo_reg[15][20]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][20]/P0001 ,
		_w24973_,
		_w24992_,
		_w25141_
	);
	LUT4 #(
		.INIT('h153f)
	) name14629 (
		\wishbone_rx_fifo_fifo_reg[12][20]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][20]/P0001 ,
		_w24976_,
		_w24995_,
		_w25142_
	);
	LUT4 #(
		.INIT('h153f)
	) name14630 (
		\wishbone_rx_fifo_fifo_reg[7][20]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][20]/P0001 ,
		_w24974_,
		_w24982_,
		_w25143_
	);
	LUT4 #(
		.INIT('h153f)
	) name14631 (
		\wishbone_rx_fifo_fifo_reg[3][20]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][20]/P0001 ,
		_w24983_,
		_w24986_,
		_w25144_
	);
	LUT4 #(
		.INIT('h8000)
	) name14632 (
		_w25141_,
		_w25142_,
		_w25143_,
		_w25144_,
		_w25145_
	);
	LUT3 #(
		.INIT('h04)
	) name14633 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[0][20]/P0001 ,
		_w25146_
	);
	LUT2 #(
		.INIT('h8)
	) name14634 (
		\wishbone_rx_fifo_fifo_reg[0][20]/P0001 ,
		_w24971_,
		_w25147_
	);
	LUT4 #(
		.INIT('hff07)
	) name14635 (
		_w25140_,
		_w25145_,
		_w25146_,
		_w25147_,
		_w25148_
	);
	LUT3 #(
		.INIT('ha8)
	) name14636 (
		\wishbone_rx_fifo_fifo_reg[0][21]/P0001 ,
		_w24970_,
		_w24971_,
		_w25149_
	);
	LUT4 #(
		.INIT('h153f)
	) name14637 (
		\wishbone_rx_fifo_fifo_reg[5][21]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][21]/P0001 ,
		_w24982_,
		_w24992_,
		_w25150_
	);
	LUT4 #(
		.INIT('h135f)
	) name14638 (
		\wishbone_rx_fifo_fifo_reg[13][21]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][21]/P0001 ,
		_w24988_,
		_w24991_,
		_w25151_
	);
	LUT4 #(
		.INIT('h153f)
	) name14639 (
		\wishbone_rx_fifo_fifo_reg[12][21]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][21]/P0001 ,
		_w24979_,
		_w24995_,
		_w25152_
	);
	LUT4 #(
		.INIT('h153f)
	) name14640 (
		\wishbone_rx_fifo_fifo_reg[11][21]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][21]/P0001 ,
		_w24974_,
		_w24989_,
		_w25153_
	);
	LUT4 #(
		.INIT('h8000)
	) name14641 (
		_w25150_,
		_w25151_,
		_w25152_,
		_w25153_,
		_w25154_
	);
	LUT2 #(
		.INIT('h8)
	) name14642 (
		\wishbone_rx_fifo_fifo_reg[3][21]/P0001 ,
		_w24986_,
		_w25155_
	);
	LUT4 #(
		.INIT('h153f)
	) name14643 (
		\wishbone_rx_fifo_fifo_reg[10][21]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][21]/P0001 ,
		_w24977_,
		_w24980_,
		_w25156_
	);
	LUT4 #(
		.INIT('h135f)
	) name14644 (
		\wishbone_rx_fifo_fifo_reg[15][21]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][21]/P0001 ,
		_w24973_,
		_w24983_,
		_w25157_
	);
	LUT4 #(
		.INIT('h153f)
	) name14645 (
		\wishbone_rx_fifo_fifo_reg[14][21]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][21]/P0001 ,
		_w24976_,
		_w24994_,
		_w25158_
	);
	LUT4 #(
		.INIT('h4000)
	) name14646 (
		_w25155_,
		_w25156_,
		_w25157_,
		_w25158_,
		_w25159_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14647 (
		_w24970_,
		_w25149_,
		_w25154_,
		_w25159_,
		_w25160_
	);
	LUT3 #(
		.INIT('ha8)
	) name14648 (
		\wishbone_rx_fifo_fifo_reg[0][22]/P0001 ,
		_w24970_,
		_w24971_,
		_w25161_
	);
	LUT4 #(
		.INIT('h153f)
	) name14649 (
		\wishbone_rx_fifo_fifo_reg[5][22]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][22]/P0001 ,
		_w24982_,
		_w24992_,
		_w25162_
	);
	LUT4 #(
		.INIT('h135f)
	) name14650 (
		\wishbone_rx_fifo_fifo_reg[13][22]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][22]/P0001 ,
		_w24988_,
		_w24991_,
		_w25163_
	);
	LUT4 #(
		.INIT('h153f)
	) name14651 (
		\wishbone_rx_fifo_fifo_reg[12][22]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][22]/P0001 ,
		_w24979_,
		_w24995_,
		_w25164_
	);
	LUT4 #(
		.INIT('h153f)
	) name14652 (
		\wishbone_rx_fifo_fifo_reg[11][22]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][22]/P0001 ,
		_w24974_,
		_w24989_,
		_w25165_
	);
	LUT4 #(
		.INIT('h8000)
	) name14653 (
		_w25162_,
		_w25163_,
		_w25164_,
		_w25165_,
		_w25166_
	);
	LUT2 #(
		.INIT('h8)
	) name14654 (
		\wishbone_rx_fifo_fifo_reg[3][22]/P0001 ,
		_w24986_,
		_w25167_
	);
	LUT4 #(
		.INIT('h153f)
	) name14655 (
		\wishbone_rx_fifo_fifo_reg[10][22]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][22]/P0001 ,
		_w24977_,
		_w24980_,
		_w25168_
	);
	LUT4 #(
		.INIT('h135f)
	) name14656 (
		\wishbone_rx_fifo_fifo_reg[15][22]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][22]/P0001 ,
		_w24973_,
		_w24983_,
		_w25169_
	);
	LUT4 #(
		.INIT('h153f)
	) name14657 (
		\wishbone_rx_fifo_fifo_reg[14][22]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][22]/P0001 ,
		_w24976_,
		_w24994_,
		_w25170_
	);
	LUT4 #(
		.INIT('h4000)
	) name14658 (
		_w25167_,
		_w25168_,
		_w25169_,
		_w25170_,
		_w25171_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14659 (
		_w24970_,
		_w25161_,
		_w25166_,
		_w25171_,
		_w25172_
	);
	LUT3 #(
		.INIT('ha8)
	) name14660 (
		\wishbone_rx_fifo_fifo_reg[0][23]/P0001 ,
		_w24970_,
		_w24971_,
		_w25173_
	);
	LUT4 #(
		.INIT('h153f)
	) name14661 (
		\wishbone_rx_fifo_fifo_reg[5][23]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][23]/P0001 ,
		_w24982_,
		_w24992_,
		_w25174_
	);
	LUT4 #(
		.INIT('h135f)
	) name14662 (
		\wishbone_rx_fifo_fifo_reg[13][23]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][23]/P0001 ,
		_w24988_,
		_w24991_,
		_w25175_
	);
	LUT4 #(
		.INIT('h153f)
	) name14663 (
		\wishbone_rx_fifo_fifo_reg[12][23]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][23]/P0001 ,
		_w24979_,
		_w24995_,
		_w25176_
	);
	LUT4 #(
		.INIT('h153f)
	) name14664 (
		\wishbone_rx_fifo_fifo_reg[11][23]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][23]/P0001 ,
		_w24974_,
		_w24989_,
		_w25177_
	);
	LUT4 #(
		.INIT('h8000)
	) name14665 (
		_w25174_,
		_w25175_,
		_w25176_,
		_w25177_,
		_w25178_
	);
	LUT2 #(
		.INIT('h8)
	) name14666 (
		\wishbone_rx_fifo_fifo_reg[3][23]/P0001 ,
		_w24986_,
		_w25179_
	);
	LUT4 #(
		.INIT('h153f)
	) name14667 (
		\wishbone_rx_fifo_fifo_reg[10][23]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][23]/P0001 ,
		_w24977_,
		_w24980_,
		_w25180_
	);
	LUT4 #(
		.INIT('h135f)
	) name14668 (
		\wishbone_rx_fifo_fifo_reg[15][23]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][23]/P0001 ,
		_w24973_,
		_w24983_,
		_w25181_
	);
	LUT4 #(
		.INIT('h153f)
	) name14669 (
		\wishbone_rx_fifo_fifo_reg[14][23]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][23]/P0001 ,
		_w24976_,
		_w24994_,
		_w25182_
	);
	LUT4 #(
		.INIT('h4000)
	) name14670 (
		_w25179_,
		_w25180_,
		_w25181_,
		_w25182_,
		_w25183_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14671 (
		_w24970_,
		_w25173_,
		_w25178_,
		_w25183_,
		_w25184_
	);
	LUT3 #(
		.INIT('ha8)
	) name14672 (
		\wishbone_rx_fifo_fifo_reg[0][24]/P0001 ,
		_w24970_,
		_w24971_,
		_w25185_
	);
	LUT4 #(
		.INIT('h153f)
	) name14673 (
		\wishbone_rx_fifo_fifo_reg[2][24]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[3][24]/P0001 ,
		_w24986_,
		_w24991_,
		_w25186_
	);
	LUT4 #(
		.INIT('h135f)
	) name14674 (
		\wishbone_rx_fifo_fifo_reg[4][24]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][24]/P0001 ,
		_w24983_,
		_w24992_,
		_w25187_
	);
	LUT4 #(
		.INIT('h153f)
	) name14675 (
		\wishbone_rx_fifo_fifo_reg[8][24]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][24]/P0001 ,
		_w24974_,
		_w24976_,
		_w25188_
	);
	LUT4 #(
		.INIT('h153f)
	) name14676 (
		\wishbone_rx_fifo_fifo_reg[12][24]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[13][24]/P0001 ,
		_w24988_,
		_w24995_,
		_w25189_
	);
	LUT4 #(
		.INIT('h8000)
	) name14677 (
		_w25186_,
		_w25187_,
		_w25188_,
		_w25189_,
		_w25190_
	);
	LUT2 #(
		.INIT('h8)
	) name14678 (
		\wishbone_rx_fifo_fifo_reg[14][24]/P0001 ,
		_w24994_,
		_w25191_
	);
	LUT4 #(
		.INIT('h135f)
	) name14679 (
		\wishbone_rx_fifo_fifo_reg[15][24]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][24]/P0001 ,
		_w24973_,
		_w24979_,
		_w25192_
	);
	LUT4 #(
		.INIT('h135f)
	) name14680 (
		\wishbone_rx_fifo_fifo_reg[10][24]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][24]/P0001 ,
		_w24980_,
		_w24982_,
		_w25193_
	);
	LUT4 #(
		.INIT('h153f)
	) name14681 (
		\wishbone_rx_fifo_fifo_reg[11][24]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][24]/P0001 ,
		_w24977_,
		_w24989_,
		_w25194_
	);
	LUT4 #(
		.INIT('h4000)
	) name14682 (
		_w25191_,
		_w25192_,
		_w25193_,
		_w25194_,
		_w25195_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14683 (
		_w24970_,
		_w25185_,
		_w25190_,
		_w25195_,
		_w25196_
	);
	LUT3 #(
		.INIT('ha8)
	) name14684 (
		\wishbone_rx_fifo_fifo_reg[0][25]/P0001 ,
		_w24970_,
		_w24971_,
		_w25197_
	);
	LUT4 #(
		.INIT('h135f)
	) name14685 (
		\wishbone_rx_fifo_fifo_reg[15][25]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][25]/P0001 ,
		_w24973_,
		_w24974_,
		_w25198_
	);
	LUT4 #(
		.INIT('h153f)
	) name14686 (
		\wishbone_rx_fifo_fifo_reg[3][25]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][25]/P0001 ,
		_w24976_,
		_w24986_,
		_w25199_
	);
	LUT4 #(
		.INIT('h153f)
	) name14687 (
		\wishbone_rx_fifo_fifo_reg[10][25]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][25]/P0001 ,
		_w24979_,
		_w24980_,
		_w25200_
	);
	LUT4 #(
		.INIT('h153f)
	) name14688 (
		\wishbone_rx_fifo_fifo_reg[4][25]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][25]/P0001 ,
		_w24982_,
		_w24983_,
		_w25201_
	);
	LUT4 #(
		.INIT('h8000)
	) name14689 (
		_w25198_,
		_w25199_,
		_w25200_,
		_w25201_,
		_w25202_
	);
	LUT2 #(
		.INIT('h8)
	) name14690 (
		\wishbone_rx_fifo_fifo_reg[1][25]/P0001 ,
		_w24977_,
		_w25203_
	);
	LUT4 #(
		.INIT('h135f)
	) name14691 (
		\wishbone_rx_fifo_fifo_reg[13][25]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][25]/P0001 ,
		_w24988_,
		_w24991_,
		_w25204_
	);
	LUT4 #(
		.INIT('h135f)
	) name14692 (
		\wishbone_rx_fifo_fifo_reg[11][25]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][25]/P0001 ,
		_w24989_,
		_w24992_,
		_w25205_
	);
	LUT4 #(
		.INIT('h153f)
	) name14693 (
		\wishbone_rx_fifo_fifo_reg[12][25]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[14][25]/P0001 ,
		_w24994_,
		_w24995_,
		_w25206_
	);
	LUT4 #(
		.INIT('h4000)
	) name14694 (
		_w25203_,
		_w25204_,
		_w25205_,
		_w25206_,
		_w25207_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14695 (
		_w24970_,
		_w25197_,
		_w25202_,
		_w25207_,
		_w25208_
	);
	LUT3 #(
		.INIT('ha8)
	) name14696 (
		\wishbone_rx_fifo_fifo_reg[0][26]/P0001 ,
		_w24970_,
		_w24971_,
		_w25209_
	);
	LUT4 #(
		.INIT('h153f)
	) name14697 (
		\wishbone_rx_fifo_fifo_reg[5][26]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][26]/P0001 ,
		_w24976_,
		_w24992_,
		_w25210_
	);
	LUT4 #(
		.INIT('h153f)
	) name14698 (
		\wishbone_rx_fifo_fifo_reg[13][26]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][26]/P0001 ,
		_w24983_,
		_w24988_,
		_w25211_
	);
	LUT4 #(
		.INIT('h153f)
	) name14699 (
		\wishbone_rx_fifo_fifo_reg[3][26]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][26]/P0001 ,
		_w24974_,
		_w24986_,
		_w25212_
	);
	LUT4 #(
		.INIT('h135f)
	) name14700 (
		\wishbone_rx_fifo_fifo_reg[15][26]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][26]/P0001 ,
		_w24973_,
		_w24979_,
		_w25213_
	);
	LUT4 #(
		.INIT('h8000)
	) name14701 (
		_w25210_,
		_w25211_,
		_w25212_,
		_w25213_,
		_w25214_
	);
	LUT2 #(
		.INIT('h8)
	) name14702 (
		\wishbone_rx_fifo_fifo_reg[11][26]/P0001 ,
		_w24989_,
		_w25215_
	);
	LUT4 #(
		.INIT('h153f)
	) name14703 (
		\wishbone_rx_fifo_fifo_reg[10][26]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][26]/P0001 ,
		_w24977_,
		_w24980_,
		_w25216_
	);
	LUT4 #(
		.INIT('h153f)
	) name14704 (
		\wishbone_rx_fifo_fifo_reg[12][26]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[14][26]/P0001 ,
		_w24994_,
		_w24995_,
		_w25217_
	);
	LUT4 #(
		.INIT('h153f)
	) name14705 (
		\wishbone_rx_fifo_fifo_reg[2][26]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][26]/P0001 ,
		_w24982_,
		_w24991_,
		_w25218_
	);
	LUT4 #(
		.INIT('h4000)
	) name14706 (
		_w25215_,
		_w25216_,
		_w25217_,
		_w25218_,
		_w25219_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14707 (
		_w24970_,
		_w25209_,
		_w25214_,
		_w25219_,
		_w25220_
	);
	LUT4 #(
		.INIT('h153f)
	) name14708 (
		\wishbone_rx_fifo_fifo_reg[11][27]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][27]/P0001 ,
		_w24974_,
		_w24989_,
		_w25221_
	);
	LUT4 #(
		.INIT('h135f)
	) name14709 (
		\wishbone_rx_fifo_fifo_reg[15][27]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][27]/P0001 ,
		_w24973_,
		_w24979_,
		_w25222_
	);
	LUT3 #(
		.INIT('h13)
	) name14710 (
		\wishbone_rx_fifo_fifo_reg[12][27]/P0001 ,
		_w24970_,
		_w24995_,
		_w25223_
	);
	LUT4 #(
		.INIT('h135f)
	) name14711 (
		\wishbone_rx_fifo_fifo_reg[1][27]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[3][27]/P0001 ,
		_w24977_,
		_w24986_,
		_w25224_
	);
	LUT4 #(
		.INIT('h8000)
	) name14712 (
		_w25221_,
		_w25222_,
		_w25223_,
		_w25224_,
		_w25225_
	);
	LUT4 #(
		.INIT('h135f)
	) name14713 (
		\wishbone_rx_fifo_fifo_reg[10][27]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][27]/P0001 ,
		_w24980_,
		_w24992_,
		_w25226_
	);
	LUT4 #(
		.INIT('h153f)
	) name14714 (
		\wishbone_rx_fifo_fifo_reg[2][27]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][27]/P0001 ,
		_w24983_,
		_w24991_,
		_w25227_
	);
	LUT4 #(
		.INIT('h153f)
	) name14715 (
		\wishbone_rx_fifo_fifo_reg[7][27]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][27]/P0001 ,
		_w24976_,
		_w24982_,
		_w25228_
	);
	LUT4 #(
		.INIT('h135f)
	) name14716 (
		\wishbone_rx_fifo_fifo_reg[13][27]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[14][27]/P0001 ,
		_w24988_,
		_w24994_,
		_w25229_
	);
	LUT4 #(
		.INIT('h8000)
	) name14717 (
		_w25226_,
		_w25227_,
		_w25228_,
		_w25229_,
		_w25230_
	);
	LUT3 #(
		.INIT('h04)
	) name14718 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[0][27]/P0001 ,
		_w25231_
	);
	LUT2 #(
		.INIT('h8)
	) name14719 (
		\wishbone_rx_fifo_fifo_reg[0][27]/P0001 ,
		_w24971_,
		_w25232_
	);
	LUT4 #(
		.INIT('hff07)
	) name14720 (
		_w25225_,
		_w25230_,
		_w25231_,
		_w25232_,
		_w25233_
	);
	LUT4 #(
		.INIT('h135f)
	) name14721 (
		\wishbone_rx_fifo_fifo_reg[13][28]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][28]/P0001 ,
		_w24988_,
		_w24992_,
		_w25234_
	);
	LUT4 #(
		.INIT('h153f)
	) name14722 (
		\wishbone_rx_fifo_fifo_reg[6][28]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][28]/P0001 ,
		_w24976_,
		_w24979_,
		_w25235_
	);
	LUT3 #(
		.INIT('h13)
	) name14723 (
		\wishbone_rx_fifo_fifo_reg[12][28]/P0001 ,
		_w24970_,
		_w24995_,
		_w25236_
	);
	LUT4 #(
		.INIT('h135f)
	) name14724 (
		\wishbone_rx_fifo_fifo_reg[15][28]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][28]/P0001 ,
		_w24973_,
		_w24991_,
		_w25237_
	);
	LUT4 #(
		.INIT('h8000)
	) name14725 (
		_w25234_,
		_w25235_,
		_w25236_,
		_w25237_,
		_w25238_
	);
	LUT4 #(
		.INIT('h135f)
	) name14726 (
		\wishbone_rx_fifo_fifo_reg[10][28]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[14][28]/P0001 ,
		_w24980_,
		_w24994_,
		_w25239_
	);
	LUT4 #(
		.INIT('h153f)
	) name14727 (
		\wishbone_rx_fifo_fifo_reg[3][28]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][28]/P0001 ,
		_w24982_,
		_w24986_,
		_w25240_
	);
	LUT4 #(
		.INIT('h153f)
	) name14728 (
		\wishbone_rx_fifo_fifo_reg[11][28]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][28]/P0001 ,
		_w24974_,
		_w24989_,
		_w25241_
	);
	LUT4 #(
		.INIT('h135f)
	) name14729 (
		\wishbone_rx_fifo_fifo_reg[1][28]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][28]/P0001 ,
		_w24977_,
		_w24983_,
		_w25242_
	);
	LUT4 #(
		.INIT('h8000)
	) name14730 (
		_w25239_,
		_w25240_,
		_w25241_,
		_w25242_,
		_w25243_
	);
	LUT3 #(
		.INIT('h04)
	) name14731 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[0][28]/P0001 ,
		_w25244_
	);
	LUT2 #(
		.INIT('h8)
	) name14732 (
		\wishbone_rx_fifo_fifo_reg[0][28]/P0001 ,
		_w24971_,
		_w25245_
	);
	LUT4 #(
		.INIT('hff07)
	) name14733 (
		_w25238_,
		_w25243_,
		_w25244_,
		_w25245_,
		_w25246_
	);
	LUT4 #(
		.INIT('h135f)
	) name14734 (
		\wishbone_rx_fifo_fifo_reg[1][29]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][29]/P0001 ,
		_w24977_,
		_w24992_,
		_w25247_
	);
	LUT4 #(
		.INIT('h153f)
	) name14735 (
		\wishbone_rx_fifo_fifo_reg[6][29]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][29]/P0001 ,
		_w24976_,
		_w24979_,
		_w25248_
	);
	LUT3 #(
		.INIT('h13)
	) name14736 (
		\wishbone_rx_fifo_fifo_reg[10][29]/P0001 ,
		_w24970_,
		_w24980_,
		_w25249_
	);
	LUT4 #(
		.INIT('h135f)
	) name14737 (
		\wishbone_rx_fifo_fifo_reg[13][29]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[14][29]/P0001 ,
		_w24988_,
		_w24994_,
		_w25250_
	);
	LUT4 #(
		.INIT('h8000)
	) name14738 (
		_w25247_,
		_w25248_,
		_w25249_,
		_w25250_,
		_w25251_
	);
	LUT4 #(
		.INIT('h135f)
	) name14739 (
		\wishbone_rx_fifo_fifo_reg[15][29]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[3][29]/P0001 ,
		_w24973_,
		_w24986_,
		_w25252_
	);
	LUT4 #(
		.INIT('h135f)
	) name14740 (
		\wishbone_rx_fifo_fifo_reg[11][29]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][29]/P0001 ,
		_w24989_,
		_w24991_,
		_w25253_
	);
	LUT4 #(
		.INIT('h153f)
	) name14741 (
		\wishbone_rx_fifo_fifo_reg[7][29]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][29]/P0001 ,
		_w24974_,
		_w24982_,
		_w25254_
	);
	LUT4 #(
		.INIT('h153f)
	) name14742 (
		\wishbone_rx_fifo_fifo_reg[12][29]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][29]/P0001 ,
		_w24983_,
		_w24995_,
		_w25255_
	);
	LUT4 #(
		.INIT('h8000)
	) name14743 (
		_w25252_,
		_w25253_,
		_w25254_,
		_w25255_,
		_w25256_
	);
	LUT3 #(
		.INIT('h04)
	) name14744 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[0][29]/P0001 ,
		_w25257_
	);
	LUT2 #(
		.INIT('h8)
	) name14745 (
		\wishbone_rx_fifo_fifo_reg[0][29]/P0001 ,
		_w24971_,
		_w25258_
	);
	LUT4 #(
		.INIT('hff07)
	) name14746 (
		_w25251_,
		_w25256_,
		_w25257_,
		_w25258_,
		_w25259_
	);
	LUT3 #(
		.INIT('ha8)
	) name14747 (
		\wishbone_rx_fifo_fifo_reg[0][2]/P0001 ,
		_w24970_,
		_w24971_,
		_w25260_
	);
	LUT4 #(
		.INIT('h153f)
	) name14748 (
		\wishbone_rx_fifo_fifo_reg[10][2]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][2]/P0001 ,
		_w24979_,
		_w24980_,
		_w25261_
	);
	LUT4 #(
		.INIT('h153f)
	) name14749 (
		\wishbone_rx_fifo_fifo_reg[12][2]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][2]/P0001 ,
		_w24983_,
		_w24995_,
		_w25262_
	);
	LUT4 #(
		.INIT('h153f)
	) name14750 (
		\wishbone_rx_fifo_fifo_reg[3][2]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][2]/P0001 ,
		_w24974_,
		_w24986_,
		_w25263_
	);
	LUT4 #(
		.INIT('h153f)
	) name14751 (
		\wishbone_rx_fifo_fifo_reg[5][2]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][2]/P0001 ,
		_w24982_,
		_w24992_,
		_w25264_
	);
	LUT4 #(
		.INIT('h8000)
	) name14752 (
		_w25261_,
		_w25262_,
		_w25263_,
		_w25264_,
		_w25265_
	);
	LUT2 #(
		.INIT('h8)
	) name14753 (
		\wishbone_rx_fifo_fifo_reg[15][2]/P0001 ,
		_w24973_,
		_w25266_
	);
	LUT4 #(
		.INIT('h153f)
	) name14754 (
		\wishbone_rx_fifo_fifo_reg[11][2]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][2]/P0001 ,
		_w24976_,
		_w24989_,
		_w25267_
	);
	LUT4 #(
		.INIT('h153f)
	) name14755 (
		\wishbone_rx_fifo_fifo_reg[13][2]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][2]/P0001 ,
		_w24977_,
		_w24988_,
		_w25268_
	);
	LUT4 #(
		.INIT('h153f)
	) name14756 (
		\wishbone_rx_fifo_fifo_reg[14][2]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][2]/P0001 ,
		_w24991_,
		_w24994_,
		_w25269_
	);
	LUT4 #(
		.INIT('h4000)
	) name14757 (
		_w25266_,
		_w25267_,
		_w25268_,
		_w25269_,
		_w25270_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14758 (
		_w24970_,
		_w25260_,
		_w25265_,
		_w25270_,
		_w25271_
	);
	LUT3 #(
		.INIT('ha8)
	) name14759 (
		\wishbone_rx_fifo_fifo_reg[0][30]/P0001 ,
		_w24970_,
		_w24971_,
		_w25272_
	);
	LUT4 #(
		.INIT('h153f)
	) name14760 (
		\wishbone_rx_fifo_fifo_reg[13][30]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][30]/P0001 ,
		_w24974_,
		_w24988_,
		_w25273_
	);
	LUT4 #(
		.INIT('h153f)
	) name14761 (
		\wishbone_rx_fifo_fifo_reg[14][30]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][30]/P0001 ,
		_w24976_,
		_w24994_,
		_w25274_
	);
	LUT4 #(
		.INIT('h135f)
	) name14762 (
		\wishbone_rx_fifo_fifo_reg[3][30]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][30]/P0001 ,
		_w24986_,
		_w24992_,
		_w25275_
	);
	LUT4 #(
		.INIT('h135f)
	) name14763 (
		\wishbone_rx_fifo_fifo_reg[15][30]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][30]/P0001 ,
		_w24973_,
		_w24991_,
		_w25276_
	);
	LUT4 #(
		.INIT('h8000)
	) name14764 (
		_w25273_,
		_w25274_,
		_w25275_,
		_w25276_,
		_w25277_
	);
	LUT2 #(
		.INIT('h8)
	) name14765 (
		\wishbone_rx_fifo_fifo_reg[1][30]/P0001 ,
		_w24977_,
		_w25278_
	);
	LUT4 #(
		.INIT('h153f)
	) name14766 (
		\wishbone_rx_fifo_fifo_reg[4][30]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][30]/P0001 ,
		_w24979_,
		_w24983_,
		_w25279_
	);
	LUT4 #(
		.INIT('h135f)
	) name14767 (
		\wishbone_rx_fifo_fifo_reg[10][30]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][30]/P0001 ,
		_w24980_,
		_w24982_,
		_w25280_
	);
	LUT4 #(
		.INIT('h135f)
	) name14768 (
		\wishbone_rx_fifo_fifo_reg[11][30]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[12][30]/P0001 ,
		_w24989_,
		_w24995_,
		_w25281_
	);
	LUT4 #(
		.INIT('h4000)
	) name14769 (
		_w25278_,
		_w25279_,
		_w25280_,
		_w25281_,
		_w25282_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14770 (
		_w24970_,
		_w25272_,
		_w25277_,
		_w25282_,
		_w25283_
	);
	LUT4 #(
		.INIT('h153f)
	) name14771 (
		\wishbone_rx_fifo_fifo_reg[11][31]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[3][31]/P0001 ,
		_w24986_,
		_w24989_,
		_w25284_
	);
	LUT4 #(
		.INIT('h153f)
	) name14772 (
		\wishbone_rx_fifo_fifo_reg[6][31]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][31]/P0001 ,
		_w24976_,
		_w24979_,
		_w25285_
	);
	LUT3 #(
		.INIT('h13)
	) name14773 (
		\wishbone_rx_fifo_fifo_reg[12][31]/P0001 ,
		_w24970_,
		_w24995_,
		_w25286_
	);
	LUT4 #(
		.INIT('h135f)
	) name14774 (
		\wishbone_rx_fifo_fifo_reg[2][31]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][31]/P0001 ,
		_w24991_,
		_w24992_,
		_w25287_
	);
	LUT4 #(
		.INIT('h8000)
	) name14775 (
		_w25284_,
		_w25285_,
		_w25286_,
		_w25287_,
		_w25288_
	);
	LUT4 #(
		.INIT('h153f)
	) name14776 (
		\wishbone_rx_fifo_fifo_reg[10][31]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][31]/P0001 ,
		_w24977_,
		_w24980_,
		_w25289_
	);
	LUT4 #(
		.INIT('h153f)
	) name14777 (
		\wishbone_rx_fifo_fifo_reg[4][31]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][31]/P0001 ,
		_w24974_,
		_w24983_,
		_w25290_
	);
	LUT4 #(
		.INIT('h153f)
	) name14778 (
		\wishbone_rx_fifo_fifo_reg[13][31]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[15][31]/P0001 ,
		_w24973_,
		_w24988_,
		_w25291_
	);
	LUT4 #(
		.INIT('h153f)
	) name14779 (
		\wishbone_rx_fifo_fifo_reg[14][31]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][31]/P0001 ,
		_w24982_,
		_w24994_,
		_w25292_
	);
	LUT4 #(
		.INIT('h8000)
	) name14780 (
		_w25289_,
		_w25290_,
		_w25291_,
		_w25292_,
		_w25293_
	);
	LUT3 #(
		.INIT('h04)
	) name14781 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[0][31]/P0001 ,
		_w25294_
	);
	LUT2 #(
		.INIT('h8)
	) name14782 (
		\wishbone_rx_fifo_fifo_reg[0][31]/P0001 ,
		_w24971_,
		_w25295_
	);
	LUT4 #(
		.INIT('hff07)
	) name14783 (
		_w25288_,
		_w25293_,
		_w25294_,
		_w25295_,
		_w25296_
	);
	LUT3 #(
		.INIT('ha8)
	) name14784 (
		\wishbone_rx_fifo_fifo_reg[0][3]/P0001 ,
		_w24970_,
		_w24971_,
		_w25297_
	);
	LUT4 #(
		.INIT('h135f)
	) name14785 (
		\wishbone_rx_fifo_fifo_reg[1][3]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][3]/P0001 ,
		_w24977_,
		_w24992_,
		_w25298_
	);
	LUT4 #(
		.INIT('h153f)
	) name14786 (
		\wishbone_rx_fifo_fifo_reg[11][3]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][3]/P0001 ,
		_w24983_,
		_w24989_,
		_w25299_
	);
	LUT4 #(
		.INIT('h153f)
	) name14787 (
		\wishbone_rx_fifo_fifo_reg[7][3]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][3]/P0001 ,
		_w24976_,
		_w24982_,
		_w25300_
	);
	LUT4 #(
		.INIT('h135f)
	) name14788 (
		\wishbone_rx_fifo_fifo_reg[10][3]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[12][3]/P0001 ,
		_w24980_,
		_w24995_,
		_w25301_
	);
	LUT4 #(
		.INIT('h8000)
	) name14789 (
		_w25298_,
		_w25299_,
		_w25300_,
		_w25301_,
		_w25302_
	);
	LUT2 #(
		.INIT('h8)
	) name14790 (
		\wishbone_rx_fifo_fifo_reg[3][3]/P0001 ,
		_w24986_,
		_w25303_
	);
	LUT4 #(
		.INIT('h153f)
	) name14791 (
		\wishbone_rx_fifo_fifo_reg[2][3]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][3]/P0001 ,
		_w24974_,
		_w24991_,
		_w25304_
	);
	LUT4 #(
		.INIT('h153f)
	) name14792 (
		\wishbone_rx_fifo_fifo_reg[13][3]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][3]/P0001 ,
		_w24979_,
		_w24988_,
		_w25305_
	);
	LUT4 #(
		.INIT('h153f)
	) name14793 (
		\wishbone_rx_fifo_fifo_reg[14][3]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[15][3]/P0001 ,
		_w24973_,
		_w24994_,
		_w25306_
	);
	LUT4 #(
		.INIT('h4000)
	) name14794 (
		_w25303_,
		_w25304_,
		_w25305_,
		_w25306_,
		_w25307_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14795 (
		_w24970_,
		_w25297_,
		_w25302_,
		_w25307_,
		_w25308_
	);
	LUT4 #(
		.INIT('h153f)
	) name14796 (
		\wishbone_rx_fifo_fifo_reg[11][4]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[3][4]/P0001 ,
		_w24986_,
		_w24989_,
		_w25309_
	);
	LUT4 #(
		.INIT('h153f)
	) name14797 (
		\wishbone_rx_fifo_fifo_reg[8][4]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][4]/P0001 ,
		_w24974_,
		_w24976_,
		_w25310_
	);
	LUT3 #(
		.INIT('h13)
	) name14798 (
		\wishbone_rx_fifo_fifo_reg[12][4]/P0001 ,
		_w24970_,
		_w24995_,
		_w25311_
	);
	LUT4 #(
		.INIT('h135f)
	) name14799 (
		\wishbone_rx_fifo_fifo_reg[2][4]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][4]/P0001 ,
		_w24991_,
		_w24992_,
		_w25312_
	);
	LUT4 #(
		.INIT('h8000)
	) name14800 (
		_w25309_,
		_w25310_,
		_w25311_,
		_w25312_,
		_w25313_
	);
	LUT4 #(
		.INIT('h153f)
	) name14801 (
		\wishbone_rx_fifo_fifo_reg[10][4]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][4]/P0001 ,
		_w24977_,
		_w24980_,
		_w25314_
	);
	LUT4 #(
		.INIT('h153f)
	) name14802 (
		\wishbone_rx_fifo_fifo_reg[4][4]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][4]/P0001 ,
		_w24979_,
		_w24983_,
		_w25315_
	);
	LUT4 #(
		.INIT('h153f)
	) name14803 (
		\wishbone_rx_fifo_fifo_reg[13][4]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[15][4]/P0001 ,
		_w24973_,
		_w24988_,
		_w25316_
	);
	LUT4 #(
		.INIT('h153f)
	) name14804 (
		\wishbone_rx_fifo_fifo_reg[14][4]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][4]/P0001 ,
		_w24982_,
		_w24994_,
		_w25317_
	);
	LUT4 #(
		.INIT('h8000)
	) name14805 (
		_w25314_,
		_w25315_,
		_w25316_,
		_w25317_,
		_w25318_
	);
	LUT3 #(
		.INIT('h04)
	) name14806 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[0][4]/P0001 ,
		_w25319_
	);
	LUT2 #(
		.INIT('h8)
	) name14807 (
		\wishbone_rx_fifo_fifo_reg[0][4]/P0001 ,
		_w24971_,
		_w25320_
	);
	LUT4 #(
		.INIT('hff07)
	) name14808 (
		_w25313_,
		_w25318_,
		_w25319_,
		_w25320_,
		_w25321_
	);
	LUT4 #(
		.INIT('h153f)
	) name14809 (
		\wishbone_rx_fifo_fifo_reg[13][5]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][5]/P0001 ,
		_w24983_,
		_w24988_,
		_w25322_
	);
	LUT4 #(
		.INIT('h153f)
	) name14810 (
		\wishbone_rx_fifo_fifo_reg[12][5]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][5]/P0001 ,
		_w24991_,
		_w24995_,
		_w25323_
	);
	LUT3 #(
		.INIT('h13)
	) name14811 (
		\wishbone_rx_fifo_fifo_reg[10][5]/P0001 ,
		_w24970_,
		_w24980_,
		_w25324_
	);
	LUT4 #(
		.INIT('h153f)
	) name14812 (
		\wishbone_rx_fifo_fifo_reg[1][5]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][5]/P0001 ,
		_w24976_,
		_w24977_,
		_w25325_
	);
	LUT4 #(
		.INIT('h8000)
	) name14813 (
		_w25322_,
		_w25323_,
		_w25324_,
		_w25325_,
		_w25326_
	);
	LUT4 #(
		.INIT('h135f)
	) name14814 (
		\wishbone_rx_fifo_fifo_reg[6][5]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][5]/P0001 ,
		_w24979_,
		_w24982_,
		_w25327_
	);
	LUT4 #(
		.INIT('h153f)
	) name14815 (
		\wishbone_rx_fifo_fifo_reg[5][5]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][5]/P0001 ,
		_w24974_,
		_w24992_,
		_w25328_
	);
	LUT4 #(
		.INIT('h135f)
	) name14816 (
		\wishbone_rx_fifo_fifo_reg[15][5]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[3][5]/P0001 ,
		_w24973_,
		_w24986_,
		_w25329_
	);
	LUT4 #(
		.INIT('h135f)
	) name14817 (
		\wishbone_rx_fifo_fifo_reg[11][5]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[14][5]/P0001 ,
		_w24989_,
		_w24994_,
		_w25330_
	);
	LUT4 #(
		.INIT('h8000)
	) name14818 (
		_w25327_,
		_w25328_,
		_w25329_,
		_w25330_,
		_w25331_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name14819 (
		\wishbone_rx_fifo_fifo_reg[0][5]/P0001 ,
		_w24971_,
		_w25326_,
		_w25331_,
		_w25332_
	);
	LUT3 #(
		.INIT('h15)
	) name14820 (
		_w24970_,
		_w25326_,
		_w25331_,
		_w25333_
	);
	LUT2 #(
		.INIT('he)
	) name14821 (
		_w25332_,
		_w25333_,
		_w25334_
	);
	LUT3 #(
		.INIT('ha8)
	) name14822 (
		\wishbone_rx_fifo_fifo_reg[0][6]/P0001 ,
		_w24970_,
		_w24971_,
		_w25335_
	);
	LUT4 #(
		.INIT('h153f)
	) name14823 (
		\wishbone_rx_fifo_fifo_reg[6][6]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][6]/P0001 ,
		_w24974_,
		_w24979_,
		_w25336_
	);
	LUT4 #(
		.INIT('h135f)
	) name14824 (
		\wishbone_rx_fifo_fifo_reg[1][6]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][6]/P0001 ,
		_w24977_,
		_w24991_,
		_w25337_
	);
	LUT4 #(
		.INIT('h153f)
	) name14825 (
		\wishbone_rx_fifo_fifo_reg[14][6]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][6]/P0001 ,
		_w24992_,
		_w24994_,
		_w25338_
	);
	LUT4 #(
		.INIT('h153f)
	) name14826 (
		\wishbone_rx_fifo_fifo_reg[12][6]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[3][6]/P0001 ,
		_w24986_,
		_w24995_,
		_w25339_
	);
	LUT4 #(
		.INIT('h8000)
	) name14827 (
		_w25336_,
		_w25337_,
		_w25338_,
		_w25339_,
		_w25340_
	);
	LUT2 #(
		.INIT('h8)
	) name14828 (
		\wishbone_rx_fifo_fifo_reg[7][6]/P0001 ,
		_w24982_,
		_w25341_
	);
	LUT4 #(
		.INIT('h153f)
	) name14829 (
		\wishbone_rx_fifo_fifo_reg[10][6]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][6]/P0001 ,
		_w24976_,
		_w24980_,
		_w25342_
	);
	LUT4 #(
		.INIT('h153f)
	) name14830 (
		\wishbone_rx_fifo_fifo_reg[11][6]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][6]/P0001 ,
		_w24983_,
		_w24989_,
		_w25343_
	);
	LUT4 #(
		.INIT('h153f)
	) name14831 (
		\wishbone_rx_fifo_fifo_reg[13][6]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[15][6]/P0001 ,
		_w24973_,
		_w24988_,
		_w25344_
	);
	LUT4 #(
		.INIT('h4000)
	) name14832 (
		_w25341_,
		_w25342_,
		_w25343_,
		_w25344_,
		_w25345_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14833 (
		_w24970_,
		_w25335_,
		_w25340_,
		_w25345_,
		_w25346_
	);
	LUT4 #(
		.INIT('h153f)
	) name14834 (
		\wishbone_rx_fifo_fifo_reg[13][7]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][7]/P0001 ,
		_w24974_,
		_w24988_,
		_w25347_
	);
	LUT4 #(
		.INIT('h153f)
	) name14835 (
		\wishbone_rx_fifo_fifo_reg[12][7]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][7]/P0001 ,
		_w24979_,
		_w24995_,
		_w25348_
	);
	LUT3 #(
		.INIT('h13)
	) name14836 (
		\wishbone_rx_fifo_fifo_reg[3][7]/P0001 ,
		_w24970_,
		_w24986_,
		_w25349_
	);
	LUT4 #(
		.INIT('h135f)
	) name14837 (
		\wishbone_rx_fifo_fifo_reg[15][7]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][7]/P0001 ,
		_w24973_,
		_w24991_,
		_w25350_
	);
	LUT4 #(
		.INIT('h8000)
	) name14838 (
		_w25347_,
		_w25348_,
		_w25349_,
		_w25350_,
		_w25351_
	);
	LUT4 #(
		.INIT('h153f)
	) name14839 (
		\wishbone_rx_fifo_fifo_reg[5][7]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][7]/P0001 ,
		_w24976_,
		_w24992_,
		_w25352_
	);
	LUT4 #(
		.INIT('h153f)
	) name14840 (
		\wishbone_rx_fifo_fifo_reg[11][7]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][7]/P0001 ,
		_w24982_,
		_w24989_,
		_w25353_
	);
	LUT4 #(
		.INIT('h135f)
	) name14841 (
		\wishbone_rx_fifo_fifo_reg[10][7]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[14][7]/P0001 ,
		_w24980_,
		_w24994_,
		_w25354_
	);
	LUT4 #(
		.INIT('h135f)
	) name14842 (
		\wishbone_rx_fifo_fifo_reg[1][7]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[4][7]/P0001 ,
		_w24977_,
		_w24983_,
		_w25355_
	);
	LUT4 #(
		.INIT('h8000)
	) name14843 (
		_w25352_,
		_w25353_,
		_w25354_,
		_w25355_,
		_w25356_
	);
	LUT3 #(
		.INIT('h04)
	) name14844 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[0][7]/P0001 ,
		_w25357_
	);
	LUT2 #(
		.INIT('h8)
	) name14845 (
		\wishbone_rx_fifo_fifo_reg[0][7]/P0001 ,
		_w24971_,
		_w25358_
	);
	LUT4 #(
		.INIT('hff07)
	) name14846 (
		_w25351_,
		_w25356_,
		_w25357_,
		_w25358_,
		_w25359_
	);
	LUT3 #(
		.INIT('ha8)
	) name14847 (
		\wishbone_rx_fifo_fifo_reg[0][8]/P0001 ,
		_w24970_,
		_w24971_,
		_w25360_
	);
	LUT4 #(
		.INIT('h135f)
	) name14848 (
		\wishbone_rx_fifo_fifo_reg[13][8]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][8]/P0001 ,
		_w24988_,
		_w24992_,
		_w25361_
	);
	LUT4 #(
		.INIT('h153f)
	) name14849 (
		\wishbone_rx_fifo_fifo_reg[7][8]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][8]/P0001 ,
		_w24974_,
		_w24982_,
		_w25362_
	);
	LUT4 #(
		.INIT('h153f)
	) name14850 (
		\wishbone_rx_fifo_fifo_reg[3][8]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][8]/P0001 ,
		_w24979_,
		_w24986_,
		_w25363_
	);
	LUT4 #(
		.INIT('h153f)
	) name14851 (
		\wishbone_rx_fifo_fifo_reg[12][8]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[2][8]/P0001 ,
		_w24991_,
		_w24995_,
		_w25364_
	);
	LUT4 #(
		.INIT('h8000)
	) name14852 (
		_w25361_,
		_w25362_,
		_w25363_,
		_w25364_,
		_w25365_
	);
	LUT2 #(
		.INIT('h8)
	) name14853 (
		\wishbone_rx_fifo_fifo_reg[1][8]/P0001 ,
		_w24977_,
		_w25366_
	);
	LUT4 #(
		.INIT('h153f)
	) name14854 (
		\wishbone_rx_fifo_fifo_reg[4][8]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][8]/P0001 ,
		_w24976_,
		_w24983_,
		_w25367_
	);
	LUT4 #(
		.INIT('h135f)
	) name14855 (
		\wishbone_rx_fifo_fifo_reg[10][8]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[14][8]/P0001 ,
		_w24980_,
		_w24994_,
		_w25368_
	);
	LUT4 #(
		.INIT('h153f)
	) name14856 (
		\wishbone_rx_fifo_fifo_reg[11][8]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[15][8]/P0001 ,
		_w24973_,
		_w24989_,
		_w25369_
	);
	LUT4 #(
		.INIT('h4000)
	) name14857 (
		_w25366_,
		_w25367_,
		_w25368_,
		_w25369_,
		_w25370_
	);
	LUT4 #(
		.INIT('hcddd)
	) name14858 (
		_w24970_,
		_w25360_,
		_w25365_,
		_w25370_,
		_w25371_
	);
	LUT4 #(
		.INIT('h153f)
	) name14859 (
		\wishbone_rx_fifo_fifo_reg[14][9]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[9][9]/P0001 ,
		_w24974_,
		_w24994_,
		_w25372_
	);
	LUT4 #(
		.INIT('h135f)
	) name14860 (
		\wishbone_rx_fifo_fifo_reg[15][9]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[6][9]/P0001 ,
		_w24973_,
		_w24979_,
		_w25373_
	);
	LUT3 #(
		.INIT('h13)
	) name14861 (
		\wishbone_rx_fifo_fifo_reg[3][9]/P0001 ,
		_w24970_,
		_w24986_,
		_w25374_
	);
	LUT4 #(
		.INIT('h153f)
	) name14862 (
		\wishbone_rx_fifo_fifo_reg[12][9]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[5][9]/P0001 ,
		_w24992_,
		_w24995_,
		_w25375_
	);
	LUT4 #(
		.INIT('h8000)
	) name14863 (
		_w25372_,
		_w25373_,
		_w25374_,
		_w25375_,
		_w25376_
	);
	LUT4 #(
		.INIT('h153f)
	) name14864 (
		\wishbone_rx_fifo_fifo_reg[10][9]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[1][9]/P0001 ,
		_w24977_,
		_w24980_,
		_w25377_
	);
	LUT4 #(
		.INIT('h153f)
	) name14865 (
		\wishbone_rx_fifo_fifo_reg[4][9]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[8][9]/P0001 ,
		_w24976_,
		_w24983_,
		_w25378_
	);
	LUT4 #(
		.INIT('h153f)
	) name14866 (
		\wishbone_rx_fifo_fifo_reg[2][9]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[7][9]/P0001 ,
		_w24982_,
		_w24991_,
		_w25379_
	);
	LUT4 #(
		.INIT('h153f)
	) name14867 (
		\wishbone_rx_fifo_fifo_reg[11][9]/P0001 ,
		\wishbone_rx_fifo_fifo_reg[13][9]/P0001 ,
		_w24988_,
		_w24989_,
		_w25380_
	);
	LUT4 #(
		.INIT('h8000)
	) name14868 (
		_w25377_,
		_w25378_,
		_w25379_,
		_w25380_,
		_w25381_
	);
	LUT3 #(
		.INIT('h04)
	) name14869 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[0][9]/P0001 ,
		_w25382_
	);
	LUT2 #(
		.INIT('h8)
	) name14870 (
		\wishbone_rx_fifo_fifo_reg[0][9]/P0001 ,
		_w24971_,
		_w25383_
	);
	LUT4 #(
		.INIT('hff07)
	) name14871 (
		_w25376_,
		_w25381_,
		_w25382_,
		_w25383_,
		_w25384_
	);
	LUT2 #(
		.INIT('h1)
	) name14872 (
		\wishbone_TxAbortPacket_reg/NET0131 ,
		\wishbone_TxRetryPacket_reg/NET0131 ,
		_w25385_
	);
	LUT4 #(
		.INIT('h0001)
	) name14873 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25386_
	);
	LUT3 #(
		.INIT('ha2)
	) name14874 (
		\wishbone_tx_fifo_fifo_reg[0][0]/P0001 ,
		_w25385_,
		_w25386_,
		_w25387_
	);
	LUT4 #(
		.INIT('h2000)
	) name14875 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25388_
	);
	LUT4 #(
		.INIT('h4000)
	) name14876 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25389_
	);
	LUT4 #(
		.INIT('h135f)
	) name14877 (
		\wishbone_tx_fifo_fifo_reg[13][0]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[14][0]/P0001 ,
		_w25388_,
		_w25389_,
		_w25390_
	);
	LUT4 #(
		.INIT('h0200)
	) name14878 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25391_
	);
	LUT2 #(
		.INIT('h8)
	) name14879 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		_w25392_
	);
	LUT4 #(
		.INIT('h0080)
	) name14880 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25393_
	);
	LUT4 #(
		.INIT('h153f)
	) name14881 (
		\wishbone_tx_fifo_fifo_reg[7][0]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][0]/P0001 ,
		_w25391_,
		_w25393_,
		_w25394_
	);
	LUT4 #(
		.INIT('h0800)
	) name14882 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25395_
	);
	LUT4 #(
		.INIT('h0020)
	) name14883 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25396_
	);
	LUT4 #(
		.INIT('h135f)
	) name14884 (
		\wishbone_tx_fifo_fifo_reg[11][0]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][0]/P0001 ,
		_w25395_,
		_w25396_,
		_w25397_
	);
	LUT4 #(
		.INIT('h0100)
	) name14885 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25398_
	);
	LUT4 #(
		.INIT('h8000)
	) name14886 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25399_
	);
	LUT4 #(
		.INIT('h153f)
	) name14887 (
		\wishbone_tx_fifo_fifo_reg[15][0]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][0]/P0001 ,
		_w25398_,
		_w25399_,
		_w25400_
	);
	LUT4 #(
		.INIT('h8000)
	) name14888 (
		_w25390_,
		_w25394_,
		_w25397_,
		_w25400_,
		_w25401_
	);
	LUT4 #(
		.INIT('h0004)
	) name14889 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25402_
	);
	LUT2 #(
		.INIT('h8)
	) name14890 (
		\wishbone_tx_fifo_fifo_reg[2][0]/P0001 ,
		_w25402_,
		_w25403_
	);
	LUT4 #(
		.INIT('h0010)
	) name14891 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25404_
	);
	LUT4 #(
		.INIT('h0400)
	) name14892 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25405_
	);
	LUT4 #(
		.INIT('h153f)
	) name14893 (
		\wishbone_tx_fifo_fifo_reg[10][0]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][0]/P0001 ,
		_w25404_,
		_w25405_,
		_w25406_
	);
	LUT4 #(
		.INIT('h0040)
	) name14894 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25407_
	);
	LUT4 #(
		.INIT('h1000)
	) name14895 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25408_
	);
	LUT4 #(
		.INIT('h153f)
	) name14896 (
		\wishbone_tx_fifo_fifo_reg[12][0]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][0]/P0001 ,
		_w25407_,
		_w25408_,
		_w25409_
	);
	LUT4 #(
		.INIT('h0002)
	) name14897 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25410_
	);
	LUT4 #(
		.INIT('h0008)
	) name14898 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25411_
	);
	LUT4 #(
		.INIT('h135f)
	) name14899 (
		\wishbone_tx_fifo_fifo_reg[1][0]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[3][0]/P0001 ,
		_w25410_,
		_w25411_,
		_w25412_
	);
	LUT4 #(
		.INIT('h4000)
	) name14900 (
		_w25403_,
		_w25406_,
		_w25409_,
		_w25412_,
		_w25413_
	);
	LUT4 #(
		.INIT('hceee)
	) name14901 (
		_w25385_,
		_w25387_,
		_w25401_,
		_w25413_,
		_w25414_
	);
	LUT3 #(
		.INIT('ha2)
	) name14902 (
		\wishbone_tx_fifo_fifo_reg[0][10]/P0001 ,
		_w25385_,
		_w25386_,
		_w25415_
	);
	LUT4 #(
		.INIT('h153f)
	) name14903 (
		\wishbone_tx_fifo_fifo_reg[3][10]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][10]/P0001 ,
		_w25393_,
		_w25411_,
		_w25416_
	);
	LUT4 #(
		.INIT('h135f)
	) name14904 (
		\wishbone_tx_fifo_fifo_reg[14][10]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[15][10]/P0001 ,
		_w25389_,
		_w25399_,
		_w25417_
	);
	LUT4 #(
		.INIT('h135f)
	) name14905 (
		\wishbone_tx_fifo_fifo_reg[13][10]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[2][10]/P0001 ,
		_w25388_,
		_w25402_,
		_w25418_
	);
	LUT4 #(
		.INIT('h135f)
	) name14906 (
		\wishbone_tx_fifo_fifo_reg[11][10]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][10]/P0001 ,
		_w25395_,
		_w25396_,
		_w25419_
	);
	LUT4 #(
		.INIT('h8000)
	) name14907 (
		_w25416_,
		_w25417_,
		_w25418_,
		_w25419_,
		_w25420_
	);
	LUT2 #(
		.INIT('h8)
	) name14908 (
		\wishbone_tx_fifo_fifo_reg[8][10]/P0001 ,
		_w25398_,
		_w25421_
	);
	LUT4 #(
		.INIT('h135f)
	) name14909 (
		\wishbone_tx_fifo_fifo_reg[10][10]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][10]/P0001 ,
		_w25405_,
		_w25407_,
		_w25422_
	);
	LUT4 #(
		.INIT('h153f)
	) name14910 (
		\wishbone_tx_fifo_fifo_reg[12][10]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][10]/P0001 ,
		_w25404_,
		_w25408_,
		_w25423_
	);
	LUT4 #(
		.INIT('h153f)
	) name14911 (
		\wishbone_tx_fifo_fifo_reg[1][10]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][10]/P0001 ,
		_w25391_,
		_w25410_,
		_w25424_
	);
	LUT4 #(
		.INIT('h4000)
	) name14912 (
		_w25421_,
		_w25422_,
		_w25423_,
		_w25424_,
		_w25425_
	);
	LUT4 #(
		.INIT('hceee)
	) name14913 (
		_w25385_,
		_w25415_,
		_w25420_,
		_w25425_,
		_w25426_
	);
	LUT3 #(
		.INIT('ha2)
	) name14914 (
		\wishbone_tx_fifo_fifo_reg[0][11]/P0001 ,
		_w25385_,
		_w25386_,
		_w25427_
	);
	LUT4 #(
		.INIT('h153f)
	) name14915 (
		\wishbone_tx_fifo_fifo_reg[10][11]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][11]/P0001 ,
		_w25396_,
		_w25405_,
		_w25428_
	);
	LUT4 #(
		.INIT('h135f)
	) name14916 (
		\wishbone_tx_fifo_fifo_reg[14][11]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][11]/P0001 ,
		_w25389_,
		_w25404_,
		_w25429_
	);
	LUT4 #(
		.INIT('h153f)
	) name14917 (
		\wishbone_tx_fifo_fifo_reg[3][11]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][11]/P0001 ,
		_w25407_,
		_w25411_,
		_w25430_
	);
	LUT4 #(
		.INIT('h135f)
	) name14918 (
		\wishbone_tx_fifo_fifo_reg[7][11]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][11]/P0001 ,
		_w25393_,
		_w25398_,
		_w25431_
	);
	LUT4 #(
		.INIT('h8000)
	) name14919 (
		_w25428_,
		_w25429_,
		_w25430_,
		_w25431_,
		_w25432_
	);
	LUT2 #(
		.INIT('h8)
	) name14920 (
		\wishbone_tx_fifo_fifo_reg[9][11]/P0001 ,
		_w25391_,
		_w25433_
	);
	LUT4 #(
		.INIT('h135f)
	) name14921 (
		\wishbone_tx_fifo_fifo_reg[11][11]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[15][11]/P0001 ,
		_w25395_,
		_w25399_,
		_w25434_
	);
	LUT4 #(
		.INIT('h135f)
	) name14922 (
		\wishbone_tx_fifo_fifo_reg[13][11]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][11]/P0001 ,
		_w25388_,
		_w25410_,
		_w25435_
	);
	LUT4 #(
		.INIT('h153f)
	) name14923 (
		\wishbone_tx_fifo_fifo_reg[12][11]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[2][11]/P0001 ,
		_w25402_,
		_w25408_,
		_w25436_
	);
	LUT4 #(
		.INIT('h4000)
	) name14924 (
		_w25433_,
		_w25434_,
		_w25435_,
		_w25436_,
		_w25437_
	);
	LUT4 #(
		.INIT('hceee)
	) name14925 (
		_w25385_,
		_w25427_,
		_w25432_,
		_w25437_,
		_w25438_
	);
	LUT3 #(
		.INIT('ha2)
	) name14926 (
		\wishbone_tx_fifo_fifo_reg[0][12]/P0001 ,
		_w25385_,
		_w25386_,
		_w25439_
	);
	LUT4 #(
		.INIT('h153f)
	) name14927 (
		\wishbone_tx_fifo_fifo_reg[5][12]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][12]/P0001 ,
		_w25391_,
		_w25396_,
		_w25440_
	);
	LUT4 #(
		.INIT('h153f)
	) name14928 (
		\wishbone_tx_fifo_fifo_reg[10][12]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[13][12]/P0001 ,
		_w25388_,
		_w25405_,
		_w25441_
	);
	LUT4 #(
		.INIT('h153f)
	) name14929 (
		\wishbone_tx_fifo_fifo_reg[12][12]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][12]/P0001 ,
		_w25407_,
		_w25408_,
		_w25442_
	);
	LUT4 #(
		.INIT('h135f)
	) name14930 (
		\wishbone_tx_fifo_fifo_reg[11][12]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][12]/P0001 ,
		_w25395_,
		_w25398_,
		_w25443_
	);
	LUT4 #(
		.INIT('h8000)
	) name14931 (
		_w25440_,
		_w25441_,
		_w25442_,
		_w25443_,
		_w25444_
	);
	LUT2 #(
		.INIT('h8)
	) name14932 (
		\wishbone_tx_fifo_fifo_reg[2][12]/P0001 ,
		_w25402_,
		_w25445_
	);
	LUT4 #(
		.INIT('h135f)
	) name14933 (
		\wishbone_tx_fifo_fifo_reg[14][12]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][12]/P0001 ,
		_w25389_,
		_w25393_,
		_w25446_
	);
	LUT4 #(
		.INIT('h135f)
	) name14934 (
		\wishbone_tx_fifo_fifo_reg[15][12]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][12]/P0001 ,
		_w25399_,
		_w25410_,
		_w25447_
	);
	LUT4 #(
		.INIT('h153f)
	) name14935 (
		\wishbone_tx_fifo_fifo_reg[3][12]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][12]/P0001 ,
		_w25404_,
		_w25411_,
		_w25448_
	);
	LUT4 #(
		.INIT('h4000)
	) name14936 (
		_w25445_,
		_w25446_,
		_w25447_,
		_w25448_,
		_w25449_
	);
	LUT4 #(
		.INIT('hceee)
	) name14937 (
		_w25385_,
		_w25439_,
		_w25444_,
		_w25449_,
		_w25450_
	);
	LUT3 #(
		.INIT('ha2)
	) name14938 (
		\wishbone_tx_fifo_fifo_reg[0][13]/P0001 ,
		_w25385_,
		_w25386_,
		_w25451_
	);
	LUT4 #(
		.INIT('h135f)
	) name14939 (
		\wishbone_tx_fifo_fifo_reg[13][13]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][13]/P0001 ,
		_w25388_,
		_w25391_,
		_w25452_
	);
	LUT4 #(
		.INIT('h135f)
	) name14940 (
		\wishbone_tx_fifo_fifo_reg[14][13]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][13]/P0001 ,
		_w25389_,
		_w25398_,
		_w25453_
	);
	LUT4 #(
		.INIT('h153f)
	) name14941 (
		\wishbone_tx_fifo_fifo_reg[3][13]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][13]/P0001 ,
		_w25396_,
		_w25411_,
		_w25454_
	);
	LUT4 #(
		.INIT('h135f)
	) name14942 (
		\wishbone_tx_fifo_fifo_reg[15][13]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[2][13]/P0001 ,
		_w25399_,
		_w25402_,
		_w25455_
	);
	LUT4 #(
		.INIT('h8000)
	) name14943 (
		_w25452_,
		_w25453_,
		_w25454_,
		_w25455_,
		_w25456_
	);
	LUT2 #(
		.INIT('h8)
	) name14944 (
		\wishbone_tx_fifo_fifo_reg[1][13]/P0001 ,
		_w25410_,
		_w25457_
	);
	LUT4 #(
		.INIT('h135f)
	) name14945 (
		\wishbone_tx_fifo_fifo_reg[4][13]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][13]/P0001 ,
		_w25404_,
		_w25407_,
		_w25458_
	);
	LUT4 #(
		.INIT('h153f)
	) name14946 (
		\wishbone_tx_fifo_fifo_reg[10][13]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][13]/P0001 ,
		_w25393_,
		_w25405_,
		_w25459_
	);
	LUT4 #(
		.INIT('h135f)
	) name14947 (
		\wishbone_tx_fifo_fifo_reg[11][13]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[12][13]/P0001 ,
		_w25395_,
		_w25408_,
		_w25460_
	);
	LUT4 #(
		.INIT('h4000)
	) name14948 (
		_w25457_,
		_w25458_,
		_w25459_,
		_w25460_,
		_w25461_
	);
	LUT4 #(
		.INIT('hceee)
	) name14949 (
		_w25385_,
		_w25451_,
		_w25456_,
		_w25461_,
		_w25462_
	);
	LUT3 #(
		.INIT('ha2)
	) name14950 (
		\wishbone_tx_fifo_fifo_reg[0][14]/P0001 ,
		_w25385_,
		_w25386_,
		_w25463_
	);
	LUT4 #(
		.INIT('h135f)
	) name14951 (
		\wishbone_tx_fifo_fifo_reg[15][14]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][14]/P0001 ,
		_w25399_,
		_w25407_,
		_w25464_
	);
	LUT4 #(
		.INIT('h135f)
	) name14952 (
		\wishbone_tx_fifo_fifo_reg[11][14]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[3][14]/P0001 ,
		_w25395_,
		_w25411_,
		_w25465_
	);
	LUT4 #(
		.INIT('h153f)
	) name14953 (
		\wishbone_tx_fifo_fifo_reg[10][14]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][14]/P0001 ,
		_w25391_,
		_w25405_,
		_w25466_
	);
	LUT4 #(
		.INIT('h153f)
	) name14954 (
		\wishbone_tx_fifo_fifo_reg[12][14]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][14]/P0001 ,
		_w25398_,
		_w25408_,
		_w25467_
	);
	LUT4 #(
		.INIT('h8000)
	) name14955 (
		_w25464_,
		_w25465_,
		_w25466_,
		_w25467_,
		_w25468_
	);
	LUT2 #(
		.INIT('h8)
	) name14956 (
		\wishbone_tx_fifo_fifo_reg[2][14]/P0001 ,
		_w25402_,
		_w25469_
	);
	LUT4 #(
		.INIT('h153f)
	) name14957 (
		\wishbone_tx_fifo_fifo_reg[1][14]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][14]/P0001 ,
		_w25404_,
		_w25410_,
		_w25470_
	);
	LUT4 #(
		.INIT('h135f)
	) name14958 (
		\wishbone_tx_fifo_fifo_reg[14][14]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][14]/P0001 ,
		_w25389_,
		_w25396_,
		_w25471_
	);
	LUT4 #(
		.INIT('h135f)
	) name14959 (
		\wishbone_tx_fifo_fifo_reg[13][14]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][14]/P0001 ,
		_w25388_,
		_w25393_,
		_w25472_
	);
	LUT4 #(
		.INIT('h4000)
	) name14960 (
		_w25469_,
		_w25470_,
		_w25471_,
		_w25472_,
		_w25473_
	);
	LUT4 #(
		.INIT('hceee)
	) name14961 (
		_w25385_,
		_w25463_,
		_w25468_,
		_w25473_,
		_w25474_
	);
	LUT3 #(
		.INIT('ha2)
	) name14962 (
		\wishbone_tx_fifo_fifo_reg[0][15]/P0001 ,
		_w25385_,
		_w25386_,
		_w25475_
	);
	LUT4 #(
		.INIT('h153f)
	) name14963 (
		\wishbone_tx_fifo_fifo_reg[2][15]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][15]/P0001 ,
		_w25393_,
		_w25402_,
		_w25476_
	);
	LUT4 #(
		.INIT('h135f)
	) name14964 (
		\wishbone_tx_fifo_fifo_reg[14][15]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[15][15]/P0001 ,
		_w25389_,
		_w25399_,
		_w25477_
	);
	LUT4 #(
		.INIT('h135f)
	) name14965 (
		\wishbone_tx_fifo_fifo_reg[13][15]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][15]/P0001 ,
		_w25388_,
		_w25410_,
		_w25478_
	);
	LUT4 #(
		.INIT('h153f)
	) name14966 (
		\wishbone_tx_fifo_fifo_reg[3][15]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][15]/P0001 ,
		_w25396_,
		_w25411_,
		_w25479_
	);
	LUT4 #(
		.INIT('h8000)
	) name14967 (
		_w25476_,
		_w25477_,
		_w25478_,
		_w25479_,
		_w25480_
	);
	LUT2 #(
		.INIT('h8)
	) name14968 (
		\wishbone_tx_fifo_fifo_reg[8][15]/P0001 ,
		_w25398_,
		_w25481_
	);
	LUT4 #(
		.INIT('h135f)
	) name14969 (
		\wishbone_tx_fifo_fifo_reg[10][15]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][15]/P0001 ,
		_w25405_,
		_w25407_,
		_w25482_
	);
	LUT4 #(
		.INIT('h153f)
	) name14970 (
		\wishbone_tx_fifo_fifo_reg[12][15]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][15]/P0001 ,
		_w25404_,
		_w25408_,
		_w25483_
	);
	LUT4 #(
		.INIT('h153f)
	) name14971 (
		\wishbone_tx_fifo_fifo_reg[11][15]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][15]/P0001 ,
		_w25391_,
		_w25395_,
		_w25484_
	);
	LUT4 #(
		.INIT('h4000)
	) name14972 (
		_w25481_,
		_w25482_,
		_w25483_,
		_w25484_,
		_w25485_
	);
	LUT4 #(
		.INIT('hceee)
	) name14973 (
		_w25385_,
		_w25475_,
		_w25480_,
		_w25485_,
		_w25486_
	);
	LUT3 #(
		.INIT('ha2)
	) name14974 (
		\wishbone_tx_fifo_fifo_reg[0][16]/P0001 ,
		_w25385_,
		_w25386_,
		_w25487_
	);
	LUT4 #(
		.INIT('h135f)
	) name14975 (
		\wishbone_tx_fifo_fifo_reg[13][16]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][16]/P0001 ,
		_w25388_,
		_w25407_,
		_w25488_
	);
	LUT4 #(
		.INIT('h135f)
	) name14976 (
		\wishbone_tx_fifo_fifo_reg[14][16]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][16]/P0001 ,
		_w25389_,
		_w25398_,
		_w25489_
	);
	LUT4 #(
		.INIT('h153f)
	) name14977 (
		\wishbone_tx_fifo_fifo_reg[2][16]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][16]/P0001 ,
		_w25396_,
		_w25402_,
		_w25490_
	);
	LUT4 #(
		.INIT('h135f)
	) name14978 (
		\wishbone_tx_fifo_fifo_reg[15][16]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][16]/P0001 ,
		_w25399_,
		_w25410_,
		_w25491_
	);
	LUT4 #(
		.INIT('h8000)
	) name14979 (
		_w25488_,
		_w25489_,
		_w25490_,
		_w25491_,
		_w25492_
	);
	LUT2 #(
		.INIT('h8)
	) name14980 (
		\wishbone_tx_fifo_fifo_reg[11][16]/P0001 ,
		_w25395_,
		_w25493_
	);
	LUT4 #(
		.INIT('h153f)
	) name14981 (
		\wishbone_tx_fifo_fifo_reg[4][16]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][16]/P0001 ,
		_w25391_,
		_w25404_,
		_w25494_
	);
	LUT4 #(
		.INIT('h153f)
	) name14982 (
		\wishbone_tx_fifo_fifo_reg[10][16]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][16]/P0001 ,
		_w25393_,
		_w25405_,
		_w25495_
	);
	LUT4 #(
		.INIT('h135f)
	) name14983 (
		\wishbone_tx_fifo_fifo_reg[12][16]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[3][16]/P0001 ,
		_w25408_,
		_w25411_,
		_w25496_
	);
	LUT4 #(
		.INIT('h4000)
	) name14984 (
		_w25493_,
		_w25494_,
		_w25495_,
		_w25496_,
		_w25497_
	);
	LUT4 #(
		.INIT('hceee)
	) name14985 (
		_w25385_,
		_w25487_,
		_w25492_,
		_w25497_,
		_w25498_
	);
	LUT3 #(
		.INIT('ha2)
	) name14986 (
		\wishbone_tx_fifo_fifo_reg[0][17]/P0001 ,
		_w25385_,
		_w25386_,
		_w25499_
	);
	LUT4 #(
		.INIT('h153f)
	) name14987 (
		\wishbone_tx_fifo_fifo_reg[2][17]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][17]/P0001 ,
		_w25393_,
		_w25402_,
		_w25500_
	);
	LUT4 #(
		.INIT('h135f)
	) name14988 (
		\wishbone_tx_fifo_fifo_reg[14][17]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[15][17]/P0001 ,
		_w25389_,
		_w25399_,
		_w25501_
	);
	LUT4 #(
		.INIT('h135f)
	) name14989 (
		\wishbone_tx_fifo_fifo_reg[13][17]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][17]/P0001 ,
		_w25388_,
		_w25410_,
		_w25502_
	);
	LUT4 #(
		.INIT('h153f)
	) name14990 (
		\wishbone_tx_fifo_fifo_reg[3][17]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][17]/P0001 ,
		_w25396_,
		_w25411_,
		_w25503_
	);
	LUT4 #(
		.INIT('h8000)
	) name14991 (
		_w25500_,
		_w25501_,
		_w25502_,
		_w25503_,
		_w25504_
	);
	LUT2 #(
		.INIT('h8)
	) name14992 (
		\wishbone_tx_fifo_fifo_reg[8][17]/P0001 ,
		_w25398_,
		_w25505_
	);
	LUT4 #(
		.INIT('h135f)
	) name14993 (
		\wishbone_tx_fifo_fifo_reg[10][17]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][17]/P0001 ,
		_w25405_,
		_w25407_,
		_w25506_
	);
	LUT4 #(
		.INIT('h153f)
	) name14994 (
		\wishbone_tx_fifo_fifo_reg[12][17]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][17]/P0001 ,
		_w25404_,
		_w25408_,
		_w25507_
	);
	LUT4 #(
		.INIT('h153f)
	) name14995 (
		\wishbone_tx_fifo_fifo_reg[11][17]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][17]/P0001 ,
		_w25391_,
		_w25395_,
		_w25508_
	);
	LUT4 #(
		.INIT('h4000)
	) name14996 (
		_w25505_,
		_w25506_,
		_w25507_,
		_w25508_,
		_w25509_
	);
	LUT4 #(
		.INIT('hceee)
	) name14997 (
		_w25385_,
		_w25499_,
		_w25504_,
		_w25509_,
		_w25510_
	);
	LUT3 #(
		.INIT('ha2)
	) name14998 (
		\wishbone_tx_fifo_fifo_reg[0][18]/P0001 ,
		_w25385_,
		_w25386_,
		_w25511_
	);
	LUT4 #(
		.INIT('h153f)
	) name14999 (
		\wishbone_tx_fifo_fifo_reg[2][18]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][18]/P0001 ,
		_w25396_,
		_w25402_,
		_w25512_
	);
	LUT4 #(
		.INIT('h153f)
	) name15000 (
		\wishbone_tx_fifo_fifo_reg[12][18]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[14][18]/P0001 ,
		_w25389_,
		_w25408_,
		_w25513_
	);
	LUT4 #(
		.INIT('h153f)
	) name15001 (
		\wishbone_tx_fifo_fifo_reg[10][18]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][18]/P0001 ,
		_w25404_,
		_w25405_,
		_w25514_
	);
	LUT4 #(
		.INIT('h135f)
	) name15002 (
		\wishbone_tx_fifo_fifo_reg[11][18]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[3][18]/P0001 ,
		_w25395_,
		_w25411_,
		_w25515_
	);
	LUT4 #(
		.INIT('h8000)
	) name15003 (
		_w25512_,
		_w25513_,
		_w25514_,
		_w25515_,
		_w25516_
	);
	LUT2 #(
		.INIT('h8)
	) name15004 (
		\wishbone_tx_fifo_fifo_reg[8][18]/P0001 ,
		_w25398_,
		_w25517_
	);
	LUT4 #(
		.INIT('h153f)
	) name15005 (
		\wishbone_tx_fifo_fifo_reg[6][18]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][18]/P0001 ,
		_w25393_,
		_w25407_,
		_w25518_
	);
	LUT4 #(
		.INIT('h135f)
	) name15006 (
		\wishbone_tx_fifo_fifo_reg[15][18]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][18]/P0001 ,
		_w25399_,
		_w25410_,
		_w25519_
	);
	LUT4 #(
		.INIT('h135f)
	) name15007 (
		\wishbone_tx_fifo_fifo_reg[13][18]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][18]/P0001 ,
		_w25388_,
		_w25391_,
		_w25520_
	);
	LUT4 #(
		.INIT('h4000)
	) name15008 (
		_w25517_,
		_w25518_,
		_w25519_,
		_w25520_,
		_w25521_
	);
	LUT4 #(
		.INIT('hceee)
	) name15009 (
		_w25385_,
		_w25511_,
		_w25516_,
		_w25521_,
		_w25522_
	);
	LUT3 #(
		.INIT('ha2)
	) name15010 (
		\wishbone_tx_fifo_fifo_reg[0][19]/P0001 ,
		_w25385_,
		_w25386_,
		_w25523_
	);
	LUT4 #(
		.INIT('h135f)
	) name15011 (
		\wishbone_tx_fifo_fifo_reg[13][19]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][19]/P0001 ,
		_w25388_,
		_w25396_,
		_w25524_
	);
	LUT4 #(
		.INIT('h153f)
	) name15012 (
		\wishbone_tx_fifo_fifo_reg[7][19]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][19]/P0001 ,
		_w25391_,
		_w25393_,
		_w25525_
	);
	LUT4 #(
		.INIT('h153f)
	) name15013 (
		\wishbone_tx_fifo_fifo_reg[3][19]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][19]/P0001 ,
		_w25407_,
		_w25411_,
		_w25526_
	);
	LUT4 #(
		.INIT('h153f)
	) name15014 (
		\wishbone_tx_fifo_fifo_reg[12][19]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[2][19]/P0001 ,
		_w25402_,
		_w25408_,
		_w25527_
	);
	LUT4 #(
		.INIT('h8000)
	) name15015 (
		_w25524_,
		_w25525_,
		_w25526_,
		_w25527_,
		_w25528_
	);
	LUT2 #(
		.INIT('h8)
	) name15016 (
		\wishbone_tx_fifo_fifo_reg[1][19]/P0001 ,
		_w25410_,
		_w25529_
	);
	LUT4 #(
		.INIT('h153f)
	) name15017 (
		\wishbone_tx_fifo_fifo_reg[4][19]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][19]/P0001 ,
		_w25398_,
		_w25404_,
		_w25530_
	);
	LUT4 #(
		.INIT('h153f)
	) name15018 (
		\wishbone_tx_fifo_fifo_reg[10][19]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[14][19]/P0001 ,
		_w25389_,
		_w25405_,
		_w25531_
	);
	LUT4 #(
		.INIT('h135f)
	) name15019 (
		\wishbone_tx_fifo_fifo_reg[11][19]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[15][19]/P0001 ,
		_w25395_,
		_w25399_,
		_w25532_
	);
	LUT4 #(
		.INIT('h4000)
	) name15020 (
		_w25529_,
		_w25530_,
		_w25531_,
		_w25532_,
		_w25533_
	);
	LUT4 #(
		.INIT('hceee)
	) name15021 (
		_w25385_,
		_w25523_,
		_w25528_,
		_w25533_,
		_w25534_
	);
	LUT3 #(
		.INIT('ha2)
	) name15022 (
		\wishbone_tx_fifo_fifo_reg[0][1]/P0001 ,
		_w25385_,
		_w25386_,
		_w25535_
	);
	LUT4 #(
		.INIT('h153f)
	) name15023 (
		\wishbone_tx_fifo_fifo_reg[6][1]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][1]/P0001 ,
		_w25391_,
		_w25407_,
		_w25536_
	);
	LUT4 #(
		.INIT('h153f)
	) name15024 (
		\wishbone_tx_fifo_fifo_reg[1][1]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[2][1]/P0001 ,
		_w25402_,
		_w25410_,
		_w25537_
	);
	LUT4 #(
		.INIT('h135f)
	) name15025 (
		\wishbone_tx_fifo_fifo_reg[14][1]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][1]/P0001 ,
		_w25389_,
		_w25396_,
		_w25538_
	);
	LUT4 #(
		.INIT('h135f)
	) name15026 (
		\wishbone_tx_fifo_fifo_reg[12][1]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[3][1]/P0001 ,
		_w25408_,
		_w25411_,
		_w25539_
	);
	LUT4 #(
		.INIT('h8000)
	) name15027 (
		_w25536_,
		_w25537_,
		_w25538_,
		_w25539_,
		_w25540_
	);
	LUT2 #(
		.INIT('h8)
	) name15028 (
		\wishbone_tx_fifo_fifo_reg[7][1]/P0001 ,
		_w25393_,
		_w25541_
	);
	LUT4 #(
		.INIT('h153f)
	) name15029 (
		\wishbone_tx_fifo_fifo_reg[10][1]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][1]/P0001 ,
		_w25398_,
		_w25405_,
		_w25542_
	);
	LUT4 #(
		.INIT('h135f)
	) name15030 (
		\wishbone_tx_fifo_fifo_reg[11][1]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][1]/P0001 ,
		_w25395_,
		_w25404_,
		_w25543_
	);
	LUT4 #(
		.INIT('h135f)
	) name15031 (
		\wishbone_tx_fifo_fifo_reg[13][1]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[15][1]/P0001 ,
		_w25388_,
		_w25399_,
		_w25544_
	);
	LUT4 #(
		.INIT('h4000)
	) name15032 (
		_w25541_,
		_w25542_,
		_w25543_,
		_w25544_,
		_w25545_
	);
	LUT4 #(
		.INIT('hceee)
	) name15033 (
		_w25385_,
		_w25535_,
		_w25540_,
		_w25545_,
		_w25546_
	);
	LUT3 #(
		.INIT('ha2)
	) name15034 (
		\wishbone_tx_fifo_fifo_reg[0][20]/P0001 ,
		_w25385_,
		_w25386_,
		_w25547_
	);
	LUT4 #(
		.INIT('h153f)
	) name15035 (
		\wishbone_tx_fifo_fifo_reg[15][20]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][20]/P0001 ,
		_w25391_,
		_w25399_,
		_w25548_
	);
	LUT4 #(
		.INIT('h153f)
	) name15036 (
		\wishbone_tx_fifo_fifo_reg[3][20]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][20]/P0001 ,
		_w25398_,
		_w25411_,
		_w25549_
	);
	LUT4 #(
		.INIT('h135f)
	) name15037 (
		\wishbone_tx_fifo_fifo_reg[10][20]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][20]/P0001 ,
		_w25405_,
		_w25407_,
		_w25550_
	);
	LUT4 #(
		.INIT('h153f)
	) name15038 (
		\wishbone_tx_fifo_fifo_reg[4][20]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][20]/P0001 ,
		_w25393_,
		_w25404_,
		_w25551_
	);
	LUT4 #(
		.INIT('h8000)
	) name15039 (
		_w25548_,
		_w25549_,
		_w25550_,
		_w25551_,
		_w25552_
	);
	LUT2 #(
		.INIT('h8)
	) name15040 (
		\wishbone_tx_fifo_fifo_reg[1][20]/P0001 ,
		_w25410_,
		_w25553_
	);
	LUT4 #(
		.INIT('h135f)
	) name15041 (
		\wishbone_tx_fifo_fifo_reg[13][20]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[2][20]/P0001 ,
		_w25388_,
		_w25402_,
		_w25554_
	);
	LUT4 #(
		.INIT('h135f)
	) name15042 (
		\wishbone_tx_fifo_fifo_reg[11][20]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][20]/P0001 ,
		_w25395_,
		_w25396_,
		_w25555_
	);
	LUT4 #(
		.INIT('h153f)
	) name15043 (
		\wishbone_tx_fifo_fifo_reg[12][20]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[14][20]/P0001 ,
		_w25389_,
		_w25408_,
		_w25556_
	);
	LUT4 #(
		.INIT('h4000)
	) name15044 (
		_w25553_,
		_w25554_,
		_w25555_,
		_w25556_,
		_w25557_
	);
	LUT4 #(
		.INIT('hceee)
	) name15045 (
		_w25385_,
		_w25547_,
		_w25552_,
		_w25557_,
		_w25558_
	);
	LUT3 #(
		.INIT('ha2)
	) name15046 (
		\wishbone_tx_fifo_fifo_reg[0][21]/P0001 ,
		_w25385_,
		_w25386_,
		_w25559_
	);
	LUT4 #(
		.INIT('h135f)
	) name15047 (
		\wishbone_tx_fifo_fifo_reg[13][21]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[14][21]/P0001 ,
		_w25388_,
		_w25389_,
		_w25560_
	);
	LUT4 #(
		.INIT('h153f)
	) name15048 (
		\wishbone_tx_fifo_fifo_reg[7][21]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][21]/P0001 ,
		_w25391_,
		_w25393_,
		_w25561_
	);
	LUT4 #(
		.INIT('h135f)
	) name15049 (
		\wishbone_tx_fifo_fifo_reg[11][21]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][21]/P0001 ,
		_w25395_,
		_w25396_,
		_w25562_
	);
	LUT4 #(
		.INIT('h153f)
	) name15050 (
		\wishbone_tx_fifo_fifo_reg[15][21]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][21]/P0001 ,
		_w25398_,
		_w25399_,
		_w25563_
	);
	LUT4 #(
		.INIT('h8000)
	) name15051 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25564_
	);
	LUT2 #(
		.INIT('h8)
	) name15052 (
		\wishbone_tx_fifo_fifo_reg[2][21]/P0001 ,
		_w25402_,
		_w25565_
	);
	LUT4 #(
		.INIT('h153f)
	) name15053 (
		\wishbone_tx_fifo_fifo_reg[10][21]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][21]/P0001 ,
		_w25404_,
		_w25405_,
		_w25566_
	);
	LUT4 #(
		.INIT('h153f)
	) name15054 (
		\wishbone_tx_fifo_fifo_reg[12][21]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][21]/P0001 ,
		_w25407_,
		_w25408_,
		_w25567_
	);
	LUT4 #(
		.INIT('h135f)
	) name15055 (
		\wishbone_tx_fifo_fifo_reg[1][21]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[3][21]/P0001 ,
		_w25410_,
		_w25411_,
		_w25568_
	);
	LUT4 #(
		.INIT('h4000)
	) name15056 (
		_w25565_,
		_w25566_,
		_w25567_,
		_w25568_,
		_w25569_
	);
	LUT4 #(
		.INIT('hceee)
	) name15057 (
		_w25385_,
		_w25559_,
		_w25564_,
		_w25569_,
		_w25570_
	);
	LUT3 #(
		.INIT('ha2)
	) name15058 (
		\wishbone_tx_fifo_fifo_reg[0][22]/P0001 ,
		_w25385_,
		_w25386_,
		_w25571_
	);
	LUT4 #(
		.INIT('h153f)
	) name15059 (
		\wishbone_tx_fifo_fifo_reg[12][22]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[13][22]/P0001 ,
		_w25388_,
		_w25408_,
		_w25572_
	);
	LUT4 #(
		.INIT('h153f)
	) name15060 (
		\wishbone_tx_fifo_fifo_reg[7][22]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][22]/P0001 ,
		_w25391_,
		_w25393_,
		_w25573_
	);
	LUT4 #(
		.INIT('h135f)
	) name15061 (
		\wishbone_tx_fifo_fifo_reg[2][22]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][22]/P0001 ,
		_w25402_,
		_w25407_,
		_w25574_
	);
	LUT4 #(
		.INIT('h135f)
	) name15062 (
		\wishbone_tx_fifo_fifo_reg[14][22]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][22]/P0001 ,
		_w25389_,
		_w25410_,
		_w25575_
	);
	LUT4 #(
		.INIT('h8000)
	) name15063 (
		_w25572_,
		_w25573_,
		_w25574_,
		_w25575_,
		_w25576_
	);
	LUT2 #(
		.INIT('h8)
	) name15064 (
		\wishbone_tx_fifo_fifo_reg[11][22]/P0001 ,
		_w25395_,
		_w25577_
	);
	LUT4 #(
		.INIT('h153f)
	) name15065 (
		\wishbone_tx_fifo_fifo_reg[4][22]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][22]/P0001 ,
		_w25398_,
		_w25404_,
		_w25578_
	);
	LUT4 #(
		.INIT('h153f)
	) name15066 (
		\wishbone_tx_fifo_fifo_reg[10][22]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][22]/P0001 ,
		_w25396_,
		_w25405_,
		_w25579_
	);
	LUT4 #(
		.INIT('h135f)
	) name15067 (
		\wishbone_tx_fifo_fifo_reg[15][22]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[3][22]/P0001 ,
		_w25399_,
		_w25411_,
		_w25580_
	);
	LUT4 #(
		.INIT('h4000)
	) name15068 (
		_w25577_,
		_w25578_,
		_w25579_,
		_w25580_,
		_w25581_
	);
	LUT4 #(
		.INIT('hceee)
	) name15069 (
		_w25385_,
		_w25571_,
		_w25576_,
		_w25581_,
		_w25582_
	);
	LUT3 #(
		.INIT('ha2)
	) name15070 (
		\wishbone_tx_fifo_fifo_reg[0][23]/P0001 ,
		_w25385_,
		_w25386_,
		_w25583_
	);
	LUT4 #(
		.INIT('h153f)
	) name15071 (
		\wishbone_tx_fifo_fifo_reg[10][23]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][23]/P0001 ,
		_w25396_,
		_w25405_,
		_w25584_
	);
	LUT4 #(
		.INIT('h135f)
	) name15072 (
		\wishbone_tx_fifo_fifo_reg[14][23]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][23]/P0001 ,
		_w25389_,
		_w25404_,
		_w25585_
	);
	LUT4 #(
		.INIT('h135f)
	) name15073 (
		\wishbone_tx_fifo_fifo_reg[2][23]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][23]/P0001 ,
		_w25402_,
		_w25407_,
		_w25586_
	);
	LUT4 #(
		.INIT('h135f)
	) name15074 (
		\wishbone_tx_fifo_fifo_reg[7][23]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][23]/P0001 ,
		_w25393_,
		_w25398_,
		_w25587_
	);
	LUT4 #(
		.INIT('h8000)
	) name15075 (
		_w25584_,
		_w25585_,
		_w25586_,
		_w25587_,
		_w25588_
	);
	LUT2 #(
		.INIT('h8)
	) name15076 (
		\wishbone_tx_fifo_fifo_reg[9][23]/P0001 ,
		_w25391_,
		_w25589_
	);
	LUT4 #(
		.INIT('h135f)
	) name15077 (
		\wishbone_tx_fifo_fifo_reg[15][23]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[3][23]/P0001 ,
		_w25399_,
		_w25411_,
		_w25590_
	);
	LUT4 #(
		.INIT('h153f)
	) name15078 (
		\wishbone_tx_fifo_fifo_reg[11][23]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[13][23]/P0001 ,
		_w25388_,
		_w25395_,
		_w25591_
	);
	LUT4 #(
		.INIT('h135f)
	) name15079 (
		\wishbone_tx_fifo_fifo_reg[12][23]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][23]/P0001 ,
		_w25408_,
		_w25410_,
		_w25592_
	);
	LUT4 #(
		.INIT('h4000)
	) name15080 (
		_w25589_,
		_w25590_,
		_w25591_,
		_w25592_,
		_w25593_
	);
	LUT4 #(
		.INIT('hceee)
	) name15081 (
		_w25385_,
		_w25583_,
		_w25588_,
		_w25593_,
		_w25594_
	);
	LUT3 #(
		.INIT('ha2)
	) name15082 (
		\wishbone_tx_fifo_fifo_reg[0][24]/P0001 ,
		_w25385_,
		_w25386_,
		_w25595_
	);
	LUT4 #(
		.INIT('h153f)
	) name15083 (
		\wishbone_tx_fifo_fifo_reg[3][24]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][24]/P0001 ,
		_w25396_,
		_w25411_,
		_w25596_
	);
	LUT4 #(
		.INIT('h135f)
	) name15084 (
		\wishbone_tx_fifo_fifo_reg[2][24]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][24]/P0001 ,
		_w25402_,
		_w25404_,
		_w25597_
	);
	LUT4 #(
		.INIT('h135f)
	) name15085 (
		\wishbone_tx_fifo_fifo_reg[7][24]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][24]/P0001 ,
		_w25393_,
		_w25398_,
		_w25598_
	);
	LUT4 #(
		.INIT('h135f)
	) name15086 (
		\wishbone_tx_fifo_fifo_reg[10][24]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[12][24]/P0001 ,
		_w25405_,
		_w25408_,
		_w25599_
	);
	LUT4 #(
		.INIT('h8000)
	) name15087 (
		_w25596_,
		_w25597_,
		_w25598_,
		_w25599_,
		_w25600_
	);
	LUT2 #(
		.INIT('h8)
	) name15088 (
		\wishbone_tx_fifo_fifo_reg[1][24]/P0001 ,
		_w25410_,
		_w25601_
	);
	LUT4 #(
		.INIT('h153f)
	) name15089 (
		\wishbone_tx_fifo_fifo_reg[11][24]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][24]/P0001 ,
		_w25391_,
		_w25395_,
		_w25602_
	);
	LUT4 #(
		.INIT('h135f)
	) name15090 (
		\wishbone_tx_fifo_fifo_reg[13][24]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][24]/P0001 ,
		_w25388_,
		_w25407_,
		_w25603_
	);
	LUT4 #(
		.INIT('h135f)
	) name15091 (
		\wishbone_tx_fifo_fifo_reg[14][24]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[15][24]/P0001 ,
		_w25389_,
		_w25399_,
		_w25604_
	);
	LUT4 #(
		.INIT('h4000)
	) name15092 (
		_w25601_,
		_w25602_,
		_w25603_,
		_w25604_,
		_w25605_
	);
	LUT4 #(
		.INIT('hceee)
	) name15093 (
		_w25385_,
		_w25595_,
		_w25600_,
		_w25605_,
		_w25606_
	);
	LUT3 #(
		.INIT('ha2)
	) name15094 (
		\wishbone_tx_fifo_fifo_reg[0][25]/P0001 ,
		_w25385_,
		_w25386_,
		_w25607_
	);
	LUT4 #(
		.INIT('h135f)
	) name15095 (
		\wishbone_tx_fifo_fifo_reg[13][25]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[3][25]/P0001 ,
		_w25388_,
		_w25411_,
		_w25608_
	);
	LUT4 #(
		.INIT('h135f)
	) name15096 (
		\wishbone_tx_fifo_fifo_reg[11][25]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][25]/P0001 ,
		_w25395_,
		_w25396_,
		_w25609_
	);
	LUT4 #(
		.INIT('h135f)
	) name15097 (
		\wishbone_tx_fifo_fifo_reg[10][25]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][25]/P0001 ,
		_w25405_,
		_w25407_,
		_w25610_
	);
	LUT4 #(
		.INIT('h153f)
	) name15098 (
		\wishbone_tx_fifo_fifo_reg[12][25]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[14][25]/P0001 ,
		_w25389_,
		_w25408_,
		_w25611_
	);
	LUT4 #(
		.INIT('h8000)
	) name15099 (
		_w25608_,
		_w25609_,
		_w25610_,
		_w25611_,
		_w25612_
	);
	LUT2 #(
		.INIT('h8)
	) name15100 (
		\wishbone_tx_fifo_fifo_reg[15][25]/P0001 ,
		_w25399_,
		_w25613_
	);
	LUT4 #(
		.INIT('h153f)
	) name15101 (
		\wishbone_tx_fifo_fifo_reg[2][25]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][25]/P0001 ,
		_w25391_,
		_w25402_,
		_w25614_
	);
	LUT4 #(
		.INIT('h153f)
	) name15102 (
		\wishbone_tx_fifo_fifo_reg[1][25]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][25]/P0001 ,
		_w25404_,
		_w25410_,
		_w25615_
	);
	LUT4 #(
		.INIT('h135f)
	) name15103 (
		\wishbone_tx_fifo_fifo_reg[7][25]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][25]/P0001 ,
		_w25393_,
		_w25398_,
		_w25616_
	);
	LUT4 #(
		.INIT('h4000)
	) name15104 (
		_w25613_,
		_w25614_,
		_w25615_,
		_w25616_,
		_w25617_
	);
	LUT4 #(
		.INIT('hceee)
	) name15105 (
		_w25385_,
		_w25607_,
		_w25612_,
		_w25617_,
		_w25618_
	);
	LUT3 #(
		.INIT('ha2)
	) name15106 (
		\wishbone_tx_fifo_fifo_reg[0][26]/P0001 ,
		_w25385_,
		_w25386_,
		_w25619_
	);
	LUT4 #(
		.INIT('h153f)
	) name15107 (
		\wishbone_tx_fifo_fifo_reg[6][26]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][26]/P0001 ,
		_w25391_,
		_w25407_,
		_w25620_
	);
	LUT4 #(
		.INIT('h153f)
	) name15108 (
		\wishbone_tx_fifo_fifo_reg[1][26]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[2][26]/P0001 ,
		_w25402_,
		_w25410_,
		_w25621_
	);
	LUT4 #(
		.INIT('h135f)
	) name15109 (
		\wishbone_tx_fifo_fifo_reg[14][26]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][26]/P0001 ,
		_w25389_,
		_w25396_,
		_w25622_
	);
	LUT4 #(
		.INIT('h135f)
	) name15110 (
		\wishbone_tx_fifo_fifo_reg[12][26]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[3][26]/P0001 ,
		_w25408_,
		_w25411_,
		_w25623_
	);
	LUT4 #(
		.INIT('h8000)
	) name15111 (
		_w25620_,
		_w25621_,
		_w25622_,
		_w25623_,
		_w25624_
	);
	LUT2 #(
		.INIT('h8)
	) name15112 (
		\wishbone_tx_fifo_fifo_reg[7][26]/P0001 ,
		_w25393_,
		_w25625_
	);
	LUT4 #(
		.INIT('h153f)
	) name15113 (
		\wishbone_tx_fifo_fifo_reg[10][26]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][26]/P0001 ,
		_w25398_,
		_w25405_,
		_w25626_
	);
	LUT4 #(
		.INIT('h135f)
	) name15114 (
		\wishbone_tx_fifo_fifo_reg[11][26]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][26]/P0001 ,
		_w25395_,
		_w25404_,
		_w25627_
	);
	LUT4 #(
		.INIT('h135f)
	) name15115 (
		\wishbone_tx_fifo_fifo_reg[13][26]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[15][26]/P0001 ,
		_w25388_,
		_w25399_,
		_w25628_
	);
	LUT4 #(
		.INIT('h4000)
	) name15116 (
		_w25625_,
		_w25626_,
		_w25627_,
		_w25628_,
		_w25629_
	);
	LUT4 #(
		.INIT('hceee)
	) name15117 (
		_w25385_,
		_w25619_,
		_w25624_,
		_w25629_,
		_w25630_
	);
	LUT3 #(
		.INIT('ha2)
	) name15118 (
		\wishbone_tx_fifo_fifo_reg[0][27]/P0001 ,
		_w25385_,
		_w25386_,
		_w25631_
	);
	LUT4 #(
		.INIT('h135f)
	) name15119 (
		\wishbone_tx_fifo_fifo_reg[12][27]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][27]/P0001 ,
		_w25408_,
		_w25410_,
		_w25632_
	);
	LUT4 #(
		.INIT('h153f)
	) name15120 (
		\wishbone_tx_fifo_fifo_reg[11][27]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][27]/P0001 ,
		_w25391_,
		_w25395_,
		_w25633_
	);
	LUT4 #(
		.INIT('h135f)
	) name15121 (
		\wishbone_tx_fifo_fifo_reg[10][27]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][27]/P0001 ,
		_w25405_,
		_w25407_,
		_w25634_
	);
	LUT4 #(
		.INIT('h153f)
	) name15122 (
		\wishbone_tx_fifo_fifo_reg[5][27]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][27]/P0001 ,
		_w25393_,
		_w25396_,
		_w25635_
	);
	LUT4 #(
		.INIT('h8000)
	) name15123 (
		_w25632_,
		_w25633_,
		_w25634_,
		_w25635_,
		_w25636_
	);
	LUT2 #(
		.INIT('h8)
	) name15124 (
		\wishbone_tx_fifo_fifo_reg[8][27]/P0001 ,
		_w25398_,
		_w25637_
	);
	LUT4 #(
		.INIT('h135f)
	) name15125 (
		\wishbone_tx_fifo_fifo_reg[15][27]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[2][27]/P0001 ,
		_w25399_,
		_w25402_,
		_w25638_
	);
	LUT4 #(
		.INIT('h153f)
	) name15126 (
		\wishbone_tx_fifo_fifo_reg[3][27]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][27]/P0001 ,
		_w25404_,
		_w25411_,
		_w25639_
	);
	LUT4 #(
		.INIT('h135f)
	) name15127 (
		\wishbone_tx_fifo_fifo_reg[13][27]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[14][27]/P0001 ,
		_w25388_,
		_w25389_,
		_w25640_
	);
	LUT4 #(
		.INIT('h4000)
	) name15128 (
		_w25637_,
		_w25638_,
		_w25639_,
		_w25640_,
		_w25641_
	);
	LUT4 #(
		.INIT('hceee)
	) name15129 (
		_w25385_,
		_w25631_,
		_w25636_,
		_w25641_,
		_w25642_
	);
	LUT3 #(
		.INIT('ha2)
	) name15130 (
		\wishbone_tx_fifo_fifo_reg[0][28]/P0001 ,
		_w25385_,
		_w25386_,
		_w25643_
	);
	LUT4 #(
		.INIT('h135f)
	) name15131 (
		\wishbone_tx_fifo_fifo_reg[14][28]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][28]/P0001 ,
		_w25389_,
		_w25407_,
		_w25644_
	);
	LUT4 #(
		.INIT('h135f)
	) name15132 (
		\wishbone_tx_fifo_fifo_reg[10][28]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][28]/P0001 ,
		_w25405_,
		_w25410_,
		_w25645_
	);
	LUT4 #(
		.INIT('h153f)
	) name15133 (
		\wishbone_tx_fifo_fifo_reg[12][28]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][28]/P0001 ,
		_w25396_,
		_w25408_,
		_w25646_
	);
	LUT4 #(
		.INIT('h153f)
	) name15134 (
		\wishbone_tx_fifo_fifo_reg[4][28]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][28]/P0001 ,
		_w25398_,
		_w25404_,
		_w25647_
	);
	LUT4 #(
		.INIT('h8000)
	) name15135 (
		_w25644_,
		_w25645_,
		_w25646_,
		_w25647_,
		_w25648_
	);
	LUT2 #(
		.INIT('h8)
	) name15136 (
		\wishbone_tx_fifo_fifo_reg[11][28]/P0001 ,
		_w25395_,
		_w25649_
	);
	LUT4 #(
		.INIT('h135f)
	) name15137 (
		\wishbone_tx_fifo_fifo_reg[15][28]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[3][28]/P0001 ,
		_w25399_,
		_w25411_,
		_w25650_
	);
	LUT4 #(
		.INIT('h153f)
	) name15138 (
		\wishbone_tx_fifo_fifo_reg[2][28]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][28]/P0001 ,
		_w25393_,
		_w25402_,
		_w25651_
	);
	LUT4 #(
		.INIT('h135f)
	) name15139 (
		\wishbone_tx_fifo_fifo_reg[13][28]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][28]/P0001 ,
		_w25388_,
		_w25391_,
		_w25652_
	);
	LUT4 #(
		.INIT('h4000)
	) name15140 (
		_w25649_,
		_w25650_,
		_w25651_,
		_w25652_,
		_w25653_
	);
	LUT4 #(
		.INIT('hceee)
	) name15141 (
		_w25385_,
		_w25643_,
		_w25648_,
		_w25653_,
		_w25654_
	);
	LUT3 #(
		.INIT('ha2)
	) name15142 (
		\wishbone_tx_fifo_fifo_reg[0][29]/P0001 ,
		_w25385_,
		_w25386_,
		_w25655_
	);
	LUT4 #(
		.INIT('h153f)
	) name15143 (
		\wishbone_tx_fifo_fifo_reg[10][29]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[11][29]/P0001 ,
		_w25395_,
		_w25405_,
		_w25656_
	);
	LUT4 #(
		.INIT('h153f)
	) name15144 (
		\wishbone_tx_fifo_fifo_reg[4][29]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][29]/P0001 ,
		_w25398_,
		_w25404_,
		_w25657_
	);
	LUT4 #(
		.INIT('h135f)
	) name15145 (
		\wishbone_tx_fifo_fifo_reg[13][29]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[3][29]/P0001 ,
		_w25388_,
		_w25411_,
		_w25658_
	);
	LUT4 #(
		.INIT('h135f)
	) name15146 (
		\wishbone_tx_fifo_fifo_reg[12][29]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][29]/P0001 ,
		_w25408_,
		_w25410_,
		_w25659_
	);
	LUT4 #(
		.INIT('h8000)
	) name15147 (
		_w25656_,
		_w25657_,
		_w25658_,
		_w25659_,
		_w25660_
	);
	LUT2 #(
		.INIT('h8)
	) name15148 (
		\wishbone_tx_fifo_fifo_reg[15][29]/P0001 ,
		_w25399_,
		_w25661_
	);
	LUT4 #(
		.INIT('h135f)
	) name15149 (
		\wishbone_tx_fifo_fifo_reg[14][29]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][29]/P0001 ,
		_w25389_,
		_w25391_,
		_w25662_
	);
	LUT4 #(
		.INIT('h153f)
	) name15150 (
		\wishbone_tx_fifo_fifo_reg[6][29]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][29]/P0001 ,
		_w25393_,
		_w25407_,
		_w25663_
	);
	LUT4 #(
		.INIT('h153f)
	) name15151 (
		\wishbone_tx_fifo_fifo_reg[2][29]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][29]/P0001 ,
		_w25396_,
		_w25402_,
		_w25664_
	);
	LUT4 #(
		.INIT('h4000)
	) name15152 (
		_w25661_,
		_w25662_,
		_w25663_,
		_w25664_,
		_w25665_
	);
	LUT4 #(
		.INIT('hceee)
	) name15153 (
		_w25385_,
		_w25655_,
		_w25660_,
		_w25665_,
		_w25666_
	);
	LUT3 #(
		.INIT('ha2)
	) name15154 (
		\wishbone_tx_fifo_fifo_reg[0][2]/P0001 ,
		_w25385_,
		_w25386_,
		_w25667_
	);
	LUT4 #(
		.INIT('h153f)
	) name15155 (
		\wishbone_tx_fifo_fifo_reg[2][2]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][2]/P0001 ,
		_w25393_,
		_w25402_,
		_w25668_
	);
	LUT4 #(
		.INIT('h135f)
	) name15156 (
		\wishbone_tx_fifo_fifo_reg[14][2]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[15][2]/P0001 ,
		_w25389_,
		_w25399_,
		_w25669_
	);
	LUT4 #(
		.INIT('h135f)
	) name15157 (
		\wishbone_tx_fifo_fifo_reg[13][2]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][2]/P0001 ,
		_w25388_,
		_w25410_,
		_w25670_
	);
	LUT4 #(
		.INIT('h153f)
	) name15158 (
		\wishbone_tx_fifo_fifo_reg[3][2]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][2]/P0001 ,
		_w25396_,
		_w25411_,
		_w25671_
	);
	LUT4 #(
		.INIT('h8000)
	) name15159 (
		_w25668_,
		_w25669_,
		_w25670_,
		_w25671_,
		_w25672_
	);
	LUT2 #(
		.INIT('h8)
	) name15160 (
		\wishbone_tx_fifo_fifo_reg[8][2]/P0001 ,
		_w25398_,
		_w25673_
	);
	LUT4 #(
		.INIT('h135f)
	) name15161 (
		\wishbone_tx_fifo_fifo_reg[10][2]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][2]/P0001 ,
		_w25405_,
		_w25407_,
		_w25674_
	);
	LUT4 #(
		.INIT('h153f)
	) name15162 (
		\wishbone_tx_fifo_fifo_reg[12][2]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][2]/P0001 ,
		_w25404_,
		_w25408_,
		_w25675_
	);
	LUT4 #(
		.INIT('h153f)
	) name15163 (
		\wishbone_tx_fifo_fifo_reg[11][2]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][2]/P0001 ,
		_w25391_,
		_w25395_,
		_w25676_
	);
	LUT4 #(
		.INIT('h4000)
	) name15164 (
		_w25673_,
		_w25674_,
		_w25675_,
		_w25676_,
		_w25677_
	);
	LUT4 #(
		.INIT('hceee)
	) name15165 (
		_w25385_,
		_w25667_,
		_w25672_,
		_w25677_,
		_w25678_
	);
	LUT3 #(
		.INIT('ha2)
	) name15166 (
		\wishbone_tx_fifo_fifo_reg[0][30]/P0001 ,
		_w25385_,
		_w25386_,
		_w25679_
	);
	LUT4 #(
		.INIT('h153f)
	) name15167 (
		\wishbone_tx_fifo_fifo_reg[5][30]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][30]/P0001 ,
		_w25391_,
		_w25396_,
		_w25680_
	);
	LUT4 #(
		.INIT('h153f)
	) name15168 (
		\wishbone_tx_fifo_fifo_reg[10][30]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[13][30]/P0001 ,
		_w25388_,
		_w25405_,
		_w25681_
	);
	LUT4 #(
		.INIT('h153f)
	) name15169 (
		\wishbone_tx_fifo_fifo_reg[12][30]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][30]/P0001 ,
		_w25407_,
		_w25408_,
		_w25682_
	);
	LUT4 #(
		.INIT('h135f)
	) name15170 (
		\wishbone_tx_fifo_fifo_reg[11][30]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][30]/P0001 ,
		_w25395_,
		_w25398_,
		_w25683_
	);
	LUT4 #(
		.INIT('h8000)
	) name15171 (
		_w25680_,
		_w25681_,
		_w25682_,
		_w25683_,
		_w25684_
	);
	LUT2 #(
		.INIT('h8)
	) name15172 (
		\wishbone_tx_fifo_fifo_reg[2][30]/P0001 ,
		_w25402_,
		_w25685_
	);
	LUT4 #(
		.INIT('h135f)
	) name15173 (
		\wishbone_tx_fifo_fifo_reg[14][30]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][30]/P0001 ,
		_w25389_,
		_w25393_,
		_w25686_
	);
	LUT4 #(
		.INIT('h135f)
	) name15174 (
		\wishbone_tx_fifo_fifo_reg[15][30]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][30]/P0001 ,
		_w25399_,
		_w25410_,
		_w25687_
	);
	LUT4 #(
		.INIT('h153f)
	) name15175 (
		\wishbone_tx_fifo_fifo_reg[3][30]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][30]/P0001 ,
		_w25404_,
		_w25411_,
		_w25688_
	);
	LUT4 #(
		.INIT('h4000)
	) name15176 (
		_w25685_,
		_w25686_,
		_w25687_,
		_w25688_,
		_w25689_
	);
	LUT4 #(
		.INIT('hceee)
	) name15177 (
		_w25385_,
		_w25679_,
		_w25684_,
		_w25689_,
		_w25690_
	);
	LUT3 #(
		.INIT('ha2)
	) name15178 (
		\wishbone_tx_fifo_fifo_reg[0][31]/P0001 ,
		_w25385_,
		_w25386_,
		_w25691_
	);
	LUT4 #(
		.INIT('h153f)
	) name15179 (
		\wishbone_tx_fifo_fifo_reg[3][31]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][31]/P0001 ,
		_w25393_,
		_w25411_,
		_w25692_
	);
	LUT4 #(
		.INIT('h135f)
	) name15180 (
		\wishbone_tx_fifo_fifo_reg[14][31]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[15][31]/P0001 ,
		_w25389_,
		_w25399_,
		_w25693_
	);
	LUT4 #(
		.INIT('h135f)
	) name15181 (
		\wishbone_tx_fifo_fifo_reg[13][31]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[2][31]/P0001 ,
		_w25388_,
		_w25402_,
		_w25694_
	);
	LUT4 #(
		.INIT('h135f)
	) name15182 (
		\wishbone_tx_fifo_fifo_reg[11][31]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][31]/P0001 ,
		_w25395_,
		_w25396_,
		_w25695_
	);
	LUT4 #(
		.INIT('h8000)
	) name15183 (
		_w25692_,
		_w25693_,
		_w25694_,
		_w25695_,
		_w25696_
	);
	LUT2 #(
		.INIT('h8)
	) name15184 (
		\wishbone_tx_fifo_fifo_reg[8][31]/P0001 ,
		_w25398_,
		_w25697_
	);
	LUT4 #(
		.INIT('h135f)
	) name15185 (
		\wishbone_tx_fifo_fifo_reg[10][31]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][31]/P0001 ,
		_w25405_,
		_w25407_,
		_w25698_
	);
	LUT4 #(
		.INIT('h153f)
	) name15186 (
		\wishbone_tx_fifo_fifo_reg[12][31]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][31]/P0001 ,
		_w25404_,
		_w25408_,
		_w25699_
	);
	LUT4 #(
		.INIT('h153f)
	) name15187 (
		\wishbone_tx_fifo_fifo_reg[1][31]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][31]/P0001 ,
		_w25391_,
		_w25410_,
		_w25700_
	);
	LUT4 #(
		.INIT('h4000)
	) name15188 (
		_w25697_,
		_w25698_,
		_w25699_,
		_w25700_,
		_w25701_
	);
	LUT4 #(
		.INIT('hceee)
	) name15189 (
		_w25385_,
		_w25691_,
		_w25696_,
		_w25701_,
		_w25702_
	);
	LUT3 #(
		.INIT('ha2)
	) name15190 (
		\wishbone_tx_fifo_fifo_reg[0][3]/P0001 ,
		_w25385_,
		_w25386_,
		_w25703_
	);
	LUT4 #(
		.INIT('h135f)
	) name15191 (
		\wishbone_tx_fifo_fifo_reg[15][3]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][3]/P0001 ,
		_w25399_,
		_w25407_,
		_w25704_
	);
	LUT4 #(
		.INIT('h135f)
	) name15192 (
		\wishbone_tx_fifo_fifo_reg[11][3]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[3][3]/P0001 ,
		_w25395_,
		_w25411_,
		_w25705_
	);
	LUT4 #(
		.INIT('h135f)
	) name15193 (
		\wishbone_tx_fifo_fifo_reg[10][3]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[12][3]/P0001 ,
		_w25405_,
		_w25408_,
		_w25706_
	);
	LUT4 #(
		.INIT('h135f)
	) name15194 (
		\wishbone_tx_fifo_fifo_reg[5][3]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][3]/P0001 ,
		_w25396_,
		_w25398_,
		_w25707_
	);
	LUT4 #(
		.INIT('h8000)
	) name15195 (
		_w25704_,
		_w25705_,
		_w25706_,
		_w25707_,
		_w25708_
	);
	LUT2 #(
		.INIT('h8)
	) name15196 (
		\wishbone_tx_fifo_fifo_reg[2][3]/P0001 ,
		_w25402_,
		_w25709_
	);
	LUT4 #(
		.INIT('h135f)
	) name15197 (
		\wishbone_tx_fifo_fifo_reg[14][3]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][3]/P0001 ,
		_w25389_,
		_w25410_,
		_w25710_
	);
	LUT4 #(
		.INIT('h135f)
	) name15198 (
		\wishbone_tx_fifo_fifo_reg[13][3]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][3]/P0001 ,
		_w25388_,
		_w25391_,
		_w25711_
	);
	LUT4 #(
		.INIT('h153f)
	) name15199 (
		\wishbone_tx_fifo_fifo_reg[4][3]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][3]/P0001 ,
		_w25393_,
		_w25404_,
		_w25712_
	);
	LUT4 #(
		.INIT('h4000)
	) name15200 (
		_w25709_,
		_w25710_,
		_w25711_,
		_w25712_,
		_w25713_
	);
	LUT4 #(
		.INIT('hceee)
	) name15201 (
		_w25385_,
		_w25703_,
		_w25708_,
		_w25713_,
		_w25714_
	);
	LUT3 #(
		.INIT('ha2)
	) name15202 (
		\wishbone_tx_fifo_fifo_reg[0][4]/P0001 ,
		_w25385_,
		_w25386_,
		_w25715_
	);
	LUT4 #(
		.INIT('h135f)
	) name15203 (
		\wishbone_tx_fifo_fifo_reg[13][4]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][4]/P0001 ,
		_w25388_,
		_w25407_,
		_w25716_
	);
	LUT4 #(
		.INIT('h135f)
	) name15204 (
		\wishbone_tx_fifo_fifo_reg[14][4]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][4]/P0001 ,
		_w25389_,
		_w25398_,
		_w25717_
	);
	LUT4 #(
		.INIT('h153f)
	) name15205 (
		\wishbone_tx_fifo_fifo_reg[3][4]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][4]/P0001 ,
		_w25396_,
		_w25411_,
		_w25718_
	);
	LUT4 #(
		.INIT('h135f)
	) name15206 (
		\wishbone_tx_fifo_fifo_reg[15][4]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[2][4]/P0001 ,
		_w25399_,
		_w25402_,
		_w25719_
	);
	LUT4 #(
		.INIT('h8000)
	) name15207 (
		_w25716_,
		_w25717_,
		_w25718_,
		_w25719_,
		_w25720_
	);
	LUT2 #(
		.INIT('h8)
	) name15208 (
		\wishbone_tx_fifo_fifo_reg[1][4]/P0001 ,
		_w25410_,
		_w25721_
	);
	LUT4 #(
		.INIT('h153f)
	) name15209 (
		\wishbone_tx_fifo_fifo_reg[4][4]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][4]/P0001 ,
		_w25391_,
		_w25404_,
		_w25722_
	);
	LUT4 #(
		.INIT('h153f)
	) name15210 (
		\wishbone_tx_fifo_fifo_reg[10][4]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][4]/P0001 ,
		_w25393_,
		_w25405_,
		_w25723_
	);
	LUT4 #(
		.INIT('h135f)
	) name15211 (
		\wishbone_tx_fifo_fifo_reg[11][4]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[12][4]/P0001 ,
		_w25395_,
		_w25408_,
		_w25724_
	);
	LUT4 #(
		.INIT('h4000)
	) name15212 (
		_w25721_,
		_w25722_,
		_w25723_,
		_w25724_,
		_w25725_
	);
	LUT4 #(
		.INIT('hceee)
	) name15213 (
		_w25385_,
		_w25715_,
		_w25720_,
		_w25725_,
		_w25726_
	);
	LUT3 #(
		.INIT('ha2)
	) name15214 (
		\wishbone_tx_fifo_fifo_reg[0][5]/P0001 ,
		_w25385_,
		_w25386_,
		_w25727_
	);
	LUT4 #(
		.INIT('h135f)
	) name15215 (
		\wishbone_tx_fifo_fifo_reg[10][5]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][5]/P0001 ,
		_w25405_,
		_w25407_,
		_w25728_
	);
	LUT4 #(
		.INIT('h153f)
	) name15216 (
		\wishbone_tx_fifo_fifo_reg[12][5]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][5]/P0001 ,
		_w25404_,
		_w25408_,
		_w25729_
	);
	LUT4 #(
		.INIT('h153f)
	) name15217 (
		\wishbone_tx_fifo_fifo_reg[3][5]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][5]/P0001 ,
		_w25391_,
		_w25411_,
		_w25730_
	);
	LUT4 #(
		.INIT('h153f)
	) name15218 (
		\wishbone_tx_fifo_fifo_reg[5][5]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][5]/P0001 ,
		_w25393_,
		_w25396_,
		_w25731_
	);
	LUT4 #(
		.INIT('h8000)
	) name15219 (
		_w25728_,
		_w25729_,
		_w25730_,
		_w25731_,
		_w25732_
	);
	LUT2 #(
		.INIT('h8)
	) name15220 (
		\wishbone_tx_fifo_fifo_reg[15][5]/P0001 ,
		_w25399_,
		_w25733_
	);
	LUT4 #(
		.INIT('h135f)
	) name15221 (
		\wishbone_tx_fifo_fifo_reg[11][5]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][5]/P0001 ,
		_w25395_,
		_w25398_,
		_w25734_
	);
	LUT4 #(
		.INIT('h135f)
	) name15222 (
		\wishbone_tx_fifo_fifo_reg[13][5]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][5]/P0001 ,
		_w25388_,
		_w25410_,
		_w25735_
	);
	LUT4 #(
		.INIT('h135f)
	) name15223 (
		\wishbone_tx_fifo_fifo_reg[14][5]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[2][5]/P0001 ,
		_w25389_,
		_w25402_,
		_w25736_
	);
	LUT4 #(
		.INIT('h4000)
	) name15224 (
		_w25733_,
		_w25734_,
		_w25735_,
		_w25736_,
		_w25737_
	);
	LUT4 #(
		.INIT('hceee)
	) name15225 (
		_w25385_,
		_w25727_,
		_w25732_,
		_w25737_,
		_w25738_
	);
	LUT3 #(
		.INIT('ha2)
	) name15226 (
		\wishbone_tx_fifo_fifo_reg[0][6]/P0001 ,
		_w25385_,
		_w25386_,
		_w25739_
	);
	LUT4 #(
		.INIT('h153f)
	) name15227 (
		\wishbone_tx_fifo_fifo_reg[6][6]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][6]/P0001 ,
		_w25391_,
		_w25407_,
		_w25740_
	);
	LUT4 #(
		.INIT('h153f)
	) name15228 (
		\wishbone_tx_fifo_fifo_reg[1][6]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[2][6]/P0001 ,
		_w25402_,
		_w25410_,
		_w25741_
	);
	LUT4 #(
		.INIT('h153f)
	) name15229 (
		\wishbone_tx_fifo_fifo_reg[12][6]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][6]/P0001 ,
		_w25396_,
		_w25408_,
		_w25742_
	);
	LUT4 #(
		.INIT('h135f)
	) name15230 (
		\wishbone_tx_fifo_fifo_reg[14][6]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[3][6]/P0001 ,
		_w25389_,
		_w25411_,
		_w25743_
	);
	LUT4 #(
		.INIT('h8000)
	) name15231 (
		_w25740_,
		_w25741_,
		_w25742_,
		_w25743_,
		_w25744_
	);
	LUT2 #(
		.INIT('h8)
	) name15232 (
		\wishbone_tx_fifo_fifo_reg[7][6]/P0001 ,
		_w25393_,
		_w25745_
	);
	LUT4 #(
		.INIT('h153f)
	) name15233 (
		\wishbone_tx_fifo_fifo_reg[10][6]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][6]/P0001 ,
		_w25398_,
		_w25405_,
		_w25746_
	);
	LUT4 #(
		.INIT('h135f)
	) name15234 (
		\wishbone_tx_fifo_fifo_reg[11][6]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][6]/P0001 ,
		_w25395_,
		_w25404_,
		_w25747_
	);
	LUT4 #(
		.INIT('h135f)
	) name15235 (
		\wishbone_tx_fifo_fifo_reg[13][6]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[15][6]/P0001 ,
		_w25388_,
		_w25399_,
		_w25748_
	);
	LUT4 #(
		.INIT('h4000)
	) name15236 (
		_w25745_,
		_w25746_,
		_w25747_,
		_w25748_,
		_w25749_
	);
	LUT4 #(
		.INIT('hceee)
	) name15237 (
		_w25385_,
		_w25739_,
		_w25744_,
		_w25749_,
		_w25750_
	);
	LUT3 #(
		.INIT('ha2)
	) name15238 (
		\wishbone_tx_fifo_fifo_reg[0][7]/P0001 ,
		_w25385_,
		_w25386_,
		_w25751_
	);
	LUT4 #(
		.INIT('h153f)
	) name15239 (
		\wishbone_tx_fifo_fifo_reg[1][7]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][7]/P0001 ,
		_w25407_,
		_w25410_,
		_w25752_
	);
	LUT4 #(
		.INIT('h135f)
	) name15240 (
		\wishbone_tx_fifo_fifo_reg[11][7]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][7]/P0001 ,
		_w25395_,
		_w25404_,
		_w25753_
	);
	LUT4 #(
		.INIT('h135f)
	) name15241 (
		\wishbone_tx_fifo_fifo_reg[14][7]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][7]/P0001 ,
		_w25389_,
		_w25391_,
		_w25754_
	);
	LUT4 #(
		.INIT('h153f)
	) name15242 (
		\wishbone_tx_fifo_fifo_reg[10][7]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[15][7]/P0001 ,
		_w25399_,
		_w25405_,
		_w25755_
	);
	LUT4 #(
		.INIT('h8000)
	) name15243 (
		_w25752_,
		_w25753_,
		_w25754_,
		_w25755_,
		_w25756_
	);
	LUT2 #(
		.INIT('h8)
	) name15244 (
		\wishbone_tx_fifo_fifo_reg[3][7]/P0001 ,
		_w25411_,
		_w25757_
	);
	LUT4 #(
		.INIT('h153f)
	) name15245 (
		\wishbone_tx_fifo_fifo_reg[2][7]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][7]/P0001 ,
		_w25398_,
		_w25402_,
		_w25758_
	);
	LUT4 #(
		.INIT('h135f)
	) name15246 (
		\wishbone_tx_fifo_fifo_reg[13][7]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][7]/P0001 ,
		_w25388_,
		_w25396_,
		_w25759_
	);
	LUT4 #(
		.INIT('h153f)
	) name15247 (
		\wishbone_tx_fifo_fifo_reg[12][7]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][7]/P0001 ,
		_w25393_,
		_w25408_,
		_w25760_
	);
	LUT4 #(
		.INIT('h4000)
	) name15248 (
		_w25757_,
		_w25758_,
		_w25759_,
		_w25760_,
		_w25761_
	);
	LUT4 #(
		.INIT('hceee)
	) name15249 (
		_w25385_,
		_w25751_,
		_w25756_,
		_w25761_,
		_w25762_
	);
	LUT3 #(
		.INIT('ha2)
	) name15250 (
		\wishbone_tx_fifo_fifo_reg[0][8]/P0001 ,
		_w25385_,
		_w25386_,
		_w25763_
	);
	LUT4 #(
		.INIT('h135f)
	) name15251 (
		\wishbone_tx_fifo_fifo_reg[5][8]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][8]/P0001 ,
		_w25396_,
		_w25398_,
		_w25764_
	);
	LUT4 #(
		.INIT('h135f)
	) name15252 (
		\wishbone_tx_fifo_fifo_reg[13][8]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][8]/P0001 ,
		_w25388_,
		_w25404_,
		_w25765_
	);
	LUT4 #(
		.INIT('h153f)
	) name15253 (
		\wishbone_tx_fifo_fifo_reg[3][8]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][8]/P0001 ,
		_w25391_,
		_w25411_,
		_w25766_
	);
	LUT4 #(
		.INIT('h135f)
	) name15254 (
		\wishbone_tx_fifo_fifo_reg[15][8]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][8]/P0001 ,
		_w25399_,
		_w25407_,
		_w25767_
	);
	LUT4 #(
		.INIT('h8000)
	) name15255 (
		_w25764_,
		_w25765_,
		_w25766_,
		_w25767_,
		_w25768_
	);
	LUT2 #(
		.INIT('h8)
	) name15256 (
		\wishbone_tx_fifo_fifo_reg[11][8]/P0001 ,
		_w25395_,
		_w25769_
	);
	LUT4 #(
		.INIT('h135f)
	) name15257 (
		\wishbone_tx_fifo_fifo_reg[10][8]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[1][8]/P0001 ,
		_w25405_,
		_w25410_,
		_w25770_
	);
	LUT4 #(
		.INIT('h153f)
	) name15258 (
		\wishbone_tx_fifo_fifo_reg[12][8]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[14][8]/P0001 ,
		_w25389_,
		_w25408_,
		_w25771_
	);
	LUT4 #(
		.INIT('h153f)
	) name15259 (
		\wishbone_tx_fifo_fifo_reg[2][8]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[7][8]/P0001 ,
		_w25393_,
		_w25402_,
		_w25772_
	);
	LUT4 #(
		.INIT('h4000)
	) name15260 (
		_w25769_,
		_w25770_,
		_w25771_,
		_w25772_,
		_w25773_
	);
	LUT4 #(
		.INIT('hceee)
	) name15261 (
		_w25385_,
		_w25763_,
		_w25768_,
		_w25773_,
		_w25774_
	);
	LUT3 #(
		.INIT('ha2)
	) name15262 (
		\wishbone_tx_fifo_fifo_reg[0][9]/P0001 ,
		_w25385_,
		_w25386_,
		_w25775_
	);
	LUT4 #(
		.INIT('h135f)
	) name15263 (
		\wishbone_tx_fifo_fifo_reg[13][9]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[14][9]/P0001 ,
		_w25388_,
		_w25389_,
		_w25776_
	);
	LUT4 #(
		.INIT('h153f)
	) name15264 (
		\wishbone_tx_fifo_fifo_reg[7][9]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[9][9]/P0001 ,
		_w25391_,
		_w25393_,
		_w25777_
	);
	LUT4 #(
		.INIT('h135f)
	) name15265 (
		\wishbone_tx_fifo_fifo_reg[11][9]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[5][9]/P0001 ,
		_w25395_,
		_w25396_,
		_w25778_
	);
	LUT4 #(
		.INIT('h153f)
	) name15266 (
		\wishbone_tx_fifo_fifo_reg[15][9]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[8][9]/P0001 ,
		_w25398_,
		_w25399_,
		_w25779_
	);
	LUT4 #(
		.INIT('h8000)
	) name15267 (
		_w25776_,
		_w25777_,
		_w25778_,
		_w25779_,
		_w25780_
	);
	LUT2 #(
		.INIT('h8)
	) name15268 (
		\wishbone_tx_fifo_fifo_reg[2][9]/P0001 ,
		_w25402_,
		_w25781_
	);
	LUT4 #(
		.INIT('h153f)
	) name15269 (
		\wishbone_tx_fifo_fifo_reg[10][9]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[4][9]/P0001 ,
		_w25404_,
		_w25405_,
		_w25782_
	);
	LUT4 #(
		.INIT('h153f)
	) name15270 (
		\wishbone_tx_fifo_fifo_reg[12][9]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[6][9]/P0001 ,
		_w25407_,
		_w25408_,
		_w25783_
	);
	LUT4 #(
		.INIT('h135f)
	) name15271 (
		\wishbone_tx_fifo_fifo_reg[1][9]/P0001 ,
		\wishbone_tx_fifo_fifo_reg[3][9]/P0001 ,
		_w25410_,
		_w25411_,
		_w25784_
	);
	LUT4 #(
		.INIT('h4000)
	) name15272 (
		_w25781_,
		_w25782_,
		_w25783_,
		_w25784_,
		_w25785_
	);
	LUT4 #(
		.INIT('hceee)
	) name15273 (
		_w25385_,
		_w25775_,
		_w25780_,
		_w25785_,
		_w25786_
	);
	LUT3 #(
		.INIT('ha8)
	) name15274 (
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		_w11882_,
		_w11884_,
		_w25787_
	);
	LUT2 #(
		.INIT('h6)
	) name15275 (
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		_w25788_
	);
	LUT4 #(
		.INIT('h8f00)
	) name15276 (
		_w11866_,
		_w11867_,
		_w11883_,
		_w25788_,
		_w25789_
	);
	LUT2 #(
		.INIT('h4)
	) name15277 (
		_w11882_,
		_w25789_,
		_w25790_
	);
	LUT3 #(
		.INIT('hf8)
	) name15278 (
		_w24535_,
		_w25787_,
		_w25790_,
		_w25791_
	);
	LUT2 #(
		.INIT('h2)
	) name15279 (
		\wishbone_ReadTxDataFromFifo_sync2_reg/NET0131 ,
		\wishbone_ReadTxDataFromFifo_sync3_reg/NET0131 ,
		_w25792_
	);
	LUT4 #(
		.INIT('h8808)
	) name15280 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_ReadTxDataFromFifo_sync2_reg/NET0131 ,
		\wishbone_ReadTxDataFromFifo_sync3_reg/NET0131 ,
		_w25793_
	);
	LUT2 #(
		.INIT('h1)
	) name15281 (
		\wishbone_tx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[1]/NET0131 ,
		_w25794_
	);
	LUT3 #(
		.INIT('h01)
	) name15282 (
		\wishbone_tx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[1]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[2]/NET0131 ,
		_w25795_
	);
	LUT2 #(
		.INIT('h1)
	) name15283 (
		\wishbone_tx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25796_
	);
	LUT4 #(
		.INIT('h0008)
	) name15284 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25797_
	);
	LUT4 #(
		.INIT('h0070)
	) name15285 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_ReadTxDataFromFifo_sync2_reg/NET0131 ,
		\wishbone_ReadTxDataFromFifo_sync3_reg/NET0131 ,
		_w25798_
	);
	LUT4 #(
		.INIT('h5999)
	) name15286 (
		_w12304_,
		_w25792_,
		_w25795_,
		_w25796_,
		_w25799_
	);
	LUT2 #(
		.INIT('h8)
	) name15287 (
		\wishbone_tx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[1]/NET0131 ,
		_w25800_
	);
	LUT4 #(
		.INIT('h8000)
	) name15288 (
		\wishbone_tx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[1]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[2]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[3]/NET0131 ,
		_w25801_
	);
	LUT4 #(
		.INIT('h0001)
	) name15289 (
		\wishbone_tx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[1]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[2]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[3]/NET0131 ,
		_w25802_
	);
	LUT4 #(
		.INIT('hf531)
	) name15290 (
		_w12304_,
		_w25792_,
		_w25801_,
		_w25802_,
		_w25803_
	);
	LUT4 #(
		.INIT('h8488)
	) name15291 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25385_,
		_w25799_,
		_w25803_,
		_w25804_
	);
	LUT3 #(
		.INIT('h1b)
	) name15292 (
		\ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131 ,
		\wishbone_RxStatusWriteLatched_sync2_reg/NET0131 ,
		_w25805_
	);
	LUT4 #(
		.INIT('hea00)
	) name15293 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131 ,
		_w11921_,
		_w24778_,
		_w25805_,
		_w25806_
	);
	LUT2 #(
		.INIT('h4)
	) name15294 (
		mdc_pad_o_pad,
		\miim1_InProgress_reg/NET0131 ,
		_w25807_
	);
	LUT3 #(
		.INIT('h80)
	) name15295 (
		_w24411_,
		_w24420_,
		_w25807_,
		_w25808_
	);
	LUT4 #(
		.INIT('h8000)
	) name15296 (
		\miim1_BitCounter_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[1]/NET0131 ,
		\miim1_BitCounter_reg[2]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w25809_
	);
	LUT3 #(
		.INIT('h6c)
	) name15297 (
		\miim1_BitCounter_reg[4]/NET0131 ,
		\miim1_BitCounter_reg[5]/NET0131 ,
		_w25809_,
		_w25810_
	);
	LUT2 #(
		.INIT('h8)
	) name15298 (
		_w25808_,
		_w25810_,
		_w25811_
	);
	LUT3 #(
		.INIT('h40)
	) name15299 (
		mdc_pad_o_pad,
		_w24411_,
		_w24420_,
		_w25812_
	);
	LUT3 #(
		.INIT('h35)
	) name15300 (
		\miim1_BitCounter_reg[5]/NET0131 ,
		_w24567_,
		_w25812_,
		_w25813_
	);
	LUT2 #(
		.INIT('hb)
	) name15301 (
		_w25811_,
		_w25813_,
		_w25814_
	);
	LUT4 #(
		.INIT('haa2a)
	) name15302 (
		\wishbone_rx_burst_en_reg/NET0131 ,
		_w11870_,
		_w11873_,
		_w11876_,
		_w25815_
	);
	LUT2 #(
		.INIT('h8)
	) name15303 (
		_w24515_,
		_w25815_,
		_w25816_
	);
	LUT3 #(
		.INIT('h08)
	) name15304 (
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w25817_
	);
	LUT3 #(
		.INIT('h07)
	) name15305 (
		_w11868_,
		_w11875_,
		_w25817_,
		_w25818_
	);
	LUT3 #(
		.INIT('h80)
	) name15306 (
		_w11870_,
		_w11873_,
		_w25818_,
		_w25819_
	);
	LUT4 #(
		.INIT('hfd00)
	) name15307 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[1]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[2]/NET0131 ,
		_w25820_
	);
	LUT2 #(
		.INIT('h2)
	) name15308 (
		_w11867_,
		_w25820_,
		_w25821_
	);
	LUT2 #(
		.INIT('h2)
	) name15309 (
		_w24505_,
		_w25821_,
		_w25822_
	);
	LUT4 #(
		.INIT('h8f03)
	) name15310 (
		_w11866_,
		_w11867_,
		_w24510_,
		_w25820_,
		_w25823_
	);
	LUT3 #(
		.INIT('h40)
	) name15311 (
		_w24504_,
		_w24513_,
		_w25823_,
		_w25824_
	);
	LUT3 #(
		.INIT('h01)
	) name15312 (
		_w25819_,
		_w25822_,
		_w25824_,
		_w25825_
	);
	LUT2 #(
		.INIT('hb)
	) name15313 (
		_w25816_,
		_w25825_,
		_w25826_
	);
	LUT2 #(
		.INIT('h2)
	) name15314 (
		\wishbone_WriteRxDataToFifoSync2_reg/NET0131 ,
		\wishbone_WriteRxDataToFifoSync3_reg/NET0131 ,
		_w25827_
	);
	LUT4 #(
		.INIT('h8808)
	) name15315 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_WriteRxDataToFifoSync2_reg/NET0131 ,
		\wishbone_WriteRxDataToFifoSync3_reg/NET0131 ,
		_w25828_
	);
	LUT2 #(
		.INIT('h4)
	) name15316 (
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[4]/NET0131 ,
		_w25829_
	);
	LUT4 #(
		.INIT('h0800)
	) name15317 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[4]/NET0131 ,
		_w25830_
	);
	LUT4 #(
		.INIT('h0070)
	) name15318 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_WriteRxDataToFifoSync2_reg/NET0131 ,
		\wishbone_WriteRxDataToFifoSync3_reg/NET0131 ,
		_w25831_
	);
	LUT4 #(
		.INIT('h63c3)
	) name15319 (
		_w11866_,
		_w13809_,
		_w25827_,
		_w25829_,
		_w25832_
	);
	LUT3 #(
		.INIT('h15)
	) name15320 (
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		_w11866_,
		_w13809_,
		_w25833_
	);
	LUT2 #(
		.INIT('h8)
	) name15321 (
		\wishbone_rx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[1]/NET0131 ,
		_w25834_
	);
	LUT3 #(
		.INIT('h70)
	) name15322 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[2]/NET0131 ,
		_w25835_
	);
	LUT3 #(
		.INIT('h2a)
	) name15323 (
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		_w25834_,
		_w25835_,
		_w25836_
	);
	LUT3 #(
		.INIT('hb0)
	) name15324 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[4]/NET0131 ,
		_w25837_
	);
	LUT4 #(
		.INIT('hfe00)
	) name15325 (
		_w25832_,
		_w25833_,
		_w25836_,
		_w25837_,
		_w25838_
	);
	LUT3 #(
		.INIT('h0b)
	) name15326 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[4]/NET0131 ,
		_w25839_
	);
	LUT4 #(
		.INIT('h0100)
	) name15327 (
		_w25832_,
		_w25833_,
		_w25836_,
		_w25839_,
		_w25840_
	);
	LUT2 #(
		.INIT('he)
	) name15328 (
		_w25838_,
		_w25840_,
		_w25841_
	);
	LUT4 #(
		.INIT('h0200)
	) name15329 (
		\maccontrol1_receivecontrol1_DlyCrcCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131 ,
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w25842_
	);
	LUT3 #(
		.INIT('h2a)
	) name15330 (
		\maccontrol1_receivecontrol1_DlyCrcCnt_reg[1]/NET0131 ,
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w25843_
	);
	LUT3 #(
		.INIT('h12)
	) name15331 (
		\maccontrol1_receivecontrol1_DlyCrcCnt_reg[1]/NET0131 ,
		_w24524_,
		_w25842_,
		_w25844_
	);
	LUT4 #(
		.INIT('h09aa)
	) name15332 (
		\maccontrol1_receivecontrol1_DlyCrcCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131 ,
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w25845_
	);
	LUT3 #(
		.INIT('h2a)
	) name15333 (
		\maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131 ,
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w25846_
	);
	LUT3 #(
		.INIT('hf8)
	) name15334 (
		_w25842_,
		_w25843_,
		_w25846_,
		_w25847_
	);
	LUT3 #(
		.INIT('h10)
	) name15335 (
		\txethmac1_txcrc_Crc_reg[28]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w25848_
	);
	LUT3 #(
		.INIT('h10)
	) name15336 (
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w25849_
	);
	LUT3 #(
		.INIT('h10)
	) name15337 (
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w25850_
	);
	LUT4 #(
		.INIT('h0103)
	) name15338 (
		_w10801_,
		_w25848_,
		_w25849_,
		_w25850_,
		_w25851_
	);
	LUT3 #(
		.INIT('h37)
	) name15339 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		_w10999_,
		_w25851_,
		_w25852_
	);
	LUT4 #(
		.INIT('h1000)
	) name15340 (
		\txethmac1_txcrc_Crc_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11787_,
		_w11790_,
		_w25853_
	);
	LUT3 #(
		.INIT('h40)
	) name15341 (
		\txethmac1_txcrc_Crc_reg[1]/NET0131 ,
		_w10913_,
		_w10914_,
		_w25854_
	);
	LUT3 #(
		.INIT('hab)
	) name15342 (
		_w25853_,
		_w25854_,
		_w11793_,
		_w25855_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name15343 (
		\wishbone_LastByteIn_reg/NET0131 ,
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		\wishbone_RxByteCnt_reg[1]/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w25856_
	);
	LUT3 #(
		.INIT('h2a)
	) name15344 (
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		\wishbone_RxByteCnt_reg[1]/NET0131 ,
		_w25857_
	);
	LUT4 #(
		.INIT('h5450)
	) name15345 (
		\RxAbort_wb_reg/NET0131 ,
		_w24427_,
		_w25856_,
		_w25857_,
		_w25858_
	);
	LUT2 #(
		.INIT('h8)
	) name15346 (
		\rxethmac1_LatchedByte_reg[4]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w25859_
	);
	LUT3 #(
		.INIT('h70)
	) name15347 (
		_w10519_,
		_w24852_,
		_w25859_,
		_w25860_
	);
	LUT2 #(
		.INIT('h8)
	) name15348 (
		\rxethmac1_DelayData_reg/NET0131 ,
		\rxethmac1_RxData_d_reg[4]/NET0131 ,
		_w25861_
	);
	LUT4 #(
		.INIT('hd500)
	) name15349 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10519_,
		_w24852_,
		_w25861_,
		_w25862_
	);
	LUT2 #(
		.INIT('he)
	) name15350 (
		_w25860_,
		_w25862_,
		_w25863_
	);
	LUT3 #(
		.INIT('h08)
	) name15351 (
		\miim1_BitCounter_reg[4]/NET0131 ,
		\miim1_BitCounter_reg[5]/NET0131 ,
		\miim1_BitCounter_reg[6]/NET0131 ,
		_w25864_
	);
	LUT2 #(
		.INIT('h8)
	) name15352 (
		_w25809_,
		_w25864_,
		_w25865_
	);
	LUT4 #(
		.INIT('h0100)
	) name15353 (
		\miim1_InProgress_q1_reg/NET0131 ,
		\miim1_InProgress_q2_reg/NET0131 ,
		\miim1_InProgress_reg/NET0131 ,
		\miim1_SyncStatMdcEn_reg/NET0131 ,
		_w25866_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name15354 (
		\miim1_RStatStart_q1_reg/NET0131 ,
		\miim1_RStatStart_q2_reg/NET0131 ,
		\miim1_WCtrlDataStart_q1_reg/NET0131 ,
		\miim1_WCtrlDataStart_q2_reg/NET0131 ,
		_w25867_
	);
	LUT2 #(
		.INIT('h4)
	) name15355 (
		_w25866_,
		_w25867_,
		_w25868_
	);
	LUT4 #(
		.INIT('h0700)
	) name15356 (
		_w25809_,
		_w25864_,
		_w25866_,
		_w25867_,
		_w25869_
	);
	LUT2 #(
		.INIT('h2)
	) name15357 (
		\miim1_InProgress_reg/NET0131 ,
		\miim1_WriteOp_reg/NET0131 ,
		_w25870_
	);
	LUT4 #(
		.INIT('hae04)
	) name15358 (
		\miim1_InProgress_reg/NET0131 ,
		\miim1_WCtrlDataStart_q1_reg/NET0131 ,
		\miim1_WCtrlDataStart_q2_reg/NET0131 ,
		\miim1_WriteOp_reg/NET0131 ,
		_w25871_
	);
	LUT3 #(
		.INIT('hb0)
	) name15359 (
		_w25866_,
		_w25867_,
		_w25871_,
		_w25872_
	);
	LUT4 #(
		.INIT('heea2)
	) name15360 (
		\miim1_WriteOp_reg/NET0131 ,
		_w25812_,
		_w25869_,
		_w25872_,
		_w25873_
	);
	LUT2 #(
		.INIT('h2)
	) name15361 (
		\ethreg1_MODER_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131 ,
		_w25874_
	);
	LUT3 #(
		.INIT('h02)
	) name15362 (
		\ethreg1_MODER_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131 ,
		\wishbone_r_RxEn_q_reg/NET0131 ,
		_w25875_
	);
	LUT4 #(
		.INIT('h8000)
	) name15363 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxStatus_reg[13]/NET0131 ,
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w25876_
	);
	LUT2 #(
		.INIT('h1)
	) name15364 (
		_w25875_,
		_w25876_,
		_w25877_
	);
	LUT3 #(
		.INIT('ha8)
	) name15365 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[3]/NET0131 ,
		_w25875_,
		_w25876_,
		_w25878_
	);
	LUT3 #(
		.INIT('h80)
	) name15366 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w25879_
	);
	LUT3 #(
		.INIT('h80)
	) name15367 (
		\wishbone_RxBDAddress_reg[1]/NET0131 ,
		\wishbone_RxBDAddress_reg[2]/NET0131 ,
		\wishbone_RxBDAddress_reg[3]/NET0131 ,
		_w25880_
	);
	LUT3 #(
		.INIT('h15)
	) name15368 (
		\wishbone_RxBDAddress_reg[4]/NET0131 ,
		_w25879_,
		_w25880_,
		_w25881_
	);
	LUT4 #(
		.INIT('h8000)
	) name15369 (
		\wishbone_RxBDAddress_reg[4]/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w25882_
	);
	LUT2 #(
		.INIT('h8)
	) name15370 (
		_w25880_,
		_w25882_,
		_w25883_
	);
	LUT4 #(
		.INIT('h0111)
	) name15371 (
		_w25875_,
		_w25876_,
		_w25880_,
		_w25882_,
		_w25884_
	);
	LUT3 #(
		.INIT('hba)
	) name15372 (
		_w25878_,
		_w25881_,
		_w25884_,
		_w25885_
	);
	LUT2 #(
		.INIT('h1)
	) name15373 (
		\wishbone_LastByteIn_reg/NET0131 ,
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w25886_
	);
	LUT4 #(
		.INIT('h80aa)
	) name15374 (
		_w24429_,
		_w24524_,
		_w24525_,
		_w25886_,
		_w25887_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name15375 (
		mdc_pad_o_pad,
		\miim1_BitCounter_reg[1]/NET0131 ,
		_w24411_,
		_w24420_,
		_w25888_
	);
	LUT2 #(
		.INIT('h6)
	) name15376 (
		\miim1_BitCounter_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[1]/NET0131 ,
		_w25889_
	);
	LUT3 #(
		.INIT('h70)
	) name15377 (
		_w24564_,
		_w24565_,
		_w25889_,
		_w25890_
	);
	LUT3 #(
		.INIT('hec)
	) name15378 (
		_w25808_,
		_w25888_,
		_w25890_,
		_w25891_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name15379 (
		mdc_pad_o_pad,
		\miim1_BitCounter_reg[2]/NET0131 ,
		_w24411_,
		_w24420_,
		_w25892_
	);
	LUT3 #(
		.INIT('h78)
	) name15380 (
		\miim1_BitCounter_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[1]/NET0131 ,
		\miim1_BitCounter_reg[2]/NET0131 ,
		_w25893_
	);
	LUT3 #(
		.INIT('h70)
	) name15381 (
		_w24564_,
		_w24565_,
		_w25893_,
		_w25894_
	);
	LUT3 #(
		.INIT('hec)
	) name15382 (
		_w25808_,
		_w25892_,
		_w25894_,
		_w25895_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name15383 (
		mdc_pad_o_pad,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w24411_,
		_w24420_,
		_w25896_
	);
	LUT4 #(
		.INIT('h7f80)
	) name15384 (
		\miim1_BitCounter_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[1]/NET0131 ,
		\miim1_BitCounter_reg[2]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w25897_
	);
	LUT4 #(
		.INIT('hf4f0)
	) name15385 (
		_w24566_,
		_w25808_,
		_w25896_,
		_w25897_,
		_w25898_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name15386 (
		mdc_pad_o_pad,
		\miim1_BitCounter_reg[4]/NET0131 ,
		_w24411_,
		_w24420_,
		_w25899_
	);
	LUT2 #(
		.INIT('h6)
	) name15387 (
		\miim1_BitCounter_reg[4]/NET0131 ,
		_w25809_,
		_w25900_
	);
	LUT4 #(
		.INIT('hf4f0)
	) name15388 (
		_w24566_,
		_w25808_,
		_w25899_,
		_w25900_,
		_w25901_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name15389 (
		mdc_pad_o_pad,
		\miim1_BitCounter_reg[6]/NET0131 ,
		_w24411_,
		_w24420_,
		_w25902_
	);
	LUT4 #(
		.INIT('h870f)
	) name15390 (
		\miim1_BitCounter_reg[4]/NET0131 ,
		\miim1_BitCounter_reg[5]/NET0131 ,
		\miim1_BitCounter_reg[6]/NET0131 ,
		_w25809_,
		_w25903_
	);
	LUT4 #(
		.INIT('hf0f4)
	) name15391 (
		_w24566_,
		_w25808_,
		_w25902_,
		_w25903_,
		_w25904_
	);
	LUT2 #(
		.INIT('h1)
	) name15392 (
		\miim1_clkgen_Counter_reg[4]/NET0131 ,
		\miim1_clkgen_Counter_reg[5]/NET0131 ,
		_w25905_
	);
	LUT3 #(
		.INIT('h2a)
	) name15393 (
		\miim1_clkgen_Counter_reg[6]/NET0131 ,
		_w24411_,
		_w25905_,
		_w25906_
	);
	LUT3 #(
		.INIT('h01)
	) name15394 (
		\ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131 ,
		_w25907_
	);
	LUT3 #(
		.INIT('h40)
	) name15395 (
		_w24415_,
		_w24416_,
		_w25907_,
		_w25908_
	);
	LUT4 #(
		.INIT('hf4f8)
	) name15396 (
		\ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131 ,
		_w24421_,
		_w25906_,
		_w25908_,
		_w25909_
	);
	LUT3 #(
		.INIT('h02)
	) name15397 (
		\rxethmac1_Multicast_reg/NET0131 ,
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		\rxethmac1_rxaddrcheck1_RxAbort_reg/NET0131 ,
		_w25910_
	);
	LUT2 #(
		.INIT('h8)
	) name15398 (
		\rxethmac1_LatchedByte_reg[0]/NET0131 ,
		_w11800_,
		_w25911_
	);
	LUT3 #(
		.INIT('hec)
	) name15399 (
		_w11797_,
		_w25910_,
		_w25911_,
		_w25912_
	);
	LUT2 #(
		.INIT('h1)
	) name15400 (
		\maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w25913_
	);
	LUT3 #(
		.INIT('h07)
	) name15401 (
		_w24444_,
		_w24445_,
		_w25913_,
		_w25914_
	);
	LUT2 #(
		.INIT('h4)
	) name15402 (
		\rxethmac1_crcrx_Crc_reg[13]/NET0131 ,
		_w10582_,
		_w25915_
	);
	LUT4 #(
		.INIT('h8f00)
	) name15403 (
		_w10554_,
		_w10573_,
		_w10581_,
		_w25915_,
		_w25916_
	);
	LUT2 #(
		.INIT('h8)
	) name15404 (
		\rxethmac1_crcrx_Crc_reg[13]/NET0131 ,
		_w10582_,
		_w25917_
	);
	LUT4 #(
		.INIT('h7000)
	) name15405 (
		_w10554_,
		_w10573_,
		_w10581_,
		_w25917_,
		_w25918_
	);
	LUT2 #(
		.INIT('h1)
	) name15406 (
		_w25916_,
		_w25918_,
		_w25919_
	);
	LUT3 #(
		.INIT('h0b)
	) name15407 (
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_q_reg/P0001 ,
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w25920_
	);
	LUT2 #(
		.INIT('h8)
	) name15408 (
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[1]/NET0131 ,
		_w25921_
	);
	LUT3 #(
		.INIT('h2a)
	) name15409 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[1]/NET0131 ,
		_w25922_
	);
	LUT4 #(
		.INIT('hc444)
	) name15410 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[1]/NET0131 ,
		_w25923_
	);
	LUT2 #(
		.INIT('h4)
	) name15411 (
		_w25920_,
		_w25923_,
		_w25924_
	);
	LUT3 #(
		.INIT('h04)
	) name15412 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w25925_
	);
	LUT4 #(
		.INIT('h1000)
	) name15413 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w25926_
	);
	LUT3 #(
		.INIT('h2a)
	) name15414 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		_w25925_,
		_w25926_,
		_w25927_
	);
	LUT4 #(
		.INIT('h2000)
	) name15415 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_q_reg/P0001 ,
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w25928_
	);
	LUT2 #(
		.INIT('h4)
	) name15416 (
		_w25922_,
		_w25928_,
		_w25929_
	);
	LUT2 #(
		.INIT('h8)
	) name15417 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w25930_
	);
	LUT4 #(
		.INIT('hf800)
	) name15418 (
		_w25924_,
		_w25927_,
		_w25929_,
		_w25930_,
		_w25931_
	);
	LUT2 #(
		.INIT('h1)
	) name15419 (
		\txethmac1_TxAbort_reg/NET0131 ,
		\txethmac1_TxDone_reg/NET0131 ,
		_w25932_
	);
	LUT4 #(
		.INIT('h00ab)
	) name15420 (
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		\txethmac1_TxAbort_reg/NET0131 ,
		\txethmac1_TxDone_reg/NET0131 ,
		wb_rst_i_pad,
		_w25933_
	);
	LUT3 #(
		.INIT('h80)
	) name15421 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		_w25934_
	);
	LUT4 #(
		.INIT('hf800)
	) name15422 (
		_w25924_,
		_w25927_,
		_w25929_,
		_w25934_,
		_w25935_
	);
	LUT4 #(
		.INIT('h00e0)
	) name15423 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		_w25931_,
		_w25933_,
		_w25935_,
		_w25936_
	);
	LUT3 #(
		.INIT('h40)
	) name15424 (
		\wishbone_LatchValidBytes_q_reg/NET0131 ,
		\wishbone_LatchValidBytes_reg/NET0131 ,
		\wishbone_TxLength_reg[0]/NET0131 ,
		_w25937_
	);
	LUT3 #(
		.INIT('h80)
	) name15425 (
		_w12314_,
		_w12316_,
		_w25937_,
		_w25938_
	);
	LUT2 #(
		.INIT('h4)
	) name15426 (
		\wishbone_TxAbort_wb_q_reg/NET0131 ,
		\wishbone_TxAbort_wb_reg/NET0131 ,
		_w25939_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name15427 (
		\wishbone_TxAbort_wb_q_reg/NET0131 ,
		\wishbone_TxAbort_wb_reg/NET0131 ,
		\wishbone_TxRetry_wb_q_reg/NET0131 ,
		\wishbone_TxRetry_wb_reg/NET0131 ,
		_w25940_
	);
	LUT2 #(
		.INIT('h4)
	) name15428 (
		\wishbone_TxDone_wb_q_reg/NET0131 ,
		\wishbone_TxDone_wb_reg/NET0131 ,
		_w25941_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name15429 (
		\wishbone_LatchValidBytes_q_reg/NET0131 ,
		\wishbone_LatchValidBytes_reg/NET0131 ,
		\wishbone_TxDone_wb_q_reg/NET0131 ,
		\wishbone_TxDone_wb_reg/NET0131 ,
		_w25942_
	);
	LUT3 #(
		.INIT('h80)
	) name15430 (
		\wishbone_TxValidBytesLatched_reg[0]/NET0131 ,
		_w25940_,
		_w25942_,
		_w25943_
	);
	LUT3 #(
		.INIT('hf8)
	) name15431 (
		_w12312_,
		_w25938_,
		_w25943_,
		_w25944_
	);
	LUT3 #(
		.INIT('h40)
	) name15432 (
		\wishbone_LatchValidBytes_q_reg/NET0131 ,
		\wishbone_LatchValidBytes_reg/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		_w25945_
	);
	LUT3 #(
		.INIT('h80)
	) name15433 (
		_w12314_,
		_w12316_,
		_w25945_,
		_w25946_
	);
	LUT3 #(
		.INIT('h80)
	) name15434 (
		\wishbone_TxValidBytesLatched_reg[1]/NET0131 ,
		_w25940_,
		_w25942_,
		_w25947_
	);
	LUT3 #(
		.INIT('hf8)
	) name15435 (
		_w12312_,
		_w25946_,
		_w25947_,
		_w25948_
	);
	LUT2 #(
		.INIT('h7)
	) name15436 (
		_w11007_,
		_w11569_,
		_w25949_
	);
	LUT2 #(
		.INIT('h7)
	) name15437 (
		_w11007_,
		_w11631_,
		_w25950_
	);
	LUT3 #(
		.INIT('h10)
	) name15438 (
		mdc_pad_o_pad,
		\miim1_BitCounter_reg[0]/NET0131 ,
		\miim1_InProgress_reg/NET0131 ,
		_w25951_
	);
	LUT3 #(
		.INIT('h80)
	) name15439 (
		_w24411_,
		_w24420_,
		_w25951_,
		_w25952_
	);
	LUT4 #(
		.INIT('hffca)
	) name15440 (
		\miim1_BitCounter_reg[0]/NET0131 ,
		_w24567_,
		_w25812_,
		_w25952_,
		_w25953_
	);
	LUT4 #(
		.INIT('h2070)
	) name15441 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_TxCtrlEndFrm_reg/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\wishbone_TxEndFrm_reg/NET0131 ,
		_w25954_
	);
	LUT4 #(
		.INIT('h3320)
	) name15442 (
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w10604_,
		_w10801_,
		_w25954_,
		_w25955_
	);
	LUT4 #(
		.INIT('h4445)
	) name15443 (
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w10779_,
		_w10936_,
		_w10937_,
		_w25956_
	);
	LUT3 #(
		.INIT('h01)
	) name15444 (
		_w10830_,
		_w25955_,
		_w25956_,
		_w25957_
	);
	LUT4 #(
		.INIT('h2aee)
	) name15445 (
		\miim1_InProgress_reg/NET0131 ,
		_w25812_,
		_w25865_,
		_w25868_,
		_w25958_
	);
	LUT3 #(
		.INIT('h1f)
	) name15446 (
		\ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131 ,
		_w25959_
	);
	LUT4 #(
		.INIT('h8a00)
	) name15447 (
		_w24411_,
		_w24415_,
		_w24416_,
		_w24420_,
		_w25960_
	);
	LUT3 #(
		.INIT('h1e)
	) name15448 (
		\miim1_clkgen_Counter_reg[0]/NET0131 ,
		\miim1_clkgen_Counter_reg[1]/NET0131 ,
		\miim1_clkgen_Counter_reg[2]/NET0131 ,
		_w25961_
	);
	LUT3 #(
		.INIT('h70)
	) name15449 (
		_w24411_,
		_w24420_,
		_w25961_,
		_w25962_
	);
	LUT3 #(
		.INIT('h07)
	) name15450 (
		_w25959_,
		_w25960_,
		_w25962_,
		_w25963_
	);
	LUT3 #(
		.INIT('h20)
	) name15451 (
		\miim1_BitCounter_reg[4]/NET0131 ,
		\miim1_BitCounter_reg[6]/NET0131 ,
		\miim1_InProgress_reg/NET0131 ,
		_w25964_
	);
	LUT2 #(
		.INIT('h8)
	) name15452 (
		\miim1_BitCounter_reg[1]/NET0131 ,
		\miim1_BitCounter_reg[2]/NET0131 ,
		_w25965_
	);
	LUT4 #(
		.INIT('h0020)
	) name15453 (
		\miim1_BitCounter_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		\miim1_BitCounter_reg[5]/NET0131 ,
		\miim1_WriteOp_reg/NET0131 ,
		_w25966_
	);
	LUT3 #(
		.INIT('h80)
	) name15454 (
		_w25964_,
		_w25965_,
		_w25966_,
		_w25967_
	);
	LUT3 #(
		.INIT('he2)
	) name15455 (
		\miim1_LatchByte1_d_reg/NET0131 ,
		_w25812_,
		_w25967_,
		_w25968_
	);
	LUT3 #(
		.INIT('h80)
	) name15456 (
		\wishbone_RxBDAddress_reg[4]/NET0131 ,
		\wishbone_RxBDAddress_reg[5]/NET0131 ,
		\wishbone_RxBDAddress_reg[6]/NET0131 ,
		_w25969_
	);
	LUT4 #(
		.INIT('h1555)
	) name15457 (
		\wishbone_RxBDAddress_reg[7]/NET0131 ,
		_w25879_,
		_w25880_,
		_w25969_,
		_w25970_
	);
	LUT4 #(
		.INIT('h8000)
	) name15458 (
		\wishbone_RxBDAddress_reg[4]/NET0131 ,
		\wishbone_RxBDAddress_reg[5]/NET0131 ,
		\wishbone_RxBDAddress_reg[6]/NET0131 ,
		\wishbone_RxBDAddress_reg[7]/NET0131 ,
		_w25971_
	);
	LUT3 #(
		.INIT('h80)
	) name15459 (
		_w25879_,
		_w25880_,
		_w25971_,
		_w25972_
	);
	LUT4 #(
		.INIT('h222e)
	) name15460 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[6]/NET0131 ,
		_w25877_,
		_w25970_,
		_w25972_,
		_w25973_
	);
	LUT3 #(
		.INIT('h20)
	) name15461 (
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_LastByteIn_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w25974_
	);
	LUT3 #(
		.INIT('h20)
	) name15462 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w25975_
	);
	LUT4 #(
		.INIT('h1000)
	) name15463 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		\wishbone_RxByteCnt_reg[1]/NET0131 ,
		\wishbone_RxEnableWindow_reg/NET0131 ,
		_w25976_
	);
	LUT4 #(
		.INIT('h1115)
	) name15464 (
		\wishbone_RxDataLatched1_reg[10]/NET0131 ,
		_w25974_,
		_w25975_,
		_w25976_,
		_w25977_
	);
	LUT4 #(
		.INIT('h0400)
	) name15465 (
		\rxethmac1_RxData_reg[2]/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_LastByteIn_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w25978_
	);
	LUT3 #(
		.INIT('he0)
	) name15466 (
		_w25975_,
		_w25976_,
		_w25978_,
		_w25979_
	);
	LUT2 #(
		.INIT('h1)
	) name15467 (
		_w25977_,
		_w25979_,
		_w25980_
	);
	LUT4 #(
		.INIT('h1115)
	) name15468 (
		\wishbone_RxDataLatched1_reg[11]/NET0131 ,
		_w25974_,
		_w25975_,
		_w25976_,
		_w25981_
	);
	LUT4 #(
		.INIT('h0400)
	) name15469 (
		\rxethmac1_RxData_reg[3]/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_LastByteIn_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w25982_
	);
	LUT3 #(
		.INIT('he0)
	) name15470 (
		_w25975_,
		_w25976_,
		_w25982_,
		_w25983_
	);
	LUT2 #(
		.INIT('h1)
	) name15471 (
		_w25981_,
		_w25983_,
		_w25984_
	);
	LUT4 #(
		.INIT('h1115)
	) name15472 (
		\wishbone_RxDataLatched1_reg[12]/NET0131 ,
		_w25974_,
		_w25975_,
		_w25976_,
		_w25985_
	);
	LUT4 #(
		.INIT('h0400)
	) name15473 (
		\rxethmac1_RxData_reg[4]/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_LastByteIn_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w25986_
	);
	LUT3 #(
		.INIT('he0)
	) name15474 (
		_w25975_,
		_w25976_,
		_w25986_,
		_w25987_
	);
	LUT2 #(
		.INIT('h1)
	) name15475 (
		_w25985_,
		_w25987_,
		_w25988_
	);
	LUT4 #(
		.INIT('h1115)
	) name15476 (
		\wishbone_RxDataLatched1_reg[13]/NET0131 ,
		_w25974_,
		_w25975_,
		_w25976_,
		_w25989_
	);
	LUT4 #(
		.INIT('h0400)
	) name15477 (
		\rxethmac1_RxData_reg[5]/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_LastByteIn_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w25990_
	);
	LUT3 #(
		.INIT('he0)
	) name15478 (
		_w25975_,
		_w25976_,
		_w25990_,
		_w25991_
	);
	LUT2 #(
		.INIT('h1)
	) name15479 (
		_w25989_,
		_w25991_,
		_w25992_
	);
	LUT4 #(
		.INIT('h1115)
	) name15480 (
		\wishbone_RxDataLatched1_reg[14]/NET0131 ,
		_w25974_,
		_w25975_,
		_w25976_,
		_w25993_
	);
	LUT4 #(
		.INIT('h0400)
	) name15481 (
		\rxethmac1_RxData_reg[6]/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_LastByteIn_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w25994_
	);
	LUT3 #(
		.INIT('he0)
	) name15482 (
		_w25975_,
		_w25976_,
		_w25994_,
		_w25995_
	);
	LUT2 #(
		.INIT('h1)
	) name15483 (
		_w25993_,
		_w25995_,
		_w25996_
	);
	LUT4 #(
		.INIT('h1115)
	) name15484 (
		\wishbone_RxDataLatched1_reg[15]/NET0131 ,
		_w25974_,
		_w25975_,
		_w25976_,
		_w25997_
	);
	LUT4 #(
		.INIT('h0400)
	) name15485 (
		\rxethmac1_RxData_reg[7]/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_LastByteIn_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w25998_
	);
	LUT3 #(
		.INIT('he0)
	) name15486 (
		_w25975_,
		_w25976_,
		_w25998_,
		_w25999_
	);
	LUT2 #(
		.INIT('h1)
	) name15487 (
		_w25997_,
		_w25999_,
		_w26000_
	);
	LUT3 #(
		.INIT('h08)
	) name15488 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w26001_
	);
	LUT4 #(
		.INIT('h0400)
	) name15489 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		\wishbone_RxByteCnt_reg[1]/NET0131 ,
		\wishbone_RxEnableWindow_reg/NET0131 ,
		_w26002_
	);
	LUT4 #(
		.INIT('h1115)
	) name15490 (
		\wishbone_RxDataLatched1_reg[16]/NET0131 ,
		_w25974_,
		_w26001_,
		_w26002_,
		_w26003_
	);
	LUT4 #(
		.INIT('h0400)
	) name15491 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_LastByteIn_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w26004_
	);
	LUT3 #(
		.INIT('he0)
	) name15492 (
		_w26001_,
		_w26002_,
		_w26004_,
		_w26005_
	);
	LUT2 #(
		.INIT('h1)
	) name15493 (
		_w26003_,
		_w26005_,
		_w26006_
	);
	LUT4 #(
		.INIT('h1115)
	) name15494 (
		\wishbone_RxDataLatched1_reg[17]/NET0131 ,
		_w25974_,
		_w26001_,
		_w26002_,
		_w26007_
	);
	LUT4 #(
		.INIT('h0400)
	) name15495 (
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_LastByteIn_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w26008_
	);
	LUT3 #(
		.INIT('he0)
	) name15496 (
		_w26001_,
		_w26002_,
		_w26008_,
		_w26009_
	);
	LUT2 #(
		.INIT('h1)
	) name15497 (
		_w26007_,
		_w26009_,
		_w26010_
	);
	LUT4 #(
		.INIT('h1115)
	) name15498 (
		\wishbone_RxDataLatched1_reg[18]/NET0131 ,
		_w25974_,
		_w26001_,
		_w26002_,
		_w26011_
	);
	LUT3 #(
		.INIT('ha8)
	) name15499 (
		_w25978_,
		_w26001_,
		_w26002_,
		_w26012_
	);
	LUT2 #(
		.INIT('h1)
	) name15500 (
		_w26011_,
		_w26012_,
		_w26013_
	);
	LUT4 #(
		.INIT('h1115)
	) name15501 (
		\wishbone_RxDataLatched1_reg[19]/NET0131 ,
		_w25974_,
		_w26001_,
		_w26002_,
		_w26014_
	);
	LUT3 #(
		.INIT('ha8)
	) name15502 (
		_w25982_,
		_w26001_,
		_w26002_,
		_w26015_
	);
	LUT2 #(
		.INIT('h1)
	) name15503 (
		_w26014_,
		_w26015_,
		_w26016_
	);
	LUT4 #(
		.INIT('h1115)
	) name15504 (
		\wishbone_RxDataLatched1_reg[20]/NET0131 ,
		_w25974_,
		_w26001_,
		_w26002_,
		_w26017_
	);
	LUT3 #(
		.INIT('ha8)
	) name15505 (
		_w25986_,
		_w26001_,
		_w26002_,
		_w26018_
	);
	LUT2 #(
		.INIT('h1)
	) name15506 (
		_w26017_,
		_w26018_,
		_w26019_
	);
	LUT4 #(
		.INIT('h1115)
	) name15507 (
		\wishbone_RxDataLatched1_reg[21]/NET0131 ,
		_w25974_,
		_w26001_,
		_w26002_,
		_w26020_
	);
	LUT3 #(
		.INIT('ha8)
	) name15508 (
		_w25990_,
		_w26001_,
		_w26002_,
		_w26021_
	);
	LUT2 #(
		.INIT('h1)
	) name15509 (
		_w26020_,
		_w26021_,
		_w26022_
	);
	LUT4 #(
		.INIT('h1115)
	) name15510 (
		\wishbone_RxDataLatched1_reg[22]/NET0131 ,
		_w25974_,
		_w26001_,
		_w26002_,
		_w26023_
	);
	LUT3 #(
		.INIT('ha8)
	) name15511 (
		_w25994_,
		_w26001_,
		_w26002_,
		_w26024_
	);
	LUT2 #(
		.INIT('h1)
	) name15512 (
		_w26023_,
		_w26024_,
		_w26025_
	);
	LUT4 #(
		.INIT('h1115)
	) name15513 (
		\wishbone_RxDataLatched1_reg[23]/NET0131 ,
		_w25974_,
		_w26001_,
		_w26002_,
		_w26026_
	);
	LUT3 #(
		.INIT('ha8)
	) name15514 (
		_w25998_,
		_w26001_,
		_w26002_,
		_w26027_
	);
	LUT2 #(
		.INIT('h1)
	) name15515 (
		_w26026_,
		_w26027_,
		_w26028_
	);
	LUT4 #(
		.INIT('h0100)
	) name15516 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		\wishbone_RxByteCnt_reg[1]/NET0131 ,
		\wishbone_RxEnableWindow_reg/NET0131 ,
		_w26029_
	);
	LUT3 #(
		.INIT('h02)
	) name15517 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w26030_
	);
	LUT4 #(
		.INIT('h1115)
	) name15518 (
		\wishbone_RxDataLatched1_reg[24]/NET0131 ,
		_w25974_,
		_w26029_,
		_w26030_,
		_w26031_
	);
	LUT3 #(
		.INIT('ha8)
	) name15519 (
		_w26004_,
		_w26029_,
		_w26030_,
		_w26032_
	);
	LUT2 #(
		.INIT('h1)
	) name15520 (
		_w26031_,
		_w26032_,
		_w26033_
	);
	LUT4 #(
		.INIT('h1115)
	) name15521 (
		\wishbone_RxDataLatched1_reg[25]/NET0131 ,
		_w25974_,
		_w26029_,
		_w26030_,
		_w26034_
	);
	LUT3 #(
		.INIT('ha8)
	) name15522 (
		_w26008_,
		_w26029_,
		_w26030_,
		_w26035_
	);
	LUT2 #(
		.INIT('h1)
	) name15523 (
		_w26034_,
		_w26035_,
		_w26036_
	);
	LUT4 #(
		.INIT('h1115)
	) name15524 (
		\wishbone_RxDataLatched1_reg[26]/NET0131 ,
		_w25974_,
		_w26029_,
		_w26030_,
		_w26037_
	);
	LUT3 #(
		.INIT('ha8)
	) name15525 (
		_w25978_,
		_w26029_,
		_w26030_,
		_w26038_
	);
	LUT2 #(
		.INIT('h1)
	) name15526 (
		_w26037_,
		_w26038_,
		_w26039_
	);
	LUT4 #(
		.INIT('h1115)
	) name15527 (
		\wishbone_RxDataLatched1_reg[27]/NET0131 ,
		_w25974_,
		_w26029_,
		_w26030_,
		_w26040_
	);
	LUT3 #(
		.INIT('ha8)
	) name15528 (
		_w25982_,
		_w26029_,
		_w26030_,
		_w26041_
	);
	LUT2 #(
		.INIT('h1)
	) name15529 (
		_w26040_,
		_w26041_,
		_w26042_
	);
	LUT4 #(
		.INIT('h1115)
	) name15530 (
		\wishbone_RxDataLatched1_reg[28]/NET0131 ,
		_w25974_,
		_w26029_,
		_w26030_,
		_w26043_
	);
	LUT3 #(
		.INIT('ha8)
	) name15531 (
		_w25986_,
		_w26029_,
		_w26030_,
		_w26044_
	);
	LUT2 #(
		.INIT('h1)
	) name15532 (
		_w26043_,
		_w26044_,
		_w26045_
	);
	LUT4 #(
		.INIT('h1115)
	) name15533 (
		\wishbone_RxDataLatched1_reg[29]/NET0131 ,
		_w25974_,
		_w26029_,
		_w26030_,
		_w26046_
	);
	LUT3 #(
		.INIT('ha8)
	) name15534 (
		_w25990_,
		_w26029_,
		_w26030_,
		_w26047_
	);
	LUT2 #(
		.INIT('h1)
	) name15535 (
		_w26046_,
		_w26047_,
		_w26048_
	);
	LUT4 #(
		.INIT('h1115)
	) name15536 (
		\wishbone_RxDataLatched1_reg[30]/NET0131 ,
		_w25974_,
		_w26029_,
		_w26030_,
		_w26049_
	);
	LUT3 #(
		.INIT('ha8)
	) name15537 (
		_w25994_,
		_w26029_,
		_w26030_,
		_w26050_
	);
	LUT2 #(
		.INIT('h1)
	) name15538 (
		_w26049_,
		_w26050_,
		_w26051_
	);
	LUT4 #(
		.INIT('h1115)
	) name15539 (
		\wishbone_RxDataLatched1_reg[31]/NET0131 ,
		_w25974_,
		_w26029_,
		_w26030_,
		_w26052_
	);
	LUT3 #(
		.INIT('ha8)
	) name15540 (
		_w25998_,
		_w26029_,
		_w26030_,
		_w26053_
	);
	LUT2 #(
		.INIT('h1)
	) name15541 (
		_w26052_,
		_w26053_,
		_w26054_
	);
	LUT4 #(
		.INIT('h1115)
	) name15542 (
		\wishbone_RxDataLatched1_reg[8]/NET0131 ,
		_w25974_,
		_w25975_,
		_w25976_,
		_w26055_
	);
	LUT3 #(
		.INIT('he0)
	) name15543 (
		_w25975_,
		_w25976_,
		_w26004_,
		_w26056_
	);
	LUT2 #(
		.INIT('h1)
	) name15544 (
		_w26055_,
		_w26056_,
		_w26057_
	);
	LUT4 #(
		.INIT('h1115)
	) name15545 (
		\wishbone_RxDataLatched1_reg[9]/NET0131 ,
		_w25974_,
		_w25975_,
		_w25976_,
		_w26058_
	);
	LUT3 #(
		.INIT('he0)
	) name15546 (
		_w25975_,
		_w25976_,
		_w26008_,
		_w26059_
	);
	LUT2 #(
		.INIT('h1)
	) name15547 (
		_w26058_,
		_w26059_,
		_w26060_
	);
	LUT3 #(
		.INIT('h80)
	) name15548 (
		_w25809_,
		_w25864_,
		_w25870_,
		_w26061_
	);
	LUT3 #(
		.INIT('he2)
	) name15549 (
		\miim1_LatchByte0_d_reg/NET0131 ,
		_w25812_,
		_w26061_,
		_w26062_
	);
	LUT4 #(
		.INIT('haa2a)
	) name15550 (
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		_w11870_,
		_w11873_,
		_w11876_,
		_w26063_
	);
	LUT2 #(
		.INIT('h6)
	) name15551 (
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		_w26064_
	);
	LUT3 #(
		.INIT('h70)
	) name15552 (
		_w11868_,
		_w11875_,
		_w26064_,
		_w26065_
	);
	LUT3 #(
		.INIT('h80)
	) name15553 (
		_w11870_,
		_w11873_,
		_w26065_,
		_w26066_
	);
	LUT3 #(
		.INIT('hf8)
	) name15554 (
		_w24515_,
		_w26063_,
		_w26066_,
		_w26067_
	);
	LUT4 #(
		.INIT('haa2a)
	) name15555 (
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w11870_,
		_w11873_,
		_w11876_,
		_w26068_
	);
	LUT3 #(
		.INIT('h87)
	) name15556 (
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w26069_
	);
	LUT3 #(
		.INIT('h07)
	) name15557 (
		_w11868_,
		_w11875_,
		_w26069_,
		_w26070_
	);
	LUT3 #(
		.INIT('h80)
	) name15558 (
		_w11870_,
		_w11873_,
		_w26070_,
		_w26071_
	);
	LUT3 #(
		.INIT('hf8)
	) name15559 (
		_w24515_,
		_w26068_,
		_w26071_,
		_w26072_
	);
	LUT2 #(
		.INIT('h4)
	) name15560 (
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26073_
	);
	LUT2 #(
		.INIT('h2)
	) name15561 (
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26074_
	);
	LUT4 #(
		.INIT('h0008)
	) name15562 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_TxAbortPacket_reg/NET0131 ,
		\wishbone_TxRetryPacket_reg/NET0131 ,
		_w26075_
	);
	LUT4 #(
		.INIT('h7000)
	) name15563 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w26074_,
		_w26075_,
		_w26076_
	);
	LUT2 #(
		.INIT('h8)
	) name15564 (
		_w26073_,
		_w26076_,
		_w26077_
	);
	LUT2 #(
		.INIT('h4)
	) name15565 (
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26078_
	);
	LUT4 #(
		.INIT('h7000)
	) name15566 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w26075_,
		_w26078_,
		_w26079_
	);
	LUT2 #(
		.INIT('h8)
	) name15567 (
		_w26073_,
		_w26079_,
		_w26080_
	);
	LUT2 #(
		.INIT('h8)
	) name15568 (
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26081_
	);
	LUT2 #(
		.INIT('h8)
	) name15569 (
		_w26079_,
		_w26081_,
		_w26082_
	);
	LUT3 #(
		.INIT('h80)
	) name15570 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		_w26083_
	);
	LUT2 #(
		.INIT('h1)
	) name15571 (
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26084_
	);
	LUT4 #(
		.INIT('h7000)
	) name15572 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w26083_,
		_w26084_,
		_w26085_
	);
	LUT3 #(
		.INIT('h01)
	) name15573 (
		\wishbone_TxAbortPacket_reg/NET0131 ,
		\wishbone_TxRetryPacket_reg/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26086_
	);
	LUT2 #(
		.INIT('h8)
	) name15574 (
		_w26085_,
		_w26086_,
		_w26087_
	);
	LUT2 #(
		.INIT('h1)
	) name15575 (
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26088_
	);
	LUT2 #(
		.INIT('h8)
	) name15576 (
		_w26076_,
		_w26088_,
		_w26089_
	);
	LUT2 #(
		.INIT('h2)
	) name15577 (
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26090_
	);
	LUT2 #(
		.INIT('h8)
	) name15578 (
		_w26076_,
		_w26090_,
		_w26091_
	);
	LUT2 #(
		.INIT('h8)
	) name15579 (
		_w26079_,
		_w26088_,
		_w26092_
	);
	LUT2 #(
		.INIT('h8)
	) name15580 (
		_w26079_,
		_w26090_,
		_w26093_
	);
	LUT4 #(
		.INIT('h0008)
	) name15581 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26094_
	);
	LUT2 #(
		.INIT('h8)
	) name15582 (
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26095_
	);
	LUT4 #(
		.INIT('h1000)
	) name15583 (
		\wishbone_TxAbortPacket_reg/NET0131 ,
		\wishbone_TxRetryPacket_reg/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26096_
	);
	LUT4 #(
		.INIT('h7000)
	) name15584 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w26094_,
		_w26096_,
		_w26097_
	);
	LUT4 #(
		.INIT('h8000)
	) name15585 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		_w26098_
	);
	LUT4 #(
		.INIT('h0010)
	) name15586 (
		\wishbone_TxAbortPacket_reg/NET0131 ,
		\wishbone_TxRetryPacket_reg/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26099_
	);
	LUT4 #(
		.INIT('h7000)
	) name15587 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w26098_,
		_w26099_,
		_w26100_
	);
	LUT4 #(
		.INIT('h0001)
	) name15588 (
		\wishbone_TxAbortPacket_reg/NET0131 ,
		\wishbone_TxRetryPacket_reg/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26101_
	);
	LUT4 #(
		.INIT('h8000)
	) name15589 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26102_
	);
	LUT4 #(
		.INIT('h7000)
	) name15590 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w26101_,
		_w26102_,
		_w26103_
	);
	LUT3 #(
		.INIT('h64)
	) name15591 (
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		_w11902_,
		_w24515_,
		_w26104_
	);
	LUT3 #(
		.INIT('h80)
	) name15592 (
		\wishbone_tx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[1]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[2]/NET0131 ,
		_w26105_
	);
	LUT4 #(
		.INIT('ha2f7)
	) name15593 (
		_w25792_,
		_w25795_,
		_w25796_,
		_w26105_,
		_w26106_
	);
	LUT4 #(
		.INIT('h8884)
	) name15594 (
		\wishbone_tx_fifo_cnt_reg[3]/NET0131 ,
		_w25385_,
		_w25799_,
		_w26106_,
		_w26107_
	);
	LUT3 #(
		.INIT('h45)
	) name15595 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		_w25922_,
		_w25928_,
		_w26108_
	);
	LUT3 #(
		.INIT('h70)
	) name15596 (
		_w25924_,
		_w25927_,
		_w26108_,
		_w26109_
	);
	LUT2 #(
		.INIT('h4)
	) name15597 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		_w25933_,
		_w26110_
	);
	LUT3 #(
		.INIT('hb0)
	) name15598 (
		_w25922_,
		_w25928_,
		_w25933_,
		_w26111_
	);
	LUT4 #(
		.INIT('h080f)
	) name15599 (
		_w25924_,
		_w25927_,
		_w26110_,
		_w26111_,
		_w26112_
	);
	LUT2 #(
		.INIT('h1)
	) name15600 (
		_w26109_,
		_w26112_,
		_w26113_
	);
	LUT2 #(
		.INIT('h1)
	) name15601 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w26114_
	);
	LUT3 #(
		.INIT('h45)
	) name15602 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w25922_,
		_w25928_,
		_w26115_
	);
	LUT4 #(
		.INIT('h080f)
	) name15603 (
		_w25924_,
		_w25927_,
		_w26114_,
		_w26115_,
		_w26116_
	);
	LUT3 #(
		.INIT('h40)
	) name15604 (
		_w25931_,
		_w25933_,
		_w26116_,
		_w26117_
	);
	LUT4 #(
		.INIT('h8000)
	) name15605 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		_w26118_
	);
	LUT4 #(
		.INIT('hf800)
	) name15606 (
		_w25924_,
		_w25927_,
		_w25929_,
		_w26118_,
		_w26119_
	);
	LUT4 #(
		.INIT('h00c8)
	) name15607 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		_w25933_,
		_w25935_,
		_w26119_,
		_w26120_
	);
	LUT4 #(
		.INIT('h1000)
	) name15608 (
		\txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		_w26121_
	);
	LUT2 #(
		.INIT('h1)
	) name15609 (
		\txethmac1_PacketFinished_q_reg/NET0131 ,
		_w26121_,
		_w26122_
	);
	LUT2 #(
		.INIT('h4)
	) name15610 (
		_w10830_,
		_w26122_,
		_w26123_
	);
	LUT4 #(
		.INIT('hfe00)
	) name15611 (
		\txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		\txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		_w26124_
	);
	LUT3 #(
		.INIT('h07)
	) name15612 (
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w10801_,
		_w26124_,
		_w26125_
	);
	LUT2 #(
		.INIT('h8)
	) name15613 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		_w26126_
	);
	LUT4 #(
		.INIT('hf800)
	) name15614 (
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w10801_,
		_w26124_,
		_w26126_,
		_w26127_
	);
	LUT3 #(
		.INIT('hc6)
	) name15615 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		_w26125_,
		_w26128_
	);
	LUT2 #(
		.INIT('h8)
	) name15616 (
		_w26123_,
		_w26128_,
		_w26129_
	);
	LUT3 #(
		.INIT('h80)
	) name15617 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		_w26130_
	);
	LUT4 #(
		.INIT('hf800)
	) name15618 (
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w10801_,
		_w26124_,
		_w26130_,
		_w26131_
	);
	LUT4 #(
		.INIT('h1020)
	) name15619 (
		\txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		_w10830_,
		_w26122_,
		_w26131_,
		_w26132_
	);
	LUT4 #(
		.INIT('hfe7f)
	) name15620 (
		\wishbone_rx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[1]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[2]/NET0131 ,
		_w13809_,
		_w26133_
	);
	LUT4 #(
		.INIT('h2221)
	) name15621 (
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		_w24970_,
		_w25832_,
		_w26133_,
		_w26134_
	);
	LUT4 #(
		.INIT('h1000)
	) name15622 (
		\wb_adr_i[10]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		wb_we_i_pad,
		_w26135_
	);
	LUT4 #(
		.INIT('h4000)
	) name15623 (
		_w18750_,
		_w18753_,
		_w24750_,
		_w26135_,
		_w26136_
	);
	LUT3 #(
		.INIT('h08)
	) name15624 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_dat_i[1]_pad ,
		_w26137_
	);
	LUT2 #(
		.INIT('h2)
	) name15625 (
		\ethreg1_MIICOMMAND1_DataOut_reg[0]/NET0131 ,
		\miim1_RStatStart_reg/NET0131 ,
		_w26138_
	);
	LUT3 #(
		.INIT('h40)
	) name15626 (
		\miim1_RStatStart_reg/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		_w26139_
	);
	LUT4 #(
		.INIT('h7270)
	) name15627 (
		_w26136_,
		_w26137_,
		_w26138_,
		_w26139_,
		_w26140_
	);
	LUT3 #(
		.INIT('h08)
	) name15628 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_dat_i[2]_pad ,
		_w26141_
	);
	LUT2 #(
		.INIT('h2)
	) name15629 (
		\ethreg1_MIICOMMAND2_DataOut_reg[0]/NET0131 ,
		\miim1_WCtrlDataStart_reg/NET0131 ,
		_w26142_
	);
	LUT3 #(
		.INIT('h40)
	) name15630 (
		\miim1_WCtrlDataStart_reg/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		_w26143_
	);
	LUT4 #(
		.INIT('h7270)
	) name15631 (
		_w26136_,
		_w26141_,
		_w26142_,
		_w26143_,
		_w26144_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name15632 (
		_w25922_,
		_w25925_,
		_w25926_,
		_w25928_,
		_w26145_
	);
	LUT4 #(
		.INIT('h60a0)
	) name15633 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		_w25924_,
		_w25933_,
		_w26145_,
		_w26146_
	);
	LUT3 #(
		.INIT('h48)
	) name15634 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w25933_,
		_w26119_,
		_w26147_
	);
	LUT2 #(
		.INIT('h1)
	) name15635 (
		_w10745_,
		_w25955_,
		_w26148_
	);
	LUT3 #(
		.INIT('h08)
	) name15636 (
		_w10749_,
		_w10754_,
		_w25955_,
		_w26149_
	);
	LUT3 #(
		.INIT('h13)
	) name15637 (
		_w10744_,
		_w26148_,
		_w26149_,
		_w26150_
	);
	LUT2 #(
		.INIT('h1)
	) name15638 (
		\txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		_w26127_,
		_w26151_
	);
	LUT3 #(
		.INIT('h04)
	) name15639 (
		_w10830_,
		_w26122_,
		_w26131_,
		_w26152_
	);
	LUT2 #(
		.INIT('h4)
	) name15640 (
		_w26151_,
		_w26152_,
		_w26153_
	);
	LUT4 #(
		.INIT('h0002)
	) name15641 (
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_TxAbortPacket_NotCleared_reg/NET0131 ,
		\wishbone_TxRetryPacket_NotCleared_reg/NET0131 ,
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w26154_
	);
	LUT2 #(
		.INIT('h8)
	) name15642 (
		_w25801_,
		_w26154_,
		_w26155_
	);
	LUT3 #(
		.INIT('he0)
	) name15643 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		\wishbone_TxLength_reg[2]/NET0131 ,
		_w26156_
	);
	LUT2 #(
		.INIT('h1)
	) name15644 (
		\wishbone_TxLength_reg[3]/NET0131 ,
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w26157_
	);
	LUT3 #(
		.INIT('h20)
	) name15645 (
		_w26154_,
		_w26156_,
		_w26157_,
		_w26158_
	);
	LUT4 #(
		.INIT('h0002)
	) name15646 (
		\wishbone_BlockReadTxDataFromMemory_reg/NET0131 ,
		\wishbone_TxAbortPacket_reg/NET0131 ,
		\wishbone_TxDonePacket_reg/NET0131 ,
		\wishbone_TxRetryPacket_reg/NET0131 ,
		_w26159_
	);
	LUT2 #(
		.INIT('h4)
	) name15647 (
		_w25792_,
		_w26159_,
		_w26160_
	);
	LUT4 #(
		.INIT('hffec)
	) name15648 (
		_w24540_,
		_w26155_,
		_w26158_,
		_w26160_,
		_w26161_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name15649 (
		mdc_pad_o_pad,
		\miim1_InProgress_q1_reg/NET0131 ,
		_w24411_,
		_w24420_,
		_w26162_
	);
	LUT2 #(
		.INIT('he)
	) name15650 (
		_w25808_,
		_w26162_,
		_w26163_
	);
	LUT3 #(
		.INIT('h45)
	) name15651 (
		\rxethmac1_RxEndFrm_d_reg/NET0131 ,
		_w10575_,
		_w11386_,
		_w26164_
	);
	LUT3 #(
		.INIT('h15)
	) name15652 (
		\rxethmac1_RxEndFrm_d_reg/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w26165_
	);
	LUT3 #(
		.INIT('h13)
	) name15653 (
		_w10519_,
		_w26164_,
		_w26165_,
		_w26166_
	);
	LUT3 #(
		.INIT('h40)
	) name15654 (
		\wb_adr_i[10]_pad ,
		\wb_adr_i[2]_pad ,
		wb_we_i_pad,
		_w26167_
	);
	LUT4 #(
		.INIT('h4000)
	) name15655 (
		_w18750_,
		_w18753_,
		_w24750_,
		_w26167_,
		_w26168_
	);
	LUT4 #(
		.INIT('h0100)
	) name15656 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		\wb_dat_i[2]_pad ,
		_w26169_
	);
	LUT4 #(
		.INIT('hceee)
	) name15657 (
		\ethreg1_irq_rxb_reg/NET0131 ,
		\wishbone_RxB_IRQ_reg/NET0131 ,
		_w26168_,
		_w26169_,
		_w26170_
	);
	LUT4 #(
		.INIT('h0100)
	) name15658 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		\wb_dat_i[6]_pad ,
		_w26171_
	);
	LUT4 #(
		.INIT('haeee)
	) name15659 (
		\ethreg1_SetRxCIrq_reg/NET0131 ,
		\ethreg1_irq_rxc_reg/NET0131 ,
		_w26168_,
		_w26171_,
		_w26172_
	);
	LUT4 #(
		.INIT('h0100)
	) name15660 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		\wb_dat_i[3]_pad ,
		_w26173_
	);
	LUT4 #(
		.INIT('hceee)
	) name15661 (
		\ethreg1_irq_rxe_reg/NET0131 ,
		\wishbone_RxE_IRQ_reg/NET0131 ,
		_w26168_,
		_w26173_,
		_w26174_
	);
	LUT4 #(
		.INIT('h0100)
	) name15662 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		\wb_dat_i[0]_pad ,
		_w26175_
	);
	LUT4 #(
		.INIT('hceee)
	) name15663 (
		\ethreg1_irq_txb_reg/NET0131 ,
		\wishbone_TxB_IRQ_reg/NET0131 ,
		_w26168_,
		_w26175_,
		_w26176_
	);
	LUT4 #(
		.INIT('h0100)
	) name15664 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		\wb_dat_i[5]_pad ,
		_w26177_
	);
	LUT4 #(
		.INIT('haeee)
	) name15665 (
		\ethreg1_SetTxCIrq_reg/NET0131 ,
		\ethreg1_irq_txc_reg/NET0131 ,
		_w26168_,
		_w26177_,
		_w26178_
	);
	LUT4 #(
		.INIT('h0100)
	) name15666 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		\wb_dat_i[1]_pad ,
		_w26179_
	);
	LUT4 #(
		.INIT('hceee)
	) name15667 (
		\ethreg1_irq_txe_reg/NET0131 ,
		\wishbone_TxE_IRQ_reg/NET0131 ,
		_w26168_,
		_w26179_,
		_w26180_
	);
	LUT4 #(
		.INIT('h002a)
	) name15668 (
		\txethmac1_ColWindow_reg/NET0131 ,
		_w10785_,
		_w10786_,
		_w10825_,
		_w26181_
	);
	LUT4 #(
		.INIT('he0a0)
	) name15669 (
		\txethmac1_TxRetry_reg/NET0131 ,
		_w10830_,
		_w11075_,
		_w26181_,
		_w26182_
	);
	LUT3 #(
		.INIT('h08)
	) name15670 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w26183_
	);
	LUT2 #(
		.INIT('h2)
	) name15671 (
		\wishbone_Busy_IRQ_rck_reg/NET0131 ,
		\wishbone_Busy_IRQ_syncb2_reg/P0001 ,
		_w26184_
	);
	LUT2 #(
		.INIT('he)
	) name15672 (
		_w26183_,
		_w26184_,
		_w26185_
	);
	LUT4 #(
		.INIT('h8000)
	) name15673 (
		\wishbone_RxBDAddress_reg[1]/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w26186_
	);
	LUT3 #(
		.INIT('h13)
	) name15674 (
		\wishbone_RxBDAddress_reg[2]/NET0131 ,
		\wishbone_RxBDAddress_reg[3]/NET0131 ,
		_w26186_,
		_w26187_
	);
	LUT4 #(
		.INIT('h0111)
	) name15675 (
		_w25875_,
		_w25876_,
		_w25879_,
		_w25880_,
		_w26188_
	);
	LUT3 #(
		.INIT('ha8)
	) name15676 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[2]/NET0131 ,
		_w25875_,
		_w25876_,
		_w26189_
	);
	LUT3 #(
		.INIT('hf4)
	) name15677 (
		_w26187_,
		_w26188_,
		_w26189_,
		_w26190_
	);
	LUT4 #(
		.INIT('h3aca)
	) name15678 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[4]/NET0131 ,
		\wishbone_RxBDAddress_reg[5]/NET0131 ,
		_w25877_,
		_w25883_,
		_w26191_
	);
	LUT3 #(
		.INIT('ha8)
	) name15679 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[5]/NET0131 ,
		_w25875_,
		_w25876_,
		_w26192_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name15680 (
		\wishbone_RxBDAddress_reg[6]/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w26193_
	);
	LUT4 #(
		.INIT('h00ea)
	) name15681 (
		\wishbone_RxStatus_reg[13]/NET0131 ,
		_w25880_,
		_w25969_,
		_w26193_,
		_w26194_
	);
	LUT4 #(
		.INIT('h5555)
	) name15682 (
		\wishbone_RxBDAddress_reg[6]/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w26195_
	);
	LUT4 #(
		.INIT('h7f00)
	) name15683 (
		\wishbone_RxBDAddress_reg[5]/NET0131 ,
		_w25880_,
		_w25882_,
		_w26195_,
		_w26196_
	);
	LUT4 #(
		.INIT('hcccd)
	) name15684 (
		_w25875_,
		_w26192_,
		_w26194_,
		_w26196_,
		_w26197_
	);
	LUT3 #(
		.INIT('h63)
	) name15685 (
		\miim1_clkgen_Counter_reg[4]/NET0131 ,
		\miim1_clkgen_Counter_reg[5]/NET0131 ,
		_w24411_,
		_w26198_
	);
	LUT4 #(
		.INIT('h0aaa)
	) name15686 (
		\ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131 ,
		_w24413_,
		_w24416_,
		_w26199_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name15687 (
		_w24421_,
		_w25908_,
		_w26198_,
		_w26199_,
		_w26200_
	);
	LUT4 #(
		.INIT('h0080)
	) name15688 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26201_
	);
	LUT3 #(
		.INIT('h70)
	) name15689 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w26201_,
		_w26202_
	);
	LUT4 #(
		.INIT('h8880)
	) name15690 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_TxAbortPacket_reg/NET0131 ,
		\wishbone_TxRetryPacket_reg/NET0131 ,
		_w26203_
	);
	LUT2 #(
		.INIT('h2)
	) name15691 (
		_w26073_,
		_w26203_,
		_w26204_
	);
	LUT4 #(
		.INIT('haccc)
	) name15692 (
		\m_wb_dat_i[14]_pad ,
		\wishbone_tx_fifo_fifo_reg[10][14]/P0001 ,
		_w26202_,
		_w26204_,
		_w26205_
	);
	LUT4 #(
		.INIT('haccc)
	) name15693 (
		\m_wb_dat_i[18]_pad ,
		\wishbone_tx_fifo_fifo_reg[10][18]/P0001 ,
		_w26202_,
		_w26204_,
		_w26206_
	);
	LUT4 #(
		.INIT('haccc)
	) name15694 (
		\m_wb_dat_i[27]_pad ,
		\wishbone_tx_fifo_fifo_reg[10][27]/P0001 ,
		_w26202_,
		_w26204_,
		_w26207_
	);
	LUT4 #(
		.INIT('haccc)
	) name15695 (
		\m_wb_dat_i[29]_pad ,
		\wishbone_tx_fifo_fifo_reg[10][29]/P0001 ,
		_w26202_,
		_w26204_,
		_w26208_
	);
	LUT4 #(
		.INIT('haccc)
	) name15696 (
		\m_wb_dat_i[3]_pad ,
		\wishbone_tx_fifo_fifo_reg[10][3]/P0001 ,
		_w26202_,
		_w26204_,
		_w26209_
	);
	LUT4 #(
		.INIT('h0800)
	) name15697 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26210_
	);
	LUT3 #(
		.INIT('h70)
	) name15698 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w26210_,
		_w26211_
	);
	LUT4 #(
		.INIT('haccc)
	) name15699 (
		\m_wb_dat_i[12]_pad ,
		\wishbone_tx_fifo_fifo_reg[12][12]/P0001 ,
		_w26204_,
		_w26211_,
		_w26212_
	);
	LUT4 #(
		.INIT('haccc)
	) name15700 (
		\m_wb_dat_i[14]_pad ,
		\wishbone_tx_fifo_fifo_reg[12][14]/P0001 ,
		_w26204_,
		_w26211_,
		_w26213_
	);
	LUT4 #(
		.INIT('haccc)
	) name15701 (
		\m_wb_dat_i[18]_pad ,
		\wishbone_tx_fifo_fifo_reg[12][18]/P0001 ,
		_w26204_,
		_w26211_,
		_w26214_
	);
	LUT4 #(
		.INIT('haccc)
	) name15702 (
		\m_wb_dat_i[22]_pad ,
		\wishbone_tx_fifo_fifo_reg[12][22]/P0001 ,
		_w26204_,
		_w26211_,
		_w26215_
	);
	LUT4 #(
		.INIT('haccc)
	) name15703 (
		\m_wb_dat_i[25]_pad ,
		\wishbone_tx_fifo_fifo_reg[12][25]/P0001 ,
		_w26204_,
		_w26211_,
		_w26216_
	);
	LUT4 #(
		.INIT('haccc)
	) name15704 (
		\m_wb_dat_i[27]_pad ,
		\wishbone_tx_fifo_fifo_reg[12][27]/P0001 ,
		_w26204_,
		_w26211_,
		_w26217_
	);
	LUT4 #(
		.INIT('haccc)
	) name15705 (
		\m_wb_dat_i[28]_pad ,
		\wishbone_tx_fifo_fifo_reg[12][28]/P0001 ,
		_w26204_,
		_w26211_,
		_w26218_
	);
	LUT4 #(
		.INIT('haccc)
	) name15706 (
		\m_wb_dat_i[30]_pad ,
		\wishbone_tx_fifo_fifo_reg[12][30]/P0001 ,
		_w26204_,
		_w26211_,
		_w26219_
	);
	LUT4 #(
		.INIT('haccc)
	) name15707 (
		\m_wb_dat_i[3]_pad ,
		\wishbone_tx_fifo_fifo_reg[12][3]/P0001 ,
		_w26204_,
		_w26211_,
		_w26220_
	);
	LUT4 #(
		.INIT('haccc)
	) name15708 (
		\m_wb_dat_i[6]_pad ,
		\wishbone_tx_fifo_fifo_reg[12][6]/P0001 ,
		_w26204_,
		_w26211_,
		_w26221_
	);
	LUT2 #(
		.INIT('h2)
	) name15709 (
		_w26090_,
		_w26203_,
		_w26222_
	);
	LUT4 #(
		.INIT('haccc)
	) name15710 (
		\m_wb_dat_i[10]_pad ,
		\wishbone_tx_fifo_fifo_reg[3][10]/P0001 ,
		_w26202_,
		_w26222_,
		_w26223_
	);
	LUT4 #(
		.INIT('haccc)
	) name15711 (
		\m_wb_dat_i[11]_pad ,
		\wishbone_tx_fifo_fifo_reg[3][11]/P0001 ,
		_w26202_,
		_w26222_,
		_w26224_
	);
	LUT4 #(
		.INIT('haccc)
	) name15712 (
		\m_wb_dat_i[13]_pad ,
		\wishbone_tx_fifo_fifo_reg[3][13]/P0001 ,
		_w26202_,
		_w26222_,
		_w26225_
	);
	LUT4 #(
		.INIT('haccc)
	) name15713 (
		\m_wb_dat_i[18]_pad ,
		\wishbone_tx_fifo_fifo_reg[3][18]/P0001 ,
		_w26202_,
		_w26222_,
		_w26226_
	);
	LUT4 #(
		.INIT('haccc)
	) name15714 (
		\m_wb_dat_i[19]_pad ,
		\wishbone_tx_fifo_fifo_reg[3][19]/P0001 ,
		_w26202_,
		_w26222_,
		_w26227_
	);
	LUT4 #(
		.INIT('haccc)
	) name15715 (
		\m_wb_dat_i[25]_pad ,
		\wishbone_tx_fifo_fifo_reg[3][25]/P0001 ,
		_w26202_,
		_w26222_,
		_w26228_
	);
	LUT4 #(
		.INIT('haccc)
	) name15716 (
		\m_wb_dat_i[29]_pad ,
		\wishbone_tx_fifo_fifo_reg[3][29]/P0001 ,
		_w26202_,
		_w26222_,
		_w26229_
	);
	LUT4 #(
		.INIT('haccc)
	) name15717 (
		\m_wb_dat_i[31]_pad ,
		\wishbone_tx_fifo_fifo_reg[3][31]/P0001 ,
		_w26202_,
		_w26222_,
		_w26230_
	);
	LUT4 #(
		.INIT('haccc)
	) name15718 (
		\m_wb_dat_i[4]_pad ,
		\wishbone_tx_fifo_fifo_reg[3][4]/P0001 ,
		_w26202_,
		_w26222_,
		_w26231_
	);
	LUT4 #(
		.INIT('haccc)
	) name15719 (
		\m_wb_dat_i[5]_pad ,
		\wishbone_tx_fifo_fifo_reg[3][5]/P0001 ,
		_w26202_,
		_w26222_,
		_w26232_
	);
	LUT4 #(
		.INIT('haccc)
	) name15720 (
		\m_wb_dat_i[8]_pad ,
		\wishbone_tx_fifo_fifo_reg[3][8]/P0001 ,
		_w26202_,
		_w26222_,
		_w26233_
	);
	LUT4 #(
		.INIT('haccc)
	) name15721 (
		\m_wb_dat_i[11]_pad ,
		\wishbone_tx_fifo_fifo_reg[5][11]/P0001 ,
		_w26211_,
		_w26222_,
		_w26234_
	);
	LUT4 #(
		.INIT('haccc)
	) name15722 (
		\m_wb_dat_i[18]_pad ,
		\wishbone_tx_fifo_fifo_reg[5][18]/P0001 ,
		_w26211_,
		_w26222_,
		_w26235_
	);
	LUT4 #(
		.INIT('haccc)
	) name15723 (
		\m_wb_dat_i[19]_pad ,
		\wishbone_tx_fifo_fifo_reg[5][19]/P0001 ,
		_w26211_,
		_w26222_,
		_w26236_
	);
	LUT4 #(
		.INIT('haccc)
	) name15724 (
		\m_wb_dat_i[1]_pad ,
		\wishbone_tx_fifo_fifo_reg[5][1]/P0001 ,
		_w26211_,
		_w26222_,
		_w26237_
	);
	LUT4 #(
		.INIT('haccc)
	) name15725 (
		\m_wb_dat_i[23]_pad ,
		\wishbone_tx_fifo_fifo_reg[5][23]/P0001 ,
		_w26211_,
		_w26222_,
		_w26238_
	);
	LUT4 #(
		.INIT('haccc)
	) name15726 (
		\m_wb_dat_i[24]_pad ,
		\wishbone_tx_fifo_fifo_reg[5][24]/P0001 ,
		_w26211_,
		_w26222_,
		_w26239_
	);
	LUT4 #(
		.INIT('haccc)
	) name15727 (
		\m_wb_dat_i[25]_pad ,
		\wishbone_tx_fifo_fifo_reg[5][25]/P0001 ,
		_w26211_,
		_w26222_,
		_w26240_
	);
	LUT4 #(
		.INIT('haccc)
	) name15728 (
		\m_wb_dat_i[26]_pad ,
		\wishbone_tx_fifo_fifo_reg[5][26]/P0001 ,
		_w26211_,
		_w26222_,
		_w26241_
	);
	LUT4 #(
		.INIT('haccc)
	) name15729 (
		\m_wb_dat_i[28]_pad ,
		\wishbone_tx_fifo_fifo_reg[5][28]/P0001 ,
		_w26211_,
		_w26222_,
		_w26242_
	);
	LUT4 #(
		.INIT('haccc)
	) name15730 (
		\m_wb_dat_i[3]_pad ,
		\wishbone_tx_fifo_fifo_reg[5][3]/P0001 ,
		_w26211_,
		_w26222_,
		_w26243_
	);
	LUT4 #(
		.INIT('haccc)
	) name15731 (
		\m_wb_dat_i[8]_pad ,
		\wishbone_tx_fifo_fifo_reg[5][8]/P0001 ,
		_w26211_,
		_w26222_,
		_w26244_
	);
	LUT3 #(
		.INIT('h70)
	) name15732 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w26094_,
		_w26245_
	);
	LUT2 #(
		.INIT('h2)
	) name15733 (
		_w26095_,
		_w26203_,
		_w26246_
	);
	LUT4 #(
		.INIT('haccc)
	) name15734 (
		\m_wb_dat_i[11]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][11]/P0001 ,
		_w26245_,
		_w26246_,
		_w26247_
	);
	LUT4 #(
		.INIT('haccc)
	) name15735 (
		\m_wb_dat_i[12]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][12]/P0001 ,
		_w26245_,
		_w26246_,
		_w26248_
	);
	LUT4 #(
		.INIT('haccc)
	) name15736 (
		\m_wb_dat_i[14]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][14]/P0001 ,
		_w26245_,
		_w26246_,
		_w26249_
	);
	LUT4 #(
		.INIT('haccc)
	) name15737 (
		\m_wb_dat_i[16]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][16]/P0001 ,
		_w26245_,
		_w26246_,
		_w26250_
	);
	LUT4 #(
		.INIT('haccc)
	) name15738 (
		\m_wb_dat_i[18]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][18]/P0001 ,
		_w26245_,
		_w26246_,
		_w26251_
	);
	LUT4 #(
		.INIT('haccc)
	) name15739 (
		\m_wb_dat_i[1]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][1]/P0001 ,
		_w26245_,
		_w26246_,
		_w26252_
	);
	LUT4 #(
		.INIT('haccc)
	) name15740 (
		\m_wb_dat_i[20]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][20]/P0001 ,
		_w26245_,
		_w26246_,
		_w26253_
	);
	LUT4 #(
		.INIT('haccc)
	) name15741 (
		\m_wb_dat_i[25]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][25]/P0001 ,
		_w26245_,
		_w26246_,
		_w26254_
	);
	LUT4 #(
		.INIT('haccc)
	) name15742 (
		\m_wb_dat_i[27]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][27]/P0001 ,
		_w26245_,
		_w26246_,
		_w26255_
	);
	LUT4 #(
		.INIT('haccc)
	) name15743 (
		\m_wb_dat_i[28]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][28]/P0001 ,
		_w26245_,
		_w26246_,
		_w26256_
	);
	LUT4 #(
		.INIT('haccc)
	) name15744 (
		\m_wb_dat_i[30]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][30]/P0001 ,
		_w26245_,
		_w26246_,
		_w26257_
	);
	LUT4 #(
		.INIT('haccc)
	) name15745 (
		\m_wb_dat_i[3]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][3]/P0001 ,
		_w26245_,
		_w26246_,
		_w26258_
	);
	LUT4 #(
		.INIT('haccc)
	) name15746 (
		\m_wb_dat_i[4]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][4]/P0001 ,
		_w26245_,
		_w26246_,
		_w26259_
	);
	LUT4 #(
		.INIT('haccc)
	) name15747 (
		\m_wb_dat_i[5]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][5]/P0001 ,
		_w26245_,
		_w26246_,
		_w26260_
	);
	LUT4 #(
		.INIT('haccc)
	) name15748 (
		\m_wb_dat_i[6]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][6]/P0001 ,
		_w26245_,
		_w26246_,
		_w26261_
	);
	LUT4 #(
		.INIT('haccc)
	) name15749 (
		\m_wb_dat_i[7]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][7]/P0001 ,
		_w26245_,
		_w26246_,
		_w26262_
	);
	LUT4 #(
		.INIT('haccc)
	) name15750 (
		\m_wb_dat_i[8]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][8]/P0001 ,
		_w26245_,
		_w26246_,
		_w26263_
	);
	LUT2 #(
		.INIT('h2)
	) name15751 (
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26203_,
		_w26264_
	);
	LUT4 #(
		.INIT('haccc)
	) name15752 (
		\m_wb_dat_i[12]_pad ,
		\wishbone_tx_fifo_fifo_reg[9][12]/P0001 ,
		_w26085_,
		_w26264_,
		_w26265_
	);
	LUT4 #(
		.INIT('haccc)
	) name15753 (
		\m_wb_dat_i[13]_pad ,
		\wishbone_tx_fifo_fifo_reg[9][13]/P0001 ,
		_w26085_,
		_w26264_,
		_w26266_
	);
	LUT4 #(
		.INIT('haccc)
	) name15754 (
		\m_wb_dat_i[14]_pad ,
		\wishbone_tx_fifo_fifo_reg[9][14]/P0001 ,
		_w26085_,
		_w26264_,
		_w26267_
	);
	LUT4 #(
		.INIT('haccc)
	) name15755 (
		\m_wb_dat_i[20]_pad ,
		\wishbone_tx_fifo_fifo_reg[9][20]/P0001 ,
		_w26085_,
		_w26264_,
		_w26268_
	);
	LUT4 #(
		.INIT('haccc)
	) name15756 (
		\m_wb_dat_i[25]_pad ,
		\wishbone_tx_fifo_fifo_reg[9][25]/P0001 ,
		_w26085_,
		_w26264_,
		_w26269_
	);
	LUT4 #(
		.INIT('haccc)
	) name15757 (
		\m_wb_dat_i[26]_pad ,
		\wishbone_tx_fifo_fifo_reg[9][26]/P0001 ,
		_w26085_,
		_w26264_,
		_w26270_
	);
	LUT4 #(
		.INIT('haccc)
	) name15758 (
		\m_wb_dat_i[30]_pad ,
		\wishbone_tx_fifo_fifo_reg[9][30]/P0001 ,
		_w26085_,
		_w26264_,
		_w26271_
	);
	LUT4 #(
		.INIT('haccc)
	) name15759 (
		\m_wb_dat_i[5]_pad ,
		\wishbone_tx_fifo_fifo_reg[9][5]/P0001 ,
		_w26085_,
		_w26264_,
		_w26272_
	);
	LUT4 #(
		.INIT('haccc)
	) name15760 (
		\m_wb_dat_i[8]_pad ,
		\wishbone_tx_fifo_fifo_reg[9][8]/P0001 ,
		_w26085_,
		_w26264_,
		_w26273_
	);
	LUT4 #(
		.INIT('haccc)
	) name15761 (
		\m_wb_dat_i[23]_pad ,
		\wishbone_tx_fifo_fifo_reg[6][23]/P0001 ,
		_w26245_,
		_w26246_,
		_w26274_
	);
	LUT4 #(
		.INIT('h0008)
	) name15762 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26275_
	);
	LUT4 #(
		.INIT('h7000)
	) name15763 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w26088_,
		_w26275_,
		_w26276_
	);
	LUT2 #(
		.INIT('he)
	) name15764 (
		_w26203_,
		_w26276_,
		_w26277_
	);
	LUT2 #(
		.INIT('h8)
	) name15765 (
		_w26076_,
		_w26081_,
		_w26278_
	);
	LUT4 #(
		.INIT('h0800)
	) name15766 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26279_
	);
	LUT4 #(
		.INIT('h7000)
	) name15767 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w26096_,
		_w26279_,
		_w26280_
	);
	LUT4 #(
		.INIT('h7000)
	) name15768 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w26096_,
		_w26102_,
		_w26281_
	);
	LUT4 #(
		.INIT('h7000)
	) name15769 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w26101_,
		_w26279_,
		_w26282_
	);
	LUT2 #(
		.INIT('h2)
	) name15770 (
		\wishbone_Busy_IRQ_sync2_reg/P0001 ,
		\wishbone_Busy_IRQ_sync3_reg/P0001 ,
		_w26283_
	);
	LUT4 #(
		.INIT('h0100)
	) name15771 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		\wb_dat_i[4]_pad ,
		_w26284_
	);
	LUT4 #(
		.INIT('hf2fa)
	) name15772 (
		\ethreg1_irq_busy_reg/NET0131 ,
		_w26168_,
		_w26283_,
		_w26284_,
		_w26285_
	);
	LUT2 #(
		.INIT('h4)
	) name15773 (
		\miim1_LatchByte_reg[0]/NET0131 ,
		\miim1_LatchByte_reg[1]/NET0131 ,
		_w26286_
	);
	LUT4 #(
		.INIT('h5700)
	) name15774 (
		_w24568_,
		_w24572_,
		_w24573_,
		_w26286_,
		_w26287_
	);
	LUT4 #(
		.INIT('h0200)
	) name15775 (
		_w24561_,
		_w24567_,
		_w24571_,
		_w26287_,
		_w26288_
	);
	LUT3 #(
		.INIT('hb0)
	) name15776 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[0]/NET0131 ,
		_w26289_
	);
	LUT2 #(
		.INIT('h9)
	) name15777 (
		_w25832_,
		_w26289_,
		_w26290_
	);
	LUT4 #(
		.INIT('h72d8)
	) name15778 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		\wishbone_LatchedRxLength_reg[13]/NET0131 ,
		_w11147_,
		_w26291_
	);
	LUT2 #(
		.INIT('h6)
	) name15779 (
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		_w11140_,
		_w26292_
	);
	LUT2 #(
		.INIT('h1)
	) name15780 (
		_w11138_,
		_w11162_,
		_w26293_
	);
	LUT2 #(
		.INIT('hd)
	) name15781 (
		_w10582_,
		_w11398_,
		_w26294_
	);
	LUT4 #(
		.INIT('h7f0f)
	) name15782 (
		_w10554_,
		_w10573_,
		_w10582_,
		_w11113_,
		_w26295_
	);
	LUT4 #(
		.INIT('h7000)
	) name15783 (
		_w10554_,
		_w10573_,
		_w10577_,
		_w10946_,
		_w26296_
	);
	LUT2 #(
		.INIT('hd)
	) name15784 (
		_w10582_,
		_w26296_,
		_w26297_
	);
	LUT4 #(
		.INIT('h0013)
	) name15785 (
		_w11866_,
		_w25828_,
		_w25830_,
		_w25834_,
		_w26298_
	);
	LUT4 #(
		.INIT('h0033)
	) name15786 (
		\wishbone_rx_fifo_cnt_reg[2]/NET0131 ,
		_w11865_,
		_w25829_,
		_w25831_,
		_w26299_
	);
	LUT4 #(
		.INIT('h2221)
	) name15787 (
		\wishbone_rx_fifo_cnt_reg[2]/NET0131 ,
		_w24970_,
		_w26298_,
		_w26299_,
		_w26300_
	);
	LUT3 #(
		.INIT('h0e)
	) name15788 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\wishbone_LatchedRxStartFrm_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		_w26301_
	);
	LUT4 #(
		.INIT('h8000)
	) name15789 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		_w26302_
	);
	LUT2 #(
		.INIT('h8)
	) name15790 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w26303_
	);
	LUT4 #(
		.INIT('h0200)
	) name15791 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131 ,
		_w26304_
	);
	LUT4 #(
		.INIT('h0006)
	) name15792 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131 ,
		_w26302_,
		_w26303_,
		_w26304_,
		_w26305_
	);
	LUT2 #(
		.INIT('h6)
	) name15793 (
		\wishbone_rx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[1]/NET0131 ,
		_w26306_
	);
	LUT4 #(
		.INIT('h00ec)
	) name15794 (
		_w11866_,
		_w25828_,
		_w25830_,
		_w26306_,
		_w26307_
	);
	LUT4 #(
		.INIT('h7000)
	) name15795 (
		_w11866_,
		_w25829_,
		_w25831_,
		_w26306_,
		_w26308_
	);
	LUT4 #(
		.INIT('h0007)
	) name15796 (
		\wishbone_rx_fifo_cnt_reg[1]/NET0131 ,
		_w25832_,
		_w26307_,
		_w26308_,
		_w26309_
	);
	LUT2 #(
		.INIT('h1)
	) name15797 (
		_w24970_,
		_w26309_,
		_w26310_
	);
	LUT2 #(
		.INIT('h8)
	) name15798 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_SlotTimer_reg[2]/NET0131 ,
		_w26311_
	);
	LUT3 #(
		.INIT('h15)
	) name15799 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[3]/NET0131 ,
		_w11279_,
		_w26311_,
		_w26312_
	);
	LUT3 #(
		.INIT('h15)
	) name15800 (
		wb_rst_i_pad,
		_w11279_,
		_w11280_,
		_w26313_
	);
	LUT2 #(
		.INIT('h4)
	) name15801 (
		_w26312_,
		_w26313_,
		_w26314_
	);
	LUT3 #(
		.INIT('h8a)
	) name15802 (
		\wishbone_StartOccured_reg/NET0131 ,
		\wishbone_TxDone_wb_q_reg/NET0131 ,
		\wishbone_TxDone_wb_reg/NET0131 ,
		_w26315_
	);
	LUT3 #(
		.INIT('hea)
	) name15803 (
		\wishbone_TxStartFrm_wb_reg/NET0131 ,
		_w25940_,
		_w26315_,
		_w26316_
	);
	LUT4 #(
		.INIT('h0001)
	) name15804 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[5]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[6]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131 ,
		_w26317_
	);
	LUT4 #(
		.INIT('h0001)
	) name15805 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[3]/NET0131 ,
		_w26318_
	);
	LUT2 #(
		.INIT('h2)
	) name15806 (
		\ethreg1_MODER_0_DataOut_reg[1]/NET0131 ,
		\wishbone_r_TxEn_q_reg/NET0131 ,
		_w26319_
	);
	LUT3 #(
		.INIT('h70)
	) name15807 (
		_w26317_,
		_w26318_,
		_w26319_,
		_w26320_
	);
	LUT4 #(
		.INIT('he000)
	) name15808 (
		\wishbone_TxAbortPacket_NotCleared_reg/NET0131 ,
		\wishbone_TxDonePacket_NotCleared_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w26321_
	);
	LUT2 #(
		.INIT('h4)
	) name15809 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		_w26321_,
		_w26322_
	);
	LUT3 #(
		.INIT('h8c)
	) name15810 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		\wishbone_TxBDAddress_reg[4]/NET0131 ,
		_w26321_,
		_w26323_
	);
	LUT2 #(
		.INIT('h1)
	) name15811 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		\wishbone_TxStatus_reg[13]/NET0131 ,
		_w26324_
	);
	LUT2 #(
		.INIT('h8)
	) name15812 (
		_w26321_,
		_w26324_,
		_w26325_
	);
	LUT4 #(
		.INIT('h8000)
	) name15813 (
		\wishbone_TxBDAddress_reg[1]/NET0131 ,
		\wishbone_TxBDAddress_reg[2]/NET0131 ,
		\wishbone_TxBDAddress_reg[3]/NET0131 ,
		\wishbone_TxBDAddress_reg[4]/NET0131 ,
		_w26326_
	);
	LUT4 #(
		.INIT('h7f80)
	) name15814 (
		\wishbone_TxBDAddress_reg[1]/NET0131 ,
		\wishbone_TxBDAddress_reg[2]/NET0131 ,
		\wishbone_TxBDAddress_reg[3]/NET0131 ,
		\wishbone_TxBDAddress_reg[4]/NET0131 ,
		_w26327_
	);
	LUT4 #(
		.INIT('h5444)
	) name15815 (
		_w26320_,
		_w26323_,
		_w26325_,
		_w26327_,
		_w26328_
	);
	LUT2 #(
		.INIT('h8)
	) name15816 (
		\wishbone_TxBDAddress_reg[5]/NET0131 ,
		\wishbone_TxBDAddress_reg[6]/NET0131 ,
		_w26329_
	);
	LUT4 #(
		.INIT('h0888)
	) name15817 (
		_w26321_,
		_w26324_,
		_w26326_,
		_w26329_,
		_w26330_
	);
	LUT4 #(
		.INIT('h2202)
	) name15818 (
		\wishbone_TxBDAddress_reg[6]/NET0131 ,
		_w26320_,
		_w26322_,
		_w26330_,
		_w26331_
	);
	LUT2 #(
		.INIT('h8)
	) name15819 (
		\wishbone_TxBDAddress_reg[5]/NET0131 ,
		_w26326_,
		_w26332_
	);
	LUT3 #(
		.INIT('h40)
	) name15820 (
		_w26320_,
		_w26330_,
		_w26332_,
		_w26333_
	);
	LUT2 #(
		.INIT('he)
	) name15821 (
		_w26331_,
		_w26333_,
		_w26334_
	);
	LUT4 #(
		.INIT('h2202)
	) name15822 (
		\wishbone_TxBDAddress_reg[7]/NET0131 ,
		_w26320_,
		_w26322_,
		_w26330_,
		_w26335_
	);
	LUT3 #(
		.INIT('h08)
	) name15823 (
		\wishbone_TxBDAddress_reg[5]/NET0131 ,
		\wishbone_TxBDAddress_reg[6]/NET0131 ,
		\wishbone_TxBDAddress_reg[7]/NET0131 ,
		_w26336_
	);
	LUT4 #(
		.INIT('h8000)
	) name15824 (
		_w26321_,
		_w26324_,
		_w26326_,
		_w26336_,
		_w26337_
	);
	LUT2 #(
		.INIT('h4)
	) name15825 (
		_w26320_,
		_w26337_,
		_w26338_
	);
	LUT2 #(
		.INIT('he)
	) name15826 (
		_w26335_,
		_w26338_,
		_w26339_
	);
	LUT3 #(
		.INIT('hb0)
	) name15827 (
		\wishbone_TxDone_wb_q_reg/NET0131 ,
		\wishbone_TxDone_wb_reg/NET0131 ,
		\wishbone_TxEndFrm_wb_reg/NET0131 ,
		_w26340_
	);
	LUT2 #(
		.INIT('h8)
	) name15828 (
		_w25940_,
		_w26340_,
		_w26341_
	);
	LUT3 #(
		.INIT('h80)
	) name15829 (
		_w12314_,
		_w12316_,
		_w14520_,
		_w26342_
	);
	LUT3 #(
		.INIT('h02)
	) name15830 (
		\wishbone_tx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[1]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[2]/NET0131 ,
		_w26343_
	);
	LUT4 #(
		.INIT('h0004)
	) name15831 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w26344_
	);
	LUT2 #(
		.INIT('h8)
	) name15832 (
		_w26343_,
		_w26344_,
		_w26345_
	);
	LUT4 #(
		.INIT('heccc)
	) name15833 (
		_w12312_,
		_w26341_,
		_w26342_,
		_w26345_,
		_w26346_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name15834 (
		mdc_pad_o_pad,
		\miim1_outctrl_Mdo_2d_reg/NET0131 ,
		_w24411_,
		_w24420_,
		_w26347_
	);
	LUT3 #(
		.INIT('h0e)
	) name15835 (
		\miim1_BitCounter_reg[4]/NET0131 ,
		\miim1_BitCounter_reg[6]/NET0131 ,
		\miim1_WriteOp_reg/NET0131 ,
		_w26348_
	);
	LUT4 #(
		.INIT('h0080)
	) name15836 (
		\miim1_BitCounter_reg[1]/NET0131 ,
		\miim1_BitCounter_reg[2]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		\miim1_WriteOp_reg/NET0131 ,
		_w26349_
	);
	LUT3 #(
		.INIT('he0)
	) name15837 (
		\miim1_BitCounter_reg[5]/NET0131 ,
		\miim1_BitCounter_reg[6]/NET0131 ,
		\miim1_InProgress_reg/NET0131 ,
		_w26350_
	);
	LUT3 #(
		.INIT('h10)
	) name15838 (
		_w26348_,
		_w26349_,
		_w26350_,
		_w26351_
	);
	LUT3 #(
		.INIT('h02)
	) name15839 (
		mdc_pad_o_pad,
		\miim1_BitCounter_reg[5]/NET0131 ,
		\miim1_BitCounter_reg[6]/NET0131 ,
		_w26352_
	);
	LUT3 #(
		.INIT('h80)
	) name15840 (
		_w24411_,
		_w24420_,
		_w26352_,
		_w26353_
	);
	LUT4 #(
		.INIT('hcdcc)
	) name15841 (
		_w24567_,
		_w26347_,
		_w26351_,
		_w26353_,
		_w26354_
	);
	LUT4 #(
		.INIT('h0200)
	) name15842 (
		\ethreg1_TXCTRL_0_DataOut_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26355_
	);
	LUT4 #(
		.INIT('hffd3)
	) name15843 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26356_
	);
	LUT3 #(
		.INIT('h8a)
	) name15844 (
		_w25925_,
		_w26355_,
		_w26356_,
		_w26357_
	);
	LUT2 #(
		.INIT('h1)
	) name15845 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		_w26358_
	);
	LUT3 #(
		.INIT('h10)
	) name15846 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w26359_
	);
	LUT4 #(
		.INIT('h0008)
	) name15847 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26360_
	);
	LUT3 #(
		.INIT('h04)
	) name15848 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26361_
	);
	LUT4 #(
		.INIT('h0200)
	) name15849 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w26362_
	);
	LUT4 #(
		.INIT('h0777)
	) name15850 (
		_w26359_,
		_w26360_,
		_w26361_,
		_w26362_,
		_w26363_
	);
	LUT2 #(
		.INIT('h4)
	) name15851 (
		_w26357_,
		_w26363_,
		_w26364_
	);
	LUT3 #(
		.INIT('h01)
	) name15852 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w26365_
	);
	LUT3 #(
		.INIT('h01)
	) name15853 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26366_
	);
	LUT4 #(
		.INIT('h0200)
	) name15854 (
		\ethreg1_TXCTRL_1_DataOut_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26367_
	);
	LUT4 #(
		.INIT('h0020)
	) name15855 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26368_
	);
	LUT4 #(
		.INIT('h000b)
	) name15856 (
		_w25922_,
		_w26366_,
		_w26367_,
		_w26368_,
		_w26369_
	);
	LUT3 #(
		.INIT('h40)
	) name15857 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w26370_
	);
	LUT4 #(
		.INIT('h0008)
	) name15858 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26371_
	);
	LUT4 #(
		.INIT('h00e0)
	) name15859 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26372_
	);
	LUT3 #(
		.INIT('ha8)
	) name15860 (
		_w26370_,
		_w26371_,
		_w26372_,
		_w26373_
	);
	LUT3 #(
		.INIT('h0d)
	) name15861 (
		_w26365_,
		_w26369_,
		_w26373_,
		_w26374_
	);
	LUT2 #(
		.INIT('h7)
	) name15862 (
		_w26364_,
		_w26374_,
		_w26375_
	);
	LUT2 #(
		.INIT('h8)
	) name15863 (
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w26376_
	);
	LUT3 #(
		.INIT('h2a)
	) name15864 (
		\txethmac1_random1_RandomLatched_reg[9]/NET0131 ,
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w26377_
	);
	LUT2 #(
		.INIT('h1)
	) name15865 (
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		_w26378_
	);
	LUT4 #(
		.INIT('h8000)
	) name15866 (
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		\txethmac1_random1_x_reg[9]/NET0131 ,
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w26379_
	);
	LUT3 #(
		.INIT('hba)
	) name15867 (
		_w26377_,
		_w26378_,
		_w26379_,
		_w26380_
	);
	LUT4 #(
		.INIT('h0100)
	) name15868 (
		\wishbone_RxEn_needed_reg/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26381_
	);
	LUT4 #(
		.INIT('hfef3)
	) name15869 (
		\wishbone_RxEn_needed_reg/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26382_
	);
	LUT2 #(
		.INIT('h2)
	) name15870 (
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26382_,
		_w26383_
	);
	LUT3 #(
		.INIT('h0d)
	) name15871 (
		\wishbone_RxEn_needed_reg/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26384_
	);
	LUT4 #(
		.INIT('h00f2)
	) name15872 (
		\wishbone_RxEn_needed_reg/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		_w26385_
	);
	LUT3 #(
		.INIT('h07)
	) name15873 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26386_
	);
	LUT2 #(
		.INIT('h4)
	) name15874 (
		_w26385_,
		_w26386_,
		_w26387_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name15875 (
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26382_,
		_w26385_,
		_w26386_,
		_w26388_
	);
	LUT4 #(
		.INIT('h0200)
	) name15876 (
		\wishbone_RxEn_needed_reg/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26389_
	);
	LUT2 #(
		.INIT('h2)
	) name15877 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		_w26389_,
		_w26390_
	);
	LUT4 #(
		.INIT('h002a)
	) name15878 (
		\wb_adr_i[2]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26391_
	);
	LUT2 #(
		.INIT('h4)
	) name15879 (
		_w26385_,
		_w26391_,
		_w26392_
	);
	LUT2 #(
		.INIT('h8)
	) name15880 (
		\wishbone_TxEn_needed_reg/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w26393_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15881 (
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w26382_,
		_w26389_,
		_w26393_,
		_w26394_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15882 (
		_w26388_,
		_w26390_,
		_w26392_,
		_w26394_,
		_w26395_
	);
	LUT2 #(
		.INIT('h2)
	) name15883 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		_w26389_,
		_w26396_
	);
	LUT4 #(
		.INIT('h002a)
	) name15884 (
		\wb_adr_i[3]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26397_
	);
	LUT2 #(
		.INIT('h4)
	) name15885 (
		_w26385_,
		_w26397_,
		_w26398_
	);
	LUT2 #(
		.INIT('h8)
	) name15886 (
		\wishbone_TxBDAddress_reg[1]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26399_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15887 (
		\wishbone_RxBDAddress_reg[1]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26399_,
		_w26400_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15888 (
		_w26388_,
		_w26396_,
		_w26398_,
		_w26400_,
		_w26401_
	);
	LUT2 #(
		.INIT('h2)
	) name15889 (
		\wishbone_ram_addr_reg[2]/NET0131 ,
		_w26389_,
		_w26402_
	);
	LUT4 #(
		.INIT('h002a)
	) name15890 (
		\wb_adr_i[4]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26403_
	);
	LUT2 #(
		.INIT('h4)
	) name15891 (
		_w26385_,
		_w26403_,
		_w26404_
	);
	LUT2 #(
		.INIT('h8)
	) name15892 (
		\wishbone_TxBDAddress_reg[2]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26405_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15893 (
		\wishbone_RxBDAddress_reg[2]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26405_,
		_w26406_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15894 (
		_w26388_,
		_w26402_,
		_w26404_,
		_w26406_,
		_w26407_
	);
	LUT2 #(
		.INIT('h2)
	) name15895 (
		\wishbone_ram_addr_reg[3]/NET0131 ,
		_w26389_,
		_w26408_
	);
	LUT4 #(
		.INIT('h002a)
	) name15896 (
		\wb_adr_i[5]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26409_
	);
	LUT2 #(
		.INIT('h4)
	) name15897 (
		_w26385_,
		_w26409_,
		_w26410_
	);
	LUT2 #(
		.INIT('h8)
	) name15898 (
		\wishbone_TxBDAddress_reg[3]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26411_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15899 (
		\wishbone_RxBDAddress_reg[3]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26411_,
		_w26412_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15900 (
		_w26388_,
		_w26408_,
		_w26410_,
		_w26412_,
		_w26413_
	);
	LUT2 #(
		.INIT('h2)
	) name15901 (
		\wishbone_ram_addr_reg[4]/NET0131 ,
		_w26389_,
		_w26414_
	);
	LUT4 #(
		.INIT('h002a)
	) name15902 (
		\wb_adr_i[6]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26415_
	);
	LUT2 #(
		.INIT('h4)
	) name15903 (
		_w26385_,
		_w26415_,
		_w26416_
	);
	LUT2 #(
		.INIT('h8)
	) name15904 (
		\wishbone_TxBDAddress_reg[4]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26417_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15905 (
		\wishbone_RxBDAddress_reg[4]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26417_,
		_w26418_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15906 (
		_w26388_,
		_w26414_,
		_w26416_,
		_w26418_,
		_w26419_
	);
	LUT2 #(
		.INIT('h2)
	) name15907 (
		\wishbone_ram_addr_reg[5]/NET0131 ,
		_w26389_,
		_w26420_
	);
	LUT4 #(
		.INIT('h002a)
	) name15908 (
		\wb_adr_i[7]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26421_
	);
	LUT2 #(
		.INIT('h4)
	) name15909 (
		_w26385_,
		_w26421_,
		_w26422_
	);
	LUT2 #(
		.INIT('h8)
	) name15910 (
		\wishbone_TxBDAddress_reg[5]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26423_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15911 (
		\wishbone_RxBDAddress_reg[5]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26423_,
		_w26424_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15912 (
		_w26388_,
		_w26420_,
		_w26422_,
		_w26424_,
		_w26425_
	);
	LUT2 #(
		.INIT('h2)
	) name15913 (
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w26389_,
		_w26426_
	);
	LUT4 #(
		.INIT('h002a)
	) name15914 (
		\wb_adr_i[8]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26427_
	);
	LUT2 #(
		.INIT('h4)
	) name15915 (
		_w26385_,
		_w26427_,
		_w26428_
	);
	LUT2 #(
		.INIT('h8)
	) name15916 (
		\wishbone_TxBDAddress_reg[6]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26429_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15917 (
		\wishbone_RxBDAddress_reg[6]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26429_,
		_w26430_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15918 (
		_w26388_,
		_w26426_,
		_w26428_,
		_w26430_,
		_w26431_
	);
	LUT2 #(
		.INIT('h2)
	) name15919 (
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w26389_,
		_w26432_
	);
	LUT4 #(
		.INIT('h002a)
	) name15920 (
		\wb_adr_i[9]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26433_
	);
	LUT2 #(
		.INIT('h4)
	) name15921 (
		_w26385_,
		_w26433_,
		_w26434_
	);
	LUT2 #(
		.INIT('h8)
	) name15922 (
		\wishbone_TxBDAddress_reg[7]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26435_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15923 (
		\wishbone_RxBDAddress_reg[7]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26435_,
		_w26436_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15924 (
		_w26388_,
		_w26432_,
		_w26434_,
		_w26436_,
		_w26437_
	);
	LUT2 #(
		.INIT('h2)
	) name15925 (
		\wishbone_ram_di_reg[0]/NET0131 ,
		_w26389_,
		_w26438_
	);
	LUT4 #(
		.INIT('h002a)
	) name15926 (
		\wb_dat_i[0]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26439_
	);
	LUT2 #(
		.INIT('h4)
	) name15927 (
		_w26385_,
		_w26439_,
		_w26440_
	);
	LUT2 #(
		.INIT('h8)
	) name15928 (
		\macstatus1_CarrierSenseLost_reg/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26441_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15929 (
		\wishbone_RxStatusInLatched_reg[0]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26441_,
		_w26442_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15930 (
		_w26388_,
		_w26438_,
		_w26440_,
		_w26442_,
		_w26443_
	);
	LUT2 #(
		.INIT('h2)
	) name15931 (
		\wishbone_ram_di_reg[13]/NET0131 ,
		_w26389_,
		_w26444_
	);
	LUT4 #(
		.INIT('h002a)
	) name15932 (
		\wb_dat_i[13]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26445_
	);
	LUT2 #(
		.INIT('h4)
	) name15933 (
		_w26385_,
		_w26445_,
		_w26446_
	);
	LUT2 #(
		.INIT('h8)
	) name15934 (
		\wishbone_TxEn_needed_reg/NET0131 ,
		\wishbone_TxStatus_reg[13]/NET0131 ,
		_w26447_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15935 (
		\wishbone_RxStatus_reg[13]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26447_,
		_w26448_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15936 (
		_w26388_,
		_w26444_,
		_w26446_,
		_w26448_,
		_w26449_
	);
	LUT2 #(
		.INIT('h2)
	) name15937 (
		\wishbone_ram_di_reg[14]/NET0131 ,
		_w26389_,
		_w26450_
	);
	LUT4 #(
		.INIT('h002a)
	) name15938 (
		\wb_dat_i[14]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26451_
	);
	LUT2 #(
		.INIT('h4)
	) name15939 (
		_w26385_,
		_w26451_,
		_w26452_
	);
	LUT2 #(
		.INIT('h8)
	) name15940 (
		\wishbone_TxEn_needed_reg/NET0131 ,
		\wishbone_TxStatus_reg[14]/NET0131 ,
		_w26453_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15941 (
		\wishbone_RxStatus_reg[14]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26453_,
		_w26454_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15942 (
		_w26388_,
		_w26450_,
		_w26452_,
		_w26454_,
		_w26455_
	);
	LUT2 #(
		.INIT('h2)
	) name15943 (
		\wishbone_ram_di_reg[16]/NET0131 ,
		_w26389_,
		_w26456_
	);
	LUT2 #(
		.INIT('h8)
	) name15944 (
		\wishbone_LatchedTxLength_reg[0]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26457_
	);
	LUT2 #(
		.INIT('h4)
	) name15945 (
		_w26382_,
		_w26457_,
		_w26458_
	);
	LUT4 #(
		.INIT('h002a)
	) name15946 (
		\wb_dat_i[16]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26459_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15947 (
		\wishbone_LatchedRxLength_reg[0]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26459_,
		_w26460_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15948 (
		_w26388_,
		_w26456_,
		_w26458_,
		_w26460_,
		_w26461_
	);
	LUT2 #(
		.INIT('h2)
	) name15949 (
		\wishbone_ram_di_reg[17]/NET0131 ,
		_w26389_,
		_w26462_
	);
	LUT2 #(
		.INIT('h8)
	) name15950 (
		\wishbone_LatchedTxLength_reg[1]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26463_
	);
	LUT2 #(
		.INIT('h4)
	) name15951 (
		_w26382_,
		_w26463_,
		_w26464_
	);
	LUT4 #(
		.INIT('h002a)
	) name15952 (
		\wb_dat_i[17]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26465_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15953 (
		\wishbone_LatchedRxLength_reg[1]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26465_,
		_w26466_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15954 (
		_w26388_,
		_w26462_,
		_w26464_,
		_w26466_,
		_w26467_
	);
	LUT2 #(
		.INIT('h2)
	) name15955 (
		\wishbone_ram_di_reg[18]/NET0131 ,
		_w26389_,
		_w26468_
	);
	LUT2 #(
		.INIT('h8)
	) name15956 (
		\wishbone_LatchedTxLength_reg[2]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26469_
	);
	LUT2 #(
		.INIT('h4)
	) name15957 (
		_w26382_,
		_w26469_,
		_w26470_
	);
	LUT4 #(
		.INIT('h002a)
	) name15958 (
		\wb_dat_i[18]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26471_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15959 (
		\wishbone_LatchedRxLength_reg[2]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26471_,
		_w26472_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15960 (
		_w26388_,
		_w26468_,
		_w26470_,
		_w26472_,
		_w26473_
	);
	LUT2 #(
		.INIT('h2)
	) name15961 (
		\wishbone_ram_di_reg[19]/NET0131 ,
		_w26389_,
		_w26474_
	);
	LUT2 #(
		.INIT('h8)
	) name15962 (
		\wishbone_LatchedTxLength_reg[3]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26475_
	);
	LUT2 #(
		.INIT('h4)
	) name15963 (
		_w26382_,
		_w26475_,
		_w26476_
	);
	LUT4 #(
		.INIT('h002a)
	) name15964 (
		\wb_dat_i[19]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26477_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15965 (
		\wishbone_LatchedRxLength_reg[3]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26477_,
		_w26478_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15966 (
		_w26388_,
		_w26474_,
		_w26476_,
		_w26478_,
		_w26479_
	);
	LUT2 #(
		.INIT('h2)
	) name15967 (
		\wishbone_ram_di_reg[1]/NET0131 ,
		_w26389_,
		_w26480_
	);
	LUT4 #(
		.INIT('h002a)
	) name15968 (
		\wb_dat_i[1]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26481_
	);
	LUT2 #(
		.INIT('h4)
	) name15969 (
		_w26385_,
		_w26481_,
		_w26482_
	);
	LUT2 #(
		.INIT('h8)
	) name15970 (
		\macstatus1_DeferLatched_reg/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26483_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15971 (
		\wishbone_RxStatusInLatched_reg[1]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26483_,
		_w26484_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15972 (
		_w26388_,
		_w26480_,
		_w26482_,
		_w26484_,
		_w26485_
	);
	LUT2 #(
		.INIT('h2)
	) name15973 (
		\wishbone_ram_di_reg[20]/NET0131 ,
		_w26389_,
		_w26486_
	);
	LUT2 #(
		.INIT('h8)
	) name15974 (
		\wishbone_LatchedTxLength_reg[4]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26487_
	);
	LUT2 #(
		.INIT('h4)
	) name15975 (
		_w26382_,
		_w26487_,
		_w26488_
	);
	LUT4 #(
		.INIT('h002a)
	) name15976 (
		\wb_dat_i[20]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26489_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15977 (
		\wishbone_LatchedRxLength_reg[4]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26489_,
		_w26490_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15978 (
		_w26388_,
		_w26486_,
		_w26488_,
		_w26490_,
		_w26491_
	);
	LUT2 #(
		.INIT('h2)
	) name15979 (
		\wishbone_ram_di_reg[21]/NET0131 ,
		_w26389_,
		_w26492_
	);
	LUT2 #(
		.INIT('h8)
	) name15980 (
		\wishbone_LatchedTxLength_reg[5]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26493_
	);
	LUT2 #(
		.INIT('h4)
	) name15981 (
		_w26382_,
		_w26493_,
		_w26494_
	);
	LUT4 #(
		.INIT('h002a)
	) name15982 (
		\wb_dat_i[21]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26495_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15983 (
		\wishbone_LatchedRxLength_reg[5]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26495_,
		_w26496_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15984 (
		_w26388_,
		_w26492_,
		_w26494_,
		_w26496_,
		_w26497_
	);
	LUT2 #(
		.INIT('h2)
	) name15985 (
		\wishbone_ram_di_reg[22]/NET0131 ,
		_w26389_,
		_w26498_
	);
	LUT2 #(
		.INIT('h8)
	) name15986 (
		\wishbone_LatchedTxLength_reg[6]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26499_
	);
	LUT2 #(
		.INIT('h4)
	) name15987 (
		_w26382_,
		_w26499_,
		_w26500_
	);
	LUT4 #(
		.INIT('h002a)
	) name15988 (
		\wb_dat_i[22]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26501_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15989 (
		\wishbone_LatchedRxLength_reg[6]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26501_,
		_w26502_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15990 (
		_w26388_,
		_w26498_,
		_w26500_,
		_w26502_,
		_w26503_
	);
	LUT2 #(
		.INIT('h2)
	) name15991 (
		\wishbone_ram_di_reg[23]/NET0131 ,
		_w26389_,
		_w26504_
	);
	LUT4 #(
		.INIT('h002a)
	) name15992 (
		\wb_dat_i[23]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26505_
	);
	LUT2 #(
		.INIT('h4)
	) name15993 (
		_w26385_,
		_w26505_,
		_w26506_
	);
	LUT2 #(
		.INIT('h8)
	) name15994 (
		\wishbone_LatchedTxLength_reg[7]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26507_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15995 (
		\wishbone_LatchedRxLength_reg[7]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26507_,
		_w26508_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name15996 (
		_w26388_,
		_w26504_,
		_w26506_,
		_w26508_,
		_w26509_
	);
	LUT2 #(
		.INIT('h2)
	) name15997 (
		\wishbone_ram_di_reg[24]/NET0131 ,
		_w26389_,
		_w26510_
	);
	LUT4 #(
		.INIT('h002a)
	) name15998 (
		\wb_dat_i[24]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26511_
	);
	LUT2 #(
		.INIT('h4)
	) name15999 (
		_w26385_,
		_w26511_,
		_w26512_
	);
	LUT2 #(
		.INIT('h8)
	) name16000 (
		\wishbone_LatchedTxLength_reg[8]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26513_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16001 (
		\wishbone_LatchedRxLength_reg[8]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26513_,
		_w26514_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name16002 (
		_w26388_,
		_w26510_,
		_w26512_,
		_w26514_,
		_w26515_
	);
	LUT2 #(
		.INIT('h2)
	) name16003 (
		\wishbone_ram_di_reg[25]/NET0131 ,
		_w26389_,
		_w26516_
	);
	LUT2 #(
		.INIT('h8)
	) name16004 (
		\wishbone_LatchedTxLength_reg[9]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26517_
	);
	LUT2 #(
		.INIT('h4)
	) name16005 (
		_w26382_,
		_w26517_,
		_w26518_
	);
	LUT4 #(
		.INIT('h002a)
	) name16006 (
		\wb_dat_i[25]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26519_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16007 (
		\wishbone_LatchedRxLength_reg[9]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26519_,
		_w26520_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name16008 (
		_w26388_,
		_w26516_,
		_w26518_,
		_w26520_,
		_w26521_
	);
	LUT2 #(
		.INIT('h2)
	) name16009 (
		\wishbone_ram_di_reg[26]/NET0131 ,
		_w26389_,
		_w26522_
	);
	LUT2 #(
		.INIT('h8)
	) name16010 (
		\wishbone_LatchedTxLength_reg[10]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26523_
	);
	LUT2 #(
		.INIT('h4)
	) name16011 (
		_w26382_,
		_w26523_,
		_w26524_
	);
	LUT4 #(
		.INIT('h002a)
	) name16012 (
		\wb_dat_i[26]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26525_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16013 (
		\wishbone_LatchedRxLength_reg[10]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26525_,
		_w26526_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name16014 (
		_w26388_,
		_w26522_,
		_w26524_,
		_w26526_,
		_w26527_
	);
	LUT2 #(
		.INIT('h2)
	) name16015 (
		\wishbone_ram_di_reg[27]/NET0131 ,
		_w26389_,
		_w26528_
	);
	LUT4 #(
		.INIT('h002a)
	) name16016 (
		\wb_dat_i[27]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26529_
	);
	LUT2 #(
		.INIT('h4)
	) name16017 (
		_w26385_,
		_w26529_,
		_w26530_
	);
	LUT2 #(
		.INIT('h8)
	) name16018 (
		\wishbone_LatchedTxLength_reg[11]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26531_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16019 (
		\wishbone_LatchedRxLength_reg[11]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26531_,
		_w26532_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name16020 (
		_w26388_,
		_w26528_,
		_w26530_,
		_w26532_,
		_w26533_
	);
	LUT2 #(
		.INIT('h2)
	) name16021 (
		\wishbone_ram_di_reg[28]/NET0131 ,
		_w26389_,
		_w26534_
	);
	LUT2 #(
		.INIT('h8)
	) name16022 (
		\wishbone_LatchedTxLength_reg[12]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26535_
	);
	LUT2 #(
		.INIT('h4)
	) name16023 (
		_w26382_,
		_w26535_,
		_w26536_
	);
	LUT4 #(
		.INIT('h002a)
	) name16024 (
		\wb_dat_i[28]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26537_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16025 (
		\wishbone_LatchedRxLength_reg[12]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26537_,
		_w26538_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name16026 (
		_w26388_,
		_w26534_,
		_w26536_,
		_w26538_,
		_w26539_
	);
	LUT2 #(
		.INIT('h2)
	) name16027 (
		\wishbone_ram_di_reg[29]/NET0131 ,
		_w26389_,
		_w26540_
	);
	LUT4 #(
		.INIT('h002a)
	) name16028 (
		\wb_dat_i[29]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26541_
	);
	LUT2 #(
		.INIT('h4)
	) name16029 (
		_w26385_,
		_w26541_,
		_w26542_
	);
	LUT2 #(
		.INIT('h8)
	) name16030 (
		\wishbone_LatchedTxLength_reg[13]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26543_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16031 (
		\wishbone_LatchedRxLength_reg[13]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26543_,
		_w26544_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name16032 (
		_w26388_,
		_w26540_,
		_w26542_,
		_w26544_,
		_w26545_
	);
	LUT2 #(
		.INIT('h2)
	) name16033 (
		\wishbone_ram_di_reg[2]/NET0131 ,
		_w26389_,
		_w26546_
	);
	LUT2 #(
		.INIT('h8)
	) name16034 (
		\macstatus1_LateCollLatched_reg/P0002 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26547_
	);
	LUT2 #(
		.INIT('h4)
	) name16035 (
		_w26382_,
		_w26547_,
		_w26548_
	);
	LUT4 #(
		.INIT('h002a)
	) name16036 (
		\wb_dat_i[2]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26549_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16037 (
		\wishbone_RxStatusInLatched_reg[2]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26549_,
		_w26550_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name16038 (
		_w26388_,
		_w26546_,
		_w26548_,
		_w26550_,
		_w26551_
	);
	LUT2 #(
		.INIT('h2)
	) name16039 (
		\wishbone_ram_di_reg[30]/NET0131 ,
		_w26389_,
		_w26552_
	);
	LUT2 #(
		.INIT('h8)
	) name16040 (
		\wishbone_LatchedTxLength_reg[14]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26553_
	);
	LUT2 #(
		.INIT('h4)
	) name16041 (
		_w26382_,
		_w26553_,
		_w26554_
	);
	LUT4 #(
		.INIT('h002a)
	) name16042 (
		\wb_dat_i[30]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26555_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16043 (
		\wishbone_LatchedRxLength_reg[14]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26555_,
		_w26556_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name16044 (
		_w26388_,
		_w26552_,
		_w26554_,
		_w26556_,
		_w26557_
	);
	LUT2 #(
		.INIT('h2)
	) name16045 (
		\wishbone_ram_di_reg[31]/NET0131 ,
		_w26389_,
		_w26558_
	);
	LUT2 #(
		.INIT('h8)
	) name16046 (
		\wishbone_LatchedTxLength_reg[15]/NET0131 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26559_
	);
	LUT2 #(
		.INIT('h4)
	) name16047 (
		_w26382_,
		_w26559_,
		_w26560_
	);
	LUT4 #(
		.INIT('h002a)
	) name16048 (
		\wb_dat_i[31]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26561_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16049 (
		\wishbone_LatchedRxLength_reg[15]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26561_,
		_w26562_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name16050 (
		_w26388_,
		_w26558_,
		_w26560_,
		_w26562_,
		_w26563_
	);
	LUT2 #(
		.INIT('h2)
	) name16051 (
		\wishbone_ram_di_reg[3]/NET0131 ,
		_w26389_,
		_w26564_
	);
	LUT4 #(
		.INIT('h002a)
	) name16052 (
		\wb_dat_i[3]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26565_
	);
	LUT2 #(
		.INIT('h4)
	) name16053 (
		_w26385_,
		_w26565_,
		_w26566_
	);
	LUT2 #(
		.INIT('h8)
	) name16054 (
		\macstatus1_RetryLimit_reg/P0002 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26567_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16055 (
		\wishbone_RxStatusInLatched_reg[3]/NET0131 ,
		_w26382_,
		_w26389_,
		_w26567_,
		_w26568_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name16056 (
		_w26388_,
		_w26564_,
		_w26566_,
		_w26568_,
		_w26569_
	);
	LUT2 #(
		.INIT('h2)
	) name16057 (
		\wishbone_ram_di_reg[4]/NET0131 ,
		_w26389_,
		_w26570_
	);
	LUT2 #(
		.INIT('h8)
	) name16058 (
		\macstatus1_RetryCntLatched_reg[0]/P0002 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26571_
	);
	LUT2 #(
		.INIT('h4)
	) name16059 (
		_w26382_,
		_w26571_,
		_w26572_
	);
	LUT4 #(
		.INIT('h002a)
	) name16060 (
		\wb_dat_i[4]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26573_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16061 (
		\wishbone_RxStatusInLatched_reg[4]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26573_,
		_w26574_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name16062 (
		_w26388_,
		_w26570_,
		_w26572_,
		_w26574_,
		_w26575_
	);
	LUT2 #(
		.INIT('h2)
	) name16063 (
		\wishbone_ram_di_reg[5]/NET0131 ,
		_w26389_,
		_w26576_
	);
	LUT2 #(
		.INIT('h8)
	) name16064 (
		\macstatus1_RetryCntLatched_reg[1]/P0002 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26577_
	);
	LUT2 #(
		.INIT('h4)
	) name16065 (
		_w26382_,
		_w26577_,
		_w26578_
	);
	LUT4 #(
		.INIT('h002a)
	) name16066 (
		\wb_dat_i[5]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26579_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16067 (
		\wishbone_RxStatusInLatched_reg[5]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26579_,
		_w26580_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name16068 (
		_w26388_,
		_w26576_,
		_w26578_,
		_w26580_,
		_w26581_
	);
	LUT2 #(
		.INIT('h2)
	) name16069 (
		\wishbone_ram_di_reg[6]/NET0131 ,
		_w26389_,
		_w26582_
	);
	LUT2 #(
		.INIT('h8)
	) name16070 (
		\macstatus1_RetryCntLatched_reg[2]/P0002 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26583_
	);
	LUT2 #(
		.INIT('h4)
	) name16071 (
		_w26382_,
		_w26583_,
		_w26584_
	);
	LUT4 #(
		.INIT('h002a)
	) name16072 (
		\wb_dat_i[6]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26585_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16073 (
		\wishbone_RxStatusInLatched_reg[6]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26585_,
		_w26586_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name16074 (
		_w26388_,
		_w26582_,
		_w26584_,
		_w26586_,
		_w26587_
	);
	LUT2 #(
		.INIT('h2)
	) name16075 (
		\wishbone_ram_di_reg[7]/NET0131 ,
		_w26389_,
		_w26588_
	);
	LUT2 #(
		.INIT('h8)
	) name16076 (
		\macstatus1_RetryCntLatched_reg[3]/P0002 ,
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w26589_
	);
	LUT2 #(
		.INIT('h4)
	) name16077 (
		_w26382_,
		_w26589_,
		_w26590_
	);
	LUT4 #(
		.INIT('h002a)
	) name16078 (
		\wb_dat_i[7]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26591_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16079 (
		\wishbone_RxStatusInLatched_reg[7]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26591_,
		_w26592_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name16080 (
		_w26388_,
		_w26588_,
		_w26590_,
		_w26592_,
		_w26593_
	);
	LUT2 #(
		.INIT('h2)
	) name16081 (
		\wishbone_ram_di_reg[8]/NET0131 ,
		_w26389_,
		_w26594_
	);
	LUT2 #(
		.INIT('h8)
	) name16082 (
		\wishbone_TxEn_needed_reg/NET0131 ,
		\wishbone_TxUnderRun_reg/NET0131 ,
		_w26595_
	);
	LUT2 #(
		.INIT('h4)
	) name16083 (
		_w26382_,
		_w26595_,
		_w26596_
	);
	LUT4 #(
		.INIT('h002a)
	) name16084 (
		\wb_dat_i[8]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26597_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16085 (
		\wishbone_RxStatusInLatched_reg[8]/NET0131 ,
		_w26385_,
		_w26389_,
		_w26597_,
		_w26598_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name16086 (
		_w26388_,
		_w26594_,
		_w26596_,
		_w26598_,
		_w26599_
	);
	LUT3 #(
		.INIT('h4c)
	) name16087 (
		_w11866_,
		_w25827_,
		_w25829_,
		_w26600_
	);
	LUT3 #(
		.INIT('hb0)
	) name16088 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		_w26601_
	);
	LUT4 #(
		.INIT('hb34c)
	) name16089 (
		_w11866_,
		_w25827_,
		_w25829_,
		_w26601_,
		_w26602_
	);
	LUT3 #(
		.INIT('h07)
	) name16090 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		_w26603_
	);
	LUT2 #(
		.INIT('h2)
	) name16091 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		_w26604_
	);
	LUT3 #(
		.INIT('h13)
	) name16092 (
		_w25802_,
		_w26603_,
		_w26604_,
		_w26605_
	);
	LUT4 #(
		.INIT('h80cc)
	) name16093 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25385_,
		_w25802_,
		_w26083_,
		_w26606_
	);
	LUT3 #(
		.INIT('hea)
	) name16094 (
		_w26203_,
		_w26605_,
		_w26606_,
		_w26607_
	);
	LUT2 #(
		.INIT('h4)
	) name16095 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26608_
	);
	LUT4 #(
		.INIT('h00b0)
	) name16096 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_WriteRxDataToFifoSync2_reg/NET0131 ,
		\wishbone_WriteRxDataToFifoSync3_reg/NET0131 ,
		_w26609_
	);
	LUT2 #(
		.INIT('h2)
	) name16097 (
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26610_
	);
	LUT4 #(
		.INIT('h7000)
	) name16098 (
		_w11866_,
		_w25829_,
		_w26609_,
		_w26610_,
		_w26611_
	);
	LUT2 #(
		.INIT('h8)
	) name16099 (
		_w26608_,
		_w26611_,
		_w26612_
	);
	LUT4 #(
		.INIT('haccc)
	) name16100 (
		\wishbone_RxDataLatched2_reg[10]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[10][10]/P0001 ,
		_w26608_,
		_w26611_,
		_w26613_
	);
	LUT4 #(
		.INIT('haccc)
	) name16101 (
		\wishbone_RxDataLatched2_reg[12]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[10][12]/P0001 ,
		_w26608_,
		_w26611_,
		_w26614_
	);
	LUT4 #(
		.INIT('haccc)
	) name16102 (
		\wishbone_RxDataLatched2_reg[14]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[10][14]/P0001 ,
		_w26608_,
		_w26611_,
		_w26615_
	);
	LUT4 #(
		.INIT('haccc)
	) name16103 (
		\wishbone_RxDataLatched2_reg[16]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[10][16]/P0001 ,
		_w26608_,
		_w26611_,
		_w26616_
	);
	LUT4 #(
		.INIT('haccc)
	) name16104 (
		\wishbone_RxDataLatched2_reg[1]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[10][1]/P0001 ,
		_w26608_,
		_w26611_,
		_w26617_
	);
	LUT4 #(
		.INIT('haccc)
	) name16105 (
		\wishbone_RxDataLatched2_reg[20]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[10][20]/P0001 ,
		_w26608_,
		_w26611_,
		_w26618_
	);
	LUT4 #(
		.INIT('haccc)
	) name16106 (
		\wishbone_RxDataLatched2_reg[27]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[10][27]/P0001 ,
		_w26608_,
		_w26611_,
		_w26619_
	);
	LUT4 #(
		.INIT('haccc)
	) name16107 (
		\wishbone_RxDataLatched2_reg[28]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[10][28]/P0001 ,
		_w26608_,
		_w26611_,
		_w26620_
	);
	LUT4 #(
		.INIT('haccc)
	) name16108 (
		\wishbone_RxDataLatched2_reg[29]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[10][29]/P0001 ,
		_w26608_,
		_w26611_,
		_w26621_
	);
	LUT4 #(
		.INIT('haccc)
	) name16109 (
		\wishbone_RxDataLatched2_reg[31]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[10][31]/P0001 ,
		_w26608_,
		_w26611_,
		_w26622_
	);
	LUT4 #(
		.INIT('haccc)
	) name16110 (
		\wishbone_RxDataLatched2_reg[4]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[10][4]/P0001 ,
		_w26608_,
		_w26611_,
		_w26623_
	);
	LUT4 #(
		.INIT('haccc)
	) name16111 (
		\wishbone_RxDataLatched2_reg[5]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[10][5]/P0001 ,
		_w26608_,
		_w26611_,
		_w26624_
	);
	LUT4 #(
		.INIT('haccc)
	) name16112 (
		\wishbone_RxDataLatched2_reg[7]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[10][7]/P0001 ,
		_w26608_,
		_w26611_,
		_w26625_
	);
	LUT4 #(
		.INIT('haccc)
	) name16113 (
		\wishbone_RxDataLatched2_reg[9]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[10][9]/P0001 ,
		_w26608_,
		_w26611_,
		_w26626_
	);
	LUT3 #(
		.INIT('h20)
	) name16114 (
		\wishbone_WriteRxDataToFifoSync2_reg/NET0131 ,
		\wishbone_WriteRxDataToFifoSync3_reg/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26627_
	);
	LUT4 #(
		.INIT('h1300)
	) name16115 (
		_w11866_,
		_w24970_,
		_w25829_,
		_w26627_,
		_w26628_
	);
	LUT3 #(
		.INIT('h10)
	) name16116 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26629_
	);
	LUT2 #(
		.INIT('h8)
	) name16117 (
		_w26628_,
		_w26629_,
		_w26630_
	);
	LUT4 #(
		.INIT('h0200)
	) name16118 (
		\wishbone_RxDataLatched2_reg[11]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26631_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16119 (
		\wishbone_rx_fifo_fifo_reg[12][11]/P0001 ,
		_w26628_,
		_w26629_,
		_w26631_,
		_w26632_
	);
	LUT4 #(
		.INIT('h0200)
	) name16120 (
		\wishbone_RxDataLatched2_reg[12]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26633_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16121 (
		\wishbone_rx_fifo_fifo_reg[12][12]/P0001 ,
		_w26628_,
		_w26629_,
		_w26633_,
		_w26634_
	);
	LUT4 #(
		.INIT('h0200)
	) name16122 (
		\wishbone_RxDataLatched2_reg[14]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26635_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16123 (
		\wishbone_rx_fifo_fifo_reg[12][14]/P0001 ,
		_w26628_,
		_w26629_,
		_w26635_,
		_w26636_
	);
	LUT4 #(
		.INIT('h0200)
	) name16124 (
		\wishbone_RxDataLatched2_reg[15]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26637_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16125 (
		\wishbone_rx_fifo_fifo_reg[12][15]/P0001 ,
		_w26628_,
		_w26629_,
		_w26637_,
		_w26638_
	);
	LUT4 #(
		.INIT('h0200)
	) name16126 (
		\wishbone_RxDataLatched2_reg[16]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26639_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16127 (
		\wishbone_rx_fifo_fifo_reg[12][16]/P0001 ,
		_w26628_,
		_w26629_,
		_w26639_,
		_w26640_
	);
	LUT4 #(
		.INIT('h0200)
	) name16128 (
		\wishbone_RxDataLatched2_reg[17]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26641_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16129 (
		\wishbone_rx_fifo_fifo_reg[12][17]/P0001 ,
		_w26628_,
		_w26629_,
		_w26641_,
		_w26642_
	);
	LUT4 #(
		.INIT('h0200)
	) name16130 (
		\wishbone_RxDataLatched2_reg[19]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26643_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16131 (
		\wishbone_rx_fifo_fifo_reg[12][19]/P0001 ,
		_w26628_,
		_w26629_,
		_w26643_,
		_w26644_
	);
	LUT4 #(
		.INIT('h0200)
	) name16132 (
		\wishbone_RxDataLatched2_reg[21]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26645_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16133 (
		\wishbone_rx_fifo_fifo_reg[12][21]/P0001 ,
		_w26628_,
		_w26629_,
		_w26645_,
		_w26646_
	);
	LUT4 #(
		.INIT('h0200)
	) name16134 (
		\wishbone_RxDataLatched2_reg[22]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26647_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16135 (
		\wishbone_rx_fifo_fifo_reg[12][22]/P0001 ,
		_w26628_,
		_w26629_,
		_w26647_,
		_w26648_
	);
	LUT4 #(
		.INIT('h0200)
	) name16136 (
		\wishbone_RxDataLatched2_reg[23]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26649_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16137 (
		\wishbone_rx_fifo_fifo_reg[12][23]/P0001 ,
		_w26628_,
		_w26629_,
		_w26649_,
		_w26650_
	);
	LUT4 #(
		.INIT('h0200)
	) name16138 (
		\wishbone_RxDataLatched2_reg[24]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26651_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16139 (
		\wishbone_rx_fifo_fifo_reg[12][24]/P0001 ,
		_w26628_,
		_w26629_,
		_w26651_,
		_w26652_
	);
	LUT4 #(
		.INIT('h0200)
	) name16140 (
		\wishbone_RxDataLatched2_reg[27]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26653_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16141 (
		\wishbone_rx_fifo_fifo_reg[12][27]/P0001 ,
		_w26628_,
		_w26629_,
		_w26653_,
		_w26654_
	);
	LUT4 #(
		.INIT('h0200)
	) name16142 (
		\wishbone_RxDataLatched2_reg[28]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26655_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16143 (
		\wishbone_rx_fifo_fifo_reg[12][28]/P0001 ,
		_w26628_,
		_w26629_,
		_w26655_,
		_w26656_
	);
	LUT4 #(
		.INIT('h0200)
	) name16144 (
		\wishbone_RxDataLatched2_reg[31]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26657_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16145 (
		\wishbone_rx_fifo_fifo_reg[12][31]/P0001 ,
		_w26628_,
		_w26629_,
		_w26657_,
		_w26658_
	);
	LUT4 #(
		.INIT('h0200)
	) name16146 (
		\wishbone_RxDataLatched2_reg[4]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26659_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16147 (
		\wishbone_rx_fifo_fifo_reg[12][4]/P0001 ,
		_w26628_,
		_w26629_,
		_w26659_,
		_w26660_
	);
	LUT4 #(
		.INIT('h0200)
	) name16148 (
		\wishbone_RxDataLatched2_reg[7]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26661_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16149 (
		\wishbone_rx_fifo_fifo_reg[12][7]/P0001 ,
		_w26628_,
		_w26629_,
		_w26661_,
		_w26662_
	);
	LUT2 #(
		.INIT('h2)
	) name16150 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26663_
	);
	LUT2 #(
		.INIT('h8)
	) name16151 (
		_w26611_,
		_w26663_,
		_w26664_
	);
	LUT4 #(
		.INIT('haccc)
	) name16152 (
		\wishbone_RxDataLatched2_reg[10]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][10]/P0001 ,
		_w26611_,
		_w26663_,
		_w26665_
	);
	LUT4 #(
		.INIT('haccc)
	) name16153 (
		\wishbone_RxDataLatched2_reg[12]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][12]/P0001 ,
		_w26611_,
		_w26663_,
		_w26666_
	);
	LUT4 #(
		.INIT('haccc)
	) name16154 (
		\wishbone_RxDataLatched2_reg[13]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][13]/P0001 ,
		_w26611_,
		_w26663_,
		_w26667_
	);
	LUT4 #(
		.INIT('haccc)
	) name16155 (
		\wishbone_RxDataLatched2_reg[14]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][14]/P0001 ,
		_w26611_,
		_w26663_,
		_w26668_
	);
	LUT4 #(
		.INIT('haccc)
	) name16156 (
		\wishbone_RxDataLatched2_reg[18]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][18]/P0001 ,
		_w26611_,
		_w26663_,
		_w26669_
	);
	LUT4 #(
		.INIT('haccc)
	) name16157 (
		\wishbone_RxDataLatched2_reg[19]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][19]/P0001 ,
		_w26611_,
		_w26663_,
		_w26670_
	);
	LUT4 #(
		.INIT('haccc)
	) name16158 (
		\wishbone_RxDataLatched2_reg[24]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][24]/P0001 ,
		_w26611_,
		_w26663_,
		_w26671_
	);
	LUT4 #(
		.INIT('haccc)
	) name16159 (
		\wishbone_RxDataLatched2_reg[26]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][26]/P0001 ,
		_w26611_,
		_w26663_,
		_w26672_
	);
	LUT4 #(
		.INIT('haccc)
	) name16160 (
		\wishbone_RxDataLatched2_reg[29]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][29]/P0001 ,
		_w26611_,
		_w26663_,
		_w26673_
	);
	LUT4 #(
		.INIT('haccc)
	) name16161 (
		\wishbone_RxDataLatched2_reg[28]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][28]/P0001 ,
		_w26611_,
		_w26663_,
		_w26674_
	);
	LUT4 #(
		.INIT('haccc)
	) name16162 (
		\wishbone_RxDataLatched2_reg[2]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][2]/P0001 ,
		_w26611_,
		_w26663_,
		_w26675_
	);
	LUT4 #(
		.INIT('haccc)
	) name16163 (
		\wishbone_RxDataLatched2_reg[30]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][30]/P0001 ,
		_w26611_,
		_w26663_,
		_w26676_
	);
	LUT4 #(
		.INIT('haccc)
	) name16164 (
		\wishbone_RxDataLatched2_reg[31]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][31]/P0001 ,
		_w26611_,
		_w26663_,
		_w26677_
	);
	LUT4 #(
		.INIT('haccc)
	) name16165 (
		\wishbone_RxDataLatched2_reg[4]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][4]/P0001 ,
		_w26611_,
		_w26663_,
		_w26678_
	);
	LUT4 #(
		.INIT('haccc)
	) name16166 (
		\wishbone_RxDataLatched2_reg[7]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][7]/P0001 ,
		_w26611_,
		_w26663_,
		_w26679_
	);
	LUT4 #(
		.INIT('haccc)
	) name16167 (
		\wishbone_RxDataLatched2_reg[8]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][8]/P0001 ,
		_w26611_,
		_w26663_,
		_w26680_
	);
	LUT4 #(
		.INIT('haccc)
	) name16168 (
		\wishbone_RxDataLatched2_reg[9]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[3][9]/P0001 ,
		_w26611_,
		_w26663_,
		_w26681_
	);
	LUT3 #(
		.INIT('h02)
	) name16169 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26682_
	);
	LUT2 #(
		.INIT('h8)
	) name16170 (
		_w26628_,
		_w26682_,
		_w26683_
	);
	LUT4 #(
		.INIT('h0008)
	) name16171 (
		\wishbone_RxDataLatched2_reg[10]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26684_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16172 (
		\wishbone_rx_fifo_fifo_reg[5][10]/P0001 ,
		_w26628_,
		_w26682_,
		_w26684_,
		_w26685_
	);
	LUT4 #(
		.INIT('h0008)
	) name16173 (
		\wishbone_RxDataLatched2_reg[13]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26686_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16174 (
		\wishbone_rx_fifo_fifo_reg[5][13]/P0001 ,
		_w26628_,
		_w26682_,
		_w26686_,
		_w26687_
	);
	LUT4 #(
		.INIT('h0008)
	) name16175 (
		\wishbone_RxDataLatched2_reg[15]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26688_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16176 (
		\wishbone_rx_fifo_fifo_reg[5][15]/P0001 ,
		_w26628_,
		_w26682_,
		_w26688_,
		_w26689_
	);
	LUT4 #(
		.INIT('h0008)
	) name16177 (
		\wishbone_RxDataLatched2_reg[17]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26690_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16178 (
		\wishbone_rx_fifo_fifo_reg[5][17]/P0001 ,
		_w26628_,
		_w26682_,
		_w26690_,
		_w26691_
	);
	LUT4 #(
		.INIT('h0008)
	) name16179 (
		\wishbone_RxDataLatched2_reg[19]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26692_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16180 (
		\wishbone_rx_fifo_fifo_reg[5][19]/P0001 ,
		_w26628_,
		_w26682_,
		_w26692_,
		_w26693_
	);
	LUT4 #(
		.INIT('h0008)
	) name16181 (
		\wishbone_RxDataLatched2_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26694_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16182 (
		\wishbone_rx_fifo_fifo_reg[5][1]/P0001 ,
		_w26628_,
		_w26682_,
		_w26694_,
		_w26695_
	);
	LUT4 #(
		.INIT('h0008)
	) name16183 (
		\wishbone_RxDataLatched2_reg[21]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26696_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16184 (
		\wishbone_rx_fifo_fifo_reg[5][21]/P0001 ,
		_w26628_,
		_w26682_,
		_w26696_,
		_w26697_
	);
	LUT4 #(
		.INIT('h0008)
	) name16185 (
		\wishbone_RxDataLatched2_reg[22]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26698_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16186 (
		\wishbone_rx_fifo_fifo_reg[5][22]/P0001 ,
		_w26628_,
		_w26682_,
		_w26698_,
		_w26699_
	);
	LUT4 #(
		.INIT('h0008)
	) name16187 (
		\wishbone_RxDataLatched2_reg[20]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26700_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16188 (
		\wishbone_rx_fifo_fifo_reg[5][20]/P0001 ,
		_w26628_,
		_w26682_,
		_w26700_,
		_w26701_
	);
	LUT4 #(
		.INIT('h0008)
	) name16189 (
		\wishbone_RxDataLatched2_reg[23]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26702_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16190 (
		\wishbone_rx_fifo_fifo_reg[5][23]/P0001 ,
		_w26628_,
		_w26682_,
		_w26702_,
		_w26703_
	);
	LUT4 #(
		.INIT('h0008)
	) name16191 (
		\wishbone_RxDataLatched2_reg[24]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26704_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16192 (
		\wishbone_rx_fifo_fifo_reg[5][24]/P0001 ,
		_w26628_,
		_w26682_,
		_w26704_,
		_w26705_
	);
	LUT4 #(
		.INIT('h0008)
	) name16193 (
		\wishbone_RxDataLatched2_reg[26]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26706_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16194 (
		\wishbone_rx_fifo_fifo_reg[5][26]/P0001 ,
		_w26628_,
		_w26682_,
		_w26706_,
		_w26707_
	);
	LUT4 #(
		.INIT('h0008)
	) name16195 (
		\wishbone_RxDataLatched2_reg[28]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26708_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16196 (
		\wishbone_rx_fifo_fifo_reg[5][28]/P0001 ,
		_w26628_,
		_w26682_,
		_w26708_,
		_w26709_
	);
	LUT4 #(
		.INIT('h0008)
	) name16197 (
		\wishbone_RxDataLatched2_reg[3]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26710_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16198 (
		\wishbone_rx_fifo_fifo_reg[5][3]/P0001 ,
		_w26628_,
		_w26682_,
		_w26710_,
		_w26711_
	);
	LUT4 #(
		.INIT('h0008)
	) name16199 (
		\wishbone_RxDataLatched2_reg[6]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26712_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16200 (
		\wishbone_rx_fifo_fifo_reg[5][6]/P0001 ,
		_w26628_,
		_w26682_,
		_w26712_,
		_w26713_
	);
	LUT4 #(
		.INIT('h0008)
	) name16201 (
		\wishbone_RxDataLatched2_reg[8]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26714_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16202 (
		\wishbone_rx_fifo_fifo_reg[5][8]/P0001 ,
		_w26628_,
		_w26682_,
		_w26714_,
		_w26715_
	);
	LUT2 #(
		.INIT('h1)
	) name16203 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26716_
	);
	LUT3 #(
		.INIT('h04)
	) name16204 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26717_
	);
	LUT2 #(
		.INIT('h8)
	) name16205 (
		_w26628_,
		_w26717_,
		_w26718_
	);
	LUT4 #(
		.INIT('h0020)
	) name16206 (
		\wishbone_RxDataLatched2_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26719_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16207 (
		\wishbone_rx_fifo_fifo_reg[6][0]/P0001 ,
		_w26628_,
		_w26717_,
		_w26719_,
		_w26720_
	);
	LUT4 #(
		.INIT('h0020)
	) name16208 (
		\wishbone_RxDataLatched2_reg[10]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26721_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16209 (
		\wishbone_rx_fifo_fifo_reg[6][10]/P0001 ,
		_w26628_,
		_w26717_,
		_w26721_,
		_w26722_
	);
	LUT4 #(
		.INIT('h0020)
	) name16210 (
		\wishbone_RxDataLatched2_reg[11]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26723_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16211 (
		\wishbone_rx_fifo_fifo_reg[6][11]/P0001 ,
		_w26628_,
		_w26717_,
		_w26723_,
		_w26724_
	);
	LUT4 #(
		.INIT('h0020)
	) name16212 (
		\wishbone_RxDataLatched2_reg[14]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26725_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16213 (
		\wishbone_rx_fifo_fifo_reg[6][14]/P0001 ,
		_w26628_,
		_w26717_,
		_w26725_,
		_w26726_
	);
	LUT4 #(
		.INIT('h0020)
	) name16214 (
		\wishbone_RxDataLatched2_reg[15]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26727_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16215 (
		\wishbone_rx_fifo_fifo_reg[6][15]/P0001 ,
		_w26628_,
		_w26717_,
		_w26727_,
		_w26728_
	);
	LUT4 #(
		.INIT('h0020)
	) name16216 (
		\wishbone_RxDataLatched2_reg[16]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26729_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16217 (
		\wishbone_rx_fifo_fifo_reg[6][16]/P0001 ,
		_w26628_,
		_w26717_,
		_w26729_,
		_w26730_
	);
	LUT4 #(
		.INIT('h0020)
	) name16218 (
		\wishbone_RxDataLatched2_reg[18]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26731_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16219 (
		\wishbone_rx_fifo_fifo_reg[6][18]/P0001 ,
		_w26628_,
		_w26717_,
		_w26731_,
		_w26732_
	);
	LUT4 #(
		.INIT('h0020)
	) name16220 (
		\wishbone_RxDataLatched2_reg[19]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26733_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16221 (
		\wishbone_rx_fifo_fifo_reg[6][19]/P0001 ,
		_w26628_,
		_w26717_,
		_w26733_,
		_w26734_
	);
	LUT4 #(
		.INIT('h0020)
	) name16222 (
		\wishbone_RxDataLatched2_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26735_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16223 (
		\wishbone_rx_fifo_fifo_reg[6][1]/P0001 ,
		_w26628_,
		_w26717_,
		_w26735_,
		_w26736_
	);
	LUT4 #(
		.INIT('h0020)
	) name16224 (
		\wishbone_RxDataLatched2_reg[21]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26737_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16225 (
		\wishbone_rx_fifo_fifo_reg[6][21]/P0001 ,
		_w26628_,
		_w26717_,
		_w26737_,
		_w26738_
	);
	LUT4 #(
		.INIT('h0020)
	) name16226 (
		\wishbone_RxDataLatched2_reg[22]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26739_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16227 (
		\wishbone_rx_fifo_fifo_reg[6][22]/P0001 ,
		_w26628_,
		_w26717_,
		_w26739_,
		_w26740_
	);
	LUT4 #(
		.INIT('h0020)
	) name16228 (
		\wishbone_RxDataLatched2_reg[23]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26741_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16229 (
		\wishbone_rx_fifo_fifo_reg[6][23]/P0001 ,
		_w26628_,
		_w26717_,
		_w26741_,
		_w26742_
	);
	LUT4 #(
		.INIT('h0020)
	) name16230 (
		\wishbone_RxDataLatched2_reg[25]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26743_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16231 (
		\wishbone_rx_fifo_fifo_reg[6][25]/P0001 ,
		_w26628_,
		_w26717_,
		_w26743_,
		_w26744_
	);
	LUT4 #(
		.INIT('h0020)
	) name16232 (
		\wishbone_RxDataLatched2_reg[26]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26745_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16233 (
		\wishbone_rx_fifo_fifo_reg[6][26]/P0001 ,
		_w26628_,
		_w26717_,
		_w26745_,
		_w26746_
	);
	LUT4 #(
		.INIT('h0020)
	) name16234 (
		\wishbone_RxDataLatched2_reg[24]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26747_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16235 (
		\wishbone_rx_fifo_fifo_reg[6][24]/P0001 ,
		_w26628_,
		_w26717_,
		_w26747_,
		_w26748_
	);
	LUT4 #(
		.INIT('h0020)
	) name16236 (
		\wishbone_RxDataLatched2_reg[27]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26749_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16237 (
		\wishbone_rx_fifo_fifo_reg[6][27]/P0001 ,
		_w26628_,
		_w26717_,
		_w26749_,
		_w26750_
	);
	LUT4 #(
		.INIT('h0020)
	) name16238 (
		\wishbone_RxDataLatched2_reg[28]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26751_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16239 (
		\wishbone_rx_fifo_fifo_reg[6][28]/P0001 ,
		_w26628_,
		_w26717_,
		_w26751_,
		_w26752_
	);
	LUT4 #(
		.INIT('h0020)
	) name16240 (
		\wishbone_RxDataLatched2_reg[2]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26753_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16241 (
		\wishbone_rx_fifo_fifo_reg[6][2]/P0001 ,
		_w26628_,
		_w26717_,
		_w26753_,
		_w26754_
	);
	LUT4 #(
		.INIT('h0020)
	) name16242 (
		\wishbone_RxDataLatched2_reg[31]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26755_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16243 (
		\wishbone_rx_fifo_fifo_reg[6][31]/P0001 ,
		_w26628_,
		_w26717_,
		_w26755_,
		_w26756_
	);
	LUT4 #(
		.INIT('h0020)
	) name16244 (
		\wishbone_RxDataLatched2_reg[5]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26757_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16245 (
		\wishbone_rx_fifo_fifo_reg[6][5]/P0001 ,
		_w26628_,
		_w26717_,
		_w26757_,
		_w26758_
	);
	LUT4 #(
		.INIT('h0020)
	) name16246 (
		\wishbone_RxDataLatched2_reg[6]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26759_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16247 (
		\wishbone_rx_fifo_fifo_reg[6][6]/P0001 ,
		_w26628_,
		_w26717_,
		_w26759_,
		_w26760_
	);
	LUT4 #(
		.INIT('h0020)
	) name16248 (
		\wishbone_RxDataLatched2_reg[7]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26761_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16249 (
		\wishbone_rx_fifo_fifo_reg[6][7]/P0001 ,
		_w26628_,
		_w26717_,
		_w26761_,
		_w26762_
	);
	LUT4 #(
		.INIT('h0020)
	) name16250 (
		\wishbone_RxDataLatched2_reg[9]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26763_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16251 (
		\wishbone_rx_fifo_fifo_reg[6][9]/P0001 ,
		_w26628_,
		_w26717_,
		_w26763_,
		_w26764_
	);
	LUT4 #(
		.INIT('h0002)
	) name16252 (
		\wishbone_WriteRxDataToFifoSync2_reg/NET0131 ,
		\wishbone_WriteRxDataToFifoSync3_reg/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26765_
	);
	LUT2 #(
		.INIT('h8)
	) name16253 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26766_
	);
	LUT4 #(
		.INIT('hb000)
	) name16254 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26767_
	);
	LUT4 #(
		.INIT('h7000)
	) name16255 (
		_w11866_,
		_w25829_,
		_w26765_,
		_w26767_,
		_w26768_
	);
	LUT3 #(
		.INIT('hac)
	) name16256 (
		\wishbone_RxDataLatched2_reg[0]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][0]/P0001 ,
		_w26768_,
		_w26769_
	);
	LUT3 #(
		.INIT('hac)
	) name16257 (
		\wishbone_RxDataLatched2_reg[10]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][10]/P0001 ,
		_w26768_,
		_w26770_
	);
	LUT3 #(
		.INIT('hac)
	) name16258 (
		\wishbone_RxDataLatched2_reg[11]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][11]/P0001 ,
		_w26768_,
		_w26771_
	);
	LUT3 #(
		.INIT('hac)
	) name16259 (
		\wishbone_RxDataLatched2_reg[13]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][13]/P0001 ,
		_w26768_,
		_w26772_
	);
	LUT3 #(
		.INIT('hac)
	) name16260 (
		\wishbone_RxDataLatched2_reg[16]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][16]/P0001 ,
		_w26768_,
		_w26773_
	);
	LUT3 #(
		.INIT('hac)
	) name16261 (
		\wishbone_RxDataLatched2_reg[17]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][17]/P0001 ,
		_w26768_,
		_w26774_
	);
	LUT3 #(
		.INIT('hac)
	) name16262 (
		\wishbone_RxDataLatched2_reg[18]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][18]/P0001 ,
		_w26768_,
		_w26775_
	);
	LUT3 #(
		.INIT('hac)
	) name16263 (
		\wishbone_RxDataLatched2_reg[19]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][19]/P0001 ,
		_w26768_,
		_w26776_
	);
	LUT3 #(
		.INIT('hac)
	) name16264 (
		\wishbone_RxDataLatched2_reg[1]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][1]/P0001 ,
		_w26768_,
		_w26777_
	);
	LUT3 #(
		.INIT('hac)
	) name16265 (
		\wishbone_RxDataLatched2_reg[20]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][20]/P0001 ,
		_w26768_,
		_w26778_
	);
	LUT3 #(
		.INIT('hac)
	) name16266 (
		\wishbone_RxDataLatched2_reg[21]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][21]/P0001 ,
		_w26768_,
		_w26779_
	);
	LUT3 #(
		.INIT('hac)
	) name16267 (
		\wishbone_RxDataLatched2_reg[22]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][22]/P0001 ,
		_w26768_,
		_w26780_
	);
	LUT3 #(
		.INIT('hac)
	) name16268 (
		\wishbone_RxDataLatched2_reg[23]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][23]/P0001 ,
		_w26768_,
		_w26781_
	);
	LUT3 #(
		.INIT('hac)
	) name16269 (
		\wishbone_RxDataLatched2_reg[24]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][24]/P0001 ,
		_w26768_,
		_w26782_
	);
	LUT3 #(
		.INIT('hac)
	) name16270 (
		\wishbone_RxDataLatched2_reg[25]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][25]/P0001 ,
		_w26768_,
		_w26783_
	);
	LUT3 #(
		.INIT('hac)
	) name16271 (
		\wishbone_RxDataLatched2_reg[26]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][26]/P0001 ,
		_w26768_,
		_w26784_
	);
	LUT3 #(
		.INIT('hac)
	) name16272 (
		\wishbone_RxDataLatched2_reg[27]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][27]/P0001 ,
		_w26768_,
		_w26785_
	);
	LUT3 #(
		.INIT('hac)
	) name16273 (
		\wishbone_RxDataLatched2_reg[29]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][29]/P0001 ,
		_w26768_,
		_w26786_
	);
	LUT3 #(
		.INIT('hac)
	) name16274 (
		\wishbone_RxDataLatched2_reg[2]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][2]/P0001 ,
		_w26768_,
		_w26787_
	);
	LUT3 #(
		.INIT('hac)
	) name16275 (
		\wishbone_RxDataLatched2_reg[30]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][30]/P0001 ,
		_w26768_,
		_w26788_
	);
	LUT3 #(
		.INIT('hac)
	) name16276 (
		\wishbone_RxDataLatched2_reg[4]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][4]/P0001 ,
		_w26768_,
		_w26789_
	);
	LUT3 #(
		.INIT('hac)
	) name16277 (
		\wishbone_RxDataLatched2_reg[5]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][5]/P0001 ,
		_w26768_,
		_w26790_
	);
	LUT3 #(
		.INIT('hac)
	) name16278 (
		\wishbone_RxDataLatched2_reg[7]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][7]/P0001 ,
		_w26768_,
		_w26791_
	);
	LUT3 #(
		.INIT('hac)
	) name16279 (
		\wishbone_RxDataLatched2_reg[9]/NET0131 ,
		\wishbone_rx_fifo_fifo_reg[9][9]/P0001 ,
		_w26768_,
		_w26792_
	);
	LUT3 #(
		.INIT('h10)
	) name16280 (
		\wishbone_TxAbortPacket_reg/NET0131 ,
		\wishbone_TxRetryPacket_reg/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[0]/NET0131 ,
		_w26793_
	);
	LUT2 #(
		.INIT('h9)
	) name16281 (
		_w25799_,
		_w26793_,
		_w26794_
	);
	LUT4 #(
		.INIT('h0001)
	) name16282 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26795_
	);
	LUT2 #(
		.INIT('h1)
	) name16283 (
		_w24970_,
		_w26795_,
		_w26796_
	);
	LUT2 #(
		.INIT('h2)
	) name16284 (
		_w26600_,
		_w26796_,
		_w26797_
	);
	LUT2 #(
		.INIT('h8)
	) name16285 (
		_w26611_,
		_w26766_,
		_w26798_
	);
	LUT3 #(
		.INIT('h20)
	) name16286 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26799_
	);
	LUT2 #(
		.INIT('h8)
	) name16287 (
		_w26628_,
		_w26799_,
		_w26800_
	);
	LUT3 #(
		.INIT('h40)
	) name16288 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26801_
	);
	LUT2 #(
		.INIT('h8)
	) name16289 (
		_w26628_,
		_w26801_,
		_w26802_
	);
	LUT3 #(
		.INIT('h80)
	) name16290 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26803_
	);
	LUT2 #(
		.INIT('h8)
	) name16291 (
		_w26628_,
		_w26803_,
		_w26804_
	);
	LUT4 #(
		.INIT('h00b0)
	) name16292 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26805_
	);
	LUT4 #(
		.INIT('h7000)
	) name16293 (
		_w11866_,
		_w25829_,
		_w26765_,
		_w26805_,
		_w26806_
	);
	LUT2 #(
		.INIT('h8)
	) name16294 (
		_w26611_,
		_w26716_,
		_w26807_
	);
	LUT3 #(
		.INIT('h01)
	) name16295 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26808_
	);
	LUT2 #(
		.INIT('h8)
	) name16296 (
		_w26628_,
		_w26808_,
		_w26809_
	);
	LUT3 #(
		.INIT('h08)
	) name16297 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26810_
	);
	LUT2 #(
		.INIT('h8)
	) name16298 (
		_w26628_,
		_w26810_,
		_w26811_
	);
	LUT4 #(
		.INIT('h0100)
	) name16299 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26812_
	);
	LUT4 #(
		.INIT('h7000)
	) name16300 (
		_w11866_,
		_w25829_,
		_w26609_,
		_w26812_,
		_w26813_
	);
	LUT4 #(
		.INIT('h222a)
	) name16301 (
		\miim1_LatchByte_reg[0]/NET0131 ,
		_w24568_,
		_w24572_,
		_w24573_,
		_w26814_
	);
	LUT4 #(
		.INIT('h0200)
	) name16302 (
		_w24561_,
		_w24567_,
		_w24571_,
		_w26814_,
		_w26815_
	);
	LUT3 #(
		.INIT('h10)
	) name16303 (
		\wishbone_TxAbortPacket_reg/NET0131 ,
		\wishbone_TxRetryPacket_reg/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		_w26816_
	);
	LUT4 #(
		.INIT('hd52a)
	) name16304 (
		_w25792_,
		_w25795_,
		_w25796_,
		_w26816_,
		_w26817_
	);
	LUT3 #(
		.INIT('h6c)
	) name16305 (
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		_w11135_,
		_w26818_
	);
	LUT4 #(
		.INIT('h0200)
	) name16306 (
		\ethreg1_TXCTRL_1_DataOut_reg[7]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26819_
	);
	LUT4 #(
		.INIT('h00e0)
	) name16307 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26820_
	);
	LUT3 #(
		.INIT('ha8)
	) name16308 (
		_w26365_,
		_w26819_,
		_w26820_,
		_w26821_
	);
	LUT3 #(
		.INIT('heb)
	) name16309 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w26822_
	);
	LUT2 #(
		.INIT('h2)
	) name16310 (
		_w26366_,
		_w26822_,
		_w26823_
	);
	LUT4 #(
		.INIT('h0200)
	) name16311 (
		\ethreg1_TXCTRL_0_DataOut_reg[7]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26824_
	);
	LUT4 #(
		.INIT('h0008)
	) name16312 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26825_
	);
	LUT4 #(
		.INIT('h135f)
	) name16313 (
		_w25925_,
		_w26359_,
		_w26824_,
		_w26825_,
		_w26826_
	);
	LUT4 #(
		.INIT('h0008)
	) name16314 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26827_
	);
	LUT4 #(
		.INIT('h0200)
	) name16315 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w26828_
	);
	LUT4 #(
		.INIT('h153f)
	) name16316 (
		_w26361_,
		_w26370_,
		_w26827_,
		_w26828_,
		_w26829_
	);
	LUT4 #(
		.INIT('h0020)
	) name16317 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w26830_
	);
	LUT4 #(
		.INIT('h0020)
	) name16318 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26831_
	);
	LUT4 #(
		.INIT('h135f)
	) name16319 (
		_w26361_,
		_w26370_,
		_w26830_,
		_w26831_,
		_w26832_
	);
	LUT4 #(
		.INIT('h4000)
	) name16320 (
		_w26823_,
		_w26826_,
		_w26829_,
		_w26832_,
		_w26833_
	);
	LUT2 #(
		.INIT('hb)
	) name16321 (
		_w26821_,
		_w26833_,
		_w26834_
	);
	LUT4 #(
		.INIT('h8000)
	) name16322 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		_w26835_
	);
	LUT4 #(
		.INIT('h2a00)
	) name16323 (
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		_w11866_,
		_w11867_,
		_w26835_,
		_w26836_
	);
	LUT3 #(
		.INIT('h12)
	) name16324 (
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w24970_,
		_w26836_,
		_w26837_
	);
	LUT4 #(
		.INIT('h008f)
	) name16325 (
		_w25795_,
		_w25796_,
		_w25798_,
		_w25800_,
		_w26838_
	);
	LUT4 #(
		.INIT('h0303)
	) name16326 (
		\wishbone_tx_fifo_cnt_reg[2]/NET0131 ,
		_w25793_,
		_w25794_,
		_w25797_,
		_w26839_
	);
	LUT4 #(
		.INIT('h8884)
	) name16327 (
		\wishbone_tx_fifo_cnt_reg[2]/NET0131 ,
		_w25385_,
		_w26838_,
		_w26839_,
		_w26840_
	);
	LUT3 #(
		.INIT('h0d)
	) name16328 (
		\wishbone_ReadTxDataFromFifo_sync2_reg/NET0131 ,
		\wishbone_ReadTxDataFromFifo_sync3_reg/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		_w26841_
	);
	LUT3 #(
		.INIT('h01)
	) name16329 (
		\wishbone_tx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		_w26842_
	);
	LUT3 #(
		.INIT('h13)
	) name16330 (
		_w25795_,
		_w26841_,
		_w26842_,
		_w26843_
	);
	LUT4 #(
		.INIT('h2002)
	) name16331 (
		\wishbone_ReadTxDataFromFifo_sync2_reg/NET0131 ,
		\wishbone_ReadTxDataFromFifo_sync3_reg/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		_w26844_
	);
	LUT4 #(
		.INIT('h80aa)
	) name16332 (
		_w25385_,
		_w25795_,
		_w25796_,
		_w26844_,
		_w26845_
	);
	LUT2 #(
		.INIT('h8)
	) name16333 (
		_w26843_,
		_w26845_,
		_w26846_
	);
	LUT3 #(
		.INIT('h20)
	) name16334 (
		\wishbone_ReadTxDataFromFifo_sync2_reg/NET0131 ,
		\wishbone_ReadTxDataFromFifo_sync3_reg/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		_w26847_
	);
	LUT4 #(
		.INIT('h2a00)
	) name16335 (
		_w25392_,
		_w25795_,
		_w25796_,
		_w26847_,
		_w26848_
	);
	LUT4 #(
		.INIT('h0888)
	) name16336 (
		_w25399_,
		_w25792_,
		_w25795_,
		_w25796_,
		_w26849_
	);
	LUT4 #(
		.INIT('h00c8)
	) name16337 (
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w25385_,
		_w26848_,
		_w26849_,
		_w26850_
	);
	LUT4 #(
		.INIT('h2000)
	) name16338 (
		\wishbone_WriteRxDataToFifoSync2_reg/NET0131 ,
		\wishbone_WriteRxDataToFifoSync3_reg/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		_w26851_
	);
	LUT3 #(
		.INIT('hb0)
	) name16339 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26852_
	);
	LUT4 #(
		.INIT('h8f00)
	) name16340 (
		_w11866_,
		_w25829_,
		_w26851_,
		_w26852_,
		_w26853_
	);
	LUT3 #(
		.INIT('h0b)
	) name16341 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26854_
	);
	LUT4 #(
		.INIT('h7000)
	) name16342 (
		_w11866_,
		_w25829_,
		_w26851_,
		_w26854_,
		_w26855_
	);
	LUT2 #(
		.INIT('he)
	) name16343 (
		_w26853_,
		_w26855_,
		_w26856_
	);
	LUT2 #(
		.INIT('h8)
	) name16344 (
		\wishbone_rx_fifo_write_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26857_
	);
	LUT4 #(
		.INIT('h7000)
	) name16345 (
		_w11866_,
		_w25829_,
		_w26851_,
		_w26857_,
		_w26858_
	);
	LUT3 #(
		.INIT('hb0)
	) name16346 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w26859_
	);
	LUT4 #(
		.INIT('h7000)
	) name16347 (
		_w11866_,
		_w25829_,
		_w26851_,
		_w26852_,
		_w26860_
	);
	LUT3 #(
		.INIT('h54)
	) name16348 (
		_w26858_,
		_w26859_,
		_w26860_,
		_w26861_
	);
	LUT3 #(
		.INIT('h10)
	) name16349 (
		\wishbone_TxAbortPacket_reg/NET0131 ,
		\wishbone_TxRetryPacket_reg/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26862_
	);
	LUT4 #(
		.INIT('h8f00)
	) name16350 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w26098_,
		_w26862_,
		_w26863_
	);
	LUT3 #(
		.INIT('h01)
	) name16351 (
		\wishbone_TxAbortPacket_reg/NET0131 ,
		\wishbone_TxRetryPacket_reg/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w26864_
	);
	LUT4 #(
		.INIT('h7000)
	) name16352 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w26098_,
		_w26864_,
		_w26865_
	);
	LUT2 #(
		.INIT('he)
	) name16353 (
		_w26863_,
		_w26865_,
		_w26866_
	);
	LUT4 #(
		.INIT('h4c00)
	) name16354 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w25802_,
		_w26098_,
		_w26867_
	);
	LUT3 #(
		.INIT('h48)
	) name16355 (
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w25385_,
		_w26867_,
		_w26868_
	);
	LUT2 #(
		.INIT('h2)
	) name16356 (
		\wishbone_TxEn_reg/NET0131 ,
		_w26389_,
		_w26869_
	);
	LUT3 #(
		.INIT('hba)
	) name16357 (
		_w26383_,
		_w26387_,
		_w26869_,
		_w26870_
	);
	LUT2 #(
		.INIT('h2)
	) name16358 (
		_w10519_,
		_w11580_,
		_w26871_
	);
	LUT3 #(
		.INIT('h70)
	) name16359 (
		_w10554_,
		_w10573_,
		_w26871_,
		_w26872_
	);
	LUT2 #(
		.INIT('h1)
	) name16360 (
		_w11390_,
		_w26872_,
		_w26873_
	);
	LUT3 #(
		.INIT('h20)
	) name16361 (
		\wishbone_WriteRxDataToFifoSync2_reg/NET0131 ,
		\wishbone_WriteRxDataToFifoSync3_reg/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		_w26874_
	);
	LUT4 #(
		.INIT('h4055)
	) name16362 (
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		_w11866_,
		_w25829_,
		_w26874_,
		_w26875_
	);
	LUT4 #(
		.INIT('h2033)
	) name16363 (
		_w11866_,
		_w24970_,
		_w25829_,
		_w26851_,
		_w26876_
	);
	LUT2 #(
		.INIT('h4)
	) name16364 (
		_w26875_,
		_w26876_,
		_w26877_
	);
	LUT2 #(
		.INIT('h6)
	) name16365 (
		\wishbone_tx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[1]/NET0131 ,
		_w26878_
	);
	LUT4 #(
		.INIT('h0070)
	) name16366 (
		_w25795_,
		_w25796_,
		_w25798_,
		_w26878_,
		_w26879_
	);
	LUT4 #(
		.INIT('hea00)
	) name16367 (
		_w25793_,
		_w25795_,
		_w25797_,
		_w26878_,
		_w26880_
	);
	LUT4 #(
		.INIT('h0007)
	) name16368 (
		\wishbone_tx_fifo_cnt_reg[1]/NET0131 ,
		_w25799_,
		_w26879_,
		_w26880_,
		_w26881_
	);
	LUT2 #(
		.INIT('h2)
	) name16369 (
		_w25385_,
		_w26881_,
		_w26882_
	);
	LUT4 #(
		.INIT('h2000)
	) name16370 (
		\wishbone_ReadTxDataFromFifo_sync2_reg/NET0131 ,
		\wishbone_ReadTxDataFromFifo_sync3_reg/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		_w26883_
	);
	LUT4 #(
		.INIT('h4055)
	) name16371 (
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		_w25795_,
		_w25796_,
		_w26883_,
		_w26884_
	);
	LUT3 #(
		.INIT('h02)
	) name16372 (
		_w25385_,
		_w26848_,
		_w26884_,
		_w26885_
	);
	LUT4 #(
		.INIT('h2033)
	) name16373 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		_w25802_,
		_w26083_,
		_w26886_
	);
	LUT4 #(
		.INIT('h80cc)
	) name16374 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25385_,
		_w25802_,
		_w26098_,
		_w26887_
	);
	LUT2 #(
		.INIT('h4)
	) name16375 (
		_w26886_,
		_w26887_,
		_w26888_
	);
	LUT2 #(
		.INIT('h2)
	) name16376 (
		\ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimerEq0_sync2_reg/NET0131 ,
		_w26889_
	);
	LUT2 #(
		.INIT('h7)
	) name16377 (
		_w11007_,
		_w11101_,
		_w26890_
	);
	LUT3 #(
		.INIT('h80)
	) name16378 (
		_w18757_,
		_w18758_,
		_w18794_,
		_w26891_
	);
	LUT4 #(
		.INIT('h4000)
	) name16379 (
		\wb_adr_i[11]_pad ,
		wb_cyc_i_pad,
		\wb_sel_i[2]_pad ,
		wb_stb_i_pad,
		_w26892_
	);
	LUT2 #(
		.INIT('h4)
	) name16380 (
		_w18750_,
		_w26892_,
		_w26893_
	);
	LUT3 #(
		.INIT('h40)
	) name16381 (
		_w18750_,
		_w24752_,
		_w26892_,
		_w26894_
	);
	LUT3 #(
		.INIT('h15)
	) name16382 (
		\ethreg1_TXCTRL_2_DataOut_reg[0]/NET0131 ,
		_w26891_,
		_w26894_,
		_w26895_
	);
	LUT4 #(
		.INIT('h0004)
	) name16383 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		\wb_dat_i[16]_pad ,
		_w26896_
	);
	LUT3 #(
		.INIT('h80)
	) name16384 (
		_w18757_,
		_w18758_,
		_w26896_,
		_w26897_
	);
	LUT3 #(
		.INIT('h15)
	) name16385 (
		\RstTxPauseRq_reg/NET0131 ,
		_w26894_,
		_w26897_,
		_w26898_
	);
	LUT2 #(
		.INIT('h4)
	) name16386 (
		_w26895_,
		_w26898_,
		_w26899_
	);
	LUT4 #(
		.INIT('hf1f0)
	) name16387 (
		\RxAbort_wb_reg/NET0131 ,
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\wishbone_RxEnableWindow_reg/NET0131 ,
		_w26900_
	);
	LUT2 #(
		.INIT('h6)
	) name16388 (
		\miim1_clkgen_Counter_reg[0]/NET0131 ,
		\miim1_clkgen_Counter_reg[1]/NET0131 ,
		_w26901_
	);
	LUT3 #(
		.INIT('h70)
	) name16389 (
		_w24411_,
		_w24420_,
		_w26901_,
		_w26902_
	);
	LUT2 #(
		.INIT('h9)
	) name16390 (
		\ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131 ,
		_w26903_
	);
	LUT2 #(
		.INIT('h1)
	) name16391 (
		\ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131 ,
		_w26904_
	);
	LUT3 #(
		.INIT('h4c)
	) name16392 (
		_w24415_,
		_w26903_,
		_w24416_,
		_w26905_
	);
	LUT3 #(
		.INIT('h31)
	) name16393 (
		_w24421_,
		_w26902_,
		_w26905_,
		_w26906_
	);
	LUT4 #(
		.INIT('h000b)
	) name16394 (
		\ethreg1_MODER_0_DataOut_reg[3]/NET0131 ,
		\rxethmac1_Broadcast_reg/NET0131 ,
		\rxethmac1_rxaddrcheck1_MulticastOK_reg/NET0131 ,
		\rxethmac1_rxaddrcheck1_UnicastOK_reg/NET0131 ,
		_w26907_
	);
	LUT2 #(
		.INIT('h8)
	) name16395 (
		\ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_AddressOK_reg/NET0131 ,
		_w26908_
	);
	LUT4 #(
		.INIT('h0080)
	) name16396 (
		_w11580_,
		_w11816_,
		_w26907_,
		_w26908_,
		_w26909_
	);
	LUT4 #(
		.INIT('hee2a)
	) name16397 (
		\rxethmac1_rxaddrcheck1_AddressMiss_reg/NET0131 ,
		_w10533_,
		_w11827_,
		_w26909_,
		_w26910_
	);
	LUT2 #(
		.INIT('h2)
	) name16398 (
		\wishbone_ram_di_reg[11]/NET0131 ,
		_w26389_,
		_w26911_
	);
	LUT4 #(
		.INIT('h002a)
	) name16399 (
		\wb_dat_i[11]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26912_
	);
	LUT2 #(
		.INIT('h8)
	) name16400 (
		\wishbone_TxEn_needed_reg/NET0131 ,
		\wishbone_TxStatus_reg[11]/NET0131 ,
		_w26913_
	);
	LUT4 #(
		.INIT('h8acf)
	) name16401 (
		_w26382_,
		_w26385_,
		_w26912_,
		_w26913_,
		_w26914_
	);
	LUT3 #(
		.INIT('h8f)
	) name16402 (
		_w26388_,
		_w26911_,
		_w26914_,
		_w26915_
	);
	LUT2 #(
		.INIT('h2)
	) name16403 (
		\wishbone_ram_di_reg[12]/NET0131 ,
		_w26389_,
		_w26916_
	);
	LUT4 #(
		.INIT('h002a)
	) name16404 (
		\wb_dat_i[12]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26917_
	);
	LUT2 #(
		.INIT('h8)
	) name16405 (
		\wishbone_TxEn_needed_reg/NET0131 ,
		\wishbone_TxStatus_reg[12]/NET0131 ,
		_w26918_
	);
	LUT4 #(
		.INIT('h8acf)
	) name16406 (
		_w26382_,
		_w26385_,
		_w26917_,
		_w26918_,
		_w26919_
	);
	LUT3 #(
		.INIT('h8f)
	) name16407 (
		_w26388_,
		_w26916_,
		_w26919_,
		_w26920_
	);
	LUT3 #(
		.INIT('h2a)
	) name16408 (
		\txethmac1_random1_RandomLatched_reg[8]/NET0131 ,
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w26921_
	);
	LUT3 #(
		.INIT('h01)
	) name16409 (
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		_w26922_
	);
	LUT4 #(
		.INIT('h8000)
	) name16410 (
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		\txethmac1_random1_x_reg[8]/NET0131 ,
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w26923_
	);
	LUT3 #(
		.INIT('hba)
	) name16411 (
		_w26921_,
		_w26922_,
		_w26923_,
		_w26924_
	);
	LUT4 #(
		.INIT('haa80)
	) name16412 (
		\wishbone_BDRead_reg/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w26925_
	);
	LUT2 #(
		.INIT('h2)
	) name16413 (
		\wishbone_BDRead_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		_w26926_
	);
	LUT3 #(
		.INIT('h23)
	) name16414 (
		_w26384_,
		_w26925_,
		_w26926_,
		_w26927_
	);
	LUT3 #(
		.INIT('h40)
	) name16415 (
		\wb_adr_i[11]_pad ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w26928_
	);
	LUT2 #(
		.INIT('h2)
	) name16416 (
		\wb_adr_i[10]_pad ,
		wb_we_i_pad,
		_w26929_
	);
	LUT3 #(
		.INIT('h40)
	) name16417 (
		_w18750_,
		_w26928_,
		_w26929_,
		_w26930_
	);
	LUT3 #(
		.INIT('hb3)
	) name16418 (
		_w26387_,
		_w26927_,
		_w26930_,
		_w26931_
	);
	LUT4 #(
		.INIT('hee0e)
	) name16419 (
		\wishbone_TxAbortPacketBlocked_reg/NET0131 ,
		\wishbone_TxAbortPacket_reg/NET0131 ,
		\wishbone_TxAbort_wb_q_reg/NET0131 ,
		\wishbone_TxAbort_wb_reg/NET0131 ,
		_w26932_
	);
	LUT4 #(
		.INIT('hee0e)
	) name16420 (
		\wishbone_TxDonePacketBlocked_reg/NET0131 ,
		\wishbone_TxDonePacket_reg/NET0131 ,
		\wishbone_TxDone_wb_q_reg/NET0131 ,
		\wishbone_TxDone_wb_reg/NET0131 ,
		_w26933_
	);
	LUT2 #(
		.INIT('h9)
	) name16421 (
		\txethmac1_random1_x_reg[2]/NET0131 ,
		\txethmac1_random1_x_reg[9]/NET0131 ,
		_w26934_
	);
	LUT2 #(
		.INIT('h2)
	) name16422 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w26935_
	);
	LUT4 #(
		.INIT('h7f00)
	) name16423 (
		_w11135_,
		_w11136_,
		_w11137_,
		_w26935_,
		_w26936_
	);
	LUT2 #(
		.INIT('h8)
	) name16424 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w26937_
	);
	LUT4 #(
		.INIT('h8000)
	) name16425 (
		_w11135_,
		_w11136_,
		_w11137_,
		_w26937_,
		_w26938_
	);
	LUT2 #(
		.INIT('h1)
	) name16426 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		\wishbone_LatchedRxLength_reg[11]/NET0131 ,
		_w26939_
	);
	LUT3 #(
		.INIT('h01)
	) name16427 (
		_w26936_,
		_w26938_,
		_w26939_,
		_w26940_
	);
	LUT3 #(
		.INIT('h07)
	) name16428 (
		\TPauseRq_reg/NET0131 ,
		\ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131 ,
		\maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131 ,
		_w26941_
	);
	LUT2 #(
		.INIT('h1)
	) name16429 (
		_w10602_,
		_w26941_,
		_w26942_
	);
	LUT3 #(
		.INIT('h4c)
	) name16430 (
		_w10744_,
		_w10745_,
		_w10755_,
		_w26943_
	);
	LUT4 #(
		.INIT('h1222)
	) name16431 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[4]/NET0131 ,
		wb_rst_i_pad,
		_w11279_,
		_w11280_,
		_w26944_
	);
	LUT3 #(
		.INIT('h15)
	) name16432 (
		\wishbone_TxBDAddress_reg[1]/NET0131 ,
		_w26321_,
		_w26324_,
		_w26945_
	);
	LUT2 #(
		.INIT('h4)
	) name16433 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		\wishbone_TxBDAddress_reg[1]/NET0131 ,
		_w26946_
	);
	LUT2 #(
		.INIT('h8)
	) name16434 (
		_w26321_,
		_w26946_,
		_w26947_
	);
	LUT3 #(
		.INIT('h01)
	) name16435 (
		_w26320_,
		_w26945_,
		_w26947_,
		_w26948_
	);
	LUT3 #(
		.INIT('h8c)
	) name16436 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		\wishbone_TxBDAddress_reg[2]/NET0131 ,
		_w26321_,
		_w26949_
	);
	LUT2 #(
		.INIT('h6)
	) name16437 (
		\wishbone_TxBDAddress_reg[1]/NET0131 ,
		\wishbone_TxBDAddress_reg[2]/NET0131 ,
		_w26950_
	);
	LUT3 #(
		.INIT('h80)
	) name16438 (
		_w26321_,
		_w26324_,
		_w26950_,
		_w26951_
	);
	LUT3 #(
		.INIT('h54)
	) name16439 (
		_w26320_,
		_w26949_,
		_w26951_,
		_w26952_
	);
	LUT3 #(
		.INIT('h8c)
	) name16440 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		\wishbone_TxBDAddress_reg[3]/NET0131 ,
		_w26321_,
		_w26953_
	);
	LUT3 #(
		.INIT('h78)
	) name16441 (
		\wishbone_TxBDAddress_reg[1]/NET0131 ,
		\wishbone_TxBDAddress_reg[2]/NET0131 ,
		\wishbone_TxBDAddress_reg[3]/NET0131 ,
		_w26954_
	);
	LUT3 #(
		.INIT('h80)
	) name16442 (
		_w26321_,
		_w26324_,
		_w26954_,
		_w26955_
	);
	LUT3 #(
		.INIT('h54)
	) name16443 (
		_w26320_,
		_w26953_,
		_w26955_,
		_w26956_
	);
	LUT3 #(
		.INIT('h8c)
	) name16444 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		\wishbone_TxBDAddress_reg[5]/NET0131 ,
		_w26321_,
		_w26957_
	);
	LUT4 #(
		.INIT('h4080)
	) name16445 (
		\wishbone_TxBDAddress_reg[5]/NET0131 ,
		_w26321_,
		_w26324_,
		_w26326_,
		_w26958_
	);
	LUT3 #(
		.INIT('h54)
	) name16446 (
		_w26320_,
		_w26957_,
		_w26958_,
		_w26959_
	);
	LUT4 #(
		.INIT('h4000)
	) name16447 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_Flop_reg/NET0131 ,
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		_w26960_
	);
	LUT4 #(
		.INIT('h000b)
	) name16448 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w26961_
	);
	LUT4 #(
		.INIT('h0004)
	) name16449 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_Flop_reg/NET0131 ,
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		_w26962_
	);
	LUT3 #(
		.INIT('h01)
	) name16450 (
		_w26960_,
		_w26961_,
		_w26962_,
		_w26963_
	);
	LUT4 #(
		.INIT('hb000)
	) name16451 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w26964_
	);
	LUT2 #(
		.INIT('h1)
	) name16452 (
		\wishbone_TxAbort_q_reg/NET0131 ,
		\wishbone_TxRetry_q_reg/NET0131 ,
		_w26965_
	);
	LUT2 #(
		.INIT('h4)
	) name16453 (
		_w26964_,
		_w26965_,
		_w26966_
	);
	LUT2 #(
		.INIT('h8)
	) name16454 (
		_w26963_,
		_w26966_,
		_w26967_
	);
	LUT3 #(
		.INIT('hb0)
	) name16455 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w26968_
	);
	LUT2 #(
		.INIT('h9)
	) name16456 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		_w26969_
	);
	LUT3 #(
		.INIT('h08)
	) name16457 (
		_w26965_,
		_w26968_,
		_w26969_,
		_w26970_
	);
	LUT2 #(
		.INIT('h8)
	) name16458 (
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		_w26960_,
		_w26971_
	);
	LUT4 #(
		.INIT('h0060)
	) name16459 (
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		_w26960_,
		_w26965_,
		_w26968_,
		_w26972_
	);
	LUT2 #(
		.INIT('he)
	) name16460 (
		_w26970_,
		_w26972_,
		_w26973_
	);
	LUT4 #(
		.INIT('h008c)
	) name16461 (
		\wishbone_TxEn_needed_reg/NET0131 ,
		\wishbone_WbEn_reg/NET0131 ,
		_w26381_,
		_w26389_,
		_w26974_
	);
	LUT3 #(
		.INIT('hdc)
	) name16462 (
		_w26383_,
		_w26387_,
		_w26974_,
		_w26975_
	);
	LUT3 #(
		.INIT('h10)
	) name16463 (
		\miim1_BitCounter_reg[5]/NET0131 ,
		\miim1_BitCounter_reg[6]/NET0131 ,
		\miim1_InProgress_reg/NET0131 ,
		_w26976_
	);
	LUT3 #(
		.INIT('hfe)
	) name16464 (
		_w24567_,
		_w26351_,
		_w26976_,
		_w26977_
	);
	LUT3 #(
		.INIT('h80)
	) name16465 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		_w26978_
	);
	LUT4 #(
		.INIT('h007f)
	) name16466 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		_w26979_
	);
	LUT4 #(
		.INIT('h0001)
	) name16467 (
		_w26302_,
		_w26303_,
		_w26304_,
		_w26979_,
		_w26980_
	);
	LUT4 #(
		.INIT('h4544)
	) name16468 (
		wb_ack_o_pad,
		\wishbone_WB_ACK_O_reg/P0001 ,
		_w18750_,
		_w18751_,
		_w26981_
	);
	LUT2 #(
		.INIT('h8)
	) name16469 (
		_w19640_,
		_w26136_,
		_w26982_
	);
	LUT4 #(
		.INIT('h060c)
	) name16470 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_SlotTimer_reg[2]/NET0131 ,
		wb_rst_i_pad,
		_w11279_,
		_w26983_
	);
	LUT2 #(
		.INIT('h8)
	) name16471 (
		_w18794_,
		_w26168_,
		_w26984_
	);
	LUT4 #(
		.INIT('h0020)
	) name16472 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w26985_
	);
	LUT2 #(
		.INIT('h8)
	) name16473 (
		_w26361_,
		_w26985_,
		_w26986_
	);
	LUT4 #(
		.INIT('h0008)
	) name16474 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26987_
	);
	LUT4 #(
		.INIT('h0200)
	) name16475 (
		\ethreg1_TXCTRL_1_DataOut_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26988_
	);
	LUT4 #(
		.INIT('h153f)
	) name16476 (
		_w26365_,
		_w26370_,
		_w26987_,
		_w26988_,
		_w26989_
	);
	LUT2 #(
		.INIT('h4)
	) name16477 (
		_w26986_,
		_w26989_,
		_w26990_
	);
	LUT4 #(
		.INIT('h0008)
	) name16478 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26991_
	);
	LUT3 #(
		.INIT('h08)
	) name16479 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26992_
	);
	LUT2 #(
		.INIT('h1)
	) name16480 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w26993_
	);
	LUT4 #(
		.INIT('h0777)
	) name16481 (
		_w26359_,
		_w26991_,
		_w26992_,
		_w26993_,
		_w26994_
	);
	LUT4 #(
		.INIT('h0020)
	) name16482 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26995_
	);
	LUT4 #(
		.INIT('h0200)
	) name16483 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w26996_
	);
	LUT4 #(
		.INIT('h153f)
	) name16484 (
		_w26361_,
		_w26370_,
		_w26995_,
		_w26996_,
		_w26997_
	);
	LUT4 #(
		.INIT('h0200)
	) name16485 (
		\ethreg1_TXCTRL_0_DataOut_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26998_
	);
	LUT4 #(
		.INIT('h0020)
	) name16486 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w26999_
	);
	LUT4 #(
		.INIT('h135f)
	) name16487 (
		_w25925_,
		_w26365_,
		_w26998_,
		_w26999_,
		_w27000_
	);
	LUT3 #(
		.INIT('h80)
	) name16488 (
		_w26994_,
		_w26997_,
		_w27000_,
		_w27001_
	);
	LUT2 #(
		.INIT('h7)
	) name16489 (
		_w26990_,
		_w27001_,
		_w27002_
	);
	LUT4 #(
		.INIT('h2322)
	) name16490 (
		\macstatus1_DribbleNibble_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w10575_,
		_w11386_,
		_w27003_
	);
	LUT2 #(
		.INIT('h4)
	) name16491 (
		\rxethmac1_crcrx_Crc_reg[28]/NET0131 ,
		_w10536_,
		_w27004_
	);
	LUT3 #(
		.INIT('h02)
	) name16492 (
		\rxethmac1_CrcHash_reg[2]/P0001 ,
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		wb_rst_i_pad,
		_w27005_
	);
	LUT4 #(
		.INIT('h7270)
	) name16493 (
		_w10533_,
		_w27004_,
		_w27005_,
		_w10540_,
		_w27006_
	);
	LUT2 #(
		.INIT('h4)
	) name16494 (
		\rxethmac1_crcrx_Crc_reg[29]/NET0131 ,
		_w10536_,
		_w27007_
	);
	LUT3 #(
		.INIT('h02)
	) name16495 (
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		wb_rst_i_pad,
		_w27008_
	);
	LUT4 #(
		.INIT('h5f08)
	) name16496 (
		_w10533_,
		_w10540_,
		_w27007_,
		_w27008_,
		_w27009_
	);
	LUT2 #(
		.INIT('h4)
	) name16497 (
		\rxethmac1_crcrx_Crc_reg[30]/NET0131 ,
		_w10536_,
		_w27010_
	);
	LUT3 #(
		.INIT('h02)
	) name16498 (
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		wb_rst_i_pad,
		_w27011_
	);
	LUT4 #(
		.INIT('h5f08)
	) name16499 (
		_w10533_,
		_w10540_,
		_w27010_,
		_w27011_,
		_w27012_
	);
	LUT2 #(
		.INIT('h4)
	) name16500 (
		\rxethmac1_crcrx_Crc_reg[31]/NET0131 ,
		_w10536_,
		_w27013_
	);
	LUT3 #(
		.INIT('h02)
	) name16501 (
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		wb_rst_i_pad,
		_w27014_
	);
	LUT4 #(
		.INIT('h5f08)
	) name16502 (
		_w10533_,
		_w10540_,
		_w27013_,
		_w27014_,
		_w27015_
	);
	LUT4 #(
		.INIT('h1555)
	) name16503 (
		\wishbone_ReadTxDataFromMemory_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w27016_
	);
	LUT2 #(
		.INIT('h2)
	) name16504 (
		_w25940_,
		_w27016_,
		_w27017_
	);
	LUT3 #(
		.INIT('h70)
	) name16505 (
		_w12312_,
		_w26342_,
		_w27017_,
		_w27018_
	);
	LUT3 #(
		.INIT('hf8)
	) name16506 (
		\wishbone_RxEn_reg/NET0131 ,
		_w26388_,
		_w26389_,
		_w27019_
	);
	LUT3 #(
		.INIT('h6a)
	) name16507 (
		mdc_pad_o_pad,
		_w24411_,
		_w24420_,
		_w27020_
	);
	LUT2 #(
		.INIT('h8)
	) name16508 (
		\rxethmac1_LatchedByte_reg[1]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w27021_
	);
	LUT3 #(
		.INIT('h70)
	) name16509 (
		_w10519_,
		_w24852_,
		_w27021_,
		_w27022_
	);
	LUT2 #(
		.INIT('h8)
	) name16510 (
		\rxethmac1_DelayData_reg/NET0131 ,
		\rxethmac1_RxData_d_reg[1]/NET0131 ,
		_w27023_
	);
	LUT4 #(
		.INIT('hd500)
	) name16511 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10519_,
		_w24852_,
		_w27023_,
		_w27024_
	);
	LUT2 #(
		.INIT('he)
	) name16512 (
		_w27022_,
		_w27024_,
		_w27025_
	);
	LUT2 #(
		.INIT('h8)
	) name16513 (
		\rxethmac1_LatchedByte_reg[2]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w27026_
	);
	LUT3 #(
		.INIT('h70)
	) name16514 (
		_w10519_,
		_w24852_,
		_w27026_,
		_w27027_
	);
	LUT2 #(
		.INIT('h8)
	) name16515 (
		\rxethmac1_DelayData_reg/NET0131 ,
		\rxethmac1_RxData_d_reg[2]/NET0131 ,
		_w27028_
	);
	LUT4 #(
		.INIT('hd500)
	) name16516 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10519_,
		_w24852_,
		_w27028_,
		_w27029_
	);
	LUT2 #(
		.INIT('he)
	) name16517 (
		_w27027_,
		_w27029_,
		_w27030_
	);
	LUT2 #(
		.INIT('h8)
	) name16518 (
		\rxethmac1_LatchedByte_reg[3]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w27031_
	);
	LUT3 #(
		.INIT('h70)
	) name16519 (
		_w10519_,
		_w24852_,
		_w27031_,
		_w27032_
	);
	LUT2 #(
		.INIT('h8)
	) name16520 (
		\rxethmac1_DelayData_reg/NET0131 ,
		\rxethmac1_RxData_d_reg[3]/NET0131 ,
		_w27033_
	);
	LUT4 #(
		.INIT('hd500)
	) name16521 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10519_,
		_w24852_,
		_w27033_,
		_w27034_
	);
	LUT2 #(
		.INIT('he)
	) name16522 (
		_w27032_,
		_w27034_,
		_w27035_
	);
	LUT2 #(
		.INIT('h8)
	) name16523 (
		\rxethmac1_LatchedByte_reg[5]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w27036_
	);
	LUT3 #(
		.INIT('h70)
	) name16524 (
		_w10519_,
		_w24852_,
		_w27036_,
		_w27037_
	);
	LUT2 #(
		.INIT('h8)
	) name16525 (
		\rxethmac1_DelayData_reg/NET0131 ,
		\rxethmac1_RxData_d_reg[5]/NET0131 ,
		_w27038_
	);
	LUT4 #(
		.INIT('hd500)
	) name16526 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10519_,
		_w24852_,
		_w27038_,
		_w27039_
	);
	LUT2 #(
		.INIT('he)
	) name16527 (
		_w27037_,
		_w27039_,
		_w27040_
	);
	LUT2 #(
		.INIT('h8)
	) name16528 (
		\rxethmac1_LatchedByte_reg[6]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w27041_
	);
	LUT3 #(
		.INIT('h70)
	) name16529 (
		_w10519_,
		_w24852_,
		_w27041_,
		_w27042_
	);
	LUT2 #(
		.INIT('h8)
	) name16530 (
		\rxethmac1_DelayData_reg/NET0131 ,
		\rxethmac1_RxData_d_reg[6]/NET0131 ,
		_w27043_
	);
	LUT4 #(
		.INIT('hd500)
	) name16531 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10519_,
		_w24852_,
		_w27043_,
		_w27044_
	);
	LUT2 #(
		.INIT('he)
	) name16532 (
		_w27042_,
		_w27044_,
		_w27045_
	);
	LUT2 #(
		.INIT('h8)
	) name16533 (
		\rxethmac1_LatchedByte_reg[7]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w27046_
	);
	LUT3 #(
		.INIT('h70)
	) name16534 (
		_w10519_,
		_w24852_,
		_w27046_,
		_w27047_
	);
	LUT2 #(
		.INIT('h8)
	) name16535 (
		\rxethmac1_DelayData_reg/NET0131 ,
		\rxethmac1_RxData_d_reg[7]/NET0131 ,
		_w27048_
	);
	LUT4 #(
		.INIT('hd500)
	) name16536 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10519_,
		_w24852_,
		_w27048_,
		_w27049_
	);
	LUT2 #(
		.INIT('he)
	) name16537 (
		_w27047_,
		_w27049_,
		_w27050_
	);
	LUT2 #(
		.INIT('h2)
	) name16538 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w27051_
	);
	LUT3 #(
		.INIT('he6)
	) name16539 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w27052_
	);
	LUT4 #(
		.INIT('h1300)
	) name16540 (
		_w10543_,
		_w26304_,
		_w27051_,
		_w27052_,
		_w27053_
	);
	LUT2 #(
		.INIT('h2)
	) name16541 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		_w27054_
	);
	LUT2 #(
		.INIT('h8)
	) name16542 (
		_w26136_,
		_w27054_,
		_w27055_
	);
	LUT3 #(
		.INIT('h04)
	) name16543 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[5]_pad ,
		_w27056_
	);
	LUT2 #(
		.INIT('h8)
	) name16544 (
		_w18753_,
		_w27056_,
		_w27057_
	);
	LUT3 #(
		.INIT('h10)
	) name16545 (
		\wb_adr_i[10]_pad ,
		\wb_adr_i[4]_pad ,
		wb_we_i_pad,
		_w27058_
	);
	LUT3 #(
		.INIT('h40)
	) name16546 (
		_w18750_,
		_w24750_,
		_w27058_,
		_w27059_
	);
	LUT2 #(
		.INIT('h8)
	) name16547 (
		_w27057_,
		_w27059_,
		_w27060_
	);
	LUT2 #(
		.INIT('h2)
	) name16548 (
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxEndFrm_wb_reg/NET0131 ,
		_w27061_
	);
	LUT2 #(
		.INIT('h8)
	) name16549 (
		_w26960_,
		_w27061_,
		_w27062_
	);
	LUT3 #(
		.INIT('hc8)
	) name16550 (
		\txethmac1_TxRetry_reg/NET0131 ,
		\wishbone_Flop_reg/NET0131 ,
		\wishbone_TxEndFrm_reg/NET0131 ,
		_w27063_
	);
	LUT4 #(
		.INIT('h0054)
	) name16551 (
		\maccontrol1_transmitcontrol1_BlockTxDone_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxAbort_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w27064_
	);
	LUT2 #(
		.INIT('h4)
	) name16552 (
		\maccontrol1_MuxedAbort_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w27065_
	);
	LUT3 #(
		.INIT('hb0)
	) name16553 (
		\maccontrol1_MuxedAbort_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\wishbone_Flop_reg/NET0131 ,
		_w27066_
	);
	LUT3 #(
		.INIT('h15)
	) name16554 (
		_w27063_,
		_w27064_,
		_w27066_,
		_w27067_
	);
	LUT3 #(
		.INIT('h15)
	) name16555 (
		\wishbone_LastWord_reg/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		_w26960_,
		_w27068_
	);
	LUT3 #(
		.INIT('h04)
	) name16556 (
		_w27062_,
		_w27067_,
		_w27068_,
		_w27069_
	);
	LUT4 #(
		.INIT('haa80)
	) name16557 (
		\wishbone_BDWrite_reg[0]/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w27070_
	);
	LUT2 #(
		.INIT('h2)
	) name16558 (
		\wishbone_BDWrite_reg[0]/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		_w27071_
	);
	LUT3 #(
		.INIT('h23)
	) name16559 (
		_w26384_,
		_w27070_,
		_w27071_,
		_w27072_
	);
	LUT2 #(
		.INIT('h8)
	) name16560 (
		\wb_adr_i[10]_pad ,
		wb_we_i_pad,
		_w27073_
	);
	LUT3 #(
		.INIT('h40)
	) name16561 (
		_w26385_,
		_w26386_,
		_w27073_,
		_w27074_
	);
	LUT3 #(
		.INIT('hb3)
	) name16562 (
		_w24751_,
		_w27072_,
		_w27074_,
		_w27075_
	);
	LUT4 #(
		.INIT('haa80)
	) name16563 (
		\wishbone_BDWrite_reg[1]/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w27076_
	);
	LUT2 #(
		.INIT('h2)
	) name16564 (
		\wishbone_BDWrite_reg[1]/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		_w27077_
	);
	LUT3 #(
		.INIT('h23)
	) name16565 (
		_w26384_,
		_w27076_,
		_w27077_,
		_w27078_
	);
	LUT4 #(
		.INIT('h4000)
	) name16566 (
		\wb_adr_i[11]_pad ,
		wb_cyc_i_pad,
		\wb_sel_i[1]_pad ,
		wb_stb_i_pad,
		_w27079_
	);
	LUT2 #(
		.INIT('h4)
	) name16567 (
		_w18750_,
		_w27079_,
		_w27080_
	);
	LUT3 #(
		.INIT('hb3)
	) name16568 (
		_w27074_,
		_w27078_,
		_w27080_,
		_w27081_
	);
	LUT4 #(
		.INIT('haa80)
	) name16569 (
		\wishbone_BDWrite_reg[2]/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w27082_
	);
	LUT2 #(
		.INIT('h2)
	) name16570 (
		\wishbone_BDWrite_reg[2]/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		_w27083_
	);
	LUT3 #(
		.INIT('h23)
	) name16571 (
		_w26384_,
		_w27082_,
		_w27083_,
		_w27084_
	);
	LUT3 #(
		.INIT('h8f)
	) name16572 (
		_w26893_,
		_w27074_,
		_w27084_,
		_w27085_
	);
	LUT2 #(
		.INIT('h4)
	) name16573 (
		\wishbone_LastWord_reg/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		_w27086_
	);
	LUT2 #(
		.INIT('h8)
	) name16574 (
		_w26960_,
		_w27086_,
		_w27087_
	);
	LUT3 #(
		.INIT('h10)
	) name16575 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w27088_
	);
	LUT3 #(
		.INIT('hd0)
	) name16576 (
		\wishbone_ReadTxDataFromFifo_syncb2_reg/NET0131 ,
		\wishbone_ReadTxDataFromFifo_syncb3_reg/NET0131 ,
		\wishbone_ReadTxDataFromFifo_tck_reg/NET0131 ,
		_w27089_
	);
	LUT4 #(
		.INIT('h0013)
	) name16577 (
		_w11658_,
		_w11666_,
		_w27088_,
		_w27089_,
		_w27090_
	);
	LUT2 #(
		.INIT('hb)
	) name16578 (
		_w27087_,
		_w27090_,
		_w27091_
	);
	LUT3 #(
		.INIT('h15)
	) name16579 (
		\ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131 ,
		_w24415_,
		_w26904_,
		_w27092_
	);
	LUT3 #(
		.INIT('hd1)
	) name16580 (
		\miim1_clkgen_Counter_reg[0]/NET0131 ,
		_w24421_,
		_w27092_,
		_w27093_
	);
	LUT3 #(
		.INIT('h2a)
	) name16581 (
		\wishbone_TxAbortPacket_NotCleared_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w27094_
	);
	LUT3 #(
		.INIT('h0e)
	) name16582 (
		m_wb_ack_i_pad,
		m_wb_err_i_pad,
		\wishbone_tx_burst_en_reg/NET0131 ,
		_w27095_
	);
	LUT4 #(
		.INIT('hf010)
	) name16583 (
		m_wb_ack_i_pad,
		m_wb_err_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_tx_burst_en_reg/NET0131 ,
		_w27096_
	);
	LUT2 #(
		.INIT('h4)
	) name16584 (
		\wishbone_TxAbortPacketBlocked_reg/NET0131 ,
		\wishbone_TxAbort_wb_reg/NET0131 ,
		_w27097_
	);
	LUT3 #(
		.INIT('h10)
	) name16585 (
		\wishbone_TxAbortPacketBlocked_reg/NET0131 ,
		\wishbone_TxAbortPacket_NotCleared_reg/NET0131 ,
		\wishbone_TxAbort_wb_reg/NET0131 ,
		_w27098_
	);
	LUT3 #(
		.INIT('hba)
	) name16586 (
		_w27094_,
		_w27096_,
		_w27098_,
		_w27099_
	);
	LUT3 #(
		.INIT('h2a)
	) name16587 (
		\wishbone_TxDonePacket_NotCleared_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w27100_
	);
	LUT2 #(
		.INIT('h4)
	) name16588 (
		\wishbone_TxDonePacketBlocked_reg/NET0131 ,
		\wishbone_TxDone_wb_reg/NET0131 ,
		_w27101_
	);
	LUT3 #(
		.INIT('h10)
	) name16589 (
		\wishbone_TxDonePacketBlocked_reg/NET0131 ,
		\wishbone_TxDonePacket_NotCleared_reg/NET0131 ,
		\wishbone_TxDone_wb_reg/NET0131 ,
		_w27102_
	);
	LUT3 #(
		.INIT('hdc)
	) name16590 (
		_w27096_,
		_w27100_,
		_w27102_,
		_w27103_
	);
	LUT4 #(
		.INIT('h0800)
	) name16591 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		_w27104_
	);
	LUT3 #(
		.INIT('h07)
	) name16592 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		_w27105_
	);
	LUT3 #(
		.INIT('h01)
	) name16593 (
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[4]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		_w27106_
	);
	LUT3 #(
		.INIT('h13)
	) name16594 (
		_w11866_,
		_w27105_,
		_w27106_,
		_w27107_
	);
	LUT3 #(
		.INIT('h80)
	) name16595 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		_w27108_
	);
	LUT4 #(
		.INIT('h080f)
	) name16596 (
		_w11866_,
		_w11867_,
		_w24970_,
		_w27108_,
		_w27109_
	);
	LUT3 #(
		.INIT('hea)
	) name16597 (
		_w27104_,
		_w27107_,
		_w27109_,
		_w27110_
	);
	LUT3 #(
		.INIT('ha8)
	) name16598 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[1]/NET0131 ,
		_w25875_,
		_w25876_,
		_w27111_
	);
	LUT4 #(
		.INIT('h0102)
	) name16599 (
		\wishbone_RxBDAddress_reg[2]/NET0131 ,
		_w25875_,
		_w25876_,
		_w26186_,
		_w27112_
	);
	LUT2 #(
		.INIT('he)
	) name16600 (
		_w27111_,
		_w27112_,
		_w27113_
	);
	LUT4 #(
		.INIT('h002a)
	) name16601 (
		\wb_dat_i[10]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w27114_
	);
	LUT2 #(
		.INIT('h4)
	) name16602 (
		_w26385_,
		_w27114_,
		_w27115_
	);
	LUT2 #(
		.INIT('h2)
	) name16603 (
		\wishbone_ram_di_reg[10]/NET0131 ,
		_w26389_,
		_w27116_
	);
	LUT3 #(
		.INIT('hec)
	) name16604 (
		_w26388_,
		_w27115_,
		_w27116_,
		_w27117_
	);
	LUT4 #(
		.INIT('h002a)
	) name16605 (
		\wb_dat_i[15]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w27118_
	);
	LUT2 #(
		.INIT('h4)
	) name16606 (
		_w26385_,
		_w27118_,
		_w27119_
	);
	LUT2 #(
		.INIT('h2)
	) name16607 (
		\wishbone_ram_di_reg[15]/NET0131 ,
		_w26389_,
		_w27120_
	);
	LUT3 #(
		.INIT('hec)
	) name16608 (
		_w26388_,
		_w27119_,
		_w27120_,
		_w27121_
	);
	LUT4 #(
		.INIT('h002a)
	) name16609 (
		\wb_dat_i[9]_pad ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w27122_
	);
	LUT2 #(
		.INIT('h4)
	) name16610 (
		_w26385_,
		_w27122_,
		_w27123_
	);
	LUT2 #(
		.INIT('h2)
	) name16611 (
		\wishbone_ram_di_reg[9]/NET0131 ,
		_w26389_,
		_w27124_
	);
	LUT3 #(
		.INIT('hec)
	) name16612 (
		_w26388_,
		_w27123_,
		_w27124_,
		_w27125_
	);
	LUT4 #(
		.INIT('hd777)
	) name16613 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w11135_,
		_w11136_,
		_w27126_
	);
	LUT2 #(
		.INIT('h4)
	) name16614 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		\wishbone_LatchedRxLength_reg[8]/NET0131 ,
		_w27127_
	);
	LUT2 #(
		.INIT('hd)
	) name16615 (
		_w27126_,
		_w27127_,
		_w27128_
	);
	LUT4 #(
		.INIT('h7ddd)
	) name16616 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		_w11135_,
		_w11168_,
		_w27129_
	);
	LUT2 #(
		.INIT('h1)
	) name16617 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		\wishbone_LatchedRxLength_reg[7]/NET0131 ,
		_w27130_
	);
	LUT2 #(
		.INIT('h2)
	) name16618 (
		_w27129_,
		_w27130_,
		_w27131_
	);
	LUT3 #(
		.INIT('h6c)
	) name16619 (
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		_w11140_,
		_w27132_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name16620 (
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w11135_,
		_w11136_,
		_w27133_
	);
	LUT2 #(
		.INIT('h6)
	) name16621 (
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w11135_,
		_w27134_
	);
	LUT4 #(
		.INIT('h00d0)
	) name16622 (
		\txethmac1_TxRetry_reg/NET0131 ,
		\wishbone_TxRetry_q_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		\wishbone_TxUsedData_q_reg/NET0131 ,
		_w27135_
	);
	LUT2 #(
		.INIT('he)
	) name16623 (
		\wishbone_TxStartFrm_sync2_reg/NET0131 ,
		_w27135_,
		_w27136_
	);
	LUT4 #(
		.INIT('h4055)
	) name16624 (
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		_w11866_,
		_w11867_,
		_w27108_,
		_w27137_
	);
	LUT4 #(
		.INIT('h080f)
	) name16625 (
		_w11866_,
		_w11867_,
		_w24970_,
		_w26835_,
		_w27138_
	);
	LUT2 #(
		.INIT('h4)
	) name16626 (
		_w27137_,
		_w27138_,
		_w27139_
	);
	LUT4 #(
		.INIT('h4000)
	) name16627 (
		_w18750_,
		_w18753_,
		_w24750_,
		_w24752_,
		_w27140_
	);
	LUT4 #(
		.INIT('h2000)
	) name16628 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w27141_
	);
	LUT2 #(
		.INIT('h8)
	) name16629 (
		_w27140_,
		_w27141_,
		_w27142_
	);
	LUT4 #(
		.INIT('h4000)
	) name16630 (
		_w18750_,
		_w18753_,
		_w24752_,
		_w27079_,
		_w27143_
	);
	LUT2 #(
		.INIT('h8)
	) name16631 (
		_w27141_,
		_w27143_,
		_w27144_
	);
	LUT4 #(
		.INIT('h0200)
	) name16632 (
		\wishbone_WriteRxDataToFifoSync2_reg/NET0131 ,
		\wishbone_WriteRxDataToFifoSync3_reg/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[4]/NET0131 ,
		_w27145_
	);
	LUT4 #(
		.INIT('h0e0a)
	) name16633 (
		\wishbone_RxOverrun_reg/NET0131 ,
		_w11866_,
		_w25879_,
		_w27145_,
		_w27146_
	);
	LUT4 #(
		.INIT('h0002)
	) name16634 (
		\wishbone_ReadTxDataFromFifo_sync2_reg/NET0131 ,
		\wishbone_ReadTxDataFromFifo_sync3_reg/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w27147_
	);
	LUT4 #(
		.INIT('h0e0a)
	) name16635 (
		\wishbone_TxUnderRun_wb_reg/NET0131 ,
		_w25795_,
		_w25939_,
		_w27147_,
		_w27148_
	);
	LUT2 #(
		.INIT('h8)
	) name16636 (
		_w19642_,
		_w24753_,
		_w27149_
	);
	LUT2 #(
		.INIT('h8)
	) name16637 (
		_w19642_,
		_w26894_,
		_w27150_
	);
	LUT4 #(
		.INIT('h4000)
	) name16638 (
		\ethreg1_MODER_0_DataOut_reg[5]/NET0131 ,
		_w11580_,
		_w11816_,
		_w26907_,
		_w27151_
	);
	LUT2 #(
		.INIT('h8)
	) name16639 (
		_w10533_,
		_w27151_,
		_w27152_
	);
	LUT3 #(
		.INIT('h80)
	) name16640 (
		_w18757_,
		_w18762_,
		_w18765_,
		_w27153_
	);
	LUT2 #(
		.INIT('h8)
	) name16641 (
		_w24753_,
		_w27153_,
		_w27154_
	);
	LUT3 #(
		.INIT('h78)
	) name16642 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		_w27155_
	);
	LUT3 #(
		.INIT('h10)
	) name16643 (
		_w26303_,
		_w26304_,
		_w27155_,
		_w27156_
	);
	LUT3 #(
		.INIT('h40)
	) name16644 (
		_w18750_,
		_w24752_,
		_w27079_,
		_w27157_
	);
	LUT2 #(
		.INIT('h8)
	) name16645 (
		_w27153_,
		_w27157_,
		_w27158_
	);
	LUT2 #(
		.INIT('h2)
	) name16646 (
		\ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_Divider2_reg/NET0131 ,
		_w27159_
	);
	LUT3 #(
		.INIT('h70)
	) name16647 (
		_w11273_,
		_w11277_,
		_w27159_,
		_w27160_
	);
	LUT3 #(
		.INIT('hb0)
	) name16648 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		_w27161_
	);
	LUT4 #(
		.INIT('h8f00)
	) name16649 (
		_w11866_,
		_w11867_,
		_w26835_,
		_w27161_,
		_w27162_
	);
	LUT3 #(
		.INIT('h0b)
	) name16650 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		_w27163_
	);
	LUT4 #(
		.INIT('h7000)
	) name16651 (
		_w11866_,
		_w11867_,
		_w26835_,
		_w27163_,
		_w27164_
	);
	LUT2 #(
		.INIT('he)
	) name16652 (
		_w27162_,
		_w27164_,
		_w27165_
	);
	LUT4 #(
		.INIT('h0010)
	) name16653 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w27166_
	);
	LUT2 #(
		.INIT('h8)
	) name16654 (
		_w27140_,
		_w27166_,
		_w27167_
	);
	LUT4 #(
		.INIT('h1333)
	) name16655 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[4]/NET0131 ,
		\maccontrol1_receivecontrol1_SlotTimer_reg[5]/NET0131 ,
		_w11279_,
		_w11280_,
		_w27168_
	);
	LUT4 #(
		.INIT('h1555)
	) name16656 (
		wb_rst_i_pad,
		_w11279_,
		_w11280_,
		_w11281_,
		_w27169_
	);
	LUT2 #(
		.INIT('h4)
	) name16657 (
		_w27168_,
		_w27169_,
		_w27170_
	);
	LUT3 #(
		.INIT('h07)
	) name16658 (
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131 ,
		_w27171_
	);
	LUT3 #(
		.INIT('hec)
	) name16659 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w27172_
	);
	LUT3 #(
		.INIT('h20)
	) name16660 (
		_w25933_,
		_w27171_,
		_w27172_,
		_w27173_
	);
	LUT2 #(
		.INIT('hd)
	) name16661 (
		_w10847_,
		_w10938_,
		_w27174_
	);
	LUT3 #(
		.INIT('h2a)
	) name16662 (
		\txethmac1_random1_RandomLatched_reg[5]/NET0131 ,
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w27175_
	);
	LUT3 #(
		.INIT('h07)
	) name16663 (
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w27176_
	);
	LUT3 #(
		.INIT('h80)
	) name16664 (
		\txethmac1_random1_x_reg[5]/NET0131 ,
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w27177_
	);
	LUT3 #(
		.INIT('hba)
	) name16665 (
		_w27175_,
		_w27176_,
		_w27177_,
		_w27178_
	);
	LUT3 #(
		.INIT('h08)
	) name16666 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[5]_pad ,
		_w27179_
	);
	LUT2 #(
		.INIT('h8)
	) name16667 (
		_w18753_,
		_w27179_,
		_w27180_
	);
	LUT2 #(
		.INIT('h8)
	) name16668 (
		_w27059_,
		_w27180_,
		_w27181_
	);
	LUT3 #(
		.INIT('hfd)
	) name16669 (
		_w11007_,
		_w11090_,
		_w11092_,
		_w27182_
	);
	LUT4 #(
		.INIT('haa80)
	) name16670 (
		\wishbone_BDWrite_reg[3]/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w27183_
	);
	LUT2 #(
		.INIT('h2)
	) name16671 (
		\wishbone_BDWrite_reg[3]/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		_w27184_
	);
	LUT3 #(
		.INIT('h23)
	) name16672 (
		_w26384_,
		_w27183_,
		_w27184_,
		_w27185_
	);
	LUT4 #(
		.INIT('h4000)
	) name16673 (
		\wb_adr_i[11]_pad ,
		wb_cyc_i_pad,
		\wb_sel_i[3]_pad ,
		wb_stb_i_pad,
		_w27186_
	);
	LUT2 #(
		.INIT('h4)
	) name16674 (
		_w18750_,
		_w27186_,
		_w27187_
	);
	LUT3 #(
		.INIT('hb3)
	) name16675 (
		_w27074_,
		_w27185_,
		_w27187_,
		_w27188_
	);
	LUT2 #(
		.INIT('h9)
	) name16676 (
		\wishbone_BlockingTxBDRead_reg/NET0131 ,
		\wishbone_TxBDReady_reg/NET0131 ,
		_w27189_
	);
	LUT2 #(
		.INIT('h1)
	) name16677 (
		\wishbone_BlockingTxBDRead_reg/NET0131 ,
		\wishbone_TxRetryPacket_NotCleared_reg/NET0131 ,
		_w27190_
	);
	LUT4 #(
		.INIT('h40f0)
	) name16678 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		_w26321_,
		_w27189_,
		_w27190_,
		_w27191_
	);
	LUT2 #(
		.INIT('h4)
	) name16679 (
		\wishbone_TxStartFrm_syncb2_reg/NET0131 ,
		\wishbone_TxStartFrm_wb_reg/NET0131 ,
		_w27192_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name16680 (
		\wishbone_StartOccured_reg/NET0131 ,
		\wishbone_TxBDReady_reg/NET0131 ,
		\wishbone_TxStartFrm_syncb2_reg/NET0131 ,
		\wishbone_TxStartFrm_wb_reg/NET0131 ,
		_w27193_
	);
	LUT3 #(
		.INIT('h07)
	) name16681 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w25802_,
		_w27192_,
		_w27194_
	);
	LUT4 #(
		.INIT('h080f)
	) name16682 (
		_w12312_,
		_w26342_,
		_w27193_,
		_w27194_,
		_w27195_
	);
	LUT4 #(
		.INIT('h1000)
	) name16683 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w27196_
	);
	LUT2 #(
		.INIT('h8)
	) name16684 (
		_w27140_,
		_w27196_,
		_w27197_
	);
	LUT2 #(
		.INIT('h8)
	) name16685 (
		_w27143_,
		_w27196_,
		_w27198_
	);
	LUT4 #(
		.INIT('h0400)
	) name16686 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w27199_
	);
	LUT2 #(
		.INIT('h8)
	) name16687 (
		_w27140_,
		_w27199_,
		_w27200_
	);
	LUT2 #(
		.INIT('h8)
	) name16688 (
		_w27143_,
		_w27199_,
		_w27201_
	);
	LUT4 #(
		.INIT('h0200)
	) name16689 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w27202_
	);
	LUT2 #(
		.INIT('h8)
	) name16690 (
		_w26361_,
		_w27202_,
		_w27203_
	);
	LUT4 #(
		.INIT('h0200)
	) name16691 (
		\ethreg1_TXCTRL_1_DataOut_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w27204_
	);
	LUT4 #(
		.INIT('h0008)
	) name16692 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w27205_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16693 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w26358_,
		_w27204_,
		_w27205_,
		_w27206_
	);
	LUT2 #(
		.INIT('h4)
	) name16694 (
		_w27203_,
		_w27206_,
		_w27207_
	);
	LUT4 #(
		.INIT('h0008)
	) name16695 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w27208_
	);
	LUT4 #(
		.INIT('h0777)
	) name16696 (
		_w26359_,
		_w26366_,
		_w26370_,
		_w27208_,
		_w27209_
	);
	LUT4 #(
		.INIT('h0020)
	) name16697 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w27210_
	);
	LUT4 #(
		.INIT('h0200)
	) name16698 (
		\ethreg1_TXCTRL_0_DataOut_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w27211_
	);
	LUT4 #(
		.INIT('h153f)
	) name16699 (
		_w25925_,
		_w26365_,
		_w27210_,
		_w27211_,
		_w27212_
	);
	LUT4 #(
		.INIT('h0020)
	) name16700 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w27213_
	);
	LUT4 #(
		.INIT('h0020)
	) name16701 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w27214_
	);
	LUT4 #(
		.INIT('h135f)
	) name16702 (
		_w26361_,
		_w26370_,
		_w27213_,
		_w27214_,
		_w27215_
	);
	LUT3 #(
		.INIT('h80)
	) name16703 (
		_w27209_,
		_w27212_,
		_w27215_,
		_w27216_
	);
	LUT2 #(
		.INIT('h7)
	) name16704 (
		_w27207_,
		_w27216_,
		_w27217_
	);
	LUT4 #(
		.INIT('h0200)
	) name16705 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w27218_
	);
	LUT2 #(
		.INIT('h8)
	) name16706 (
		_w26361_,
		_w27218_,
		_w27219_
	);
	LUT4 #(
		.INIT('h0200)
	) name16707 (
		\ethreg1_TXCTRL_1_DataOut_reg[6]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w27220_
	);
	LUT4 #(
		.INIT('h0008)
	) name16708 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w27221_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16709 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w26358_,
		_w27220_,
		_w27221_,
		_w27222_
	);
	LUT2 #(
		.INIT('h4)
	) name16710 (
		_w27219_,
		_w27222_,
		_w27223_
	);
	LUT4 #(
		.INIT('h0008)
	) name16711 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w27224_
	);
	LUT4 #(
		.INIT('h0777)
	) name16712 (
		_w26359_,
		_w26366_,
		_w26370_,
		_w27224_,
		_w27225_
	);
	LUT4 #(
		.INIT('h0020)
	) name16713 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w27226_
	);
	LUT4 #(
		.INIT('h0200)
	) name16714 (
		\ethreg1_TXCTRL_0_DataOut_reg[6]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w27227_
	);
	LUT4 #(
		.INIT('h153f)
	) name16715 (
		_w25925_,
		_w26365_,
		_w27226_,
		_w27227_,
		_w27228_
	);
	LUT4 #(
		.INIT('h0020)
	) name16716 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w27229_
	);
	LUT4 #(
		.INIT('h0020)
	) name16717 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w27230_
	);
	LUT4 #(
		.INIT('h135f)
	) name16718 (
		_w26361_,
		_w26370_,
		_w27229_,
		_w27230_,
		_w27231_
	);
	LUT3 #(
		.INIT('h80)
	) name16719 (
		_w27225_,
		_w27228_,
		_w27231_,
		_w27232_
	);
	LUT2 #(
		.INIT('h7)
	) name16720 (
		_w27223_,
		_w27232_,
		_w27233_
	);
	LUT2 #(
		.INIT('h8)
	) name16721 (
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		\txethmac1_random1_x_reg[6]/NET0131 ,
		_w27234_
	);
	LUT4 #(
		.INIT('h8000)
	) name16722 (
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		\txethmac1_random1_x_reg[6]/NET0131 ,
		_w27235_
	);
	LUT4 #(
		.INIT('heee2)
	) name16723 (
		\txethmac1_random1_RandomLatched_reg[6]/NET0131 ,
		_w26376_,
		_w27234_,
		_w27235_,
		_w27236_
	);
	LUT2 #(
		.INIT('h4)
	) name16724 (
		\wishbone_BlockingTxBDRead_reg/NET0131 ,
		\wishbone_TxRetryPacket_NotCleared_reg/NET0131 ,
		_w27237_
	);
	LUT2 #(
		.INIT('h1)
	) name16725 (
		\wishbone_BlockingTxBDRead_reg/NET0131 ,
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		_w27238_
	);
	LUT4 #(
		.INIT('h0105)
	) name16726 (
		\wishbone_TxBDRead_reg/NET0131 ,
		_w26321_,
		_w27237_,
		_w27238_,
		_w27239_
	);
	LUT2 #(
		.INIT('h1)
	) name16727 (
		\wishbone_TxBDReady_reg/NET0131 ,
		_w27239_,
		_w27240_
	);
	LUT4 #(
		.INIT('h5450)
	) name16728 (
		\wishbone_TxBDReady_reg/NET0131 ,
		_w26321_,
		_w27237_,
		_w27238_,
		_w27241_
	);
	LUT2 #(
		.INIT('h4)
	) name16729 (
		\wishbone_TxRetryPacketBlocked_reg/NET0131 ,
		\wishbone_TxRetry_wb_reg/NET0131 ,
		_w27242_
	);
	LUT3 #(
		.INIT('h23)
	) name16730 (
		\wishbone_TxRetryPacketBlocked_reg/NET0131 ,
		\wishbone_TxRetryPacket_NotCleared_reg/NET0131 ,
		\wishbone_TxRetry_wb_reg/NET0131 ,
		_w27243_
	);
	LUT2 #(
		.INIT('h2)
	) name16731 (
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_TxRetryPacket_NotCleared_reg/NET0131 ,
		_w27244_
	);
	LUT3 #(
		.INIT('h23)
	) name16732 (
		_w27095_,
		_w27243_,
		_w27244_,
		_w27245_
	);
	LUT2 #(
		.INIT('h4)
	) name16733 (
		_w27241_,
		_w27245_,
		_w27246_
	);
	LUT4 #(
		.INIT('h0208)
	) name16734 (
		\wishbone_LastWord_reg/NET0131 ,
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxEndFrm_reg/NET0131 ,
		\wishbone_TxValidBytesLatched_reg[0]/NET0131 ,
		_w27247_
	);
	LUT4 #(
		.INIT('h7dd7)
	) name16735 (
		\wishbone_Flop_reg/NET0131 ,
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		\wishbone_TxValidBytesLatched_reg[1]/NET0131 ,
		_w27248_
	);
	LUT3 #(
		.INIT('hd0)
	) name16736 (
		\wishbone_Flop_reg/NET0131 ,
		_w27247_,
		_w27248_,
		_w27249_
	);
	LUT2 #(
		.INIT('h2)
	) name16737 (
		_w27064_,
		_w27065_,
		_w27250_
	);
	LUT3 #(
		.INIT('h0e)
	) name16738 (
		\wishbone_Flop_reg/NET0131 ,
		\wishbone_TxEndFrm_reg/NET0131 ,
		\wishbone_TxRetry_q_reg/NET0131 ,
		_w27251_
	);
	LUT3 #(
		.INIT('hd0)
	) name16739 (
		_w27064_,
		_w27065_,
		_w27251_,
		_w27252_
	);
	LUT2 #(
		.INIT('h8)
	) name16740 (
		_w27249_,
		_w27252_,
		_w27253_
	);
	LUT2 #(
		.INIT('h8)
	) name16741 (
		\wishbone_WbEn_q_reg/NET0131 ,
		\wishbone_WbEn_reg/NET0131 ,
		_w27254_
	);
	LUT3 #(
		.INIT('h80)
	) name16742 (
		\wishbone_BDWrite_reg[1]/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		\wishbone_WbEn_reg/NET0131 ,
		_w27255_
	);
	LUT4 #(
		.INIT('h0023)
	) name16743 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		_w25879_,
		_w26321_,
		_w27255_,
		_w27256_
	);
	LUT4 #(
		.INIT('h0200)
	) name16744 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27257_
	);
	LUT4 #(
		.INIT('h0020)
	) name16745 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27258_
	);
	LUT2 #(
		.INIT('h8)
	) name16746 (
		_w27257_,
		_w27258_,
		_w27259_
	);
	LUT2 #(
		.INIT('h4)
	) name16747 (
		_w27256_,
		_w27259_,
		_w27260_
	);
	LUT3 #(
		.INIT('h80)
	) name16748 (
		\wishbone_BDWrite_reg[2]/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		\wishbone_WbEn_reg/NET0131 ,
		_w27261_
	);
	LUT4 #(
		.INIT('h0023)
	) name16749 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		_w25879_,
		_w26321_,
		_w27261_,
		_w27262_
	);
	LUT4 #(
		.INIT('h0040)
	) name16750 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27263_
	);
	LUT2 #(
		.INIT('h8)
	) name16751 (
		_w27257_,
		_w27263_,
		_w27264_
	);
	LUT2 #(
		.INIT('h4)
	) name16752 (
		_w27262_,
		_w27264_,
		_w27265_
	);
	LUT4 #(
		.INIT('h0080)
	) name16753 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27266_
	);
	LUT4 #(
		.INIT('h0100)
	) name16754 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27267_
	);
	LUT2 #(
		.INIT('h8)
	) name16755 (
		_w27266_,
		_w27267_,
		_w27268_
	);
	LUT2 #(
		.INIT('h4)
	) name16756 (
		_w27262_,
		_w27268_,
		_w27269_
	);
	LUT4 #(
		.INIT('h0800)
	) name16757 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27270_
	);
	LUT4 #(
		.INIT('h0010)
	) name16758 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27271_
	);
	LUT2 #(
		.INIT('h8)
	) name16759 (
		_w27270_,
		_w27271_,
		_w27272_
	);
	LUT2 #(
		.INIT('h4)
	) name16760 (
		_w27262_,
		_w27272_,
		_w27273_
	);
	LUT4 #(
		.INIT('h0400)
	) name16761 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27274_
	);
	LUT2 #(
		.INIT('h8)
	) name16762 (
		_w27258_,
		_w27274_,
		_w27275_
	);
	LUT2 #(
		.INIT('h4)
	) name16763 (
		_w27262_,
		_w27275_,
		_w27276_
	);
	LUT2 #(
		.INIT('h8)
	) name16764 (
		_w27263_,
		_w27274_,
		_w27277_
	);
	LUT2 #(
		.INIT('h4)
	) name16765 (
		_w27262_,
		_w27277_,
		_w27278_
	);
	LUT3 #(
		.INIT('h80)
	) name16766 (
		\wishbone_BDWrite_reg[0]/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		\wishbone_WbEn_reg/NET0131 ,
		_w27279_
	);
	LUT4 #(
		.INIT('h0023)
	) name16767 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		_w25879_,
		_w26321_,
		_w27279_,
		_w27280_
	);
	LUT4 #(
		.INIT('h0002)
	) name16768 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27281_
	);
	LUT4 #(
		.INIT('h8000)
	) name16769 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27282_
	);
	LUT2 #(
		.INIT('h8)
	) name16770 (
		_w27281_,
		_w27282_,
		_w27283_
	);
	LUT2 #(
		.INIT('h4)
	) name16771 (
		_w27280_,
		_w27283_,
		_w27284_
	);
	LUT4 #(
		.INIT('h2000)
	) name16772 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27285_
	);
	LUT2 #(
		.INIT('h8)
	) name16773 (
		_w27271_,
		_w27285_,
		_w27286_
	);
	LUT2 #(
		.INIT('h4)
	) name16774 (
		_w27262_,
		_w27286_,
		_w27287_
	);
	LUT4 #(
		.INIT('h1000)
	) name16775 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27288_
	);
	LUT2 #(
		.INIT('h8)
	) name16776 (
		_w27258_,
		_w27288_,
		_w27289_
	);
	LUT2 #(
		.INIT('h4)
	) name16777 (
		_w27262_,
		_w27289_,
		_w27290_
	);
	LUT2 #(
		.INIT('h8)
	) name16778 (
		_w27263_,
		_w27288_,
		_w27291_
	);
	LUT2 #(
		.INIT('h4)
	) name16779 (
		_w27262_,
		_w27291_,
		_w27292_
	);
	LUT4 #(
		.INIT('h4000)
	) name16780 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27293_
	);
	LUT2 #(
		.INIT('h8)
	) name16781 (
		_w27271_,
		_w27293_,
		_w27294_
	);
	LUT2 #(
		.INIT('h4)
	) name16782 (
		_w27262_,
		_w27294_,
		_w27295_
	);
	LUT2 #(
		.INIT('h8)
	) name16783 (
		_w27271_,
		_w27282_,
		_w27296_
	);
	LUT2 #(
		.INIT('h4)
	) name16784 (
		_w27262_,
		_w27296_,
		_w27297_
	);
	LUT4 #(
		.INIT('h0800)
	) name16785 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27298_
	);
	LUT4 #(
		.INIT('h0001)
	) name16786 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27299_
	);
	LUT2 #(
		.INIT('h8)
	) name16787 (
		_w27298_,
		_w27299_,
		_w27300_
	);
	LUT2 #(
		.INIT('h4)
	) name16788 (
		_w27262_,
		_w27300_,
		_w27301_
	);
	LUT4 #(
		.INIT('h0002)
	) name16789 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27302_
	);
	LUT2 #(
		.INIT('h8)
	) name16790 (
		_w27298_,
		_w27302_,
		_w27303_
	);
	LUT2 #(
		.INIT('h4)
	) name16791 (
		_w27262_,
		_w27303_,
		_w27304_
	);
	LUT4 #(
		.INIT('h0200)
	) name16792 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27305_
	);
	LUT4 #(
		.INIT('h0008)
	) name16793 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27306_
	);
	LUT2 #(
		.INIT('h8)
	) name16794 (
		_w27305_,
		_w27306_,
		_w27307_
	);
	LUT2 #(
		.INIT('h4)
	) name16795 (
		_w27262_,
		_w27307_,
		_w27308_
	);
	LUT4 #(
		.INIT('h0400)
	) name16796 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27309_
	);
	LUT2 #(
		.INIT('h8)
	) name16797 (
		_w27306_,
		_w27309_,
		_w27310_
	);
	LUT2 #(
		.INIT('h4)
	) name16798 (
		_w27262_,
		_w27310_,
		_w27311_
	);
	LUT4 #(
		.INIT('h0004)
	) name16799 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27312_
	);
	LUT2 #(
		.INIT('h8)
	) name16800 (
		_w27298_,
		_w27312_,
		_w27313_
	);
	LUT2 #(
		.INIT('h4)
	) name16801 (
		_w27262_,
		_w27313_,
		_w27314_
	);
	LUT4 #(
		.INIT('h0020)
	) name16802 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27315_
	);
	LUT2 #(
		.INIT('h8)
	) name16803 (
		_w27305_,
		_w27315_,
		_w27316_
	);
	LUT2 #(
		.INIT('h4)
	) name16804 (
		_w27262_,
		_w27316_,
		_w27317_
	);
	LUT2 #(
		.INIT('h8)
	) name16805 (
		_w27309_,
		_w27315_,
		_w27318_
	);
	LUT2 #(
		.INIT('h4)
	) name16806 (
		_w27262_,
		_w27318_,
		_w27319_
	);
	LUT4 #(
		.INIT('h0010)
	) name16807 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27320_
	);
	LUT2 #(
		.INIT('h8)
	) name16808 (
		_w27298_,
		_w27320_,
		_w27321_
	);
	LUT2 #(
		.INIT('h4)
	) name16809 (
		_w27262_,
		_w27321_,
		_w27322_
	);
	LUT2 #(
		.INIT('h4)
	) name16810 (
		_w27256_,
		_w27300_,
		_w27323_
	);
	LUT4 #(
		.INIT('h0100)
	) name16811 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27324_
	);
	LUT4 #(
		.INIT('h0080)
	) name16812 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27325_
	);
	LUT2 #(
		.INIT('h8)
	) name16813 (
		_w27324_,
		_w27325_,
		_w27326_
	);
	LUT2 #(
		.INIT('h4)
	) name16814 (
		_w27262_,
		_w27326_,
		_w27327_
	);
	LUT4 #(
		.INIT('h0040)
	) name16815 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w27328_
	);
	LUT2 #(
		.INIT('h8)
	) name16816 (
		_w27305_,
		_w27328_,
		_w27329_
	);
	LUT2 #(
		.INIT('h4)
	) name16817 (
		_w27262_,
		_w27329_,
		_w27330_
	);
	LUT2 #(
		.INIT('h8)
	) name16818 (
		_w27309_,
		_w27328_,
		_w27331_
	);
	LUT2 #(
		.INIT('h4)
	) name16819 (
		_w27262_,
		_w27331_,
		_w27332_
	);
	LUT4 #(
		.INIT('h0008)
	) name16820 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27333_
	);
	LUT2 #(
		.INIT('h8)
	) name16821 (
		_w27306_,
		_w27333_,
		_w27334_
	);
	LUT2 #(
		.INIT('h4)
	) name16822 (
		_w27262_,
		_w27334_,
		_w27335_
	);
	LUT4 #(
		.INIT('h2000)
	) name16823 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27336_
	);
	LUT2 #(
		.INIT('h8)
	) name16824 (
		_w27299_,
		_w27336_,
		_w27337_
	);
	LUT2 #(
		.INIT('h4)
	) name16825 (
		_w27262_,
		_w27337_,
		_w27338_
	);
	LUT2 #(
		.INIT('h8)
	) name16826 (
		_w27302_,
		_w27336_,
		_w27339_
	);
	LUT2 #(
		.INIT('h4)
	) name16827 (
		_w27262_,
		_w27339_,
		_w27340_
	);
	LUT4 #(
		.INIT('h4000)
	) name16828 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27341_
	);
	LUT2 #(
		.INIT('h8)
	) name16829 (
		_w27299_,
		_w27341_,
		_w27342_
	);
	LUT2 #(
		.INIT('h4)
	) name16830 (
		_w27262_,
		_w27342_,
		_w27343_
	);
	LUT2 #(
		.INIT('h8)
	) name16831 (
		_w27302_,
		_w27341_,
		_w27344_
	);
	LUT2 #(
		.INIT('h4)
	) name16832 (
		_w27262_,
		_w27344_,
		_w27345_
	);
	LUT4 #(
		.INIT('h8000)
	) name16833 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27346_
	);
	LUT2 #(
		.INIT('h8)
	) name16834 (
		_w27299_,
		_w27346_,
		_w27347_
	);
	LUT2 #(
		.INIT('h4)
	) name16835 (
		_w27262_,
		_w27347_,
		_w27348_
	);
	LUT2 #(
		.INIT('h8)
	) name16836 (
		_w27302_,
		_w27346_,
		_w27349_
	);
	LUT2 #(
		.INIT('h4)
	) name16837 (
		_w27262_,
		_w27349_,
		_w27350_
	);
	LUT4 #(
		.INIT('h1000)
	) name16838 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27351_
	);
	LUT2 #(
		.INIT('h8)
	) name16839 (
		_w27306_,
		_w27351_,
		_w27352_
	);
	LUT2 #(
		.INIT('h4)
	) name16840 (
		_w27262_,
		_w27352_,
		_w27353_
	);
	LUT2 #(
		.INIT('h8)
	) name16841 (
		_w27312_,
		_w27336_,
		_w27354_
	);
	LUT2 #(
		.INIT('h4)
	) name16842 (
		_w27262_,
		_w27354_,
		_w27355_
	);
	LUT2 #(
		.INIT('h8)
	) name16843 (
		_w27312_,
		_w27341_,
		_w27356_
	);
	LUT2 #(
		.INIT('h4)
	) name16844 (
		_w27262_,
		_w27356_,
		_w27357_
	);
	LUT2 #(
		.INIT('h8)
	) name16845 (
		_w27312_,
		_w27346_,
		_w27358_
	);
	LUT2 #(
		.INIT('h4)
	) name16846 (
		_w27262_,
		_w27358_,
		_w27359_
	);
	LUT2 #(
		.INIT('h8)
	) name16847 (
		_w27315_,
		_w27351_,
		_w27360_
	);
	LUT2 #(
		.INIT('h4)
	) name16848 (
		_w27262_,
		_w27360_,
		_w27361_
	);
	LUT2 #(
		.INIT('h8)
	) name16849 (
		_w27320_,
		_w27336_,
		_w27362_
	);
	LUT2 #(
		.INIT('h4)
	) name16850 (
		_w27262_,
		_w27362_,
		_w27363_
	);
	LUT2 #(
		.INIT('h8)
	) name16851 (
		_w27320_,
		_w27341_,
		_w27364_
	);
	LUT2 #(
		.INIT('h4)
	) name16852 (
		_w27262_,
		_w27364_,
		_w27365_
	);
	LUT2 #(
		.INIT('h8)
	) name16853 (
		_w27320_,
		_w27346_,
		_w27366_
	);
	LUT2 #(
		.INIT('h4)
	) name16854 (
		_w27262_,
		_w27366_,
		_w27367_
	);
	LUT2 #(
		.INIT('h8)
	) name16855 (
		_w27328_,
		_w27351_,
		_w27368_
	);
	LUT2 #(
		.INIT('h4)
	) name16856 (
		_w27262_,
		_w27368_,
		_w27369_
	);
	LUT2 #(
		.INIT('h8)
	) name16857 (
		_w27257_,
		_w27305_,
		_w27370_
	);
	LUT2 #(
		.INIT('h4)
	) name16858 (
		_w27262_,
		_w27370_,
		_w27371_
	);
	LUT2 #(
		.INIT('h8)
	) name16859 (
		_w27257_,
		_w27309_,
		_w27372_
	);
	LUT2 #(
		.INIT('h4)
	) name16860 (
		_w27262_,
		_w27372_,
		_w27373_
	);
	LUT2 #(
		.INIT('h8)
	) name16861 (
		_w27267_,
		_w27298_,
		_w27374_
	);
	LUT2 #(
		.INIT('h4)
	) name16862 (
		_w27262_,
		_w27374_,
		_w27375_
	);
	LUT2 #(
		.INIT('h8)
	) name16863 (
		_w27270_,
		_w27324_,
		_w27376_
	);
	LUT2 #(
		.INIT('h4)
	) name16864 (
		_w27262_,
		_w27376_,
		_w27377_
	);
	LUT2 #(
		.INIT('h8)
	) name16865 (
		_w27274_,
		_w27305_,
		_w27378_
	);
	LUT2 #(
		.INIT('h4)
	) name16866 (
		_w27262_,
		_w27378_,
		_w27379_
	);
	LUT2 #(
		.INIT('h8)
	) name16867 (
		_w27274_,
		_w27309_,
		_w27380_
	);
	LUT2 #(
		.INIT('h4)
	) name16868 (
		_w27262_,
		_w27380_,
		_w27381_
	);
	LUT2 #(
		.INIT('h8)
	) name16869 (
		_w27285_,
		_w27324_,
		_w27382_
	);
	LUT2 #(
		.INIT('h4)
	) name16870 (
		_w27262_,
		_w27382_,
		_w27383_
	);
	LUT2 #(
		.INIT('h8)
	) name16871 (
		_w27288_,
		_w27305_,
		_w27384_
	);
	LUT2 #(
		.INIT('h4)
	) name16872 (
		_w27262_,
		_w27384_,
		_w27385_
	);
	LUT2 #(
		.INIT('h8)
	) name16873 (
		_w27288_,
		_w27309_,
		_w27386_
	);
	LUT2 #(
		.INIT('h4)
	) name16874 (
		_w27262_,
		_w27386_,
		_w27387_
	);
	LUT2 #(
		.INIT('h8)
	) name16875 (
		_w27293_,
		_w27324_,
		_w27388_
	);
	LUT2 #(
		.INIT('h4)
	) name16876 (
		_w27262_,
		_w27388_,
		_w27389_
	);
	LUT2 #(
		.INIT('h8)
	) name16877 (
		_w27282_,
		_w27324_,
		_w27390_
	);
	LUT2 #(
		.INIT('h4)
	) name16878 (
		_w27262_,
		_w27390_,
		_w27391_
	);
	LUT2 #(
		.INIT('h4)
	) name16879 (
		_w27256_,
		_w27303_,
		_w27392_
	);
	LUT2 #(
		.INIT('h8)
	) name16880 (
		_w27257_,
		_w27351_,
		_w27393_
	);
	LUT2 #(
		.INIT('h4)
	) name16881 (
		_w27262_,
		_w27393_,
		_w27394_
	);
	LUT2 #(
		.INIT('h8)
	) name16882 (
		_w27267_,
		_w27336_,
		_w27395_
	);
	LUT2 #(
		.INIT('h4)
	) name16883 (
		_w27262_,
		_w27395_,
		_w27396_
	);
	LUT2 #(
		.INIT('h2)
	) name16884 (
		_w27264_,
		_w27280_,
		_w27397_
	);
	LUT2 #(
		.INIT('h8)
	) name16885 (
		_w27267_,
		_w27341_,
		_w27398_
	);
	LUT2 #(
		.INIT('h4)
	) name16886 (
		_w27262_,
		_w27398_,
		_w27399_
	);
	LUT2 #(
		.INIT('h2)
	) name16887 (
		_w27268_,
		_w27280_,
		_w27400_
	);
	LUT2 #(
		.INIT('h8)
	) name16888 (
		_w27267_,
		_w27346_,
		_w27401_
	);
	LUT2 #(
		.INIT('h4)
	) name16889 (
		_w27262_,
		_w27401_,
		_w27402_
	);
	LUT2 #(
		.INIT('h8)
	) name16890 (
		_w27274_,
		_w27351_,
		_w27403_
	);
	LUT2 #(
		.INIT('h4)
	) name16891 (
		_w27262_,
		_w27403_,
		_w27404_
	);
	LUT2 #(
		.INIT('h2)
	) name16892 (
		_w27272_,
		_w27280_,
		_w27405_
	);
	LUT2 #(
		.INIT('h2)
	) name16893 (
		_w27275_,
		_w27280_,
		_w27406_
	);
	LUT2 #(
		.INIT('h8)
	) name16894 (
		_w27315_,
		_w27333_,
		_w27407_
	);
	LUT2 #(
		.INIT('h4)
	) name16895 (
		_w27262_,
		_w27407_,
		_w27408_
	);
	LUT2 #(
		.INIT('h2)
	) name16896 (
		_w27277_,
		_w27280_,
		_w27409_
	);
	LUT2 #(
		.INIT('h8)
	) name16897 (
		_w27288_,
		_w27351_,
		_w27410_
	);
	LUT2 #(
		.INIT('h4)
	) name16898 (
		_w27262_,
		_w27410_,
		_w27411_
	);
	LUT2 #(
		.INIT('h4)
	) name16899 (
		_w27280_,
		_w27286_,
		_w27412_
	);
	LUT4 #(
		.INIT('h0004)
	) name16900 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27413_
	);
	LUT2 #(
		.INIT('h8)
	) name16901 (
		_w27270_,
		_w27413_,
		_w27414_
	);
	LUT2 #(
		.INIT('h4)
	) name16902 (
		_w27280_,
		_w27414_,
		_w27415_
	);
	LUT2 #(
		.INIT('h4)
	) name16903 (
		_w27280_,
		_w27289_,
		_w27416_
	);
	LUT4 #(
		.INIT('h0001)
	) name16904 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w27417_
	);
	LUT2 #(
		.INIT('h8)
	) name16905 (
		_w27325_,
		_w27417_,
		_w27418_
	);
	LUT2 #(
		.INIT('h4)
	) name16906 (
		_w27262_,
		_w27418_,
		_w27419_
	);
	LUT2 #(
		.INIT('h4)
	) name16907 (
		_w27280_,
		_w27291_,
		_w27420_
	);
	LUT2 #(
		.INIT('h8)
	) name16908 (
		_w27281_,
		_w27325_,
		_w27421_
	);
	LUT2 #(
		.INIT('h4)
	) name16909 (
		_w27262_,
		_w27421_,
		_w27422_
	);
	LUT2 #(
		.INIT('h8)
	) name16910 (
		_w27325_,
		_w27413_,
		_w27423_
	);
	LUT2 #(
		.INIT('h4)
	) name16911 (
		_w27262_,
		_w27423_,
		_w27424_
	);
	LUT2 #(
		.INIT('h8)
	) name16912 (
		_w27328_,
		_w27333_,
		_w27425_
	);
	LUT2 #(
		.INIT('h4)
	) name16913 (
		_w27262_,
		_w27425_,
		_w27426_
	);
	LUT2 #(
		.INIT('h4)
	) name16914 (
		_w27280_,
		_w27294_,
		_w27427_
	);
	LUT2 #(
		.INIT('h4)
	) name16915 (
		_w27280_,
		_w27296_,
		_w27428_
	);
	LUT2 #(
		.INIT('h8)
	) name16916 (
		_w27266_,
		_w27299_,
		_w27429_
	);
	LUT2 #(
		.INIT('h4)
	) name16917 (
		_w27262_,
		_w27429_,
		_w27430_
	);
	LUT2 #(
		.INIT('h8)
	) name16918 (
		_w27266_,
		_w27302_,
		_w27431_
	);
	LUT2 #(
		.INIT('h4)
	) name16919 (
		_w27262_,
		_w27431_,
		_w27432_
	);
	LUT2 #(
		.INIT('h8)
	) name16920 (
		_w27258_,
		_w27306_,
		_w27433_
	);
	LUT2 #(
		.INIT('h4)
	) name16921 (
		_w27262_,
		_w27433_,
		_w27434_
	);
	LUT2 #(
		.INIT('h8)
	) name16922 (
		_w27263_,
		_w27306_,
		_w27435_
	);
	LUT2 #(
		.INIT('h4)
	) name16923 (
		_w27262_,
		_w27435_,
		_w27436_
	);
	LUT2 #(
		.INIT('h8)
	) name16924 (
		_w27266_,
		_w27312_,
		_w27437_
	);
	LUT2 #(
		.INIT('h4)
	) name16925 (
		_w27262_,
		_w27437_,
		_w27438_
	);
	LUT2 #(
		.INIT('h8)
	) name16926 (
		_w27258_,
		_w27315_,
		_w27439_
	);
	LUT2 #(
		.INIT('h4)
	) name16927 (
		_w27262_,
		_w27439_,
		_w27440_
	);
	LUT2 #(
		.INIT('h8)
	) name16928 (
		_w27263_,
		_w27315_,
		_w27441_
	);
	LUT2 #(
		.INIT('h4)
	) name16929 (
		_w27262_,
		_w27441_,
		_w27442_
	);
	LUT2 #(
		.INIT('h8)
	) name16930 (
		_w27266_,
		_w27320_,
		_w27443_
	);
	LUT2 #(
		.INIT('h4)
	) name16931 (
		_w27262_,
		_w27443_,
		_w27444_
	);
	LUT2 #(
		.INIT('h8)
	) name16932 (
		_w27271_,
		_w27325_,
		_w27445_
	);
	LUT2 #(
		.INIT('h4)
	) name16933 (
		_w27262_,
		_w27445_,
		_w27446_
	);
	LUT2 #(
		.INIT('h8)
	) name16934 (
		_w27258_,
		_w27328_,
		_w27447_
	);
	LUT2 #(
		.INIT('h4)
	) name16935 (
		_w27262_,
		_w27447_,
		_w27448_
	);
	LUT2 #(
		.INIT('h8)
	) name16936 (
		_w27263_,
		_w27328_,
		_w27449_
	);
	LUT2 #(
		.INIT('h4)
	) name16937 (
		_w27262_,
		_w27449_,
		_w27450_
	);
	LUT2 #(
		.INIT('h4)
	) name16938 (
		_w27280_,
		_w27300_,
		_w27451_
	);
	LUT2 #(
		.INIT('h4)
	) name16939 (
		_w27280_,
		_w27303_,
		_w27452_
	);
	LUT2 #(
		.INIT('h8)
	) name16940 (
		_w27257_,
		_w27333_,
		_w27453_
	);
	LUT2 #(
		.INIT('h4)
	) name16941 (
		_w27262_,
		_w27453_,
		_w27454_
	);
	LUT2 #(
		.INIT('h4)
	) name16942 (
		_w27280_,
		_w27307_,
		_w27455_
	);
	LUT2 #(
		.INIT('h8)
	) name16943 (
		_w27270_,
		_w27417_,
		_w27456_
	);
	LUT2 #(
		.INIT('h4)
	) name16944 (
		_w27262_,
		_w27456_,
		_w27457_
	);
	LUT2 #(
		.INIT('h8)
	) name16945 (
		_w27270_,
		_w27281_,
		_w27458_
	);
	LUT2 #(
		.INIT('h4)
	) name16946 (
		_w27262_,
		_w27458_,
		_w27459_
	);
	LUT2 #(
		.INIT('h4)
	) name16947 (
		_w27262_,
		_w27414_,
		_w27460_
	);
	LUT2 #(
		.INIT('h8)
	) name16948 (
		_w27274_,
		_w27333_,
		_w27461_
	);
	LUT2 #(
		.INIT('h4)
	) name16949 (
		_w27262_,
		_w27461_,
		_w27462_
	);
	LUT2 #(
		.INIT('h4)
	) name16950 (
		_w27280_,
		_w27310_,
		_w27463_
	);
	LUT2 #(
		.INIT('h4)
	) name16951 (
		_w27280_,
		_w27313_,
		_w27464_
	);
	LUT2 #(
		.INIT('h8)
	) name16952 (
		_w27285_,
		_w27417_,
		_w27465_
	);
	LUT2 #(
		.INIT('h4)
	) name16953 (
		_w27262_,
		_w27465_,
		_w27466_
	);
	LUT2 #(
		.INIT('h8)
	) name16954 (
		_w27281_,
		_w27285_,
		_w27467_
	);
	LUT2 #(
		.INIT('h4)
	) name16955 (
		_w27262_,
		_w27467_,
		_w27468_
	);
	LUT2 #(
		.INIT('h8)
	) name16956 (
		_w27285_,
		_w27413_,
		_w27469_
	);
	LUT2 #(
		.INIT('h4)
	) name16957 (
		_w27262_,
		_w27469_,
		_w27470_
	);
	LUT2 #(
		.INIT('h8)
	) name16958 (
		_w27288_,
		_w27333_,
		_w27471_
	);
	LUT2 #(
		.INIT('h4)
	) name16959 (
		_w27262_,
		_w27471_,
		_w27472_
	);
	LUT2 #(
		.INIT('h8)
	) name16960 (
		_w27293_,
		_w27417_,
		_w27473_
	);
	LUT2 #(
		.INIT('h4)
	) name16961 (
		_w27262_,
		_w27473_,
		_w27474_
	);
	LUT2 #(
		.INIT('h8)
	) name16962 (
		_w27282_,
		_w27417_,
		_w27475_
	);
	LUT2 #(
		.INIT('h4)
	) name16963 (
		_w27262_,
		_w27475_,
		_w27476_
	);
	LUT2 #(
		.INIT('h4)
	) name16964 (
		_w27280_,
		_w27316_,
		_w27477_
	);
	LUT2 #(
		.INIT('h8)
	) name16965 (
		_w27281_,
		_w27293_,
		_w27478_
	);
	LUT2 #(
		.INIT('h4)
	) name16966 (
		_w27262_,
		_w27478_,
		_w27479_
	);
	LUT2 #(
		.INIT('h4)
	) name16967 (
		_w27262_,
		_w27283_,
		_w27480_
	);
	LUT2 #(
		.INIT('h8)
	) name16968 (
		_w27293_,
		_w27413_,
		_w27481_
	);
	LUT2 #(
		.INIT('h4)
	) name16969 (
		_w27262_,
		_w27481_,
		_w27482_
	);
	LUT2 #(
		.INIT('h4)
	) name16970 (
		_w27280_,
		_w27318_,
		_w27483_
	);
	LUT2 #(
		.INIT('h8)
	) name16971 (
		_w27282_,
		_w27413_,
		_w27484_
	);
	LUT2 #(
		.INIT('h4)
	) name16972 (
		_w27262_,
		_w27484_,
		_w27485_
	);
	LUT2 #(
		.INIT('h4)
	) name16973 (
		_w27280_,
		_w27321_,
		_w27486_
	);
	LUT2 #(
		.INIT('h2)
	) name16974 (
		_w27259_,
		_w27262_,
		_w27487_
	);
	LUT2 #(
		.INIT('h4)
	) name16975 (
		_w27280_,
		_w27326_,
		_w27488_
	);
	LUT3 #(
		.INIT('h80)
	) name16976 (
		\wishbone_BDWrite_reg[3]/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		\wishbone_WbEn_reg/NET0131 ,
		_w27489_
	);
	LUT4 #(
		.INIT('h0023)
	) name16977 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		_w25879_,
		_w26321_,
		_w27489_,
		_w27490_
	);
	LUT2 #(
		.INIT('h2)
	) name16978 (
		_w27264_,
		_w27490_,
		_w27491_
	);
	LUT2 #(
		.INIT('h2)
	) name16979 (
		_w27268_,
		_w27490_,
		_w27492_
	);
	LUT2 #(
		.INIT('h4)
	) name16980 (
		_w27280_,
		_w27329_,
		_w27493_
	);
	LUT2 #(
		.INIT('h2)
	) name16981 (
		_w27272_,
		_w27490_,
		_w27494_
	);
	LUT2 #(
		.INIT('h2)
	) name16982 (
		_w27275_,
		_w27490_,
		_w27495_
	);
	LUT2 #(
		.INIT('h4)
	) name16983 (
		_w27280_,
		_w27331_,
		_w27496_
	);
	LUT2 #(
		.INIT('h2)
	) name16984 (
		_w27277_,
		_w27490_,
		_w27497_
	);
	LUT2 #(
		.INIT('h2)
	) name16985 (
		_w27286_,
		_w27490_,
		_w27498_
	);
	LUT2 #(
		.INIT('h4)
	) name16986 (
		_w27280_,
		_w27334_,
		_w27499_
	);
	LUT2 #(
		.INIT('h2)
	) name16987 (
		_w27289_,
		_w27490_,
		_w27500_
	);
	LUT2 #(
		.INIT('h2)
	) name16988 (
		_w27291_,
		_w27490_,
		_w27501_
	);
	LUT2 #(
		.INIT('h4)
	) name16989 (
		_w27280_,
		_w27337_,
		_w27502_
	);
	LUT2 #(
		.INIT('h2)
	) name16990 (
		_w27294_,
		_w27490_,
		_w27503_
	);
	LUT2 #(
		.INIT('h2)
	) name16991 (
		_w27296_,
		_w27490_,
		_w27504_
	);
	LUT2 #(
		.INIT('h4)
	) name16992 (
		_w27280_,
		_w27339_,
		_w27505_
	);
	LUT2 #(
		.INIT('h4)
	) name16993 (
		_w27280_,
		_w27342_,
		_w27506_
	);
	LUT2 #(
		.INIT('h4)
	) name16994 (
		_w27280_,
		_w27344_,
		_w27507_
	);
	LUT2 #(
		.INIT('h4)
	) name16995 (
		_w27280_,
		_w27347_,
		_w27508_
	);
	LUT2 #(
		.INIT('h4)
	) name16996 (
		_w27280_,
		_w27349_,
		_w27509_
	);
	LUT2 #(
		.INIT('h4)
	) name16997 (
		_w27280_,
		_w27352_,
		_w27510_
	);
	LUT2 #(
		.INIT('h2)
	) name16998 (
		_w27300_,
		_w27490_,
		_w27511_
	);
	LUT2 #(
		.INIT('h2)
	) name16999 (
		_w27303_,
		_w27490_,
		_w27512_
	);
	LUT2 #(
		.INIT('h4)
	) name17000 (
		_w27280_,
		_w27354_,
		_w27513_
	);
	LUT2 #(
		.INIT('h2)
	) name17001 (
		_w27307_,
		_w27490_,
		_w27514_
	);
	LUT2 #(
		.INIT('h4)
	) name17002 (
		_w27280_,
		_w27356_,
		_w27515_
	);
	LUT2 #(
		.INIT('h2)
	) name17003 (
		_w27310_,
		_w27490_,
		_w27516_
	);
	LUT2 #(
		.INIT('h2)
	) name17004 (
		_w27313_,
		_w27490_,
		_w27517_
	);
	LUT2 #(
		.INIT('h4)
	) name17005 (
		_w27280_,
		_w27358_,
		_w27518_
	);
	LUT2 #(
		.INIT('h2)
	) name17006 (
		_w27316_,
		_w27490_,
		_w27519_
	);
	LUT2 #(
		.INIT('h2)
	) name17007 (
		_w27318_,
		_w27490_,
		_w27520_
	);
	LUT2 #(
		.INIT('h4)
	) name17008 (
		_w27280_,
		_w27360_,
		_w27521_
	);
	LUT2 #(
		.INIT('h2)
	) name17009 (
		_w27321_,
		_w27490_,
		_w27522_
	);
	LUT2 #(
		.INIT('h4)
	) name17010 (
		_w27280_,
		_w27362_,
		_w27523_
	);
	LUT2 #(
		.INIT('h2)
	) name17011 (
		_w27326_,
		_w27490_,
		_w27524_
	);
	LUT2 #(
		.INIT('h2)
	) name17012 (
		_w27329_,
		_w27490_,
		_w27525_
	);
	LUT2 #(
		.INIT('h2)
	) name17013 (
		_w27331_,
		_w27490_,
		_w27526_
	);
	LUT2 #(
		.INIT('h4)
	) name17014 (
		_w27280_,
		_w27364_,
		_w27527_
	);
	LUT2 #(
		.INIT('h2)
	) name17015 (
		_w27334_,
		_w27490_,
		_w27528_
	);
	LUT2 #(
		.INIT('h4)
	) name17016 (
		_w27280_,
		_w27366_,
		_w27529_
	);
	LUT2 #(
		.INIT('h2)
	) name17017 (
		_w27337_,
		_w27490_,
		_w27530_
	);
	LUT2 #(
		.INIT('h2)
	) name17018 (
		_w27339_,
		_w27490_,
		_w27531_
	);
	LUT2 #(
		.INIT('h2)
	) name17019 (
		_w27342_,
		_w27490_,
		_w27532_
	);
	LUT2 #(
		.INIT('h4)
	) name17020 (
		_w27280_,
		_w27368_,
		_w27533_
	);
	LUT2 #(
		.INIT('h2)
	) name17021 (
		_w27344_,
		_w27490_,
		_w27534_
	);
	LUT2 #(
		.INIT('h2)
	) name17022 (
		_w27347_,
		_w27490_,
		_w27535_
	);
	LUT2 #(
		.INIT('h2)
	) name17023 (
		_w27349_,
		_w27490_,
		_w27536_
	);
	LUT2 #(
		.INIT('h2)
	) name17024 (
		_w27352_,
		_w27490_,
		_w27537_
	);
	LUT2 #(
		.INIT('h2)
	) name17025 (
		_w27354_,
		_w27490_,
		_w27538_
	);
	LUT2 #(
		.INIT('h2)
	) name17026 (
		_w27356_,
		_w27490_,
		_w27539_
	);
	LUT2 #(
		.INIT('h2)
	) name17027 (
		_w27358_,
		_w27490_,
		_w27540_
	);
	LUT2 #(
		.INIT('h2)
	) name17028 (
		_w27360_,
		_w27490_,
		_w27541_
	);
	LUT2 #(
		.INIT('h2)
	) name17029 (
		_w27362_,
		_w27490_,
		_w27542_
	);
	LUT2 #(
		.INIT('h2)
	) name17030 (
		_w27364_,
		_w27490_,
		_w27543_
	);
	LUT2 #(
		.INIT('h2)
	) name17031 (
		_w27366_,
		_w27490_,
		_w27544_
	);
	LUT2 #(
		.INIT('h2)
	) name17032 (
		_w27368_,
		_w27490_,
		_w27545_
	);
	LUT2 #(
		.INIT('h4)
	) name17033 (
		_w27280_,
		_w27370_,
		_w27546_
	);
	LUT2 #(
		.INIT('h4)
	) name17034 (
		_w27280_,
		_w27372_,
		_w27547_
	);
	LUT2 #(
		.INIT('h4)
	) name17035 (
		_w27280_,
		_w27374_,
		_w27548_
	);
	LUT2 #(
		.INIT('h2)
	) name17036 (
		_w27370_,
		_w27490_,
		_w27549_
	);
	LUT2 #(
		.INIT('h2)
	) name17037 (
		_w27372_,
		_w27490_,
		_w27550_
	);
	LUT2 #(
		.INIT('h2)
	) name17038 (
		_w27374_,
		_w27490_,
		_w27551_
	);
	LUT2 #(
		.INIT('h4)
	) name17039 (
		_w27280_,
		_w27376_,
		_w27552_
	);
	LUT2 #(
		.INIT('h2)
	) name17040 (
		_w27376_,
		_w27490_,
		_w27553_
	);
	LUT2 #(
		.INIT('h4)
	) name17041 (
		_w27280_,
		_w27378_,
		_w27554_
	);
	LUT2 #(
		.INIT('h2)
	) name17042 (
		_w27378_,
		_w27490_,
		_w27555_
	);
	LUT2 #(
		.INIT('h2)
	) name17043 (
		_w27380_,
		_w27490_,
		_w27556_
	);
	LUT2 #(
		.INIT('h4)
	) name17044 (
		_w27280_,
		_w27380_,
		_w27557_
	);
	LUT2 #(
		.INIT('h2)
	) name17045 (
		_w27382_,
		_w27490_,
		_w27558_
	);
	LUT2 #(
		.INIT('h2)
	) name17046 (
		_w27384_,
		_w27490_,
		_w27559_
	);
	LUT2 #(
		.INIT('h2)
	) name17047 (
		_w27386_,
		_w27490_,
		_w27560_
	);
	LUT2 #(
		.INIT('h4)
	) name17048 (
		_w27280_,
		_w27382_,
		_w27561_
	);
	LUT2 #(
		.INIT('h2)
	) name17049 (
		_w27388_,
		_w27490_,
		_w27562_
	);
	LUT2 #(
		.INIT('h2)
	) name17050 (
		_w27390_,
		_w27490_,
		_w27563_
	);
	LUT2 #(
		.INIT('h4)
	) name17051 (
		_w27280_,
		_w27384_,
		_w27564_
	);
	LUT2 #(
		.INIT('h4)
	) name17052 (
		_w27280_,
		_w27386_,
		_w27565_
	);
	LUT2 #(
		.INIT('h2)
	) name17053 (
		_w27393_,
		_w27490_,
		_w27566_
	);
	LUT2 #(
		.INIT('h2)
	) name17054 (
		_w27395_,
		_w27490_,
		_w27567_
	);
	LUT2 #(
		.INIT('h2)
	) name17055 (
		_w27398_,
		_w27490_,
		_w27568_
	);
	LUT2 #(
		.INIT('h4)
	) name17056 (
		_w27280_,
		_w27388_,
		_w27569_
	);
	LUT2 #(
		.INIT('h2)
	) name17057 (
		_w27401_,
		_w27490_,
		_w27570_
	);
	LUT2 #(
		.INIT('h4)
	) name17058 (
		_w27280_,
		_w27390_,
		_w27571_
	);
	LUT2 #(
		.INIT('h2)
	) name17059 (
		_w27403_,
		_w27490_,
		_w27572_
	);
	LUT2 #(
		.INIT('h2)
	) name17060 (
		_w27407_,
		_w27490_,
		_w27573_
	);
	LUT2 #(
		.INIT('h2)
	) name17061 (
		_w27410_,
		_w27490_,
		_w27574_
	);
	LUT2 #(
		.INIT('h4)
	) name17062 (
		_w27280_,
		_w27393_,
		_w27575_
	);
	LUT2 #(
		.INIT('h4)
	) name17063 (
		_w27280_,
		_w27395_,
		_w27576_
	);
	LUT2 #(
		.INIT('h4)
	) name17064 (
		_w27280_,
		_w27398_,
		_w27577_
	);
	LUT2 #(
		.INIT('h2)
	) name17065 (
		_w27418_,
		_w27490_,
		_w27578_
	);
	LUT2 #(
		.INIT('h2)
	) name17066 (
		_w27421_,
		_w27490_,
		_w27579_
	);
	LUT2 #(
		.INIT('h4)
	) name17067 (
		_w27280_,
		_w27401_,
		_w27580_
	);
	LUT2 #(
		.INIT('h2)
	) name17068 (
		_w27423_,
		_w27490_,
		_w27581_
	);
	LUT2 #(
		.INIT('h2)
	) name17069 (
		_w27425_,
		_w27490_,
		_w27582_
	);
	LUT2 #(
		.INIT('h4)
	) name17070 (
		_w27280_,
		_w27403_,
		_w27583_
	);
	LUT2 #(
		.INIT('h2)
	) name17071 (
		_w27429_,
		_w27490_,
		_w27584_
	);
	LUT2 #(
		.INIT('h2)
	) name17072 (
		_w27431_,
		_w27490_,
		_w27585_
	);
	LUT2 #(
		.INIT('h2)
	) name17073 (
		_w27433_,
		_w27490_,
		_w27586_
	);
	LUT2 #(
		.INIT('h2)
	) name17074 (
		_w27435_,
		_w27490_,
		_w27587_
	);
	LUT2 #(
		.INIT('h2)
	) name17075 (
		_w27437_,
		_w27490_,
		_w27588_
	);
	LUT2 #(
		.INIT('h4)
	) name17076 (
		_w27280_,
		_w27407_,
		_w27589_
	);
	LUT2 #(
		.INIT('h4)
	) name17077 (
		_w27280_,
		_w27410_,
		_w27590_
	);
	LUT2 #(
		.INIT('h2)
	) name17078 (
		_w27439_,
		_w27490_,
		_w27591_
	);
	LUT2 #(
		.INIT('h2)
	) name17079 (
		_w27441_,
		_w27490_,
		_w27592_
	);
	LUT2 #(
		.INIT('h2)
	) name17080 (
		_w27443_,
		_w27490_,
		_w27593_
	);
	LUT2 #(
		.INIT('h2)
	) name17081 (
		_w27445_,
		_w27490_,
		_w27594_
	);
	LUT2 #(
		.INIT('h2)
	) name17082 (
		_w27447_,
		_w27490_,
		_w27595_
	);
	LUT2 #(
		.INIT('h2)
	) name17083 (
		_w27449_,
		_w27490_,
		_w27596_
	);
	LUT2 #(
		.INIT('h2)
	) name17084 (
		_w27453_,
		_w27490_,
		_w27597_
	);
	LUT2 #(
		.INIT('h2)
	) name17085 (
		_w27456_,
		_w27490_,
		_w27598_
	);
	LUT2 #(
		.INIT('h2)
	) name17086 (
		_w27458_,
		_w27490_,
		_w27599_
	);
	LUT2 #(
		.INIT('h2)
	) name17087 (
		_w27414_,
		_w27490_,
		_w27600_
	);
	LUT2 #(
		.INIT('h2)
	) name17088 (
		_w27461_,
		_w27490_,
		_w27601_
	);
	LUT2 #(
		.INIT('h4)
	) name17089 (
		_w27280_,
		_w27418_,
		_w27602_
	);
	LUT2 #(
		.INIT('h2)
	) name17090 (
		_w27465_,
		_w27490_,
		_w27603_
	);
	LUT2 #(
		.INIT('h2)
	) name17091 (
		_w27467_,
		_w27490_,
		_w27604_
	);
	LUT2 #(
		.INIT('h4)
	) name17092 (
		_w27280_,
		_w27421_,
		_w27605_
	);
	LUT2 #(
		.INIT('h2)
	) name17093 (
		_w27469_,
		_w27490_,
		_w27606_
	);
	LUT2 #(
		.INIT('h2)
	) name17094 (
		_w27471_,
		_w27490_,
		_w27607_
	);
	LUT2 #(
		.INIT('h2)
	) name17095 (
		_w27473_,
		_w27490_,
		_w27608_
	);
	LUT2 #(
		.INIT('h4)
	) name17096 (
		_w27280_,
		_w27423_,
		_w27609_
	);
	LUT2 #(
		.INIT('h2)
	) name17097 (
		_w27475_,
		_w27490_,
		_w27610_
	);
	LUT2 #(
		.INIT('h2)
	) name17098 (
		_w27478_,
		_w27490_,
		_w27611_
	);
	LUT2 #(
		.INIT('h2)
	) name17099 (
		_w27283_,
		_w27490_,
		_w27612_
	);
	LUT2 #(
		.INIT('h4)
	) name17100 (
		_w27280_,
		_w27425_,
		_w27613_
	);
	LUT2 #(
		.INIT('h2)
	) name17101 (
		_w27481_,
		_w27490_,
		_w27614_
	);
	LUT2 #(
		.INIT('h2)
	) name17102 (
		_w27484_,
		_w27490_,
		_w27615_
	);
	LUT2 #(
		.INIT('h2)
	) name17103 (
		_w27259_,
		_w27490_,
		_w27616_
	);
	LUT2 #(
		.INIT('h4)
	) name17104 (
		_w27280_,
		_w27429_,
		_w27617_
	);
	LUT2 #(
		.INIT('h4)
	) name17105 (
		_w27280_,
		_w27431_,
		_w27618_
	);
	LUT2 #(
		.INIT('h4)
	) name17106 (
		_w27280_,
		_w27469_,
		_w27619_
	);
	LUT2 #(
		.INIT('h4)
	) name17107 (
		_w27280_,
		_w27433_,
		_w27620_
	);
	LUT2 #(
		.INIT('h4)
	) name17108 (
		_w27280_,
		_w27435_,
		_w27621_
	);
	LUT2 #(
		.INIT('h4)
	) name17109 (
		_w27280_,
		_w27437_,
		_w27622_
	);
	LUT2 #(
		.INIT('h4)
	) name17110 (
		_w27256_,
		_w27296_,
		_w27623_
	);
	LUT2 #(
		.INIT('h4)
	) name17111 (
		_w27280_,
		_w27439_,
		_w27624_
	);
	LUT2 #(
		.INIT('h4)
	) name17112 (
		_w27280_,
		_w27441_,
		_w27625_
	);
	LUT2 #(
		.INIT('h4)
	) name17113 (
		_w27280_,
		_w27443_,
		_w27626_
	);
	LUT2 #(
		.INIT('h4)
	) name17114 (
		_w27280_,
		_w27445_,
		_w27627_
	);
	LUT2 #(
		.INIT('h4)
	) name17115 (
		_w27280_,
		_w27447_,
		_w27628_
	);
	LUT2 #(
		.INIT('h4)
	) name17116 (
		_w27280_,
		_w27449_,
		_w27629_
	);
	LUT2 #(
		.INIT('h4)
	) name17117 (
		_w27280_,
		_w27453_,
		_w27630_
	);
	LUT2 #(
		.INIT('h4)
	) name17118 (
		_w27280_,
		_w27456_,
		_w27631_
	);
	LUT2 #(
		.INIT('h4)
	) name17119 (
		_w27280_,
		_w27481_,
		_w27632_
	);
	LUT2 #(
		.INIT('h4)
	) name17120 (
		_w27280_,
		_w27458_,
		_w27633_
	);
	LUT2 #(
		.INIT('h4)
	) name17121 (
		_w27280_,
		_w27461_,
		_w27634_
	);
	LUT2 #(
		.INIT('h4)
	) name17122 (
		_w27280_,
		_w27465_,
		_w27635_
	);
	LUT2 #(
		.INIT('h4)
	) name17123 (
		_w27280_,
		_w27467_,
		_w27636_
	);
	LUT2 #(
		.INIT('h4)
	) name17124 (
		_w27280_,
		_w27471_,
		_w27637_
	);
	LUT2 #(
		.INIT('h4)
	) name17125 (
		_w27280_,
		_w27473_,
		_w27638_
	);
	LUT2 #(
		.INIT('h4)
	) name17126 (
		_w27280_,
		_w27475_,
		_w27639_
	);
	LUT2 #(
		.INIT('h4)
	) name17127 (
		_w27280_,
		_w27478_,
		_w27640_
	);
	LUT2 #(
		.INIT('h4)
	) name17128 (
		_w27280_,
		_w27484_,
		_w27641_
	);
	LUT2 #(
		.INIT('h2)
	) name17129 (
		_w27259_,
		_w27280_,
		_w27642_
	);
	LUT2 #(
		.INIT('h4)
	) name17130 (
		_w27256_,
		_w27264_,
		_w27643_
	);
	LUT2 #(
		.INIT('h4)
	) name17131 (
		_w27256_,
		_w27268_,
		_w27644_
	);
	LUT2 #(
		.INIT('h4)
	) name17132 (
		_w27256_,
		_w27272_,
		_w27645_
	);
	LUT2 #(
		.INIT('h4)
	) name17133 (
		_w27256_,
		_w27275_,
		_w27646_
	);
	LUT2 #(
		.INIT('h4)
	) name17134 (
		_w27256_,
		_w27277_,
		_w27647_
	);
	LUT2 #(
		.INIT('h4)
	) name17135 (
		_w27256_,
		_w27294_,
		_w27648_
	);
	LUT2 #(
		.INIT('h4)
	) name17136 (
		_w27256_,
		_w27286_,
		_w27649_
	);
	LUT2 #(
		.INIT('h4)
	) name17137 (
		_w27256_,
		_w27289_,
		_w27650_
	);
	LUT2 #(
		.INIT('h4)
	) name17138 (
		_w27256_,
		_w27291_,
		_w27651_
	);
	LUT2 #(
		.INIT('h4)
	) name17139 (
		_w27256_,
		_w27307_,
		_w27652_
	);
	LUT2 #(
		.INIT('h4)
	) name17140 (
		_w27256_,
		_w27310_,
		_w27653_
	);
	LUT2 #(
		.INIT('h4)
	) name17141 (
		_w27256_,
		_w27313_,
		_w27654_
	);
	LUT2 #(
		.INIT('h4)
	) name17142 (
		_w27256_,
		_w27316_,
		_w27655_
	);
	LUT2 #(
		.INIT('h4)
	) name17143 (
		_w27256_,
		_w27318_,
		_w27656_
	);
	LUT2 #(
		.INIT('h4)
	) name17144 (
		_w27256_,
		_w27321_,
		_w27657_
	);
	LUT2 #(
		.INIT('h4)
	) name17145 (
		_w27256_,
		_w27326_,
		_w27658_
	);
	LUT2 #(
		.INIT('h4)
	) name17146 (
		_w27256_,
		_w27329_,
		_w27659_
	);
	LUT2 #(
		.INIT('h4)
	) name17147 (
		_w27256_,
		_w27331_,
		_w27660_
	);
	LUT2 #(
		.INIT('h4)
	) name17148 (
		_w27256_,
		_w27334_,
		_w27661_
	);
	LUT2 #(
		.INIT('h4)
	) name17149 (
		_w27256_,
		_w27337_,
		_w27662_
	);
	LUT2 #(
		.INIT('h4)
	) name17150 (
		_w27256_,
		_w27339_,
		_w27663_
	);
	LUT2 #(
		.INIT('h4)
	) name17151 (
		_w27256_,
		_w27342_,
		_w27664_
	);
	LUT2 #(
		.INIT('h4)
	) name17152 (
		_w27256_,
		_w27344_,
		_w27665_
	);
	LUT2 #(
		.INIT('h4)
	) name17153 (
		_w27256_,
		_w27347_,
		_w27666_
	);
	LUT2 #(
		.INIT('h4)
	) name17154 (
		_w27256_,
		_w27349_,
		_w27667_
	);
	LUT2 #(
		.INIT('h4)
	) name17155 (
		_w27256_,
		_w27352_,
		_w27668_
	);
	LUT2 #(
		.INIT('h4)
	) name17156 (
		_w27256_,
		_w27354_,
		_w27669_
	);
	LUT2 #(
		.INIT('h4)
	) name17157 (
		_w27256_,
		_w27356_,
		_w27670_
	);
	LUT2 #(
		.INIT('h4)
	) name17158 (
		_w27256_,
		_w27358_,
		_w27671_
	);
	LUT2 #(
		.INIT('h4)
	) name17159 (
		_w27256_,
		_w27360_,
		_w27672_
	);
	LUT2 #(
		.INIT('h4)
	) name17160 (
		_w27256_,
		_w27362_,
		_w27673_
	);
	LUT2 #(
		.INIT('h4)
	) name17161 (
		_w27256_,
		_w27364_,
		_w27674_
	);
	LUT2 #(
		.INIT('h4)
	) name17162 (
		_w27256_,
		_w27366_,
		_w27675_
	);
	LUT2 #(
		.INIT('h4)
	) name17163 (
		_w27256_,
		_w27368_,
		_w27676_
	);
	LUT2 #(
		.INIT('h4)
	) name17164 (
		_w27256_,
		_w27370_,
		_w27677_
	);
	LUT2 #(
		.INIT('h4)
	) name17165 (
		_w27256_,
		_w27372_,
		_w27678_
	);
	LUT2 #(
		.INIT('h4)
	) name17166 (
		_w27256_,
		_w27374_,
		_w27679_
	);
	LUT2 #(
		.INIT('h4)
	) name17167 (
		_w27256_,
		_w27376_,
		_w27680_
	);
	LUT2 #(
		.INIT('h4)
	) name17168 (
		_w27256_,
		_w27378_,
		_w27681_
	);
	LUT2 #(
		.INIT('h4)
	) name17169 (
		_w27256_,
		_w27380_,
		_w27682_
	);
	LUT2 #(
		.INIT('h4)
	) name17170 (
		_w27256_,
		_w27382_,
		_w27683_
	);
	LUT2 #(
		.INIT('h4)
	) name17171 (
		_w27256_,
		_w27384_,
		_w27684_
	);
	LUT2 #(
		.INIT('h4)
	) name17172 (
		_w27256_,
		_w27386_,
		_w27685_
	);
	LUT2 #(
		.INIT('h4)
	) name17173 (
		_w27256_,
		_w27388_,
		_w27686_
	);
	LUT2 #(
		.INIT('h4)
	) name17174 (
		_w27256_,
		_w27390_,
		_w27687_
	);
	LUT2 #(
		.INIT('h4)
	) name17175 (
		_w27256_,
		_w27393_,
		_w27688_
	);
	LUT2 #(
		.INIT('h4)
	) name17176 (
		_w27256_,
		_w27395_,
		_w27689_
	);
	LUT2 #(
		.INIT('h4)
	) name17177 (
		_w27256_,
		_w27398_,
		_w27690_
	);
	LUT2 #(
		.INIT('h4)
	) name17178 (
		_w27256_,
		_w27401_,
		_w27691_
	);
	LUT2 #(
		.INIT('h4)
	) name17179 (
		_w27256_,
		_w27403_,
		_w27692_
	);
	LUT2 #(
		.INIT('h4)
	) name17180 (
		_w27256_,
		_w27407_,
		_w27693_
	);
	LUT2 #(
		.INIT('h4)
	) name17181 (
		_w27256_,
		_w27410_,
		_w27694_
	);
	LUT2 #(
		.INIT('h4)
	) name17182 (
		_w27256_,
		_w27418_,
		_w27695_
	);
	LUT2 #(
		.INIT('h4)
	) name17183 (
		_w27256_,
		_w27421_,
		_w27696_
	);
	LUT2 #(
		.INIT('h4)
	) name17184 (
		_w27256_,
		_w27423_,
		_w27697_
	);
	LUT2 #(
		.INIT('h4)
	) name17185 (
		_w27256_,
		_w27425_,
		_w27698_
	);
	LUT2 #(
		.INIT('h4)
	) name17186 (
		_w27256_,
		_w27429_,
		_w27699_
	);
	LUT2 #(
		.INIT('h4)
	) name17187 (
		_w27256_,
		_w27431_,
		_w27700_
	);
	LUT2 #(
		.INIT('h4)
	) name17188 (
		_w27256_,
		_w27433_,
		_w27701_
	);
	LUT2 #(
		.INIT('h4)
	) name17189 (
		_w27256_,
		_w27435_,
		_w27702_
	);
	LUT2 #(
		.INIT('h4)
	) name17190 (
		_w27256_,
		_w27437_,
		_w27703_
	);
	LUT2 #(
		.INIT('h4)
	) name17191 (
		_w27256_,
		_w27439_,
		_w27704_
	);
	LUT2 #(
		.INIT('h4)
	) name17192 (
		_w27256_,
		_w27441_,
		_w27705_
	);
	LUT2 #(
		.INIT('h4)
	) name17193 (
		_w27256_,
		_w27443_,
		_w27706_
	);
	LUT2 #(
		.INIT('h4)
	) name17194 (
		_w27256_,
		_w27445_,
		_w27707_
	);
	LUT2 #(
		.INIT('h4)
	) name17195 (
		_w27256_,
		_w27447_,
		_w27708_
	);
	LUT2 #(
		.INIT('h4)
	) name17196 (
		_w27256_,
		_w27449_,
		_w27709_
	);
	LUT2 #(
		.INIT('h4)
	) name17197 (
		_w27256_,
		_w27453_,
		_w27710_
	);
	LUT2 #(
		.INIT('h4)
	) name17198 (
		_w27256_,
		_w27456_,
		_w27711_
	);
	LUT2 #(
		.INIT('h4)
	) name17199 (
		_w27256_,
		_w27458_,
		_w27712_
	);
	LUT2 #(
		.INIT('h4)
	) name17200 (
		_w27256_,
		_w27414_,
		_w27713_
	);
	LUT2 #(
		.INIT('h4)
	) name17201 (
		_w27256_,
		_w27461_,
		_w27714_
	);
	LUT2 #(
		.INIT('h4)
	) name17202 (
		_w27256_,
		_w27465_,
		_w27715_
	);
	LUT2 #(
		.INIT('h4)
	) name17203 (
		_w27256_,
		_w27467_,
		_w27716_
	);
	LUT2 #(
		.INIT('h4)
	) name17204 (
		_w27256_,
		_w27469_,
		_w27717_
	);
	LUT2 #(
		.INIT('h4)
	) name17205 (
		_w27256_,
		_w27471_,
		_w27718_
	);
	LUT2 #(
		.INIT('h4)
	) name17206 (
		_w27256_,
		_w27473_,
		_w27719_
	);
	LUT2 #(
		.INIT('h4)
	) name17207 (
		_w27256_,
		_w27475_,
		_w27720_
	);
	LUT2 #(
		.INIT('h4)
	) name17208 (
		_w27256_,
		_w27478_,
		_w27721_
	);
	LUT2 #(
		.INIT('h4)
	) name17209 (
		_w27256_,
		_w27283_,
		_w27722_
	);
	LUT2 #(
		.INIT('h4)
	) name17210 (
		_w27256_,
		_w27481_,
		_w27723_
	);
	LUT2 #(
		.INIT('h4)
	) name17211 (
		_w27256_,
		_w27484_,
		_w27724_
	);
	LUT2 #(
		.INIT('h8)
	) name17212 (
		_w27306_,
		_w27417_,
		_w27725_
	);
	LUT2 #(
		.INIT('h4)
	) name17213 (
		_w27256_,
		_w27725_,
		_w27726_
	);
	LUT2 #(
		.INIT('h8)
	) name17214 (
		_w27258_,
		_w27285_,
		_w27727_
	);
	LUT2 #(
		.INIT('h4)
	) name17215 (
		_w27256_,
		_w27727_,
		_w27728_
	);
	LUT2 #(
		.INIT('h8)
	) name17216 (
		_w27299_,
		_w27417_,
		_w27729_
	);
	LUT2 #(
		.INIT('h4)
	) name17217 (
		_w27262_,
		_w27729_,
		_w27730_
	);
	LUT2 #(
		.INIT('h8)
	) name17218 (
		_w27263_,
		_w27267_,
		_w27731_
	);
	LUT2 #(
		.INIT('h4)
	) name17219 (
		_w27262_,
		_w27731_,
		_w27732_
	);
	LUT2 #(
		.INIT('h8)
	) name17220 (
		_w27257_,
		_w27266_,
		_w27733_
	);
	LUT2 #(
		.INIT('h4)
	) name17221 (
		_w27262_,
		_w27733_,
		_w27734_
	);
	LUT2 #(
		.INIT('h8)
	) name17222 (
		_w27271_,
		_w27274_,
		_w27735_
	);
	LUT2 #(
		.INIT('h4)
	) name17223 (
		_w27262_,
		_w27735_,
		_w27736_
	);
	LUT2 #(
		.INIT('h8)
	) name17224 (
		_w27258_,
		_w27270_,
		_w27737_
	);
	LUT2 #(
		.INIT('h4)
	) name17225 (
		_w27262_,
		_w27737_,
		_w27738_
	);
	LUT2 #(
		.INIT('h8)
	) name17226 (
		_w27263_,
		_w27270_,
		_w27739_
	);
	LUT2 #(
		.INIT('h4)
	) name17227 (
		_w27262_,
		_w27739_,
		_w27740_
	);
	LUT2 #(
		.INIT('h8)
	) name17228 (
		_w27281_,
		_w27312_,
		_w27741_
	);
	LUT2 #(
		.INIT('h4)
	) name17229 (
		_w27262_,
		_w27741_,
		_w27742_
	);
	LUT2 #(
		.INIT('h8)
	) name17230 (
		_w27266_,
		_w27274_,
		_w27743_
	);
	LUT2 #(
		.INIT('h4)
	) name17231 (
		_w27262_,
		_w27743_,
		_w27744_
	);
	LUT2 #(
		.INIT('h8)
	) name17232 (
		_w27266_,
		_w27270_,
		_w27745_
	);
	LUT2 #(
		.INIT('h4)
	) name17233 (
		_w27262_,
		_w27745_,
		_w27746_
	);
	LUT2 #(
		.INIT('h8)
	) name17234 (
		_w27271_,
		_w27288_,
		_w27747_
	);
	LUT2 #(
		.INIT('h4)
	) name17235 (
		_w27262_,
		_w27747_,
		_w27748_
	);
	LUT2 #(
		.INIT('h4)
	) name17236 (
		_w27262_,
		_w27727_,
		_w27749_
	);
	LUT2 #(
		.INIT('h8)
	) name17237 (
		_w27263_,
		_w27285_,
		_w27750_
	);
	LUT2 #(
		.INIT('h4)
	) name17238 (
		_w27262_,
		_w27750_,
		_w27751_
	);
	LUT2 #(
		.INIT('h8)
	) name17239 (
		_w27266_,
		_w27288_,
		_w27752_
	);
	LUT2 #(
		.INIT('h4)
	) name17240 (
		_w27262_,
		_w27752_,
		_w27753_
	);
	LUT2 #(
		.INIT('h8)
	) name17241 (
		_w27263_,
		_w27312_,
		_w27754_
	);
	LUT2 #(
		.INIT('h4)
	) name17242 (
		_w27280_,
		_w27754_,
		_w27755_
	);
	LUT2 #(
		.INIT('h8)
	) name17243 (
		_w27266_,
		_w27285_,
		_w27756_
	);
	LUT2 #(
		.INIT('h4)
	) name17244 (
		_w27262_,
		_w27756_,
		_w27757_
	);
	LUT2 #(
		.INIT('h8)
	) name17245 (
		_w27281_,
		_w27306_,
		_w27758_
	);
	LUT2 #(
		.INIT('h4)
	) name17246 (
		_w27262_,
		_w27758_,
		_w27759_
	);
	LUT2 #(
		.INIT('h8)
	) name17247 (
		_w27258_,
		_w27293_,
		_w27760_
	);
	LUT2 #(
		.INIT('h4)
	) name17248 (
		_w27262_,
		_w27760_,
		_w27761_
	);
	LUT2 #(
		.INIT('h8)
	) name17249 (
		_w27258_,
		_w27282_,
		_w27762_
	);
	LUT2 #(
		.INIT('h4)
	) name17250 (
		_w27262_,
		_w27762_,
		_w27763_
	);
	LUT2 #(
		.INIT('h8)
	) name17251 (
		_w27263_,
		_w27293_,
		_w27764_
	);
	LUT2 #(
		.INIT('h4)
	) name17252 (
		_w27262_,
		_w27764_,
		_w27765_
	);
	LUT2 #(
		.INIT('h8)
	) name17253 (
		_w27263_,
		_w27282_,
		_w27766_
	);
	LUT2 #(
		.INIT('h4)
	) name17254 (
		_w27262_,
		_w27766_,
		_w27767_
	);
	LUT2 #(
		.INIT('h8)
	) name17255 (
		_w27266_,
		_w27293_,
		_w27768_
	);
	LUT2 #(
		.INIT('h4)
	) name17256 (
		_w27262_,
		_w27768_,
		_w27769_
	);
	LUT2 #(
		.INIT('h8)
	) name17257 (
		_w27266_,
		_w27282_,
		_w27770_
	);
	LUT2 #(
		.INIT('h4)
	) name17258 (
		_w27262_,
		_w27770_,
		_w27771_
	);
	LUT2 #(
		.INIT('h8)
	) name17259 (
		_w27299_,
		_w27324_,
		_w27772_
	);
	LUT2 #(
		.INIT('h4)
	) name17260 (
		_w27262_,
		_w27772_,
		_w27773_
	);
	LUT2 #(
		.INIT('h8)
	) name17261 (
		_w27302_,
		_w27324_,
		_w27774_
	);
	LUT2 #(
		.INIT('h4)
	) name17262 (
		_w27262_,
		_w27774_,
		_w27775_
	);
	LUT2 #(
		.INIT('h8)
	) name17263 (
		_w27312_,
		_w27413_,
		_w27776_
	);
	LUT2 #(
		.INIT('h4)
	) name17264 (
		_w27262_,
		_w27776_,
		_w27777_
	);
	LUT2 #(
		.INIT('h8)
	) name17265 (
		_w27299_,
		_w27305_,
		_w27778_
	);
	LUT2 #(
		.INIT('h4)
	) name17266 (
		_w27262_,
		_w27778_,
		_w27779_
	);
	LUT2 #(
		.INIT('h8)
	) name17267 (
		_w27302_,
		_w27305_,
		_w27780_
	);
	LUT2 #(
		.INIT('h4)
	) name17268 (
		_w27262_,
		_w27780_,
		_w27781_
	);
	LUT2 #(
		.INIT('h8)
	) name17269 (
		_w27299_,
		_w27309_,
		_w27782_
	);
	LUT2 #(
		.INIT('h4)
	) name17270 (
		_w27262_,
		_w27782_,
		_w27783_
	);
	LUT2 #(
		.INIT('h8)
	) name17271 (
		_w27302_,
		_w27309_,
		_w27784_
	);
	LUT2 #(
		.INIT('h4)
	) name17272 (
		_w27262_,
		_w27784_,
		_w27785_
	);
	LUT2 #(
		.INIT('h8)
	) name17273 (
		_w27312_,
		_w27324_,
		_w27786_
	);
	LUT2 #(
		.INIT('h4)
	) name17274 (
		_w27262_,
		_w27786_,
		_w27787_
	);
	LUT2 #(
		.INIT('h8)
	) name17275 (
		_w27306_,
		_w27324_,
		_w27788_
	);
	LUT2 #(
		.INIT('h4)
	) name17276 (
		_w27262_,
		_w27788_,
		_w27789_
	);
	LUT2 #(
		.INIT('h8)
	) name17277 (
		_w27305_,
		_w27312_,
		_w27790_
	);
	LUT2 #(
		.INIT('h4)
	) name17278 (
		_w27262_,
		_w27790_,
		_w27791_
	);
	LUT2 #(
		.INIT('h8)
	) name17279 (
		_w27306_,
		_w27413_,
		_w27792_
	);
	LUT2 #(
		.INIT('h4)
	) name17280 (
		_w27262_,
		_w27792_,
		_w27793_
	);
	LUT2 #(
		.INIT('h8)
	) name17281 (
		_w27309_,
		_w27312_,
		_w27794_
	);
	LUT2 #(
		.INIT('h4)
	) name17282 (
		_w27262_,
		_w27794_,
		_w27795_
	);
	LUT2 #(
		.INIT('h8)
	) name17283 (
		_w27298_,
		_w27306_,
		_w27796_
	);
	LUT2 #(
		.INIT('h4)
	) name17284 (
		_w27262_,
		_w27796_,
		_w27797_
	);
	LUT2 #(
		.INIT('h8)
	) name17285 (
		_w27320_,
		_w27324_,
		_w27798_
	);
	LUT2 #(
		.INIT('h4)
	) name17286 (
		_w27262_,
		_w27798_,
		_w27799_
	);
	LUT2 #(
		.INIT('h4)
	) name17287 (
		_w27256_,
		_w27774_,
		_w27800_
	);
	LUT2 #(
		.INIT('h4)
	) name17288 (
		_w27256_,
		_w27784_,
		_w27801_
	);
	LUT2 #(
		.INIT('h8)
	) name17289 (
		_w27315_,
		_w27324_,
		_w27802_
	);
	LUT2 #(
		.INIT('h4)
	) name17290 (
		_w27262_,
		_w27802_,
		_w27803_
	);
	LUT2 #(
		.INIT('h8)
	) name17291 (
		_w27305_,
		_w27320_,
		_w27804_
	);
	LUT2 #(
		.INIT('h4)
	) name17292 (
		_w27262_,
		_w27804_,
		_w27805_
	);
	LUT2 #(
		.INIT('h4)
	) name17293 (
		_w27256_,
		_w27770_,
		_w27806_
	);
	LUT2 #(
		.INIT('h8)
	) name17294 (
		_w27309_,
		_w27320_,
		_w27807_
	);
	LUT2 #(
		.INIT('h4)
	) name17295 (
		_w27262_,
		_w27807_,
		_w27808_
	);
	LUT2 #(
		.INIT('h8)
	) name17296 (
		_w27312_,
		_w27333_,
		_w27809_
	);
	LUT2 #(
		.INIT('h4)
	) name17297 (
		_w27262_,
		_w27809_,
		_w27810_
	);
	LUT2 #(
		.INIT('h4)
	) name17298 (
		_w27256_,
		_w27786_,
		_w27811_
	);
	LUT2 #(
		.INIT('h8)
	) name17299 (
		_w27298_,
		_w27315_,
		_w27812_
	);
	LUT2 #(
		.INIT('h4)
	) name17300 (
		_w27262_,
		_w27812_,
		_w27813_
	);
	LUT2 #(
		.INIT('h8)
	) name17301 (
		_w27324_,
		_w27328_,
		_w27814_
	);
	LUT2 #(
		.INIT('h4)
	) name17302 (
		_w27262_,
		_w27814_,
		_w27815_
	);
	LUT2 #(
		.INIT('h8)
	) name17303 (
		_w27305_,
		_w27325_,
		_w27816_
	);
	LUT2 #(
		.INIT('h4)
	) name17304 (
		_w27262_,
		_w27816_,
		_w27817_
	);
	LUT2 #(
		.INIT('h8)
	) name17305 (
		_w27309_,
		_w27325_,
		_w27818_
	);
	LUT2 #(
		.INIT('h4)
	) name17306 (
		_w27262_,
		_w27818_,
		_w27819_
	);
	LUT2 #(
		.INIT('h8)
	) name17307 (
		_w27298_,
		_w27328_,
		_w27820_
	);
	LUT2 #(
		.INIT('h4)
	) name17308 (
		_w27262_,
		_w27820_,
		_w27821_
	);
	LUT2 #(
		.INIT('h4)
	) name17309 (
		_w27256_,
		_w27778_,
		_w27822_
	);
	LUT2 #(
		.INIT('h8)
	) name17310 (
		_w27298_,
		_w27325_,
		_w27823_
	);
	LUT2 #(
		.INIT('h4)
	) name17311 (
		_w27262_,
		_w27823_,
		_w27824_
	);
	LUT2 #(
		.INIT('h8)
	) name17312 (
		_w27299_,
		_w27351_,
		_w27825_
	);
	LUT2 #(
		.INIT('h4)
	) name17313 (
		_w27262_,
		_w27825_,
		_w27826_
	);
	LUT2 #(
		.INIT('h8)
	) name17314 (
		_w27302_,
		_w27351_,
		_w27827_
	);
	LUT2 #(
		.INIT('h4)
	) name17315 (
		_w27262_,
		_w27827_,
		_w27828_
	);
	LUT2 #(
		.INIT('h4)
	) name17316 (
		_w27256_,
		_w27776_,
		_w27829_
	);
	LUT2 #(
		.INIT('h4)
	) name17317 (
		_w27256_,
		_w27792_,
		_w27830_
	);
	LUT2 #(
		.INIT('h8)
	) name17318 (
		_w27312_,
		_w27351_,
		_w27831_
	);
	LUT2 #(
		.INIT('h4)
	) name17319 (
		_w27262_,
		_w27831_,
		_w27832_
	);
	LUT2 #(
		.INIT('h8)
	) name17320 (
		_w27320_,
		_w27417_,
		_w27833_
	);
	LUT2 #(
		.INIT('h4)
	) name17321 (
		_w27262_,
		_w27833_,
		_w27834_
	);
	LUT2 #(
		.INIT('h8)
	) name17322 (
		_w27306_,
		_w27336_,
		_w27835_
	);
	LUT2 #(
		.INIT('h4)
	) name17323 (
		_w27262_,
		_w27835_,
		_w27836_
	);
	LUT2 #(
		.INIT('h8)
	) name17324 (
		_w27306_,
		_w27341_,
		_w27837_
	);
	LUT2 #(
		.INIT('h4)
	) name17325 (
		_w27262_,
		_w27837_,
		_w27838_
	);
	LUT2 #(
		.INIT('h4)
	) name17326 (
		_w27256_,
		_w27790_,
		_w27839_
	);
	LUT2 #(
		.INIT('h8)
	) name17327 (
		_w27306_,
		_w27346_,
		_w27840_
	);
	LUT2 #(
		.INIT('h4)
	) name17328 (
		_w27262_,
		_w27840_,
		_w27841_
	);
	LUT2 #(
		.INIT('h8)
	) name17329 (
		_w27320_,
		_w27351_,
		_w27842_
	);
	LUT2 #(
		.INIT('h4)
	) name17330 (
		_w27262_,
		_w27842_,
		_w27843_
	);
	LUT2 #(
		.INIT('h4)
	) name17331 (
		_w27256_,
		_w27782_,
		_w27844_
	);
	LUT2 #(
		.INIT('h8)
	) name17332 (
		_w27315_,
		_w27336_,
		_w27845_
	);
	LUT2 #(
		.INIT('h4)
	) name17333 (
		_w27262_,
		_w27845_,
		_w27846_
	);
	LUT2 #(
		.INIT('h8)
	) name17334 (
		_w27315_,
		_w27417_,
		_w27847_
	);
	LUT2 #(
		.INIT('h4)
	) name17335 (
		_w27262_,
		_w27847_,
		_w27848_
	);
	LUT2 #(
		.INIT('h4)
	) name17336 (
		_w27256_,
		_w27768_,
		_w27849_
	);
	LUT2 #(
		.INIT('h8)
	) name17337 (
		_w27267_,
		_w27417_,
		_w27850_
	);
	LUT2 #(
		.INIT('h4)
	) name17338 (
		_w27280_,
		_w27850_,
		_w27851_
	);
	LUT2 #(
		.INIT('h8)
	) name17339 (
		_w27315_,
		_w27341_,
		_w27852_
	);
	LUT2 #(
		.INIT('h4)
	) name17340 (
		_w27262_,
		_w27852_,
		_w27853_
	);
	LUT2 #(
		.INIT('h8)
	) name17341 (
		_w27315_,
		_w27346_,
		_w27854_
	);
	LUT2 #(
		.INIT('h4)
	) name17342 (
		_w27262_,
		_w27854_,
		_w27855_
	);
	LUT2 #(
		.INIT('h8)
	) name17343 (
		_w27325_,
		_w27351_,
		_w27856_
	);
	LUT2 #(
		.INIT('h4)
	) name17344 (
		_w27262_,
		_w27856_,
		_w27857_
	);
	LUT2 #(
		.INIT('h8)
	) name17345 (
		_w27328_,
		_w27336_,
		_w27858_
	);
	LUT2 #(
		.INIT('h4)
	) name17346 (
		_w27262_,
		_w27858_,
		_w27859_
	);
	LUT2 #(
		.INIT('h8)
	) name17347 (
		_w27325_,
		_w27336_,
		_w27860_
	);
	LUT2 #(
		.INIT('h4)
	) name17348 (
		_w27262_,
		_w27860_,
		_w27861_
	);
	LUT2 #(
		.INIT('h8)
	) name17349 (
		_w27328_,
		_w27341_,
		_w27862_
	);
	LUT2 #(
		.INIT('h4)
	) name17350 (
		_w27262_,
		_w27862_,
		_w27863_
	);
	LUT2 #(
		.INIT('h8)
	) name17351 (
		_w27325_,
		_w27341_,
		_w27864_
	);
	LUT2 #(
		.INIT('h4)
	) name17352 (
		_w27262_,
		_w27864_,
		_w27865_
	);
	LUT2 #(
		.INIT('h4)
	) name17353 (
		_w27256_,
		_w27731_,
		_w27866_
	);
	LUT2 #(
		.INIT('h8)
	) name17354 (
		_w27281_,
		_w27320_,
		_w27867_
	);
	LUT2 #(
		.INIT('h4)
	) name17355 (
		_w27262_,
		_w27867_,
		_w27868_
	);
	LUT2 #(
		.INIT('h8)
	) name17356 (
		_w27328_,
		_w27346_,
		_w27869_
	);
	LUT2 #(
		.INIT('h4)
	) name17357 (
		_w27262_,
		_w27869_,
		_w27870_
	);
	LUT2 #(
		.INIT('h8)
	) name17358 (
		_w27325_,
		_w27346_,
		_w27871_
	);
	LUT2 #(
		.INIT('h4)
	) name17359 (
		_w27262_,
		_w27871_,
		_w27872_
	);
	LUT2 #(
		.INIT('h8)
	) name17360 (
		_w27267_,
		_w27324_,
		_w27873_
	);
	LUT2 #(
		.INIT('h4)
	) name17361 (
		_w27262_,
		_w27873_,
		_w27874_
	);
	LUT2 #(
		.INIT('h8)
	) name17362 (
		_w27257_,
		_w27324_,
		_w27875_
	);
	LUT2 #(
		.INIT('h4)
	) name17363 (
		_w27262_,
		_w27875_,
		_w27876_
	);
	LUT2 #(
		.INIT('h8)
	) name17364 (
		_w27267_,
		_w27305_,
		_w27877_
	);
	LUT2 #(
		.INIT('h4)
	) name17365 (
		_w27262_,
		_w27877_,
		_w27878_
	);
	LUT2 #(
		.INIT('h8)
	) name17366 (
		_w27267_,
		_w27309_,
		_w27879_
	);
	LUT2 #(
		.INIT('h4)
	) name17367 (
		_w27262_,
		_w27879_,
		_w27880_
	);
	LUT2 #(
		.INIT('h8)
	) name17368 (
		_w27257_,
		_w27298_,
		_w27881_
	);
	LUT2 #(
		.INIT('h4)
	) name17369 (
		_w27262_,
		_w27881_,
		_w27882_
	);
	LUT2 #(
		.INIT('h8)
	) name17370 (
		_w27281_,
		_w27315_,
		_w27883_
	);
	LUT2 #(
		.INIT('h4)
	) name17371 (
		_w27262_,
		_w27883_,
		_w27884_
	);
	LUT2 #(
		.INIT('h8)
	) name17372 (
		_w27302_,
		_w27417_,
		_w27885_
	);
	LUT2 #(
		.INIT('h4)
	) name17373 (
		_w27262_,
		_w27885_,
		_w27886_
	);
	LUT2 #(
		.INIT('h8)
	) name17374 (
		_w27274_,
		_w27324_,
		_w27887_
	);
	LUT2 #(
		.INIT('h4)
	) name17375 (
		_w27262_,
		_w27887_,
		_w27888_
	);
	LUT2 #(
		.INIT('h4)
	) name17376 (
		_w27256_,
		_w27766_,
		_w27889_
	);
	LUT2 #(
		.INIT('h8)
	) name17377 (
		_w27270_,
		_w27305_,
		_w27890_
	);
	LUT2 #(
		.INIT('h4)
	) name17378 (
		_w27262_,
		_w27890_,
		_w27891_
	);
	LUT2 #(
		.INIT('h8)
	) name17379 (
		_w27270_,
		_w27309_,
		_w27892_
	);
	LUT2 #(
		.INIT('h4)
	) name17380 (
		_w27262_,
		_w27892_,
		_w27893_
	);
	LUT2 #(
		.INIT('h8)
	) name17381 (
		_w27274_,
		_w27298_,
		_w27894_
	);
	LUT2 #(
		.INIT('h4)
	) name17382 (
		_w27262_,
		_w27894_,
		_w27895_
	);
	LUT2 #(
		.INIT('h8)
	) name17383 (
		_w27270_,
		_w27298_,
		_w27896_
	);
	LUT2 #(
		.INIT('h4)
	) name17384 (
		_w27262_,
		_w27896_,
		_w27897_
	);
	LUT2 #(
		.INIT('h8)
	) name17385 (
		_w27288_,
		_w27324_,
		_w27898_
	);
	LUT2 #(
		.INIT('h4)
	) name17386 (
		_w27262_,
		_w27898_,
		_w27899_
	);
	LUT2 #(
		.INIT('h8)
	) name17387 (
		_w27320_,
		_w27413_,
		_w27900_
	);
	LUT2 #(
		.INIT('h4)
	) name17388 (
		_w27262_,
		_w27900_,
		_w27901_
	);
	LUT2 #(
		.INIT('h8)
	) name17389 (
		_w27285_,
		_w27305_,
		_w27902_
	);
	LUT2 #(
		.INIT('h4)
	) name17390 (
		_w27262_,
		_w27902_,
		_w27903_
	);
	LUT2 #(
		.INIT('h8)
	) name17391 (
		_w27285_,
		_w27309_,
		_w27904_
	);
	LUT2 #(
		.INIT('h4)
	) name17392 (
		_w27262_,
		_w27904_,
		_w27905_
	);
	LUT2 #(
		.INIT('h8)
	) name17393 (
		_w27288_,
		_w27298_,
		_w27906_
	);
	LUT2 #(
		.INIT('h4)
	) name17394 (
		_w27262_,
		_w27906_,
		_w27907_
	);
	LUT2 #(
		.INIT('h8)
	) name17395 (
		_w27285_,
		_w27298_,
		_w27908_
	);
	LUT2 #(
		.INIT('h4)
	) name17396 (
		_w27262_,
		_w27908_,
		_w27909_
	);
	LUT2 #(
		.INIT('h8)
	) name17397 (
		_w27281_,
		_w27288_,
		_w27910_
	);
	LUT2 #(
		.INIT('h4)
	) name17398 (
		_w27280_,
		_w27910_,
		_w27911_
	);
	LUT2 #(
		.INIT('h8)
	) name17399 (
		_w27293_,
		_w27305_,
		_w27912_
	);
	LUT2 #(
		.INIT('h4)
	) name17400 (
		_w27262_,
		_w27912_,
		_w27913_
	);
	LUT2 #(
		.INIT('h8)
	) name17401 (
		_w27282_,
		_w27305_,
		_w27914_
	);
	LUT2 #(
		.INIT('h4)
	) name17402 (
		_w27262_,
		_w27914_,
		_w27915_
	);
	LUT2 #(
		.INIT('h8)
	) name17403 (
		_w27315_,
		_w27413_,
		_w27916_
	);
	LUT2 #(
		.INIT('h4)
	) name17404 (
		_w27262_,
		_w27916_,
		_w27917_
	);
	LUT2 #(
		.INIT('h8)
	) name17405 (
		_w27293_,
		_w27309_,
		_w27918_
	);
	LUT2 #(
		.INIT('h4)
	) name17406 (
		_w27262_,
		_w27918_,
		_w27919_
	);
	LUT2 #(
		.INIT('h8)
	) name17407 (
		_w27282_,
		_w27309_,
		_w27920_
	);
	LUT2 #(
		.INIT('h4)
	) name17408 (
		_w27262_,
		_w27920_,
		_w27921_
	);
	LUT2 #(
		.INIT('h4)
	) name17409 (
		_w27280_,
		_w27729_,
		_w27922_
	);
	LUT2 #(
		.INIT('h8)
	) name17410 (
		_w27293_,
		_w27298_,
		_w27923_
	);
	LUT2 #(
		.INIT('h4)
	) name17411 (
		_w27262_,
		_w27923_,
		_w27924_
	);
	LUT2 #(
		.INIT('h8)
	) name17412 (
		_w27282_,
		_w27298_,
		_w27925_
	);
	LUT2 #(
		.INIT('h4)
	) name17413 (
		_w27262_,
		_w27925_,
		_w27926_
	);
	LUT2 #(
		.INIT('h8)
	) name17414 (
		_w27267_,
		_w27351_,
		_w27927_
	);
	LUT2 #(
		.INIT('h4)
	) name17415 (
		_w27262_,
		_w27927_,
		_w27928_
	);
	LUT2 #(
		.INIT('h4)
	) name17416 (
		_w27280_,
		_w27731_,
		_w27929_
	);
	LUT2 #(
		.INIT('h8)
	) name17417 (
		_w27257_,
		_w27336_,
		_w27930_
	);
	LUT2 #(
		.INIT('h4)
	) name17418 (
		_w27262_,
		_w27930_,
		_w27931_
	);
	LUT2 #(
		.INIT('h8)
	) name17419 (
		_w27257_,
		_w27341_,
		_w27932_
	);
	LUT2 #(
		.INIT('h4)
	) name17420 (
		_w27262_,
		_w27932_,
		_w27933_
	);
	LUT2 #(
		.INIT('h8)
	) name17421 (
		_w27320_,
		_w27333_,
		_w27934_
	);
	LUT2 #(
		.INIT('h4)
	) name17422 (
		_w27262_,
		_w27934_,
		_w27935_
	);
	LUT2 #(
		.INIT('h4)
	) name17423 (
		_w27280_,
		_w27733_,
		_w27936_
	);
	LUT2 #(
		.INIT('h8)
	) name17424 (
		_w27257_,
		_w27346_,
		_w27937_
	);
	LUT2 #(
		.INIT('h4)
	) name17425 (
		_w27262_,
		_w27937_,
		_w27938_
	);
	LUT2 #(
		.INIT('h4)
	) name17426 (
		_w27280_,
		_w27735_,
		_w27939_
	);
	LUT2 #(
		.INIT('h8)
	) name17427 (
		_w27270_,
		_w27351_,
		_w27940_
	);
	LUT2 #(
		.INIT('h4)
	) name17428 (
		_w27262_,
		_w27940_,
		_w27941_
	);
	LUT2 #(
		.INIT('h8)
	) name17429 (
		_w27274_,
		_w27336_,
		_w27942_
	);
	LUT2 #(
		.INIT('h4)
	) name17430 (
		_w27262_,
		_w27942_,
		_w27943_
	);
	LUT2 #(
		.INIT('h8)
	) name17431 (
		_w27270_,
		_w27336_,
		_w27944_
	);
	LUT2 #(
		.INIT('h4)
	) name17432 (
		_w27262_,
		_w27944_,
		_w27945_
	);
	LUT2 #(
		.INIT('h8)
	) name17433 (
		_w27274_,
		_w27341_,
		_w27946_
	);
	LUT2 #(
		.INIT('h4)
	) name17434 (
		_w27262_,
		_w27946_,
		_w27947_
	);
	LUT2 #(
		.INIT('h8)
	) name17435 (
		_w27270_,
		_w27341_,
		_w27948_
	);
	LUT2 #(
		.INIT('h4)
	) name17436 (
		_w27262_,
		_w27948_,
		_w27949_
	);
	LUT2 #(
		.INIT('h8)
	) name17437 (
		_w27274_,
		_w27346_,
		_w27950_
	);
	LUT2 #(
		.INIT('h4)
	) name17438 (
		_w27262_,
		_w27950_,
		_w27951_
	);
	LUT2 #(
		.INIT('h4)
	) name17439 (
		_w27280_,
		_w27737_,
		_w27952_
	);
	LUT2 #(
		.INIT('h8)
	) name17440 (
		_w27270_,
		_w27346_,
		_w27953_
	);
	LUT2 #(
		.INIT('h4)
	) name17441 (
		_w27262_,
		_w27953_,
		_w27954_
	);
	LUT2 #(
		.INIT('h8)
	) name17442 (
		_w27302_,
		_w27333_,
		_w27955_
	);
	LUT2 #(
		.INIT('h4)
	) name17443 (
		_w27280_,
		_w27955_,
		_w27956_
	);
	LUT2 #(
		.INIT('h8)
	) name17444 (
		_w27285_,
		_w27351_,
		_w27957_
	);
	LUT2 #(
		.INIT('h4)
	) name17445 (
		_w27262_,
		_w27957_,
		_w27958_
	);
	LUT2 #(
		.INIT('h4)
	) name17446 (
		_w27280_,
		_w27739_,
		_w27959_
	);
	LUT2 #(
		.INIT('h8)
	) name17447 (
		_w27288_,
		_w27336_,
		_w27960_
	);
	LUT2 #(
		.INIT('h4)
	) name17448 (
		_w27262_,
		_w27960_,
		_w27961_
	);
	LUT2 #(
		.INIT('h8)
	) name17449 (
		_w27285_,
		_w27336_,
		_w27962_
	);
	LUT2 #(
		.INIT('h4)
	) name17450 (
		_w27262_,
		_w27962_,
		_w27963_
	);
	LUT2 #(
		.INIT('h4)
	) name17451 (
		_w27280_,
		_w27741_,
		_w27964_
	);
	LUT2 #(
		.INIT('h8)
	) name17452 (
		_w27288_,
		_w27341_,
		_w27965_
	);
	LUT2 #(
		.INIT('h4)
	) name17453 (
		_w27262_,
		_w27965_,
		_w27966_
	);
	LUT2 #(
		.INIT('h8)
	) name17454 (
		_w27285_,
		_w27341_,
		_w27967_
	);
	LUT2 #(
		.INIT('h4)
	) name17455 (
		_w27262_,
		_w27967_,
		_w27968_
	);
	LUT2 #(
		.INIT('h4)
	) name17456 (
		_w27280_,
		_w27743_,
		_w27969_
	);
	LUT2 #(
		.INIT('h8)
	) name17457 (
		_w27288_,
		_w27346_,
		_w27970_
	);
	LUT2 #(
		.INIT('h4)
	) name17458 (
		_w27262_,
		_w27970_,
		_w27971_
	);
	LUT2 #(
		.INIT('h8)
	) name17459 (
		_w27285_,
		_w27346_,
		_w27972_
	);
	LUT2 #(
		.INIT('h4)
	) name17460 (
		_w27262_,
		_w27972_,
		_w27973_
	);
	LUT2 #(
		.INIT('h4)
	) name17461 (
		_w27280_,
		_w27745_,
		_w27974_
	);
	LUT2 #(
		.INIT('h8)
	) name17462 (
		_w27293_,
		_w27351_,
		_w27975_
	);
	LUT2 #(
		.INIT('h4)
	) name17463 (
		_w27262_,
		_w27975_,
		_w27976_
	);
	LUT2 #(
		.INIT('h8)
	) name17464 (
		_w27282_,
		_w27351_,
		_w27977_
	);
	LUT2 #(
		.INIT('h4)
	) name17465 (
		_w27262_,
		_w27977_,
		_w27978_
	);
	LUT2 #(
		.INIT('h4)
	) name17466 (
		_w27280_,
		_w27747_,
		_w27979_
	);
	LUT2 #(
		.INIT('h8)
	) name17467 (
		_w27328_,
		_w27417_,
		_w27980_
	);
	LUT2 #(
		.INIT('h4)
	) name17468 (
		_w27262_,
		_w27980_,
		_w27981_
	);
	LUT2 #(
		.INIT('h8)
	) name17469 (
		_w27293_,
		_w27336_,
		_w27982_
	);
	LUT2 #(
		.INIT('h4)
	) name17470 (
		_w27262_,
		_w27982_,
		_w27983_
	);
	LUT2 #(
		.INIT('h8)
	) name17471 (
		_w27282_,
		_w27336_,
		_w27984_
	);
	LUT2 #(
		.INIT('h4)
	) name17472 (
		_w27262_,
		_w27984_,
		_w27985_
	);
	LUT2 #(
		.INIT('h8)
	) name17473 (
		_w27293_,
		_w27341_,
		_w27986_
	);
	LUT2 #(
		.INIT('h4)
	) name17474 (
		_w27262_,
		_w27986_,
		_w27987_
	);
	LUT2 #(
		.INIT('h8)
	) name17475 (
		_w27282_,
		_w27341_,
		_w27988_
	);
	LUT2 #(
		.INIT('h4)
	) name17476 (
		_w27262_,
		_w27988_,
		_w27989_
	);
	LUT2 #(
		.INIT('h4)
	) name17477 (
		_w27256_,
		_w27764_,
		_w27990_
	);
	LUT2 #(
		.INIT('h8)
	) name17478 (
		_w27293_,
		_w27346_,
		_w27991_
	);
	LUT2 #(
		.INIT('h4)
	) name17479 (
		_w27262_,
		_w27991_,
		_w27992_
	);
	LUT2 #(
		.INIT('h4)
	) name17480 (
		_w27280_,
		_w27727_,
		_w27993_
	);
	LUT2 #(
		.INIT('h8)
	) name17481 (
		_w27282_,
		_w27346_,
		_w27994_
	);
	LUT2 #(
		.INIT('h4)
	) name17482 (
		_w27262_,
		_w27994_,
		_w27995_
	);
	LUT2 #(
		.INIT('h8)
	) name17483 (
		_w27281_,
		_w27328_,
		_w27996_
	);
	LUT2 #(
		.INIT('h4)
	) name17484 (
		_w27262_,
		_w27996_,
		_w27997_
	);
	LUT2 #(
		.INIT('h4)
	) name17485 (
		_w27280_,
		_w27750_,
		_w27998_
	);
	LUT2 #(
		.INIT('h8)
	) name17486 (
		_w27328_,
		_w27413_,
		_w27999_
	);
	LUT2 #(
		.INIT('h4)
	) name17487 (
		_w27262_,
		_w27999_,
		_w28000_
	);
	LUT2 #(
		.INIT('h8)
	) name17488 (
		_w27281_,
		_w27299_,
		_w28001_
	);
	LUT2 #(
		.INIT('h4)
	) name17489 (
		_w27262_,
		_w28001_,
		_w28002_
	);
	LUT2 #(
		.INIT('h4)
	) name17490 (
		_w27280_,
		_w27752_,
		_w28003_
	);
	LUT2 #(
		.INIT('h4)
	) name17491 (
		_w27280_,
		_w27756_,
		_w28004_
	);
	LUT2 #(
		.INIT('h8)
	) name17492 (
		_w27325_,
		_w27333_,
		_w28005_
	);
	LUT2 #(
		.INIT('h4)
	) name17493 (
		_w27262_,
		_w28005_,
		_w28006_
	);
	LUT2 #(
		.INIT('h8)
	) name17494 (
		_w27271_,
		_w27299_,
		_w28007_
	);
	LUT2 #(
		.INIT('h4)
	) name17495 (
		_w27262_,
		_w28007_,
		_w28008_
	);
	LUT2 #(
		.INIT('h4)
	) name17496 (
		_w27280_,
		_w27758_,
		_w28009_
	);
	LUT2 #(
		.INIT('h8)
	) name17497 (
		_w27271_,
		_w27302_,
		_w28010_
	);
	LUT2 #(
		.INIT('h4)
	) name17498 (
		_w27262_,
		_w28010_,
		_w28011_
	);
	LUT2 #(
		.INIT('h8)
	) name17499 (
		_w27258_,
		_w27299_,
		_w28012_
	);
	LUT2 #(
		.INIT('h4)
	) name17500 (
		_w27262_,
		_w28012_,
		_w28013_
	);
	LUT2 #(
		.INIT('h8)
	) name17501 (
		_w27258_,
		_w27302_,
		_w28014_
	);
	LUT2 #(
		.INIT('h4)
	) name17502 (
		_w27262_,
		_w28014_,
		_w28015_
	);
	LUT2 #(
		.INIT('h8)
	) name17503 (
		_w27263_,
		_w27299_,
		_w28016_
	);
	LUT2 #(
		.INIT('h4)
	) name17504 (
		_w27262_,
		_w28016_,
		_w28017_
	);
	LUT2 #(
		.INIT('h8)
	) name17505 (
		_w27263_,
		_w27302_,
		_w28018_
	);
	LUT2 #(
		.INIT('h4)
	) name17506 (
		_w27262_,
		_w28018_,
		_w28019_
	);
	LUT2 #(
		.INIT('h4)
	) name17507 (
		_w27280_,
		_w27760_,
		_w28020_
	);
	LUT2 #(
		.INIT('h8)
	) name17508 (
		_w27281_,
		_w27302_,
		_w28021_
	);
	LUT2 #(
		.INIT('h4)
	) name17509 (
		_w27262_,
		_w28021_,
		_w28022_
	);
	LUT2 #(
		.INIT('h8)
	) name17510 (
		_w27271_,
		_w27312_,
		_w28023_
	);
	LUT2 #(
		.INIT('h4)
	) name17511 (
		_w27262_,
		_w28023_,
		_w28024_
	);
	LUT2 #(
		.INIT('h4)
	) name17512 (
		_w27280_,
		_w27762_,
		_w28025_
	);
	LUT2 #(
		.INIT('h8)
	) name17513 (
		_w27271_,
		_w27306_,
		_w28026_
	);
	LUT2 #(
		.INIT('h4)
	) name17514 (
		_w27262_,
		_w28026_,
		_w28027_
	);
	LUT2 #(
		.INIT('h8)
	) name17515 (
		_w27258_,
		_w27312_,
		_w28028_
	);
	LUT2 #(
		.INIT('h4)
	) name17516 (
		_w27262_,
		_w28028_,
		_w28029_
	);
	LUT2 #(
		.INIT('h4)
	) name17517 (
		_w27280_,
		_w27764_,
		_w28030_
	);
	LUT2 #(
		.INIT('h4)
	) name17518 (
		_w27262_,
		_w27754_,
		_w28031_
	);
	LUT2 #(
		.INIT('h4)
	) name17519 (
		_w27280_,
		_w27766_,
		_w28032_
	);
	LUT2 #(
		.INIT('h4)
	) name17520 (
		_w27280_,
		_w27768_,
		_w28033_
	);
	LUT2 #(
		.INIT('h8)
	) name17521 (
		_w27266_,
		_w27306_,
		_w28034_
	);
	LUT2 #(
		.INIT('h4)
	) name17522 (
		_w27262_,
		_w28034_,
		_w28035_
	);
	LUT2 #(
		.INIT('h8)
	) name17523 (
		_w27271_,
		_w27320_,
		_w28036_
	);
	LUT2 #(
		.INIT('h4)
	) name17524 (
		_w27262_,
		_w28036_,
		_w28037_
	);
	LUT2 #(
		.INIT('h4)
	) name17525 (
		_w27280_,
		_w27770_,
		_w28038_
	);
	LUT2 #(
		.INIT('h8)
	) name17526 (
		_w27271_,
		_w27315_,
		_w28039_
	);
	LUT2 #(
		.INIT('h4)
	) name17527 (
		_w27262_,
		_w28039_,
		_w28040_
	);
	LUT2 #(
		.INIT('h8)
	) name17528 (
		_w27299_,
		_w27413_,
		_w28041_
	);
	LUT2 #(
		.INIT('h4)
	) name17529 (
		_w27262_,
		_w28041_,
		_w28042_
	);
	LUT2 #(
		.INIT('h4)
	) name17530 (
		_w27280_,
		_w27772_,
		_w28043_
	);
	LUT2 #(
		.INIT('h8)
	) name17531 (
		_w27258_,
		_w27320_,
		_w28044_
	);
	LUT2 #(
		.INIT('h4)
	) name17532 (
		_w27262_,
		_w28044_,
		_w28045_
	);
	LUT2 #(
		.INIT('h4)
	) name17533 (
		_w27280_,
		_w27774_,
		_w28046_
	);
	LUT2 #(
		.INIT('h8)
	) name17534 (
		_w27263_,
		_w27320_,
		_w28047_
	);
	LUT2 #(
		.INIT('h4)
	) name17535 (
		_w27262_,
		_w28047_,
		_w28048_
	);
	LUT2 #(
		.INIT('h4)
	) name17536 (
		_w27280_,
		_w27776_,
		_w28049_
	);
	LUT2 #(
		.INIT('h8)
	) name17537 (
		_w27266_,
		_w27315_,
		_w28050_
	);
	LUT2 #(
		.INIT('h4)
	) name17538 (
		_w27262_,
		_w28050_,
		_w28051_
	);
	LUT2 #(
		.INIT('h4)
	) name17539 (
		_w27280_,
		_w27778_,
		_w28052_
	);
	LUT2 #(
		.INIT('h8)
	) name17540 (
		_w27271_,
		_w27328_,
		_w28053_
	);
	LUT2 #(
		.INIT('h4)
	) name17541 (
		_w27262_,
		_w28053_,
		_w28054_
	);
	LUT2 #(
		.INIT('h4)
	) name17542 (
		_w27280_,
		_w27780_,
		_w28055_
	);
	LUT2 #(
		.INIT('h8)
	) name17543 (
		_w27258_,
		_w27325_,
		_w28056_
	);
	LUT2 #(
		.INIT('h4)
	) name17544 (
		_w27262_,
		_w28056_,
		_w28057_
	);
	LUT2 #(
		.INIT('h4)
	) name17545 (
		_w27280_,
		_w27782_,
		_w28058_
	);
	LUT2 #(
		.INIT('h8)
	) name17546 (
		_w27302_,
		_w27413_,
		_w28059_
	);
	LUT2 #(
		.INIT('h4)
	) name17547 (
		_w27262_,
		_w28059_,
		_w28060_
	);
	LUT2 #(
		.INIT('h4)
	) name17548 (
		_w27280_,
		_w27784_,
		_w28061_
	);
	LUT2 #(
		.INIT('h8)
	) name17549 (
		_w27263_,
		_w27325_,
		_w28062_
	);
	LUT2 #(
		.INIT('h4)
	) name17550 (
		_w27262_,
		_w28062_,
		_w28063_
	);
	LUT2 #(
		.INIT('h8)
	) name17551 (
		_w27266_,
		_w27328_,
		_w28064_
	);
	LUT2 #(
		.INIT('h4)
	) name17552 (
		_w27262_,
		_w28064_,
		_w28065_
	);
	LUT2 #(
		.INIT('h8)
	) name17553 (
		_w27266_,
		_w27325_,
		_w28066_
	);
	LUT2 #(
		.INIT('h4)
	) name17554 (
		_w27262_,
		_w28066_,
		_w28067_
	);
	LUT2 #(
		.INIT('h4)
	) name17555 (
		_w27262_,
		_w27850_,
		_w28068_
	);
	LUT2 #(
		.INIT('h8)
	) name17556 (
		_w27257_,
		_w27417_,
		_w28069_
	);
	LUT2 #(
		.INIT('h4)
	) name17557 (
		_w27262_,
		_w28069_,
		_w28070_
	);
	LUT2 #(
		.INIT('h4)
	) name17558 (
		_w27280_,
		_w28062_,
		_w28071_
	);
	LUT2 #(
		.INIT('h8)
	) name17559 (
		_w27267_,
		_w27281_,
		_w28072_
	);
	LUT2 #(
		.INIT('h4)
	) name17560 (
		_w27262_,
		_w28072_,
		_w28073_
	);
	LUT2 #(
		.INIT('h8)
	) name17561 (
		_w27257_,
		_w27281_,
		_w28074_
	);
	LUT2 #(
		.INIT('h4)
	) name17562 (
		_w27262_,
		_w28074_,
		_w28075_
	);
	LUT2 #(
		.INIT('h4)
	) name17563 (
		_w27280_,
		_w27786_,
		_w28076_
	);
	LUT2 #(
		.INIT('h8)
	) name17564 (
		_w27267_,
		_w27413_,
		_w28077_
	);
	LUT2 #(
		.INIT('h4)
	) name17565 (
		_w27262_,
		_w28077_,
		_w28078_
	);
	LUT2 #(
		.INIT('h8)
	) name17566 (
		_w27257_,
		_w27413_,
		_w28079_
	);
	LUT2 #(
		.INIT('h4)
	) name17567 (
		_w27262_,
		_w28079_,
		_w28080_
	);
	LUT2 #(
		.INIT('h4)
	) name17568 (
		_w27280_,
		_w27788_,
		_w28081_
	);
	LUT2 #(
		.INIT('h8)
	) name17569 (
		_w27299_,
		_w27333_,
		_w28082_
	);
	LUT2 #(
		.INIT('h4)
	) name17570 (
		_w27262_,
		_w28082_,
		_w28083_
	);
	LUT2 #(
		.INIT('h8)
	) name17571 (
		_w27267_,
		_w27333_,
		_w28084_
	);
	LUT2 #(
		.INIT('h4)
	) name17572 (
		_w27262_,
		_w28084_,
		_w28085_
	);
	LUT2 #(
		.INIT('h4)
	) name17573 (
		_w27280_,
		_w27790_,
		_w28086_
	);
	LUT2 #(
		.INIT('h8)
	) name17574 (
		_w27274_,
		_w27417_,
		_w28087_
	);
	LUT2 #(
		.INIT('h4)
	) name17575 (
		_w27262_,
		_w28087_,
		_w28088_
	);
	LUT2 #(
		.INIT('h8)
	) name17576 (
		_w27274_,
		_w27281_,
		_w28089_
	);
	LUT2 #(
		.INIT('h4)
	) name17577 (
		_w27262_,
		_w28089_,
		_w28090_
	);
	LUT2 #(
		.INIT('h4)
	) name17578 (
		_w27280_,
		_w27792_,
		_w28091_
	);
	LUT2 #(
		.INIT('h8)
	) name17579 (
		_w27274_,
		_w27413_,
		_w28092_
	);
	LUT2 #(
		.INIT('h4)
	) name17580 (
		_w27262_,
		_w28092_,
		_w28093_
	);
	LUT2 #(
		.INIT('h4)
	) name17581 (
		_w27280_,
		_w27794_,
		_w28094_
	);
	LUT2 #(
		.INIT('h8)
	) name17582 (
		_w27270_,
		_w27333_,
		_w28095_
	);
	LUT2 #(
		.INIT('h4)
	) name17583 (
		_w27262_,
		_w28095_,
		_w28096_
	);
	LUT2 #(
		.INIT('h4)
	) name17584 (
		_w27262_,
		_w27955_,
		_w28097_
	);
	LUT2 #(
		.INIT('h8)
	) name17585 (
		_w27288_,
		_w27417_,
		_w28098_
	);
	LUT2 #(
		.INIT('h4)
	) name17586 (
		_w27262_,
		_w28098_,
		_w28099_
	);
	LUT2 #(
		.INIT('h4)
	) name17587 (
		_w27280_,
		_w27796_,
		_w28100_
	);
	LUT2 #(
		.INIT('h4)
	) name17588 (
		_w27262_,
		_w27910_,
		_w28101_
	);
	LUT2 #(
		.INIT('h4)
	) name17589 (
		_w27280_,
		_w27798_,
		_w28102_
	);
	LUT2 #(
		.INIT('h8)
	) name17590 (
		_w27288_,
		_w27413_,
		_w28103_
	);
	LUT2 #(
		.INIT('h4)
	) name17591 (
		_w27262_,
		_w28103_,
		_w28104_
	);
	LUT2 #(
		.INIT('h8)
	) name17592 (
		_w27282_,
		_w27333_,
		_w28105_
	);
	LUT2 #(
		.INIT('h4)
	) name17593 (
		_w27490_,
		_w28105_,
		_w28106_
	);
	LUT2 #(
		.INIT('h4)
	) name17594 (
		_w27280_,
		_w27802_,
		_w28107_
	);
	LUT2 #(
		.INIT('h8)
	) name17595 (
		_w27285_,
		_w27333_,
		_w28108_
	);
	LUT2 #(
		.INIT('h4)
	) name17596 (
		_w27262_,
		_w28108_,
		_w28109_
	);
	LUT2 #(
		.INIT('h4)
	) name17597 (
		_w27280_,
		_w27804_,
		_w28110_
	);
	LUT2 #(
		.INIT('h8)
	) name17598 (
		_w27312_,
		_w27417_,
		_w28111_
	);
	LUT2 #(
		.INIT('h4)
	) name17599 (
		_w27262_,
		_w28111_,
		_w28112_
	);
	LUT2 #(
		.INIT('h4)
	) name17600 (
		_w27280_,
		_w27807_,
		_w28113_
	);
	LUT2 #(
		.INIT('h8)
	) name17601 (
		_w27293_,
		_w27333_,
		_w28114_
	);
	LUT2 #(
		.INIT('h4)
	) name17602 (
		_w27262_,
		_w28114_,
		_w28115_
	);
	LUT2 #(
		.INIT('h4)
	) name17603 (
		_w27280_,
		_w27809_,
		_w28116_
	);
	LUT2 #(
		.INIT('h4)
	) name17604 (
		_w27262_,
		_w28105_,
		_w28117_
	);
	LUT2 #(
		.INIT('h4)
	) name17605 (
		_w27490_,
		_w28114_,
		_w28118_
	);
	LUT2 #(
		.INIT('h8)
	) name17606 (
		_w27267_,
		_w27271_,
		_w28119_
	);
	LUT2 #(
		.INIT('h4)
	) name17607 (
		_w27262_,
		_w28119_,
		_w28120_
	);
	LUT2 #(
		.INIT('h8)
	) name17608 (
		_w27257_,
		_w27271_,
		_w28121_
	);
	LUT2 #(
		.INIT('h4)
	) name17609 (
		_w27262_,
		_w28121_,
		_w28122_
	);
	LUT2 #(
		.INIT('h8)
	) name17610 (
		_w27258_,
		_w27267_,
		_w28123_
	);
	LUT2 #(
		.INIT('h4)
	) name17611 (
		_w27262_,
		_w28123_,
		_w28124_
	);
	LUT2 #(
		.INIT('h4)
	) name17612 (
		_w27280_,
		_w27812_,
		_w28125_
	);
	LUT2 #(
		.INIT('h4)
	) name17613 (
		_w27262_,
		_w27725_,
		_w28126_
	);
	LUT2 #(
		.INIT('h4)
	) name17614 (
		_w27280_,
		_w27814_,
		_w28127_
	);
	LUT2 #(
		.INIT('h4)
	) name17615 (
		_w27490_,
		_w27729_,
		_w28128_
	);
	LUT2 #(
		.INIT('h4)
	) name17616 (
		_w27490_,
		_w27731_,
		_w28129_
	);
	LUT2 #(
		.INIT('h4)
	) name17617 (
		_w27280_,
		_w28059_,
		_w28130_
	);
	LUT2 #(
		.INIT('h4)
	) name17618 (
		_w27490_,
		_w27733_,
		_w28131_
	);
	LUT2 #(
		.INIT('h4)
	) name17619 (
		_w27256_,
		_w27772_,
		_w28132_
	);
	LUT2 #(
		.INIT('h4)
	) name17620 (
		_w27490_,
		_w27735_,
		_w28133_
	);
	LUT2 #(
		.INIT('h4)
	) name17621 (
		_w27280_,
		_w27816_,
		_w28134_
	);
	LUT2 #(
		.INIT('h4)
	) name17622 (
		_w27490_,
		_w27737_,
		_w28135_
	);
	LUT2 #(
		.INIT('h4)
	) name17623 (
		_w27280_,
		_w27818_,
		_w28136_
	);
	LUT2 #(
		.INIT('h4)
	) name17624 (
		_w27490_,
		_w27739_,
		_w28137_
	);
	LUT2 #(
		.INIT('h4)
	) name17625 (
		_w27490_,
		_w27741_,
		_w28138_
	);
	LUT2 #(
		.INIT('h4)
	) name17626 (
		_w27280_,
		_w27820_,
		_w28139_
	);
	LUT2 #(
		.INIT('h4)
	) name17627 (
		_w27490_,
		_w27743_,
		_w28140_
	);
	LUT2 #(
		.INIT('h4)
	) name17628 (
		_w27490_,
		_w27745_,
		_w28141_
	);
	LUT2 #(
		.INIT('h4)
	) name17629 (
		_w27280_,
		_w27823_,
		_w28142_
	);
	LUT2 #(
		.INIT('h4)
	) name17630 (
		_w27490_,
		_w27747_,
		_w28143_
	);
	LUT2 #(
		.INIT('h4)
	) name17631 (
		_w27490_,
		_w27727_,
		_w28144_
	);
	LUT2 #(
		.INIT('h4)
	) name17632 (
		_w27280_,
		_w27825_,
		_w28145_
	);
	LUT2 #(
		.INIT('h4)
	) name17633 (
		_w27490_,
		_w27750_,
		_w28146_
	);
	LUT2 #(
		.INIT('h4)
	) name17634 (
		_w27490_,
		_w27752_,
		_w28147_
	);
	LUT2 #(
		.INIT('h4)
	) name17635 (
		_w27280_,
		_w27827_,
		_w28148_
	);
	LUT2 #(
		.INIT('h4)
	) name17636 (
		_w27490_,
		_w27756_,
		_w28149_
	);
	LUT2 #(
		.INIT('h4)
	) name17637 (
		_w27490_,
		_w27758_,
		_w28150_
	);
	LUT2 #(
		.INIT('h4)
	) name17638 (
		_w27490_,
		_w27760_,
		_w28151_
	);
	LUT2 #(
		.INIT('h4)
	) name17639 (
		_w27490_,
		_w27762_,
		_w28152_
	);
	LUT2 #(
		.INIT('h4)
	) name17640 (
		_w27490_,
		_w27764_,
		_w28153_
	);
	LUT2 #(
		.INIT('h4)
	) name17641 (
		_w27490_,
		_w27766_,
		_w28154_
	);
	LUT2 #(
		.INIT('h4)
	) name17642 (
		_w27490_,
		_w27768_,
		_w28155_
	);
	LUT2 #(
		.INIT('h4)
	) name17643 (
		_w27490_,
		_w27770_,
		_w28156_
	);
	LUT2 #(
		.INIT('h4)
	) name17644 (
		_w27490_,
		_w27772_,
		_w28157_
	);
	LUT2 #(
		.INIT('h4)
	) name17645 (
		_w27490_,
		_w27774_,
		_w28158_
	);
	LUT2 #(
		.INIT('h4)
	) name17646 (
		_w27490_,
		_w27776_,
		_w28159_
	);
	LUT2 #(
		.INIT('h4)
	) name17647 (
		_w27490_,
		_w27778_,
		_w28160_
	);
	LUT2 #(
		.INIT('h4)
	) name17648 (
		_w27280_,
		_w27831_,
		_w28161_
	);
	LUT2 #(
		.INIT('h4)
	) name17649 (
		_w27490_,
		_w27780_,
		_w28162_
	);
	LUT2 #(
		.INIT('h4)
	) name17650 (
		_w27490_,
		_w27782_,
		_w28163_
	);
	LUT2 #(
		.INIT('h4)
	) name17651 (
		_w27490_,
		_w27784_,
		_w28164_
	);
	LUT2 #(
		.INIT('h4)
	) name17652 (
		_w27280_,
		_w27833_,
		_w28165_
	);
	LUT2 #(
		.INIT('h4)
	) name17653 (
		_w27490_,
		_w27786_,
		_w28166_
	);
	LUT2 #(
		.INIT('h4)
	) name17654 (
		_w27490_,
		_w27788_,
		_w28167_
	);
	LUT2 #(
		.INIT('h4)
	) name17655 (
		_w27490_,
		_w27790_,
		_w28168_
	);
	LUT2 #(
		.INIT('h4)
	) name17656 (
		_w27280_,
		_w28056_,
		_w28169_
	);
	LUT2 #(
		.INIT('h4)
	) name17657 (
		_w27280_,
		_w27835_,
		_w28170_
	);
	LUT2 #(
		.INIT('h4)
	) name17658 (
		_w27256_,
		_w27747_,
		_w28171_
	);
	LUT2 #(
		.INIT('h4)
	) name17659 (
		_w27490_,
		_w27792_,
		_w28172_
	);
	LUT2 #(
		.INIT('h4)
	) name17660 (
		_w27490_,
		_w27794_,
		_w28173_
	);
	LUT2 #(
		.INIT('h4)
	) name17661 (
		_w27280_,
		_w27837_,
		_w28174_
	);
	LUT2 #(
		.INIT('h4)
	) name17662 (
		_w27490_,
		_w27796_,
		_w28175_
	);
	LUT2 #(
		.INIT('h4)
	) name17663 (
		_w27490_,
		_w27798_,
		_w28176_
	);
	LUT2 #(
		.INIT('h4)
	) name17664 (
		_w27490_,
		_w27802_,
		_w28177_
	);
	LUT2 #(
		.INIT('h4)
	) name17665 (
		_w27280_,
		_w27840_,
		_w28178_
	);
	LUT2 #(
		.INIT('h4)
	) name17666 (
		_w27490_,
		_w27804_,
		_w28179_
	);
	LUT2 #(
		.INIT('h4)
	) name17667 (
		_w27280_,
		_w27842_,
		_w28180_
	);
	LUT2 #(
		.INIT('h4)
	) name17668 (
		_w27490_,
		_w27807_,
		_w28181_
	);
	LUT2 #(
		.INIT('h4)
	) name17669 (
		_w27490_,
		_w27809_,
		_w28182_
	);
	LUT2 #(
		.INIT('h4)
	) name17670 (
		_w27490_,
		_w27812_,
		_w28183_
	);
	LUT2 #(
		.INIT('h4)
	) name17671 (
		_w27490_,
		_w27814_,
		_w28184_
	);
	LUT2 #(
		.INIT('h4)
	) name17672 (
		_w27280_,
		_w27845_,
		_w28185_
	);
	LUT2 #(
		.INIT('h4)
	) name17673 (
		_w27280_,
		_w27847_,
		_w28186_
	);
	LUT2 #(
		.INIT('h4)
	) name17674 (
		_w27490_,
		_w27816_,
		_w28187_
	);
	LUT2 #(
		.INIT('h4)
	) name17675 (
		_w27490_,
		_w27818_,
		_w28188_
	);
	LUT2 #(
		.INIT('h4)
	) name17676 (
		_w27490_,
		_w27820_,
		_w28189_
	);
	LUT2 #(
		.INIT('h4)
	) name17677 (
		_w27280_,
		_w27852_,
		_w28190_
	);
	LUT2 #(
		.INIT('h4)
	) name17678 (
		_w27490_,
		_w27823_,
		_w28191_
	);
	LUT2 #(
		.INIT('h4)
	) name17679 (
		_w27490_,
		_w27825_,
		_w28192_
	);
	LUT2 #(
		.INIT('h4)
	) name17680 (
		_w27490_,
		_w27827_,
		_w28193_
	);
	LUT2 #(
		.INIT('h4)
	) name17681 (
		_w27280_,
		_w27854_,
		_w28194_
	);
	LUT2 #(
		.INIT('h4)
	) name17682 (
		_w27280_,
		_w27856_,
		_w28195_
	);
	LUT2 #(
		.INIT('h4)
	) name17683 (
		_w27490_,
		_w27831_,
		_w28196_
	);
	LUT2 #(
		.INIT('h4)
	) name17684 (
		_w27280_,
		_w27858_,
		_w28197_
	);
	LUT2 #(
		.INIT('h4)
	) name17685 (
		_w27490_,
		_w27833_,
		_w28198_
	);
	LUT2 #(
		.INIT('h4)
	) name17686 (
		_w27280_,
		_w27860_,
		_w28199_
	);
	LUT2 #(
		.INIT('h4)
	) name17687 (
		_w27490_,
		_w27835_,
		_w28200_
	);
	LUT2 #(
		.INIT('h4)
	) name17688 (
		_w27280_,
		_w27862_,
		_w28201_
	);
	LUT2 #(
		.INIT('h4)
	) name17689 (
		_w27490_,
		_w27837_,
		_w28202_
	);
	LUT2 #(
		.INIT('h4)
	) name17690 (
		_w27280_,
		_w27864_,
		_w28203_
	);
	LUT2 #(
		.INIT('h4)
	) name17691 (
		_w27490_,
		_w27840_,
		_w28204_
	);
	LUT2 #(
		.INIT('h4)
	) name17692 (
		_w27280_,
		_w27867_,
		_w28205_
	);
	LUT2 #(
		.INIT('h4)
	) name17693 (
		_w27490_,
		_w27842_,
		_w28206_
	);
	LUT2 #(
		.INIT('h4)
	) name17694 (
		_w27280_,
		_w27869_,
		_w28207_
	);
	LUT2 #(
		.INIT('h4)
	) name17695 (
		_w27490_,
		_w27845_,
		_w28208_
	);
	LUT2 #(
		.INIT('h4)
	) name17696 (
		_w27280_,
		_w27871_,
		_w28209_
	);
	LUT2 #(
		.INIT('h4)
	) name17697 (
		_w27490_,
		_w27847_,
		_w28210_
	);
	LUT2 #(
		.INIT('h4)
	) name17698 (
		_w27280_,
		_w27873_,
		_w28211_
	);
	LUT2 #(
		.INIT('h4)
	) name17699 (
		_w27490_,
		_w27852_,
		_w28212_
	);
	LUT2 #(
		.INIT('h4)
	) name17700 (
		_w27280_,
		_w27875_,
		_w28213_
	);
	LUT2 #(
		.INIT('h4)
	) name17701 (
		_w27490_,
		_w27854_,
		_w28214_
	);
	LUT2 #(
		.INIT('h4)
	) name17702 (
		_w27280_,
		_w27877_,
		_w28215_
	);
	LUT2 #(
		.INIT('h4)
	) name17703 (
		_w27490_,
		_w27856_,
		_w28216_
	);
	LUT2 #(
		.INIT('h4)
	) name17704 (
		_w27490_,
		_w27858_,
		_w28217_
	);
	LUT2 #(
		.INIT('h4)
	) name17705 (
		_w27490_,
		_w27860_,
		_w28218_
	);
	LUT2 #(
		.INIT('h4)
	) name17706 (
		_w27490_,
		_w27862_,
		_w28219_
	);
	LUT2 #(
		.INIT('h4)
	) name17707 (
		_w27280_,
		_w27879_,
		_w28220_
	);
	LUT2 #(
		.INIT('h4)
	) name17708 (
		_w27490_,
		_w27864_,
		_w28221_
	);
	LUT2 #(
		.INIT('h4)
	) name17709 (
		_w27490_,
		_w27867_,
		_w28222_
	);
	LUT2 #(
		.INIT('h4)
	) name17710 (
		_w27490_,
		_w27869_,
		_w28223_
	);
	LUT2 #(
		.INIT('h4)
	) name17711 (
		_w27490_,
		_w27871_,
		_w28224_
	);
	LUT2 #(
		.INIT('h4)
	) name17712 (
		_w27490_,
		_w27873_,
		_w28225_
	);
	LUT2 #(
		.INIT('h4)
	) name17713 (
		_w27490_,
		_w27875_,
		_w28226_
	);
	LUT2 #(
		.INIT('h4)
	) name17714 (
		_w27280_,
		_w27881_,
		_w28227_
	);
	LUT2 #(
		.INIT('h4)
	) name17715 (
		_w27490_,
		_w27877_,
		_w28228_
	);
	LUT2 #(
		.INIT('h4)
	) name17716 (
		_w27280_,
		_w27883_,
		_w28229_
	);
	LUT2 #(
		.INIT('h4)
	) name17717 (
		_w27490_,
		_w27879_,
		_w28230_
	);
	LUT2 #(
		.INIT('h4)
	) name17718 (
		_w27280_,
		_w27885_,
		_w28231_
	);
	LUT2 #(
		.INIT('h4)
	) name17719 (
		_w27490_,
		_w27881_,
		_w28232_
	);
	LUT2 #(
		.INIT('h4)
	) name17720 (
		_w27280_,
		_w27887_,
		_w28233_
	);
	LUT2 #(
		.INIT('h4)
	) name17721 (
		_w27490_,
		_w27883_,
		_w28234_
	);
	LUT2 #(
		.INIT('h4)
	) name17722 (
		_w27490_,
		_w27885_,
		_w28235_
	);
	LUT2 #(
		.INIT('h4)
	) name17723 (
		_w27490_,
		_w27887_,
		_w28236_
	);
	LUT2 #(
		.INIT('h4)
	) name17724 (
		_w27490_,
		_w27890_,
		_w28237_
	);
	LUT2 #(
		.INIT('h4)
	) name17725 (
		_w27280_,
		_w27890_,
		_w28238_
	);
	LUT2 #(
		.INIT('h4)
	) name17726 (
		_w27490_,
		_w27892_,
		_w28239_
	);
	LUT2 #(
		.INIT('h4)
	) name17727 (
		_w27490_,
		_w27894_,
		_w28240_
	);
	LUT2 #(
		.INIT('h4)
	) name17728 (
		_w27490_,
		_w27896_,
		_w28241_
	);
	LUT2 #(
		.INIT('h4)
	) name17729 (
		_w27490_,
		_w27898_,
		_w28242_
	);
	LUT2 #(
		.INIT('h4)
	) name17730 (
		_w27280_,
		_w27892_,
		_w28243_
	);
	LUT2 #(
		.INIT('h4)
	) name17731 (
		_w27490_,
		_w28095_,
		_w28244_
	);
	LUT2 #(
		.INIT('h4)
	) name17732 (
		_w27490_,
		_w27900_,
		_w28245_
	);
	LUT2 #(
		.INIT('h4)
	) name17733 (
		_w27280_,
		_w27894_,
		_w28246_
	);
	LUT2 #(
		.INIT('h4)
	) name17734 (
		_w27490_,
		_w27902_,
		_w28247_
	);
	LUT2 #(
		.INIT('h4)
	) name17735 (
		_w27280_,
		_w27896_,
		_w28248_
	);
	LUT2 #(
		.INIT('h4)
	) name17736 (
		_w27490_,
		_w27904_,
		_w28249_
	);
	LUT2 #(
		.INIT('h4)
	) name17737 (
		_w27280_,
		_w27898_,
		_w28250_
	);
	LUT2 #(
		.INIT('h4)
	) name17738 (
		_w27490_,
		_w27906_,
		_w28251_
	);
	LUT2 #(
		.INIT('h4)
	) name17739 (
		_w27490_,
		_w27908_,
		_w28252_
	);
	LUT2 #(
		.INIT('h4)
	) name17740 (
		_w27280_,
		_w28050_,
		_w28253_
	);
	LUT2 #(
		.INIT('h4)
	) name17741 (
		_w27280_,
		_w27900_,
		_w28254_
	);
	LUT2 #(
		.INIT('h4)
	) name17742 (
		_w27490_,
		_w27912_,
		_w28255_
	);
	LUT2 #(
		.INIT('h4)
	) name17743 (
		_w27490_,
		_w27914_,
		_w28256_
	);
	LUT2 #(
		.INIT('h4)
	) name17744 (
		_w27490_,
		_w27916_,
		_w28257_
	);
	LUT2 #(
		.INIT('h4)
	) name17745 (
		_w27490_,
		_w27918_,
		_w28258_
	);
	LUT2 #(
		.INIT('h4)
	) name17746 (
		_w27280_,
		_w27902_,
		_w28259_
	);
	LUT2 #(
		.INIT('h4)
	) name17747 (
		_w27490_,
		_w27920_,
		_w28260_
	);
	LUT2 #(
		.INIT('h4)
	) name17748 (
		_w27280_,
		_w27991_,
		_w28261_
	);
	LUT2 #(
		.INIT('h4)
	) name17749 (
		_w27490_,
		_w27923_,
		_w28262_
	);
	LUT2 #(
		.INIT('h4)
	) name17750 (
		_w27490_,
		_w27925_,
		_w28263_
	);
	LUT2 #(
		.INIT('h4)
	) name17751 (
		_w27490_,
		_w27927_,
		_w28264_
	);
	LUT2 #(
		.INIT('h4)
	) name17752 (
		_w27280_,
		_w27904_,
		_w28265_
	);
	LUT2 #(
		.INIT('h4)
	) name17753 (
		_w27490_,
		_w28092_,
		_w28266_
	);
	LUT2 #(
		.INIT('h4)
	) name17754 (
		_w27280_,
		_w27906_,
		_w28267_
	);
	LUT2 #(
		.INIT('h4)
	) name17755 (
		_w27490_,
		_w27930_,
		_w28268_
	);
	LUT2 #(
		.INIT('h4)
	) name17756 (
		_w27280_,
		_w27908_,
		_w28269_
	);
	LUT2 #(
		.INIT('h4)
	) name17757 (
		_w27490_,
		_w27932_,
		_w28270_
	);
	LUT2 #(
		.INIT('h4)
	) name17758 (
		_w27490_,
		_w27934_,
		_w28271_
	);
	LUT2 #(
		.INIT('h4)
	) name17759 (
		_w27490_,
		_w27937_,
		_w28272_
	);
	LUT2 #(
		.INIT('h4)
	) name17760 (
		_w27490_,
		_w27940_,
		_w28273_
	);
	LUT2 #(
		.INIT('h4)
	) name17761 (
		_w27280_,
		_w27912_,
		_w28274_
	);
	LUT2 #(
		.INIT('h4)
	) name17762 (
		_w27490_,
		_w27942_,
		_w28275_
	);
	LUT2 #(
		.INIT('h4)
	) name17763 (
		_w27490_,
		_w27944_,
		_w28276_
	);
	LUT2 #(
		.INIT('h4)
	) name17764 (
		_w27280_,
		_w27914_,
		_w28277_
	);
	LUT2 #(
		.INIT('h4)
	) name17765 (
		_w27490_,
		_w27946_,
		_w28278_
	);
	LUT2 #(
		.INIT('h4)
	) name17766 (
		_w27490_,
		_w27948_,
		_w28279_
	);
	LUT2 #(
		.INIT('h4)
	) name17767 (
		_w27280_,
		_w27916_,
		_w28280_
	);
	LUT2 #(
		.INIT('h4)
	) name17768 (
		_w27490_,
		_w27950_,
		_w28281_
	);
	LUT2 #(
		.INIT('h4)
	) name17769 (
		_w27490_,
		_w27953_,
		_w28282_
	);
	LUT2 #(
		.INIT('h4)
	) name17770 (
		_w27280_,
		_w27918_,
		_w28283_
	);
	LUT2 #(
		.INIT('h4)
	) name17771 (
		_w27280_,
		_w27920_,
		_w28284_
	);
	LUT2 #(
		.INIT('h4)
	) name17772 (
		_w27490_,
		_w27957_,
		_w28285_
	);
	LUT2 #(
		.INIT('h4)
	) name17773 (
		_w27490_,
		_w27960_,
		_w28286_
	);
	LUT2 #(
		.INIT('h4)
	) name17774 (
		_w27280_,
		_w28092_,
		_w28287_
	);
	LUT2 #(
		.INIT('h4)
	) name17775 (
		_w27280_,
		_w27923_,
		_w28288_
	);
	LUT2 #(
		.INIT('h4)
	) name17776 (
		_w27490_,
		_w27962_,
		_w28289_
	);
	LUT2 #(
		.INIT('h4)
	) name17777 (
		_w27490_,
		_w27965_,
		_w28290_
	);
	LUT2 #(
		.INIT('h4)
	) name17778 (
		_w27280_,
		_w27925_,
		_w28291_
	);
	LUT2 #(
		.INIT('h4)
	) name17779 (
		_w27490_,
		_w27967_,
		_w28292_
	);
	LUT2 #(
		.INIT('h4)
	) name17780 (
		_w27490_,
		_w27970_,
		_w28293_
	);
	LUT2 #(
		.INIT('h4)
	) name17781 (
		_w27280_,
		_w27927_,
		_w28294_
	);
	LUT2 #(
		.INIT('h4)
	) name17782 (
		_w27490_,
		_w27972_,
		_w28295_
	);
	LUT2 #(
		.INIT('h4)
	) name17783 (
		_w27490_,
		_w27975_,
		_w28296_
	);
	LUT2 #(
		.INIT('h4)
	) name17784 (
		_w27490_,
		_w27977_,
		_w28297_
	);
	LUT2 #(
		.INIT('h4)
	) name17785 (
		_w27490_,
		_w27980_,
		_w28298_
	);
	LUT2 #(
		.INIT('h4)
	) name17786 (
		_w27490_,
		_w27982_,
		_w28299_
	);
	LUT2 #(
		.INIT('h4)
	) name17787 (
		_w27490_,
		_w27984_,
		_w28300_
	);
	LUT2 #(
		.INIT('h4)
	) name17788 (
		_w27280_,
		_w27930_,
		_w28301_
	);
	LUT2 #(
		.INIT('h4)
	) name17789 (
		_w27490_,
		_w27986_,
		_w28302_
	);
	LUT2 #(
		.INIT('h4)
	) name17790 (
		_w27490_,
		_w27988_,
		_w28303_
	);
	LUT2 #(
		.INIT('h4)
	) name17791 (
		_w27490_,
		_w27991_,
		_w28304_
	);
	LUT2 #(
		.INIT('h4)
	) name17792 (
		_w27490_,
		_w27994_,
		_w28305_
	);
	LUT2 #(
		.INIT('h4)
	) name17793 (
		_w27280_,
		_w27932_,
		_w28306_
	);
	LUT2 #(
		.INIT('h4)
	) name17794 (
		_w27490_,
		_w27996_,
		_w28307_
	);
	LUT2 #(
		.INIT('h4)
	) name17795 (
		_w27280_,
		_w27934_,
		_w28308_
	);
	LUT2 #(
		.INIT('h4)
	) name17796 (
		_w27490_,
		_w27999_,
		_w28309_
	);
	LUT2 #(
		.INIT('h4)
	) name17797 (
		_w27490_,
		_w28001_,
		_w28310_
	);
	LUT2 #(
		.INIT('h4)
	) name17798 (
		_w27280_,
		_w27937_,
		_w28311_
	);
	LUT2 #(
		.INIT('h4)
	) name17799 (
		_w27490_,
		_w28005_,
		_w28312_
	);
	LUT2 #(
		.INIT('h4)
	) name17800 (
		_w27490_,
		_w28007_,
		_w28313_
	);
	LUT2 #(
		.INIT('h4)
	) name17801 (
		_w27490_,
		_w28010_,
		_w28314_
	);
	LUT2 #(
		.INIT('h4)
	) name17802 (
		_w27490_,
		_w28012_,
		_w28315_
	);
	LUT2 #(
		.INIT('h4)
	) name17803 (
		_w27280_,
		_w27940_,
		_w28316_
	);
	LUT2 #(
		.INIT('h4)
	) name17804 (
		_w27490_,
		_w28014_,
		_w28317_
	);
	LUT2 #(
		.INIT('h4)
	) name17805 (
		_w27490_,
		_w28016_,
		_w28318_
	);
	LUT2 #(
		.INIT('h4)
	) name17806 (
		_w27280_,
		_w27942_,
		_w28319_
	);
	LUT2 #(
		.INIT('h4)
	) name17807 (
		_w27490_,
		_w28018_,
		_w28320_
	);
	LUT2 #(
		.INIT('h4)
	) name17808 (
		_w27280_,
		_w27944_,
		_w28321_
	);
	LUT2 #(
		.INIT('h4)
	) name17809 (
		_w27490_,
		_w28021_,
		_w28322_
	);
	LUT2 #(
		.INIT('h4)
	) name17810 (
		_w27280_,
		_w27946_,
		_w28323_
	);
	LUT2 #(
		.INIT('h4)
	) name17811 (
		_w27490_,
		_w28023_,
		_w28324_
	);
	LUT2 #(
		.INIT('h4)
	) name17812 (
		_w27490_,
		_w28026_,
		_w28325_
	);
	LUT2 #(
		.INIT('h4)
	) name17813 (
		_w27280_,
		_w27948_,
		_w28326_
	);
	LUT2 #(
		.INIT('h4)
	) name17814 (
		_w27490_,
		_w28028_,
		_w28327_
	);
	LUT2 #(
		.INIT('h4)
	) name17815 (
		_w27280_,
		_w27950_,
		_w28328_
	);
	LUT2 #(
		.INIT('h4)
	) name17816 (
		_w27490_,
		_w28079_,
		_w28329_
	);
	LUT2 #(
		.INIT('h4)
	) name17817 (
		_w27490_,
		_w27754_,
		_w28330_
	);
	LUT2 #(
		.INIT('h4)
	) name17818 (
		_w27280_,
		_w27953_,
		_w28331_
	);
	LUT2 #(
		.INIT('h4)
	) name17819 (
		_w27490_,
		_w28034_,
		_w28332_
	);
	LUT2 #(
		.INIT('h4)
	) name17820 (
		_w27490_,
		_w28036_,
		_w28333_
	);
	LUT2 #(
		.INIT('h4)
	) name17821 (
		_w27490_,
		_w28077_,
		_w28334_
	);
	LUT2 #(
		.INIT('h4)
	) name17822 (
		_w27490_,
		_w28039_,
		_w28335_
	);
	LUT2 #(
		.INIT('h4)
	) name17823 (
		_w27490_,
		_w28041_,
		_w28336_
	);
	LUT2 #(
		.INIT('h4)
	) name17824 (
		_w27490_,
		_w28044_,
		_w28337_
	);
	LUT2 #(
		.INIT('h4)
	) name17825 (
		_w27280_,
		_w27957_,
		_w28338_
	);
	LUT2 #(
		.INIT('h4)
	) name17826 (
		_w27490_,
		_w28047_,
		_w28339_
	);
	LUT2 #(
		.INIT('h4)
	) name17827 (
		_w27490_,
		_w28074_,
		_w28340_
	);
	LUT2 #(
		.INIT('h4)
	) name17828 (
		_w27280_,
		_w27960_,
		_w28341_
	);
	LUT2 #(
		.INIT('h4)
	) name17829 (
		_w27280_,
		_w27962_,
		_w28342_
	);
	LUT2 #(
		.INIT('h4)
	) name17830 (
		_w27490_,
		_w28050_,
		_w28343_
	);
	LUT2 #(
		.INIT('h4)
	) name17831 (
		_w27490_,
		_w28053_,
		_w28344_
	);
	LUT2 #(
		.INIT('h4)
	) name17832 (
		_w27280_,
		_w27965_,
		_w28345_
	);
	LUT2 #(
		.INIT('h4)
	) name17833 (
		_w27280_,
		_w27967_,
		_w28346_
	);
	LUT2 #(
		.INIT('h4)
	) name17834 (
		_w27490_,
		_w28056_,
		_w28347_
	);
	LUT2 #(
		.INIT('h4)
	) name17835 (
		_w27490_,
		_w28059_,
		_w28348_
	);
	LUT2 #(
		.INIT('h4)
	) name17836 (
		_w27280_,
		_w27970_,
		_w28349_
	);
	LUT2 #(
		.INIT('h4)
	) name17837 (
		_w27490_,
		_w28062_,
		_w28350_
	);
	LUT2 #(
		.INIT('h4)
	) name17838 (
		_w27490_,
		_w28072_,
		_w28351_
	);
	LUT2 #(
		.INIT('h4)
	) name17839 (
		_w27280_,
		_w27972_,
		_w28352_
	);
	LUT2 #(
		.INIT('h4)
	) name17840 (
		_w27490_,
		_w28064_,
		_w28353_
	);
	LUT2 #(
		.INIT('h4)
	) name17841 (
		_w27490_,
		_w28066_,
		_w28354_
	);
	LUT2 #(
		.INIT('h4)
	) name17842 (
		_w27280_,
		_w27975_,
		_w28355_
	);
	LUT2 #(
		.INIT('h4)
	) name17843 (
		_w27490_,
		_w27850_,
		_w28356_
	);
	LUT2 #(
		.INIT('h4)
	) name17844 (
		_w27490_,
		_w28069_,
		_w28357_
	);
	LUT2 #(
		.INIT('h4)
	) name17845 (
		_w27280_,
		_w27977_,
		_w28358_
	);
	LUT2 #(
		.INIT('h4)
	) name17846 (
		_w27280_,
		_w27980_,
		_w28359_
	);
	LUT2 #(
		.INIT('h4)
	) name17847 (
		_w27280_,
		_w27982_,
		_w28360_
	);
	LUT2 #(
		.INIT('h4)
	) name17848 (
		_w27490_,
		_w28082_,
		_w28361_
	);
	LUT2 #(
		.INIT('h4)
	) name17849 (
		_w27490_,
		_w28084_,
		_w28362_
	);
	LUT2 #(
		.INIT('h4)
	) name17850 (
		_w27280_,
		_w27984_,
		_w28363_
	);
	LUT2 #(
		.INIT('h4)
	) name17851 (
		_w27490_,
		_w28087_,
		_w28364_
	);
	LUT2 #(
		.INIT('h4)
	) name17852 (
		_w27280_,
		_w27986_,
		_w28365_
	);
	LUT2 #(
		.INIT('h4)
	) name17853 (
		_w27490_,
		_w28089_,
		_w28366_
	);
	LUT2 #(
		.INIT('h4)
	) name17854 (
		_w27280_,
		_w27988_,
		_w28367_
	);
	LUT2 #(
		.INIT('h4)
	) name17855 (
		_w27280_,
		_w27994_,
		_w28368_
	);
	LUT2 #(
		.INIT('h4)
	) name17856 (
		_w27490_,
		_w27955_,
		_w28369_
	);
	LUT2 #(
		.INIT('h4)
	) name17857 (
		_w27490_,
		_w28098_,
		_w28370_
	);
	LUT2 #(
		.INIT('h4)
	) name17858 (
		_w27280_,
		_w27996_,
		_w28371_
	);
	LUT2 #(
		.INIT('h4)
	) name17859 (
		_w27490_,
		_w27910_,
		_w28372_
	);
	LUT2 #(
		.INIT('h4)
	) name17860 (
		_w27490_,
		_w28103_,
		_w28373_
	);
	LUT2 #(
		.INIT('h4)
	) name17861 (
		_w27280_,
		_w27999_,
		_w28374_
	);
	LUT2 #(
		.INIT('h4)
	) name17862 (
		_w27490_,
		_w28108_,
		_w28375_
	);
	LUT2 #(
		.INIT('h4)
	) name17863 (
		_w27490_,
		_w28111_,
		_w28376_
	);
	LUT2 #(
		.INIT('h4)
	) name17864 (
		_w27280_,
		_w28001_,
		_w28377_
	);
	LUT2 #(
		.INIT('h4)
	) name17865 (
		_w27280_,
		_w28005_,
		_w28378_
	);
	LUT2 #(
		.INIT('h4)
	) name17866 (
		_w27280_,
		_w28007_,
		_w28379_
	);
	LUT2 #(
		.INIT('h4)
	) name17867 (
		_w27490_,
		_w28119_,
		_w28380_
	);
	LUT2 #(
		.INIT('h4)
	) name17868 (
		_w27490_,
		_w28121_,
		_w28381_
	);
	LUT2 #(
		.INIT('h4)
	) name17869 (
		_w27280_,
		_w28010_,
		_w28382_
	);
	LUT2 #(
		.INIT('h4)
	) name17870 (
		_w27490_,
		_w28123_,
		_w28383_
	);
	LUT2 #(
		.INIT('h4)
	) name17871 (
		_w27280_,
		_w28012_,
		_w28384_
	);
	LUT2 #(
		.INIT('h4)
	) name17872 (
		_w27490_,
		_w27725_,
		_w28385_
	);
	LUT2 #(
		.INIT('h4)
	) name17873 (
		_w27280_,
		_w28014_,
		_w28386_
	);
	LUT2 #(
		.INIT('h4)
	) name17874 (
		_w27280_,
		_w28016_,
		_w28387_
	);
	LUT2 #(
		.INIT('h4)
	) name17875 (
		_w27280_,
		_w28111_,
		_w28388_
	);
	LUT2 #(
		.INIT('h4)
	) name17876 (
		_w27256_,
		_w27743_,
		_w28389_
	);
	LUT2 #(
		.INIT('h4)
	) name17877 (
		_w27280_,
		_w28018_,
		_w28390_
	);
	LUT2 #(
		.INIT('h4)
	) name17878 (
		_w27256_,
		_w27741_,
		_w28391_
	);
	LUT2 #(
		.INIT('h4)
	) name17879 (
		_w27256_,
		_w27760_,
		_w28392_
	);
	LUT2 #(
		.INIT('h4)
	) name17880 (
		_w27280_,
		_w28021_,
		_w28393_
	);
	LUT2 #(
		.INIT('h4)
	) name17881 (
		_w27280_,
		_w28023_,
		_w28394_
	);
	LUT2 #(
		.INIT('h4)
	) name17882 (
		_w27256_,
		_w27788_,
		_w28395_
	);
	LUT2 #(
		.INIT('h4)
	) name17883 (
		_w27280_,
		_w28026_,
		_w28396_
	);
	LUT2 #(
		.INIT('h4)
	) name17884 (
		_w27280_,
		_w28028_,
		_w28397_
	);
	LUT2 #(
		.INIT('h4)
	) name17885 (
		_w27280_,
		_w28034_,
		_w28398_
	);
	LUT2 #(
		.INIT('h4)
	) name17886 (
		_w27280_,
		_w28036_,
		_w28399_
	);
	LUT2 #(
		.INIT('h4)
	) name17887 (
		_w27280_,
		_w28039_,
		_w28400_
	);
	LUT2 #(
		.INIT('h4)
	) name17888 (
		_w27280_,
		_w28041_,
		_w28401_
	);
	LUT2 #(
		.INIT('h4)
	) name17889 (
		_w27280_,
		_w28044_,
		_w28402_
	);
	LUT2 #(
		.INIT('h4)
	) name17890 (
		_w27280_,
		_w28047_,
		_w28403_
	);
	LUT2 #(
		.INIT('h4)
	) name17891 (
		_w27280_,
		_w28053_,
		_w28404_
	);
	LUT2 #(
		.INIT('h4)
	) name17892 (
		_w27256_,
		_w27733_,
		_w28405_
	);
	LUT2 #(
		.INIT('h4)
	) name17893 (
		_w27280_,
		_w28064_,
		_w28406_
	);
	LUT2 #(
		.INIT('h4)
	) name17894 (
		_w27280_,
		_w28066_,
		_w28407_
	);
	LUT2 #(
		.INIT('h4)
	) name17895 (
		_w27280_,
		_w28069_,
		_w28408_
	);
	LUT2 #(
		.INIT('h4)
	) name17896 (
		_w27280_,
		_w28072_,
		_w28409_
	);
	LUT2 #(
		.INIT('h4)
	) name17897 (
		_w27280_,
		_w28074_,
		_w28410_
	);
	LUT2 #(
		.INIT('h4)
	) name17898 (
		_w27280_,
		_w28077_,
		_w28411_
	);
	LUT2 #(
		.INIT('h4)
	) name17899 (
		_w27280_,
		_w28079_,
		_w28412_
	);
	LUT2 #(
		.INIT('h4)
	) name17900 (
		_w27280_,
		_w28082_,
		_w28413_
	);
	LUT2 #(
		.INIT('h4)
	) name17901 (
		_w27280_,
		_w28084_,
		_w28414_
	);
	LUT2 #(
		.INIT('h4)
	) name17902 (
		_w27280_,
		_w28087_,
		_w28415_
	);
	LUT2 #(
		.INIT('h4)
	) name17903 (
		_w27280_,
		_w28089_,
		_w28416_
	);
	LUT2 #(
		.INIT('h4)
	) name17904 (
		_w27280_,
		_w28095_,
		_w28417_
	);
	LUT2 #(
		.INIT('h4)
	) name17905 (
		_w27280_,
		_w28098_,
		_w28418_
	);
	LUT2 #(
		.INIT('h4)
	) name17906 (
		_w27280_,
		_w28103_,
		_w28419_
	);
	LUT2 #(
		.INIT('h4)
	) name17907 (
		_w27280_,
		_w28108_,
		_w28420_
	);
	LUT2 #(
		.INIT('h4)
	) name17908 (
		_w27256_,
		_w27752_,
		_w28421_
	);
	LUT2 #(
		.INIT('h4)
	) name17909 (
		_w27280_,
		_w28114_,
		_w28422_
	);
	LUT2 #(
		.INIT('h4)
	) name17910 (
		_w27280_,
		_w28105_,
		_w28423_
	);
	LUT2 #(
		.INIT('h4)
	) name17911 (
		_w27256_,
		_w27750_,
		_w28424_
	);
	LUT2 #(
		.INIT('h4)
	) name17912 (
		_w27280_,
		_w28119_,
		_w28425_
	);
	LUT2 #(
		.INIT('h4)
	) name17913 (
		_w27280_,
		_w28121_,
		_w28426_
	);
	LUT2 #(
		.INIT('h4)
	) name17914 (
		_w27280_,
		_w28123_,
		_w28427_
	);
	LUT2 #(
		.INIT('h4)
	) name17915 (
		_w27280_,
		_w27725_,
		_w28428_
	);
	LUT2 #(
		.INIT('h4)
	) name17916 (
		_w27256_,
		_w27729_,
		_w28429_
	);
	LUT2 #(
		.INIT('h4)
	) name17917 (
		_w27256_,
		_w27735_,
		_w28430_
	);
	LUT2 #(
		.INIT('h4)
	) name17918 (
		_w27256_,
		_w27737_,
		_w28431_
	);
	LUT2 #(
		.INIT('h4)
	) name17919 (
		_w27256_,
		_w27739_,
		_w28432_
	);
	LUT2 #(
		.INIT('h4)
	) name17920 (
		_w27256_,
		_w27745_,
		_w28433_
	);
	LUT2 #(
		.INIT('h4)
	) name17921 (
		_w27256_,
		_w27756_,
		_w28434_
	);
	LUT2 #(
		.INIT('h4)
	) name17922 (
		_w27256_,
		_w27758_,
		_w28435_
	);
	LUT2 #(
		.INIT('h4)
	) name17923 (
		_w27256_,
		_w27762_,
		_w28436_
	);
	LUT2 #(
		.INIT('h4)
	) name17924 (
		_w27256_,
		_w27780_,
		_w28437_
	);
	LUT2 #(
		.INIT('h4)
	) name17925 (
		_w27256_,
		_w27794_,
		_w28438_
	);
	LUT2 #(
		.INIT('h4)
	) name17926 (
		_w27256_,
		_w27796_,
		_w28439_
	);
	LUT2 #(
		.INIT('h4)
	) name17927 (
		_w27256_,
		_w27798_,
		_w28440_
	);
	LUT2 #(
		.INIT('h4)
	) name17928 (
		_w27256_,
		_w27802_,
		_w28441_
	);
	LUT2 #(
		.INIT('h4)
	) name17929 (
		_w27256_,
		_w27804_,
		_w28442_
	);
	LUT2 #(
		.INIT('h4)
	) name17930 (
		_w27256_,
		_w27807_,
		_w28443_
	);
	LUT2 #(
		.INIT('h4)
	) name17931 (
		_w27256_,
		_w27809_,
		_w28444_
	);
	LUT2 #(
		.INIT('h4)
	) name17932 (
		_w27256_,
		_w27812_,
		_w28445_
	);
	LUT2 #(
		.INIT('h4)
	) name17933 (
		_w27256_,
		_w27814_,
		_w28446_
	);
	LUT2 #(
		.INIT('h4)
	) name17934 (
		_w27256_,
		_w27816_,
		_w28447_
	);
	LUT2 #(
		.INIT('h4)
	) name17935 (
		_w27256_,
		_w27818_,
		_w28448_
	);
	LUT2 #(
		.INIT('h4)
	) name17936 (
		_w27256_,
		_w27820_,
		_w28449_
	);
	LUT2 #(
		.INIT('h4)
	) name17937 (
		_w27256_,
		_w27823_,
		_w28450_
	);
	LUT2 #(
		.INIT('h4)
	) name17938 (
		_w27256_,
		_w27825_,
		_w28451_
	);
	LUT2 #(
		.INIT('h4)
	) name17939 (
		_w27256_,
		_w27827_,
		_w28452_
	);
	LUT2 #(
		.INIT('h4)
	) name17940 (
		_w27256_,
		_w27831_,
		_w28453_
	);
	LUT2 #(
		.INIT('h4)
	) name17941 (
		_w27256_,
		_w27833_,
		_w28454_
	);
	LUT2 #(
		.INIT('h4)
	) name17942 (
		_w27256_,
		_w27835_,
		_w28455_
	);
	LUT2 #(
		.INIT('h4)
	) name17943 (
		_w27256_,
		_w27837_,
		_w28456_
	);
	LUT2 #(
		.INIT('h4)
	) name17944 (
		_w27256_,
		_w27840_,
		_w28457_
	);
	LUT2 #(
		.INIT('h4)
	) name17945 (
		_w27256_,
		_w27842_,
		_w28458_
	);
	LUT2 #(
		.INIT('h4)
	) name17946 (
		_w27256_,
		_w27845_,
		_w28459_
	);
	LUT2 #(
		.INIT('h4)
	) name17947 (
		_w27256_,
		_w27847_,
		_w28460_
	);
	LUT2 #(
		.INIT('h4)
	) name17948 (
		_w27256_,
		_w27852_,
		_w28461_
	);
	LUT2 #(
		.INIT('h4)
	) name17949 (
		_w27256_,
		_w27854_,
		_w28462_
	);
	LUT2 #(
		.INIT('h4)
	) name17950 (
		_w27256_,
		_w27856_,
		_w28463_
	);
	LUT2 #(
		.INIT('h4)
	) name17951 (
		_w27256_,
		_w27858_,
		_w28464_
	);
	LUT2 #(
		.INIT('h4)
	) name17952 (
		_w27256_,
		_w27860_,
		_w28465_
	);
	LUT2 #(
		.INIT('h4)
	) name17953 (
		_w27256_,
		_w27862_,
		_w28466_
	);
	LUT2 #(
		.INIT('h4)
	) name17954 (
		_w27256_,
		_w27864_,
		_w28467_
	);
	LUT2 #(
		.INIT('h4)
	) name17955 (
		_w27256_,
		_w27867_,
		_w28468_
	);
	LUT2 #(
		.INIT('h4)
	) name17956 (
		_w27256_,
		_w27869_,
		_w28469_
	);
	LUT2 #(
		.INIT('h4)
	) name17957 (
		_w27256_,
		_w27871_,
		_w28470_
	);
	LUT2 #(
		.INIT('h4)
	) name17958 (
		_w27256_,
		_w27873_,
		_w28471_
	);
	LUT2 #(
		.INIT('h4)
	) name17959 (
		_w27256_,
		_w27875_,
		_w28472_
	);
	LUT2 #(
		.INIT('h4)
	) name17960 (
		_w27256_,
		_w27877_,
		_w28473_
	);
	LUT2 #(
		.INIT('h4)
	) name17961 (
		_w27256_,
		_w27879_,
		_w28474_
	);
	LUT2 #(
		.INIT('h4)
	) name17962 (
		_w27256_,
		_w27881_,
		_w28475_
	);
	LUT2 #(
		.INIT('h4)
	) name17963 (
		_w27256_,
		_w27883_,
		_w28476_
	);
	LUT2 #(
		.INIT('h4)
	) name17964 (
		_w27256_,
		_w27885_,
		_w28477_
	);
	LUT2 #(
		.INIT('h4)
	) name17965 (
		_w27256_,
		_w27887_,
		_w28478_
	);
	LUT2 #(
		.INIT('h4)
	) name17966 (
		_w27256_,
		_w27890_,
		_w28479_
	);
	LUT2 #(
		.INIT('h4)
	) name17967 (
		_w27256_,
		_w27892_,
		_w28480_
	);
	LUT2 #(
		.INIT('h4)
	) name17968 (
		_w27256_,
		_w27894_,
		_w28481_
	);
	LUT2 #(
		.INIT('h4)
	) name17969 (
		_w27256_,
		_w27896_,
		_w28482_
	);
	LUT2 #(
		.INIT('h4)
	) name17970 (
		_w27256_,
		_w27898_,
		_w28483_
	);
	LUT2 #(
		.INIT('h4)
	) name17971 (
		_w27256_,
		_w27900_,
		_w28484_
	);
	LUT2 #(
		.INIT('h4)
	) name17972 (
		_w27256_,
		_w27902_,
		_w28485_
	);
	LUT2 #(
		.INIT('h4)
	) name17973 (
		_w27256_,
		_w27904_,
		_w28486_
	);
	LUT2 #(
		.INIT('h4)
	) name17974 (
		_w27256_,
		_w27906_,
		_w28487_
	);
	LUT2 #(
		.INIT('h4)
	) name17975 (
		_w27256_,
		_w27908_,
		_w28488_
	);
	LUT2 #(
		.INIT('h4)
	) name17976 (
		_w27256_,
		_w27912_,
		_w28489_
	);
	LUT2 #(
		.INIT('h4)
	) name17977 (
		_w27256_,
		_w27914_,
		_w28490_
	);
	LUT2 #(
		.INIT('h4)
	) name17978 (
		_w27256_,
		_w27916_,
		_w28491_
	);
	LUT2 #(
		.INIT('h4)
	) name17979 (
		_w27256_,
		_w27918_,
		_w28492_
	);
	LUT2 #(
		.INIT('h4)
	) name17980 (
		_w27256_,
		_w27920_,
		_w28493_
	);
	LUT2 #(
		.INIT('h4)
	) name17981 (
		_w27256_,
		_w27923_,
		_w28494_
	);
	LUT2 #(
		.INIT('h4)
	) name17982 (
		_w27256_,
		_w27925_,
		_w28495_
	);
	LUT2 #(
		.INIT('h4)
	) name17983 (
		_w27256_,
		_w27927_,
		_w28496_
	);
	LUT2 #(
		.INIT('h4)
	) name17984 (
		_w27256_,
		_w27930_,
		_w28497_
	);
	LUT2 #(
		.INIT('h4)
	) name17985 (
		_w27256_,
		_w27932_,
		_w28498_
	);
	LUT2 #(
		.INIT('h4)
	) name17986 (
		_w27256_,
		_w27934_,
		_w28499_
	);
	LUT2 #(
		.INIT('h4)
	) name17987 (
		_w27256_,
		_w27937_,
		_w28500_
	);
	LUT2 #(
		.INIT('h4)
	) name17988 (
		_w27256_,
		_w27940_,
		_w28501_
	);
	LUT2 #(
		.INIT('h4)
	) name17989 (
		_w27256_,
		_w27942_,
		_w28502_
	);
	LUT2 #(
		.INIT('h4)
	) name17990 (
		_w27256_,
		_w27944_,
		_w28503_
	);
	LUT2 #(
		.INIT('h4)
	) name17991 (
		_w27256_,
		_w27946_,
		_w28504_
	);
	LUT2 #(
		.INIT('h4)
	) name17992 (
		_w27256_,
		_w27948_,
		_w28505_
	);
	LUT2 #(
		.INIT('h4)
	) name17993 (
		_w27256_,
		_w27950_,
		_w28506_
	);
	LUT2 #(
		.INIT('h4)
	) name17994 (
		_w27256_,
		_w27953_,
		_w28507_
	);
	LUT2 #(
		.INIT('h4)
	) name17995 (
		_w27256_,
		_w27957_,
		_w28508_
	);
	LUT2 #(
		.INIT('h4)
	) name17996 (
		_w27256_,
		_w27960_,
		_w28509_
	);
	LUT2 #(
		.INIT('h4)
	) name17997 (
		_w27256_,
		_w27962_,
		_w28510_
	);
	LUT2 #(
		.INIT('h4)
	) name17998 (
		_w27256_,
		_w27965_,
		_w28511_
	);
	LUT2 #(
		.INIT('h4)
	) name17999 (
		_w27256_,
		_w27967_,
		_w28512_
	);
	LUT2 #(
		.INIT('h4)
	) name18000 (
		_w27256_,
		_w27970_,
		_w28513_
	);
	LUT2 #(
		.INIT('h4)
	) name18001 (
		_w27256_,
		_w27972_,
		_w28514_
	);
	LUT2 #(
		.INIT('h4)
	) name18002 (
		_w27256_,
		_w27975_,
		_w28515_
	);
	LUT2 #(
		.INIT('h4)
	) name18003 (
		_w27256_,
		_w27977_,
		_w28516_
	);
	LUT2 #(
		.INIT('h4)
	) name18004 (
		_w27256_,
		_w27980_,
		_w28517_
	);
	LUT2 #(
		.INIT('h4)
	) name18005 (
		_w27256_,
		_w27982_,
		_w28518_
	);
	LUT2 #(
		.INIT('h4)
	) name18006 (
		_w27256_,
		_w27984_,
		_w28519_
	);
	LUT2 #(
		.INIT('h4)
	) name18007 (
		_w27256_,
		_w27986_,
		_w28520_
	);
	LUT2 #(
		.INIT('h4)
	) name18008 (
		_w27256_,
		_w27988_,
		_w28521_
	);
	LUT2 #(
		.INIT('h4)
	) name18009 (
		_w27256_,
		_w27991_,
		_w28522_
	);
	LUT2 #(
		.INIT('h4)
	) name18010 (
		_w27256_,
		_w27994_,
		_w28523_
	);
	LUT2 #(
		.INIT('h4)
	) name18011 (
		_w27256_,
		_w27996_,
		_w28524_
	);
	LUT2 #(
		.INIT('h4)
	) name18012 (
		_w27256_,
		_w27999_,
		_w28525_
	);
	LUT2 #(
		.INIT('h4)
	) name18013 (
		_w27256_,
		_w28001_,
		_w28526_
	);
	LUT2 #(
		.INIT('h4)
	) name18014 (
		_w27256_,
		_w28005_,
		_w28527_
	);
	LUT2 #(
		.INIT('h4)
	) name18015 (
		_w27256_,
		_w28007_,
		_w28528_
	);
	LUT2 #(
		.INIT('h4)
	) name18016 (
		_w27256_,
		_w28010_,
		_w28529_
	);
	LUT2 #(
		.INIT('h4)
	) name18017 (
		_w27256_,
		_w28012_,
		_w28530_
	);
	LUT2 #(
		.INIT('h4)
	) name18018 (
		_w27256_,
		_w28014_,
		_w28531_
	);
	LUT2 #(
		.INIT('h4)
	) name18019 (
		_w27256_,
		_w28016_,
		_w28532_
	);
	LUT2 #(
		.INIT('h4)
	) name18020 (
		_w27256_,
		_w28018_,
		_w28533_
	);
	LUT2 #(
		.INIT('h4)
	) name18021 (
		_w27256_,
		_w28021_,
		_w28534_
	);
	LUT2 #(
		.INIT('h4)
	) name18022 (
		_w27256_,
		_w28023_,
		_w28535_
	);
	LUT2 #(
		.INIT('h4)
	) name18023 (
		_w27256_,
		_w28026_,
		_w28536_
	);
	LUT2 #(
		.INIT('h4)
	) name18024 (
		_w27256_,
		_w28028_,
		_w28537_
	);
	LUT2 #(
		.INIT('h4)
	) name18025 (
		_w27256_,
		_w27754_,
		_w28538_
	);
	LUT2 #(
		.INIT('h4)
	) name18026 (
		_w27256_,
		_w28034_,
		_w28539_
	);
	LUT2 #(
		.INIT('h4)
	) name18027 (
		_w27256_,
		_w28036_,
		_w28540_
	);
	LUT2 #(
		.INIT('h4)
	) name18028 (
		_w27256_,
		_w28039_,
		_w28541_
	);
	LUT2 #(
		.INIT('h4)
	) name18029 (
		_w27256_,
		_w28041_,
		_w28542_
	);
	LUT2 #(
		.INIT('h4)
	) name18030 (
		_w27256_,
		_w28044_,
		_w28543_
	);
	LUT2 #(
		.INIT('h4)
	) name18031 (
		_w27256_,
		_w28047_,
		_w28544_
	);
	LUT2 #(
		.INIT('h4)
	) name18032 (
		_w27256_,
		_w28050_,
		_w28545_
	);
	LUT2 #(
		.INIT('h4)
	) name18033 (
		_w27256_,
		_w28053_,
		_w28546_
	);
	LUT2 #(
		.INIT('h4)
	) name18034 (
		_w27256_,
		_w28056_,
		_w28547_
	);
	LUT2 #(
		.INIT('h4)
	) name18035 (
		_w27256_,
		_w28059_,
		_w28548_
	);
	LUT2 #(
		.INIT('h4)
	) name18036 (
		_w27256_,
		_w28062_,
		_w28549_
	);
	LUT2 #(
		.INIT('h4)
	) name18037 (
		_w27256_,
		_w28064_,
		_w28550_
	);
	LUT2 #(
		.INIT('h4)
	) name18038 (
		_w27256_,
		_w28066_,
		_w28551_
	);
	LUT2 #(
		.INIT('h4)
	) name18039 (
		_w27256_,
		_w27850_,
		_w28552_
	);
	LUT2 #(
		.INIT('h4)
	) name18040 (
		_w27256_,
		_w28069_,
		_w28553_
	);
	LUT2 #(
		.INIT('h4)
	) name18041 (
		_w27256_,
		_w28072_,
		_w28554_
	);
	LUT2 #(
		.INIT('h4)
	) name18042 (
		_w27256_,
		_w28074_,
		_w28555_
	);
	LUT2 #(
		.INIT('h4)
	) name18043 (
		_w27256_,
		_w28077_,
		_w28556_
	);
	LUT2 #(
		.INIT('h4)
	) name18044 (
		_w27256_,
		_w28079_,
		_w28557_
	);
	LUT2 #(
		.INIT('h4)
	) name18045 (
		_w27256_,
		_w28082_,
		_w28558_
	);
	LUT2 #(
		.INIT('h4)
	) name18046 (
		_w27256_,
		_w28084_,
		_w28559_
	);
	LUT2 #(
		.INIT('h4)
	) name18047 (
		_w27256_,
		_w28087_,
		_w28560_
	);
	LUT2 #(
		.INIT('h4)
	) name18048 (
		_w27256_,
		_w28089_,
		_w28561_
	);
	LUT2 #(
		.INIT('h4)
	) name18049 (
		_w27256_,
		_w28092_,
		_w28562_
	);
	LUT2 #(
		.INIT('h4)
	) name18050 (
		_w27256_,
		_w28095_,
		_w28563_
	);
	LUT2 #(
		.INIT('h4)
	) name18051 (
		_w27256_,
		_w27955_,
		_w28564_
	);
	LUT2 #(
		.INIT('h4)
	) name18052 (
		_w27256_,
		_w28098_,
		_w28565_
	);
	LUT2 #(
		.INIT('h4)
	) name18053 (
		_w27256_,
		_w27910_,
		_w28566_
	);
	LUT2 #(
		.INIT('h4)
	) name18054 (
		_w27256_,
		_w28103_,
		_w28567_
	);
	LUT2 #(
		.INIT('h4)
	) name18055 (
		_w27256_,
		_w28108_,
		_w28568_
	);
	LUT2 #(
		.INIT('h4)
	) name18056 (
		_w27256_,
		_w28111_,
		_w28569_
	);
	LUT2 #(
		.INIT('h4)
	) name18057 (
		_w27256_,
		_w28114_,
		_w28570_
	);
	LUT2 #(
		.INIT('h4)
	) name18058 (
		_w27256_,
		_w28105_,
		_w28571_
	);
	LUT2 #(
		.INIT('h4)
	) name18059 (
		_w27256_,
		_w28119_,
		_w28572_
	);
	LUT2 #(
		.INIT('h4)
	) name18060 (
		_w27256_,
		_w28121_,
		_w28573_
	);
	LUT2 #(
		.INIT('h4)
	) name18061 (
		_w27256_,
		_w28123_,
		_w28574_
	);
	LUT3 #(
		.INIT('h6c)
	) name18062 (
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		_w11138_,
		_w28575_
	);
	LUT2 #(
		.INIT('h4)
	) name18063 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		_w11800_,
		_w28576_
	);
	LUT3 #(
		.INIT('h10)
	) name18064 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w28577_
	);
	LUT2 #(
		.INIT('h8)
	) name18065 (
		_w26978_,
		_w28577_,
		_w28578_
	);
	LUT3 #(
		.INIT('hf8)
	) name18066 (
		_w11797_,
		_w28576_,
		_w28578_,
		_w28579_
	);
	LUT3 #(
		.INIT('h80)
	) name18067 (
		\wishbone_TxBDReady_reg/NET0131 ,
		_w12314_,
		_w12316_,
		_w28580_
	);
	LUT2 #(
		.INIT('h8)
	) name18068 (
		_w12312_,
		_w28580_,
		_w28581_
	);
	LUT3 #(
		.INIT('h80)
	) name18069 (
		_w18757_,
		_w18758_,
		_w18765_,
		_w28582_
	);
	LUT2 #(
		.INIT('h8)
	) name18070 (
		_w24753_,
		_w28582_,
		_w28583_
	);
	LUT2 #(
		.INIT('h4)
	) name18071 (
		_w27096_,
		_w27097_,
		_w28584_
	);
	LUT3 #(
		.INIT('h13)
	) name18072 (
		_w11658_,
		_w11666_,
		_w27088_,
		_w28585_
	);
	LUT2 #(
		.INIT('hb)
	) name18073 (
		_w26971_,
		_w28585_,
		_w28586_
	);
	LUT2 #(
		.INIT('h8)
	) name18074 (
		_w18802_,
		_w24753_,
		_w28587_
	);
	LUT2 #(
		.INIT('h4)
	) name18075 (
		_w27096_,
		_w27101_,
		_w28588_
	);
	LUT2 #(
		.INIT('h8)
	) name18076 (
		_w18802_,
		_w27157_,
		_w28589_
	);
	LUT2 #(
		.INIT('h8)
	) name18077 (
		_w27157_,
		_w28582_,
		_w28590_
	);
	LUT2 #(
		.INIT('h8)
	) name18078 (
		_w18802_,
		_w26894_,
		_w28591_
	);
	LUT2 #(
		.INIT('h8)
	) name18079 (
		_w18755_,
		_w24753_,
		_w28592_
	);
	LUT2 #(
		.INIT('h8)
	) name18080 (
		_w24753_,
		_w26891_,
		_w28593_
	);
	LUT2 #(
		.INIT('h8)
	) name18081 (
		_w18755_,
		_w27157_,
		_w28594_
	);
	LUT2 #(
		.INIT('h8)
	) name18082 (
		_w26891_,
		_w27157_,
		_w28595_
	);
	LUT2 #(
		.INIT('h8)
	) name18083 (
		_w26894_,
		_w28582_,
		_w28596_
	);
	LUT2 #(
		.INIT('h8)
	) name18084 (
		_w18755_,
		_w26894_,
		_w28597_
	);
	LUT3 #(
		.INIT('h40)
	) name18085 (
		_w18750_,
		_w24752_,
		_w27186_,
		_w28598_
	);
	LUT2 #(
		.INIT('h8)
	) name18086 (
		_w18755_,
		_w28598_,
		_w28599_
	);
	LUT2 #(
		.INIT('h8)
	) name18087 (
		_w28582_,
		_w28598_,
		_w28600_
	);
	LUT3 #(
		.INIT('h80)
	) name18088 (
		_w18757_,
		_w18758_,
		_w18759_,
		_w28601_
	);
	LUT2 #(
		.INIT('h8)
	) name18089 (
		_w27157_,
		_w28601_,
		_w28602_
	);
	LUT2 #(
		.INIT('h8)
	) name18090 (
		_w26894_,
		_w28601_,
		_w28603_
	);
	LUT2 #(
		.INIT('h8)
	) name18091 (
		_w28598_,
		_w28601_,
		_w28604_
	);
	LUT2 #(
		.INIT('h8)
	) name18092 (
		_w24753_,
		_w28601_,
		_w28605_
	);
	LUT3 #(
		.INIT('h80)
	) name18093 (
		_w18757_,
		_w18759_,
		_w18762_,
		_w28606_
	);
	LUT2 #(
		.INIT('h8)
	) name18094 (
		_w24753_,
		_w28606_,
		_w28607_
	);
	LUT2 #(
		.INIT('h8)
	) name18095 (
		_w27157_,
		_w28606_,
		_w28608_
	);
	LUT2 #(
		.INIT('h8)
	) name18096 (
		_w26894_,
		_w28606_,
		_w28609_
	);
	LUT2 #(
		.INIT('h8)
	) name18097 (
		_w28598_,
		_w28606_,
		_w28610_
	);
	LUT3 #(
		.INIT('h10)
	) name18098 (
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w28611_
	);
	LUT4 #(
		.INIT('h1110)
	) name18099 (
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w28612_
	);
	LUT3 #(
		.INIT('h54)
	) name18100 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		_w28611_,
		_w28612_,
		_w28613_
	);
	LUT2 #(
		.INIT('hd)
	) name18101 (
		_w11004_,
		_w28613_,
		_w28614_
	);
	LUT2 #(
		.INIT('h8)
	) name18102 (
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		\txethmac1_random1_x_reg[7]/NET0131 ,
		_w28615_
	);
	LUT3 #(
		.INIT('hd0)
	) name18103 (
		\wishbone_RxBDRead_reg/NET0131 ,
		\wishbone_RxBDReady_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w28616_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name18104 (
		\wishbone_RxAbortSync3_reg/NET0131 ,
		\wishbone_RxAbortSync4_reg/NET0131 ,
		\wishbone_RxBDRead_reg/NET0131 ,
		\wishbone_RxBDReady_reg/NET0131 ,
		_w28617_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name18105 (
		_w25875_,
		_w25879_,
		_w28616_,
		_w28617_,
		_w28618_
	);
	LUT3 #(
		.INIT('h2a)
	) name18106 (
		\txethmac1_random1_RandomLatched_reg[2]/NET0131 ,
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w28619_
	);
	LUT2 #(
		.INIT('h1)
	) name18107 (
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w28620_
	);
	LUT4 #(
		.INIT('h0007)
	) name18108 (
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w28621_
	);
	LUT3 #(
		.INIT('h80)
	) name18109 (
		\txethmac1_random1_x_reg[2]/NET0131 ,
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w28622_
	);
	LUT3 #(
		.INIT('hba)
	) name18110 (
		_w28619_,
		_w28621_,
		_w28622_,
		_w28623_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name18111 (
		\wishbone_RxBDAddress_reg[1]/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w28624_
	);
	LUT4 #(
		.INIT('haba8)
	) name18112 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[0]/NET0131 ,
		_w25875_,
		_w25876_,
		_w28624_,
		_w28625_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name18113 (
		\wishbone_TxEn_needed_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w28626_
	);
	LUT2 #(
		.INIT('h4)
	) name18114 (
		\wishbone_WbEn_q_reg/NET0131 ,
		\wishbone_WbEn_reg/NET0131 ,
		_w28627_
	);
	LUT4 #(
		.INIT('h0200)
	) name18115 (
		\ethreg1_MODER_0_DataOut_reg[1]/NET0131 ,
		\wishbone_TxBDReady_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		\wishbone_WbEn_reg/NET0131 ,
		_w28628_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name18116 (
		_w26317_,
		_w26318_,
		_w28626_,
		_w28628_,
		_w28629_
	);
	LUT4 #(
		.INIT('h0008)
	) name18117 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28630_
	);
	LUT4 #(
		.INIT('h0008)
	) name18118 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28631_
	);
	LUT4 #(
		.INIT('h135f)
	) name18119 (
		_w26359_,
		_w26370_,
		_w28630_,
		_w28631_,
		_w28632_
	);
	LUT4 #(
		.INIT('h0200)
	) name18120 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w28633_
	);
	LUT4 #(
		.INIT('h0200)
	) name18121 (
		\ethreg1_TXCTRL_0_DataOut_reg[2]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28634_
	);
	LUT4 #(
		.INIT('h153f)
	) name18122 (
		_w25925_,
		_w26361_,
		_w28633_,
		_w28634_,
		_w28635_
	);
	LUT4 #(
		.INIT('h0020)
	) name18123 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28636_
	);
	LUT4 #(
		.INIT('h0200)
	) name18124 (
		\ethreg1_TXCTRL_1_DataOut_reg[2]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28637_
	);
	LUT4 #(
		.INIT('h153f)
	) name18125 (
		_w26365_,
		_w26370_,
		_w28636_,
		_w28637_,
		_w28638_
	);
	LUT4 #(
		.INIT('h0020)
	) name18126 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w28639_
	);
	LUT4 #(
		.INIT('h0020)
	) name18127 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28640_
	);
	LUT4 #(
		.INIT('h135f)
	) name18128 (
		_w26361_,
		_w26365_,
		_w28639_,
		_w28640_,
		_w28641_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18129 (
		_w28632_,
		_w28635_,
		_w28638_,
		_w28641_,
		_w28642_
	);
	LUT4 #(
		.INIT('h0008)
	) name18130 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28643_
	);
	LUT4 #(
		.INIT('h0008)
	) name18131 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28644_
	);
	LUT4 #(
		.INIT('h135f)
	) name18132 (
		_w26359_,
		_w26370_,
		_w28643_,
		_w28644_,
		_w28645_
	);
	LUT4 #(
		.INIT('h0200)
	) name18133 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w28646_
	);
	LUT4 #(
		.INIT('h0200)
	) name18134 (
		\ethreg1_TXCTRL_0_DataOut_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28647_
	);
	LUT4 #(
		.INIT('h153f)
	) name18135 (
		_w25925_,
		_w26361_,
		_w28646_,
		_w28647_,
		_w28648_
	);
	LUT4 #(
		.INIT('h0020)
	) name18136 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28649_
	);
	LUT4 #(
		.INIT('h0200)
	) name18137 (
		\ethreg1_TXCTRL_1_DataOut_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28650_
	);
	LUT4 #(
		.INIT('h153f)
	) name18138 (
		_w26365_,
		_w26370_,
		_w28649_,
		_w28650_,
		_w28651_
	);
	LUT4 #(
		.INIT('h0020)
	) name18139 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w28652_
	);
	LUT4 #(
		.INIT('h0020)
	) name18140 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28653_
	);
	LUT4 #(
		.INIT('h135f)
	) name18141 (
		_w26361_,
		_w26365_,
		_w28652_,
		_w28653_,
		_w28654_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18142 (
		_w28645_,
		_w28648_,
		_w28651_,
		_w28654_,
		_w28655_
	);
	LUT4 #(
		.INIT('h0008)
	) name18143 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28656_
	);
	LUT4 #(
		.INIT('h0008)
	) name18144 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28657_
	);
	LUT4 #(
		.INIT('h135f)
	) name18145 (
		_w26359_,
		_w26370_,
		_w28656_,
		_w28657_,
		_w28658_
	);
	LUT4 #(
		.INIT('h0200)
	) name18146 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w28659_
	);
	LUT4 #(
		.INIT('h0200)
	) name18147 (
		\ethreg1_TXCTRL_0_DataOut_reg[5]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28660_
	);
	LUT4 #(
		.INIT('h153f)
	) name18148 (
		_w25925_,
		_w26361_,
		_w28659_,
		_w28660_,
		_w28661_
	);
	LUT4 #(
		.INIT('h0020)
	) name18149 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28662_
	);
	LUT4 #(
		.INIT('h0200)
	) name18150 (
		\ethreg1_TXCTRL_1_DataOut_reg[5]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28663_
	);
	LUT4 #(
		.INIT('h153f)
	) name18151 (
		_w26365_,
		_w26370_,
		_w28662_,
		_w28663_,
		_w28664_
	);
	LUT4 #(
		.INIT('h0020)
	) name18152 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w28665_
	);
	LUT4 #(
		.INIT('h0020)
	) name18153 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28666_
	);
	LUT4 #(
		.INIT('h135f)
	) name18154 (
		_w26361_,
		_w26365_,
		_w28665_,
		_w28666_,
		_w28667_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18155 (
		_w28658_,
		_w28661_,
		_w28664_,
		_w28667_,
		_w28668_
	);
	LUT2 #(
		.INIT('h1)
	) name18156 (
		\wishbone_TxAbort_wb_reg/NET0131 ,
		\wishbone_TxDone_wb_reg/NET0131 ,
		_w28669_
	);
	LUT3 #(
		.INIT('h0e)
	) name18157 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		_w26321_,
		_w28669_,
		_w28670_
	);
	LUT4 #(
		.INIT('hf531)
	) name18158 (
		\Collision_Tx2_reg/NET0131 ,
		\ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		_w28671_
	);
	LUT4 #(
		.INIT('hf531)
	) name18159 (
		\ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		_w28672_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name18160 (
		\ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		_w28673_
	);
	LUT3 #(
		.INIT('h80)
	) name18161 (
		_w28671_,
		_w28672_,
		_w28673_,
		_w28674_
	);
	LUT2 #(
		.INIT('h4)
	) name18162 (
		\ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		_w28675_
	);
	LUT4 #(
		.INIT('haf23)
	) name18163 (
		\ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w28676_
	);
	LUT4 #(
		.INIT('h8caf)
	) name18164 (
		\ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w28677_
	);
	LUT4 #(
		.INIT('haf23)
	) name18165 (
		\ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		_w28678_
	);
	LUT4 #(
		.INIT('h4000)
	) name18166 (
		_w28675_,
		_w28676_,
		_w28677_,
		_w28678_,
		_w28679_
	);
	LUT3 #(
		.INIT('h01)
	) name18167 (
		\txethmac1_ColWindow_reg/NET0131 ,
		\txethmac1_txstatem1_StateIPG_reg/NET0131 ,
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		_w28680_
	);
	LUT4 #(
		.INIT('h00bf)
	) name18168 (
		_w13021_,
		_w28674_,
		_w28679_,
		_w28680_,
		_w28681_
	);
	LUT2 #(
		.INIT('h8)
	) name18169 (
		_w10533_,
		_w10536_,
		_w28682_
	);
	LUT4 #(
		.INIT('h0100)
	) name18170 (
		\txethmac1_txcrc_Crc_reg[30]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w28683_
	);
	LUT4 #(
		.INIT('hfefc)
	) name18171 (
		_w11026_,
		_w11028_,
		_w28683_,
		_w11027_,
		_w28684_
	);
	LUT3 #(
		.INIT('h12)
	) name18172 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131 ,
		wb_rst_i_pad,
		_w11279_,
		_w28685_
	);
	LUT3 #(
		.INIT('hd0)
	) name18173 (
		\ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131 ,
		_w28686_
	);
	LUT4 #(
		.INIT('h8000)
	) name18174 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxStatus_reg[14]/NET0131 ,
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w28687_
	);
	LUT4 #(
		.INIT('h0001)
	) name18175 (
		\wishbone_RxStatusInLatched_reg[3]/NET0131 ,
		\wishbone_RxStatusInLatched_reg[4]/NET0131 ,
		\wishbone_RxStatusInLatched_reg[5]/NET0131 ,
		\wishbone_RxStatusInLatched_reg[6]/NET0131 ,
		_w28688_
	);
	LUT2 #(
		.INIT('h1)
	) name18176 (
		\wishbone_RxStatusInLatched_reg[0]/NET0131 ,
		\wishbone_RxStatusInLatched_reg[1]/NET0131 ,
		_w28689_
	);
	LUT3 #(
		.INIT('h01)
	) name18177 (
		\macstatus1_LatchedCrcError_reg/NET0131 ,
		\wishbone_RxStatusInLatched_reg[0]/NET0131 ,
		\wishbone_RxStatusInLatched_reg[1]/NET0131 ,
		_w28690_
	);
	LUT4 #(
		.INIT('h4000)
	) name18178 (
		_w28686_,
		_w28687_,
		_w28688_,
		_w28690_,
		_w28691_
	);
	LUT4 #(
		.INIT('h0444)
	) name18179 (
		_w28686_,
		_w28687_,
		_w28688_,
		_w28689_,
		_w28692_
	);
	LUT4 #(
		.INIT('h4454)
	) name18180 (
		\miim1_EndBusy_reg/NET0131 ,
		\miim1_RStatStart_reg/NET0131 ,
		\miim1_RStat_q2_reg/NET0131 ,
		\miim1_RStat_q3_reg/NET0131 ,
		_w28693_
	);
	LUT4 #(
		.INIT('h0800)
	) name18181 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w28694_
	);
	LUT2 #(
		.INIT('h1)
	) name18182 (
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[1]/NET0131 ,
		_w28694_,
		_w28695_
	);
	LUT3 #(
		.INIT('h20)
	) name18183 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w28696_
	);
	LUT3 #(
		.INIT('h4c)
	) name18184 (
		_w25921_,
		_w25933_,
		_w28696_,
		_w28697_
	);
	LUT2 #(
		.INIT('h4)
	) name18185 (
		_w28695_,
		_w28697_,
		_w28698_
	);
	LUT3 #(
		.INIT('h10)
	) name18186 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w28699_
	);
	LUT2 #(
		.INIT('h8)
	) name18187 (
		_w25925_,
		_w28699_,
		_w28700_
	);
	LUT3 #(
		.INIT('hea)
	) name18188 (
		\maccontrol1_transmitcontrol1_ControlEnd_q_reg/P0001 ,
		_w25925_,
		_w28699_,
		_w28701_
	);
	LUT3 #(
		.INIT('h70)
	) name18189 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w28702_
	);
	LUT3 #(
		.INIT('h02)
	) name18190 (
		\wishbone_rx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[1]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[2]/NET0131 ,
		_w28703_
	);
	LUT2 #(
		.INIT('h2)
	) name18191 (
		\wishbone_ShiftEndedSync3_reg/NET0131 ,
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w28704_
	);
	LUT4 #(
		.INIT('h0008)
	) name18192 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[4]/NET0131 ,
		_w28705_
	);
	LUT4 #(
		.INIT('heaaa)
	) name18193 (
		_w28702_,
		_w28703_,
		_w28704_,
		_w28705_,
		_w28706_
	);
	LUT3 #(
		.INIT('h2a)
	) name18194 (
		\txethmac1_random1_RandomLatched_reg[4]/NET0131 ,
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w28707_
	);
	LUT4 #(
		.INIT('h001f)
	) name18195 (
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w28708_
	);
	LUT3 #(
		.INIT('h80)
	) name18196 (
		\txethmac1_random1_x_reg[4]/NET0131 ,
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w28709_
	);
	LUT3 #(
		.INIT('hba)
	) name18197 (
		_w28707_,
		_w28708_,
		_w28709_,
		_w28710_
	);
	LUT4 #(
		.INIT('h007f)
	) name18198 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxPointerRead_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w28711_
	);
	LUT3 #(
		.INIT('hd0)
	) name18199 (
		\ethreg1_MODER_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131 ,
		\wishbone_r_RxEn_q_reg/NET0131 ,
		_w28712_
	);
	LUT3 #(
		.INIT('h0d)
	) name18200 (
		\wishbone_RxAbortSync2_reg/NET0131 ,
		\wishbone_RxAbortSync3_reg/NET0131 ,
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w28713_
	);
	LUT3 #(
		.INIT('h10)
	) name18201 (
		_w28711_,
		_w28712_,
		_w28713_,
		_w28714_
	);
	LUT3 #(
		.INIT('h70)
	) name18202 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		\macstatus1_CarrierSenseLost_reg/NET0131 ,
		_w28715_
	);
	LUT4 #(
		.INIT('h0001)
	) name18203 (
		\CarrierSense_Tx2_reg/NET0131 ,
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		mcoll_pad_i_pad,
		_w28716_
	);
	LUT4 #(
		.INIT('h7350)
	) name18204 (
		_w10835_,
		_w10845_,
		_w28715_,
		_w28716_,
		_w28717_
	);
	LUT3 #(
		.INIT('h51)
	) name18205 (
		\wishbone_TxRetry_q_reg/NET0131 ,
		_w27064_,
		_w27065_,
		_w28718_
	);
	LUT2 #(
		.INIT('h4)
	) name18206 (
		\maccontrol1_MuxedDone_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w28719_
	);
	LUT4 #(
		.INIT('h0054)
	) name18207 (
		\maccontrol1_transmitcontrol1_BlockTxDone_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxDone_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w28720_
	);
	LUT2 #(
		.INIT('h4)
	) name18208 (
		_w28719_,
		_w28720_,
		_w28721_
	);
	LUT3 #(
		.INIT('hb4)
	) name18209 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		\wishbone_Flop_reg/NET0131 ,
		_w28722_
	);
	LUT3 #(
		.INIT('hb0)
	) name18210 (
		_w28719_,
		_w28720_,
		_w28722_,
		_w28723_
	);
	LUT2 #(
		.INIT('h8)
	) name18211 (
		_w28718_,
		_w28723_,
		_w28724_
	);
	LUT4 #(
		.INIT('h7f80)
	) name18212 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		_w28725_
	);
	LUT3 #(
		.INIT('h10)
	) name18213 (
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w28726_
	);
	LUT4 #(
		.INIT('h0100)
	) name18214 (
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w28727_
	);
	LUT3 #(
		.INIT('h54)
	) name18215 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		_w28726_,
		_w28727_,
		_w28728_
	);
	LUT2 #(
		.INIT('hd)
	) name18216 (
		_w11014_,
		_w28728_,
		_w28729_
	);
	LUT3 #(
		.INIT('h2a)
	) name18217 (
		\ethreg1_MODER_0_DataOut_reg[1]/NET0131 ,
		_w26317_,
		_w26318_,
		_w28730_
	);
	LUT2 #(
		.INIT('h4)
	) name18218 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		\wishbone_TxStatus_reg[14]/NET0131 ,
		_w28731_
	);
	LUT4 #(
		.INIT('h0001)
	) name18219 (
		\macstatus1_CarrierSenseLost_reg/NET0131 ,
		\macstatus1_LateCollLatched_reg/P0002 ,
		\macstatus1_RetryLimit_reg/P0002 ,
		\wishbone_TxUnderRun_reg/NET0131 ,
		_w28732_
	);
	LUT3 #(
		.INIT('h80)
	) name18220 (
		_w26321_,
		_w28731_,
		_w28732_,
		_w28733_
	);
	LUT3 #(
		.INIT('h08)
	) name18221 (
		_w26321_,
		_w28731_,
		_w28732_,
		_w28734_
	);
	LUT4 #(
		.INIT('h3133)
	) name18222 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w28735_
	);
	LUT3 #(
		.INIT('h02)
	) name18223 (
		_w25933_,
		_w28694_,
		_w28735_,
		_w28736_
	);
	LUT4 #(
		.INIT('h007f)
	) name18224 (
		\ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_Divider2_reg/NET0131 ,
		\maccontrol1_receivecontrol1_Pause_reg/NET0131 ,
		\maccontrol1_receivecontrol1_SlotTimer_reg[0]/NET0131 ,
		_w28737_
	);
	LUT3 #(
		.INIT('h01)
	) name18225 (
		wb_rst_i_pad,
		_w11279_,
		_w28737_,
		_w28738_
	);
	LUT3 #(
		.INIT('h51)
	) name18226 (
		\miim1_Nvalid_reg/NET0131 ,
		\miim1_ScanStat_q2_reg/NET0131 ,
		\miim1_SyncStatMdcEn_reg/NET0131 ,
		_w28739_
	);
	LUT2 #(
		.INIT('h4)
	) name18227 (
		\miim1_InProgress_q2_reg/NET0131 ,
		\miim1_InProgress_q3_reg/NET0131 ,
		_w28740_
	);
	LUT2 #(
		.INIT('h1)
	) name18228 (
		_w28739_,
		_w28740_,
		_w28741_
	);
	LUT2 #(
		.INIT('h2)
	) name18229 (
		\TxPauseRq_sync2_reg/NET0131 ,
		\TxPauseRq_sync3_reg/NET0131 ,
		_w28742_
	);
	LUT2 #(
		.INIT('h8)
	) name18230 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_TxUsedDataIn_q_reg/NET0131 ,
		_w28743_
	);
	LUT3 #(
		.INIT('h8c)
	) name18231 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w28744_
	);
	LUT4 #(
		.INIT('h0002)
	) name18232 (
		\maccontrol1_TxUsedDataOutDetected_reg/NET0131 ,
		\txethmac1_TxAbort_reg/NET0131 ,
		\txethmac1_TxDone_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w28745_
	);
	LUT4 #(
		.INIT('h2232)
	) name18233 (
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		_w28743_,
		_w28744_,
		_w28745_,
		_w28746_
	);
	LUT3 #(
		.INIT('ha2)
	) name18234 (
		\macstatus1_DeferLatched_reg/NET0131 ,
		\wishbone_BlockingTxStatusWrite_sync2_reg/NET0131 ,
		\wishbone_BlockingTxStatusWrite_sync3_reg/NET0131 ,
		_w28747_
	);
	LUT2 #(
		.INIT('he)
	) name18235 (
		_w10811_,
		_w28747_,
		_w28748_
	);
	LUT3 #(
		.INIT('h2a)
	) name18236 (
		\txethmac1_random1_RandomLatched_reg[3]/NET0131 ,
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w28749_
	);
	LUT3 #(
		.INIT('h80)
	) name18237 (
		\txethmac1_random1_x_reg[3]/NET0131 ,
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w28750_
	);
	LUT3 #(
		.INIT('hdc)
	) name18238 (
		_w28620_,
		_w28749_,
		_w28750_,
		_w28751_
	);
	LUT2 #(
		.INIT('h2)
	) name18239 (
		\wishbone_RxStatusWriteLatched_reg/NET0131 ,
		\wishbone_RxStatusWriteLatched_syncb2_reg/NET0131 ,
		_w28752_
	);
	LUT4 #(
		.INIT('h0800)
	) name18240 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxStatusWriteLatched_syncb2_reg/NET0131 ,
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w28753_
	);
	LUT2 #(
		.INIT('he)
	) name18241 (
		_w28752_,
		_w28753_,
		_w28754_
	);
	LUT4 #(
		.INIT('h4454)
	) name18242 (
		\miim1_EndBusy_reg/NET0131 ,
		\miim1_WCtrlDataStart_reg/NET0131 ,
		\miim1_WCtrlData_q2_reg/NET0131 ,
		\miim1_WCtrlData_q3_reg/NET0131 ,
		_w28755_
	);
	LUT3 #(
		.INIT('h01)
	) name18243 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[2]/NET0131 ,
		\ethreg1_MIIADDRESS_1_DataOut_reg[3]/NET0131 ,
		\ethreg1_MIIADDRESS_1_DataOut_reg[4]/NET0131 ,
		_w28756_
	);
	LUT2 #(
		.INIT('h2)
	) name18244 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[0]/NET0131 ,
		\ethreg1_MIIADDRESS_1_DataOut_reg[1]/NET0131 ,
		_w28757_
	);
	LUT4 #(
		.INIT('h3aaa)
	) name18245 (
		\miim1_shftrg_LinkFail_reg/NET0131 ,
		\miim1_shftrg_ShiftReg_reg[1]/NET0131 ,
		_w28756_,
		_w28757_,
		_w28758_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name18246 (
		\wishbone_RxEn_needed_reg/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w28759_
	);
	LUT3 #(
		.INIT('h02)
	) name18247 (
		\ethreg1_MODER_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w28760_
	);
	LUT3 #(
		.INIT('hec)
	) name18248 (
		_w28627_,
		_w28759_,
		_w28760_,
		_w28761_
	);
	LUT3 #(
		.INIT('h20)
	) name18249 (
		wb_cyc_i_pad,
		wb_err_o_pad,
		wb_stb_i_pad,
		_w28762_
	);
	LUT3 #(
		.INIT('he0)
	) name18250 (
		\wb_adr_i[11]_pad ,
		_w18750_,
		_w28762_,
		_w28763_
	);
	LUT2 #(
		.INIT('h2)
	) name18251 (
		\maccontrol1_MuxedDone_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w28764_
	);
	LUT4 #(
		.INIT('h0040)
	) name18252 (
		\maccontrol1_TxDoneInLatched_reg/NET0131 ,
		\maccontrol1_TxUsedDataOutDetected_reg/NET0131 ,
		\txethmac1_TxDone_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w28765_
	);
	LUT2 #(
		.INIT('he)
	) name18253 (
		_w28764_,
		_w28765_,
		_w28766_
	);
	LUT2 #(
		.INIT('h2)
	) name18254 (
		\maccontrol1_MuxedAbort_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w28767_
	);
	LUT4 #(
		.INIT('h0040)
	) name18255 (
		\maccontrol1_TxAbortInLatched_reg/NET0131 ,
		\maccontrol1_TxUsedDataOutDetected_reg/NET0131 ,
		\txethmac1_TxAbort_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w28768_
	);
	LUT2 #(
		.INIT('he)
	) name18256 (
		_w28767_,
		_w28768_,
		_w28769_
	);
	LUT2 #(
		.INIT('h4)
	) name18257 (
		_w27096_,
		_w27242_,
		_w28770_
	);
	LUT2 #(
		.INIT('h2)
	) name18258 (
		\ethreg1_SetTxCIrq_sync2_reg/NET0131 ,
		\ethreg1_SetTxCIrq_sync3_reg/NET0131 ,
		_w28771_
	);
	LUT2 #(
		.INIT('h2)
	) name18259 (
		\ethreg1_SetRxCIrq_sync2_reg/NET0131 ,
		\ethreg1_SetRxCIrq_sync3_reg/NET0131 ,
		_w28772_
	);
	LUT3 #(
		.INIT('h20)
	) name18260 (
		\wishbone_BDRead_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		\wishbone_WbEn_reg/NET0131 ,
		_w28773_
	);
	LUT4 #(
		.INIT('h0001)
	) name18261 (
		\wishbone_BDWrite_reg[0]/NET0131 ,
		\wishbone_BDWrite_reg[1]/NET0131 ,
		\wishbone_BDWrite_reg[2]/NET0131 ,
		\wishbone_BDWrite_reg[3]/NET0131 ,
		_w28774_
	);
	LUT3 #(
		.INIT('hce)
	) name18262 (
		_w27254_,
		_w28773_,
		_w28774_,
		_w28775_
	);
	LUT3 #(
		.INIT('h02)
	) name18263 (
		\maccontrol1_TxUsedDataOutDetected_reg/NET0131 ,
		\txethmac1_TxAbort_reg/NET0131 ,
		\txethmac1_TxDone_reg/NET0131 ,
		_w28776_
	);
	LUT2 #(
		.INIT('h2)
	) name18264 (
		_w10836_,
		_w28776_,
		_w28777_
	);
	LUT2 #(
		.INIT('h2)
	) name18265 (
		\WillSendControlFrame_sync2_reg/NET0131 ,
		\WillSendControlFrame_sync3_reg/NET0131 ,
		_w28778_
	);
	LUT3 #(
		.INIT('h2a)
	) name18266 (
		\txethmac1_random1_RandomLatched_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w28779_
	);
	LUT3 #(
		.INIT('h01)
	) name18267 (
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w28780_
	);
	LUT3 #(
		.INIT('h80)
	) name18268 (
		\txethmac1_random1_x_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w28781_
	);
	LUT3 #(
		.INIT('hba)
	) name18269 (
		_w28779_,
		_w28780_,
		_w28781_,
		_w28782_
	);
	LUT4 #(
		.INIT('h4500)
	) name18270 (
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\ethreg1_MODER_2_DataOut_reg[0]/NET0131 ,
		\macstatus1_RxColWindow_reg/NET0131 ,
		mcoll_pad_i_pad,
		_w28783_
	);
	LUT3 #(
		.INIT('h54)
	) name18271 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		\macstatus1_RxLateCollision_reg/NET0131 ,
		_w28783_,
		_w28784_
	);
	LUT2 #(
		.INIT('h1)
	) name18272 (
		\Collision_Tx1_reg/NET0131 ,
		\Collision_Tx2_reg/NET0131 ,
		_w28785_
	);
	LUT3 #(
		.INIT('h07)
	) name18273 (
		_w10827_,
		_w10845_,
		_w28785_,
		_w28786_
	);
	LUT3 #(
		.INIT('h70)
	) name18274 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w28787_
	);
	LUT2 #(
		.INIT('h8)
	) name18275 (
		\wishbone_RxBDRead_reg/NET0131 ,
		\wishbone_RxBDReady_reg/NET0131 ,
		_w28788_
	);
	LUT2 #(
		.INIT('he)
	) name18276 (
		_w28787_,
		_w28788_,
		_w28789_
	);
	LUT3 #(
		.INIT('h45)
	) name18277 (
		\maccontrol1_TxUsedDataOutDetected_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w28790_
	);
	LUT2 #(
		.INIT('h2)
	) name18278 (
		_w25932_,
		_w28790_,
		_w28791_
	);
	LUT4 #(
		.INIT('h22f2)
	) name18279 (
		\wishbone_ShiftEndedSync1_reg/NET0131 ,
		\wishbone_ShiftEndedSync2_reg/NET0131 ,
		\wishbone_ShiftEndedSync3_reg/NET0131 ,
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w28792_
	);
	LUT3 #(
		.INIT('h01)
	) name18280 (
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\txethmac1_txstatem1_Rule1_reg/NET0131 ,
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w28793_
	);
	LUT2 #(
		.INIT('h1)
	) name18281 (
		\txethmac1_txstatem1_StateBackOff_reg/NET0131 ,
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		_w28794_
	);
	LUT2 #(
		.INIT('h4)
	) name18282 (
		_w28793_,
		_w28794_,
		_w28795_
	);
	LUT4 #(
		.INIT('hee0e)
	) name18283 (
		\wishbone_TxRetryPacketBlocked_reg/NET0131 ,
		\wishbone_TxRetryPacket_reg/NET0131 ,
		\wishbone_TxRetry_wb_q_reg/NET0131 ,
		\wishbone_TxRetry_wb_reg/NET0131 ,
		_w28796_
	);
	LUT3 #(
		.INIT('h0e)
	) name18284 (
		\RxAbort_wb_reg/NET0131 ,
		\wishbone_RxAbortLatched_reg/NET0131 ,
		\wishbone_RxAbortSyncb2_reg/NET0131 ,
		_w28797_
	);
	LUT4 #(
		.INIT('h8ace)
	) name18285 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131 ,
		\txethmac1_TxDone_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w28798_
	);
	LUT4 #(
		.INIT('h8f88)
	) name18286 (
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxBDReady_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w28799_
	);
	LUT4 #(
		.INIT('haa0c)
	) name18287 (
		\RxEnSync_reg/NET0131 ,
		\ethreg1_MODER_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131 ,
		mrxdv_pad_i_pad,
		_w28800_
	);
	LUT4 #(
		.INIT('h1110)
	) name18288 (
		m_wb_ack_i_pad,
		m_wb_err_i_pad,
		\wishbone_BlockingIncrementTxPointer_reg/NET0131 ,
		\wishbone_IncrTxPointer_reg/NET0131 ,
		_w28801_
	);
	LUT3 #(
		.INIT('hf4)
	) name18289 (
		\wishbone_BlockingTxStatusWrite_sync2_reg/NET0131 ,
		\wishbone_TxUnderRun_sync1_reg/NET0131 ,
		\wishbone_TxUnderRun_wb_reg/NET0131 ,
		_w28802_
	);
	LUT2 #(
		.INIT('h2)
	) name18290 (
		\miim1_EndBusy_reg/NET0131 ,
		\miim1_WCtrlDataStart_q_reg/NET0131 ,
		_w28803_
	);
	LUT3 #(
		.INIT('hd8)
	) name18291 (
		\miim1_EndBusy_reg/NET0131 ,
		\miim1_WCtrlDataStart_q_reg/NET0131 ,
		\miim1_WCtrlDataStart_reg/NET0131 ,
		_w28804_
	);
	LUT3 #(
		.INIT('hce)
	) name18292 (
		\maccontrol1_transmitcontrol1_BlockTxDone_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w28805_
	);
	LUT3 #(
		.INIT('h54)
	) name18293 (
		\wishbone_BlockingTxStatusWrite_sync2_reg/NET0131 ,
		\wishbone_TxUnderRun_reg/NET0131 ,
		\wishbone_TxUnderRun_sync1_reg/NET0131 ,
		_w28806_
	);
	LUT4 #(
		.INIT('hc0ea)
	) name18294 (
		\maccontrol1_transmitcontrol1_SendingCtrlFrm_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131 ,
		\txethmac1_TxDone_reg/NET0131 ,
		_w28807_
	);
	LUT2 #(
		.INIT('he)
	) name18295 (
		\miim1_outctrl_Mdo_2d_reg/NET0131 ,
		\miim1_shftrg_ShiftReg_reg[7]/NET0131 ,
		_w28808_
	);
	LUT2 #(
		.INIT('h8)
	) name18296 (
		\ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_TXCTRL_2_DataOut_reg[0]/NET0131 ,
		_w28809_
	);
	LUT3 #(
		.INIT('hea)
	) name18297 (
		wb_rst_i_pad,
		_w13016_,
		_w13397_,
		_w28810_
	);
	LUT3 #(
		.INIT('hea)
	) name18298 (
		wb_rst_i_pad,
		_w14512_,
		_w14872_,
		_w28811_
	);
	LUT4 #(
		.INIT('h0111)
	) name18299 (
		wb_rst_i_pad,
		_w15775_,
		_w16122_,
		_w16814_,
		_w28812_
	);
	LUT3 #(
		.INIT('hea)
	) name18300 (
		wb_rst_i_pad,
		_w12301_,
		_w12668_,
		_w28813_
	);
	LUT4 #(
		.INIT('h0800)
	) name18301 (
		_w28810_,
		_w28811_,
		_w28812_,
		_w28813_,
		_w28814_
	);
	LUT4 #(
		.INIT('heaaa)
	) name18302 (
		wb_rst_i_pad,
		_w18058_,
		_w18401_,
		_w18746_,
		_w28815_
	);
	LUT3 #(
		.INIT('hea)
	) name18303 (
		wb_rst_i_pad,
		_w15222_,
		_w16469_,
		_w28816_
	);
	LUT3 #(
		.INIT('hea)
	) name18304 (
		wb_rst_i_pad,
		_w17356_,
		_w17713_,
		_w28817_
	);
	LUT3 #(
		.INIT('h80)
	) name18305 (
		_w28815_,
		_w28816_,
		_w28817_,
		_w28818_
	);
	LUT2 #(
		.INIT('h2)
	) name18306 (
		_w12303_,
		_w13800_,
		_w28819_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name18307 (
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxBDReady_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w28820_
	);
	LUT3 #(
		.INIT('h20)
	) name18308 (
		_w25940_,
		_w25941_,
		_w28820_,
		_w28821_
	);
	LUT4 #(
		.INIT('hff70)
	) name18309 (
		_w28814_,
		_w28818_,
		_w28819_,
		_w28821_,
		_w28822_
	);
	LUT2 #(
		.INIT('h1)
	) name18310 (
		wb_rst_i_pad,
		_w23950_,
		_w28823_
	);
	LUT2 #(
		.INIT('h1)
	) name18311 (
		wb_rst_i_pad,
		_w23589_,
		_w28824_
	);
	LUT2 #(
		.INIT('h1)
	) name18312 (
		wb_rst_i_pad,
		_w22213_,
		_w28825_
	);
	LUT4 #(
		.INIT('h070f)
	) name18313 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w28826_
	);
	LUT3 #(
		.INIT('h02)
	) name18314 (
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		_w13807_,
		_w13809_,
		_w28827_
	);
	LUT3 #(
		.INIT('h01)
	) name18315 (
		wb_rst_i_pad,
		_w13809_,
		_w28826_,
		_w28828_
	);
	LUT3 #(
		.INIT('hdc)
	) name18316 (
		_w19524_,
		_w28827_,
		_w28828_,
		_w28829_
	);
	LUT2 #(
		.INIT('h1)
	) name18317 (
		wb_rst_i_pad,
		_w19149_,
		_w28830_
	);
	LUT4 #(
		.INIT('h0002)
	) name18318 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w28831_
	);
	LUT3 #(
		.INIT('h80)
	) name18319 (
		_w18757_,
		_w18762_,
		_w28831_,
		_w28832_
	);
	LUT3 #(
		.INIT('h80)
	) name18320 (
		\ethreg1_MIIRX_DATA_DataOut_reg[10]/NET0131 ,
		_w18785_,
		_w18786_,
		_w28833_
	);
	LUT4 #(
		.INIT('h0008)
	) name18321 (
		\ethreg1_RXHASH0_1_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w28834_
	);
	LUT3 #(
		.INIT('h80)
	) name18322 (
		_w18757_,
		_w18758_,
		_w28834_,
		_w28835_
	);
	LUT4 #(
		.INIT('h0008)
	) name18323 (
		\ethreg1_RXHASH1_1_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w28836_
	);
	LUT3 #(
		.INIT('h80)
	) name18324 (
		_w18757_,
		_w18762_,
		_w28836_,
		_w28837_
	);
	LUT4 #(
		.INIT('h0001)
	) name18325 (
		_w28832_,
		_w28833_,
		_w28835_,
		_w28837_,
		_w28838_
	);
	LUT4 #(
		.INIT('h0002)
	) name18326 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w28839_
	);
	LUT4 #(
		.INIT('h0020)
	) name18327 (
		\ethreg1_TXCTRL_1_DataOut_reg[2]/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w28840_
	);
	LUT4 #(
		.INIT('h777f)
	) name18328 (
		_w18757_,
		_w18758_,
		_w28839_,
		_w28840_,
		_w28841_
	);
	LUT2 #(
		.INIT('h8)
	) name18329 (
		_w18752_,
		_w28841_,
		_w28842_
	);
	LUT3 #(
		.INIT('h80)
	) name18330 (
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		_w18800_,
		_w18801_,
		_w28843_
	);
	LUT3 #(
		.INIT('h80)
	) name18331 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[2]/NET0131 ,
		_w18785_,
		_w18798_,
		_w28844_
	);
	LUT3 #(
		.INIT('h80)
	) name18332 (
		\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 ,
		_w18753_,
		_w18754_,
		_w28845_
	);
	LUT3 #(
		.INIT('h80)
	) name18333 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[2]/NET0131 ,
		_w18798_,
		_w18805_,
		_w28846_
	);
	LUT4 #(
		.INIT('h0001)
	) name18334 (
		_w28843_,
		_w28844_,
		_w28845_,
		_w28846_,
		_w28847_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name18335 (
		_w18752_,
		_w28838_,
		_w28841_,
		_w28847_,
		_w28848_
	);
	LUT4 #(
		.INIT('h1555)
	) name18336 (
		wb_rst_i_pad,
		_w28838_,
		_w28842_,
		_w28847_,
		_w28849_
	);
	LUT3 #(
		.INIT('hdc)
	) name18337 (
		_w24382_,
		_w28848_,
		_w28849_,
		_w28850_
	);
	LUT4 #(
		.INIT('h1555)
	) name18338 (
		\wishbone_RxPointerMSB_reg[10]/NET0131 ,
		_w15283_,
		_w15284_,
		_w23169_,
		_w28851_
	);
	LUT4 #(
		.INIT('h1555)
	) name18339 (
		_w13807_,
		_w15283_,
		_w15284_,
		_w15285_,
		_w28852_
	);
	LUT2 #(
		.INIT('h4)
	) name18340 (
		_w28851_,
		_w28852_,
		_w28853_
	);
	LUT3 #(
		.INIT('hf2)
	) name18341 (
		_w15282_,
		_w24382_,
		_w28853_,
		_w28854_
	);
	LUT2 #(
		.INIT('h8)
	) name18342 (
		\ethreg1_INT_MASK_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_irq_rxe_reg/NET0131 ,
		_w28855_
	);
	LUT4 #(
		.INIT('h135f)
	) name18343 (
		\ethreg1_INT_MASK_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_INT_MASK_0_DataOut_reg[6]/NET0131 ,
		\ethreg1_irq_rxb_reg/NET0131 ,
		\ethreg1_irq_rxc_reg/NET0131 ,
		_w28856_
	);
	LUT4 #(
		.INIT('h135f)
	) name18344 (
		\ethreg1_INT_MASK_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_INT_MASK_0_DataOut_reg[5]/NET0131 ,
		\ethreg1_irq_busy_reg/NET0131 ,
		\ethreg1_irq_txc_reg/NET0131 ,
		_w28857_
	);
	LUT4 #(
		.INIT('h135f)
	) name18345 (
		\ethreg1_INT_MASK_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_INT_MASK_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_irq_txb_reg/NET0131 ,
		\ethreg1_irq_txe_reg/NET0131 ,
		_w28858_
	);
	LUT4 #(
		.INIT('hbfff)
	) name18346 (
		_w28855_,
		_w28856_,
		_w28857_,
		_w28858_,
		_w28859_
	);
	LUT4 #(
		.INIT('haccc)
	) name18347 (
		\m_wb_dat_i[15]_pad ,
		\wishbone_tx_fifo_fifo_reg[2][15]/P0001 ,
		_w26076_,
		_w26088_,
		_w28860_
	);
	LUT4 #(
		.INIT('haccc)
	) name18348 (
		\m_wb_dat_i[16]_pad ,
		\wishbone_tx_fifo_fifo_reg[2][16]/P0001 ,
		_w26076_,
		_w26088_,
		_w28861_
	);
	LUT4 #(
		.INIT('haccc)
	) name18349 (
		\m_wb_dat_i[17]_pad ,
		\wishbone_tx_fifo_fifo_reg[2][17]/P0001 ,
		_w26076_,
		_w26088_,
		_w28862_
	);
	LUT4 #(
		.INIT('haccc)
	) name18350 (
		\m_wb_dat_i[22]_pad ,
		\wishbone_tx_fifo_fifo_reg[2][22]/P0001 ,
		_w26076_,
		_w26088_,
		_w28863_
	);
	LUT4 #(
		.INIT('haccc)
	) name18351 (
		\m_wb_dat_i[23]_pad ,
		\wishbone_tx_fifo_fifo_reg[2][23]/P0001 ,
		_w26076_,
		_w26088_,
		_w28864_
	);
	LUT4 #(
		.INIT('haccc)
	) name18352 (
		\m_wb_dat_i[25]_pad ,
		\wishbone_tx_fifo_fifo_reg[2][25]/P0001 ,
		_w26076_,
		_w26088_,
		_w28865_
	);
	LUT4 #(
		.INIT('haccc)
	) name18353 (
		\m_wb_dat_i[2]_pad ,
		\wishbone_tx_fifo_fifo_reg[2][2]/P0001 ,
		_w26076_,
		_w26088_,
		_w28866_
	);
	assign \_al_n1  = 1'b1;
	assign \g215539/_0_  = _w10532_ ;
	assign \g215543/_0_  = _w10541_ ;
	assign \g215547/_0_  = _w10545_ ;
	assign \g215551/_0_  = _w10587_ ;
	assign \g215552/_0_  = _w10596_ ;
	assign \g215578/_0_  = _w10599_ ;
	assign \g215587/_1_  = _w10852_ ;
	assign \g215589/_1_  = _w10859_ ;
	assign \g215591/_1_  = _w10864_ ;
	assign \g215593/_1_  = _w10866_ ;
	assign \g215595/_1_  = _w10868_ ;
	assign \g215597/_1_  = _w10872_ ;
	assign \g215599/_1_  = _w10876_ ;
	assign \g215601/_1_  = _w10881_ ;
	assign \g215603/_1_  = _w10887_ ;
	assign \g215605/_1_  = _w10893_ ;
	assign \g215607/_1_  = _w10900_ ;
	assign \g215609/_1_  = _w10904_ ;
	assign \g215611/_1_  = _w10906_ ;
	assign \g215613/_1_  = _w10908_ ;
	assign \g215615/_1_  = _w10910_ ;
	assign \g215617/_1_  = _w10912_ ;
	assign \g215618/_0_  = _w10916_ ;
	assign \g215619/_0_  = _w10918_ ;
	assign \g215620/_0_  = _w10940_ ;
	assign \g215632/_1_  = _w10942_ ;
	assign \g215634/_0_  = _w10952_ ;
	assign \g215635/_0_  = _w10959_ ;
	assign \g215636/_0_  = _w10961_ ;
	assign \g215637/_0_  = _w10963_ ;
	assign \g215638/_0_  = _w10969_ ;
	assign \g215639/_0_  = _w10974_ ;
	assign \g215655/_1_  = _w10984_ ;
	assign \g215657/_1_  = _w10988_ ;
	assign \g215659/_1_  = _w10993_ ;
	assign \g215661/_1_  = _w10995_ ;
	assign \g215662/_0_  = _w11010_ ;
	assign \g215663/_0_  = _w11025_ ;
	assign \g215664/_0_  = _w11039_ ;
	assign \g215665/_0_  = _w11042_ ;
	assign \g215668/_0_  = _w11044_ ;
	assign \g215674/_0_  = _w11050_ ;
	assign \g215677/_0_  = _w11061_ ;
	assign \g215686/_0_  = _w11071_ ;
	assign \g215695/_0_  = _w11076_ ;
	assign \g215696/_0_  = _w11080_ ;
	assign \g215702/_1__syn_2  = _w11071_ ;
	assign \g215705/_0_  = _w11086_ ;
	assign \g215706/_0_  = _w11088_ ;
	assign \g215716/_0_  = _w11099_ ;
	assign \g215717/_0_  = _w11104_ ;
	assign \g215718/_0_  = _w11112_ ;
	assign \g215726/_0_  = _w11118_ ;
	assign \g215727/_0_  = _w11123_ ;
	assign \g215728/_0_  = _w11127_ ;
	assign \g215760/_0_  = _w11132_ ;
	assign \g215764/_0_  = _w11270_ ;
	assign \g215765/_0_  = _w11291_ ;
	assign \g215766/_0_  = _w11296_ ;
	assign \g215767/_3_  = _w11304_ ;
	assign \g215768/_3_  = _w11310_ ;
	assign \g215769/_3_  = _w11317_ ;
	assign \g215770/_3_  = _w11322_ ;
	assign \g215771/_3_  = _w11326_ ;
	assign \g215772/_3_  = _w11330_ ;
	assign \g215773/_3_  = _w11334_ ;
	assign \g215774/_3_  = _w11338_ ;
	assign \g215775/_3_  = _w11344_ ;
	assign \g215776/_3_  = _w11348_ ;
	assign \g215777/_3_  = _w11352_ ;
	assign \g215778/_3_  = _w11356_ ;
	assign \g215779/_3_  = _w11361_ ;
	assign \g215780/_3_  = _w11365_ ;
	assign \g215790/_0_  = _w11369_ ;
	assign \g215791/_0_  = _w11376_ ;
	assign \g215792/_0_  = _w11383_ ;
	assign \g215793/_0_  = _w11385_ ;
	assign \g215801/_0_  = _w11396_ ;
	assign \g215802/_0_  = _w11399_ ;
	assign \g215803/_0_  = _w11404_ ;
	assign \g215804/_0_  = _w11406_ ;
	assign \g215812/_0_  = _w11410_ ;
	assign \g215813/_0_  = _w11417_ ;
	assign \g215821/_0_  = _w11421_ ;
	assign \g215823/_0_  = _w11428_ ;
	assign \g215831/_0_  = _w11432_ ;
	assign \g215832/_0_  = _w11435_ ;
	assign \g215833/_0_  = _w11442_ ;
	assign \g215845/_0_  = _w11448_ ;
	assign \g215846/_0_  = _w11449_ ;
	assign \g215847/_0_  = _w11541_ ;
	assign \g215872/_0_  = _w11546_ ;
	assign \g215873/_0_  = _w11568_ ;
	assign \g215874/_0_  = _w11572_ ;
	assign \g215904/_0_  = _w11575_ ;
	assign \g215905/_0_  = _w11589_ ;
	assign \g215906/_0_  = _w11595_ ;
	assign \g215907/_0_  = _w11596_ ;
	assign \g215908/_0_  = _w11599_ ;
	assign \g215909/_0_  = _w11602_ ;
	assign \g215910/_0_  = _w11607_ ;
	assign \g215911/_0_  = _w11608_ ;
	assign \g215912/_0_  = _w11609_ ;
	assign \g215913/_0_  = _w11611_ ;
	assign \g215914/_0_  = _w11613_ ;
	assign \g215915/_0_  = _w11617_ ;
	assign \g215916/_0_  = _w11622_ ;
	assign \g215917/_0_  = _w11623_ ;
	assign \g215918/_0_  = _w11626_ ;
	assign \g215919/_0_  = _w11629_ ;
	assign \g215920/_0_  = _w11630_ ;
	assign \g215923/_0_  = _w11634_ ;
	assign \g215926/_0_  = _w11637_ ;
	assign \g215941/_0_  = _w11645_ ;
	assign \g215942/_0_  = _w11647_ ;
	assign \g215943/_0_  = _w11650_ ;
	assign \g215944/_0_  = _w11654_ ;
	assign \g215945/_0_  = _w11673_ ;
	assign \g215946/_0_  = _w11686_ ;
	assign \g215947/_0_  = _w11699_ ;
	assign \g215948/_0_  = _w11712_ ;
	assign \g215949/_0_  = _w11725_ ;
	assign \g215950/_0_  = _w11738_ ;
	assign \g215951/_0_  = _w11751_ ;
	assign \g215952/_0_  = _w11764_ ;
	assign \g215953/_0_  = _w11765_ ;
	assign \g215954/_0_  = _w11770_ ;
	assign \g215955/_0_  = _w11772_ ;
	assign \g215956/_0_  = _w11783_ ;
	assign \g215957/_0_  = _w11794_ ;
	assign \g215959/_00_  = _w11807_ ;
	assign \g215960/_0_  = _w11810_ ;
	assign \g215962/_0_  = _w11813_ ;
	assign \g215964/_0_  = _w11837_ ;
	assign \g215966/_0_  = _w11840_ ;
	assign \g215972/_0_  = _w11844_ ;
	assign \g216035/_0_  = _w11918_ ;
	assign \g216037/_0_  = _w11928_ ;
	assign \g216038/_0_  = _w12327_ ;
	assign \g216039/_0_  = _w12675_ ;
	assign \g216040/_0_  = _w13018_ ;
	assign \g216041/_0_  = _w13019_ ;
	assign \g216042/_0_  = _w13020_ ;
	assign \g216046/_0_  = _w13045_ ;
	assign \g216048/_0_  = _w13056_ ;
	assign \g216057/_0_  = _w13405_ ;
	assign \g216263/_0_  = _w13418_ ;
	assign \g216264/_0_  = _w13431_ ;
	assign \g216265/_0_  = _w13435_ ;
	assign \g216266/_0_  = _w13439_ ;
	assign \g216267/_0_  = _w13443_ ;
	assign \g216268/_0_  = _w13447_ ;
	assign \g216269/_0_  = _w13451_ ;
	assign \g216270/_0_  = _w13455_ ;
	assign \g216271/_0_  = _w13802_ ;
	assign \g216272/_0_  = _w13806_ ;
	assign \g216273/_0_  = _w14153_ ;
	assign \g216284/_0_  = _w14157_ ;
	assign \g216289/_0_  = _w14160_ ;
	assign \g216290/_0_  = _w14171_ ;
	assign \g216292/_0_  = _w14531_ ;
	assign \g216296/_0_  = _w14881_ ;
	assign \g216297/_0_  = _w15233_ ;
	assign \g216300/_0_  = _w15239_ ;
	assign \g216301/_0_  = _w15245_ ;
	assign \g216302/_0_  = _w15251_ ;
	assign \g216303/_0_  = _w15257_ ;
	assign \g216304/_0_  = _w15263_ ;
	assign \g216305/_0_  = _w15269_ ;
	assign \g216306/_0_  = _w15275_ ;
	assign \g216307/_0_  = _w15281_ ;
	assign \g216310/_3_  = _w15302_ ;
	assign \g216311/_3_  = _w15329_ ;
	assign \g216314/u3_syn_7  = _w13429_ ;
	assign \g216322/_3_  = _w15331_ ;
	assign \g216323/_3_  = _w15333_ ;
	assign \g216324/_3_  = _w15335_ ;
	assign \g216325/_3_  = _w15337_ ;
	assign \g216326/_3_  = _w15339_ ;
	assign \g216327/_3_  = _w15341_ ;
	assign \g216328/_3_  = _w15343_ ;
	assign \g216329/_3_  = _w15345_ ;
	assign \g216369/_0_  = _w15357_ ;
	assign \g216370/_0_  = _w15368_ ;
	assign \g216371/_0_  = _w15376_ ;
	assign \g216372/_0_  = _w15386_ ;
	assign \g216373/_0_  = _w15395_ ;
	assign \g216374/_0_  = _w15403_ ;
	assign \g216375/_0_  = _w15414_ ;
	assign \g216376/_0_  = _w15423_ ;
	assign \g216379/_0_  = _w15434_ ;
	assign \g216380/_0_  = _w15780_ ;
	assign \g216381/_0_  = _w15781_ ;
	assign \g216385/_0_  = _w16128_ ;
	assign \g216389/_0_  = _w16473_ ;
	assign \g216390/_0_  = _w16820_ ;
	assign \g216402/_0_  = _w16823_ ;
	assign \g216404/_0_  = _w16828_ ;
	assign \g216405/_0_  = _w16838_ ;
	assign \g216406/_0_  = _w16848_ ;
	assign \g216407/_0_  = _w16858_ ;
	assign \g216408/_0_  = _w16868_ ;
	assign \g216409/_0_  = _w16877_ ;
	assign \g216410/_0_  = _w16888_ ;
	assign \g216411/_0_  = _w16896_ ;
	assign \g216412/_0_  = _w16908_ ;
	assign \g216413/_0_  = _w16915_ ;
	assign \g216414/_0_  = _w16926_ ;
	assign \g216415/_0_  = _w16947_ ;
	assign \g216416/_0_  = _w16959_ ;
	assign \g216417/_0_  = _w16970_ ;
	assign \g216418/_0_  = _w16978_ ;
	assign \g216419/_0_  = _w16986_ ;
	assign \g216420/_0_  = _w16994_ ;
	assign \g216421/_0_  = _w17002_ ;
	assign \g216422/_0_  = _w17010_ ;
	assign \g216423/_0_  = _w17012_ ;
	assign \g216424/_0_  = _w17014_ ;
	assign \g216425/_0_  = _w17357_ ;
	assign \g216426/_0_  = _w17359_ ;
	assign \g216427/_0_  = _w17361_ ;
	assign \g216428/_0_  = _w17363_ ;
	assign \g216429/_0_  = _w17367_ ;
	assign \g216430/_0_  = _w17369_ ;
	assign \g216431/_0_  = _w17371_ ;
	assign \g216432/_0_  = _w17714_ ;
	assign \g216433/_0_  = _w17716_ ;
	assign \g216434/_0_  = _w18059_ ;
	assign \g216435/_0_  = _w18402_ ;
	assign \g216436/_0_  = _w18404_ ;
	assign \g216437/_0_  = _w18747_ ;
	assign \g216438/_0_  = _w18749_ ;
	assign \g216439/_3_  = _w18771_ ;
	assign \g216447/_3_  = _w18782_ ;
	assign \g216448/_3_  = _w19151_ ;
	assign \g216452/_0_  = _w19162_ ;
	assign \g216453/_0_  = _w19178_ ;
	assign \g216454/_0_  = _w19181_ ;
	assign \g216455/_0_  = _w19525_ ;
	assign \g216456/_0_  = _w19527_ ;
	assign \g216457/_0_  = _w19530_ ;
	assign \g216458/_3_  = _w19541_ ;
	assign \g216459/_3_  = _w19552_ ;
	assign \g216461/_3_  = _w19563_ ;
	assign \g216462/_3_  = _w19574_ ;
	assign \g216463/_3_  = _w19585_ ;
	assign \g216464/_3_  = _w19596_ ;
	assign \g216465/_3_  = _w19607_ ;
	assign \g216466/_0_  = _w19609_ ;
	assign \g216467/_3_  = _w19620_ ;
	assign \g216468/_3_  = _w19631_ ;
	assign \g216469/_3_  = _w20010_ ;
	assign \g216470/_3_  = _w20384_ ;
	assign \g216471/_3_  = _w20756_ ;
	assign \g216473/_3_  = _w21119_ ;
	assign \g216474/_3_  = _w21482_ ;
	assign \g216475/_3_  = _w21843_ ;
	assign \g216476/_3_  = _w21854_ ;
	assign \g216477/_3_  = _w22215_ ;
	assign \g216478/_0_  = _w22220_ ;
	assign \g216479/_3_  = _w22596_ ;
	assign \g216480/_3_  = _w22632_ ;
	assign \g216481/_3_  = _w22672_ ;
	assign \g216492/_0_  = _w22675_ ;
	assign \g216494/_0_  = _w22691_ ;
	assign \g216495/_3_  = _w22707_ ;
	assign \g216496/_3_  = _w23077_ ;
	assign \g216498/_3_  = _w23090_ ;
	assign \g216499/_3_  = _w23103_ ;
	assign \g216500/_3_  = _w23116_ ;
	assign \g216513/_3_  = _w23122_ ;
	assign \g216514/_3_  = _w23126_ ;
	assign \g216515/_3_  = _w23128_ ;
	assign \g216516/_3_  = _w23132_ ;
	assign \g216517/_3_  = _w23137_ ;
	assign \g216518/_3_  = _w23141_ ;
	assign \g216519/_3_  = _w23147_ ;
	assign \g216520/_3_  = _w23153_ ;
	assign \g216521/_3_  = _w23157_ ;
	assign \g216522/_3_  = _w23161_ ;
	assign \g216523/_3_  = _w23163_ ;
	assign \g216524/_3_  = _w23166_ ;
	assign \g216525/_3_  = _w23172_ ;
	assign \g216526/_3_  = _w23179_ ;
	assign \g216527/_3_  = _w23183_ ;
	assign \g216528/_3_  = _w23188_ ;
	assign \g216529/_3_  = _w23192_ ;
	assign \g216530/_3_  = _w23198_ ;
	assign \g216531/_3_  = _w23200_ ;
	assign \g216532/_3_  = _w23207_ ;
	assign \g216533/_3_  = _w23211_ ;
	assign \g216534/_3_  = _w23216_ ;
	assign \g216535/_3_  = _w23218_ ;
	assign \g216536/_3_  = _w23220_ ;
	assign \g216537/_3_  = _w23225_ ;
	assign \g216538/_3_  = _w23230_ ;
	assign \g216555/_3_  = _w23591_ ;
	assign \g216556/_3_  = _w23952_ ;
	assign \g216557/_3_  = _w23972_ ;
	assign \g216560/_3_  = _w23976_ ;
	assign \g216561/_3_  = _w23980_ ;
	assign \g216562/_3_  = _w23982_ ;
	assign \g216563/_3_  = _w23985_ ;
	assign \g216564/_3_  = _w23987_ ;
	assign \g216565/_3_  = _w23991_ ;
	assign \g216566/_3_  = _w23995_ ;
	assign \g216567/_3_  = _w23997_ ;
	assign \g216568/_3_  = _w23999_ ;
	assign \g216569/_3_  = _w24002_ ;
	assign \g216570/_3_  = _w24006_ ;
	assign \g216571/_3_  = _w24008_ ;
	assign \g216575/_3_  = _w24014_ ;
	assign \g216576/_3_  = _w24016_ ;
	assign \g216577/_3_  = _w24018_ ;
	assign \g216578/_3_  = _w24021_ ;
	assign \g216579/_3_  = _w24025_ ;
	assign \g216580/_3_  = _w24027_ ;
	assign \g216581/_3_  = _w24029_ ;
	assign \g216582/_3_  = _w24032_ ;
	assign \g216583/_3_  = _w24036_ ;
	assign \g216586/_3_  = _w24383_ ;
	assign \g216587/_3_  = _w24385_ ;
	assign \g216588/_3_  = _w24387_ ;
	assign \g216589/_3_  = _w24390_ ;
	assign \g216590/_3_  = _w24395_ ;
	assign \g216591/_3_  = _w24399_ ;
	assign \g216592/_3_  = _w24401_ ;
	assign \g216593/_3_  = _w24403_ ;
	assign \g216594/_3_  = _w24406_ ;
	assign \g216595/_3_  = _w24410_ ;
	assign \g216600/_3_  = _w24422_ ;
	assign \g216683/_0_  = _w24431_ ;
	assign \g216689/_0_  = _w24432_ ;
	assign \g216693/_0_  = _w24439_ ;
	assign \g216694/_0_  = _w24443_ ;
	assign \g216727/_0_  = _w24448_ ;
	assign \g216728/_0_  = _w24449_ ;
	assign \g216729/_0_  = _w24452_ ;
	assign \g216732/_0_  = _w24453_ ;
	assign \g216733/_0_  = _w24457_ ;
	assign \g216734/_0_  = _w24460_ ;
	assign \g216735/_0_  = _w24465_ ;
	assign \g216736/_0_  = _w24467_ ;
	assign \g216737/_0_  = _w24468_ ;
	assign \g216738/_0_  = _w24473_ ;
	assign \g216739/_0_  = _w24475_ ;
	assign \g216740/_0_  = _w24479_ ;
	assign \g216741/_0_  = _w24480_ ;
	assign \g216742/_0_  = _w24483_ ;
	assign \g216743/_0_  = _w24487_ ;
	assign \g216744/_0_  = _w24492_ ;
	assign \g216745/_0_  = _w24495_ ;
	assign \g216746/_0_  = _w24500_ ;
	assign \g216748/_0_  = _w24517_ ;
	assign \g216751/_0_  = _w24522_ ;
	assign \g216754/_0_  = _w24528_ ;
	assign \g216762/_0_  = _w24529_ ;
	assign \g216934/_2_  = _w24531_ ;
	assign \g216952/_0_  = _w24543_ ;
	assign \g216955/_0_  = _w24544_ ;
	assign \g216969/_0_  = _w24550_ ;
	assign \g216979/_0_  = _w24552_ ;
	assign \g216984/_0_  = _w24554_ ;
	assign \g216996/_0_  = _w24557_ ;
	assign \g217002/_0_  = _w24560_ ;
	assign \g217014/_0_  = _w24579_ ;
	assign \g217015/_0_  = _w24591_ ;
	assign \g217016/_0_  = _w24603_ ;
	assign \g217017/_0_  = _w24615_ ;
	assign \g217018/_0_  = _w24627_ ;
	assign \g217019/_0_  = _w24636_ ;
	assign \g217023/_0_  = _w24639_ ;
	assign \g217116/_0_  = _w24749_ ;
	assign \g217146/_3_  = _w24770_ ;
	assign \g217149/_0_  = _w24772_ ;
	assign \g217151/_0_  = _w24776_ ;
	assign \g217160/_0_  = _w24780_ ;
	assign \g217167/_0_  = _w24783_ ;
	assign \g217168/_0_  = _w24787_ ;
	assign \g217169/_0_  = _w24791_ ;
	assign \g217170/_0_  = _w24794_ ;
	assign \g217171/_0_  = _w24797_ ;
	assign \g217172/_0_  = _w24800_ ;
	assign \g217173/_0_  = _w24803_ ;
	assign \g217174/_0_  = _w24806_ ;
	assign \g217175/_0_  = _w24809_ ;
	assign \g217176/_0_  = _w24811_ ;
	assign \g217177/_0_  = _w24813_ ;
	assign \g217178/_0_  = _w24815_ ;
	assign \g217179/_0_  = _w24817_ ;
	assign \g217180/_0_  = _w24819_ ;
	assign \g217181/_0_  = _w24821_ ;
	assign \g217182/_0_  = _w24823_ ;
	assign \g217183/_0_  = _w24825_ ;
	assign \g217187/_0_  = _w24829_ ;
	assign \g217188/_0_  = _w24832_ ;
	assign \g217189/_0_  = _w24836_ ;
	assign \g217193/_0_  = _w24839_ ;
	assign \g217194/_0_  = _w24841_ ;
	assign \g217195/_0_  = _w24850_ ;
	assign \g217196/_0_  = _w24858_ ;
	assign \g217202/_0_  = _w24860_ ;
	assign \g217205/_0_  = _w24865_ ;
	assign \g217206/_0_  = _w24870_ ;
	assign \g217207/_0_  = _w24875_ ;
	assign \g217208/_0_  = _w24880_ ;
	assign \g217209/_0_  = _w24885_ ;
	assign \g217210/_0_  = _w24890_ ;
	assign \g217211/_0_  = _w24895_ ;
	assign \g217212/_0_  = _w24900_ ;
	assign \g217213/_0_  = _w24905_ ;
	assign \g217214/_0_  = _w24910_ ;
	assign \g217215/_0_  = _w24915_ ;
	assign \g217216/_0_  = _w24920_ ;
	assign \g217217/_0_  = _w24925_ ;
	assign \g217218/_0_  = _w24930_ ;
	assign \g217219/_0_  = _w24935_ ;
	assign \g217220/_0_  = _w24940_ ;
	assign \g217223/_0_  = _w24942_ ;
	assign \g217231/_0_  = _w24945_ ;
	assign \g217237/_0_  = _w24954_ ;
	assign \g217238/_0_  = _w24963_ ;
	assign \g217242/_0_  = _w24964_ ;
	assign \g217243/_0_  = _w24969_ ;
	assign \g217250/_3_  = _w24998_ ;
	assign \g217251/_3_  = _w25011_ ;
	assign \g217252/_3_  = _w25023_ ;
	assign \g217253/_3_  = _w25036_ ;
	assign \g217254/_3_  = _w25048_ ;
	assign \g217255/_3_  = _w25061_ ;
	assign \g217256/_3_  = _w25073_ ;
	assign \g217257/_3_  = _w25086_ ;
	assign \g217258/_3_  = _w25098_ ;
	assign \g217259/_3_  = _w25110_ ;
	assign \g217260/_3_  = _w25122_ ;
	assign \g217261/_3_  = _w25135_ ;
	assign \g217262/_3_  = _w25148_ ;
	assign \g217263/_3_  = _w25160_ ;
	assign \g217264/_3_  = _w25172_ ;
	assign \g217265/_3_  = _w25184_ ;
	assign \g217266/_3_  = _w25196_ ;
	assign \g217267/_3_  = _w25208_ ;
	assign \g217268/_3_  = _w25220_ ;
	assign \g217269/_3_  = _w25233_ ;
	assign \g217270/_3_  = _w25246_ ;
	assign \g217271/_3_  = _w25259_ ;
	assign \g217272/_3_  = _w25271_ ;
	assign \g217273/_3_  = _w25283_ ;
	assign \g217274/_3_  = _w25296_ ;
	assign \g217275/_3_  = _w25308_ ;
	assign \g217276/_3_  = _w25321_ ;
	assign \g217277/_3_  = _w25334_ ;
	assign \g217278/_3_  = _w25346_ ;
	assign \g217279/_3_  = _w25359_ ;
	assign \g217280/_3_  = _w25371_ ;
	assign \g217281/_3_  = _w25384_ ;
	assign \g217282/_3_  = _w25414_ ;
	assign \g217283/_3_  = _w25426_ ;
	assign \g217284/_3_  = _w25438_ ;
	assign \g217285/_3_  = _w25450_ ;
	assign \g217286/_3_  = _w25462_ ;
	assign \g217287/_3_  = _w25474_ ;
	assign \g217288/_3_  = _w25486_ ;
	assign \g217289/_3_  = _w25498_ ;
	assign \g217290/_3_  = _w25510_ ;
	assign \g217291/_3_  = _w25522_ ;
	assign \g217292/_3_  = _w25534_ ;
	assign \g217293/_3_  = _w25546_ ;
	assign \g217294/_3_  = _w25558_ ;
	assign \g217295/_3_  = _w25570_ ;
	assign \g217296/_3_  = _w25582_ ;
	assign \g217297/_3_  = _w25594_ ;
	assign \g217298/_3_  = _w25606_ ;
	assign \g217299/_3_  = _w25618_ ;
	assign \g217300/_3_  = _w25630_ ;
	assign \g217301/_3_  = _w25642_ ;
	assign \g217302/_3_  = _w25654_ ;
	assign \g217303/_3_  = _w25666_ ;
	assign \g217304/_3_  = _w25678_ ;
	assign \g217305/_3_  = _w25690_ ;
	assign \g217306/_3_  = _w25702_ ;
	assign \g217307/_3_  = _w25714_ ;
	assign \g217308/_3_  = _w25726_ ;
	assign \g217309/_3_  = _w25738_ ;
	assign \g217310/_3_  = _w25750_ ;
	assign \g217311/_3_  = _w25762_ ;
	assign \g217312/_3_  = _w25774_ ;
	assign \g217313/_3_  = _w25786_ ;
	assign \g217318/_0_  = _w25791_ ;
	assign \g217662/_0_  = _w25804_ ;
	assign \g217663/_0_  = _w25806_ ;
	assign \g217682/_0_  = _w25814_ ;
	assign \g217697/_0_  = _w25826_ ;
	assign \g217698/_0_  = _w25841_ ;
	assign \g217699/_0_  = _w25844_ ;
	assign \g217700/_0_  = _w25845_ ;
	assign \g217701/_0_  = _w25847_ ;
	assign \g217705/_0_  = _w25852_ ;
	assign \g217711/_0_  = _w25855_ ;
	assign \g217747/_0_  = _w25858_ ;
	assign \g217753/_00_  = _w25863_ ;
	assign \g217775/_0_  = _w25873_ ;
	assign \g217781/_0_  = _w25885_ ;
	assign \g217784/_0_  = _w25887_ ;
	assign \g217785/_0_  = _w25891_ ;
	assign \g217786/_0_  = _w25895_ ;
	assign \g217787/_0_  = _w25898_ ;
	assign \g217788/_0_  = _w25901_ ;
	assign \g217790/_0_  = _w25904_ ;
	assign \g217815/_0_  = _w25909_ ;
	assign \g217817/_0_  = _w25912_ ;
	assign \g218145/_0_  = _w25914_ ;
	assign \g218148/_0_  = _w25919_ ;
	assign \g218150/_0_  = _w25936_ ;
	assign \g218167/_0_  = _w25944_ ;
	assign \g218168/_0_  = _w25948_ ;
	assign \g218234/_0_  = _w25949_ ;
	assign \g218235/_0_  = _w25950_ ;
	assign \g218236/_0_  = _w25953_ ;
	assign \g218238/_0_  = _w25957_ ;
	assign \g218242/_0_  = _w25958_ ;
	assign \g218332/_0_  = _w25963_ ;
	assign \g218335/_0_  = _w25968_ ;
	assign \g218336/_0_  = _w25973_ ;
	assign \g218337/_0_  = _w25980_ ;
	assign \g218338/_0_  = _w25984_ ;
	assign \g218339/_0_  = _w25988_ ;
	assign \g218340/_0_  = _w25992_ ;
	assign \g218341/_0_  = _w25996_ ;
	assign \g218342/_0_  = _w26000_ ;
	assign \g218343/_0_  = _w26006_ ;
	assign \g218344/_0_  = _w26010_ ;
	assign \g218345/_0_  = _w26013_ ;
	assign \g218346/_0_  = _w26016_ ;
	assign \g218347/_0_  = _w26019_ ;
	assign \g218348/_0_  = _w26022_ ;
	assign \g218349/_0_  = _w26025_ ;
	assign \g218350/_0_  = _w26028_ ;
	assign \g218351/_0_  = _w26033_ ;
	assign \g218352/_0_  = _w26036_ ;
	assign \g218353/_0_  = _w26039_ ;
	assign \g218354/_0_  = _w26042_ ;
	assign \g218355/_0_  = _w26045_ ;
	assign \g218356/_0_  = _w26048_ ;
	assign \g218357/_0_  = _w26051_ ;
	assign \g218358/_0_  = _w26054_ ;
	assign \g218359/_0_  = _w26057_ ;
	assign \g218360/_0_  = _w26060_ ;
	assign \g218398/_3_  = _w26062_ ;
	assign \g218430/_0_  = _w26067_ ;
	assign \g218440/_0_  = _w26072_ ;
	assign \g218452/u3_syn_4  = _w26077_ ;
	assign \g218495/u3_syn_4  = _w26080_ ;
	assign \g218517/u3_syn_4  = _w26082_ ;
	assign \g218554/u3_syn_4  = _w26087_ ;
	assign \g218575/u3_syn_4  = _w26089_ ;
	assign \g218600/u3_syn_4  = _w26091_ ;
	assign \g218621/u3_syn_4  = _w26092_ ;
	assign \g218638/u3_syn_4  = _w26093_ ;
	assign \g218659/u3_syn_4  = _w26097_ ;
	assign \g218673/u3_syn_4  = _w26100_ ;
	assign \g218707/u3_syn_4  = _w26103_ ;
	assign \g218735/_3_  = _w26104_ ;
	assign \g219186/_0_  = _w26107_ ;
	assign \g219187/_0_  = _w26113_ ;
	assign \g219188/_0_  = _w26117_ ;
	assign \g219189/_0_  = _w26120_ ;
	assign \g219190/_0_  = _w26129_ ;
	assign \g219196/_0_  = _w26132_ ;
	assign \g219198/_0_  = _w26134_ ;
	assign \g219199/_0_  = _w26140_ ;
	assign \g219200/_0_  = _w26144_ ;
	assign \g219308/_0_  = _w26146_ ;
	assign \g219314/_0_  = _w26147_ ;
	assign \g219326/_0_  = _w26150_ ;
	assign \g219328/_0_  = _w26153_ ;
	assign \g219348/_0_  = _w26161_ ;
	assign \g219351/_0_  = _w26163_ ;
	assign \g219363/_0_  = _w26166_ ;
	assign \g219364/_0_  = _w26170_ ;
	assign \g219365/_0_  = _w26172_ ;
	assign \g219366/_0_  = _w26174_ ;
	assign \g219367/_0_  = _w26176_ ;
	assign \g219368/_0_  = _w26178_ ;
	assign \g219369/_0_  = _w26180_ ;
	assign \g219376/_0_  = _w26182_ ;
	assign \g219381/_0_  = _w26185_ ;
	assign \g219382/_0_  = _w26190_ ;
	assign \g219384/_0_  = _w26191_ ;
	assign \g219385/_0_  = _w26197_ ;
	assign \g219391/_0_  = _w26200_ ;
	assign \g219394/_0_  = _w26205_ ;
	assign \g219395/_0_  = _w26206_ ;
	assign \g219396/_0_  = _w26207_ ;
	assign \g219397/_0_  = _w26208_ ;
	assign \g219398/_0_  = _w26209_ ;
	assign \g219399/_0_  = _w26212_ ;
	assign \g219400/_0_  = _w26213_ ;
	assign \g219401/_0_  = _w26214_ ;
	assign \g219402/_0_  = _w26215_ ;
	assign \g219403/_0_  = _w26216_ ;
	assign \g219404/_0_  = _w26217_ ;
	assign \g219405/_0_  = _w26218_ ;
	assign \g219406/_0_  = _w26219_ ;
	assign \g219407/_0_  = _w26220_ ;
	assign \g219408/_0_  = _w26221_ ;
	assign \g219409/_0_  = _w26223_ ;
	assign \g219410/_0_  = _w26224_ ;
	assign \g219411/_0_  = _w26225_ ;
	assign \g219412/_0_  = _w26226_ ;
	assign \g219413/_0_  = _w26227_ ;
	assign \g219414/_0_  = _w26228_ ;
	assign \g219415/_0_  = _w26229_ ;
	assign \g219416/_0_  = _w26230_ ;
	assign \g219417/_0_  = _w26231_ ;
	assign \g219418/_0_  = _w26232_ ;
	assign \g219419/_0_  = _w26233_ ;
	assign \g219420/_0_  = _w26234_ ;
	assign \g219421/_0_  = _w26235_ ;
	assign \g219422/_0_  = _w26236_ ;
	assign \g219423/_0_  = _w26237_ ;
	assign \g219424/_0_  = _w26238_ ;
	assign \g219425/_0_  = _w26239_ ;
	assign \g219426/_0_  = _w26240_ ;
	assign \g219427/_0_  = _w26241_ ;
	assign \g219428/_0_  = _w26242_ ;
	assign \g219429/_0_  = _w26243_ ;
	assign \g219430/_0_  = _w26244_ ;
	assign \g219431/_0_  = _w26247_ ;
	assign \g219432/_0_  = _w26248_ ;
	assign \g219433/_0_  = _w26249_ ;
	assign \g219434/_0_  = _w26250_ ;
	assign \g219435/_0_  = _w26251_ ;
	assign \g219436/_0_  = _w26252_ ;
	assign \g219437/_0_  = _w26253_ ;
	assign \g219438/_0_  = _w26254_ ;
	assign \g219439/_0_  = _w26255_ ;
	assign \g219440/_0_  = _w26256_ ;
	assign \g219441/_0_  = _w26257_ ;
	assign \g219442/_0_  = _w26258_ ;
	assign \g219443/_0_  = _w26259_ ;
	assign \g219444/_0_  = _w26260_ ;
	assign \g219445/_0_  = _w26261_ ;
	assign \g219446/_0_  = _w26262_ ;
	assign \g219447/_0_  = _w26263_ ;
	assign \g219449/_0_  = _w26265_ ;
	assign \g219450/_0_  = _w26266_ ;
	assign \g219451/_0_  = _w26267_ ;
	assign \g219452/_0_  = _w26268_ ;
	assign \g219453/_0_  = _w26269_ ;
	assign \g219454/_0_  = _w26270_ ;
	assign \g219455/_0_  = _w26271_ ;
	assign \g219456/_0_  = _w26272_ ;
	assign \g219457/_0_  = _w26273_ ;
	assign \g219458/_0_  = _w26274_ ;
	assign \g219464/u3_syn_7  = _w26277_ ;
	assign \g219496/u3_syn_4  = _w26278_ ;
	assign \g219512/u3_syn_4  = _w26082_ ;
	assign \g219526/u3_syn_4  = _w26280_ ;
	assign \g219549/u3_syn_4  = _w26281_ ;
	assign \g219571/u3_syn_4  = _w26087_ ;
	assign \g219588/u3_syn_4  = _w26092_ ;
	assign \g219603/u3_syn_4  = _w26100_ ;
	assign \g219621/u3_syn_4  = _w26282_ ;
	assign \g219636/_3_  = _w26285_ ;
	assign \g219652/u3_syn_4  = _w26288_ ;
	assign \g219676/_3_  = _w26290_ ;
	assign \g219686/_0_  = _w26291_ ;
	assign \g219689/_0_  = _w26292_ ;
	assign \g219694/_3_  = _w26293_ ;
	assign \g220062/_0_  = _w26294_ ;
	assign \g220068/_0_  = _w26295_ ;
	assign \g220069/_0_  = _w26297_ ;
	assign \g220072/_0_  = _w26300_ ;
	assign \g220084/_0_  = _w26301_ ;
	assign \g220149/_0_  = _w26305_ ;
	assign \g220162/_0_  = _w26310_ ;
	assign \g220317/_0_  = _w26314_ ;
	assign \g220360/_2_  = _w11392_ ;
	assign \g220368/_2_  = _w26316_ ;
	assign \g220369/_0_  = _w26328_ ;
	assign \g220370/_0_  = _w26334_ ;
	assign \g220371/_0_  = _w26339_ ;
	assign \g220372/_0_  = _w26346_ ;
	assign \g220376/_0_  = _w26354_ ;
	assign \g220390/_0_  = _w26375_ ;
	assign \g220395/_0_  = _w26380_ ;
	assign \g220499/_0_  = _w26395_ ;
	assign \g220500/_0_  = _w26401_ ;
	assign \g220501/_0_  = _w26407_ ;
	assign \g220502/_0_  = _w26413_ ;
	assign \g220503/_0_  = _w26419_ ;
	assign \g220504/_0_  = _w26425_ ;
	assign \g220505/_0_  = _w26431_ ;
	assign \g220506/_0_  = _w26437_ ;
	assign \g220507/_0_  = _w26443_ ;
	assign \g220508/_0_  = _w26449_ ;
	assign \g220509/_0_  = _w26455_ ;
	assign \g220510/_0_  = _w26461_ ;
	assign \g220511/_0_  = _w26467_ ;
	assign \g220512/_0_  = _w26473_ ;
	assign \g220513/_0_  = _w26479_ ;
	assign \g220514/_0_  = _w26485_ ;
	assign \g220515/_0_  = _w26491_ ;
	assign \g220516/_0_  = _w26497_ ;
	assign \g220517/_0_  = _w26503_ ;
	assign \g220518/_0_  = _w26509_ ;
	assign \g220519/_0_  = _w26515_ ;
	assign \g220520/_0_  = _w26521_ ;
	assign \g220521/_0_  = _w26527_ ;
	assign \g220522/_0_  = _w26533_ ;
	assign \g220523/_0_  = _w26539_ ;
	assign \g220524/_0_  = _w26545_ ;
	assign \g220525/_0_  = _w26551_ ;
	assign \g220526/_0_  = _w26557_ ;
	assign \g220527/_0_  = _w26563_ ;
	assign \g220528/_0_  = _w26569_ ;
	assign \g220529/_0_  = _w26575_ ;
	assign \g220530/_0_  = _w26581_ ;
	assign \g220531/_0_  = _w26587_ ;
	assign \g220532/_0_  = _w26593_ ;
	assign \g220533/_0_  = _w26599_ ;
	assign \g220534/_0_  = _w26602_ ;
	assign \g220535/_0_  = _w26607_ ;
	assign \g220557/_0_  = _w26613_ ;
	assign \g220558/_0_  = _w26614_ ;
	assign \g220559/_0_  = _w26615_ ;
	assign \g220560/_0_  = _w26616_ ;
	assign \g220561/_0_  = _w26617_ ;
	assign \g220562/_0_  = _w26618_ ;
	assign \g220563/_0_  = _w26619_ ;
	assign \g220564/_0_  = _w26620_ ;
	assign \g220565/_0_  = _w26621_ ;
	assign \g220566/_0_  = _w26622_ ;
	assign \g220567/_0_  = _w26623_ ;
	assign \g220568/_0_  = _w26624_ ;
	assign \g220569/_0_  = _w26625_ ;
	assign \g220570/_0_  = _w26626_ ;
	assign \g220571/_0_  = _w26632_ ;
	assign \g220572/_0_  = _w26634_ ;
	assign \g220573/_0_  = _w26636_ ;
	assign \g220574/_0_  = _w26638_ ;
	assign \g220575/_0_  = _w26640_ ;
	assign \g220576/_0_  = _w26642_ ;
	assign \g220577/_0_  = _w26644_ ;
	assign \g220578/_0_  = _w26646_ ;
	assign \g220579/_0_  = _w26648_ ;
	assign \g220580/_0_  = _w26650_ ;
	assign \g220581/_0_  = _w26652_ ;
	assign \g220582/_0_  = _w26654_ ;
	assign \g220583/_0_  = _w26656_ ;
	assign \g220584/_0_  = _w26658_ ;
	assign \g220585/_0_  = _w26660_ ;
	assign \g220586/_0_  = _w26662_ ;
	assign \g220587/_0_  = _w26665_ ;
	assign \g220588/_0_  = _w26666_ ;
	assign \g220589/_0_  = _w26667_ ;
	assign \g220590/_0_  = _w26668_ ;
	assign \g220591/_0_  = _w26669_ ;
	assign \g220592/_0_  = _w26670_ ;
	assign \g220593/_0_  = _w26671_ ;
	assign \g220594/_0_  = _w26672_ ;
	assign \g220595/_0_  = _w26673_ ;
	assign \g220596/_0_  = _w26674_ ;
	assign \g220597/_0_  = _w26675_ ;
	assign \g220598/_0_  = _w26676_ ;
	assign \g220599/_0_  = _w26677_ ;
	assign \g220600/_0_  = _w26678_ ;
	assign \g220601/_0_  = _w26679_ ;
	assign \g220602/_0_  = _w26680_ ;
	assign \g220603/_0_  = _w26681_ ;
	assign \g220604/_0_  = _w26685_ ;
	assign \g220605/_0_  = _w26687_ ;
	assign \g220606/_0_  = _w26689_ ;
	assign \g220607/_0_  = _w26691_ ;
	assign \g220608/_0_  = _w26693_ ;
	assign \g220609/_0_  = _w26695_ ;
	assign \g220610/_0_  = _w26697_ ;
	assign \g220611/_0_  = _w26699_ ;
	assign \g220612/_0_  = _w26701_ ;
	assign \g220613/_0_  = _w26703_ ;
	assign \g220614/_0_  = _w26705_ ;
	assign \g220615/_0_  = _w26707_ ;
	assign \g220616/_0_  = _w26709_ ;
	assign \g220617/_0_  = _w26711_ ;
	assign \g220618/_0_  = _w26713_ ;
	assign \g220619/_0_  = _w26715_ ;
	assign \g220620/_0_  = _w26720_ ;
	assign \g220621/_0_  = _w26722_ ;
	assign \g220622/_0_  = _w26724_ ;
	assign \g220623/_0_  = _w26726_ ;
	assign \g220624/_0_  = _w26728_ ;
	assign \g220625/_0_  = _w26730_ ;
	assign \g220626/_0_  = _w26732_ ;
	assign \g220627/_0_  = _w26734_ ;
	assign \g220628/_0_  = _w26736_ ;
	assign \g220629/_0_  = _w26738_ ;
	assign \g220630/_0_  = _w26740_ ;
	assign \g220631/_0_  = _w26742_ ;
	assign \g220632/_0_  = _w26744_ ;
	assign \g220633/_0_  = _w26746_ ;
	assign \g220634/_0_  = _w26748_ ;
	assign \g220635/_0_  = _w26750_ ;
	assign \g220636/_0_  = _w26752_ ;
	assign \g220637/_0_  = _w26754_ ;
	assign \g220638/_0_  = _w26756_ ;
	assign \g220639/_0_  = _w26758_ ;
	assign \g220640/_0_  = _w26760_ ;
	assign \g220641/_0_  = _w26762_ ;
	assign \g220642/_0_  = _w26764_ ;
	assign \g220643/_0_  = _w26769_ ;
	assign \g220644/_0_  = _w26770_ ;
	assign \g220645/_0_  = _w26771_ ;
	assign \g220646/_0_  = _w26772_ ;
	assign \g220647/_0_  = _w26773_ ;
	assign \g220648/_0_  = _w26774_ ;
	assign \g220649/_0_  = _w26775_ ;
	assign \g220650/_0_  = _w26776_ ;
	assign \g220651/_0_  = _w26777_ ;
	assign \g220652/_0_  = _w26778_ ;
	assign \g220653/_0_  = _w26779_ ;
	assign \g220654/_0_  = _w26780_ ;
	assign \g220655/_0_  = _w26781_ ;
	assign \g220656/_0_  = _w26782_ ;
	assign \g220657/_0_  = _w26783_ ;
	assign \g220658/_0_  = _w26784_ ;
	assign \g220659/_0_  = _w26785_ ;
	assign \g220660/_0_  = _w26786_ ;
	assign \g220661/_0_  = _w26787_ ;
	assign \g220662/_0_  = _w26788_ ;
	assign \g220663/_0_  = _w26789_ ;
	assign \g220664/_0_  = _w26790_ ;
	assign \g220665/_0_  = _w26791_ ;
	assign \g220666/_0_  = _w26792_ ;
	assign \g220674/_0_  = _w26794_ ;
	assign \g220679/u3_syn_7  = _w26797_ ;
	assign \g220711/u3_syn_4  = _w26798_ ;
	assign \g220726/u3_syn_4  = _w26800_ ;
	assign \g220739/u3_syn_4  = _w26802_ ;
	assign \g220751/u3_syn_4  = _w26804_ ;
	assign \g220759/u3_syn_4  = _w26806_ ;
	assign \g220773/u3_syn_4  = _w26807_ ;
	assign \g220782/u3_syn_4  = _w26809_ ;
	assign \g220805/u3_syn_4  = _w26811_ ;
	assign \g220828/u3_syn_4  = _w26813_ ;
	assign \g220921/_0_  = _w25955_ ;
	assign \g220930/u3_syn_4  = _w26815_ ;
	assign \g220949/_3_  = _w26817_ ;
	assign \g220994/_3_  = _w26818_ ;
	assign \g221207/_0_  = _w26834_ ;
	assign \g221213/_0_  = _w11063_ ;
	assign \g221223/_0_  = _w26837_ ;
	assign \g221224/_0_  = _w26840_ ;
	assign \g221225/_0_  = _w26846_ ;
	assign \g221226/_0_  = _w26850_ ;
	assign \g221231/_0_  = _w26856_ ;
	assign \g221232/_0_  = _w26861_ ;
	assign \g221234/_0_  = _w26866_ ;
	assign \g221235/_0_  = _w26868_ ;
	assign \g221246/_2_  = _w11065_ ;
	assign \g221249/_2_  = _w11067_ ;
	assign \g221265/_0_  = _w26870_ ;
	assign \g221287/_0_  = _w26873_ ;
	assign \g221325/_0_  = _w26877_ ;
	assign \g221326/_0_  = _w26882_ ;
	assign \g221447/_0_  = _w26885_ ;
	assign \g221449/_0_  = _w26888_ ;
	assign \g221452/_0_  = _w26889_ ;
	assign \g221469/_0_  = _w26890_ ;
	assign \g221473/_0_  = _w26899_ ;
	assign \g221503/_0_  = _w26900_ ;
	assign \g221510/_0_  = _w26906_ ;
	assign \g221512/_0_  = _w26910_ ;
	assign \g221516/_0_  = _w26915_ ;
	assign \g221517/_0_  = _w26920_ ;
	assign \g221524/_0_  = _w26924_ ;
	assign \g221530/_0_  = _w26931_ ;
	assign \g221592/_0_  = _w26932_ ;
	assign \g221593/_0_  = _w26933_ ;
	assign \g221634/u3_syn_4  = _w26612_ ;
	assign \g221669/u3_syn_4  = _w26630_ ;
	assign \g221789/u3_syn_4  = _w26664_ ;
	assign \g221813/u3_syn_4  = _w26683_ ;
	assign \g221829/u3_syn_4  = _w26718_ ;
	assign \g221861/u3_syn_4  = _w26768_ ;
	assign \g221876/_0_  = _w26934_ ;
	assign \g221935/_0_  = _w26940_ ;
	assign \g221944/_3_  = _w11046_ ;
	assign \g230200/_0_  = _w26942_ ;
	assign \g230201/_0_  = _w26943_ ;
	assign \g230205/_0_  = _w26944_ ;
	assign \g230295/_0_  = _w26948_ ;
	assign \g230297/_0_  = _w26952_ ;
	assign \g230298/_0_  = _w26956_ ;
	assign \g230300/_0_  = _w26959_ ;
	assign \g230302/_0_  = _w26967_ ;
	assign \g230303/_0_  = _w26973_ ;
	assign \g230343/_0_  = _w26975_ ;
	assign \g230368/_0_  = _w26977_ ;
	assign \g230511/_0_  = _w26980_ ;
	assign \g230531/_0_  = _w26981_ ;
	assign \g230635/_2_  = _w26982_ ;
	assign \g230661/_0_  = _w26983_ ;
	assign \g230715/_1__syn_2  = _w26984_ ;
	assign \g230731/_0_  = _w27002_ ;
	assign \g230766/_0_  = _w27003_ ;
	assign \g230784/_0_  = _w27006_ ;
	assign \g230785/_0_  = _w27009_ ;
	assign \g230786/_0_  = _w27012_ ;
	assign \g230787/_0_  = _w27015_ ;
	assign \g230797/_0_  = _w27018_ ;
	assign \g230798/_0_  = _w27019_ ;
	assign \g230803/_0_  = _w27020_ ;
	assign \g230804/_00_  = _w27025_ ;
	assign \g230805/_00_  = _w27030_ ;
	assign \g230806/_00_  = _w27035_ ;
	assign \g230807/_00_  = _w27040_ ;
	assign \g230808/_00_  = _w27045_ ;
	assign \g230809/_00_  = _w27050_ ;
	assign \g230815/_0_  = _w27053_ ;
	assign \g230816/_2_  = _w27055_ ;
	assign \g230817/_2_  = _w27060_ ;
	assign \g230829/_0_  = _w27069_ ;
	assign \g230834/_0_  = _w27075_ ;
	assign \g230835/_0_  = _w27081_ ;
	assign \g230836/_0_  = _w27085_ ;
	assign \g230837/_0_  = _w27091_ ;
	assign \g230844/_0_  = _w27093_ ;
	assign \g230863/_3_  = _w27099_ ;
	assign \g230864/_3_  = _w27103_ ;
	assign \g230870/_0_  = _w27110_ ;
	assign \g230988/_3_  = _w27113_ ;
	assign \g231010/_3_  = _w27117_ ;
	assign \g231016/_3_  = _w27121_ ;
	assign \g231042/_3_  = _w27125_ ;
	assign \g231471/_0_  = _w27128_ ;
	assign \g231472/_0_  = _w27131_ ;
	assign \g231476/_3_  = _w27132_ ;
	assign \g231480/_3_  = _w27133_ ;
	assign \g231484/_3_  = _w27134_ ;
	assign \g231504/_0_  = _w27136_ ;
	assign \g231532/_0_  = _w24561_ ;
	assign \g231542/_0_  = _w27139_ ;
	assign \g231560/_1_  = _w27142_ ;
	assign \g231578/_1_  = _w27144_ ;
	assign \g231580/_0_  = _w27146_ ;
	assign \g231590/_1__syn_2  = _w25812_ ;
	assign \g231615/_0_  = _w27148_ ;
	assign \g231623/_1_  = _w27149_ ;
	assign \g231634/_2_  = _w27150_ ;
	assign \g231635/_0_  = _w27152_ ;
	assign \g231638/_2_  = _w27154_ ;
	assign \g231640/_0_  = _w27156_ ;
	assign \g231653/_2_  = _w27158_ ;
	assign \g231787/_0_  = _w27160_ ;
	assign \g231931/_0_  = _w27165_ ;
	assign \g231939/_3_  = _w27167_ ;
	assign \g231940/_0_  = _w27170_ ;
	assign \g231951/_0_  = _w27173_ ;
	assign \g231955/_0_  = _w27174_ ;
	assign \g231956/_0_  = _w27178_ ;
	assign \g231959/_2_  = _w27181_ ;
	assign \g231960/_0_  = _w27182_ ;
	assign \g231964/_0_  = _w27188_ ;
	assign \g231965/_0_  = _w27191_ ;
	assign \g231975/_0_  = _w27195_ ;
	assign \g231986/_1_  = _w27197_ ;
	assign \g231987/_1_  = _w27198_ ;
	assign \g231989/_1_  = _w27200_ ;
	assign \g231990/_1_  = _w27201_ ;
	assign \g231991/_0_  = _w27217_ ;
	assign \g231992/_0_  = _w27233_ ;
	assign \g231995/_0_  = _w27236_ ;
	assign \g231998/_0_  = _w27240_ ;
	assign \g231999/_0_  = _w27246_ ;
	assign \g232002/_3_  = _w27253_ ;
	assign \g232035/u3_syn_4  = _w27260_ ;
	assign \g232038/u3_syn_4  = _w27265_ ;
	assign \g232046/u3_syn_4  = _w27269_ ;
	assign \g232054/u3_syn_4  = _w27273_ ;
	assign \g232062/u3_syn_4  = _w27276_ ;
	assign \g232070/u3_syn_4  = _w27278_ ;
	assign \g232078/u3_syn_4  = _w27284_ ;
	assign \g232079/u3_syn_4  = _w27287_ ;
	assign \g232087/u3_syn_4  = _w27290_ ;
	assign \g232096/u3_syn_4  = _w27292_ ;
	assign \g232104/u3_syn_4  = _w27295_ ;
	assign \g232112/u3_syn_4  = _w27297_ ;
	assign \g232120/u3_syn_4  = _w27301_ ;
	assign \g232128/u3_syn_4  = _w27304_ ;
	assign \g232136/u3_syn_4  = _w27308_ ;
	assign \g232144/u3_syn_4  = _w27311_ ;
	assign \g232152/u3_syn_4  = _w27314_ ;
	assign \g232161/u3_syn_4  = _w27317_ ;
	assign \g232169/u3_syn_4  = _w27319_ ;
	assign \g232177/u3_syn_4  = _w27322_ ;
	assign \g232185/u3_syn_4  = _w27323_ ;
	assign \g232186/u3_syn_4  = _w27327_ ;
	assign \g232194/u3_syn_4  = _w27330_ ;
	assign \g232202/u3_syn_4  = _w27332_ ;
	assign \g232210/u3_syn_4  = _w27335_ ;
	assign \g232218/u3_syn_4  = _w27338_ ;
	assign \g232226/u3_syn_4  = _w27340_ ;
	assign \g232234/u3_syn_4  = _w27343_ ;
	assign \g232242/u3_syn_4  = _w27345_ ;
	assign \g232251/u3_syn_4  = _w27348_ ;
	assign \g232259/u3_syn_4  = _w27350_ ;
	assign \g232267/u3_syn_4  = _w27353_ ;
	assign \g232275/u3_syn_4  = _w27355_ ;
	assign \g232283/u3_syn_4  = _w27357_ ;
	assign \g232291/u3_syn_4  = _w27359_ ;
	assign \g232299/u3_syn_4  = _w27361_ ;
	assign \g232307/u3_syn_4  = _w27363_ ;
	assign \g232315/u3_syn_4  = _w27365_ ;
	assign \g232324/u3_syn_4  = _w27367_ ;
	assign \g232332/u3_syn_4  = _w27369_ ;
	assign \g232341/u3_syn_4  = _w27371_ ;
	assign \g232349/u3_syn_4  = _w27373_ ;
	assign \g232357/u3_syn_4  = _w27375_ ;
	assign \g232366/u3_syn_4  = _w27377_ ;
	assign \g232374/u3_syn_4  = _w27379_ ;
	assign \g232382/u3_syn_4  = _w27381_ ;
	assign \g232390/u3_syn_4  = _w27383_ ;
	assign \g232398/u3_syn_4  = _w27385_ ;
	assign \g232406/u3_syn_4  = _w27387_ ;
	assign \g232414/u3_syn_4  = _w27389_ ;
	assign \g232422/u3_syn_4  = _w27391_ ;
	assign \g232427/u3_syn_4  = _w27392_ ;
	assign \g232431/u3_syn_4  = _w27394_ ;
	assign \g232439/u3_syn_4  = _w27396_ ;
	assign \g232444/u3_syn_4  = _w27397_ ;
	assign \g232452/u3_syn_4  = _w27399_ ;
	assign \g232461/u3_syn_4  = _w27400_ ;
	assign \g232471/u3_syn_4  = _w27402_ ;
	assign \g232479/u3_syn_4  = _w27404_ ;
	assign \g232487/u3_syn_4  = _w27405_ ;
	assign \g232495/u3_syn_4  = _w27406_ ;
	assign \g232503/u3_syn_4  = _w27408_ ;
	assign \g232506/u3_syn_4  = _w27409_ ;
	assign \g232514/u3_syn_4  = _w27411_ ;
	assign \g232527/u3_syn_4  = _w27412_ ;
	assign \g232530/u3_syn_4  = _w27415_ ;
	assign \g232536/u3_syn_4  = _w27416_ ;
	assign \g232544/u3_syn_4  = _w27419_ ;
	assign \g232551/u3_syn_4  = _w27420_ ;
	assign \g232557/u3_syn_4  = _w27422_ ;
	assign \g232568/u3_syn_4  = _w27424_ ;
	assign \g232576/u3_syn_4  = _w27426_ ;
	assign \g232585/u3_syn_4  = _w27427_ ;
	assign \g232593/u3_syn_4  = _w27428_ ;
	assign \g232597/u3_syn_4  = _w27430_ ;
	assign \g232609/u3_syn_4  = _w27432_ ;
	assign \g232617/u3_syn_4  = _w27434_ ;
	assign \g232625/u3_syn_4  = _w27436_ ;
	assign \g232633/u3_syn_4  = _w27438_ ;
	assign \g232641/u3_syn_4  = _w27440_ ;
	assign \g232649/u3_syn_4  = _w27442_ ;
	assign \g232657/u3_syn_4  = _w27444_ ;
	assign \g232665/u3_syn_4  = _w27446_ ;
	assign \g232673/u3_syn_4  = _w27448_ ;
	assign \g232681/u3_syn_4  = _w27450_ ;
	assign \g232689/u3_syn_4  = _w27451_ ;
	assign \g232697/u3_syn_4  = _w27452_ ;
	assign \g232705/u3_syn_4  = _w27454_ ;
	assign \g232713/u3_syn_4  = _w27455_ ;
	assign \g232717/u3_syn_4  = _w27457_ ;
	assign \g232729/u3_syn_4  = _w27459_ ;
	assign \g232737/u3_syn_4  = _w27460_ ;
	assign \g232745/u3_syn_4  = _w27462_ ;
	assign \g232749/u3_syn_4  = _w27463_ ;
	assign \g232761/u3_syn_4  = _w27464_ ;
	assign \g232768/u3_syn_4  = _w27466_ ;
	assign \g232777/u3_syn_4  = _w27468_ ;
	assign \g232785/u3_syn_4  = _w27470_ ;
	assign \g232793/u3_syn_4  = _w27472_ ;
	assign \g232801/u3_syn_4  = _w27474_ ;
	assign \g232809/u3_syn_4  = _w27476_ ;
	assign \g232815/u3_syn_4  = _w27477_ ;
	assign \g232823/u3_syn_4  = _w27479_ ;
	assign \g232833/u3_syn_4  = _w27480_ ;
	assign \g232841/u3_syn_4  = _w27482_ ;
	assign \g232846/u3_syn_4  = _w27483_ ;
	assign \g232851/u3_syn_4  = _w27485_ ;
	assign \g232865/u3_syn_4  = _w27486_ ;
	assign \g232873/u3_syn_4  = _w27487_ ;
	assign \g232881/u3_syn_4  = _w27488_ ;
	assign \g232882/u3_syn_4  = _w27491_ ;
	assign \g232895/u3_syn_4  = _w27492_ ;
	assign \g232904/u3_syn_4  = _w27493_ ;
	assign \g232913/u3_syn_4  = _w27494_ ;
	assign \g232921/u3_syn_4  = _w27495_ ;
	assign \g232928/u3_syn_4  = _w27496_ ;
	assign \g232934/u3_syn_4  = _w27497_ ;
	assign \g232945/u3_syn_4  = _w27498_ ;
	assign \g232953/u3_syn_4  = _w27499_ ;
	assign \g232954/u3_syn_4  = _w27500_ ;
	assign \g232969/u3_syn_4  = _w27501_ ;
	assign \g232977/u3_syn_4  = _w27502_ ;
	assign \g232981/u3_syn_4  = _w27503_ ;
	assign \g232993/u3_syn_4  = _w27504_ ;
	assign \g232995/u3_syn_4  = _w27505_ ;
	assign \g233009/u3_syn_4  = _w27506_ ;
	assign \g233017/u3_syn_4  = _w27507_ ;
	assign \g233025/u3_syn_4  = _w27508_ ;
	assign \g233033/u3_syn_4  = _w27509_ ;
	assign \g233041/u3_syn_4  = _w27510_ ;
	assign \g233047/u3_syn_4  = _w27511_ ;
	assign \g233057/u3_syn_4  = _w27512_ ;
	assign \g233065/u3_syn_4  = _w27513_ ;
	assign \g233073/u3_syn_4  = _w27514_ ;
	assign \g233081/u3_syn_4  = _w27515_ ;
	assign \g233087/u3_syn_4  = _w27516_ ;
	assign \g233097/u3_syn_4  = _w27517_ ;
	assign \g233105/u3_syn_4  = _w27518_ ;
	assign \g233113/u3_syn_4  = _w27519_ ;
	assign \g233121/u3_syn_4  = _w27520_ ;
	assign \g233128/u3_syn_4  = _w27521_ ;
	assign \g233134/u3_syn_4  = _w27522_ ;
	assign \g233144/u3_syn_4  = _w27523_ ;
	assign \g233153/u3_syn_4  = _w27524_ ;
	assign \g233161/u3_syn_4  = _w27525_ ;
	assign \g233169/u3_syn_4  = _w27526_ ;
	assign \g233177/u3_syn_4  = _w27527_ ;
	assign \g233185/u3_syn_4  = _w27528_ ;
	assign \g233193/u3_syn_4  = _w27529_ ;
	assign \g233201/u3_syn_4  = _w27530_ ;
	assign \g233209/u3_syn_4  = _w27531_ ;
	assign \g233217/u3_syn_4  = _w27532_ ;
	assign \g233219/u3_syn_4  = _w27533_ ;
	assign \g233229/u3_syn_4  = _w27534_ ;
	assign \g233241/u3_syn_4  = _w27535_ ;
	assign \g233249/u3_syn_4  = _w27536_ ;
	assign \g233257/u3_syn_4  = _w27537_ ;
	assign \g233265/u3_syn_4  = _w27538_ ;
	assign \g233273/u3_syn_4  = _w27539_ ;
	assign \g233281/u3_syn_4  = _w27540_ ;
	assign \g233289/u3_syn_4  = _w27541_ ;
	assign \g233297/u3_syn_4  = _w27542_ ;
	assign \g233305/u3_syn_4  = _w27543_ ;
	assign \g233313/u3_syn_4  = _w27544_ ;
	assign \g233321/u3_syn_4  = _w27545_ ;
	assign \g233329/u3_syn_4  = _w27546_ ;
	assign \g233337/u3_syn_4  = _w27547_ ;
	assign \g233345/u3_syn_4  = _w27548_ ;
	assign \g233353/u3_syn_4  = _w27549_ ;
	assign \g233361/u3_syn_4  = _w27550_ ;
	assign \g233369/u3_syn_4  = _w27551_ ;
	assign \g233377/u3_syn_4  = _w27552_ ;
	assign \g233382/u3_syn_4  = _w27553_ ;
	assign \g233392/u3_syn_4  = _w27554_ ;
	assign \g233394/u3_syn_4  = _w27555_ ;
	assign \g233409/u3_syn_4  = _w27556_ ;
	assign \g233417/u3_syn_4  = _w27557_ ;
	assign \g233425/u3_syn_4  = _w27558_ ;
	assign \g233433/u3_syn_4  = _w27559_ ;
	assign \g233441/u3_syn_4  = _w27560_ ;
	assign \g233449/u3_syn_4  = _w27561_ ;
	assign \g233453/u3_syn_4  = _w27562_ ;
	assign \g233465/u3_syn_4  = _w27563_ ;
	assign \g233473/u3_syn_4  = _w27564_ ;
	assign \g233481/u3_syn_4  = _w27565_ ;
	assign \g233489/u3_syn_4  = _w27566_ ;
	assign \g233497/u3_syn_4  = _w27567_ ;
	assign \g233505/u3_syn_4  = _w27568_ ;
	assign \g233513/u3_syn_4  = _w27569_ ;
	assign \g233516/u3_syn_4  = _w27570_ ;
	assign \g233529/u3_syn_4  = _w27571_ ;
	assign \g233531/u3_syn_4  = _w27572_ ;
	assign \g233546/u3_syn_4  = _w27573_ ;
	assign \g233554/u3_syn_4  = _w27574_ ;
	assign \g233562/u3_syn_4  = _w27575_ ;
	assign \g233570/u3_syn_4  = _w27576_ ;
	assign \g233578/u3_syn_4  = _w27577_ ;
	assign \g233586/u3_syn_4  = _w27578_ ;
	assign \g233594/u3_syn_4  = _w27579_ ;
	assign \g233602/u3_syn_4  = _w27580_ ;
	assign \g233603/u3_syn_4  = _w27581_ ;
	assign \g233618/u3_syn_4  = _w27582_ ;
	assign \g233626/u3_syn_4  = _w27583_ ;
	assign \g233634/u3_syn_4  = _w27584_ ;
	assign \g233642/u3_syn_4  = _w27585_ ;
	assign \g233650/u3_syn_4  = _w27586_ ;
	assign \g233658/u3_syn_4  = _w27587_ ;
	assign \g233666/u3_syn_4  = _w27588_ ;
	assign \g233674/u3_syn_4  = _w27589_ ;
	assign \g233682/u3_syn_4  = _w27590_ ;
	assign \g233690/u3_syn_4  = _w27591_ ;
	assign \g233698/u3_syn_4  = _w27592_ ;
	assign \g233706/u3_syn_4  = _w27593_ ;
	assign \g233714/u3_syn_4  = _w27594_ ;
	assign \g233722/u3_syn_4  = _w27595_ ;
	assign \g233730/u3_syn_4  = _w27596_ ;
	assign \g233738/u3_syn_4  = _w27597_ ;
	assign \g233746/u3_syn_4  = _w27598_ ;
	assign \g233754/u3_syn_4  = _w27599_ ;
	assign \g233762/u3_syn_4  = _w27600_ ;
	assign \g233770/u3_syn_4  = _w27601_ ;
	assign \g233778/u3_syn_4  = _w27602_ ;
	assign \g233783/u3_syn_4  = _w27603_ ;
	assign \g233794/u3_syn_4  = _w27604_ ;
	assign \g233802/u3_syn_4  = _w27605_ ;
	assign \g233806/u3_syn_4  = _w27606_ ;
	assign \g233818/u3_syn_4  = _w27607_ ;
	assign \g233826/u3_syn_4  = _w27608_ ;
	assign \g233828/u3_syn_4  = _w27609_ ;
	assign \g233838/u3_syn_4  = _w27610_ ;
	assign \g233850/u3_syn_4  = _w27611_ ;
	assign \g233858/u3_syn_4  = _w27612_ ;
	assign \g233860/u3_syn_4  = _w27613_ ;
	assign \g233870/u3_syn_4  = _w27614_ ;
	assign \g233881/u3_syn_4  = _w27615_ ;
	assign \g233890/u3_syn_4  = _w27616_ ;
	assign \g233899/u3_syn_4  = _w27617_ ;
	assign \g233908/u3_syn_4  = _w27618_ ;
	assign \g233917/u3_syn_4  = _w27619_ ;
	assign \g233919/u3_syn_4  = _w27620_ ;
	assign \g233927/u3_syn_4  = _w27621_ ;
	assign \g233935/u3_syn_4  = _w27622_ ;
	assign \g233943/u3_syn_4  = _w27623_ ;
	assign \g233945/u3_syn_4  = _w27624_ ;
	assign \g233953/u3_syn_4  = _w27625_ ;
	assign \g233961/u3_syn_4  = _w27626_ ;
	assign \g233969/u3_syn_4  = _w27627_ ;
	assign \g233977/u3_syn_4  = _w27628_ ;
	assign \g233985/u3_syn_4  = _w27629_ ;
	assign \g233993/u3_syn_4  = _w27630_ ;
	assign \g234001/u3_syn_4  = _w27631_ ;
	assign \g234008/u3_syn_4  = _w27632_ ;
	assign \g234009/u3_syn_4  = _w27633_ ;
	assign \g234024/u3_syn_4  = _w27634_ ;
	assign \g234032/u3_syn_4  = _w27635_ ;
	assign \g234038/u3_syn_4  = _w27636_ ;
	assign \g234056/u3_syn_4  = _w27637_ ;
	assign \g234063/u3_syn_4  = _w27638_ ;
	assign \g234071/u3_syn_4  = _w27639_ ;
	assign \g234079/u3_syn_4  = _w27640_ ;
	assign \g234098/u3_syn_4  = _w27641_ ;
	assign \g234106/u3_syn_4  = _w27642_ ;
	assign \g234114/u3_syn_4  = _w27643_ ;
	assign \g234122/u3_syn_4  = _w27644_ ;
	assign \g234130/u3_syn_4  = _w27645_ ;
	assign \g234138/u3_syn_4  = _w27646_ ;
	assign \g234145/u3_syn_4  = _w27647_ ;
	assign \g234156/u3_syn_4  = _w27648_ ;
	assign \g234162/u3_syn_4  = _w27649_ ;
	assign \g234171/u3_syn_4  = _w27650_ ;
	assign \g234183/u3_syn_4  = _w27651_ ;
	assign \g234248/u3_syn_4  = _w27652_ ;
	assign \g234265/u3_syn_4  = _w27653_ ;
	assign \g234273/u3_syn_4  = _w27654_ ;
	assign \g234281/u3_syn_4  = _w27655_ ;
	assign \g234289/u3_syn_4  = _w27656_ ;
	assign \g234297/u3_syn_4  = _w27657_ ;
	assign \g234306/u3_syn_4  = _w27658_ ;
	assign \g234314/u3_syn_4  = _w27659_ ;
	assign \g234322/u3_syn_4  = _w27660_ ;
	assign \g234331/u3_syn_4  = _w27661_ ;
	assign \g234339/u3_syn_4  = _w27662_ ;
	assign \g234347/u3_syn_4  = _w27663_ ;
	assign \g234355/u3_syn_4  = _w27664_ ;
	assign \g234363/u3_syn_4  = _w27665_ ;
	assign \g234371/u3_syn_4  = _w27666_ ;
	assign \g234379/u3_syn_4  = _w27667_ ;
	assign \g234387/u3_syn_4  = _w27668_ ;
	assign \g234395/u3_syn_4  = _w27669_ ;
	assign \g234403/u3_syn_4  = _w27670_ ;
	assign \g234411/u3_syn_4  = _w27671_ ;
	assign \g234419/u3_syn_4  = _w27672_ ;
	assign \g234427/u3_syn_4  = _w27673_ ;
	assign \g234435/u3_syn_4  = _w27674_ ;
	assign \g234443/u3_syn_4  = _w27675_ ;
	assign \g234451/u3_syn_4  = _w27676_ ;
	assign \g234459/u3_syn_4  = _w27677_ ;
	assign \g234467/u3_syn_4  = _w27678_ ;
	assign \g234475/u3_syn_4  = _w27679_ ;
	assign \g234483/u3_syn_4  = _w27680_ ;
	assign \g234491/u3_syn_4  = _w27681_ ;
	assign \g234499/u3_syn_4  = _w27682_ ;
	assign \g234507/u3_syn_4  = _w27683_ ;
	assign \g234515/u3_syn_4  = _w27684_ ;
	assign \g234523/u3_syn_4  = _w27685_ ;
	assign \g234531/u3_syn_4  = _w27686_ ;
	assign \g234539/u3_syn_4  = _w27687_ ;
	assign \g234547/u3_syn_4  = _w27688_ ;
	assign \g234555/u3_syn_4  = _w27689_ ;
	assign \g234563/u3_syn_4  = _w27690_ ;
	assign \g234571/u3_syn_4  = _w27691_ ;
	assign \g234579/u3_syn_4  = _w27692_ ;
	assign \g234587/u3_syn_4  = _w27693_ ;
	assign \g234595/u3_syn_4  = _w27694_ ;
	assign \g234604/u3_syn_4  = _w27695_ ;
	assign \g234612/u3_syn_4  = _w27696_ ;
	assign \g234620/u3_syn_4  = _w27697_ ;
	assign \g234628/u3_syn_4  = _w27698_ ;
	assign \g234636/u3_syn_4  = _w27699_ ;
	assign \g234644/u3_syn_4  = _w27700_ ;
	assign \g234652/u3_syn_4  = _w27701_ ;
	assign \g234660/u3_syn_4  = _w27702_ ;
	assign \g234668/u3_syn_4  = _w27703_ ;
	assign \g234676/u3_syn_4  = _w27704_ ;
	assign \g234684/u3_syn_4  = _w27705_ ;
	assign \g234692/u3_syn_4  = _w27706_ ;
	assign \g234700/u3_syn_4  = _w27707_ ;
	assign \g234708/u3_syn_4  = _w27708_ ;
	assign \g234716/u3_syn_4  = _w27709_ ;
	assign \g234725/u3_syn_4  = _w27710_ ;
	assign \g234733/u3_syn_4  = _w27711_ ;
	assign \g234741/u3_syn_4  = _w27712_ ;
	assign \g234749/u3_syn_4  = _w27713_ ;
	assign \g234757/u3_syn_4  = _w27714_ ;
	assign \g234765/u3_syn_4  = _w27715_ ;
	assign \g234773/u3_syn_4  = _w27716_ ;
	assign \g234781/u3_syn_4  = _w27717_ ;
	assign \g234789/u3_syn_4  = _w27718_ ;
	assign \g234798/u3_syn_4  = _w27719_ ;
	assign \g234806/u3_syn_4  = _w27720_ ;
	assign \g234814/u3_syn_4  = _w27721_ ;
	assign \g234822/u3_syn_4  = _w27722_ ;
	assign \g234830/u3_syn_4  = _w27723_ ;
	assign \g234838/u3_syn_4  = _w27724_ ;
	assign \g235911/u3_syn_4  = _w27726_ ;
	assign \g235912/u3_syn_4  = _w27728_ ;
	assign \g235920/u3_syn_4  = _w27730_ ;
	assign \g235928/u3_syn_4  = _w27732_ ;
	assign \g235936/u3_syn_4  = _w27734_ ;
	assign \g235944/u3_syn_4  = _w27736_ ;
	assign \g235952/u3_syn_4  = _w27738_ ;
	assign \g235960/u3_syn_4  = _w27740_ ;
	assign \g235968/u3_syn_4  = _w27742_ ;
	assign \g235976/u3_syn_4  = _w27744_ ;
	assign \g235984/u3_syn_4  = _w27746_ ;
	assign \g235992/u3_syn_4  = _w27748_ ;
	assign \g236000/u3_syn_4  = _w27749_ ;
	assign \g236008/u3_syn_4  = _w27751_ ;
	assign \g236016/u3_syn_4  = _w27753_ ;
	assign \g236021/u3_syn_4  = _w27755_ ;
	assign \g236025/u3_syn_4  = _w27757_ ;
	assign \g236033/u3_syn_4  = _w27759_ ;
	assign \g236041/u3_syn_4  = _w27761_ ;
	assign \g236049/u3_syn_4  = _w27763_ ;
	assign \g236057/u3_syn_4  = _w27765_ ;
	assign \g236065/u3_syn_4  = _w27767_ ;
	assign \g236073/u3_syn_4  = _w27769_ ;
	assign \g236081/u3_syn_4  = _w27771_ ;
	assign \g236089/u3_syn_4  = _w27773_ ;
	assign \g236097/u3_syn_4  = _w27775_ ;
	assign \g236105/u3_syn_4  = _w27777_ ;
	assign \g236113/u3_syn_4  = _w27779_ ;
	assign \g236121/u3_syn_4  = _w27781_ ;
	assign \g236129/u3_syn_4  = _w27783_ ;
	assign \g236137/u3_syn_4  = _w27785_ ;
	assign \g236145/u3_syn_4  = _w27787_ ;
	assign \g236153/u3_syn_4  = _w27789_ ;
	assign \g236161/u3_syn_4  = _w27791_ ;
	assign \g236169/u3_syn_4  = _w27793_ ;
	assign \g236177/u3_syn_4  = _w27795_ ;
	assign \g236185/u3_syn_4  = _w27797_ ;
	assign \g236193/u3_syn_4  = _w27799_ ;
	assign \g236196/u3_syn_4  = _w27800_ ;
	assign \g236198/u3_syn_4  = _w27801_ ;
	assign \g236203/u3_syn_4  = _w27803_ ;
	assign \g236211/u3_syn_4  = _w27805_ ;
	assign \g236219/u3_syn_4  = _w27806_ ;
	assign \g236220/u3_syn_4  = _w27808_ ;
	assign \g236229/u3_syn_4  = _w27810_ ;
	assign \g236232/u3_syn_4  = _w27811_ ;
	assign \g236238/u3_syn_4  = _w27813_ ;
	assign \g236246/u3_syn_4  = _w27815_ ;
	assign \g236255/u3_syn_4  = _w27817_ ;
	assign \g236263/u3_syn_4  = _w27819_ ;
	assign \g236271/u3_syn_4  = _w27821_ ;
	assign \g236275/u3_syn_4  = _w27822_ ;
	assign \g236280/u3_syn_4  = _w27824_ ;
	assign \g236288/u3_syn_4  = _w27826_ ;
	assign \g236296/u3_syn_4  = _w27828_ ;
	assign \g236304/u3_syn_4  = _w27829_ ;
	assign \g236305/u3_syn_4  = _w27830_ ;
	assign \g236306/u3_syn_4  = _w27832_ ;
	assign \g236315/u3_syn_4  = _w27834_ ;
	assign \g236323/u3_syn_4  = _w27836_ ;
	assign \g236331/u3_syn_4  = _w27838_ ;
	assign \g236334/u3_syn_4  = _w27839_ ;
	assign \g236340/u3_syn_4  = _w27841_ ;
	assign \g236348/u3_syn_4  = _w27843_ ;
	assign \g236357/u3_syn_4  = _w27844_ ;
	assign \g236359/u3_syn_4  = _w27846_ ;
	assign \g236367/u3_syn_4  = _w27848_ ;
	assign \g236374/u3_syn_4  = _w27849_ ;
	assign \g236376/u3_syn_4  = _w27851_ ;
	assign \g236377/u3_syn_4  = _w27853_ ;
	assign \g236385/u3_syn_4  = _w27855_ ;
	assign \g236393/u3_syn_4  = _w27857_ ;
	assign \g236402/u3_syn_4  = _w27859_ ;
	assign \g236410/u3_syn_4  = _w27861_ ;
	assign \g236419/u3_syn_4  = _w27863_ ;
	assign \g236427/u3_syn_4  = _w27865_ ;
	assign \g236433/u3_syn_4  = _w27866_ ;
	assign \g236436/u3_syn_4  = _w27868_ ;
	assign \g236444/u3_syn_4  = _w27870_ ;
	assign \g236452/u3_syn_4  = _w27872_ ;
	assign \g236460/u3_syn_4  = _w27874_ ;
	assign \g236468/u3_syn_4  = _w27876_ ;
	assign \g236476/u3_syn_4  = _w27878_ ;
	assign \g236484/u3_syn_4  = _w27880_ ;
	assign \g236492/u3_syn_4  = _w27882_ ;
	assign \g236500/u3_syn_4  = _w27884_ ;
	assign \g236508/u3_syn_4  = _w27886_ ;
	assign \g236516/u3_syn_4  = _w27888_ ;
	assign \g236518/u3_syn_4  = _w27889_ ;
	assign \g236525/u3_syn_4  = _w27891_ ;
	assign \g236533/u3_syn_4  = _w27893_ ;
	assign \g236542/u3_syn_4  = _w27895_ ;
	assign \g236550/u3_syn_4  = _w27897_ ;
	assign \g236559/u3_syn_4  = _w27899_ ;
	assign \g236567/u3_syn_4  = _w27901_ ;
	assign \g236575/u3_syn_4  = _w27903_ ;
	assign \g236583/u3_syn_4  = _w27905_ ;
	assign \g236591/u3_syn_4  = _w27907_ ;
	assign \g236599/u3_syn_4  = _w27909_ ;
	assign \g236607/u3_syn_4  = _w27911_ ;
	assign \g236608/u3_syn_4  = _w27913_ ;
	assign \g236616/u3_syn_4  = _w27915_ ;
	assign \g236624/u3_syn_4  = _w27917_ ;
	assign \g236632/u3_syn_4  = _w27919_ ;
	assign \g236640/u3_syn_4  = _w27921_ ;
	assign \g236647/u3_syn_4  = _w27922_ ;
	assign \g236649/u3_syn_4  = _w27924_ ;
	assign \g236659/u3_syn_4  = _w27926_ ;
	assign \g236671/u3_syn_4  = _w27928_ ;
	assign \g236677/u3_syn_4  = _w27929_ ;
	assign \g236688/u3_syn_4  = _w27931_ ;
	assign \g236696/u3_syn_4  = _w27933_ ;
	assign \g236705/u3_syn_4  = _w27935_ ;
	assign \g236712/u3_syn_4  = _w27936_ ;
	assign \g236718/u3_syn_4  = _w27938_ ;
	assign \g236729/u3_syn_4  = _w27939_ ;
	assign \g236732/u3_syn_4  = _w27941_ ;
	assign \g236745/u3_syn_4  = _w27943_ ;
	assign \g236753/u3_syn_4  = _w27945_ ;
	assign \g236761/u3_syn_4  = _w27947_ ;
	assign \g236769/u3_syn_4  = _w27949_ ;
	assign \g236777/u3_syn_4  = _w27951_ ;
	assign \g236779/u3_syn_4  = _w27952_ ;
	assign \g236788/u3_syn_4  = _w27954_ ;
	assign \g236800/u3_syn_4  = _w27956_ ;
	assign \g236802/u3_syn_4  = _w27958_ ;
	assign \g236805/u3_syn_4  = _w27959_ ;
	assign \g236813/u3_syn_4  = _w27961_ ;
	assign \g236825/u3_syn_4  = _w27963_ ;
	assign \g236829/u3_syn_4  = _w27964_ ;
	assign \g236837/u3_syn_4  = _w27966_ ;
	assign \g236849/u3_syn_4  = _w27968_ ;
	assign \g236854/u3_syn_4  = _w27969_ ;
	assign \g236860/u3_syn_4  = _w27971_ ;
	assign \g236872/u3_syn_4  = _w27973_ ;
	assign \g236878/u3_syn_4  = _w27974_ ;
	assign \g236884/u3_syn_4  = _w27976_ ;
	assign \g236896/u3_syn_4  = _w27978_ ;
	assign \g236903/u3_syn_4  = _w27979_ ;
	assign \g236908/u3_syn_4  = _w27981_ ;
	assign \g236920/u3_syn_4  = _w27983_ ;
	assign \g236930/u3_syn_4  = _w27985_ ;
	assign \g236939/u3_syn_4  = _w27987_ ;
	assign \g236947/u3_syn_4  = _w27989_ ;
	assign \g236949/u3_syn_4  = _w27990_ ;
	assign \g236956/u3_syn_4  = _w27992_ ;
	assign \g236962/u3_syn_4  = _w27993_ ;
	assign \g236965/u3_syn_4  = _w27995_ ;
	assign \g236980/u3_syn_4  = _w27997_ ;
	assign \g236988/u3_syn_4  = _w27998_ ;
	assign \g236989/u3_syn_4  = _w28000_ ;
	assign \g237004/u3_syn_4  = _w28002_ ;
	assign \g237005/u3_syn_4  = _w28003_ ;
	assign \g237020/u3_syn_4  = _w28004_ ;
	assign \g237021/u3_syn_4  = _w28006_ ;
	assign \g237033/u3_syn_4  = _w28008_ ;
	assign \g237044/u3_syn_4  = _w28009_ ;
	assign \g237045/u3_syn_4  = _w28011_ ;
	assign \g237056/u3_syn_4  = _w28013_ ;
	assign \g237068/u3_syn_4  = _w28015_ ;
	assign \g237076/u3_syn_4  = _w28017_ ;
	assign \g237084/u3_syn_4  = _w28019_ ;
	assign \g237092/u3_syn_4  = _w28020_ ;
	assign \g237095/u3_syn_4  = _w28022_ ;
	assign \g237107/u3_syn_4  = _w28024_ ;
	assign \g237110/u3_syn_4  = _w28025_ ;
	assign \g237119/u3_syn_4  = _w28027_ ;
	assign \g237131/u3_syn_4  = _w28029_ ;
	assign \g237135/u3_syn_4  = _w28030_ ;
	assign \g237148/u3_syn_4  = _w28031_ ;
	assign \g237152/u3_syn_4  = _w28032_ ;
	assign \g237165/u3_syn_4  = _w28033_ ;
	assign \g237168/u3_syn_4  = _w28035_ ;
	assign \g237180/u3_syn_4  = _w28037_ ;
	assign \g237185/u3_syn_4  = _w28038_ ;
	assign \g237192/u3_syn_4  = _w28040_ ;
	assign \g237204/u3_syn_4  = _w28042_ ;
	assign \g237209/u3_syn_4  = _w28043_ ;
	assign \g237215/u3_syn_4  = _w28045_ ;
	assign \g237229/u3_syn_4  = _w28046_ ;
	assign \g237231/u3_syn_4  = _w28048_ ;
	assign \g237245/u3_syn_4  = _w28049_ ;
	assign \g237251/u3_syn_4  = _w28051_ ;
	assign \g237260/u3_syn_4  = _w28052_ ;
	assign \g237262/u3_syn_4  = _w28054_ ;
	assign \g237277/u3_syn_4  = _w28055_ ;
	assign \g237281/u3_syn_4  = _w28057_ ;
	assign \g237293/u3_syn_4  = _w28058_ ;
	assign \g237294/u3_syn_4  = _w28060_ ;
	assign \g237310/u3_syn_4  = _w28061_ ;
	assign \g237311/u3_syn_4  = _w28063_ ;
	assign \g237323/u3_syn_4  = _w28065_ ;
	assign \g237334/u3_syn_4  = _w28067_ ;
	assign \g237342/u3_syn_4  = _w28068_ ;
	assign \g237350/u3_syn_4  = _w28070_ ;
	assign \g237353/u3_syn_4  = _w28071_ ;
	assign \g237359/u3_syn_4  = _w28073_ ;
	assign \g237367/u3_syn_4  = _w28075_ ;
	assign \g237368/u3_syn_4  = _w28076_ ;
	assign \g237378/u3_syn_4  = _w28078_ ;
	assign \g237391/u3_syn_4  = _w28080_ ;
	assign \g237392/u3_syn_4  = _w28081_ ;
	assign \g237403/u3_syn_4  = _w28083_ ;
	assign \g237415/u3_syn_4  = _w28085_ ;
	assign \g237417/u3_syn_4  = _w28086_ ;
	assign \g237431/u3_syn_4  = _w28088_ ;
	assign \g237439/u3_syn_4  = _w28090_ ;
	assign \g237440/u3_syn_4  = _w28091_ ;
	assign \g237454/u3_syn_4  = _w28093_ ;
	assign \g237457/u3_syn_4  = _w28094_ ;
	assign \g237472/u3_syn_4  = _w28096_ ;
	assign \g237480/u3_syn_4  = _w28097_ ;
	assign \g237488/u3_syn_4  = _w28099_ ;
	assign \g237496/u3_syn_4  = _w28100_ ;
	assign \g237499/u3_syn_4  = _w28101_ ;
	assign \g237512/u3_syn_4  = _w28102_ ;
	assign \g237515/u3_syn_4  = _w28104_ ;
	assign \g237525/u3_syn_4  = _w28106_ ;
	assign \g237529/u3_syn_4  = _w28107_ ;
	assign \g237535/u3_syn_4  = _w28109_ ;
	assign \g237541/u3_syn_4  = _w28110_ ;
	assign \g237553/u3_syn_4  = _w28112_ ;
	assign \g237561/u3_syn_4  = _w28113_ ;
	assign \g237569/u3_syn_4  = _w28115_ ;
	assign \g237575/u3_syn_4  = _w28116_ ;
	assign \g237578/u3_syn_4  = _w28117_ ;
	assign \g237581/u3_syn_4  = _w28118_ ;
	assign \g237591/u3_syn_4  = _w28120_ ;
	assign \g237602/u3_syn_4  = _w28122_ ;
	assign \g237610/u3_syn_4  = _w28124_ ;
	assign \g237617/u3_syn_4  = _w28125_ ;
	assign \g237623/u3_syn_4  = _w28126_ ;
	assign \g237633/u3_syn_4  = _w28127_ ;
	assign \g237635/u3_syn_4  = _w28128_ ;
	assign \g237648/u3_syn_4  = _w28129_ ;
	assign \g237658/u3_syn_4  = _w28130_ ;
	assign \g237659/u3_syn_4  = _w28131_ ;
	assign \g237660/u3_syn_4  = _w28132_ ;
	assign \g237668/u3_syn_4  = _w28133_ ;
	assign \g237675/u3_syn_4  = _w28134_ ;
	assign \g237684/u3_syn_4  = _w28135_ ;
	assign \g237692/u3_syn_4  = _w28136_ ;
	assign \g237693/u3_syn_4  = _w28137_ ;
	assign \g237705/u3_syn_4  = _w28138_ ;
	assign \g237716/u3_syn_4  = _w28139_ ;
	assign \g237717/u3_syn_4  = _w28140_ ;
	assign \g237729/u3_syn_4  = _w28141_ ;
	assign \g237740/u3_syn_4  = _w28142_ ;
	assign \g237741/u3_syn_4  = _w28143_ ;
	assign \g237756/u3_syn_4  = _w28144_ ;
	assign \g237764/u3_syn_4  = _w28145_ ;
	assign \g237768/u3_syn_4  = _w28146_ ;
	assign \g237780/u3_syn_4  = _w28147_ ;
	assign \g237782/u3_syn_4  = _w28148_ ;
	assign \g237792/u3_syn_4  = _w28149_ ;
	assign \g237804/u3_syn_4  = _w28150_ ;
	assign \g237812/u3_syn_4  = _w28151_ ;
	assign \g237820/u3_syn_4  = _w28152_ ;
	assign \g237828/u3_syn_4  = _w28153_ ;
	assign \g237836/u3_syn_4  = _w28154_ ;
	assign \g237844/u3_syn_4  = _w28155_ ;
	assign \g237852/u3_syn_4  = _w28156_ ;
	assign \g237860/u3_syn_4  = _w28157_ ;
	assign \g237868/u3_syn_4  = _w28158_ ;
	assign \g237876/u3_syn_4  = _w28159_ ;
	assign \g237884/u3_syn_4  = _w28160_ ;
	assign \g237888/u3_syn_4  = _w28161_ ;
	assign \g237895/u3_syn_4  = _w28162_ ;
	assign \g237907/u3_syn_4  = _w28163_ ;
	assign \g237916/u3_syn_4  = _w28164_ ;
	assign \g237924/u3_syn_4  = _w28165_ ;
	assign \g237931/u3_syn_4  = _w28166_ ;
	assign \g237940/u3_syn_4  = _w28167_ ;
	assign \g237949/u3_syn_4  = _w28168_ ;
	assign \g237950/u3_syn_4  = _w28169_ ;
	assign \g237955/u3_syn_4  = _w28170_ ;
	assign \g237961/u3_syn_4  = _w28171_ ;
	assign \g237965/u3_syn_4  = _w28172_ ;
	assign \g237975/u3_syn_4  = _w28173_ ;
	assign \g237983/u3_syn_4  = _w28174_ ;
	assign \g237989/u3_syn_4  = _w28175_ ;
	assign \g237999/u3_syn_4  = _w28176_ ;
	assign \g238007/u3_syn_4  = _w28177_ ;
	assign \g238015/u3_syn_4  = _w28178_ ;
	assign \g238017/u3_syn_4  = _w28179_ ;
	assign \g238033/u3_syn_4  = _w28180_ ;
	assign \g238035/u3_syn_4  = _w28181_ ;
	assign \g238049/u3_syn_4  = _w28182_ ;
	assign \g238057/u3_syn_4  = _w28183_ ;
	assign \g238065/u3_syn_4  = _w28184_ ;
	assign \g238072/u3_syn_4  = _w28185_ ;
	assign \g238081/u3_syn_4  = _w28186_ ;
	assign \g238082/u3_syn_4  = _w28187_ ;
	assign \g238097/u3_syn_4  = _w28188_ ;
	assign \g238105/u3_syn_4  = _w28189_ ;
	assign \g238113/u3_syn_4  = _w28190_ ;
	assign \g238114/u3_syn_4  = _w28191_ ;
	assign \g238129/u3_syn_4  = _w28192_ ;
	assign \g238137/u3_syn_4  = _w28193_ ;
	assign \g238145/u3_syn_4  = _w28194_ ;
	assign \g238153/u3_syn_4  = _w28195_ ;
	assign \g238161/u3_syn_4  = _w28196_ ;
	assign \g238163/u3_syn_4  = _w28197_ ;
	assign \g238177/u3_syn_4  = _w28198_ ;
	assign \g238179/u3_syn_4  = _w28199_ ;
	assign \g238194/u3_syn_4  = _w28200_ ;
	assign \g238197/u3_syn_4  = _w28201_ ;
	assign \g238209/u3_syn_4  = _w28202_ ;
	assign \g238213/u3_syn_4  = _w28203_ ;
	assign \g238225/u3_syn_4  = _w28204_ ;
	assign \g238229/u3_syn_4  = _w28205_ ;
	assign \g238237/u3_syn_4  = _w28206_ ;
	assign \g238250/u3_syn_4  = _w28207_ ;
	assign \g238257/u3_syn_4  = _w28208_ ;
	assign \g238263/u3_syn_4  = _w28209_ ;
	assign \g238269/u3_syn_4  = _w28210_ ;
	assign \g238282/u3_syn_4  = _w28211_ ;
	assign \g238285/u3_syn_4  = _w28212_ ;
	assign \g238298/u3_syn_4  = _w28213_ ;
	assign \g238301/u3_syn_4  = _w28214_ ;
	assign \g238314/u3_syn_4  = _w28215_ ;
	assign \g238316/u3_syn_4  = _w28216_ ;
	assign \g238329/u3_syn_4  = _w28217_ ;
	assign \g238338/u3_syn_4  = _w28218_ ;
	assign \g238346/u3_syn_4  = _w28219_ ;
	assign \g238351/u3_syn_4  = _w28220_ ;
	assign \g238356/u3_syn_4  = _w28221_ ;
	assign \g238368/u3_syn_4  = _w28222_ ;
	assign \g238378/u3_syn_4  = _w28223_ ;
	assign \g238386/u3_syn_4  = _w28224_ ;
	assign \g238394/u3_syn_4  = _w28225_ ;
	assign \g238402/u3_syn_4  = _w28226_ ;
	assign \g238409/u3_syn_4  = _w28227_ ;
	assign \g238412/u3_syn_4  = _w28228_ ;
	assign \g238427/u3_syn_4  = _w28229_ ;
	assign \g238429/u3_syn_4  = _w28230_ ;
	assign \g238443/u3_syn_4  = _w28231_ ;
	assign \g238448/u3_syn_4  = _w28232_ ;
	assign \g238457/u3_syn_4  = _w28233_ ;
	assign \g238460/u3_syn_4  = _w28234_ ;
	assign \g238472/u3_syn_4  = _w28235_ ;
	assign \g238484/u3_syn_4  = _w28236_ ;
	assign \g238492/u3_syn_4  = _w28237_ ;
	assign \g238500/u3_syn_4  = _w28238_ ;
	assign \g238505/u3_syn_4  = _w28239_ ;
	assign \g238516/u3_syn_4  = _w28240_ ;
	assign \g238524/u3_syn_4  = _w28241_ ;
	assign \g238532/u3_syn_4  = _w28242_ ;
	assign \g238534/u3_syn_4  = _w28243_ ;
	assign \g238544/u3_syn_4  = _w28244_ ;
	assign \g238549/u3_syn_4  = _w28245_ ;
	assign \g238550/u3_syn_4  = _w28246_ ;
	assign \g238565/u3_syn_4  = _w28247_ ;
	assign \g238566/u3_syn_4  = _w28248_ ;
	assign \g238582/u3_syn_4  = _w28249_ ;
	assign \g238583/u3_syn_4  = _w28250_ ;
	assign \g238594/u3_syn_4  = _w28251_ ;
	assign \g238606/u3_syn_4  = _w28252_ ;
	assign \g238614/u3_syn_4  = _w28253_ ;
	assign \g238615/u3_syn_4  = _w28254_ ;
	assign \g238619/u3_syn_4  = _w28255_ ;
	assign \g238631/u3_syn_4  = _w28256_ ;
	assign \g238639/u3_syn_4  = _w28257_ ;
	assign \g238647/u3_syn_4  = _w28258_ ;
	assign \g238649/u3_syn_4  = _w28259_ ;
	assign \g238659/u3_syn_4  = _w28260_ ;
	assign \g238670/u3_syn_4  = _w28261_ ;
	assign \g238671/u3_syn_4  = _w28262_ ;
	assign \g238680/u3_syn_4  = _w28263_ ;
	assign \g238688/u3_syn_4  = _w28264_ ;
	assign \g238691/u3_syn_4  = _w28265_ ;
	assign \g238696/u3_syn_4  = _w28266_ ;
	assign \g238705/u3_syn_4  = _w28267_ ;
	assign \g238708/u3_syn_4  = _w28268_ ;
	assign \g238721/u3_syn_4  = _w28269_ ;
	assign \g238724/u3_syn_4  = _w28270_ ;
	assign \g238736/u3_syn_4  = _w28271_ ;
	assign \g238745/u3_syn_4  = _w28272_ ;
	assign \g238753/u3_syn_4  = _w28273_ ;
	assign \g238757/u3_syn_4  = _w28274_ ;
	assign \g238764/u3_syn_4  = _w28275_ ;
	assign \g238776/u3_syn_4  = _w28276_ ;
	assign \g238781/u3_syn_4  = _w28277_ ;
	assign \g238787/u3_syn_4  = _w28278_ ;
	assign \g238799/u3_syn_4  = _w28279_ ;
	assign \g238807/u3_syn_4  = _w28280_ ;
	assign \g238811/u3_syn_4  = _w28281_ ;
	assign \g238824/u3_syn_4  = _w28282_ ;
	assign \g238830/u3_syn_4  = _w28283_ ;
	assign \g238841/u3_syn_4  = _w28284_ ;
	assign \g238843/u3_syn_4  = _w28285_ ;
	assign \g238855/u3_syn_4  = _w28286_ ;
	assign \g238859/u3_syn_4  = _w28287_ ;
	assign \g238863/u3_syn_4  = _w28288_ ;
	assign \g238868/u3_syn_4  = _w28289_ ;
	assign \g238880/u3_syn_4  = _w28290_ ;
	assign \g238888/u3_syn_4  = _w28291_ ;
	assign \g238892/u3_syn_4  = _w28292_ ;
	assign \g238903/u3_syn_4  = _w28293_ ;
	assign \g238911/u3_syn_4  = _w28294_ ;
	assign \g238915/u3_syn_4  = _w28295_ ;
	assign \g238927/u3_syn_4  = _w28296_ ;
	assign \g238937/u3_syn_4  = _w28297_ ;
	assign \g238945/u3_syn_4  = _w28298_ ;
	assign \g238953/u3_syn_4  = _w28299_ ;
	assign \g238961/u3_syn_4  = _w28300_ ;
	assign \g238970/u3_syn_4  = _w28301_ ;
	assign \g238971/u3_syn_4  = _w28302_ ;
	assign \g238983/u3_syn_4  = _w28303_ ;
	assign \g238994/u3_syn_4  = _w28304_ ;
	assign \g239002/u3_syn_4  = _w28305_ ;
	assign \g239009/u3_syn_4  = _w28306_ ;
	assign \g239015/u3_syn_4  = _w28307_ ;
	assign \g239025/u3_syn_4  = _w28308_ ;
	assign \g239030/u3_syn_4  = _w28309_ ;
	assign \g239041/u3_syn_4  = _w28310_ ;
	assign \g239048/u3_syn_4  = _w28311_ ;
	assign \g239053/u3_syn_4  = _w28312_ ;
	assign \g239065/u3_syn_4  = _w28313_ ;
	assign \g239073/u3_syn_4  = _w28314_ ;
	assign \g239081/u3_syn_4  = _w28315_ ;
	assign \g239082/u3_syn_4  = _w28316_ ;
	assign \g239093/u3_syn_4  = _w28317_ ;
	assign \g239105/u3_syn_4  = _w28318_ ;
	assign \g239108/u3_syn_4  = _w28319_ ;
	assign \g239117/u3_syn_4  = _w28320_ ;
	assign \g239129/u3_syn_4  = _w28321_ ;
	assign \g239137/u3_syn_4  = _w28322_ ;
	assign \g239139/u3_syn_4  = _w28323_ ;
	assign \g239148/u3_syn_4  = _w28324_ ;
	assign \g239160/u3_syn_4  = _w28325_ ;
	assign \g239162/u3_syn_4  = _w28326_ ;
	assign \g239172/u3_syn_4  = _w28327_ ;
	assign \g239184/u3_syn_4  = _w28328_ ;
	assign \g239187/u3_syn_4  = _w28329_ ;
	assign \g239189/u3_syn_4  = _w28330_ ;
	assign \g239201/u3_syn_4  = _w28331_ ;
	assign \g239208/u3_syn_4  = _w28332_ ;
	assign \g239217/u3_syn_4  = _w28333_ ;
	assign \g239219/u3_syn_4  = _w28334_ ;
	assign \g239226/u3_syn_4  = _w28335_ ;
	assign \g239234/u3_syn_4  = _w28336_ ;
	assign \g239242/u3_syn_4  = _w28337_ ;
	assign \g239246/u3_syn_4  = _w28338_ ;
	assign \g239257/u3_syn_4  = _w28339_ ;
	assign \g239258/u3_syn_4  = _w28340_ ;
	assign \g239263/u3_syn_4  = _w28341_ ;
	assign \g239275/u3_syn_4  = _w28342_ ;
	assign \g239277/u3_syn_4  = _w28343_ ;
	assign \g239291/u3_syn_4  = _w28344_ ;
	assign \g239296/u3_syn_4  = _w28345_ ;
	assign \g239308/u3_syn_4  = _w28346_ ;
	assign \g239311/u3_syn_4  = _w28347_ ;
	assign \g239322/u3_syn_4  = _w28348_ ;
	assign \g239329/u3_syn_4  = _w28349_ ;
	assign \g239338/u3_syn_4  = _w28350_ ;
	assign \g239339/u3_syn_4  = _w28351_ ;
	assign \g239346/u3_syn_4  = _w28352_ ;
	assign \g239351/u3_syn_4  = _w28353_ ;
	assign \g239363/u3_syn_4  = _w28354_ ;
	assign \g239370/u3_syn_4  = _w28355_ ;
	assign \g239375/u3_syn_4  = _w28356_ ;
	assign \g239387/u3_syn_4  = _w28357_ ;
	assign \g239395/u3_syn_4  = _w28358_ ;
	assign \g239418/u3_syn_4  = _w28359_ ;
	assign \g239439/u3_syn_4  = _w28360_ ;
	assign \g239442/u3_syn_4  = _w28361_ ;
	assign \g239454/u3_syn_4  = _w28362_ ;
	assign \g239464/u3_syn_4  = _w28363_ ;
	assign \g239470/u3_syn_4  = _w28364_ ;
	assign \g239481/u3_syn_4  = _w28365_ ;
	assign \g239487/u3_syn_4  = _w28366_ ;
	assign \g239497/u3_syn_4  = _w28367_ ;
	assign \g239520/u3_syn_4  = _w28368_ ;
	assign \g239532/u3_syn_4  = _w28369_ ;
	assign \g239543/u3_syn_4  = _w28370_ ;
	assign \g239551/u3_syn_4  = _w28371_ ;
	assign \g239552/u3_syn_4  = _w28372_ ;
	assign \g239567/u3_syn_4  = _w28373_ ;
	assign \g239575/u3_syn_4  = _w28374_ ;
	assign \g239579/u3_syn_4  = _w28375_ ;
	assign \g239592/u3_syn_4  = _w28376_ ;
	assign \g239594/u3_syn_4  = _w28377_ ;
	assign \g239608/u3_syn_4  = _w28378_ ;
	assign \g239626/u3_syn_4  = _w28379_ ;
	assign \g239634/u3_syn_4  = _w28380_ ;
	assign \g239646/u3_syn_4  = _w28381_ ;
	assign \g239649/u3_syn_4  = _w28382_ ;
	assign \g239657/u3_syn_4  = _w28383_ ;
	assign \g239670/u3_syn_4  = _w28384_ ;
	assign \g239673/u3_syn_4  = _w28385_ ;
	assign \g239686/u3_syn_4  = _w28386_ ;
	assign \g239694/u3_syn_4  = _w28387_ ;
	assign \g239695/u3_syn_4  = _w28388_ ;
	assign \g239701/u3_syn_4  = _w28389_ ;
	assign \g239705/u3_syn_4  = _w28390_ ;
	assign \g239709/u3_syn_4  = _w28391_ ;
	assign \g239715/u3_syn_4  = _w28392_ ;
	assign \g239717/u3_syn_4  = _w28393_ ;
	assign \g239726/u3_syn_4  = _w28394_ ;
	assign \g239734/u3_syn_4  = _w28395_ ;
	assign \g239735/u3_syn_4  = _w28396_ ;
	assign \g239743/u3_syn_4  = _w28397_ ;
	assign \g239760/u3_syn_4  = _w28398_ ;
	assign \g239768/u3_syn_4  = _w28399_ ;
	assign \g239776/u3_syn_4  = _w28400_ ;
	assign \g239784/u3_syn_4  = _w28401_ ;
	assign \g239793/u3_syn_4  = _w28402_ ;
	assign \g239801/u3_syn_4  = _w28403_ ;
	assign \g239817/u3_syn_4  = _w28404_ ;
	assign \g239818/u3_syn_4  = _w28405_ ;
	assign \g239848/u3_syn_4  = _w28406_ ;
	assign \g239856/u3_syn_4  = _w28407_ ;
	assign \g239872/u3_syn_4  = _w28408_ ;
	assign \g239880/u3_syn_4  = _w28409_ ;
	assign \g239888/u3_syn_4  = _w28410_ ;
	assign \g239896/u3_syn_4  = _w28411_ ;
	assign \g239904/u3_syn_4  = _w28412_ ;
	assign \g239912/u3_syn_4  = _w28413_ ;
	assign \g239920/u3_syn_4  = _w28414_ ;
	assign \g239928/u3_syn_4  = _w28415_ ;
	assign \g239936/u3_syn_4  = _w28416_ ;
	assign \g239951/u3_syn_4  = _w28417_ ;
	assign \g239963/u3_syn_4  = _w28418_ ;
	assign \g239979/u3_syn_4  = _w28419_ ;
	assign \g239986/u3_syn_4  = _w28420_ ;
	assign \g239999/u3_syn_4  = _w28421_ ;
	assign \g240000/u3_syn_4  = _w28422_ ;
	assign \g240008/u3_syn_4  = _w28423_ ;
	assign \g240012/u3_syn_4  = _w28424_ ;
	assign \g240018/u3_syn_4  = _w28425_ ;
	assign \g240026/u3_syn_4  = _w28426_ ;
	assign \g240034/u3_syn_4  = _w28427_ ;
	assign \g240042/u3_syn_4  = _w28428_ ;
	assign \g240050/u3_syn_4  = _w28429_ ;
	assign \g240074/u3_syn_4  = _w28430_ ;
	assign \g240091/u3_syn_4  = _w28431_ ;
	assign \g240122/u3_syn_4  = _w28432_ ;
	assign \g240147/u3_syn_4  = _w28433_ ;
	assign \g240209/u3_syn_4  = _w28434_ ;
	assign \g240219/u3_syn_4  = _w28435_ ;
	assign \g240259/u3_syn_4  = _w28436_ ;
	assign \g240334/u3_syn_4  = _w28437_ ;
	assign \g240406/u3_syn_4  = _w28438_ ;
	assign \g240416/u3_syn_4  = _w28439_ ;
	assign \g240424/u3_syn_4  = _w28440_ ;
	assign \g240432/u3_syn_4  = _w28441_ ;
	assign \g240440/u3_syn_4  = _w28442_ ;
	assign \g240448/u3_syn_4  = _w28443_ ;
	assign \g240456/u3_syn_4  = _w28444_ ;
	assign \g240464/u3_syn_4  = _w28445_ ;
	assign \g240472/u3_syn_4  = _w28446_ ;
	assign \g240480/u3_syn_4  = _w28447_ ;
	assign \g240488/u3_syn_4  = _w28448_ ;
	assign \g240496/u3_syn_4  = _w28449_ ;
	assign \g240504/u3_syn_4  = _w28450_ ;
	assign \g240512/u3_syn_4  = _w28451_ ;
	assign \g240520/u3_syn_4  = _w28452_ ;
	assign \g240530/u3_syn_4  = _w28453_ ;
	assign \g240538/u3_syn_4  = _w28454_ ;
	assign \g240547/u3_syn_4  = _w28455_ ;
	assign \g240555/u3_syn_4  = _w28456_ ;
	assign \g240563/u3_syn_4  = _w28457_ ;
	assign \g240571/u3_syn_4  = _w28458_ ;
	assign \g240579/u3_syn_4  = _w28459_ ;
	assign \g240587/u3_syn_4  = _w28460_ ;
	assign \g240595/u3_syn_4  = _w28461_ ;
	assign \g240603/u3_syn_4  = _w28462_ ;
	assign \g240611/u3_syn_4  = _w28463_ ;
	assign \g240619/u3_syn_4  = _w28464_ ;
	assign \g240627/u3_syn_4  = _w28465_ ;
	assign \g240635/u3_syn_4  = _w28466_ ;
	assign \g240643/u3_syn_4  = _w28467_ ;
	assign \g240651/u3_syn_4  = _w28468_ ;
	assign \g240659/u3_syn_4  = _w28469_ ;
	assign \g240667/u3_syn_4  = _w28470_ ;
	assign \g240675/u3_syn_4  = _w28471_ ;
	assign \g240683/u3_syn_4  = _w28472_ ;
	assign \g240691/u3_syn_4  = _w28473_ ;
	assign \g240699/u3_syn_4  = _w28474_ ;
	assign \g240707/u3_syn_4  = _w28475_ ;
	assign \g240715/u3_syn_4  = _w28476_ ;
	assign \g240723/u3_syn_4  = _w28477_ ;
	assign \g240731/u3_syn_4  = _w28478_ ;
	assign \g240739/u3_syn_4  = _w28479_ ;
	assign \g240747/u3_syn_4  = _w28480_ ;
	assign \g240755/u3_syn_4  = _w28481_ ;
	assign \g240763/u3_syn_4  = _w28482_ ;
	assign \g240771/u3_syn_4  = _w28483_ ;
	assign \g240779/u3_syn_4  = _w28484_ ;
	assign \g240787/u3_syn_4  = _w28485_ ;
	assign \g240795/u3_syn_4  = _w28486_ ;
	assign \g240803/u3_syn_4  = _w28487_ ;
	assign \g240811/u3_syn_4  = _w28488_ ;
	assign \g240819/u3_syn_4  = _w28489_ ;
	assign \g240827/u3_syn_4  = _w28490_ ;
	assign \g240835/u3_syn_4  = _w28491_ ;
	assign \g240843/u3_syn_4  = _w28492_ ;
	assign \g240851/u3_syn_4  = _w28493_ ;
	assign \g240859/u3_syn_4  = _w28494_ ;
	assign \g240867/u3_syn_4  = _w28495_ ;
	assign \g240875/u3_syn_4  = _w28496_ ;
	assign \g240883/u3_syn_4  = _w28497_ ;
	assign \g240891/u3_syn_4  = _w28498_ ;
	assign \g240899/u3_syn_4  = _w28499_ ;
	assign \g240907/u3_syn_4  = _w28500_ ;
	assign \g240915/u3_syn_4  = _w28501_ ;
	assign \g240923/u3_syn_4  = _w28502_ ;
	assign \g240931/u3_syn_4  = _w28503_ ;
	assign \g240939/u3_syn_4  = _w28504_ ;
	assign \g240947/u3_syn_4  = _w28505_ ;
	assign \g240955/u3_syn_4  = _w28506_ ;
	assign \g240963/u3_syn_4  = _w28507_ ;
	assign \g240971/u3_syn_4  = _w28508_ ;
	assign \g240979/u3_syn_4  = _w28509_ ;
	assign \g240987/u3_syn_4  = _w28510_ ;
	assign \g240995/u3_syn_4  = _w28511_ ;
	assign \g241003/u3_syn_4  = _w28512_ ;
	assign \g241011/u3_syn_4  = _w28513_ ;
	assign \g241019/u3_syn_4  = _w28514_ ;
	assign \g241027/u3_syn_4  = _w28515_ ;
	assign \g241036/u3_syn_4  = _w28516_ ;
	assign \g241044/u3_syn_4  = _w28517_ ;
	assign \g241052/u3_syn_4  = _w28518_ ;
	assign \g241060/u3_syn_4  = _w28519_ ;
	assign \g241068/u3_syn_4  = _w28520_ ;
	assign \g241076/u3_syn_4  = _w28521_ ;
	assign \g241084/u3_syn_4  = _w28522_ ;
	assign \g241092/u3_syn_4  = _w28523_ ;
	assign \g241100/u3_syn_4  = _w28524_ ;
	assign \g241108/u3_syn_4  = _w28525_ ;
	assign \g241116/u3_syn_4  = _w28526_ ;
	assign \g241124/u3_syn_4  = _w28527_ ;
	assign \g241132/u3_syn_4  = _w28528_ ;
	assign \g241140/u3_syn_4  = _w28529_ ;
	assign \g241148/u3_syn_4  = _w28530_ ;
	assign \g241156/u3_syn_4  = _w28531_ ;
	assign \g241164/u3_syn_4  = _w28532_ ;
	assign \g241172/u3_syn_4  = _w28533_ ;
	assign \g241180/u3_syn_4  = _w28534_ ;
	assign \g241188/u3_syn_4  = _w28535_ ;
	assign \g241196/u3_syn_4  = _w28536_ ;
	assign \g241205/u3_syn_4  = _w28537_ ;
	assign \g241213/u3_syn_4  = _w28538_ ;
	assign \g241221/u3_syn_4  = _w28539_ ;
	assign \g241229/u3_syn_4  = _w28540_ ;
	assign \g241237/u3_syn_4  = _w28541_ ;
	assign \g241245/u3_syn_4  = _w28542_ ;
	assign \g241253/u3_syn_4  = _w28543_ ;
	assign \g241261/u3_syn_4  = _w28544_ ;
	assign \g241269/u3_syn_4  = _w28545_ ;
	assign \g241277/u3_syn_4  = _w28546_ ;
	assign \g241285/u3_syn_4  = _w28547_ ;
	assign \g241293/u3_syn_4  = _w28548_ ;
	assign \g241301/u3_syn_4  = _w28549_ ;
	assign \g241309/u3_syn_4  = _w28550_ ;
	assign \g241317/u3_syn_4  = _w28551_ ;
	assign \g241325/u3_syn_4  = _w28552_ ;
	assign \g241333/u3_syn_4  = _w28553_ ;
	assign \g241341/u3_syn_4  = _w28554_ ;
	assign \g241349/u3_syn_4  = _w28555_ ;
	assign \g241358/u3_syn_4  = _w28556_ ;
	assign \g241366/u3_syn_4  = _w28557_ ;
	assign \g241374/u3_syn_4  = _w28558_ ;
	assign \g241382/u3_syn_4  = _w28559_ ;
	assign \g241390/u3_syn_4  = _w28560_ ;
	assign \g241398/u3_syn_4  = _w28561_ ;
	assign \g241406/u3_syn_4  = _w28562_ ;
	assign \g241415/u3_syn_4  = _w28563_ ;
	assign \g241424/u3_syn_4  = _w28564_ ;
	assign \g241433/u3_syn_4  = _w28565_ ;
	assign \g241441/u3_syn_4  = _w28566_ ;
	assign \g241449/u3_syn_4  = _w28567_ ;
	assign \g241459/u3_syn_4  = _w28568_ ;
	assign \g241470/u3_syn_4  = _w28569_ ;
	assign \g241480/u3_syn_4  = _w28570_ ;
	assign \g241489/u3_syn_4  = _w28571_ ;
	assign \g241497/u3_syn_4  = _w28572_ ;
	assign \g241505/u3_syn_4  = _w28573_ ;
	assign \g241513/u3_syn_4  = _w28574_ ;
	assign \g241545/_3_  = _w28575_ ;
	assign \g241580/_00_  = _w28579_ ;
	assign \g241737/_0_  = _w28581_ ;
	assign \g241752/_0_  = _w28583_ ;
	assign \g241755/_0_  = _w28584_ ;
	assign \g241767/_2__syn_2  = _w28586_ ;
	assign \g241781/_1__syn_2  = _w28587_ ;
	assign \g241782/_0_  = _w28588_ ;
	assign \g241803/_1__syn_2  = _w28589_ ;
	assign \g241805/_0_  = _w28590_ ;
	assign \g241812/_1__syn_2  = _w28591_ ;
	assign \g241814/_1__syn_2  = _w28592_ ;
	assign \g241816/_1__syn_2  = _w28593_ ;
	assign \g241819/_1__syn_2  = _w28594_ ;
	assign \g241822/_1__syn_2  = _w28595_ ;
	assign \g241823/_0_  = _w28596_ ;
	assign \g241833/_1__syn_2  = _w28597_ ;
	assign \g241843/_1__syn_2  = _w28599_ ;
	assign \g241844/_1__syn_2  = _w28600_ ;
	assign \g241848/_1__syn_2  = _w28602_ ;
	assign \g241855/_1__syn_2  = _w28603_ ;
	assign \g241868/_1__syn_2  = _w28604_ ;
	assign \g242013/_1__syn_2  = _w28605_ ;
	assign \g242015/_1__syn_2  = _w28607_ ;
	assign \g242017/_1__syn_2  = _w28608_ ;
	assign \g242021/_1__syn_2  = _w28609_ ;
	assign \g242039/_1__syn_2  = _w28610_ ;
	assign \g242081/_0_  = _w28614_ ;
	assign \g242086/_0_  = _w28615_ ;
	assign \g242101/_3_  = _w11278_ ;
	assign \g242116/_0_  = _w28618_ ;
	assign \g242135/_2_  = _w24853_ ;
	assign \g242147/_0_  = _w28623_ ;
	assign \g242158/_0_  = _w28625_ ;
	assign \g242196/_0_  = _w28629_ ;
	assign \g242202/_0_  = _w28642_ ;
	assign \g242203/_0_  = _w28655_ ;
	assign \g242204/_0_  = _w28668_ ;
	assign \g242212/_0_  = _w28670_ ;
	assign \g242226/_01_  = _w28681_ ;
	assign \g242281/_0_  = _w28682_ ;
	assign \g242407/_0_  = _w28684_ ;
	assign \g242410/_0_  = _w28685_ ;
	assign \g242426/_0_  = _w28691_ ;
	assign \g242438/_2_  = _w28692_ ;
	assign \g242466/_0_  = _w28693_ ;
	assign \g242530/_0_  = _w28698_ ;
	assign \g242532/_0_  = _w28701_ ;
	assign \g243397/_0_  = _w28706_ ;
	assign \g245925/_0_  = _w28710_ ;
	assign \g245932/_0_  = _w28714_ ;
	assign \g245933/_0_  = _w28717_ ;
	assign \g245986/_3_  = _w28724_ ;
	assign \g250157/_3_  = _w28725_ ;
	assign \g250202/_0_  = _w28729_ ;
	assign \g250246/_1_  = _w28730_ ;
	assign \g250248/_0_  = _w28733_ ;
	assign \g250250/_0_  = _w28734_ ;
	assign \g250305/_0_  = _w28736_ ;
	assign \g250323/_0_  = _w28738_ ;
	assign \g250373/_0_  = _w28741_ ;
	assign \g250377/_0_  = _w28742_ ;
	assign \g250412/_0_  = _w28746_ ;
	assign \g250413/_0_  = _w28748_ ;
	assign \g250418/_0_  = _w28751_ ;
	assign \g250419/_0_  = _w28754_ ;
	assign \g250421/_0_  = _w28755_ ;
	assign \g250433/_0_  = _w28758_ ;
	assign \g250448/_3_  = _w28761_ ;
	assign \g250567/_3_  = _w11178_ ;
	assign \g258965/_0_  = _w28763_ ;
	assign \g259006/_0_  = _w28766_ ;
	assign \g259471/_0_  = _w28769_ ;
	assign \g259473/_2_  = _w28770_ ;
	assign \g260557/_0_  = _w28771_ ;
	assign \g261035/_0_  = _w28772_ ;
	assign \g261095/_3_  = _w28775_ ;
	assign \g261207/_2__syn_2  = _w28777_ ;
	assign \g261754/_0_  = _w28778_ ;
	assign \g262017/_0_  = _w28782_ ;
	assign \g262045/_0_  = _w28784_ ;
	assign \g262046/_0_  = _w28786_ ;
	assign \g262100/_3_  = _w28789_ ;
	assign \g263539/_1_  = _w13456_ ;
	assign \g263574/_0_  = _w12302_ ;
	assign \g263858/_0_  = _w10848_ ;
	assign \g264104/_1_  = _w28721_ ;
	assign \g264107/_1_  = _w27250_ ;
	assign \g264117/_0_  = _w28791_ ;
	assign \g264282/_0_  = _w28700_ ;
	assign \g264511/_0_  = _w28792_ ;
	assign \g264541/_0_  = _w28795_ ;
	assign \g264562/_0_  = _w28796_ ;
	assign \g264618/_0_  = _w28797_ ;
	assign \g264660/_0_  = _w28798_ ;
	assign \g264681/_3_  = _w28799_ ;
	assign \g264727/_0_  = _w28800_ ;
	assign \g265013/_0_  = _w28801_ ;
	assign \g265084/_0_  = _w28802_ ;
	assign \g265378/_0_  = _w28804_ ;
	assign \g265413/_0_  = _w28805_ ;
	assign \g265446/_0_  = _w28806_ ;
	assign \g265486/_0_  = _w28807_ ;
	assign \g265524/_3_  = _w10589_ ;
	assign \g265528/_3_  = _w10944_ ;
	assign \g265548/_3_  = _w10579_ ;
	assign \g265579/_0_  = _w11174_ ;
	assign \g265768/_0_  = _w28740_ ;
	assign \g265801/_0_  = _w11656_ ;
	assign \g265819/_1_  = _w25874_ ;
	assign \g265853/_0_  = _w28803_ ;
	assign \g265933/_0_  = _w28808_ ;
	assign \g266022/_0_  = _w28809_ ;
	assign \g266183/_1_  = _w26376_ ;
	assign \g281909/_0_  = _w28822_ ;
	assign \g281965/_1_  = _w28823_ ;
	assign \g282284/_1_  = _w28824_ ;
	assign \g282639/_1_  = _w28825_ ;
	assign \g283047/_0_  = _w28829_ ;
	assign \g283157/_1_  = _w28830_ ;
	assign \g283184/_0_  = _w28850_ ;
	assign \g283334/_3_  = _w28854_ ;
	assign int_o_pad = _w28859_ ;
	assign \m_wb_adr_o[0]_pad  = 1'b0;
	assign \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131_syn_2  = _w460_ ;
	assign \wishbone_tx_fifo_fifo_reg[2][15]/P0001_reg_syn_3  = _w28860_ ;
	assign \wishbone_tx_fifo_fifo_reg[2][16]/P0001_reg_syn_3  = _w28861_ ;
	assign \wishbone_tx_fifo_fifo_reg[2][17]/P0001_reg_syn_3  = _w28862_ ;
	assign \wishbone_tx_fifo_fifo_reg[2][22]/P0001_reg_syn_3  = _w28863_ ;
	assign \wishbone_tx_fifo_fifo_reg[2][23]/P0001_reg_syn_3  = _w28864_ ;
	assign \wishbone_tx_fifo_fifo_reg[2][25]/P0001_reg_syn_3  = _w28865_ ;
	assign \wishbone_tx_fifo_fifo_reg[2][2]/P0001_reg_syn_3  = _w28866_ ;
endmodule;