module top( \ahb_mst0_hsizeo_reg[0]/NET0131  , \ahb_mst0_hsizeo_reg[1]/NET0131  , \ahb_mst0_hsizeo_reg[2]/NET0131  , \ahb_mst0_m0_m1_diff_tx_reg/NET0131  , \ahb_mst0_mx_cmd_st_reg[0]/NET0131  , \ahb_mst0_mx_cmd_st_reg[1]/NET0131  , \ahb_mst0_mx_dtp_reg/NET0131  , \ahb_mst1_mx_cmd_st_reg[0]/NET0131  , \ahb_mst1_mx_cmd_st_reg[1]/NET0131  , \ahb_mst1_mx_dtp_reg/NET0131  , \ahb_slv_br_st_reg[0]/NET0131  , \ahb_slv_br_st_reg[1]/NET0131  , \ahb_slv_br_st_reg[2]/NET0131  , \ahb_slv_slv_ad_d1o_reg[2]/NET0131  , \ahb_slv_slv_ad_d1o_reg[3]/NET0131  , \ahb_slv_slv_ad_d1o_reg[4]/NET0131  , \ahb_slv_slv_ad_d1o_reg[5]/NET0131  , \ahb_slv_slv_ad_d1o_reg[6]/NET0131  , \ahb_slv_slv_ad_d1o_reg[7]/NET0131  , \ahb_slv_slv_ad_d1o_reg[8]/NET0131  , \ahb_slv_slv_br_req_reg/NET0131  , \ahb_slv_slv_pt_d1o_reg[0]/NET0131  , \ahb_slv_slv_pt_d1o_reg[1]/NET0131  , \ahb_slv_slv_pt_d1o_reg[2]/NET0131  , \ahb_slv_slv_pt_d1o_reg[3]/NET0131  , \ahb_slv_slv_sz_d1o_reg[0]/NET0131  , \ahb_slv_slv_sz_d1o_reg[1]/NET0131  , \ahb_slv_slv_sz_d1o_reg[2]/NET0131  , \ahb_slv_slv_wr_d1o_reg/NET0131  , \ch_sel_arb_ch_sel_reg[0]/P0000_reg_syn_2  , \ch_sel_arb_ch_sel_reg[1]/P0000_reg_syn_2  , \ch_sel_arb_ch_sel_reg[2]/P0000_reg_syn_2  , \ch_sel_arb_chcsr_reg_reg[10]/NET0131  , \ch_sel_arb_chcsr_reg_reg[11]/NET0131  , \ch_sel_arb_chcsr_reg_reg[12]/NET0131  , \ch_sel_arb_chcsr_reg_reg[13]/NET0131  , \ch_sel_arb_chcsr_reg_reg[15]/NET0131  , \ch_sel_arb_chcsr_reg_reg[16]/NET0131  , \ch_sel_arb_chcsr_reg_reg[17]/NET0131  , \ch_sel_arb_chcsr_reg_reg[18]/NET0131  , \ch_sel_arb_chcsr_reg_reg[19]/NET0131  , \ch_sel_arb_chcsr_reg_reg[1]/NET0131  , \ch_sel_arb_chcsr_reg_reg[20]/NET0131  , \ch_sel_arb_chcsr_reg_reg[2]/NET0131  , \ch_sel_arb_chcsr_reg_reg[3]/NET0131  , \ch_sel_arb_chcsr_reg_reg[4]/NET0131  , \ch_sel_arb_chcsr_reg_reg[5]/NET0131  , \ch_sel_arb_chcsr_reg_reg[6]/NET0131  , \ch_sel_arb_chcsr_reg_reg[8]/NET0131  , \ch_sel_arb_chcsr_reg_reg[9]/NET0131  , \ch_sel_arb_req_reg/NET0131  , \ch_sel_de_stup_d1_reg/NET0131  , \ch_sel_dma_reqd1_reg[0]/NET0131  , \ch_sel_dma_reqd1_reg[1]/NET0131  , \ch_sel_dma_reqd1_reg[2]/NET0131  , \ch_sel_dma_reqd1_reg[3]/NET0131  , \ch_sel_dma_reqd1_reg[4]/NET0131  , \ch_sel_dma_reqd1_reg[5]/NET0131  , \ch_sel_dma_reqd1_reg[6]/NET0131  , \ch_sel_dma_reqd1_reg[7]/NET0131  , \ch_sel_dma_reqd2_reg[0]/NET0131  , \ch_sel_dma_reqd2_reg[1]/P0001  , \ch_sel_dma_reqd2_reg[2]/P0001  , \ch_sel_dma_reqd2_reg[3]/P0001  , \ch_sel_dma_reqd2_reg[4]/NET0131  , \ch_sel_dma_reqd2_reg[5]/NET0131  , \ch_sel_dma_reqd2_reg[6]/NET0131  , \ch_sel_dma_reqd2_reg[7]/NET0131  , \ch_sel_dma_rrarb0_state_reg[0]/NET0131  , \ch_sel_dma_rrarb0_state_reg[1]/NET0131  , \ch_sel_dma_rrarb0_state_reg[2]/NET0131  , \ch_sel_dma_rrarb1_state_reg[0]/NET0131  , \ch_sel_dma_rrarb1_state_reg[1]/NET0131  , \ch_sel_dma_rrarb1_state_reg[2]/NET0131  , \ch_sel_dma_rrarb2_state_reg[0]/NET0131  , \ch_sel_dma_rrarb2_state_reg[1]/NET0131  , \ch_sel_dma_rrarb2_state_reg[2]/NET0131  , \ch_sel_dma_rrarb3_state_reg[0]/NET0131  , \ch_sel_dma_rrarb3_state_reg[1]/NET0131  , \ch_sel_dma_rrarb3_state_reg[2]/NET0131  , \ch_sel_fix_pri_sel_reg[0]/NET0131  , \ch_sel_fix_pri_sel_reg[1]/NET0131  , \ch_sel_vld_req_any_d1_reg/NET0131  , \ctl_rf_abt_reg[0]/NET0131  , \ctl_rf_abt_reg[1]/NET0131  , \ctl_rf_abt_reg[2]/NET0131  , \ctl_rf_abt_reg[3]/NET0131  , \ctl_rf_abt_reg[4]/NET0131  , \ctl_rf_abt_reg[5]/NET0131  , \ctl_rf_abt_reg[6]/NET0131  , \ctl_rf_abt_reg[7]/NET0131  , \ctl_rf_be_d1_reg[0]/P0001  , \ctl_rf_be_d1_reg[1]/P0001  , \ctl_rf_be_d1_reg[2]/P0001  , \ctl_rf_be_d1_reg[3]/P0001  , \ctl_rf_c0_rf_autold_reg/NET0131  , \ctl_rf_c0_rf_ch_en_reg/NET0131  , \ctl_rf_c0_rf_chabt_reg/NET0131  , \ctl_rf_c0_rf_chdad_reg[0]/NET0131  , \ctl_rf_c0_rf_chdad_reg[10]/P0002  , \ctl_rf_c0_rf_chdad_reg[11]/NET0131  , \ctl_rf_c0_rf_chdad_reg[12]/NET0131  , \ctl_rf_c0_rf_chdad_reg[13]/P0002  , \ctl_rf_c0_rf_chdad_reg[14]/NET0131  , \ctl_rf_c0_rf_chdad_reg[15]/NET0131  , \ctl_rf_c0_rf_chdad_reg[16]/NET0131  , \ctl_rf_c0_rf_chdad_reg[17]/NET0131  , \ctl_rf_c0_rf_chdad_reg[18]/NET0131  , \ctl_rf_c0_rf_chdad_reg[19]/NET0131  , \ctl_rf_c0_rf_chdad_reg[1]/NET0131  , \ctl_rf_c0_rf_chdad_reg[20]/P0002  , \ctl_rf_c0_rf_chdad_reg[21]/P0002  , \ctl_rf_c0_rf_chdad_reg[22]/P0002  , \ctl_rf_c0_rf_chdad_reg[23]/P0002  , \ctl_rf_c0_rf_chdad_reg[24]/P0002  , \ctl_rf_c0_rf_chdad_reg[25]/P0002  , \ctl_rf_c0_rf_chdad_reg[26]/P0002  , \ctl_rf_c0_rf_chdad_reg[27]/P0002  , \ctl_rf_c0_rf_chdad_reg[28]/P0002  , \ctl_rf_c0_rf_chdad_reg[29]/P0002  , \ctl_rf_c0_rf_chdad_reg[2]/NET0131  , \ctl_rf_c0_rf_chdad_reg[30]/P0002  , \ctl_rf_c0_rf_chdad_reg[31]/P0002  , \ctl_rf_c0_rf_chdad_reg[3]/P0002  , \ctl_rf_c0_rf_chdad_reg[4]/P0002  , \ctl_rf_c0_rf_chdad_reg[5]/P0002  , \ctl_rf_c0_rf_chdad_reg[6]/P0002  , \ctl_rf_c0_rf_chdad_reg[7]/P0002  , \ctl_rf_c0_rf_chdad_reg[8]/NET0131  , \ctl_rf_c0_rf_chdad_reg[9]/P0002  , \ctl_rf_c0_rf_chllp_cnt_reg[0]/NET0131  , \ctl_rf_c0_rf_chllp_cnt_reg[1]/NET0131  , \ctl_rf_c0_rf_chllp_cnt_reg[2]/NET0131  , \ctl_rf_c0_rf_chllp_cnt_reg[3]/NET0131  , \ctl_rf_c0_rf_chllp_on_reg/NET0131  , \ctl_rf_c0_rf_chllp_reg[0]/P0002  , \ctl_rf_c0_rf_chllp_reg[10]/NET0131  , \ctl_rf_c0_rf_chllp_reg[11]/NET0131  , \ctl_rf_c0_rf_chllp_reg[12]/NET0131  , \ctl_rf_c0_rf_chllp_reg[13]/NET0131  , \ctl_rf_c0_rf_chllp_reg[14]/NET0131  , \ctl_rf_c0_rf_chllp_reg[15]/NET0131  , \ctl_rf_c0_rf_chllp_reg[16]/NET0131  , \ctl_rf_c0_rf_chllp_reg[17]/NET0131  , \ctl_rf_c0_rf_chllp_reg[18]/NET0131  , \ctl_rf_c0_rf_chllp_reg[19]/NET0131  , \ctl_rf_c0_rf_chllp_reg[1]/P0002  , \ctl_rf_c0_rf_chllp_reg[20]/NET0131  , \ctl_rf_c0_rf_chllp_reg[21]/NET0131  , \ctl_rf_c0_rf_chllp_reg[22]/NET0131  , \ctl_rf_c0_rf_chllp_reg[23]/NET0131  , \ctl_rf_c0_rf_chllp_reg[24]/NET0131  , \ctl_rf_c0_rf_chllp_reg[25]/NET0131  , \ctl_rf_c0_rf_chllp_reg[26]/NET0131  , \ctl_rf_c0_rf_chllp_reg[27]/NET0131  , \ctl_rf_c0_rf_chllp_reg[28]/NET0131  , \ctl_rf_c0_rf_chllp_reg[29]/NET0131  , \ctl_rf_c0_rf_chllp_reg[2]/NET0131  , \ctl_rf_c0_rf_chllp_reg[30]/NET0131  , \ctl_rf_c0_rf_chllp_reg[31]/NET0131  , \ctl_rf_c0_rf_chllp_reg[3]/NET0131  , \ctl_rf_c0_rf_chllp_reg[4]/NET0131  , \ctl_rf_c0_rf_chllp_reg[5]/NET0131  , \ctl_rf_c0_rf_chllp_reg[6]/NET0131  , \ctl_rf_c0_rf_chllp_reg[7]/NET0131  , \ctl_rf_c0_rf_chllp_reg[8]/NET0131  , \ctl_rf_c0_rf_chllp_reg[9]/NET0131  , \ctl_rf_c0_rf_chllpen_reg/NET0131  , \ctl_rf_c0_rf_chpri_reg[0]/NET0131  , \ctl_rf_c0_rf_chpri_reg[1]/NET0131  , \ctl_rf_c0_rf_chsad_reg[0]/NET0131  , \ctl_rf_c0_rf_chsad_reg[10]/NET0131  , \ctl_rf_c0_rf_chsad_reg[11]/P0002  , \ctl_rf_c0_rf_chsad_reg[12]/P0002  , \ctl_rf_c0_rf_chsad_reg[13]/NET0131  , \ctl_rf_c0_rf_chsad_reg[14]/P0002  , \ctl_rf_c0_rf_chsad_reg[15]/P0002  , \ctl_rf_c0_rf_chsad_reg[16]/NET0131  , \ctl_rf_c0_rf_chsad_reg[17]/NET0131  , \ctl_rf_c0_rf_chsad_reg[18]/NET0131  , \ctl_rf_c0_rf_chsad_reg[19]/NET0131  , \ctl_rf_c0_rf_chsad_reg[1]/NET0131  , \ctl_rf_c0_rf_chsad_reg[20]/NET0131  , \ctl_rf_c0_rf_chsad_reg[21]/NET0131  , \ctl_rf_c0_rf_chsad_reg[22]/NET0131  , \ctl_rf_c0_rf_chsad_reg[23]/NET0131  , \ctl_rf_c0_rf_chsad_reg[24]/NET0131  , \ctl_rf_c0_rf_chsad_reg[25]/P0002  , \ctl_rf_c0_rf_chsad_reg[26]/P0002  , \ctl_rf_c0_rf_chsad_reg[27]/P0002  , \ctl_rf_c0_rf_chsad_reg[28]/P0002  , \ctl_rf_c0_rf_chsad_reg[29]/P0002  , \ctl_rf_c0_rf_chsad_reg[2]/NET0131  , \ctl_rf_c0_rf_chsad_reg[30]/P0002  , \ctl_rf_c0_rf_chsad_reg[31]/NET0131  , \ctl_rf_c0_rf_chsad_reg[3]/NET0131  , \ctl_rf_c0_rf_chsad_reg[4]/NET0131  , \ctl_rf_c0_rf_chsad_reg[5]/NET0131  , \ctl_rf_c0_rf_chsad_reg[6]/NET0131  , \ctl_rf_c0_rf_chsad_reg[7]/NET0131  , \ctl_rf_c0_rf_chsad_reg[8]/P0002  , \ctl_rf_c0_rf_chsad_reg[9]/NET0131  , \ctl_rf_c0_rf_chtsz_reg[0]/P0002  , \ctl_rf_c0_rf_chtsz_reg[10]/P0002  , \ctl_rf_c0_rf_chtsz_reg[11]/P0002  , \ctl_rf_c0_rf_chtsz_reg[1]/P0002  , \ctl_rf_c0_rf_chtsz_reg[2]/P0002  , \ctl_rf_c0_rf_chtsz_reg[3]/P0002  , \ctl_rf_c0_rf_chtsz_reg[4]/NET0131  , \ctl_rf_c0_rf_chtsz_reg[5]/NET0131  , \ctl_rf_c0_rf_chtsz_reg[6]/NET0131  , \ctl_rf_c0_rf_chtsz_reg[7]/NET0131  , \ctl_rf_c0_rf_chtsz_reg[8]/P0002  , \ctl_rf_c0_rf_chtsz_reg[9]/P0002  , \ctl_rf_c0_rf_dad_ctl0_reg/NET0131  , \ctl_rf_c0_rf_dad_ctl1_reg/NET0131  , \ctl_rf_c0_rf_dreqmode_reg/NET0131  , \ctl_rf_c0_rf_dst_sel_reg/NET0131  , \ctl_rf_c0_rf_dwidth_reg[0]/NET0131  , \ctl_rf_c0_rf_dwidth_reg[1]/NET0131  , \ctl_rf_c0_rf_dwidth_reg[2]/NET0131  , \ctl_rf_c0_rf_int_abt_msk_reg/NET0131  , \ctl_rf_c0_rf_int_err_msk_reg/NET0131  , \ctl_rf_c0_rf_int_tc1_msk_reg/NET0131  , \ctl_rf_c0_rf_int_tc_msk_reg/NET0131  , \ctl_rf_c0_rf_mode_reg/NET0131  , \ctl_rf_c0_rf_prot1_reg/NET0131  , \ctl_rf_c0_rf_prot2_reg/NET0131  , \ctl_rf_c0_rf_prot3_reg/NET0131  , \ctl_rf_c0_rf_sad_ctl0_reg/NET0131  , \ctl_rf_c0_rf_sad_ctl1_reg/NET0131  , \ctl_rf_c0_rf_src_sel_reg/NET0131  , \ctl_rf_c0_rf_src_sz_reg[0]/NET0131  , \ctl_rf_c0_rf_src_sz_reg[1]/NET0131  , \ctl_rf_c0_rf_src_sz_reg[2]/NET0131  , \ctl_rf_c0_rf_swidth_reg[0]/NET0131  , \ctl_rf_c0_rf_swidth_reg[1]/NET0131  , \ctl_rf_c0_rf_swidth_reg[2]/NET0131  , \ctl_rf_c0brbs_reg[16]/NET0131  , \ctl_rf_c0brbs_reg[17]/NET0131  , \ctl_rf_c0brbs_reg[18]/NET0131  , \ctl_rf_c0brbs_reg[19]/NET0131  , \ctl_rf_c0brbs_reg[20]/NET0131  , \ctl_rf_c0brbs_reg[21]/NET0131  , \ctl_rf_c0brbs_reg[22]/NET0131  , \ctl_rf_c0brbs_reg[23]/NET0131  , \ctl_rf_c0brbs_reg[24]/NET0131  , \ctl_rf_c0brbs_reg[25]/NET0131  , \ctl_rf_c0brbs_reg[26]/NET0131  , \ctl_rf_c0brbs_reg[27]/NET0131  , \ctl_rf_c0brbs_reg[28]/NET0131  , \ctl_rf_c0brbs_reg[29]/NET0131  , \ctl_rf_c0brbs_reg[30]/NET0131  , \ctl_rf_c0brbs_reg[31]/NET0131  , \ctl_rf_c0dmabs_reg[16]/NET0131  , \ctl_rf_c0dmabs_reg[17]/NET0131  , \ctl_rf_c0dmabs_reg[18]/NET0131  , \ctl_rf_c0dmabs_reg[19]/NET0131  , \ctl_rf_c0dmabs_reg[20]/NET0131  , \ctl_rf_c0dmabs_reg[21]/NET0131  , \ctl_rf_c0dmabs_reg[22]/NET0131  , \ctl_rf_c0dmabs_reg[23]/NET0131  , \ctl_rf_c0dmabs_reg[24]/NET0131  , \ctl_rf_c0dmabs_reg[25]/NET0131  , \ctl_rf_c0dmabs_reg[26]/NET0131  , \ctl_rf_c0dmabs_reg[27]/NET0131  , \ctl_rf_c0dmabs_reg[28]/NET0131  , \ctl_rf_c0dmabs_reg[29]/NET0131  , \ctl_rf_c0dmabs_reg[30]/NET0131  , \ctl_rf_c0dmabs_reg[31]/NET0131  , \ctl_rf_c1_rf_autold_reg/NET0131  , \ctl_rf_c1_rf_ch_en_reg/NET0131  , \ctl_rf_c1_rf_chabt_reg/NET0131  , \ctl_rf_c1_rf_chdad_reg[0]/NET0131  , \ctl_rf_c1_rf_chdad_reg[10]/NET0131  , \ctl_rf_c1_rf_chdad_reg[11]/P0002  , \ctl_rf_c1_rf_chdad_reg[12]/NET0131  , \ctl_rf_c1_rf_chdad_reg[13]/NET0131  , \ctl_rf_c1_rf_chdad_reg[14]/NET0131  , \ctl_rf_c1_rf_chdad_reg[15]/NET0131  , \ctl_rf_c1_rf_chdad_reg[16]/NET0131  , \ctl_rf_c1_rf_chdad_reg[17]/NET0131  , \ctl_rf_c1_rf_chdad_reg[18]/NET0131  , \ctl_rf_c1_rf_chdad_reg[19]/NET0131  , \ctl_rf_c1_rf_chdad_reg[1]/NET0131  , \ctl_rf_c1_rf_chdad_reg[20]/P0002  , \ctl_rf_c1_rf_chdad_reg[21]/P0002  , \ctl_rf_c1_rf_chdad_reg[22]/P0002  , \ctl_rf_c1_rf_chdad_reg[23]/P0002  , \ctl_rf_c1_rf_chdad_reg[24]/P0002  , \ctl_rf_c1_rf_chdad_reg[25]/P0002  , \ctl_rf_c1_rf_chdad_reg[26]/P0002  , \ctl_rf_c1_rf_chdad_reg[27]/P0002  , \ctl_rf_c1_rf_chdad_reg[28]/P0002  , \ctl_rf_c1_rf_chdad_reg[29]/P0002  , \ctl_rf_c1_rf_chdad_reg[2]/NET0131  , \ctl_rf_c1_rf_chdad_reg[30]/P0002  , \ctl_rf_c1_rf_chdad_reg[31]/P0002  , \ctl_rf_c1_rf_chdad_reg[3]/P0002  , \ctl_rf_c1_rf_chdad_reg[4]/P0002  , \ctl_rf_c1_rf_chdad_reg[5]/P0002  , \ctl_rf_c1_rf_chdad_reg[6]/P0002  , \ctl_rf_c1_rf_chdad_reg[7]/P0002  , \ctl_rf_c1_rf_chdad_reg[8]/NET0131  , \ctl_rf_c1_rf_chdad_reg[9]/P0002  , \ctl_rf_c1_rf_chllp_cnt_reg[0]/NET0131  , \ctl_rf_c1_rf_chllp_cnt_reg[1]/NET0131  , \ctl_rf_c1_rf_chllp_cnt_reg[2]/NET0131  , \ctl_rf_c1_rf_chllp_cnt_reg[3]/NET0131  , \ctl_rf_c1_rf_chllp_on_reg/NET0131  , \ctl_rf_c1_rf_chllp_reg[0]/P0002  , \ctl_rf_c1_rf_chllp_reg[10]/NET0131  , \ctl_rf_c1_rf_chllp_reg[11]/NET0131  , \ctl_rf_c1_rf_chllp_reg[12]/NET0131  , \ctl_rf_c1_rf_chllp_reg[13]/NET0131  , \ctl_rf_c1_rf_chllp_reg[14]/NET0131  , \ctl_rf_c1_rf_chllp_reg[15]/NET0131  , \ctl_rf_c1_rf_chllp_reg[16]/NET0131  , \ctl_rf_c1_rf_chllp_reg[17]/NET0131  , \ctl_rf_c1_rf_chllp_reg[18]/NET0131  , \ctl_rf_c1_rf_chllp_reg[19]/NET0131  , \ctl_rf_c1_rf_chllp_reg[1]/P0002  , \ctl_rf_c1_rf_chllp_reg[20]/NET0131  , \ctl_rf_c1_rf_chllp_reg[21]/NET0131  , \ctl_rf_c1_rf_chllp_reg[22]/NET0131  , \ctl_rf_c1_rf_chllp_reg[23]/NET0131  , \ctl_rf_c1_rf_chllp_reg[24]/NET0131  , \ctl_rf_c1_rf_chllp_reg[25]/NET0131  , \ctl_rf_c1_rf_chllp_reg[26]/NET0131  , \ctl_rf_c1_rf_chllp_reg[27]/NET0131  , \ctl_rf_c1_rf_chllp_reg[28]/NET0131  , \ctl_rf_c1_rf_chllp_reg[29]/NET0131  , \ctl_rf_c1_rf_chllp_reg[2]/NET0131  , \ctl_rf_c1_rf_chllp_reg[30]/NET0131  , \ctl_rf_c1_rf_chllp_reg[31]/NET0131  , \ctl_rf_c1_rf_chllp_reg[3]/NET0131  , \ctl_rf_c1_rf_chllp_reg[4]/NET0131  , \ctl_rf_c1_rf_chllp_reg[5]/NET0131  , \ctl_rf_c1_rf_chllp_reg[6]/NET0131  , \ctl_rf_c1_rf_chllp_reg[7]/NET0131  , \ctl_rf_c1_rf_chllp_reg[8]/NET0131  , \ctl_rf_c1_rf_chllp_reg[9]/NET0131  , \ctl_rf_c1_rf_chllpen_reg/NET0131  , \ctl_rf_c1_rf_chpri_reg[0]/NET0131  , \ctl_rf_c1_rf_chpri_reg[1]/NET0131  , \ctl_rf_c1_rf_chsad_reg[0]/NET0131  , \ctl_rf_c1_rf_chsad_reg[10]/P0002  , \ctl_rf_c1_rf_chsad_reg[11]/NET0131  , \ctl_rf_c1_rf_chsad_reg[12]/P0002  , \ctl_rf_c1_rf_chsad_reg[13]/P0002  , \ctl_rf_c1_rf_chsad_reg[14]/P0002  , \ctl_rf_c1_rf_chsad_reg[15]/P0002  , \ctl_rf_c1_rf_chsad_reg[16]/NET0131  , \ctl_rf_c1_rf_chsad_reg[17]/NET0131  , \ctl_rf_c1_rf_chsad_reg[18]/NET0131  , \ctl_rf_c1_rf_chsad_reg[19]/NET0131  , \ctl_rf_c1_rf_chsad_reg[1]/NET0131  , \ctl_rf_c1_rf_chsad_reg[20]/NET0131  , \ctl_rf_c1_rf_chsad_reg[21]/NET0131  , \ctl_rf_c1_rf_chsad_reg[22]/NET0131  , \ctl_rf_c1_rf_chsad_reg[23]/NET0131  , \ctl_rf_c1_rf_chsad_reg[24]/NET0131  , \ctl_rf_c1_rf_chsad_reg[25]/P0002  , \ctl_rf_c1_rf_chsad_reg[26]/P0002  , \ctl_rf_c1_rf_chsad_reg[27]/P0002  , \ctl_rf_c1_rf_chsad_reg[28]/P0002  , \ctl_rf_c1_rf_chsad_reg[29]/P0002  , \ctl_rf_c1_rf_chsad_reg[2]/NET0131  , \ctl_rf_c1_rf_chsad_reg[30]/P0002  , \ctl_rf_c1_rf_chsad_reg[31]/NET0131  , \ctl_rf_c1_rf_chsad_reg[3]/NET0131  , \ctl_rf_c1_rf_chsad_reg[4]/NET0131  , \ctl_rf_c1_rf_chsad_reg[5]/NET0131  , \ctl_rf_c1_rf_chsad_reg[6]/NET0131  , \ctl_rf_c1_rf_chsad_reg[7]/NET0131  , \ctl_rf_c1_rf_chsad_reg[8]/P0002  , \ctl_rf_c1_rf_chsad_reg[9]/NET0131  , \ctl_rf_c1_rf_chtsz_reg[0]/P0002  , \ctl_rf_c1_rf_chtsz_reg[10]/P0002  , \ctl_rf_c1_rf_chtsz_reg[11]/P0002  , \ctl_rf_c1_rf_chtsz_reg[1]/P0002  , \ctl_rf_c1_rf_chtsz_reg[2]/P0002  , \ctl_rf_c1_rf_chtsz_reg[3]/P0002  , \ctl_rf_c1_rf_chtsz_reg[4]/NET0131  , \ctl_rf_c1_rf_chtsz_reg[5]/NET0131  , \ctl_rf_c1_rf_chtsz_reg[6]/NET0131  , \ctl_rf_c1_rf_chtsz_reg[7]/NET0131  , \ctl_rf_c1_rf_chtsz_reg[8]/P0002  , \ctl_rf_c1_rf_chtsz_reg[9]/P0002  , \ctl_rf_c1_rf_dad_ctl0_reg/NET0131  , \ctl_rf_c1_rf_dad_ctl1_reg/NET0131  , \ctl_rf_c1_rf_dreqmode_reg/NET0131  , \ctl_rf_c1_rf_dst_sel_reg/NET0131  , \ctl_rf_c1_rf_dwidth_reg[0]/NET0131  , \ctl_rf_c1_rf_dwidth_reg[1]/NET0131  , \ctl_rf_c1_rf_dwidth_reg[2]/NET0131  , \ctl_rf_c1_rf_int_abt_msk_reg/NET0131  , \ctl_rf_c1_rf_int_err_msk_reg/NET0131  , \ctl_rf_c1_rf_int_tc1_msk_reg/NET0131  , \ctl_rf_c1_rf_int_tc_msk_reg/NET0131  , \ctl_rf_c1_rf_mode_reg/NET0131  , \ctl_rf_c1_rf_prot1_reg/NET0131  , \ctl_rf_c1_rf_prot2_reg/NET0131  , \ctl_rf_c1_rf_prot3_reg/NET0131  , \ctl_rf_c1_rf_sad_ctl0_reg/NET0131  , \ctl_rf_c1_rf_sad_ctl1_reg/NET0131  , \ctl_rf_c1_rf_src_sel_reg/NET0131  , \ctl_rf_c1_rf_src_sz_reg[0]/NET0131  , \ctl_rf_c1_rf_src_sz_reg[1]/NET0131  , \ctl_rf_c1_rf_src_sz_reg[2]/NET0131  , \ctl_rf_c1_rf_swidth_reg[0]/NET0131  , \ctl_rf_c1_rf_swidth_reg[1]/NET0131  , \ctl_rf_c1_rf_swidth_reg[2]/NET0131  , \ctl_rf_c1brbs_reg[16]/NET0131  , \ctl_rf_c1brbs_reg[17]/NET0131  , \ctl_rf_c1brbs_reg[18]/NET0131  , \ctl_rf_c1brbs_reg[19]/NET0131  , \ctl_rf_c1brbs_reg[20]/NET0131  , \ctl_rf_c1brbs_reg[21]/NET0131  , \ctl_rf_c1brbs_reg[22]/NET0131  , \ctl_rf_c1brbs_reg[23]/NET0131  , \ctl_rf_c1brbs_reg[24]/NET0131  , \ctl_rf_c1brbs_reg[25]/NET0131  , \ctl_rf_c1brbs_reg[26]/NET0131  , \ctl_rf_c1brbs_reg[27]/NET0131  , \ctl_rf_c1brbs_reg[28]/NET0131  , \ctl_rf_c1brbs_reg[29]/NET0131  , \ctl_rf_c1brbs_reg[30]/NET0131  , \ctl_rf_c1brbs_reg[31]/NET0131  , \ctl_rf_c1dmabs_reg[16]/NET0131  , \ctl_rf_c1dmabs_reg[17]/NET0131  , \ctl_rf_c1dmabs_reg[18]/NET0131  , \ctl_rf_c1dmabs_reg[19]/NET0131  , \ctl_rf_c1dmabs_reg[20]/NET0131  , \ctl_rf_c1dmabs_reg[21]/NET0131  , \ctl_rf_c1dmabs_reg[22]/NET0131  , \ctl_rf_c1dmabs_reg[23]/NET0131  , \ctl_rf_c1dmabs_reg[24]/NET0131  , \ctl_rf_c1dmabs_reg[25]/NET0131  , \ctl_rf_c1dmabs_reg[26]/NET0131  , \ctl_rf_c1dmabs_reg[27]/NET0131  , \ctl_rf_c1dmabs_reg[28]/NET0131  , \ctl_rf_c1dmabs_reg[29]/NET0131  , \ctl_rf_c1dmabs_reg[30]/NET0131  , \ctl_rf_c1dmabs_reg[31]/NET0131  , \ctl_rf_c2_rf_autold_reg/NET0131  , \ctl_rf_c2_rf_ch_en_reg/NET0131  , \ctl_rf_c2_rf_chabt_reg/NET0131  , \ctl_rf_c2_rf_chdad_reg[0]/NET0131  , \ctl_rf_c2_rf_chdad_reg[10]/P0002  , \ctl_rf_c2_rf_chdad_reg[11]/P0002  , \ctl_rf_c2_rf_chdad_reg[12]/P0002  , \ctl_rf_c2_rf_chdad_reg[13]/P0002  , \ctl_rf_c2_rf_chdad_reg[14]/P0002  , \ctl_rf_c2_rf_chdad_reg[15]/P0002  , \ctl_rf_c2_rf_chdad_reg[16]/NET0131  , \ctl_rf_c2_rf_chdad_reg[17]/NET0131  , \ctl_rf_c2_rf_chdad_reg[18]/NET0131  , \ctl_rf_c2_rf_chdad_reg[19]/NET0131  , \ctl_rf_c2_rf_chdad_reg[1]/NET0131  , \ctl_rf_c2_rf_chdad_reg[20]/P0002  , \ctl_rf_c2_rf_chdad_reg[21]/P0002  , \ctl_rf_c2_rf_chdad_reg[22]/P0002  , \ctl_rf_c2_rf_chdad_reg[23]/P0002  , \ctl_rf_c2_rf_chdad_reg[24]/P0002  , \ctl_rf_c2_rf_chdad_reg[25]/P0002  , \ctl_rf_c2_rf_chdad_reg[26]/P0002  , \ctl_rf_c2_rf_chdad_reg[27]/P0002  , \ctl_rf_c2_rf_chdad_reg[28]/P0002  , \ctl_rf_c2_rf_chdad_reg[29]/P0002  , \ctl_rf_c2_rf_chdad_reg[2]/NET0131  , \ctl_rf_c2_rf_chdad_reg[30]/P0002  , \ctl_rf_c2_rf_chdad_reg[31]/P0002  , \ctl_rf_c2_rf_chdad_reg[3]/P0002  , \ctl_rf_c2_rf_chdad_reg[4]/P0002  , \ctl_rf_c2_rf_chdad_reg[5]/P0002  , \ctl_rf_c2_rf_chdad_reg[6]/P0002  , \ctl_rf_c2_rf_chdad_reg[7]/P0002  , \ctl_rf_c2_rf_chdad_reg[8]/NET0131  , \ctl_rf_c2_rf_chdad_reg[9]/P0002  , \ctl_rf_c2_rf_chllp_cnt_reg[0]/NET0131  , \ctl_rf_c2_rf_chllp_cnt_reg[1]/NET0131  , \ctl_rf_c2_rf_chllp_cnt_reg[2]/NET0131  , \ctl_rf_c2_rf_chllp_cnt_reg[3]/NET0131  , \ctl_rf_c2_rf_chllp_on_reg/NET0131  , \ctl_rf_c2_rf_chllp_reg[0]/P0002  , \ctl_rf_c2_rf_chllp_reg[10]/NET0131  , \ctl_rf_c2_rf_chllp_reg[11]/NET0131  , \ctl_rf_c2_rf_chllp_reg[12]/NET0131  , \ctl_rf_c2_rf_chllp_reg[13]/NET0131  , \ctl_rf_c2_rf_chllp_reg[14]/NET0131  , \ctl_rf_c2_rf_chllp_reg[15]/NET0131  , \ctl_rf_c2_rf_chllp_reg[16]/NET0131  , \ctl_rf_c2_rf_chllp_reg[17]/NET0131  , \ctl_rf_c2_rf_chllp_reg[18]/NET0131  , \ctl_rf_c2_rf_chllp_reg[19]/NET0131  , \ctl_rf_c2_rf_chllp_reg[1]/P0002  , \ctl_rf_c2_rf_chllp_reg[20]/NET0131  , \ctl_rf_c2_rf_chllp_reg[21]/NET0131  , \ctl_rf_c2_rf_chllp_reg[22]/NET0131  , \ctl_rf_c2_rf_chllp_reg[23]/NET0131  , \ctl_rf_c2_rf_chllp_reg[24]/NET0131  , \ctl_rf_c2_rf_chllp_reg[25]/NET0131  , \ctl_rf_c2_rf_chllp_reg[26]/NET0131  , \ctl_rf_c2_rf_chllp_reg[27]/NET0131  , \ctl_rf_c2_rf_chllp_reg[28]/NET0131  , \ctl_rf_c2_rf_chllp_reg[29]/NET0131  , \ctl_rf_c2_rf_chllp_reg[2]/NET0131  , \ctl_rf_c2_rf_chllp_reg[30]/NET0131  , \ctl_rf_c2_rf_chllp_reg[31]/NET0131  , \ctl_rf_c2_rf_chllp_reg[3]/NET0131  , \ctl_rf_c2_rf_chllp_reg[4]/NET0131  , \ctl_rf_c2_rf_chllp_reg[5]/NET0131  , \ctl_rf_c2_rf_chllp_reg[6]/NET0131  , \ctl_rf_c2_rf_chllp_reg[7]/NET0131  , \ctl_rf_c2_rf_chllp_reg[8]/NET0131  , \ctl_rf_c2_rf_chllp_reg[9]/NET0131  , \ctl_rf_c2_rf_chllpen_reg/NET0131  , \ctl_rf_c2_rf_chpri_reg[0]/NET0131  , \ctl_rf_c2_rf_chpri_reg[1]/NET0131  , \ctl_rf_c2_rf_chsad_reg[0]/NET0131  , \ctl_rf_c2_rf_chsad_reg[10]/NET0131  , \ctl_rf_c2_rf_chsad_reg[11]/NET0131  , \ctl_rf_c2_rf_chsad_reg[12]/NET0131  , \ctl_rf_c2_rf_chsad_reg[13]/NET0131  , \ctl_rf_c2_rf_chsad_reg[14]/NET0131  , \ctl_rf_c2_rf_chsad_reg[15]/NET0131  , \ctl_rf_c2_rf_chsad_reg[16]/NET0131  , \ctl_rf_c2_rf_chsad_reg[17]/NET0131  , \ctl_rf_c2_rf_chsad_reg[18]/NET0131  , \ctl_rf_c2_rf_chsad_reg[19]/NET0131  , \ctl_rf_c2_rf_chsad_reg[1]/NET0131  , \ctl_rf_c2_rf_chsad_reg[20]/NET0131  , \ctl_rf_c2_rf_chsad_reg[21]/NET0131  , \ctl_rf_c2_rf_chsad_reg[22]/NET0131  , \ctl_rf_c2_rf_chsad_reg[23]/NET0131  , \ctl_rf_c2_rf_chsad_reg[24]/NET0131  , \ctl_rf_c2_rf_chsad_reg[25]/P0002  , \ctl_rf_c2_rf_chsad_reg[26]/P0002  , \ctl_rf_c2_rf_chsad_reg[27]/P0002  , \ctl_rf_c2_rf_chsad_reg[28]/P0002  , \ctl_rf_c2_rf_chsad_reg[29]/P0002  , \ctl_rf_c2_rf_chsad_reg[2]/NET0131  , \ctl_rf_c2_rf_chsad_reg[30]/P0002  , \ctl_rf_c2_rf_chsad_reg[31]/NET0131  , \ctl_rf_c2_rf_chsad_reg[3]/NET0131  , \ctl_rf_c2_rf_chsad_reg[4]/NET0131  , \ctl_rf_c2_rf_chsad_reg[5]/NET0131  , \ctl_rf_c2_rf_chsad_reg[6]/NET0131  , \ctl_rf_c2_rf_chsad_reg[7]/NET0131  , \ctl_rf_c2_rf_chsad_reg[8]/P0002  , \ctl_rf_c2_rf_chsad_reg[9]/NET0131  , \ctl_rf_c2_rf_chtsz_reg[0]/P0002  , \ctl_rf_c2_rf_chtsz_reg[10]/P0002  , \ctl_rf_c2_rf_chtsz_reg[11]/P0002  , \ctl_rf_c2_rf_chtsz_reg[1]/P0002  , \ctl_rf_c2_rf_chtsz_reg[2]/P0002  , \ctl_rf_c2_rf_chtsz_reg[3]/P0002  , \ctl_rf_c2_rf_chtsz_reg[4]/NET0131  , \ctl_rf_c2_rf_chtsz_reg[5]/NET0131  , \ctl_rf_c2_rf_chtsz_reg[6]/NET0131  , \ctl_rf_c2_rf_chtsz_reg[7]/NET0131  , \ctl_rf_c2_rf_chtsz_reg[8]/P0002  , \ctl_rf_c2_rf_chtsz_reg[9]/P0002  , \ctl_rf_c2_rf_dad_ctl0_reg/NET0131  , \ctl_rf_c2_rf_dad_ctl1_reg/NET0131  , \ctl_rf_c2_rf_dreqmode_reg/NET0131  , \ctl_rf_c2_rf_dst_sel_reg/NET0131  , \ctl_rf_c2_rf_dwidth_reg[0]/NET0131  , \ctl_rf_c2_rf_dwidth_reg[1]/NET0131  , \ctl_rf_c2_rf_dwidth_reg[2]/NET0131  , \ctl_rf_c2_rf_int_abt_msk_reg/NET0131  , \ctl_rf_c2_rf_int_err_msk_reg/NET0131  , \ctl_rf_c2_rf_int_tc1_msk_reg/NET0131  , \ctl_rf_c2_rf_int_tc_msk_reg/NET0131  , \ctl_rf_c2_rf_mode_reg/NET0131  , \ctl_rf_c2_rf_prot1_reg/NET0131  , \ctl_rf_c2_rf_prot2_reg/NET0131  , \ctl_rf_c2_rf_prot3_reg/NET0131  , \ctl_rf_c2_rf_sad_ctl0_reg/NET0131  , \ctl_rf_c2_rf_sad_ctl1_reg/NET0131  , \ctl_rf_c2_rf_src_sel_reg/NET0131  , \ctl_rf_c2_rf_src_sz_reg[0]/NET0131  , \ctl_rf_c2_rf_src_sz_reg[1]/NET0131  , \ctl_rf_c2_rf_src_sz_reg[2]/NET0131  , \ctl_rf_c2_rf_swidth_reg[0]/NET0131  , \ctl_rf_c2_rf_swidth_reg[1]/NET0131  , \ctl_rf_c2_rf_swidth_reg[2]/NET0131  , \ctl_rf_c2brbs_reg[16]/NET0131  , \ctl_rf_c2brbs_reg[17]/NET0131  , \ctl_rf_c2brbs_reg[18]/NET0131  , \ctl_rf_c2brbs_reg[19]/NET0131  , \ctl_rf_c2brbs_reg[20]/NET0131  , \ctl_rf_c2brbs_reg[21]/NET0131  , \ctl_rf_c2brbs_reg[22]/NET0131  , \ctl_rf_c2brbs_reg[23]/NET0131  , \ctl_rf_c2brbs_reg[24]/NET0131  , \ctl_rf_c2brbs_reg[25]/NET0131  , \ctl_rf_c2brbs_reg[26]/NET0131  , \ctl_rf_c2brbs_reg[27]/NET0131  , \ctl_rf_c2brbs_reg[28]/NET0131  , \ctl_rf_c2brbs_reg[29]/NET0131  , \ctl_rf_c2brbs_reg[30]/NET0131  , \ctl_rf_c2brbs_reg[31]/NET0131  , \ctl_rf_c2dmabs_reg[16]/NET0131  , \ctl_rf_c2dmabs_reg[17]/NET0131  , \ctl_rf_c2dmabs_reg[18]/NET0131  , \ctl_rf_c2dmabs_reg[19]/NET0131  , \ctl_rf_c2dmabs_reg[20]/NET0131  , \ctl_rf_c2dmabs_reg[21]/NET0131  , \ctl_rf_c2dmabs_reg[22]/NET0131  , \ctl_rf_c2dmabs_reg[23]/NET0131  , \ctl_rf_c2dmabs_reg[24]/NET0131  , \ctl_rf_c2dmabs_reg[25]/NET0131  , \ctl_rf_c2dmabs_reg[26]/NET0131  , \ctl_rf_c2dmabs_reg[27]/NET0131  , \ctl_rf_c2dmabs_reg[28]/NET0131  , \ctl_rf_c2dmabs_reg[29]/NET0131  , \ctl_rf_c2dmabs_reg[30]/NET0131  , \ctl_rf_c2dmabs_reg[31]/NET0131  , \ctl_rf_c3_rf_autold_reg/NET0131  , \ctl_rf_c3_rf_ch_en_reg/NET0131  , \ctl_rf_c3_rf_chabt_reg/NET0131  , \ctl_rf_c3_rf_chdad_reg[0]/NET0131  , \ctl_rf_c3_rf_chdad_reg[10]/NET0131  , \ctl_rf_c3_rf_chdad_reg[11]/NET0131  , \ctl_rf_c3_rf_chdad_reg[12]/NET0131  , \ctl_rf_c3_rf_chdad_reg[13]/P0002  , \ctl_rf_c3_rf_chdad_reg[14]/P0002  , \ctl_rf_c3_rf_chdad_reg[15]/NET0131  , \ctl_rf_c3_rf_chdad_reg[16]/NET0131  , \ctl_rf_c3_rf_chdad_reg[17]/NET0131  , \ctl_rf_c3_rf_chdad_reg[18]/NET0131  , \ctl_rf_c3_rf_chdad_reg[19]/NET0131  , \ctl_rf_c3_rf_chdad_reg[1]/NET0131  , \ctl_rf_c3_rf_chdad_reg[20]/P0002  , \ctl_rf_c3_rf_chdad_reg[21]/P0002  , \ctl_rf_c3_rf_chdad_reg[22]/P0002  , \ctl_rf_c3_rf_chdad_reg[23]/P0002  , \ctl_rf_c3_rf_chdad_reg[24]/P0002  , \ctl_rf_c3_rf_chdad_reg[25]/P0002  , \ctl_rf_c3_rf_chdad_reg[26]/P0002  , \ctl_rf_c3_rf_chdad_reg[27]/P0002  , \ctl_rf_c3_rf_chdad_reg[28]/P0002  , \ctl_rf_c3_rf_chdad_reg[29]/P0002  , \ctl_rf_c3_rf_chdad_reg[2]/NET0131  , \ctl_rf_c3_rf_chdad_reg[30]/P0002  , \ctl_rf_c3_rf_chdad_reg[31]/P0002  , \ctl_rf_c3_rf_chdad_reg[3]/P0002  , \ctl_rf_c3_rf_chdad_reg[4]/P0002  , \ctl_rf_c3_rf_chdad_reg[5]/P0002  , \ctl_rf_c3_rf_chdad_reg[6]/P0002  , \ctl_rf_c3_rf_chdad_reg[7]/P0002  , \ctl_rf_c3_rf_chdad_reg[8]/NET0131  , \ctl_rf_c3_rf_chdad_reg[9]/P0002  , \ctl_rf_c3_rf_chllp_cnt_reg[0]/NET0131  , \ctl_rf_c3_rf_chllp_cnt_reg[1]/NET0131  , \ctl_rf_c3_rf_chllp_cnt_reg[2]/NET0131  , \ctl_rf_c3_rf_chllp_cnt_reg[3]/NET0131  , \ctl_rf_c3_rf_chllp_on_reg/NET0131  , \ctl_rf_c3_rf_chllp_reg[0]/P0002  , \ctl_rf_c3_rf_chllp_reg[10]/NET0131  , \ctl_rf_c3_rf_chllp_reg[11]/NET0131  , \ctl_rf_c3_rf_chllp_reg[12]/NET0131  , \ctl_rf_c3_rf_chllp_reg[13]/NET0131  , \ctl_rf_c3_rf_chllp_reg[14]/NET0131  , \ctl_rf_c3_rf_chllp_reg[15]/NET0131  , \ctl_rf_c3_rf_chllp_reg[16]/NET0131  , \ctl_rf_c3_rf_chllp_reg[17]/NET0131  , \ctl_rf_c3_rf_chllp_reg[18]/NET0131  , \ctl_rf_c3_rf_chllp_reg[19]/NET0131  , \ctl_rf_c3_rf_chllp_reg[1]/P0002  , \ctl_rf_c3_rf_chllp_reg[20]/NET0131  , \ctl_rf_c3_rf_chllp_reg[21]/NET0131  , \ctl_rf_c3_rf_chllp_reg[22]/NET0131  , \ctl_rf_c3_rf_chllp_reg[23]/NET0131  , \ctl_rf_c3_rf_chllp_reg[24]/NET0131  , \ctl_rf_c3_rf_chllp_reg[25]/NET0131  , \ctl_rf_c3_rf_chllp_reg[26]/NET0131  , \ctl_rf_c3_rf_chllp_reg[27]/NET0131  , \ctl_rf_c3_rf_chllp_reg[28]/NET0131  , \ctl_rf_c3_rf_chllp_reg[29]/NET0131  , \ctl_rf_c3_rf_chllp_reg[2]/NET0131  , \ctl_rf_c3_rf_chllp_reg[30]/NET0131  , \ctl_rf_c3_rf_chllp_reg[31]/NET0131  , \ctl_rf_c3_rf_chllp_reg[3]/NET0131  , \ctl_rf_c3_rf_chllp_reg[4]/NET0131  , \ctl_rf_c3_rf_chllp_reg[5]/NET0131  , \ctl_rf_c3_rf_chllp_reg[6]/NET0131  , \ctl_rf_c3_rf_chllp_reg[7]/NET0131  , \ctl_rf_c3_rf_chllp_reg[8]/NET0131  , \ctl_rf_c3_rf_chllp_reg[9]/NET0131  , \ctl_rf_c3_rf_chllpen_reg/NET0131  , \ctl_rf_c3_rf_chpri_reg[0]/NET0131  , \ctl_rf_c3_rf_chpri_reg[1]/NET0131  , \ctl_rf_c3_rf_chsad_reg[0]/NET0131  , \ctl_rf_c3_rf_chsad_reg[10]/P0002  , \ctl_rf_c3_rf_chsad_reg[11]/P0002  , \ctl_rf_c3_rf_chsad_reg[12]/P0002  , \ctl_rf_c3_rf_chsad_reg[13]/NET0131  , \ctl_rf_c3_rf_chsad_reg[14]/NET0131  , \ctl_rf_c3_rf_chsad_reg[15]/P0002  , \ctl_rf_c3_rf_chsad_reg[16]/NET0131  , \ctl_rf_c3_rf_chsad_reg[17]/NET0131  , \ctl_rf_c3_rf_chsad_reg[18]/NET0131  , \ctl_rf_c3_rf_chsad_reg[19]/NET0131  , \ctl_rf_c3_rf_chsad_reg[1]/NET0131  , \ctl_rf_c3_rf_chsad_reg[20]/NET0131  , \ctl_rf_c3_rf_chsad_reg[21]/NET0131  , \ctl_rf_c3_rf_chsad_reg[22]/NET0131  , \ctl_rf_c3_rf_chsad_reg[23]/NET0131  , \ctl_rf_c3_rf_chsad_reg[24]/NET0131  , \ctl_rf_c3_rf_chsad_reg[25]/P0002  , \ctl_rf_c3_rf_chsad_reg[26]/P0002  , \ctl_rf_c3_rf_chsad_reg[27]/P0002  , \ctl_rf_c3_rf_chsad_reg[28]/P0002  , \ctl_rf_c3_rf_chsad_reg[29]/P0002  , \ctl_rf_c3_rf_chsad_reg[2]/NET0131  , \ctl_rf_c3_rf_chsad_reg[30]/P0002  , \ctl_rf_c3_rf_chsad_reg[31]/NET0131  , \ctl_rf_c3_rf_chsad_reg[3]/NET0131  , \ctl_rf_c3_rf_chsad_reg[4]/NET0131  , \ctl_rf_c3_rf_chsad_reg[5]/NET0131  , \ctl_rf_c3_rf_chsad_reg[6]/NET0131  , \ctl_rf_c3_rf_chsad_reg[7]/NET0131  , \ctl_rf_c3_rf_chsad_reg[8]/P0002  , \ctl_rf_c3_rf_chsad_reg[9]/NET0131  , \ctl_rf_c3_rf_chtsz_reg[0]/P0002  , \ctl_rf_c3_rf_chtsz_reg[10]/P0002  , \ctl_rf_c3_rf_chtsz_reg[11]/P0002  , \ctl_rf_c3_rf_chtsz_reg[1]/P0002  , \ctl_rf_c3_rf_chtsz_reg[2]/P0002  , \ctl_rf_c3_rf_chtsz_reg[3]/P0002  , \ctl_rf_c3_rf_chtsz_reg[4]/NET0131  , \ctl_rf_c3_rf_chtsz_reg[5]/NET0131  , \ctl_rf_c3_rf_chtsz_reg[6]/NET0131  , \ctl_rf_c3_rf_chtsz_reg[7]/NET0131  , \ctl_rf_c3_rf_chtsz_reg[8]/P0002  , \ctl_rf_c3_rf_chtsz_reg[9]/P0002  , \ctl_rf_c3_rf_dad_ctl0_reg/NET0131  , \ctl_rf_c3_rf_dad_ctl1_reg/NET0131  , \ctl_rf_c3_rf_dreqmode_reg/NET0131  , \ctl_rf_c3_rf_dst_sel_reg/NET0131  , \ctl_rf_c3_rf_dwidth_reg[0]/NET0131  , \ctl_rf_c3_rf_dwidth_reg[1]/NET0131  , \ctl_rf_c3_rf_dwidth_reg[2]/NET0131  , \ctl_rf_c3_rf_int_abt_msk_reg/NET0131  , \ctl_rf_c3_rf_int_err_msk_reg/NET0131  , \ctl_rf_c3_rf_int_tc1_msk_reg/NET0131  , \ctl_rf_c3_rf_int_tc_msk_reg/NET0131  , \ctl_rf_c3_rf_mode_reg/NET0131  , \ctl_rf_c3_rf_prot1_reg/NET0131  , \ctl_rf_c3_rf_prot2_reg/NET0131  , \ctl_rf_c3_rf_prot3_reg/NET0131  , \ctl_rf_c3_rf_sad_ctl0_reg/NET0131  , \ctl_rf_c3_rf_sad_ctl1_reg/NET0131  , \ctl_rf_c3_rf_src_sel_reg/NET0131  , \ctl_rf_c3_rf_src_sz_reg[0]/NET0131  , \ctl_rf_c3_rf_src_sz_reg[1]/NET0131  , \ctl_rf_c3_rf_src_sz_reg[2]/NET0131  , \ctl_rf_c3_rf_swidth_reg[0]/NET0131  , \ctl_rf_c3_rf_swidth_reg[1]/NET0131  , \ctl_rf_c3_rf_swidth_reg[2]/NET0131  , \ctl_rf_c3brbs_reg[16]/NET0131  , \ctl_rf_c3brbs_reg[17]/NET0131  , \ctl_rf_c3brbs_reg[18]/NET0131  , \ctl_rf_c3brbs_reg[19]/NET0131  , \ctl_rf_c3brbs_reg[20]/NET0131  , \ctl_rf_c3brbs_reg[21]/NET0131  , \ctl_rf_c3brbs_reg[22]/NET0131  , \ctl_rf_c3brbs_reg[23]/NET0131  , \ctl_rf_c3brbs_reg[24]/NET0131  , \ctl_rf_c3brbs_reg[25]/NET0131  , \ctl_rf_c3brbs_reg[26]/NET0131  , \ctl_rf_c3brbs_reg[27]/NET0131  , \ctl_rf_c3brbs_reg[28]/NET0131  , \ctl_rf_c3brbs_reg[29]/NET0131  , \ctl_rf_c3brbs_reg[30]/NET0131  , \ctl_rf_c3brbs_reg[31]/NET0131  , \ctl_rf_c3dmabs_reg[16]/NET0131  , \ctl_rf_c3dmabs_reg[17]/NET0131  , \ctl_rf_c3dmabs_reg[18]/NET0131  , \ctl_rf_c3dmabs_reg[19]/NET0131  , \ctl_rf_c3dmabs_reg[20]/NET0131  , \ctl_rf_c3dmabs_reg[21]/NET0131  , \ctl_rf_c3dmabs_reg[22]/NET0131  , \ctl_rf_c3dmabs_reg[23]/NET0131  , \ctl_rf_c3dmabs_reg[24]/NET0131  , \ctl_rf_c3dmabs_reg[25]/NET0131  , \ctl_rf_c3dmabs_reg[26]/NET0131  , \ctl_rf_c3dmabs_reg[27]/NET0131  , \ctl_rf_c3dmabs_reg[28]/NET0131  , \ctl_rf_c3dmabs_reg[29]/NET0131  , \ctl_rf_c3dmabs_reg[30]/NET0131  , \ctl_rf_c3dmabs_reg[31]/NET0131  , \ctl_rf_c4_rf_autold_reg/NET0131  , \ctl_rf_c4_rf_ch_en_reg/NET0131  , \ctl_rf_c4_rf_chabt_reg/NET0131  , \ctl_rf_c4_rf_chdad_reg[0]/NET0131  , \ctl_rf_c4_rf_chdad_reg[10]/P0002  , \ctl_rf_c4_rf_chdad_reg[11]/P0002  , \ctl_rf_c4_rf_chdad_reg[12]/P0002  , \ctl_rf_c4_rf_chdad_reg[13]/P0002  , \ctl_rf_c4_rf_chdad_reg[14]/P0002  , \ctl_rf_c4_rf_chdad_reg[15]/P0002  , \ctl_rf_c4_rf_chdad_reg[16]/NET0131  , \ctl_rf_c4_rf_chdad_reg[17]/NET0131  , \ctl_rf_c4_rf_chdad_reg[18]/NET0131  , \ctl_rf_c4_rf_chdad_reg[19]/NET0131  , \ctl_rf_c4_rf_chdad_reg[1]/NET0131  , \ctl_rf_c4_rf_chdad_reg[20]/P0002  , \ctl_rf_c4_rf_chdad_reg[21]/P0002  , \ctl_rf_c4_rf_chdad_reg[22]/P0002  , \ctl_rf_c4_rf_chdad_reg[23]/P0002  , \ctl_rf_c4_rf_chdad_reg[24]/P0002  , \ctl_rf_c4_rf_chdad_reg[25]/P0002  , \ctl_rf_c4_rf_chdad_reg[26]/P0002  , \ctl_rf_c4_rf_chdad_reg[27]/P0002  , \ctl_rf_c4_rf_chdad_reg[28]/P0002  , \ctl_rf_c4_rf_chdad_reg[29]/P0002  , \ctl_rf_c4_rf_chdad_reg[2]/NET0131  , \ctl_rf_c4_rf_chdad_reg[30]/P0002  , \ctl_rf_c4_rf_chdad_reg[31]/P0002  , \ctl_rf_c4_rf_chdad_reg[3]/P0002  , \ctl_rf_c4_rf_chdad_reg[4]/P0002  , \ctl_rf_c4_rf_chdad_reg[5]/P0002  , \ctl_rf_c4_rf_chdad_reg[6]/P0002  , \ctl_rf_c4_rf_chdad_reg[7]/P0002  , \ctl_rf_c4_rf_chdad_reg[8]/NET0131  , \ctl_rf_c4_rf_chdad_reg[9]/P0002  , \ctl_rf_c4_rf_chllp_cnt_reg[0]/NET0131  , \ctl_rf_c4_rf_chllp_cnt_reg[1]/NET0131  , \ctl_rf_c4_rf_chllp_cnt_reg[2]/NET0131  , \ctl_rf_c4_rf_chllp_cnt_reg[3]/NET0131  , \ctl_rf_c4_rf_chllp_on_reg/NET0131  , \ctl_rf_c4_rf_chllp_reg[0]/P0002  , \ctl_rf_c4_rf_chllp_reg[10]/NET0131  , \ctl_rf_c4_rf_chllp_reg[11]/NET0131  , \ctl_rf_c4_rf_chllp_reg[12]/NET0131  , \ctl_rf_c4_rf_chllp_reg[13]/NET0131  , \ctl_rf_c4_rf_chllp_reg[14]/NET0131  , \ctl_rf_c4_rf_chllp_reg[15]/NET0131  , \ctl_rf_c4_rf_chllp_reg[16]/NET0131  , \ctl_rf_c4_rf_chllp_reg[17]/NET0131  , \ctl_rf_c4_rf_chllp_reg[18]/NET0131  , \ctl_rf_c4_rf_chllp_reg[19]/NET0131  , \ctl_rf_c4_rf_chllp_reg[1]/P0002  , \ctl_rf_c4_rf_chllp_reg[20]/NET0131  , \ctl_rf_c4_rf_chllp_reg[21]/NET0131  , \ctl_rf_c4_rf_chllp_reg[22]/NET0131  , \ctl_rf_c4_rf_chllp_reg[23]/NET0131  , \ctl_rf_c4_rf_chllp_reg[24]/NET0131  , \ctl_rf_c4_rf_chllp_reg[25]/NET0131  , \ctl_rf_c4_rf_chllp_reg[26]/NET0131  , \ctl_rf_c4_rf_chllp_reg[27]/NET0131  , \ctl_rf_c4_rf_chllp_reg[28]/NET0131  , \ctl_rf_c4_rf_chllp_reg[29]/NET0131  , \ctl_rf_c4_rf_chllp_reg[2]/NET0131  , \ctl_rf_c4_rf_chllp_reg[30]/NET0131  , \ctl_rf_c4_rf_chllp_reg[31]/NET0131  , \ctl_rf_c4_rf_chllp_reg[3]/NET0131  , \ctl_rf_c4_rf_chllp_reg[4]/NET0131  , \ctl_rf_c4_rf_chllp_reg[5]/NET0131  , \ctl_rf_c4_rf_chllp_reg[6]/NET0131  , \ctl_rf_c4_rf_chllp_reg[7]/NET0131  , \ctl_rf_c4_rf_chllp_reg[8]/NET0131  , \ctl_rf_c4_rf_chllp_reg[9]/NET0131  , \ctl_rf_c4_rf_chllpen_reg/NET0131  , \ctl_rf_c4_rf_chpri_reg[0]/NET0131  , \ctl_rf_c4_rf_chpri_reg[1]/NET0131  , \ctl_rf_c4_rf_chsad_reg[0]/NET0131  , \ctl_rf_c4_rf_chsad_reg[10]/NET0131  , \ctl_rf_c4_rf_chsad_reg[11]/NET0131  , \ctl_rf_c4_rf_chsad_reg[12]/NET0131  , \ctl_rf_c4_rf_chsad_reg[13]/NET0131  , \ctl_rf_c4_rf_chsad_reg[14]/NET0131  , \ctl_rf_c4_rf_chsad_reg[15]/NET0131  , \ctl_rf_c4_rf_chsad_reg[16]/NET0131  , \ctl_rf_c4_rf_chsad_reg[17]/NET0131  , \ctl_rf_c4_rf_chsad_reg[18]/NET0131  , \ctl_rf_c4_rf_chsad_reg[19]/NET0131  , \ctl_rf_c4_rf_chsad_reg[1]/NET0131  , \ctl_rf_c4_rf_chsad_reg[20]/NET0131  , \ctl_rf_c4_rf_chsad_reg[21]/NET0131  , \ctl_rf_c4_rf_chsad_reg[22]/NET0131  , \ctl_rf_c4_rf_chsad_reg[23]/NET0131  , \ctl_rf_c4_rf_chsad_reg[24]/NET0131  , \ctl_rf_c4_rf_chsad_reg[25]/P0002  , \ctl_rf_c4_rf_chsad_reg[26]/P0002  , \ctl_rf_c4_rf_chsad_reg[27]/P0002  , \ctl_rf_c4_rf_chsad_reg[28]/P0002  , \ctl_rf_c4_rf_chsad_reg[29]/P0002  , \ctl_rf_c4_rf_chsad_reg[2]/NET0131  , \ctl_rf_c4_rf_chsad_reg[30]/P0002  , \ctl_rf_c4_rf_chsad_reg[31]/NET0131  , \ctl_rf_c4_rf_chsad_reg[3]/NET0131  , \ctl_rf_c4_rf_chsad_reg[4]/NET0131  , \ctl_rf_c4_rf_chsad_reg[5]/NET0131  , \ctl_rf_c4_rf_chsad_reg[6]/NET0131  , \ctl_rf_c4_rf_chsad_reg[7]/NET0131  , \ctl_rf_c4_rf_chsad_reg[8]/P0002  , \ctl_rf_c4_rf_chsad_reg[9]/NET0131  , \ctl_rf_c4_rf_chtsz_reg[0]/P0002  , \ctl_rf_c4_rf_chtsz_reg[10]/P0002  , \ctl_rf_c4_rf_chtsz_reg[11]/P0002  , \ctl_rf_c4_rf_chtsz_reg[1]/P0002  , \ctl_rf_c4_rf_chtsz_reg[2]/P0002  , \ctl_rf_c4_rf_chtsz_reg[3]/P0002  , \ctl_rf_c4_rf_chtsz_reg[4]/NET0131  , \ctl_rf_c4_rf_chtsz_reg[5]/NET0131  , \ctl_rf_c4_rf_chtsz_reg[6]/NET0131  , \ctl_rf_c4_rf_chtsz_reg[7]/NET0131  , \ctl_rf_c4_rf_chtsz_reg[8]/P0002  , \ctl_rf_c4_rf_chtsz_reg[9]/P0002  , \ctl_rf_c4_rf_dad_ctl0_reg/NET0131  , \ctl_rf_c4_rf_dad_ctl1_reg/NET0131  , \ctl_rf_c4_rf_dreqmode_reg/NET0131  , \ctl_rf_c4_rf_dst_sel_reg/NET0131  , \ctl_rf_c4_rf_dwidth_reg[0]/NET0131  , \ctl_rf_c4_rf_dwidth_reg[1]/NET0131  , \ctl_rf_c4_rf_dwidth_reg[2]/NET0131  , \ctl_rf_c4_rf_int_abt_msk_reg/NET0131  , \ctl_rf_c4_rf_int_err_msk_reg/NET0131  , \ctl_rf_c4_rf_int_tc1_msk_reg/NET0131  , \ctl_rf_c4_rf_int_tc_msk_reg/NET0131  , \ctl_rf_c4_rf_mode_reg/NET0131  , \ctl_rf_c4_rf_prot1_reg/NET0131  , \ctl_rf_c4_rf_prot2_reg/NET0131  , \ctl_rf_c4_rf_prot3_reg/NET0131  , \ctl_rf_c4_rf_sad_ctl0_reg/NET0131  , \ctl_rf_c4_rf_sad_ctl1_reg/NET0131  , \ctl_rf_c4_rf_src_sel_reg/NET0131  , \ctl_rf_c4_rf_src_sz_reg[0]/NET0131  , \ctl_rf_c4_rf_src_sz_reg[1]/NET0131  , \ctl_rf_c4_rf_src_sz_reg[2]/NET0131  , \ctl_rf_c4_rf_swidth_reg[0]/NET0131  , \ctl_rf_c4_rf_swidth_reg[1]/NET0131  , \ctl_rf_c4_rf_swidth_reg[2]/NET0131  , \ctl_rf_c4brbs_reg[16]/NET0131  , \ctl_rf_c4brbs_reg[17]/NET0131  , \ctl_rf_c4brbs_reg[18]/NET0131  , \ctl_rf_c4brbs_reg[19]/NET0131  , \ctl_rf_c4brbs_reg[20]/NET0131  , \ctl_rf_c4brbs_reg[21]/NET0131  , \ctl_rf_c4brbs_reg[22]/NET0131  , \ctl_rf_c4brbs_reg[23]/NET0131  , \ctl_rf_c4brbs_reg[24]/NET0131  , \ctl_rf_c4brbs_reg[25]/NET0131  , \ctl_rf_c4brbs_reg[26]/NET0131  , \ctl_rf_c4brbs_reg[27]/NET0131  , \ctl_rf_c4brbs_reg[28]/NET0131  , \ctl_rf_c4brbs_reg[29]/NET0131  , \ctl_rf_c4brbs_reg[30]/NET0131  , \ctl_rf_c4brbs_reg[31]/NET0131  , \ctl_rf_c4dmabs_reg[16]/NET0131  , \ctl_rf_c4dmabs_reg[17]/NET0131  , \ctl_rf_c4dmabs_reg[18]/NET0131  , \ctl_rf_c4dmabs_reg[19]/NET0131  , \ctl_rf_c4dmabs_reg[20]/NET0131  , \ctl_rf_c4dmabs_reg[21]/NET0131  , \ctl_rf_c4dmabs_reg[22]/NET0131  , \ctl_rf_c4dmabs_reg[23]/NET0131  , \ctl_rf_c4dmabs_reg[24]/NET0131  , \ctl_rf_c4dmabs_reg[25]/NET0131  , \ctl_rf_c4dmabs_reg[26]/NET0131  , \ctl_rf_c4dmabs_reg[27]/NET0131  , \ctl_rf_c4dmabs_reg[28]/NET0131  , \ctl_rf_c4dmabs_reg[29]/NET0131  , \ctl_rf_c4dmabs_reg[30]/NET0131  , \ctl_rf_c4dmabs_reg[31]/NET0131  , \ctl_rf_c5_rf_autold_reg/NET0131  , \ctl_rf_c5_rf_ch_en_reg/NET0131  , \ctl_rf_c5_rf_chabt_reg/NET0131  , \ctl_rf_c5_rf_chdad_reg[0]/NET0131  , \ctl_rf_c5_rf_chdad_reg[10]/P0002  , \ctl_rf_c5_rf_chdad_reg[11]/P0002  , \ctl_rf_c5_rf_chdad_reg[12]/P0002  , \ctl_rf_c5_rf_chdad_reg[13]/NET0131  , \ctl_rf_c5_rf_chdad_reg[14]/P0002  , \ctl_rf_c5_rf_chdad_reg[15]/P0002  , \ctl_rf_c5_rf_chdad_reg[16]/NET0131  , \ctl_rf_c5_rf_chdad_reg[17]/NET0131  , \ctl_rf_c5_rf_chdad_reg[18]/NET0131  , \ctl_rf_c5_rf_chdad_reg[19]/NET0131  , \ctl_rf_c5_rf_chdad_reg[1]/NET0131  , \ctl_rf_c5_rf_chdad_reg[20]/P0002  , \ctl_rf_c5_rf_chdad_reg[21]/P0002  , \ctl_rf_c5_rf_chdad_reg[22]/P0002  , \ctl_rf_c5_rf_chdad_reg[23]/P0002  , \ctl_rf_c5_rf_chdad_reg[24]/P0002  , \ctl_rf_c5_rf_chdad_reg[25]/P0002  , \ctl_rf_c5_rf_chdad_reg[26]/P0002  , \ctl_rf_c5_rf_chdad_reg[27]/P0002  , \ctl_rf_c5_rf_chdad_reg[28]/P0002  , \ctl_rf_c5_rf_chdad_reg[29]/P0002  , \ctl_rf_c5_rf_chdad_reg[2]/NET0131  , \ctl_rf_c5_rf_chdad_reg[30]/P0002  , \ctl_rf_c5_rf_chdad_reg[31]/P0002  , \ctl_rf_c5_rf_chdad_reg[3]/P0002  , \ctl_rf_c5_rf_chdad_reg[4]/P0002  , \ctl_rf_c5_rf_chdad_reg[5]/P0002  , \ctl_rf_c5_rf_chdad_reg[6]/P0002  , \ctl_rf_c5_rf_chdad_reg[7]/P0002  , \ctl_rf_c5_rf_chdad_reg[8]/NET0131  , \ctl_rf_c5_rf_chdad_reg[9]/P0002  , \ctl_rf_c5_rf_chllp_cnt_reg[0]/NET0131  , \ctl_rf_c5_rf_chllp_cnt_reg[1]/NET0131  , \ctl_rf_c5_rf_chllp_cnt_reg[2]/NET0131  , \ctl_rf_c5_rf_chllp_cnt_reg[3]/NET0131  , \ctl_rf_c5_rf_chllp_on_reg/NET0131  , \ctl_rf_c5_rf_chllp_reg[0]/P0002  , \ctl_rf_c5_rf_chllp_reg[10]/NET0131  , \ctl_rf_c5_rf_chllp_reg[11]/NET0131  , \ctl_rf_c5_rf_chllp_reg[12]/NET0131  , \ctl_rf_c5_rf_chllp_reg[13]/NET0131  , \ctl_rf_c5_rf_chllp_reg[14]/NET0131  , \ctl_rf_c5_rf_chllp_reg[15]/NET0131  , \ctl_rf_c5_rf_chllp_reg[16]/NET0131  , \ctl_rf_c5_rf_chllp_reg[17]/NET0131  , \ctl_rf_c5_rf_chllp_reg[18]/NET0131  , \ctl_rf_c5_rf_chllp_reg[19]/NET0131  , \ctl_rf_c5_rf_chllp_reg[1]/P0002  , \ctl_rf_c5_rf_chllp_reg[20]/NET0131  , \ctl_rf_c5_rf_chllp_reg[21]/NET0131  , \ctl_rf_c5_rf_chllp_reg[22]/NET0131  , \ctl_rf_c5_rf_chllp_reg[23]/NET0131  , \ctl_rf_c5_rf_chllp_reg[24]/NET0131  , \ctl_rf_c5_rf_chllp_reg[25]/NET0131  , \ctl_rf_c5_rf_chllp_reg[26]/NET0131  , \ctl_rf_c5_rf_chllp_reg[27]/NET0131  , \ctl_rf_c5_rf_chllp_reg[28]/NET0131  , \ctl_rf_c5_rf_chllp_reg[29]/NET0131  , \ctl_rf_c5_rf_chllp_reg[2]/NET0131  , \ctl_rf_c5_rf_chllp_reg[30]/NET0131  , \ctl_rf_c5_rf_chllp_reg[31]/NET0131  , \ctl_rf_c5_rf_chllp_reg[3]/NET0131  , \ctl_rf_c5_rf_chllp_reg[4]/NET0131  , \ctl_rf_c5_rf_chllp_reg[5]/NET0131  , \ctl_rf_c5_rf_chllp_reg[6]/NET0131  , \ctl_rf_c5_rf_chllp_reg[7]/NET0131  , \ctl_rf_c5_rf_chllp_reg[8]/NET0131  , \ctl_rf_c5_rf_chllp_reg[9]/NET0131  , \ctl_rf_c5_rf_chllpen_reg/NET0131  , \ctl_rf_c5_rf_chpri_reg[0]/NET0131  , \ctl_rf_c5_rf_chpri_reg[1]/NET0131  , \ctl_rf_c5_rf_chsad_reg[0]/NET0131  , \ctl_rf_c5_rf_chsad_reg[10]/NET0131  , \ctl_rf_c5_rf_chsad_reg[11]/NET0131  , \ctl_rf_c5_rf_chsad_reg[12]/NET0131  , \ctl_rf_c5_rf_chsad_reg[13]/P0002  , \ctl_rf_c5_rf_chsad_reg[14]/NET0131  , \ctl_rf_c5_rf_chsad_reg[15]/NET0131  , \ctl_rf_c5_rf_chsad_reg[16]/NET0131  , \ctl_rf_c5_rf_chsad_reg[17]/NET0131  , \ctl_rf_c5_rf_chsad_reg[18]/NET0131  , \ctl_rf_c5_rf_chsad_reg[19]/NET0131  , \ctl_rf_c5_rf_chsad_reg[1]/NET0131  , \ctl_rf_c5_rf_chsad_reg[20]/NET0131  , \ctl_rf_c5_rf_chsad_reg[21]/NET0131  , \ctl_rf_c5_rf_chsad_reg[22]/NET0131  , \ctl_rf_c5_rf_chsad_reg[23]/NET0131  , \ctl_rf_c5_rf_chsad_reg[24]/NET0131  , \ctl_rf_c5_rf_chsad_reg[25]/P0002  , \ctl_rf_c5_rf_chsad_reg[26]/P0002  , \ctl_rf_c5_rf_chsad_reg[27]/P0002  , \ctl_rf_c5_rf_chsad_reg[28]/P0002  , \ctl_rf_c5_rf_chsad_reg[29]/P0002  , \ctl_rf_c5_rf_chsad_reg[2]/NET0131  , \ctl_rf_c5_rf_chsad_reg[30]/P0002  , \ctl_rf_c5_rf_chsad_reg[31]/NET0131  , \ctl_rf_c5_rf_chsad_reg[3]/NET0131  , \ctl_rf_c5_rf_chsad_reg[4]/NET0131  , \ctl_rf_c5_rf_chsad_reg[5]/NET0131  , \ctl_rf_c5_rf_chsad_reg[6]/NET0131  , \ctl_rf_c5_rf_chsad_reg[7]/NET0131  , \ctl_rf_c5_rf_chsad_reg[8]/P0002  , \ctl_rf_c5_rf_chsad_reg[9]/NET0131  , \ctl_rf_c5_rf_chtsz_reg[0]/P0002  , \ctl_rf_c5_rf_chtsz_reg[10]/P0002  , \ctl_rf_c5_rf_chtsz_reg[11]/P0002  , \ctl_rf_c5_rf_chtsz_reg[1]/P0002  , \ctl_rf_c5_rf_chtsz_reg[2]/P0002  , \ctl_rf_c5_rf_chtsz_reg[3]/P0002  , \ctl_rf_c5_rf_chtsz_reg[4]/NET0131  , \ctl_rf_c5_rf_chtsz_reg[5]/NET0131  , \ctl_rf_c5_rf_chtsz_reg[6]/NET0131  , \ctl_rf_c5_rf_chtsz_reg[7]/NET0131  , \ctl_rf_c5_rf_chtsz_reg[8]/P0002  , \ctl_rf_c5_rf_chtsz_reg[9]/P0002  , \ctl_rf_c5_rf_dad_ctl0_reg/NET0131  , \ctl_rf_c5_rf_dad_ctl1_reg/NET0131  , \ctl_rf_c5_rf_dreqmode_reg/NET0131  , \ctl_rf_c5_rf_dst_sel_reg/NET0131  , \ctl_rf_c5_rf_dwidth_reg[0]/NET0131  , \ctl_rf_c5_rf_dwidth_reg[1]/NET0131  , \ctl_rf_c5_rf_dwidth_reg[2]/NET0131  , \ctl_rf_c5_rf_int_abt_msk_reg/NET0131  , \ctl_rf_c5_rf_int_err_msk_reg/NET0131  , \ctl_rf_c5_rf_int_tc1_msk_reg/NET0131  , \ctl_rf_c5_rf_int_tc_msk_reg/NET0131  , \ctl_rf_c5_rf_mode_reg/NET0131  , \ctl_rf_c5_rf_prot1_reg/NET0131  , \ctl_rf_c5_rf_prot2_reg/NET0131  , \ctl_rf_c5_rf_prot3_reg/NET0131  , \ctl_rf_c5_rf_sad_ctl0_reg/NET0131  , \ctl_rf_c5_rf_sad_ctl1_reg/NET0131  , \ctl_rf_c5_rf_src_sel_reg/NET0131  , \ctl_rf_c5_rf_src_sz_reg[0]/NET0131  , \ctl_rf_c5_rf_src_sz_reg[1]/NET0131  , \ctl_rf_c5_rf_src_sz_reg[2]/NET0131  , \ctl_rf_c5_rf_swidth_reg[0]/NET0131  , \ctl_rf_c5_rf_swidth_reg[1]/NET0131  , \ctl_rf_c5_rf_swidth_reg[2]/NET0131  , \ctl_rf_c5brbs_reg[16]/NET0131  , \ctl_rf_c5brbs_reg[17]/NET0131  , \ctl_rf_c5brbs_reg[18]/NET0131  , \ctl_rf_c5brbs_reg[19]/NET0131  , \ctl_rf_c5brbs_reg[20]/NET0131  , \ctl_rf_c5brbs_reg[21]/NET0131  , \ctl_rf_c5brbs_reg[22]/NET0131  , \ctl_rf_c5brbs_reg[23]/NET0131  , \ctl_rf_c5brbs_reg[24]/NET0131  , \ctl_rf_c5brbs_reg[25]/NET0131  , \ctl_rf_c5brbs_reg[26]/NET0131  , \ctl_rf_c5brbs_reg[27]/NET0131  , \ctl_rf_c5brbs_reg[28]/NET0131  , \ctl_rf_c5brbs_reg[29]/NET0131  , \ctl_rf_c5brbs_reg[30]/NET0131  , \ctl_rf_c5brbs_reg[31]/NET0131  , \ctl_rf_c5dmabs_reg[16]/NET0131  , \ctl_rf_c5dmabs_reg[17]/NET0131  , \ctl_rf_c5dmabs_reg[18]/NET0131  , \ctl_rf_c5dmabs_reg[19]/NET0131  , \ctl_rf_c5dmabs_reg[20]/NET0131  , \ctl_rf_c5dmabs_reg[21]/NET0131  , \ctl_rf_c5dmabs_reg[22]/NET0131  , \ctl_rf_c5dmabs_reg[23]/NET0131  , \ctl_rf_c5dmabs_reg[24]/NET0131  , \ctl_rf_c5dmabs_reg[25]/NET0131  , \ctl_rf_c5dmabs_reg[26]/NET0131  , \ctl_rf_c5dmabs_reg[27]/NET0131  , \ctl_rf_c5dmabs_reg[28]/NET0131  , \ctl_rf_c5dmabs_reg[29]/NET0131  , \ctl_rf_c5dmabs_reg[30]/NET0131  , \ctl_rf_c5dmabs_reg[31]/NET0131  , \ctl_rf_c6_rf_autold_reg/NET0131  , \ctl_rf_c6_rf_ch_en_reg/NET0131  , \ctl_rf_c6_rf_chabt_reg/NET0131  , \ctl_rf_c6_rf_chdad_reg[0]/NET0131  , \ctl_rf_c6_rf_chdad_reg[10]/NET0131  , \ctl_rf_c6_rf_chdad_reg[11]/P0002  , \ctl_rf_c6_rf_chdad_reg[12]/P0002  , \ctl_rf_c6_rf_chdad_reg[13]/NET0131  , \ctl_rf_c6_rf_chdad_reg[14]/P0002  , \ctl_rf_c6_rf_chdad_reg[15]/P0002  , \ctl_rf_c6_rf_chdad_reg[16]/NET0131  , \ctl_rf_c6_rf_chdad_reg[17]/NET0131  , \ctl_rf_c6_rf_chdad_reg[18]/NET0131  , \ctl_rf_c6_rf_chdad_reg[19]/NET0131  , \ctl_rf_c6_rf_chdad_reg[1]/NET0131  , \ctl_rf_c6_rf_chdad_reg[20]/P0002  , \ctl_rf_c6_rf_chdad_reg[21]/P0002  , \ctl_rf_c6_rf_chdad_reg[22]/P0002  , \ctl_rf_c6_rf_chdad_reg[23]/P0002  , \ctl_rf_c6_rf_chdad_reg[24]/P0002  , \ctl_rf_c6_rf_chdad_reg[25]/P0002  , \ctl_rf_c6_rf_chdad_reg[26]/P0002  , \ctl_rf_c6_rf_chdad_reg[27]/P0002  , \ctl_rf_c6_rf_chdad_reg[28]/P0002  , \ctl_rf_c6_rf_chdad_reg[29]/P0002  , \ctl_rf_c6_rf_chdad_reg[2]/NET0131  , \ctl_rf_c6_rf_chdad_reg[30]/P0002  , \ctl_rf_c6_rf_chdad_reg[31]/P0002  , \ctl_rf_c6_rf_chdad_reg[3]/P0002  , \ctl_rf_c6_rf_chdad_reg[4]/P0002  , \ctl_rf_c6_rf_chdad_reg[5]/P0002  , \ctl_rf_c6_rf_chdad_reg[6]/P0002  , \ctl_rf_c6_rf_chdad_reg[7]/P0002  , \ctl_rf_c6_rf_chdad_reg[8]/NET0131  , \ctl_rf_c6_rf_chdad_reg[9]/P0002  , \ctl_rf_c6_rf_chllp_cnt_reg[0]/NET0131  , \ctl_rf_c6_rf_chllp_cnt_reg[1]/NET0131  , \ctl_rf_c6_rf_chllp_cnt_reg[2]/NET0131  , \ctl_rf_c6_rf_chllp_cnt_reg[3]/NET0131  , \ctl_rf_c6_rf_chllp_on_reg/NET0131  , \ctl_rf_c6_rf_chllp_reg[0]/P0002  , \ctl_rf_c6_rf_chllp_reg[10]/NET0131  , \ctl_rf_c6_rf_chllp_reg[11]/NET0131  , \ctl_rf_c6_rf_chllp_reg[12]/NET0131  , \ctl_rf_c6_rf_chllp_reg[13]/NET0131  , \ctl_rf_c6_rf_chllp_reg[14]/NET0131  , \ctl_rf_c6_rf_chllp_reg[15]/NET0131  , \ctl_rf_c6_rf_chllp_reg[16]/NET0131  , \ctl_rf_c6_rf_chllp_reg[17]/NET0131  , \ctl_rf_c6_rf_chllp_reg[18]/NET0131  , \ctl_rf_c6_rf_chllp_reg[19]/NET0131  , \ctl_rf_c6_rf_chllp_reg[1]/P0002  , \ctl_rf_c6_rf_chllp_reg[20]/NET0131  , \ctl_rf_c6_rf_chllp_reg[21]/NET0131  , \ctl_rf_c6_rf_chllp_reg[22]/NET0131  , \ctl_rf_c6_rf_chllp_reg[23]/NET0131  , \ctl_rf_c6_rf_chllp_reg[24]/NET0131  , \ctl_rf_c6_rf_chllp_reg[25]/NET0131  , \ctl_rf_c6_rf_chllp_reg[26]/NET0131  , \ctl_rf_c6_rf_chllp_reg[27]/NET0131  , \ctl_rf_c6_rf_chllp_reg[28]/NET0131  , \ctl_rf_c6_rf_chllp_reg[29]/NET0131  , \ctl_rf_c6_rf_chllp_reg[2]/NET0131  , \ctl_rf_c6_rf_chllp_reg[30]/NET0131  , \ctl_rf_c6_rf_chllp_reg[31]/NET0131  , \ctl_rf_c6_rf_chllp_reg[3]/NET0131  , \ctl_rf_c6_rf_chllp_reg[4]/NET0131  , \ctl_rf_c6_rf_chllp_reg[5]/NET0131  , \ctl_rf_c6_rf_chllp_reg[6]/NET0131  , \ctl_rf_c6_rf_chllp_reg[7]/NET0131  , \ctl_rf_c6_rf_chllp_reg[8]/NET0131  , \ctl_rf_c6_rf_chllp_reg[9]/NET0131  , \ctl_rf_c6_rf_chllpen_reg/NET0131  , \ctl_rf_c6_rf_chpri_reg[0]/NET0131  , \ctl_rf_c6_rf_chpri_reg[1]/NET0131  , \ctl_rf_c6_rf_chsad_reg[0]/NET0131  , \ctl_rf_c6_rf_chsad_reg[10]/P0002  , \ctl_rf_c6_rf_chsad_reg[11]/NET0131  , \ctl_rf_c6_rf_chsad_reg[12]/NET0131  , \ctl_rf_c6_rf_chsad_reg[13]/P0002  , \ctl_rf_c6_rf_chsad_reg[14]/NET0131  , \ctl_rf_c6_rf_chsad_reg[15]/NET0131  , \ctl_rf_c6_rf_chsad_reg[16]/NET0131  , \ctl_rf_c6_rf_chsad_reg[17]/NET0131  , \ctl_rf_c6_rf_chsad_reg[18]/NET0131  , \ctl_rf_c6_rf_chsad_reg[19]/NET0131  , \ctl_rf_c6_rf_chsad_reg[1]/NET0131  , \ctl_rf_c6_rf_chsad_reg[20]/NET0131  , \ctl_rf_c6_rf_chsad_reg[21]/NET0131  , \ctl_rf_c6_rf_chsad_reg[22]/NET0131  , \ctl_rf_c6_rf_chsad_reg[23]/NET0131  , \ctl_rf_c6_rf_chsad_reg[24]/NET0131  , \ctl_rf_c6_rf_chsad_reg[25]/P0002  , \ctl_rf_c6_rf_chsad_reg[26]/P0002  , \ctl_rf_c6_rf_chsad_reg[27]/P0002  , \ctl_rf_c6_rf_chsad_reg[28]/P0002  , \ctl_rf_c6_rf_chsad_reg[29]/P0002  , \ctl_rf_c6_rf_chsad_reg[2]/NET0131  , \ctl_rf_c6_rf_chsad_reg[30]/P0002  , \ctl_rf_c6_rf_chsad_reg[31]/NET0131  , \ctl_rf_c6_rf_chsad_reg[3]/NET0131  , \ctl_rf_c6_rf_chsad_reg[4]/NET0131  , \ctl_rf_c6_rf_chsad_reg[5]/NET0131  , \ctl_rf_c6_rf_chsad_reg[6]/NET0131  , \ctl_rf_c6_rf_chsad_reg[7]/NET0131  , \ctl_rf_c6_rf_chsad_reg[8]/P0002  , \ctl_rf_c6_rf_chsad_reg[9]/NET0131  , \ctl_rf_c6_rf_chtsz_reg[0]/P0002  , \ctl_rf_c6_rf_chtsz_reg[10]/P0002  , \ctl_rf_c6_rf_chtsz_reg[11]/P0002  , \ctl_rf_c6_rf_chtsz_reg[1]/P0002  , \ctl_rf_c6_rf_chtsz_reg[2]/P0002  , \ctl_rf_c6_rf_chtsz_reg[3]/P0002  , \ctl_rf_c6_rf_chtsz_reg[4]/NET0131  , \ctl_rf_c6_rf_chtsz_reg[5]/NET0131  , \ctl_rf_c6_rf_chtsz_reg[6]/NET0131  , \ctl_rf_c6_rf_chtsz_reg[7]/NET0131  , \ctl_rf_c6_rf_chtsz_reg[8]/P0002  , \ctl_rf_c6_rf_chtsz_reg[9]/P0002  , \ctl_rf_c6_rf_dad_ctl0_reg/NET0131  , \ctl_rf_c6_rf_dad_ctl1_reg/NET0131  , \ctl_rf_c6_rf_dreqmode_reg/NET0131  , \ctl_rf_c6_rf_dst_sel_reg/NET0131  , \ctl_rf_c6_rf_dwidth_reg[0]/NET0131  , \ctl_rf_c6_rf_dwidth_reg[1]/NET0131  , \ctl_rf_c6_rf_dwidth_reg[2]/NET0131  , \ctl_rf_c6_rf_int_abt_msk_reg/NET0131  , \ctl_rf_c6_rf_int_err_msk_reg/NET0131  , \ctl_rf_c6_rf_int_tc1_msk_reg/NET0131  , \ctl_rf_c6_rf_int_tc_msk_reg/NET0131  , \ctl_rf_c6_rf_mode_reg/NET0131  , \ctl_rf_c6_rf_prot1_reg/NET0131  , \ctl_rf_c6_rf_prot2_reg/NET0131  , \ctl_rf_c6_rf_prot3_reg/NET0131  , \ctl_rf_c6_rf_sad_ctl0_reg/NET0131  , \ctl_rf_c6_rf_sad_ctl1_reg/NET0131  , \ctl_rf_c6_rf_src_sel_reg/NET0131  , \ctl_rf_c6_rf_src_sz_reg[0]/NET0131  , \ctl_rf_c6_rf_src_sz_reg[1]/NET0131  , \ctl_rf_c6_rf_src_sz_reg[2]/NET0131  , \ctl_rf_c6_rf_swidth_reg[0]/NET0131  , \ctl_rf_c6_rf_swidth_reg[1]/NET0131  , \ctl_rf_c6_rf_swidth_reg[2]/NET0131  , \ctl_rf_c6brbs_reg[16]/NET0131  , \ctl_rf_c6brbs_reg[17]/NET0131  , \ctl_rf_c6brbs_reg[18]/NET0131  , \ctl_rf_c6brbs_reg[19]/NET0131  , \ctl_rf_c6brbs_reg[20]/NET0131  , \ctl_rf_c6brbs_reg[21]/NET0131  , \ctl_rf_c6brbs_reg[22]/NET0131  , \ctl_rf_c6brbs_reg[23]/NET0131  , \ctl_rf_c6brbs_reg[24]/NET0131  , \ctl_rf_c6brbs_reg[25]/NET0131  , \ctl_rf_c6brbs_reg[26]/NET0131  , \ctl_rf_c6brbs_reg[27]/NET0131  , \ctl_rf_c6brbs_reg[28]/NET0131  , \ctl_rf_c6brbs_reg[29]/NET0131  , \ctl_rf_c6brbs_reg[30]/NET0131  , \ctl_rf_c6brbs_reg[31]/NET0131  , \ctl_rf_c6dmabs_reg[16]/NET0131  , \ctl_rf_c6dmabs_reg[17]/NET0131  , \ctl_rf_c6dmabs_reg[18]/NET0131  , \ctl_rf_c6dmabs_reg[19]/NET0131  , \ctl_rf_c6dmabs_reg[20]/NET0131  , \ctl_rf_c6dmabs_reg[21]/NET0131  , \ctl_rf_c6dmabs_reg[22]/NET0131  , \ctl_rf_c6dmabs_reg[23]/NET0131  , \ctl_rf_c6dmabs_reg[24]/NET0131  , \ctl_rf_c6dmabs_reg[25]/NET0131  , \ctl_rf_c6dmabs_reg[26]/NET0131  , \ctl_rf_c6dmabs_reg[27]/NET0131  , \ctl_rf_c6dmabs_reg[28]/NET0131  , \ctl_rf_c6dmabs_reg[29]/NET0131  , \ctl_rf_c6dmabs_reg[30]/NET0131  , \ctl_rf_c6dmabs_reg[31]/NET0131  , \ctl_rf_c7_rf_autold_reg/NET0131  , \ctl_rf_c7_rf_ch_en_reg/NET0131  , \ctl_rf_c7_rf_chabt_reg/NET0131  , \ctl_rf_c7_rf_chdad_reg[0]/NET0131  , \ctl_rf_c7_rf_chdad_reg[10]/P0002  , \ctl_rf_c7_rf_chdad_reg[11]/NET0131  , \ctl_rf_c7_rf_chdad_reg[12]/P0002  , \ctl_rf_c7_rf_chdad_reg[13]/NET0131  , \ctl_rf_c7_rf_chdad_reg[14]/NET0131  , \ctl_rf_c7_rf_chdad_reg[15]/NET0131  , \ctl_rf_c7_rf_chdad_reg[16]/NET0131  , \ctl_rf_c7_rf_chdad_reg[17]/NET0131  , \ctl_rf_c7_rf_chdad_reg[18]/NET0131  , \ctl_rf_c7_rf_chdad_reg[19]/NET0131  , \ctl_rf_c7_rf_chdad_reg[1]/NET0131  , \ctl_rf_c7_rf_chdad_reg[20]/P0002  , \ctl_rf_c7_rf_chdad_reg[21]/P0002  , \ctl_rf_c7_rf_chdad_reg[22]/P0002  , \ctl_rf_c7_rf_chdad_reg[23]/P0002  , \ctl_rf_c7_rf_chdad_reg[24]/P0002  , \ctl_rf_c7_rf_chdad_reg[25]/P0002  , \ctl_rf_c7_rf_chdad_reg[26]/P0002  , \ctl_rf_c7_rf_chdad_reg[27]/P0002  , \ctl_rf_c7_rf_chdad_reg[28]/P0002  , \ctl_rf_c7_rf_chdad_reg[29]/P0002  , \ctl_rf_c7_rf_chdad_reg[2]/NET0131  , \ctl_rf_c7_rf_chdad_reg[30]/P0002  , \ctl_rf_c7_rf_chdad_reg[31]/P0002  , \ctl_rf_c7_rf_chdad_reg[3]/P0002  , \ctl_rf_c7_rf_chdad_reg[4]/P0002  , \ctl_rf_c7_rf_chdad_reg[5]/P0002  , \ctl_rf_c7_rf_chdad_reg[6]/P0002  , \ctl_rf_c7_rf_chdad_reg[7]/P0002  , \ctl_rf_c7_rf_chdad_reg[8]/NET0131  , \ctl_rf_c7_rf_chdad_reg[9]/P0002  , \ctl_rf_c7_rf_chllp_cnt_reg[0]/NET0131  , \ctl_rf_c7_rf_chllp_cnt_reg[1]/NET0131  , \ctl_rf_c7_rf_chllp_cnt_reg[2]/NET0131  , \ctl_rf_c7_rf_chllp_cnt_reg[3]/NET0131  , \ctl_rf_c7_rf_chllp_on_reg/NET0131  , \ctl_rf_c7_rf_chllp_reg[0]/P0002  , \ctl_rf_c7_rf_chllp_reg[10]/NET0131  , \ctl_rf_c7_rf_chllp_reg[11]/NET0131  , \ctl_rf_c7_rf_chllp_reg[12]/NET0131  , \ctl_rf_c7_rf_chllp_reg[13]/NET0131  , \ctl_rf_c7_rf_chllp_reg[14]/NET0131  , \ctl_rf_c7_rf_chllp_reg[15]/NET0131  , \ctl_rf_c7_rf_chllp_reg[16]/NET0131  , \ctl_rf_c7_rf_chllp_reg[17]/NET0131  , \ctl_rf_c7_rf_chllp_reg[18]/NET0131  , \ctl_rf_c7_rf_chllp_reg[19]/NET0131  , \ctl_rf_c7_rf_chllp_reg[1]/P0002  , \ctl_rf_c7_rf_chllp_reg[20]/NET0131  , \ctl_rf_c7_rf_chllp_reg[21]/NET0131  , \ctl_rf_c7_rf_chllp_reg[22]/NET0131  , \ctl_rf_c7_rf_chllp_reg[23]/NET0131  , \ctl_rf_c7_rf_chllp_reg[24]/NET0131  , \ctl_rf_c7_rf_chllp_reg[25]/NET0131  , \ctl_rf_c7_rf_chllp_reg[26]/NET0131  , \ctl_rf_c7_rf_chllp_reg[27]/NET0131  , \ctl_rf_c7_rf_chllp_reg[28]/NET0131  , \ctl_rf_c7_rf_chllp_reg[29]/NET0131  , \ctl_rf_c7_rf_chllp_reg[2]/NET0131  , \ctl_rf_c7_rf_chllp_reg[30]/NET0131  , \ctl_rf_c7_rf_chllp_reg[31]/NET0131  , \ctl_rf_c7_rf_chllp_reg[3]/NET0131  , \ctl_rf_c7_rf_chllp_reg[4]/NET0131  , \ctl_rf_c7_rf_chllp_reg[5]/NET0131  , \ctl_rf_c7_rf_chllp_reg[6]/NET0131  , \ctl_rf_c7_rf_chllp_reg[7]/NET0131  , \ctl_rf_c7_rf_chllp_reg[8]/NET0131  , \ctl_rf_c7_rf_chllp_reg[9]/NET0131  , \ctl_rf_c7_rf_chllpen_reg/NET0131  , \ctl_rf_c7_rf_chpri_reg[0]/NET0131  , \ctl_rf_c7_rf_chpri_reg[1]/NET0131  , \ctl_rf_c7_rf_chsad_reg[0]/NET0131  , \ctl_rf_c7_rf_chsad_reg[10]/NET0131  , \ctl_rf_c7_rf_chsad_reg[11]/P0002  , \ctl_rf_c7_rf_chsad_reg[12]/NET0131  , \ctl_rf_c7_rf_chsad_reg[13]/P0002  , \ctl_rf_c7_rf_chsad_reg[14]/P0002  , \ctl_rf_c7_rf_chsad_reg[15]/P0002  , \ctl_rf_c7_rf_chsad_reg[16]/NET0131  , \ctl_rf_c7_rf_chsad_reg[17]/NET0131  , \ctl_rf_c7_rf_chsad_reg[18]/NET0131  , \ctl_rf_c7_rf_chsad_reg[19]/NET0131  , \ctl_rf_c7_rf_chsad_reg[1]/NET0131  , \ctl_rf_c7_rf_chsad_reg[20]/NET0131  , \ctl_rf_c7_rf_chsad_reg[21]/NET0131  , \ctl_rf_c7_rf_chsad_reg[22]/NET0131  , \ctl_rf_c7_rf_chsad_reg[23]/NET0131  , \ctl_rf_c7_rf_chsad_reg[24]/NET0131  , \ctl_rf_c7_rf_chsad_reg[25]/P0002  , \ctl_rf_c7_rf_chsad_reg[26]/P0002  , \ctl_rf_c7_rf_chsad_reg[27]/P0002  , \ctl_rf_c7_rf_chsad_reg[28]/P0002  , \ctl_rf_c7_rf_chsad_reg[29]/P0002  , \ctl_rf_c7_rf_chsad_reg[2]/NET0131  , \ctl_rf_c7_rf_chsad_reg[30]/P0002  , \ctl_rf_c7_rf_chsad_reg[31]/NET0131  , \ctl_rf_c7_rf_chsad_reg[3]/NET0131  , \ctl_rf_c7_rf_chsad_reg[4]/NET0131  , \ctl_rf_c7_rf_chsad_reg[5]/NET0131  , \ctl_rf_c7_rf_chsad_reg[6]/NET0131  , \ctl_rf_c7_rf_chsad_reg[7]/NET0131  , \ctl_rf_c7_rf_chsad_reg[8]/P0002  , \ctl_rf_c7_rf_chsad_reg[9]/NET0131  , \ctl_rf_c7_rf_chtsz_reg[0]/P0002  , \ctl_rf_c7_rf_chtsz_reg[10]/P0002  , \ctl_rf_c7_rf_chtsz_reg[11]/P0002  , \ctl_rf_c7_rf_chtsz_reg[1]/P0002  , \ctl_rf_c7_rf_chtsz_reg[2]/P0002  , \ctl_rf_c7_rf_chtsz_reg[3]/P0002  , \ctl_rf_c7_rf_chtsz_reg[4]/NET0131  , \ctl_rf_c7_rf_chtsz_reg[5]/NET0131  , \ctl_rf_c7_rf_chtsz_reg[6]/NET0131  , \ctl_rf_c7_rf_chtsz_reg[7]/NET0131  , \ctl_rf_c7_rf_chtsz_reg[8]/P0002  , \ctl_rf_c7_rf_chtsz_reg[9]/P0002  , \ctl_rf_c7_rf_dad_ctl0_reg/NET0131  , \ctl_rf_c7_rf_dad_ctl1_reg/NET0131  , \ctl_rf_c7_rf_dreqmode_reg/NET0131  , \ctl_rf_c7_rf_dst_sel_reg/NET0131  , \ctl_rf_c7_rf_dwidth_reg[0]/NET0131  , \ctl_rf_c7_rf_dwidth_reg[1]/NET0131  , \ctl_rf_c7_rf_dwidth_reg[2]/NET0131  , \ctl_rf_c7_rf_int_abt_msk_reg/NET0131  , \ctl_rf_c7_rf_int_err_msk_reg/NET0131  , \ctl_rf_c7_rf_int_tc1_msk_reg/NET0131  , \ctl_rf_c7_rf_int_tc_msk_reg/NET0131  , \ctl_rf_c7_rf_mode_reg/NET0131  , \ctl_rf_c7_rf_prot1_reg/NET0131  , \ctl_rf_c7_rf_prot2_reg/NET0131  , \ctl_rf_c7_rf_prot3_reg/NET0131  , \ctl_rf_c7_rf_sad_ctl0_reg/NET0131  , \ctl_rf_c7_rf_sad_ctl1_reg/NET0131  , \ctl_rf_c7_rf_src_sel_reg/NET0131  , \ctl_rf_c7_rf_src_sz_reg[0]/NET0131  , \ctl_rf_c7_rf_src_sz_reg[1]/NET0131  , \ctl_rf_c7_rf_src_sz_reg[2]/NET0131  , \ctl_rf_c7_rf_swidth_reg[0]/NET0131  , \ctl_rf_c7_rf_swidth_reg[1]/NET0131  , \ctl_rf_c7_rf_swidth_reg[2]/NET0131  , \ctl_rf_c7brbs_reg[16]/NET0131  , \ctl_rf_c7brbs_reg[17]/NET0131  , \ctl_rf_c7brbs_reg[18]/NET0131  , \ctl_rf_c7brbs_reg[19]/NET0131  , \ctl_rf_c7brbs_reg[20]/NET0131  , \ctl_rf_c7brbs_reg[21]/NET0131  , \ctl_rf_c7brbs_reg[22]/NET0131  , \ctl_rf_c7brbs_reg[23]/NET0131  , \ctl_rf_c7brbs_reg[24]/NET0131  , \ctl_rf_c7brbs_reg[25]/NET0131  , \ctl_rf_c7brbs_reg[26]/NET0131  , \ctl_rf_c7brbs_reg[27]/NET0131  , \ctl_rf_c7brbs_reg[28]/NET0131  , \ctl_rf_c7brbs_reg[29]/NET0131  , \ctl_rf_c7brbs_reg[30]/NET0131  , \ctl_rf_c7brbs_reg[31]/NET0131  , \ctl_rf_c7dmabs_reg[16]/NET0131  , \ctl_rf_c7dmabs_reg[17]/NET0131  , \ctl_rf_c7dmabs_reg[18]/NET0131  , \ctl_rf_c7dmabs_reg[19]/NET0131  , \ctl_rf_c7dmabs_reg[20]/NET0131  , \ctl_rf_c7dmabs_reg[21]/NET0131  , \ctl_rf_c7dmabs_reg[22]/NET0131  , \ctl_rf_c7dmabs_reg[23]/NET0131  , \ctl_rf_c7dmabs_reg[24]/NET0131  , \ctl_rf_c7dmabs_reg[25]/NET0131  , \ctl_rf_c7dmabs_reg[26]/NET0131  , \ctl_rf_c7dmabs_reg[27]/NET0131  , \ctl_rf_c7dmabs_reg[28]/NET0131  , \ctl_rf_c7dmabs_reg[29]/NET0131  , \ctl_rf_c7dmabs_reg[30]/NET0131  , \ctl_rf_c7dmabs_reg[31]/NET0131  , \ctl_rf_dmacen_reg/NET0131  , \ctl_rf_m0end_reg/NET0131  , \ctl_rf_m1end_reg/NET0131  , \ctl_rf_rf_sel_d1_reg/NET0131  , \ctl_rf_sync_reg[0]/NET0131  , \ctl_rf_sync_reg[1]/NET0131  , \ctl_rf_sync_reg[2]/NET0131  , \ctl_rf_sync_reg[3]/NET0131  , \ctl_rf_sync_reg[4]/NET0131  , \ctl_rf_sync_reg[5]/NET0131  , \ctl_rf_sync_reg[6]/NET0131  , \ctl_rf_sync_reg[7]/NET0131  , \ctl_rf_tc_reg[0]/NET0131  , \ctl_rf_tc_reg[1]/NET0131  , \ctl_rf_tc_reg[2]/NET0131  , \ctl_rf_tc_reg[3]/NET0131  , \ctl_rf_tc_reg[4]/NET0131  , \ctl_rf_tc_reg[5]/NET0131  , \ctl_rf_tc_reg[6]/NET0131  , \ctl_rf_tc_reg[7]/NET0131  , \de_bst_cnt_reg[0]/NET0131  , \de_bst_cnt_reg[2]/NET0131  , \de_bst_cnt_reg[3]/NET0131  , \de_bst_cnt_reg[4]/NET0131  , \de_bst_cnt_reg[5]/NET0131  , \de_bst_cnt_reg[6]/NET0131  , \de_bst_cnt_reg[7]/NET0131  , \de_bst_cnt_reg[8]/NET0131  , \de_de_st_reg[0]/NET0131  , \de_de_st_reg[1]/NET0131  , \de_de_st_reg[2]/NET0131  , \de_de_st_reg[5]/NET0131  , \de_de_st_reg[6]/NET0131  , \de_m0_arb_st_reg/NET0131  , \de_m0_is_llp_reg/NET0131  , \de_m1_arb_st_reg[0]/NET0131  , \de_m1_arb_st_reg[1]/NET0131  , \de_m1_is_llp_reg/NET0131  , \de_st_rd_msk_reg/NET0131  , \de_tsz_cnt_reg[0]/NET0131  , \de_tsz_cnt_reg[10]/NET0131  , \de_tsz_cnt_reg[11]/NET0131  , \de_tsz_cnt_reg[1]/NET0131  , \de_tsz_cnt_reg[2]/NET0131  , \de_tsz_cnt_reg[3]/NET0131  , \de_tsz_cnt_reg[4]/NET0131  , \de_tsz_cnt_reg[5]/NET0131  , \de_tsz_cnt_reg[6]/NET0131  , \de_tsz_cnt_reg[7]/NET0131  , \de_tsz_cnt_reg[8]/NET0131  , \de_tsz_cnt_reg[9]/NET0131  , \dma_ack[0]_pad  , \dma_ack[1]_pad  , \dma_ack[2]_pad  , \dma_ack[3]_pad  , \dma_ack[4]_pad  , \dma_ack[5]_pad  , \dma_ack[6]_pad  , \dma_ack[7]_pad  , \dma_tc[0]_pad  , \dma_tc[1]_pad  , \dma_tc[2]_pad  , \dma_tc[3]_pad  , \dma_tc[4]_pad  , \dma_tc[5]_pad  , \dma_tc[6]_pad  , \dma_tc[7]_pad  , \h0burst[0]_pad  , \h0grant_pad  , \h0readyin_pad  , \h0req_pad  , \h0resp[0]_pad  , \h0resp[1]_pad  , \h0write_pad  , \h1burst[0]_pad  , \h1prot[0]_pad  , \h1rdt0_br[0]_pad  , \h1rdt0_br[10]_pad  , \h1rdt0_br[11]_pad  , \h1rdt0_br[12]_pad  , \h1rdt0_br[13]_pad  , \h1rdt0_br[14]_pad  , \h1rdt0_br[15]_pad  , \h1rdt0_br[16]_pad  , \h1rdt0_br[17]_pad  , \h1rdt0_br[18]_pad  , \h1rdt0_br[19]_pad  , \h1rdt0_br[1]_pad  , \h1rdt0_br[20]_pad  , \h1rdt0_br[21]_pad  , \h1rdt0_br[22]_pad  , \h1rdt0_br[23]_pad  , \h1rdt0_br[24]_pad  , \h1rdt0_br[25]_pad  , \h1rdt0_br[26]_pad  , \h1rdt0_br[27]_pad  , \h1rdt0_br[28]_pad  , \h1rdt0_br[29]_pad  , \h1rdt0_br[2]_pad  , \h1rdt0_br[30]_pad  , \h1rdt0_br[31]_pad  , \h1rdt0_br[3]_pad  , \h1rdt0_br[4]_pad  , \h1rdt0_br[5]_pad  , \h1rdt0_br[6]_pad  , \h1rdt0_br[7]_pad  , \h1rdt0_br[8]_pad  , \h1rdt0_br[9]_pad  , \h1rdt0_dma[0]_pad  , \h1rdt0_dma[10]_pad  , \h1rdt0_dma[11]_pad  , \h1rdt0_dma[12]_pad  , \h1rdt0_dma[13]_pad  , \h1rdt0_dma[14]_pad  , \h1rdt0_dma[15]_pad  , \h1rdt0_dma[16]_pad  , \h1rdt0_dma[17]_pad  , \h1rdt0_dma[18]_pad  , \h1rdt0_dma[19]_pad  , \h1rdt0_dma[1]_pad  , \h1rdt0_dma[20]_pad  , \h1rdt0_dma[21]_pad  , \h1rdt0_dma[22]_pad  , \h1rdt0_dma[23]_pad  , \h1rdt0_dma[24]_pad  , \h1rdt0_dma[25]_pad  , \h1rdt0_dma[26]_pad  , \h1rdt0_dma[27]_pad  , \h1rdt0_dma[28]_pad  , \h1rdt0_dma[29]_pad  , \h1rdt0_dma[2]_pad  , \h1rdt0_dma[30]_pad  , \h1rdt0_dma[31]_pad  , \h1rdt0_dma[3]_pad  , \h1rdt0_dma[4]_pad  , \h1rdt0_dma[5]_pad  , \h1rdt0_dma[6]_pad  , \h1rdt0_dma[7]_pad  , \h1rdt0_dma[8]_pad  , \h1rdt0_dma[9]_pad  , \h1rdt1_br[0]_pad  , \h1rdt1_br[10]_pad  , \h1rdt1_br[11]_pad  , \h1rdt1_br[12]_pad  , \h1rdt1_br[13]_pad  , \h1rdt1_br[14]_pad  , \h1rdt1_br[15]_pad  , \h1rdt1_br[16]_pad  , \h1rdt1_br[17]_pad  , \h1rdt1_br[18]_pad  , \h1rdt1_br[19]_pad  , \h1rdt1_br[1]_pad  , \h1rdt1_br[20]_pad  , \h1rdt1_br[21]_pad  , \h1rdt1_br[22]_pad  , \h1rdt1_br[23]_pad  , \h1rdt1_br[24]_pad  , \h1rdt1_br[25]_pad  , \h1rdt1_br[26]_pad  , \h1rdt1_br[27]_pad  , \h1rdt1_br[28]_pad  , \h1rdt1_br[29]_pad  , \h1rdt1_br[2]_pad  , \h1rdt1_br[30]_pad  , \h1rdt1_br[31]_pad  , \h1rdt1_br[3]_pad  , \h1rdt1_br[4]_pad  , \h1rdt1_br[5]_pad  , \h1rdt1_br[6]_pad  , \h1rdt1_br[7]_pad  , \h1rdt1_br[8]_pad  , \h1rdt1_br[9]_pad  , \h1rdt1_dma[0]_pad  , \h1rdt1_dma[10]_pad  , \h1rdt1_dma[11]_pad  , \h1rdt1_dma[12]_pad  , \h1rdt1_dma[13]_pad  , \h1rdt1_dma[14]_pad  , \h1rdt1_dma[15]_pad  , \h1rdt1_dma[16]_pad  , \h1rdt1_dma[17]_pad  , \h1rdt1_dma[18]_pad  , \h1rdt1_dma[19]_pad  , \h1rdt1_dma[1]_pad  , \h1rdt1_dma[20]_pad  , \h1rdt1_dma[21]_pad  , \h1rdt1_dma[22]_pad  , \h1rdt1_dma[23]_pad  , \h1rdt1_dma[24]_pad  , \h1rdt1_dma[25]_pad  , \h1rdt1_dma[26]_pad  , \h1rdt1_dma[27]_pad  , \h1rdt1_dma[28]_pad  , \h1rdt1_dma[29]_pad  , \h1rdt1_dma[2]_pad  , \h1rdt1_dma[30]_pad  , \h1rdt1_dma[31]_pad  , \h1rdt1_dma[3]_pad  , \h1rdt1_dma[4]_pad  , \h1rdt1_dma[5]_pad  , \h1rdt1_dma[6]_pad  , \h1rdt1_dma[7]_pad  , \h1rdt1_dma[8]_pad  , \h1rdt1_dma[9]_pad  , \h1rdt2_br[0]_pad  , \h1rdt2_br[10]_pad  , \h1rdt2_br[11]_pad  , \h1rdt2_br[12]_pad  , \h1rdt2_br[13]_pad  , \h1rdt2_br[14]_pad  , \h1rdt2_br[15]_pad  , \h1rdt2_br[16]_pad  , \h1rdt2_br[17]_pad  , \h1rdt2_br[18]_pad  , \h1rdt2_br[19]_pad  , \h1rdt2_br[1]_pad  , \h1rdt2_br[20]_pad  , \h1rdt2_br[21]_pad  , \h1rdt2_br[22]_pad  , \h1rdt2_br[23]_pad  , \h1rdt2_br[24]_pad  , \h1rdt2_br[25]_pad  , \h1rdt2_br[26]_pad  , \h1rdt2_br[27]_pad  , \h1rdt2_br[28]_pad  , \h1rdt2_br[29]_pad  , \h1rdt2_br[2]_pad  , \h1rdt2_br[30]_pad  , \h1rdt2_br[31]_pad  , \h1rdt2_br[3]_pad  , \h1rdt2_br[4]_pad  , \h1rdt2_br[5]_pad  , \h1rdt2_br[6]_pad  , \h1rdt2_br[7]_pad  , \h1rdt2_br[8]_pad  , \h1rdt2_br[9]_pad  , \h1rdt2_dma[0]_pad  , \h1rdt2_dma[10]_pad  , \h1rdt2_dma[11]_pad  , \h1rdt2_dma[12]_pad  , \h1rdt2_dma[13]_pad  , \h1rdt2_dma[14]_pad  , \h1rdt2_dma[15]_pad  , \h1rdt2_dma[16]_pad  , \h1rdt2_dma[17]_pad  , \h1rdt2_dma[18]_pad  , \h1rdt2_dma[19]_pad  , \h1rdt2_dma[1]_pad  , \h1rdt2_dma[20]_pad  , \h1rdt2_dma[21]_pad  , \h1rdt2_dma[22]_pad  , \h1rdt2_dma[23]_pad  , \h1rdt2_dma[24]_pad  , \h1rdt2_dma[25]_pad  , \h1rdt2_dma[26]_pad  , \h1rdt2_dma[27]_pad  , \h1rdt2_dma[28]_pad  , \h1rdt2_dma[29]_pad  , \h1rdt2_dma[2]_pad  , \h1rdt2_dma[30]_pad  , \h1rdt2_dma[31]_pad  , \h1rdt2_dma[3]_pad  , \h1rdt2_dma[4]_pad  , \h1rdt2_dma[5]_pad  , \h1rdt2_dma[6]_pad  , \h1rdt2_dma[7]_pad  , \h1rdt2_dma[8]_pad  , \h1rdt2_dma[9]_pad  , \h1rdt3_br[0]_pad  , \h1rdt3_br[10]_pad  , \h1rdt3_br[11]_pad  , \h1rdt3_br[12]_pad  , \h1rdt3_br[13]_pad  , \h1rdt3_br[14]_pad  , \h1rdt3_br[15]_pad  , \h1rdt3_br[16]_pad  , \h1rdt3_br[17]_pad  , \h1rdt3_br[18]_pad  , \h1rdt3_br[19]_pad  , \h1rdt3_br[1]_pad  , \h1rdt3_br[20]_pad  , \h1rdt3_br[21]_pad  , \h1rdt3_br[22]_pad  , \h1rdt3_br[23]_pad  , \h1rdt3_br[24]_pad  , \h1rdt3_br[25]_pad  , \h1rdt3_br[26]_pad  , \h1rdt3_br[27]_pad  , \h1rdt3_br[28]_pad  , \h1rdt3_br[29]_pad  , \h1rdt3_br[2]_pad  , \h1rdt3_br[30]_pad  , \h1rdt3_br[31]_pad  , \h1rdt3_br[3]_pad  , \h1rdt3_br[4]_pad  , \h1rdt3_br[5]_pad  , \h1rdt3_br[6]_pad  , \h1rdt3_br[7]_pad  , \h1rdt3_br[8]_pad  , \h1rdt3_br[9]_pad  , \h1rdt3_dma[0]_pad  , \h1rdt3_dma[10]_pad  , \h1rdt3_dma[11]_pad  , \h1rdt3_dma[12]_pad  , \h1rdt3_dma[13]_pad  , \h1rdt3_dma[14]_pad  , \h1rdt3_dma[15]_pad  , \h1rdt3_dma[16]_pad  , \h1rdt3_dma[17]_pad  , \h1rdt3_dma[18]_pad  , \h1rdt3_dma[19]_pad  , \h1rdt3_dma[1]_pad  , \h1rdt3_dma[20]_pad  , \h1rdt3_dma[21]_pad  , \h1rdt3_dma[22]_pad  , \h1rdt3_dma[23]_pad  , \h1rdt3_dma[24]_pad  , \h1rdt3_dma[25]_pad  , \h1rdt3_dma[26]_pad  , \h1rdt3_dma[27]_pad  , \h1rdt3_dma[28]_pad  , \h1rdt3_dma[29]_pad  , \h1rdt3_dma[2]_pad  , \h1rdt3_dma[30]_pad  , \h1rdt3_dma[31]_pad  , \h1rdt3_dma[3]_pad  , \h1rdt3_dma[4]_pad  , \h1rdt3_dma[5]_pad  , \h1rdt3_dma[6]_pad  , \h1rdt3_dma[7]_pad  , \h1rdt3_dma[8]_pad  , \h1rdt3_dma[9]_pad  , \h1rdt4_br[0]_pad  , \h1rdt4_br[10]_pad  , \h1rdt4_br[11]_pad  , \h1rdt4_br[12]_pad  , \h1rdt4_br[13]_pad  , \h1rdt4_br[14]_pad  , \h1rdt4_br[15]_pad  , \h1rdt4_br[16]_pad  , \h1rdt4_br[17]_pad  , \h1rdt4_br[18]_pad  , \h1rdt4_br[19]_pad  , \h1rdt4_br[1]_pad  , \h1rdt4_br[20]_pad  , \h1rdt4_br[21]_pad  , \h1rdt4_br[22]_pad  , \h1rdt4_br[23]_pad  , \h1rdt4_br[24]_pad  , \h1rdt4_br[25]_pad  , \h1rdt4_br[26]_pad  , \h1rdt4_br[27]_pad  , \h1rdt4_br[28]_pad  , \h1rdt4_br[29]_pad  , \h1rdt4_br[2]_pad  , \h1rdt4_br[30]_pad  , \h1rdt4_br[31]_pad  , \h1rdt4_br[3]_pad  , \h1rdt4_br[4]_pad  , \h1rdt4_br[5]_pad  , \h1rdt4_br[6]_pad  , \h1rdt4_br[7]_pad  , \h1rdt4_br[8]_pad  , \h1rdt4_br[9]_pad  , \h1rdt4_dma[0]_pad  , \h1rdt4_dma[10]_pad  , \h1rdt4_dma[11]_pad  , \h1rdt4_dma[12]_pad  , \h1rdt4_dma[13]_pad  , \h1rdt4_dma[14]_pad  , \h1rdt4_dma[15]_pad  , \h1rdt4_dma[16]_pad  , \h1rdt4_dma[17]_pad  , \h1rdt4_dma[18]_pad  , \h1rdt4_dma[19]_pad  , \h1rdt4_dma[1]_pad  , \h1rdt4_dma[20]_pad  , \h1rdt4_dma[21]_pad  , \h1rdt4_dma[22]_pad  , \h1rdt4_dma[23]_pad  , \h1rdt4_dma[24]_pad  , \h1rdt4_dma[25]_pad  , \h1rdt4_dma[26]_pad  , \h1rdt4_dma[27]_pad  , \h1rdt4_dma[28]_pad  , \h1rdt4_dma[29]_pad  , \h1rdt4_dma[2]_pad  , \h1rdt4_dma[30]_pad  , \h1rdt4_dma[31]_pad  , \h1rdt4_dma[3]_pad  , \h1rdt4_dma[4]_pad  , \h1rdt4_dma[5]_pad  , \h1rdt4_dma[6]_pad  , \h1rdt4_dma[7]_pad  , \h1rdt4_dma[8]_pad  , \h1rdt4_dma[9]_pad  , \h1rdt5_br[0]_pad  , \h1rdt5_br[10]_pad  , \h1rdt5_br[11]_pad  , \h1rdt5_br[12]_pad  , \h1rdt5_br[13]_pad  , \h1rdt5_br[14]_pad  , \h1rdt5_br[15]_pad  , \h1rdt5_br[16]_pad  , \h1rdt5_br[17]_pad  , \h1rdt5_br[18]_pad  , \h1rdt5_br[19]_pad  , \h1rdt5_br[1]_pad  , \h1rdt5_br[20]_pad  , \h1rdt5_br[21]_pad  , \h1rdt5_br[22]_pad  , \h1rdt5_br[23]_pad  , \h1rdt5_br[24]_pad  , \h1rdt5_br[25]_pad  , \h1rdt5_br[26]_pad  , \h1rdt5_br[27]_pad  , \h1rdt5_br[28]_pad  , \h1rdt5_br[29]_pad  , \h1rdt5_br[2]_pad  , \h1rdt5_br[30]_pad  , \h1rdt5_br[31]_pad  , \h1rdt5_br[3]_pad  , \h1rdt5_br[4]_pad  , \h1rdt5_br[5]_pad  , \h1rdt5_br[6]_pad  , \h1rdt5_br[7]_pad  , \h1rdt5_br[8]_pad  , \h1rdt5_br[9]_pad  , \h1rdt5_dma[0]_pad  , \h1rdt5_dma[10]_pad  , \h1rdt5_dma[11]_pad  , \h1rdt5_dma[12]_pad  , \h1rdt5_dma[13]_pad  , \h1rdt5_dma[14]_pad  , \h1rdt5_dma[15]_pad  , \h1rdt5_dma[16]_pad  , \h1rdt5_dma[17]_pad  , \h1rdt5_dma[18]_pad  , \h1rdt5_dma[19]_pad  , \h1rdt5_dma[1]_pad  , \h1rdt5_dma[20]_pad  , \h1rdt5_dma[21]_pad  , \h1rdt5_dma[22]_pad  , \h1rdt5_dma[23]_pad  , \h1rdt5_dma[24]_pad  , \h1rdt5_dma[25]_pad  , \h1rdt5_dma[26]_pad  , \h1rdt5_dma[27]_pad  , \h1rdt5_dma[28]_pad  , \h1rdt5_dma[29]_pad  , \h1rdt5_dma[2]_pad  , \h1rdt5_dma[30]_pad  , \h1rdt5_dma[31]_pad  , \h1rdt5_dma[3]_pad  , \h1rdt5_dma[4]_pad  , \h1rdt5_dma[5]_pad  , \h1rdt5_dma[6]_pad  , \h1rdt5_dma[7]_pad  , \h1rdt5_dma[8]_pad  , \h1rdt5_dma[9]_pad  , \h1rdt6_br[0]_pad  , \h1rdt6_br[10]_pad  , \h1rdt6_br[11]_pad  , \h1rdt6_br[12]_pad  , \h1rdt6_br[13]_pad  , \h1rdt6_br[14]_pad  , \h1rdt6_br[15]_pad  , \h1rdt6_br[16]_pad  , \h1rdt6_br[17]_pad  , \h1rdt6_br[18]_pad  , \h1rdt6_br[19]_pad  , \h1rdt6_br[1]_pad  , \h1rdt6_br[20]_pad  , \h1rdt6_br[21]_pad  , \h1rdt6_br[22]_pad  , \h1rdt6_br[23]_pad  , \h1rdt6_br[24]_pad  , \h1rdt6_br[25]_pad  , \h1rdt6_br[26]_pad  , \h1rdt6_br[27]_pad  , \h1rdt6_br[28]_pad  , \h1rdt6_br[29]_pad  , \h1rdt6_br[2]_pad  , \h1rdt6_br[30]_pad  , \h1rdt6_br[31]_pad  , \h1rdt6_br[3]_pad  , \h1rdt6_br[4]_pad  , \h1rdt6_br[5]_pad  , \h1rdt6_br[6]_pad  , \h1rdt6_br[7]_pad  , \h1rdt6_br[8]_pad  , \h1rdt6_br[9]_pad  , \h1rdt6_dma[0]_pad  , \h1rdt6_dma[10]_pad  , \h1rdt6_dma[11]_pad  , \h1rdt6_dma[12]_pad  , \h1rdt6_dma[13]_pad  , \h1rdt6_dma[14]_pad  , \h1rdt6_dma[15]_pad  , \h1rdt6_dma[16]_pad  , \h1rdt6_dma[17]_pad  , \h1rdt6_dma[18]_pad  , \h1rdt6_dma[19]_pad  , \h1rdt6_dma[1]_pad  , \h1rdt6_dma[20]_pad  , \h1rdt6_dma[21]_pad  , \h1rdt6_dma[22]_pad  , \h1rdt6_dma[23]_pad  , \h1rdt6_dma[24]_pad  , \h1rdt6_dma[25]_pad  , \h1rdt6_dma[26]_pad  , \h1rdt6_dma[27]_pad  , \h1rdt6_dma[28]_pad  , \h1rdt6_dma[29]_pad  , \h1rdt6_dma[2]_pad  , \h1rdt6_dma[30]_pad  , \h1rdt6_dma[31]_pad  , \h1rdt6_dma[3]_pad  , \h1rdt6_dma[4]_pad  , \h1rdt6_dma[5]_pad  , \h1rdt6_dma[6]_pad  , \h1rdt6_dma[7]_pad  , \h1rdt6_dma[8]_pad  , \h1rdt6_dma[9]_pad  , \h1rdt7_br[0]_pad  , \h1rdt7_br[10]_pad  , \h1rdt7_br[11]_pad  , \h1rdt7_br[12]_pad  , \h1rdt7_br[13]_pad  , \h1rdt7_br[14]_pad  , \h1rdt7_br[15]_pad  , \h1rdt7_br[16]_pad  , \h1rdt7_br[17]_pad  , \h1rdt7_br[18]_pad  , \h1rdt7_br[19]_pad  , \h1rdt7_br[1]_pad  , \h1rdt7_br[20]_pad  , \h1rdt7_br[21]_pad  , \h1rdt7_br[22]_pad  , \h1rdt7_br[23]_pad  , \h1rdt7_br[24]_pad  , \h1rdt7_br[25]_pad  , \h1rdt7_br[26]_pad  , \h1rdt7_br[27]_pad  , \h1rdt7_br[28]_pad  , \h1rdt7_br[29]_pad  , \h1rdt7_br[2]_pad  , \h1rdt7_br[30]_pad  , \h1rdt7_br[31]_pad  , \h1rdt7_br[3]_pad  , \h1rdt7_br[4]_pad  , \h1rdt7_br[5]_pad  , \h1rdt7_br[6]_pad  , \h1rdt7_br[7]_pad  , \h1rdt7_br[8]_pad  , \h1rdt7_br[9]_pad  , \h1rdt7_dma[0]_pad  , \h1rdt7_dma[10]_pad  , \h1rdt7_dma[11]_pad  , \h1rdt7_dma[12]_pad  , \h1rdt7_dma[13]_pad  , \h1rdt7_dma[14]_pad  , \h1rdt7_dma[15]_pad  , \h1rdt7_dma[16]_pad  , \h1rdt7_dma[17]_pad  , \h1rdt7_dma[18]_pad  , \h1rdt7_dma[19]_pad  , \h1rdt7_dma[1]_pad  , \h1rdt7_dma[20]_pad  , \h1rdt7_dma[21]_pad  , \h1rdt7_dma[22]_pad  , \h1rdt7_dma[23]_pad  , \h1rdt7_dma[24]_pad  , \h1rdt7_dma[25]_pad  , \h1rdt7_dma[26]_pad  , \h1rdt7_dma[27]_pad  , \h1rdt7_dma[28]_pad  , \h1rdt7_dma[29]_pad  , \h1rdt7_dma[2]_pad  , \h1rdt7_dma[30]_pad  , \h1rdt7_dma[31]_pad  , \h1rdt7_dma[3]_pad  , \h1rdt7_dma[4]_pad  , \h1rdt7_dma[5]_pad  , \h1rdt7_dma[6]_pad  , \h1rdt7_dma[7]_pad  , \h1rdt7_dma[8]_pad  , \h1rdt7_dma[9]_pad  , \h1rdy0_br_pad  , \h1rdy0_dma_pad  , \h1rdy1_br_pad  , \h1rdy1_dma_pad  , \h1rdy2_br_pad  , \h1rdy2_dma_pad  , \h1rdy3_br_pad  , \h1rdy3_dma_pad  , \h1rdy4_br_pad  , \h1rdy4_dma_pad  , \h1rdy5_br_pad  , \h1rdy5_dma_pad  , \h1rdy6_br_pad  , \h1rdy6_dma_pad  , \h1rdy7_br_pad  , \h1rdy7_dma_pad  , \h1rp0_br[0]_pad  , \h1rp0_br[1]_pad  , \h1rp0_dma[0]_pad  , \h1rp0_dma[1]_pad  , \h1rp1_br[0]_pad  , \h1rp1_br[1]_pad  , \h1rp1_dma[0]_pad  , \h1rp1_dma[1]_pad  , \h1rp2_br[0]_pad  , \h1rp2_br[1]_pad  , \h1rp2_dma[0]_pad  , \h1rp2_dma[1]_pad  , \h1rp3_br[0]_pad  , \h1rp3_br[1]_pad  , \h1rp3_dma[0]_pad  , \h1rp3_dma[1]_pad  , \h1rp4_br[0]_pad  , \h1rp4_br[1]_pad  , \h1rp4_dma[0]_pad  , \h1rp4_dma[1]_pad  , \h1rp5_br[0]_pad  , \h1rp5_br[1]_pad  , \h1rp5_dma[0]_pad  , \h1rp5_dma[1]_pad  , \h1rp6_br[0]_pad  , \h1rp6_br[1]_pad  , \h1rp6_dma[0]_pad  , \h1rp6_dma[1]_pad  , \h1rp7_br[0]_pad  , \h1rp7_br[1]_pad  , \h1rp7_dma[0]_pad  , \h1rp7_dma[1]_pad  , \h1size[0]_pad  , \h1size[1]_pad  , \h1size[2]_pad  , \h1write_pad  , \haddr[0]_pad  , \haddr[1]_pad  , \haddr[2]_pad  , \haddr[3]_pad  , \haddr[4]_pad  , \haddr[5]_pad  , \haddr[6]_pad  , \haddr[7]_pad  , \haddr[8]_pad  , \hrdata_reg[0]_pad  , \hrdata_reg[10]_pad  , \hrdata_reg[11]_pad  , \hrdata_reg[12]_pad  , \hrdata_reg[13]_pad  , \hrdata_reg[14]_pad  , \hrdata_reg[15]_pad  , \hrdata_reg[16]_pad  , \hrdata_reg[17]_pad  , \hrdata_reg[18]_pad  , \hrdata_reg[19]_pad  , \hrdata_reg[1]_pad  , \hrdata_reg[20]_pad  , \hrdata_reg[21]_pad  , \hrdata_reg[22]_pad  , \hrdata_reg[23]_pad  , \hrdata_reg[24]_pad  , \hrdata_reg[25]_pad  , \hrdata_reg[26]_pad  , \hrdata_reg[27]_pad  , \hrdata_reg[28]_pad  , \hrdata_reg[29]_pad  , \hrdata_reg[2]_pad  , \hrdata_reg[30]_pad  , \hrdata_reg[31]_pad  , \hrdata_reg[3]_pad  , \hrdata_reg[4]_pad  , \hrdata_reg[5]_pad  , \hrdata_reg[6]_pad  , \hrdata_reg[7]_pad  , \hrdata_reg[8]_pad  , \hrdata_reg[9]_pad  , hreadyin_pad , hreadyout_br_pad , \hresp_br[0]_pad  , \hresp_br[1]_pad  , hsel_br_pad , hsel_reg_pad , \hsize[0]_pad  , \hsize[1]_pad  , \hsize[2]_pad  , \htrans[0]_pad  , \htrans[1]_pad  , \hwdata[0]_pad  , \hwdata[10]_pad  , \hwdata[11]_pad  , \hwdata[12]_pad  , \hwdata[13]_pad  , \hwdata[14]_pad  , \hwdata[15]_pad  , \hwdata[16]_pad  , \hwdata[17]_pad  , \hwdata[18]_pad  , \hwdata[19]_pad  , \hwdata[1]_pad  , \hwdata[20]_pad  , \hwdata[21]_pad  , \hwdata[22]_pad  , \hwdata[23]_pad  , \hwdata[24]_pad  , \hwdata[25]_pad  , \hwdata[26]_pad  , \hwdata[27]_pad  , \hwdata[28]_pad  , \hwdata[29]_pad  , \hwdata[2]_pad  , \hwdata[30]_pad  , \hwdata[31]_pad  , \hwdata[3]_pad  , \hwdata[4]_pad  , \hwdata[5]_pad  , \hwdata[6]_pad  , \hwdata[7]_pad  , \hwdata[8]_pad  , \hwdata[9]_pad  , hwrite_pad , \m1_mux_hrdy_df_reg/NET0131  , \m1_mux_hrmxnof_reg/NET0131  , \m1_mux_hrp_df_reg[0]/NET0131  , \m1_mux_mux_no_reg[0]/NET0131  , \m1_mux_mux_no_reg[1]/NET0131  , \m1_mux_mux_no_reg[2]/NET0131  , \m1_mux_mux_no_reg[3]/NET0131  , \_al_n1  , \g16/_0_  , \g58487/_0_  , \g58489/_0_  , \g58491/_0_  , \g58493/_0_  , \g58495/_0_  , \g58497/_0_  , \g58499/_0_  , \g58500/_0_  , \g58501/_0_  , \g58502/_0_  , \g58504/_0_  , \g58505/_0_  , \g58507/_0_  , \g58508/_0_  , \g58509/_0_  , \g58510/_0_  , \g58556/_0_  , \g58557/_0_  , \g58558/_0_  , \g58559/_0_  , \g58560/_0_  , \g58561/_0_  , \g58562/_0_  , \g58563/_0_  , \g58566/_0_  , \g58567/_0_  , \g58568/_0_  , \g58569/_0_  , \g58570/_0_  , \g58571/_0_  , \g58572/_0_  , \g58573/_0_  , \g58574/_0_  , \g58575/_0_  , \g58576/_0_  , \g58577/_0_  , \g58578/_0_  , \g58579/_0_  , \g58580/_0_  , \g58581/_0_  , \g58584/_0_  , \g58585/_0_  , \g58586/_0_  , \g58587/_0_  , \g58588/_0_  , \g58589/_0_  , \g58590/_0_  , \g58591/_0_  , \g58592/_0_  , \g58593/_0_  , \g58594/_0_  , \g58595/_0_  , \g58596/_0_  , \g58597/_0_  , \g58598/_0_  , \g58599/_0_  , \g58600/_0_  , \g58601/_0_  , \g58602/_0_  , \g58603/_0_  , \g58604/_0_  , \g58605/_0_  , \g58606/_0_  , \g58607/_0_  , \g58608/_0_  , \g58609/_0_  , \g58610/_0_  , \g58611/_0_  , \g58612/_0_  , \g58613/_0_  , \g58614/_0_  , \g58615/_0_  , \g58616/_0_  , \g58617/_0_  , \g58618/_0_  , \g58619/_0_  , \g58620/_0_  , \g58621/_0_  , \g58622/_0_  , \g58623/_0_  , \g58624/_0_  , \g58625/_0_  , \g58626/_0_  , \g58627/_0_  , \g58723/_0_  , \g58734/_0_  , \g58737/_0_  , \g58741/_0_  , \g58749/_0_  , \g58754/_0_  , \g58762/_0_  , \g58763/_0_  , \g58764/_0_  , \g58765/_0_  , \g58766/_0_  , \g58767/_0_  , \g58768/_0_  , \g58769/_0_  , \g58770/_0_  , \g58771/_0_  , \g59788/_0_  , \g59832/_0_  , \g59873/_0_  , \g59874/_0_  , \g59893/_0_  , \g59894/_0_  , \g59895/_0_  , \g59896/_0_  , \g59923/_0_  , \g60031/_0_  , \g60032/_0_  , \g60033/_0_  , \g60036/_0_  , \g60037/_0_  , \g60038/_0_  , \g60165/_0_  , \g60186/_2__syn_2  , \g60187/_0_  , \g60188/_0_  , \g60258/_0_  , \g60259/_0_  , \g60260/_0_  , \g60261/_0_  , \g60263/_0_  , \g60264/_0_  , \g60265/_0_  , \g60266/_0_  , \g60267/_0_  , \g60303/_3_  , \g60360/_0_  , \g60361/_0_  , \g60401/_00_  , \g60428/_0_  , \g60429/_0_  , \g60448/_0_  , \g60449/_0_  , \g60974/_0_  , \g61072/_0_  , \g61073/_0_  , \g61074/_0_  , \g61075/_0_  , \g61076/_0_  , \g61077/_0_  , \g61078/_0_  , \g61079/_0_  , \g61486/_0_  , \g61502/_3_  , \g61879/_0_  , \g62077/_0_  , \g62078/_0_  , \g62079/_0_  , \g62080/_0_  , \g62081/_0_  , \g62082/_0_  , \g62083/_0_  , \g62084/_0_  , \g62085/_0_  , \g62086/_0_  , \g62087/_0_  , \g62088/_0_  , \g62089/_0_  , \g62090/_0_  , \g62091/_0_  , \g62629/_0_  , \g62630/_0_  , \g62631/_0_  , \g62632/_0_  , \g62633/_0_  , \g62634/_0_  , \g62635/_0_  , \g62637/_0_  , \g62638/_0_  , \g62639/_0_  , \g62641/_0_  , \g62643/_0_  , \g62645/_0_  , \g62646/_0_  , \g62647/_0_  , \g62648/_0_  , \g62649/_0_  , \g62650/_0_  , \g62651/_0_  , \g62652/_0_  , \g62655/_0_  , \g62656/_0_  , \g62657/_0_  , \g62658/_0_  , \g62659/_0_  , \g62660/_0_  , \g62661/_0_  , \g62662/_0_  , \g62663/_0_  , \g62664/_0_  , \g62665/_0_  , \g62667/_0_  , \g62668/_0_  , \g62669/_0_  , \g62670/_0_  , \g62671/_0_  , \g62672/_0_  , \g62673/_0_  , \g62674/_0_  , \g62675/_0_  , \g62676/_0_  , \g62677/_0_  , \g62678/_0_  , \g62679/_0_  , \g62680/_0_  , \g62681/_0_  , \g62682/_0_  , \g62683/_0_  , \g62684/_0_  , \g62685/_0_  , \g62686/_0_  , \g62687/_0_  , \g62688/_0_  , \g62689/_0_  , \g62690/_0_  , \g62691/_0_  , \g62692/_0_  , \g62693/_0_  , \g62694/_0_  , \g62695/_0_  , \g62696/_0_  , \g62697/_0_  , \g62698/_0_  , \g62699/_0_  , \g62700/_0_  , \g62701/_0_  , \g62702/_0_  , \g62703/_0_  , \g62704/_0_  , \g62705/_0_  , \g62706/_0_  , \g62707/_0_  , \g62708/_0_  , \g62709/_0_  , \g62710/_0_  , \g62711/_0_  , \g62712/_0_  , \g62713/_0_  , \g62714/_0_  , \g62715/_0_  , \g62716/_0_  , \g62721/_0_  , \g62722/_0_  , \g62723/_0_  , \g62725/_0_  , \g62726/_0_  , \g62727/_0_  , \g62728/_0_  , \g62729/_0_  , \g62730/_0_  , \g62731/_0_  , \g62732/_0_  , \g62733/_0_  , \g62734/_0_  , \g62735/_0_  , \g62736/_0_  , \g62737/_0_  , \g62738/_0_  , \g62739/_0_  , \g62740/_0_  , \g62741/_0_  , \g62742/_0_  , \g62743/_0_  , \g62744/_0_  , \g62745/_0_  , \g62746/_0_  , \g62747/_0_  , \g62748/_0_  , \g62749/_0_  , \g62750/_0_  , \g62751/_0_  , \g62752/_0_  , \g62753/_0_  , \g62754/_0_  , \g62755/_0_  , \g62756/_0_  , \g62757/_0_  , \g62758/_0_  , \g62759/_0_  , \g62760/_0_  , \g62761/_0_  , \g62762/_0_  , \g62763/_0_  , \g62764/_0_  , \g62765/_0_  , \g62766/_0_  , \g62767/_0_  , \g62768/_0_  , \g62769/_0_  , \g62770/_0_  , \g62771/_0_  , \g62772/_0_  , \g62773/_0_  , \g62774/_0_  , \g62775/_0_  , \g62776/_0_  , \g62777/_0_  , \g62778/_0_  , \g62779/_0_  , \g62780/_0_  , \g62781/_0_  , \g62783/_0_  , \g62784/_0_  , \g62785/_0_  , \g62786/_0_  , \g62787/_0_  , \g62788/_0_  , \g62789/_0_  , \g62790/_0_  , \g62791/_0_  , \g62792/_0_  , \g62793/_0_  , \g62794/_0_  , \g62795/_0_  , \g62797/_0_  , \g62798/_0_  , \g62799/_0_  , \g62800/_0_  , \g62801/_0_  , \g62802/_0_  , \g62803/_0_  , \g62804/_0_  , \g62805/_0_  , \g62806/_0_  , \g62807/_0_  , \g62808/_0_  , \g62809/_0_  , \g62810/_0_  , \g62811/_0_  , \g62812/_0_  , \g62813/_0_  , \g62814/_0_  , \g62815/_0_  , \g62816/_0_  , \g62817/_0_  , \g62818/_0_  , \g63108/_0_  , \g63117/_0_  , \g63125/_0_  , \g63126/_0_  , \g63127/_0_  , \g63128/_0_  , \g63129/_0_  , \g63130/_0_  , \g63131/_0_  , \g63132/_0_  , \g63133/_0_  , \g63134/_0_  , \g63135/_0_  , \g63136/_0_  , \g63137/_0_  , \g63138/_0_  , \g63139/_0_  , \g63140/_0_  , \g63141/_0_  , \g63142/_0_  , \g63143/_0_  , \g63144/_0_  , \g63145/_0_  , \g63146/_0_  , \g63147/_0_  , \g63148/_0_  , \g63149/_0_  , \g63150/_0_  , \g63151/_0_  , \g63152/_0_  , \g63153/_0_  , \g63154/_0_  , \g63155/_0_  , \g63156/_0_  , \g63157/_0_  , \g63159/_0_  , \g63160/_0_  , \g63161/_0_  , \g63162/_0_  , \g63163/_0_  , \g63164/_0_  , \g63165/_0_  , \g63166/_0_  , \g63167/_0_  , \g63168/_0_  , \g63169/_0_  , \g63170/_0_  , \g63171/_0_  , \g63172/_0_  , \g63173/_0_  , \g63174/_0_  , \g63175/_0_  , \g63176/_0_  , \g63177/_0_  , \g63178/_0_  , \g63179/_0_  , \g63180/_0_  , \g63181/_0_  , \g63182/_0_  , \g63183/_0_  , \g63184/_0_  , \g63185/_0_  , \g63186/_0_  , \g63187/_0_  , \g63188/_0_  , \g63189/_0_  , \g63190/_0_  , \g63191/_0_  , \g63192/_0_  , \g63193/_0_  , \g63194/_0_  , \g63195/_0_  , \g63196/_0_  , \g63197/_0_  , \g63198/_0_  , \g63199/_0_  , \g63200/_0_  , \g63201/_0_  , \g63202/_0_  , \g63203/_0_  , \g63204/_0_  , \g63205/_0_  , \g63206/_0_  , \g63207/_0_  , \g63208/_0_  , \g63209/_0_  , \g63210/_0_  , \g63211/_0_  , \g63212/_0_  , \g63213/_0_  , \g63214/_0_  , \g63215/_0_  , \g63216/_0_  , \g63217/_0_  , \g63218/_0_  , \g63219/_0_  , \g63220/_0_  , \g63221/_0_  , \g63222/_0_  , \g63223/_0_  , \g63224/_0_  , \g63225/_0_  , \g63226/_0_  , \g63228/_0_  , \g63229/_0_  , \g63231/_0_  , \g63232/_0_  , \g63233/_0_  , \g63234/_0_  , \g63235/_0_  , \g63236/_0_  , \g63237/_0_  , \g63238/_0_  , \g63239/_0_  , \g63240/_0_  , \g63241/_0_  , \g63242/_0_  , \g63244/_0_  , \g63246/_0_  , \g63247/_0_  , \g63248/_0_  , \g63249/_0_  , \g63250/_0_  , \g63251/_0_  , \g63252/_0_  , \g63253/_0_  , \g63254/_0_  , \g63255/_0_  , \g63256/_0_  , \g63257/_0_  , \g63258/_0_  , \g63259/_0_  , \g63260/_0_  , \g63261/_0_  , \g63262/_0_  , \g63263/_0_  , \g63264/_0_  , \g63265/_0_  , \g63266/_0_  , \g63267/_0_  , \g63268/_0_  , \g63269/_0_  , \g63270/_0_  , \g63272/_0_  , \g63291/_0_  , \g63292/_0_  , \g63293/_0_  , \g63294/_0_  , \g63295/_0_  , \g63298/_0_  , \g63299/_0_  , \g63300/_0_  , \g63301/_0_  , \g63302/_0_  , \g63303/_0_  , \g63304/_0_  , \g63305/_0_  , \g63306/_0_  , \g63307/_0_  , \g63308/_0_  , \g63309/_0_  , \g63310/_0_  , \g63311/_0_  , \g63312/_0_  , \g63313/_0_  , \g63314/_0_  , \g63315/_0_  , \g63316/_0_  , \g63317/_0_  , \g63318/_0_  , \g63320/_0_  , \g63322/_0_  , \g63323/_0_  , \g63324/_0_  , \g63325/_0_  , \g63326/_0_  , \g63327/_0_  , \g63328/_0_  , \g63329/_0_  , \g63330/_0_  , \g63331/_0_  , \g63332/_0_  , \g63333/_0_  , \g63334/_0_  , \g63335/_0_  , \g63336/_0_  , \g63337/_0_  , \g63338/_0_  , \g63339/_0_  , \g63340/_0_  , \g63341/_0_  , \g63342/_0_  , \g63343/_0_  , \g63344/_0_  , \g63345/_0_  , \g63346/_0_  , \g63347/_0_  , \g63348/_0_  , \g63349/_0_  , \g63350/_0_  , \g63351/_0_  , \g63352/_0_  , \g63353/_0_  , \g63354/_0_  , \g63355/_0_  , \g63356/_0_  , \g63357/_0_  , \g63358/_0_  , \g63359/_0_  , \g63360/_0_  , \g63361/_0_  , \g63362/_0_  , \g63363/_0_  , \g63364/_0_  , \g63365/_0_  , \g63366/_0_  , \g63367/_0_  , \g63368/_0_  , \g63369/_0_  , \g63370/_0_  , \g63371/_0_  , \g63372/_0_  , \g63373/_0_  , \g63374/_0_  , \g63375/_0_  , \g63376/_0_  , \g63377/_0_  , \g63378/_0_  , \g63379/_0_  , \g63380/_0_  , \g63383/_3_  , \g63386/_0_  , \g63387/_0_  , \g63388/_0_  , \g63389/_0_  , \g63390/_0_  , \g63391/_0_  , \g63392/_0_  , \g63419/_0_  , \g63421/_0_  , \g63422/_0_  , \g63423/_0_  , \g63424/_0_  , \g63425/_0_  , \g63536/_3_  , \g63625/_0_  , \g63628/_0_  , \g63871/_0_  , \g63874/_0_  , \g63889/_0_  , \g63933/_0_  , \g63945/_0_  , \g63959/_0_  , \g63962/_0_  , \g63974/_0_  , \g63977/_0_  , \g64035/_0_  , \g64435/_3_  , \g64939/_0_  , \g65149/_0_  , \g65632/_3_  , \g65633/_0_  , \g65634/_0_  , \g65635/_0_  , \g65636/_0_  , \g65638/_3_  , \g65640/_3_  , \g65999/_0_  , \g66912/_0_  , \g66914/_0_  , \g67555/_3_  , \g67564/_3_  , \g67567/_3_  , \g67735/_0_  , \g67736/_0_  , \g67737/_0_  , \g67738/_0_  , \g67758/_0_  , \g67760/_0_  , \g67761/_0_  , \g67763/_0_  , \g67766/_0_  , \g67810/_0_  , \g67816/_0_  , \g67902/_0_  , \g67927/_0_  , \g67936/_0_  , \g68067/_0_  , \g68068/_0_  , \g68069/_0_  , \g68070/_0_  , \g68071/_0_  , \g68072/_0_  , \g68073/_0_  , \g68074/_0_  , \g68075/_0_  , \g68076/_0_  , \g68077/_0_  , \g68078/_0_  , \g68079/_0_  , \g68080/_0_  , \g68081/_0_  , \g68082/_0_  , \g68083/_0_  , \g68084/_0_  , \g68085/_0_  , \g68086/_0_  , \g68087/_0_  , \g68088/_0_  , \g68089/_0_  , \g68090/_0_  , \g68091/_0_  , \g68096/_0_  , \g68160/_0_  , \g68218/_0_  , \g68219/_0_  , \g68220/_0_  , \g68221/_0_  , \g68222/_0_  , \g68226/_0_  , \g68247/_0_  , \g68252/_0_  , \g68632/_0_  , \g68633/_0_  , \g68635/_0_  , \g68640/_0_  , \g68642/_0_  , \g68643/_0_  , \g68644/_0_  , \g68645/_0_  , \g68649/_0_  , \g68668/_2_  , \g68670/_0_  , \g68681/_3_  , \g68689/_0_  , \g68690/_0_  , \g68691/_0_  , \g68692/_0_  , \g68693/_0_  , \g68694/_0_  , \g68695/_0_  , \g68737/_0_  , \g68742/_0_  , \g68745/_0_  , \g68750/_0_  , \g68759/_0_  , \g68761/_0_  , \g68774/_0_  , \g68775/_0_  , \g68776/_0_  , \g68777/_0_  , \g68778/_0_  , \g68780/_0_  , \g68781/_0_  , \g68782/_0_  , \g68783/_0_  , \g68784/_0_  , \g68785/_0_  , \g68786/_0_  , \g68787/_0_  , \g68790/_0_  , \g68791/_0_  , \g68793/_0_  , \g68794/_0_  , \g68795/_0_  , \g68796/_0_  , \g68797/_0_  , \g68804/_0_  , \g68805/_0_  , \g68807/_0_  , \g68809/_0_  , \g68864/_3_  , \g68865/_3_  , \g68866/_3_  , \g68867/_3_  , \g68868/_3_  , \g68869/_3_  , \g68870/_3_  , \g68871/_3_  , \g68872/_3_  , \g68873/_3_  , \g68874/_3_  , \g68875/_3_  , \g68876/_3_  , \g68877/_3_  , \g68878/_3_  , \g68879/_3_  , \g68880/_3_  , \g68881/_3_  , \g68882/_3_  , \g68883/_3_  , \g68884/_3_  , \g68885/_3_  , \g68886/_3_  , \g68887/_3_  , \g68888/_3_  , \g68889/_3_  , \g68890/_3_  , \g68891/_3_  , \g68892/_3_  , \g68893/_3_  , \g68894/_3_  , \g68895/_3_  , \g69037/_1__syn_2  , \g69077/_0_  , \g69081/_0_  , \g69084/_0_  , \g69085/_0_  , \g69086/_0_  , \g69088/_0_  , \g69094/_0_  , \g69095/_0_  , \g69097/_0_  , \g69114/_3_  , \g69116/_3_  , \g69118/_3_  , \g69120/_3_  , \g69122/_3_  , \g69124/_3_  , \g69126/_3_  , \g69128/_3_  , \g69581/_3_  , \g70303/_1__syn_2  , \g70304/_1__syn_2  , \g70305/_1__syn_2  , \g70306/_1__syn_2  , \g70353/_1__syn_2  , \g70359/_2_  , \g70364/_1__syn_2  , \g70375/_1__syn_2  , \g70380/_2_  , \g70383/_1__syn_2  , \g70394/_2_  , \g70395/_2_  , \g70396/_1__syn_2  , \g70398/_1__syn_2  , \g70407/_1_  , \g70416/_1__syn_2  , \g70418/_1__syn_2  , \g70419/_2_  , \g70424/_1_  , \g70465/_2_  , \g70511/_1_  , \g70512/_1_  , \g70513/_2_  , \g70514/_2_  , \g70516/_2_  , \g70518/_2_  , \g70519/_2_  , \g70520/_2_  , \g70530/_2_  , \g70534/_3_  , \g70536/_3_  , \g70540/_3_  , \g70541/_2_  , \g70545/_3_  , \g70546/_2_  , \g70547/_2_  , \g70550/_3_  , \g70551/_2_  , \g70552/_2_  , \g70558/_3_  , \g70559/_2_  , \g70560/_2_  , \g70562/_3_  , \g70564/_3_  , \g70567/_3_  , \g70568/_2_  , \g70571/_3_  , \g70577/_0_  , \g70578/_2_  , \g70585/_3_  , \g70586/_2_  , \g70587/_2_  , \g70588/_3_  , \g70602/_3_  , \g70841/_0_  , \g70842/_0_  , \g70843/_0_  , \g70844/_0_  , \g70845/_0_  , \g70846/_0_  , \g70847/_0_  , \g70848/_0_  , \g70849/_0_  , \g70850/_0_  , \g70851/_0_  , \g70852/_0_  , \g70853/_0_  , \g70854/_0_  , \g70855/_0_  , \g70856/_0_  , \g70857/_0_  , \g70858/_0_  , \g70859/_0_  , \g70860/_0_  , \g70861/_0_  , \g70862/_0_  , \g70863/_0_  , \g70864/_0_  , \g70865/_0_  , \g70866/_0_  , \g70867/_0_  , \g70868/_0_  , \g70869/_0_  , \g70870/_0_  , \g70871/_0_  , \g70872/_0_  , \g70944/_1__syn_2  , \g71042/_1__syn_2  , \g71064/_1__syn_2  , \g71065/_1__syn_2  , \g71076/_1__syn_2  , \g71077/_1__syn_2  , \g71202/_1__syn_2  , \g71204/_1__syn_2  , \g71236/_0_  , \g71237/_0_  , \g71241/_0_  , \g71242/_0_  , \g71245/_0_  , \g71246/_0_  , \g71306/_0_  , \g71308/_0_  , \g71309/_0_  , \g71310/_0_  , \g71355/_0_  , \g71416/_0_  , \g71417/_0_  , \g71420/_0_  , \g71432/_0_  , \g71434/_0_  , \g71435/_0_  , \g71436/_0_  , \g71446/_0_  , \g71449/_0_  , \g71451/_0_  , \g71452/_0_  , \g71485/_0_  , \g71494/_0_  , \g71499/_0_  , \g71500/_0_  , \g71501/_0_  , \g71502/_0_  , \g71503/_0_  , \g71504/_0_  , \g71505/_0_  , \g71506/_0_  , \g71815/_0_  , \g71823/_0_  , \g71832/_0_  , \g71833/_0__syn_2  , \g71837/_0_  , \g71838/_0_  , \g71846/_1__syn_2  , \g71847/_1__syn_2  , \g71849/_0_  , \g71854/_0_  , \g71858/_1__syn_2  , \g71859/_1__syn_2  , \g71863/_0_  , \g71867/_0_  , \g71869/_0_  , \g71872/_1_  , \g71873/_1__syn_2  , \g71874/_1__syn_2  , \g71875/_0_  , \g71877/_1__syn_2  , \g71881/_0_  , \g71906/_0_  , \g71907/_1__syn_2  , \g71910/_0_  , \g71911/_0_  , \g71912/_1__syn_2  , \g71913/_1__syn_2  , \g71914/_1__syn_2  , \g71918/_0_  , \g71921/_0_  , \g71922/_0_  , \g71929/_1__syn_2  , \g71931/_1__syn_2  , \g71938/_1__syn_2  , \g71942/_0_  , \g71946/_1__syn_2  , \g71947/_0_  , \g71951/_0_  , \g71958/_1__syn_2  , \g71965/_0_  , \g71970/_1__syn_2  , \g71972/_1__syn_2  , \g71973/_1__syn_2  , \g71986/_1__syn_2  , \g71987/_1__syn_2  , \g71990/_1__syn_2  , \g71991/_1__syn_2  , \g71992/_1__syn_2  , \g71994/_1__syn_2  , \g71997/_1__syn_2  , \g72001/_1__syn_2  , \g72013/_1__syn_2  , \g72021/_1__syn_2  , \g72030/_0_  , \g72031/_0__syn_2  , \g72036/_1__syn_2  , \g72038/_0_  , \g72042/_1__syn_2  , \g72047/_1__syn_2  , \g72048/_1__syn_2  , \g72049/_1__syn_2  , \g72056/_0_  , \g72064/_1__syn_2  , \g72073/_1__syn_2  , \g72075/_0_  , \g72078/_0_  , \g72081/_0_  , \g72091/_0_  , \g72096/_0_  , \g72100/_1__syn_2  , \g72113/_0_  , \g72118/_0_  , \g72121/_1__syn_2  , \g72122/_1__syn_2  , \g72125/_1__syn_2  , \g72128/_0_  , \g72140/_0_  , \g72144/_1__syn_2  , \g72154/_1__syn_2  , \g72159/_0_  , \g72164/_1__syn_2  , \g72165/_1__syn_2  , \g72167/_1__syn_2  , \g72170/_1__syn_2  , \g72172/_1__syn_2  , \g72173/_0_  , \g72177/_1__syn_2  , \g72189/_0_  , \g72194/_0_  , \g72196/_0_  , \g72198/_0_  , \g72206/_1__syn_2  , \g72209/_1__syn_2  , \g72210/_1__syn_2  , \g72211/_0_  , \g72215/_0_  , \g72227/_1__syn_2  , \g72229/_1__syn_2  , \g72230/_0_  , \g72239/_0_  , \g72250/_3_  , \g72251/_3_  , \g72252/_3_  , \g72253/_3_  , \g72254/_3_  , \g72255/_3_  , \g72256/_3_  , \g72257/_3_  , \g72259/_3_  , \g72260/_3_  , \g72261/_3_  , \g72262/_3_  , \g72263/_3_  , \g72264/_3_  , \g72265/_3_  , \g72266/_3_  , \g72267/_3_  , \g72273/_3_  , \g72275/_3_  , \g72282/_3_  , \g72285/_3_  , \g72293/_3_  , \g72304/_3_  , \g72305/_3_  , \g72306/_3_  , \g72307/_3_  , \g72309/_3_  , \g72310/_3_  , \g72324/_3_  , \g72325/_3_  , \g72326/_3_  , \g72327/_3_  , \g72711/_0_  , \g72763/_0_  , \g72966/_0_  , \g72967/_0_  , \g73018/_0_  , \g73058/_0_  , \g73062/_0_  , \g73067/_0_  , \g73068/_0_  , \g73207/_0_  , \g75007/_1__syn_2  , \g75568/_1_  , \g75792/_0_  , \g75836/_0_  , \g76027/_0_  , \g76034/_0_  , \g76108/_0_  , \g76130/_0_  , \g76266/_0_  , \g76315/_0_  , \g76569/_0_  , \g76714/_0_  , \g77122/_1__syn_2  , \g77709/_1_  , \g81909/_0_  , \g81922/_0_  , \g81926/_1__syn_2  , \g82197/_1_  , \g82272/_0_  , \g82291/_0_  , \g82716/_0_  , \g82718/_0_  , \g82738/_0_  , \g82769/_0_  , \g82775/_0_  , \g82779/_1__syn_2  , \g82804/_0_  , \g82810/_0_  , \g82817/_0_  , \g82823/_0_  , \g82835/_0_  , \g82841/_0_  , \g82847/_0_  , \g82853/_0_  , \g82859/_0_  , \g82862/_1__syn_2  , \g82956/_0_  , \g82959/_1_  , \g83020/_0_  , \g83025/_0_  , \g83078/_0_  , \g83083/_0_  , \g83121/_0_  , \g83135/_0_  , \g83205/_0_  , \g83240/_0_  , \g83509/_1__syn_2  , \g83769/_0_  , \h0lock_pad  , \h1sel_br[7]_pad  , \h1sel_dma[0]_pad  , \h1sel_dma[4]_pad  , \h1sel_dma[7]_pad  );
  input \ahb_mst0_hsizeo_reg[0]/NET0131  ;
  input \ahb_mst0_hsizeo_reg[1]/NET0131  ;
  input \ahb_mst0_hsizeo_reg[2]/NET0131  ;
  input \ahb_mst0_m0_m1_diff_tx_reg/NET0131  ;
  input \ahb_mst0_mx_cmd_st_reg[0]/NET0131  ;
  input \ahb_mst0_mx_cmd_st_reg[1]/NET0131  ;
  input \ahb_mst0_mx_dtp_reg/NET0131  ;
  input \ahb_mst1_mx_cmd_st_reg[0]/NET0131  ;
  input \ahb_mst1_mx_cmd_st_reg[1]/NET0131  ;
  input \ahb_mst1_mx_dtp_reg/NET0131  ;
  input \ahb_slv_br_st_reg[0]/NET0131  ;
  input \ahb_slv_br_st_reg[1]/NET0131  ;
  input \ahb_slv_br_st_reg[2]/NET0131  ;
  input \ahb_slv_slv_ad_d1o_reg[2]/NET0131  ;
  input \ahb_slv_slv_ad_d1o_reg[3]/NET0131  ;
  input \ahb_slv_slv_ad_d1o_reg[4]/NET0131  ;
  input \ahb_slv_slv_ad_d1o_reg[5]/NET0131  ;
  input \ahb_slv_slv_ad_d1o_reg[6]/NET0131  ;
  input \ahb_slv_slv_ad_d1o_reg[7]/NET0131  ;
  input \ahb_slv_slv_ad_d1o_reg[8]/NET0131  ;
  input \ahb_slv_slv_br_req_reg/NET0131  ;
  input \ahb_slv_slv_pt_d1o_reg[0]/NET0131  ;
  input \ahb_slv_slv_pt_d1o_reg[1]/NET0131  ;
  input \ahb_slv_slv_pt_d1o_reg[2]/NET0131  ;
  input \ahb_slv_slv_pt_d1o_reg[3]/NET0131  ;
  input \ahb_slv_slv_sz_d1o_reg[0]/NET0131  ;
  input \ahb_slv_slv_sz_d1o_reg[1]/NET0131  ;
  input \ahb_slv_slv_sz_d1o_reg[2]/NET0131  ;
  input \ahb_slv_slv_wr_d1o_reg/NET0131  ;
  input \ch_sel_arb_ch_sel_reg[0]/P0000_reg_syn_2  ;
  input \ch_sel_arb_ch_sel_reg[1]/P0000_reg_syn_2  ;
  input \ch_sel_arb_ch_sel_reg[2]/P0000_reg_syn_2  ;
  input \ch_sel_arb_chcsr_reg_reg[10]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[11]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[12]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[13]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[15]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[16]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[17]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[18]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[19]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[1]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[20]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[2]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[3]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[4]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[5]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[6]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[8]/NET0131  ;
  input \ch_sel_arb_chcsr_reg_reg[9]/NET0131  ;
  input \ch_sel_arb_req_reg/NET0131  ;
  input \ch_sel_de_stup_d1_reg/NET0131  ;
  input \ch_sel_dma_reqd1_reg[0]/NET0131  ;
  input \ch_sel_dma_reqd1_reg[1]/NET0131  ;
  input \ch_sel_dma_reqd1_reg[2]/NET0131  ;
  input \ch_sel_dma_reqd1_reg[3]/NET0131  ;
  input \ch_sel_dma_reqd1_reg[4]/NET0131  ;
  input \ch_sel_dma_reqd1_reg[5]/NET0131  ;
  input \ch_sel_dma_reqd1_reg[6]/NET0131  ;
  input \ch_sel_dma_reqd1_reg[7]/NET0131  ;
  input \ch_sel_dma_reqd2_reg[0]/NET0131  ;
  input \ch_sel_dma_reqd2_reg[1]/P0001  ;
  input \ch_sel_dma_reqd2_reg[2]/P0001  ;
  input \ch_sel_dma_reqd2_reg[3]/P0001  ;
  input \ch_sel_dma_reqd2_reg[4]/NET0131  ;
  input \ch_sel_dma_reqd2_reg[5]/NET0131  ;
  input \ch_sel_dma_reqd2_reg[6]/NET0131  ;
  input \ch_sel_dma_reqd2_reg[7]/NET0131  ;
  input \ch_sel_dma_rrarb0_state_reg[0]/NET0131  ;
  input \ch_sel_dma_rrarb0_state_reg[1]/NET0131  ;
  input \ch_sel_dma_rrarb0_state_reg[2]/NET0131  ;
  input \ch_sel_dma_rrarb1_state_reg[0]/NET0131  ;
  input \ch_sel_dma_rrarb1_state_reg[1]/NET0131  ;
  input \ch_sel_dma_rrarb1_state_reg[2]/NET0131  ;
  input \ch_sel_dma_rrarb2_state_reg[0]/NET0131  ;
  input \ch_sel_dma_rrarb2_state_reg[1]/NET0131  ;
  input \ch_sel_dma_rrarb2_state_reg[2]/NET0131  ;
  input \ch_sel_dma_rrarb3_state_reg[0]/NET0131  ;
  input \ch_sel_dma_rrarb3_state_reg[1]/NET0131  ;
  input \ch_sel_dma_rrarb3_state_reg[2]/NET0131  ;
  input \ch_sel_fix_pri_sel_reg[0]/NET0131  ;
  input \ch_sel_fix_pri_sel_reg[1]/NET0131  ;
  input \ch_sel_vld_req_any_d1_reg/NET0131  ;
  input \ctl_rf_abt_reg[0]/NET0131  ;
  input \ctl_rf_abt_reg[1]/NET0131  ;
  input \ctl_rf_abt_reg[2]/NET0131  ;
  input \ctl_rf_abt_reg[3]/NET0131  ;
  input \ctl_rf_abt_reg[4]/NET0131  ;
  input \ctl_rf_abt_reg[5]/NET0131  ;
  input \ctl_rf_abt_reg[6]/NET0131  ;
  input \ctl_rf_abt_reg[7]/NET0131  ;
  input \ctl_rf_be_d1_reg[0]/P0001  ;
  input \ctl_rf_be_d1_reg[1]/P0001  ;
  input \ctl_rf_be_d1_reg[2]/P0001  ;
  input \ctl_rf_be_d1_reg[3]/P0001  ;
  input \ctl_rf_c0_rf_autold_reg/NET0131  ;
  input \ctl_rf_c0_rf_ch_en_reg/NET0131  ;
  input \ctl_rf_c0_rf_chabt_reg/NET0131  ;
  input \ctl_rf_c0_rf_chdad_reg[0]/NET0131  ;
  input \ctl_rf_c0_rf_chdad_reg[10]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[11]/NET0131  ;
  input \ctl_rf_c0_rf_chdad_reg[12]/NET0131  ;
  input \ctl_rf_c0_rf_chdad_reg[13]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[14]/NET0131  ;
  input \ctl_rf_c0_rf_chdad_reg[15]/NET0131  ;
  input \ctl_rf_c0_rf_chdad_reg[16]/NET0131  ;
  input \ctl_rf_c0_rf_chdad_reg[17]/NET0131  ;
  input \ctl_rf_c0_rf_chdad_reg[18]/NET0131  ;
  input \ctl_rf_c0_rf_chdad_reg[19]/NET0131  ;
  input \ctl_rf_c0_rf_chdad_reg[1]/NET0131  ;
  input \ctl_rf_c0_rf_chdad_reg[20]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[21]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[22]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[23]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[24]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[25]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[26]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[27]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[28]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[29]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[2]/NET0131  ;
  input \ctl_rf_c0_rf_chdad_reg[30]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[31]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[3]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[4]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[5]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[6]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[7]/P0002  ;
  input \ctl_rf_c0_rf_chdad_reg[8]/NET0131  ;
  input \ctl_rf_c0_rf_chdad_reg[9]/P0002  ;
  input \ctl_rf_c0_rf_chllp_cnt_reg[0]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_cnt_reg[1]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_cnt_reg[2]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_cnt_reg[3]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_on_reg/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[0]/P0002  ;
  input \ctl_rf_c0_rf_chllp_reg[10]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[11]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[12]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[13]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[14]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[15]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[16]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[17]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[18]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[19]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[1]/P0002  ;
  input \ctl_rf_c0_rf_chllp_reg[20]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[21]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[22]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[23]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[24]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[25]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[26]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[27]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[28]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[29]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[2]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[30]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[31]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[3]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[4]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[5]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[6]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[7]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[8]/NET0131  ;
  input \ctl_rf_c0_rf_chllp_reg[9]/NET0131  ;
  input \ctl_rf_c0_rf_chllpen_reg/NET0131  ;
  input \ctl_rf_c0_rf_chpri_reg[0]/NET0131  ;
  input \ctl_rf_c0_rf_chpri_reg[1]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[0]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[10]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[11]/P0002  ;
  input \ctl_rf_c0_rf_chsad_reg[12]/P0002  ;
  input \ctl_rf_c0_rf_chsad_reg[13]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[14]/P0002  ;
  input \ctl_rf_c0_rf_chsad_reg[15]/P0002  ;
  input \ctl_rf_c0_rf_chsad_reg[16]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[17]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[18]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[19]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[1]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[20]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[21]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[22]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[23]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[24]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[25]/P0002  ;
  input \ctl_rf_c0_rf_chsad_reg[26]/P0002  ;
  input \ctl_rf_c0_rf_chsad_reg[27]/P0002  ;
  input \ctl_rf_c0_rf_chsad_reg[28]/P0002  ;
  input \ctl_rf_c0_rf_chsad_reg[29]/P0002  ;
  input \ctl_rf_c0_rf_chsad_reg[2]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[30]/P0002  ;
  input \ctl_rf_c0_rf_chsad_reg[31]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[3]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[4]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[5]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[6]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[7]/NET0131  ;
  input \ctl_rf_c0_rf_chsad_reg[8]/P0002  ;
  input \ctl_rf_c0_rf_chsad_reg[9]/NET0131  ;
  input \ctl_rf_c0_rf_chtsz_reg[0]/P0002  ;
  input \ctl_rf_c0_rf_chtsz_reg[10]/P0002  ;
  input \ctl_rf_c0_rf_chtsz_reg[11]/P0002  ;
  input \ctl_rf_c0_rf_chtsz_reg[1]/P0002  ;
  input \ctl_rf_c0_rf_chtsz_reg[2]/P0002  ;
  input \ctl_rf_c0_rf_chtsz_reg[3]/P0002  ;
  input \ctl_rf_c0_rf_chtsz_reg[4]/NET0131  ;
  input \ctl_rf_c0_rf_chtsz_reg[5]/NET0131  ;
  input \ctl_rf_c0_rf_chtsz_reg[6]/NET0131  ;
  input \ctl_rf_c0_rf_chtsz_reg[7]/NET0131  ;
  input \ctl_rf_c0_rf_chtsz_reg[8]/P0002  ;
  input \ctl_rf_c0_rf_chtsz_reg[9]/P0002  ;
  input \ctl_rf_c0_rf_dad_ctl0_reg/NET0131  ;
  input \ctl_rf_c0_rf_dad_ctl1_reg/NET0131  ;
  input \ctl_rf_c0_rf_dreqmode_reg/NET0131  ;
  input \ctl_rf_c0_rf_dst_sel_reg/NET0131  ;
  input \ctl_rf_c0_rf_dwidth_reg[0]/NET0131  ;
  input \ctl_rf_c0_rf_dwidth_reg[1]/NET0131  ;
  input \ctl_rf_c0_rf_dwidth_reg[2]/NET0131  ;
  input \ctl_rf_c0_rf_int_abt_msk_reg/NET0131  ;
  input \ctl_rf_c0_rf_int_err_msk_reg/NET0131  ;
  input \ctl_rf_c0_rf_int_tc1_msk_reg/NET0131  ;
  input \ctl_rf_c0_rf_int_tc_msk_reg/NET0131  ;
  input \ctl_rf_c0_rf_mode_reg/NET0131  ;
  input \ctl_rf_c0_rf_prot1_reg/NET0131  ;
  input \ctl_rf_c0_rf_prot2_reg/NET0131  ;
  input \ctl_rf_c0_rf_prot3_reg/NET0131  ;
  input \ctl_rf_c0_rf_sad_ctl0_reg/NET0131  ;
  input \ctl_rf_c0_rf_sad_ctl1_reg/NET0131  ;
  input \ctl_rf_c0_rf_src_sel_reg/NET0131  ;
  input \ctl_rf_c0_rf_src_sz_reg[0]/NET0131  ;
  input \ctl_rf_c0_rf_src_sz_reg[1]/NET0131  ;
  input \ctl_rf_c0_rf_src_sz_reg[2]/NET0131  ;
  input \ctl_rf_c0_rf_swidth_reg[0]/NET0131  ;
  input \ctl_rf_c0_rf_swidth_reg[1]/NET0131  ;
  input \ctl_rf_c0_rf_swidth_reg[2]/NET0131  ;
  input \ctl_rf_c0brbs_reg[16]/NET0131  ;
  input \ctl_rf_c0brbs_reg[17]/NET0131  ;
  input \ctl_rf_c0brbs_reg[18]/NET0131  ;
  input \ctl_rf_c0brbs_reg[19]/NET0131  ;
  input \ctl_rf_c0brbs_reg[20]/NET0131  ;
  input \ctl_rf_c0brbs_reg[21]/NET0131  ;
  input \ctl_rf_c0brbs_reg[22]/NET0131  ;
  input \ctl_rf_c0brbs_reg[23]/NET0131  ;
  input \ctl_rf_c0brbs_reg[24]/NET0131  ;
  input \ctl_rf_c0brbs_reg[25]/NET0131  ;
  input \ctl_rf_c0brbs_reg[26]/NET0131  ;
  input \ctl_rf_c0brbs_reg[27]/NET0131  ;
  input \ctl_rf_c0brbs_reg[28]/NET0131  ;
  input \ctl_rf_c0brbs_reg[29]/NET0131  ;
  input \ctl_rf_c0brbs_reg[30]/NET0131  ;
  input \ctl_rf_c0brbs_reg[31]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[16]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[17]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[18]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[19]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[20]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[21]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[22]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[23]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[24]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[25]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[26]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[27]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[28]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[29]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[30]/NET0131  ;
  input \ctl_rf_c0dmabs_reg[31]/NET0131  ;
  input \ctl_rf_c1_rf_autold_reg/NET0131  ;
  input \ctl_rf_c1_rf_ch_en_reg/NET0131  ;
  input \ctl_rf_c1_rf_chabt_reg/NET0131  ;
  input \ctl_rf_c1_rf_chdad_reg[0]/NET0131  ;
  input \ctl_rf_c1_rf_chdad_reg[10]/NET0131  ;
  input \ctl_rf_c1_rf_chdad_reg[11]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[12]/NET0131  ;
  input \ctl_rf_c1_rf_chdad_reg[13]/NET0131  ;
  input \ctl_rf_c1_rf_chdad_reg[14]/NET0131  ;
  input \ctl_rf_c1_rf_chdad_reg[15]/NET0131  ;
  input \ctl_rf_c1_rf_chdad_reg[16]/NET0131  ;
  input \ctl_rf_c1_rf_chdad_reg[17]/NET0131  ;
  input \ctl_rf_c1_rf_chdad_reg[18]/NET0131  ;
  input \ctl_rf_c1_rf_chdad_reg[19]/NET0131  ;
  input \ctl_rf_c1_rf_chdad_reg[1]/NET0131  ;
  input \ctl_rf_c1_rf_chdad_reg[20]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[21]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[22]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[23]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[24]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[25]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[26]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[27]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[28]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[29]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[2]/NET0131  ;
  input \ctl_rf_c1_rf_chdad_reg[30]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[31]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[3]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[4]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[5]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[6]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[7]/P0002  ;
  input \ctl_rf_c1_rf_chdad_reg[8]/NET0131  ;
  input \ctl_rf_c1_rf_chdad_reg[9]/P0002  ;
  input \ctl_rf_c1_rf_chllp_cnt_reg[0]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_cnt_reg[1]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_cnt_reg[2]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_cnt_reg[3]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_on_reg/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[0]/P0002  ;
  input \ctl_rf_c1_rf_chllp_reg[10]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[11]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[12]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[13]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[14]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[15]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[16]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[17]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[18]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[19]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[1]/P0002  ;
  input \ctl_rf_c1_rf_chllp_reg[20]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[21]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[22]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[23]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[24]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[25]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[26]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[27]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[28]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[29]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[2]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[30]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[31]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[3]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[4]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[5]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[6]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[7]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[8]/NET0131  ;
  input \ctl_rf_c1_rf_chllp_reg[9]/NET0131  ;
  input \ctl_rf_c1_rf_chllpen_reg/NET0131  ;
  input \ctl_rf_c1_rf_chpri_reg[0]/NET0131  ;
  input \ctl_rf_c1_rf_chpri_reg[1]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[0]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[10]/P0002  ;
  input \ctl_rf_c1_rf_chsad_reg[11]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[12]/P0002  ;
  input \ctl_rf_c1_rf_chsad_reg[13]/P0002  ;
  input \ctl_rf_c1_rf_chsad_reg[14]/P0002  ;
  input \ctl_rf_c1_rf_chsad_reg[15]/P0002  ;
  input \ctl_rf_c1_rf_chsad_reg[16]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[17]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[18]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[19]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[1]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[20]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[21]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[22]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[23]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[24]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[25]/P0002  ;
  input \ctl_rf_c1_rf_chsad_reg[26]/P0002  ;
  input \ctl_rf_c1_rf_chsad_reg[27]/P0002  ;
  input \ctl_rf_c1_rf_chsad_reg[28]/P0002  ;
  input \ctl_rf_c1_rf_chsad_reg[29]/P0002  ;
  input \ctl_rf_c1_rf_chsad_reg[2]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[30]/P0002  ;
  input \ctl_rf_c1_rf_chsad_reg[31]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[3]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[4]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[5]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[6]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[7]/NET0131  ;
  input \ctl_rf_c1_rf_chsad_reg[8]/P0002  ;
  input \ctl_rf_c1_rf_chsad_reg[9]/NET0131  ;
  input \ctl_rf_c1_rf_chtsz_reg[0]/P0002  ;
  input \ctl_rf_c1_rf_chtsz_reg[10]/P0002  ;
  input \ctl_rf_c1_rf_chtsz_reg[11]/P0002  ;
  input \ctl_rf_c1_rf_chtsz_reg[1]/P0002  ;
  input \ctl_rf_c1_rf_chtsz_reg[2]/P0002  ;
  input \ctl_rf_c1_rf_chtsz_reg[3]/P0002  ;
  input \ctl_rf_c1_rf_chtsz_reg[4]/NET0131  ;
  input \ctl_rf_c1_rf_chtsz_reg[5]/NET0131  ;
  input \ctl_rf_c1_rf_chtsz_reg[6]/NET0131  ;
  input \ctl_rf_c1_rf_chtsz_reg[7]/NET0131  ;
  input \ctl_rf_c1_rf_chtsz_reg[8]/P0002  ;
  input \ctl_rf_c1_rf_chtsz_reg[9]/P0002  ;
  input \ctl_rf_c1_rf_dad_ctl0_reg/NET0131  ;
  input \ctl_rf_c1_rf_dad_ctl1_reg/NET0131  ;
  input \ctl_rf_c1_rf_dreqmode_reg/NET0131  ;
  input \ctl_rf_c1_rf_dst_sel_reg/NET0131  ;
  input \ctl_rf_c1_rf_dwidth_reg[0]/NET0131  ;
  input \ctl_rf_c1_rf_dwidth_reg[1]/NET0131  ;
  input \ctl_rf_c1_rf_dwidth_reg[2]/NET0131  ;
  input \ctl_rf_c1_rf_int_abt_msk_reg/NET0131  ;
  input \ctl_rf_c1_rf_int_err_msk_reg/NET0131  ;
  input \ctl_rf_c1_rf_int_tc1_msk_reg/NET0131  ;
  input \ctl_rf_c1_rf_int_tc_msk_reg/NET0131  ;
  input \ctl_rf_c1_rf_mode_reg/NET0131  ;
  input \ctl_rf_c1_rf_prot1_reg/NET0131  ;
  input \ctl_rf_c1_rf_prot2_reg/NET0131  ;
  input \ctl_rf_c1_rf_prot3_reg/NET0131  ;
  input \ctl_rf_c1_rf_sad_ctl0_reg/NET0131  ;
  input \ctl_rf_c1_rf_sad_ctl1_reg/NET0131  ;
  input \ctl_rf_c1_rf_src_sel_reg/NET0131  ;
  input \ctl_rf_c1_rf_src_sz_reg[0]/NET0131  ;
  input \ctl_rf_c1_rf_src_sz_reg[1]/NET0131  ;
  input \ctl_rf_c1_rf_src_sz_reg[2]/NET0131  ;
  input \ctl_rf_c1_rf_swidth_reg[0]/NET0131  ;
  input \ctl_rf_c1_rf_swidth_reg[1]/NET0131  ;
  input \ctl_rf_c1_rf_swidth_reg[2]/NET0131  ;
  input \ctl_rf_c1brbs_reg[16]/NET0131  ;
  input \ctl_rf_c1brbs_reg[17]/NET0131  ;
  input \ctl_rf_c1brbs_reg[18]/NET0131  ;
  input \ctl_rf_c1brbs_reg[19]/NET0131  ;
  input \ctl_rf_c1brbs_reg[20]/NET0131  ;
  input \ctl_rf_c1brbs_reg[21]/NET0131  ;
  input \ctl_rf_c1brbs_reg[22]/NET0131  ;
  input \ctl_rf_c1brbs_reg[23]/NET0131  ;
  input \ctl_rf_c1brbs_reg[24]/NET0131  ;
  input \ctl_rf_c1brbs_reg[25]/NET0131  ;
  input \ctl_rf_c1brbs_reg[26]/NET0131  ;
  input \ctl_rf_c1brbs_reg[27]/NET0131  ;
  input \ctl_rf_c1brbs_reg[28]/NET0131  ;
  input \ctl_rf_c1brbs_reg[29]/NET0131  ;
  input \ctl_rf_c1brbs_reg[30]/NET0131  ;
  input \ctl_rf_c1brbs_reg[31]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[16]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[17]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[18]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[19]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[20]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[21]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[22]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[23]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[24]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[25]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[26]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[27]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[28]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[29]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[30]/NET0131  ;
  input \ctl_rf_c1dmabs_reg[31]/NET0131  ;
  input \ctl_rf_c2_rf_autold_reg/NET0131  ;
  input \ctl_rf_c2_rf_ch_en_reg/NET0131  ;
  input \ctl_rf_c2_rf_chabt_reg/NET0131  ;
  input \ctl_rf_c2_rf_chdad_reg[0]/NET0131  ;
  input \ctl_rf_c2_rf_chdad_reg[10]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[11]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[12]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[13]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[14]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[15]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[16]/NET0131  ;
  input \ctl_rf_c2_rf_chdad_reg[17]/NET0131  ;
  input \ctl_rf_c2_rf_chdad_reg[18]/NET0131  ;
  input \ctl_rf_c2_rf_chdad_reg[19]/NET0131  ;
  input \ctl_rf_c2_rf_chdad_reg[1]/NET0131  ;
  input \ctl_rf_c2_rf_chdad_reg[20]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[21]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[22]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[23]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[24]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[25]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[26]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[27]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[28]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[29]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[2]/NET0131  ;
  input \ctl_rf_c2_rf_chdad_reg[30]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[31]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[3]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[4]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[5]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[6]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[7]/P0002  ;
  input \ctl_rf_c2_rf_chdad_reg[8]/NET0131  ;
  input \ctl_rf_c2_rf_chdad_reg[9]/P0002  ;
  input \ctl_rf_c2_rf_chllp_cnt_reg[0]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_cnt_reg[1]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_cnt_reg[2]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_cnt_reg[3]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_on_reg/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[0]/P0002  ;
  input \ctl_rf_c2_rf_chllp_reg[10]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[11]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[12]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[13]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[14]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[15]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[16]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[17]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[18]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[19]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[1]/P0002  ;
  input \ctl_rf_c2_rf_chllp_reg[20]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[21]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[22]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[23]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[24]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[25]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[26]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[27]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[28]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[29]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[2]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[30]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[31]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[3]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[4]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[5]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[6]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[7]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[8]/NET0131  ;
  input \ctl_rf_c2_rf_chllp_reg[9]/NET0131  ;
  input \ctl_rf_c2_rf_chllpen_reg/NET0131  ;
  input \ctl_rf_c2_rf_chpri_reg[0]/NET0131  ;
  input \ctl_rf_c2_rf_chpri_reg[1]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[0]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[10]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[11]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[12]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[13]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[14]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[15]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[16]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[17]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[18]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[19]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[1]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[20]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[21]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[22]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[23]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[24]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[25]/P0002  ;
  input \ctl_rf_c2_rf_chsad_reg[26]/P0002  ;
  input \ctl_rf_c2_rf_chsad_reg[27]/P0002  ;
  input \ctl_rf_c2_rf_chsad_reg[28]/P0002  ;
  input \ctl_rf_c2_rf_chsad_reg[29]/P0002  ;
  input \ctl_rf_c2_rf_chsad_reg[2]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[30]/P0002  ;
  input \ctl_rf_c2_rf_chsad_reg[31]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[3]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[4]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[5]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[6]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[7]/NET0131  ;
  input \ctl_rf_c2_rf_chsad_reg[8]/P0002  ;
  input \ctl_rf_c2_rf_chsad_reg[9]/NET0131  ;
  input \ctl_rf_c2_rf_chtsz_reg[0]/P0002  ;
  input \ctl_rf_c2_rf_chtsz_reg[10]/P0002  ;
  input \ctl_rf_c2_rf_chtsz_reg[11]/P0002  ;
  input \ctl_rf_c2_rf_chtsz_reg[1]/P0002  ;
  input \ctl_rf_c2_rf_chtsz_reg[2]/P0002  ;
  input \ctl_rf_c2_rf_chtsz_reg[3]/P0002  ;
  input \ctl_rf_c2_rf_chtsz_reg[4]/NET0131  ;
  input \ctl_rf_c2_rf_chtsz_reg[5]/NET0131  ;
  input \ctl_rf_c2_rf_chtsz_reg[6]/NET0131  ;
  input \ctl_rf_c2_rf_chtsz_reg[7]/NET0131  ;
  input \ctl_rf_c2_rf_chtsz_reg[8]/P0002  ;
  input \ctl_rf_c2_rf_chtsz_reg[9]/P0002  ;
  input \ctl_rf_c2_rf_dad_ctl0_reg/NET0131  ;
  input \ctl_rf_c2_rf_dad_ctl1_reg/NET0131  ;
  input \ctl_rf_c2_rf_dreqmode_reg/NET0131  ;
  input \ctl_rf_c2_rf_dst_sel_reg/NET0131  ;
  input \ctl_rf_c2_rf_dwidth_reg[0]/NET0131  ;
  input \ctl_rf_c2_rf_dwidth_reg[1]/NET0131  ;
  input \ctl_rf_c2_rf_dwidth_reg[2]/NET0131  ;
  input \ctl_rf_c2_rf_int_abt_msk_reg/NET0131  ;
  input \ctl_rf_c2_rf_int_err_msk_reg/NET0131  ;
  input \ctl_rf_c2_rf_int_tc1_msk_reg/NET0131  ;
  input \ctl_rf_c2_rf_int_tc_msk_reg/NET0131  ;
  input \ctl_rf_c2_rf_mode_reg/NET0131  ;
  input \ctl_rf_c2_rf_prot1_reg/NET0131  ;
  input \ctl_rf_c2_rf_prot2_reg/NET0131  ;
  input \ctl_rf_c2_rf_prot3_reg/NET0131  ;
  input \ctl_rf_c2_rf_sad_ctl0_reg/NET0131  ;
  input \ctl_rf_c2_rf_sad_ctl1_reg/NET0131  ;
  input \ctl_rf_c2_rf_src_sel_reg/NET0131  ;
  input \ctl_rf_c2_rf_src_sz_reg[0]/NET0131  ;
  input \ctl_rf_c2_rf_src_sz_reg[1]/NET0131  ;
  input \ctl_rf_c2_rf_src_sz_reg[2]/NET0131  ;
  input \ctl_rf_c2_rf_swidth_reg[0]/NET0131  ;
  input \ctl_rf_c2_rf_swidth_reg[1]/NET0131  ;
  input \ctl_rf_c2_rf_swidth_reg[2]/NET0131  ;
  input \ctl_rf_c2brbs_reg[16]/NET0131  ;
  input \ctl_rf_c2brbs_reg[17]/NET0131  ;
  input \ctl_rf_c2brbs_reg[18]/NET0131  ;
  input \ctl_rf_c2brbs_reg[19]/NET0131  ;
  input \ctl_rf_c2brbs_reg[20]/NET0131  ;
  input \ctl_rf_c2brbs_reg[21]/NET0131  ;
  input \ctl_rf_c2brbs_reg[22]/NET0131  ;
  input \ctl_rf_c2brbs_reg[23]/NET0131  ;
  input \ctl_rf_c2brbs_reg[24]/NET0131  ;
  input \ctl_rf_c2brbs_reg[25]/NET0131  ;
  input \ctl_rf_c2brbs_reg[26]/NET0131  ;
  input \ctl_rf_c2brbs_reg[27]/NET0131  ;
  input \ctl_rf_c2brbs_reg[28]/NET0131  ;
  input \ctl_rf_c2brbs_reg[29]/NET0131  ;
  input \ctl_rf_c2brbs_reg[30]/NET0131  ;
  input \ctl_rf_c2brbs_reg[31]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[16]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[17]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[18]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[19]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[20]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[21]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[22]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[23]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[24]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[25]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[26]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[27]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[28]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[29]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[30]/NET0131  ;
  input \ctl_rf_c2dmabs_reg[31]/NET0131  ;
  input \ctl_rf_c3_rf_autold_reg/NET0131  ;
  input \ctl_rf_c3_rf_ch_en_reg/NET0131  ;
  input \ctl_rf_c3_rf_chabt_reg/NET0131  ;
  input \ctl_rf_c3_rf_chdad_reg[0]/NET0131  ;
  input \ctl_rf_c3_rf_chdad_reg[10]/NET0131  ;
  input \ctl_rf_c3_rf_chdad_reg[11]/NET0131  ;
  input \ctl_rf_c3_rf_chdad_reg[12]/NET0131  ;
  input \ctl_rf_c3_rf_chdad_reg[13]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[14]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[15]/NET0131  ;
  input \ctl_rf_c3_rf_chdad_reg[16]/NET0131  ;
  input \ctl_rf_c3_rf_chdad_reg[17]/NET0131  ;
  input \ctl_rf_c3_rf_chdad_reg[18]/NET0131  ;
  input \ctl_rf_c3_rf_chdad_reg[19]/NET0131  ;
  input \ctl_rf_c3_rf_chdad_reg[1]/NET0131  ;
  input \ctl_rf_c3_rf_chdad_reg[20]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[21]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[22]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[23]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[24]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[25]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[26]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[27]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[28]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[29]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[2]/NET0131  ;
  input \ctl_rf_c3_rf_chdad_reg[30]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[31]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[3]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[4]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[5]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[6]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[7]/P0002  ;
  input \ctl_rf_c3_rf_chdad_reg[8]/NET0131  ;
  input \ctl_rf_c3_rf_chdad_reg[9]/P0002  ;
  input \ctl_rf_c3_rf_chllp_cnt_reg[0]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_cnt_reg[1]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_cnt_reg[2]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_cnt_reg[3]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_on_reg/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[0]/P0002  ;
  input \ctl_rf_c3_rf_chllp_reg[10]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[11]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[12]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[13]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[14]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[15]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[16]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[17]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[18]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[19]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[1]/P0002  ;
  input \ctl_rf_c3_rf_chllp_reg[20]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[21]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[22]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[23]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[24]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[25]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[26]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[27]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[28]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[29]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[2]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[30]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[31]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[3]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[4]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[5]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[6]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[7]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[8]/NET0131  ;
  input \ctl_rf_c3_rf_chllp_reg[9]/NET0131  ;
  input \ctl_rf_c3_rf_chllpen_reg/NET0131  ;
  input \ctl_rf_c3_rf_chpri_reg[0]/NET0131  ;
  input \ctl_rf_c3_rf_chpri_reg[1]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[0]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[10]/P0002  ;
  input \ctl_rf_c3_rf_chsad_reg[11]/P0002  ;
  input \ctl_rf_c3_rf_chsad_reg[12]/P0002  ;
  input \ctl_rf_c3_rf_chsad_reg[13]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[14]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[15]/P0002  ;
  input \ctl_rf_c3_rf_chsad_reg[16]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[17]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[18]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[19]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[1]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[20]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[21]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[22]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[23]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[24]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[25]/P0002  ;
  input \ctl_rf_c3_rf_chsad_reg[26]/P0002  ;
  input \ctl_rf_c3_rf_chsad_reg[27]/P0002  ;
  input \ctl_rf_c3_rf_chsad_reg[28]/P0002  ;
  input \ctl_rf_c3_rf_chsad_reg[29]/P0002  ;
  input \ctl_rf_c3_rf_chsad_reg[2]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[30]/P0002  ;
  input \ctl_rf_c3_rf_chsad_reg[31]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[3]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[4]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[5]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[6]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[7]/NET0131  ;
  input \ctl_rf_c3_rf_chsad_reg[8]/P0002  ;
  input \ctl_rf_c3_rf_chsad_reg[9]/NET0131  ;
  input \ctl_rf_c3_rf_chtsz_reg[0]/P0002  ;
  input \ctl_rf_c3_rf_chtsz_reg[10]/P0002  ;
  input \ctl_rf_c3_rf_chtsz_reg[11]/P0002  ;
  input \ctl_rf_c3_rf_chtsz_reg[1]/P0002  ;
  input \ctl_rf_c3_rf_chtsz_reg[2]/P0002  ;
  input \ctl_rf_c3_rf_chtsz_reg[3]/P0002  ;
  input \ctl_rf_c3_rf_chtsz_reg[4]/NET0131  ;
  input \ctl_rf_c3_rf_chtsz_reg[5]/NET0131  ;
  input \ctl_rf_c3_rf_chtsz_reg[6]/NET0131  ;
  input \ctl_rf_c3_rf_chtsz_reg[7]/NET0131  ;
  input \ctl_rf_c3_rf_chtsz_reg[8]/P0002  ;
  input \ctl_rf_c3_rf_chtsz_reg[9]/P0002  ;
  input \ctl_rf_c3_rf_dad_ctl0_reg/NET0131  ;
  input \ctl_rf_c3_rf_dad_ctl1_reg/NET0131  ;
  input \ctl_rf_c3_rf_dreqmode_reg/NET0131  ;
  input \ctl_rf_c3_rf_dst_sel_reg/NET0131  ;
  input \ctl_rf_c3_rf_dwidth_reg[0]/NET0131  ;
  input \ctl_rf_c3_rf_dwidth_reg[1]/NET0131  ;
  input \ctl_rf_c3_rf_dwidth_reg[2]/NET0131  ;
  input \ctl_rf_c3_rf_int_abt_msk_reg/NET0131  ;
  input \ctl_rf_c3_rf_int_err_msk_reg/NET0131  ;
  input \ctl_rf_c3_rf_int_tc1_msk_reg/NET0131  ;
  input \ctl_rf_c3_rf_int_tc_msk_reg/NET0131  ;
  input \ctl_rf_c3_rf_mode_reg/NET0131  ;
  input \ctl_rf_c3_rf_prot1_reg/NET0131  ;
  input \ctl_rf_c3_rf_prot2_reg/NET0131  ;
  input \ctl_rf_c3_rf_prot3_reg/NET0131  ;
  input \ctl_rf_c3_rf_sad_ctl0_reg/NET0131  ;
  input \ctl_rf_c3_rf_sad_ctl1_reg/NET0131  ;
  input \ctl_rf_c3_rf_src_sel_reg/NET0131  ;
  input \ctl_rf_c3_rf_src_sz_reg[0]/NET0131  ;
  input \ctl_rf_c3_rf_src_sz_reg[1]/NET0131  ;
  input \ctl_rf_c3_rf_src_sz_reg[2]/NET0131  ;
  input \ctl_rf_c3_rf_swidth_reg[0]/NET0131  ;
  input \ctl_rf_c3_rf_swidth_reg[1]/NET0131  ;
  input \ctl_rf_c3_rf_swidth_reg[2]/NET0131  ;
  input \ctl_rf_c3brbs_reg[16]/NET0131  ;
  input \ctl_rf_c3brbs_reg[17]/NET0131  ;
  input \ctl_rf_c3brbs_reg[18]/NET0131  ;
  input \ctl_rf_c3brbs_reg[19]/NET0131  ;
  input \ctl_rf_c3brbs_reg[20]/NET0131  ;
  input \ctl_rf_c3brbs_reg[21]/NET0131  ;
  input \ctl_rf_c3brbs_reg[22]/NET0131  ;
  input \ctl_rf_c3brbs_reg[23]/NET0131  ;
  input \ctl_rf_c3brbs_reg[24]/NET0131  ;
  input \ctl_rf_c3brbs_reg[25]/NET0131  ;
  input \ctl_rf_c3brbs_reg[26]/NET0131  ;
  input \ctl_rf_c3brbs_reg[27]/NET0131  ;
  input \ctl_rf_c3brbs_reg[28]/NET0131  ;
  input \ctl_rf_c3brbs_reg[29]/NET0131  ;
  input \ctl_rf_c3brbs_reg[30]/NET0131  ;
  input \ctl_rf_c3brbs_reg[31]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[16]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[17]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[18]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[19]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[20]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[21]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[22]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[23]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[24]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[25]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[26]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[27]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[28]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[29]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[30]/NET0131  ;
  input \ctl_rf_c3dmabs_reg[31]/NET0131  ;
  input \ctl_rf_c4_rf_autold_reg/NET0131  ;
  input \ctl_rf_c4_rf_ch_en_reg/NET0131  ;
  input \ctl_rf_c4_rf_chabt_reg/NET0131  ;
  input \ctl_rf_c4_rf_chdad_reg[0]/NET0131  ;
  input \ctl_rf_c4_rf_chdad_reg[10]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[11]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[12]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[13]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[14]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[15]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[16]/NET0131  ;
  input \ctl_rf_c4_rf_chdad_reg[17]/NET0131  ;
  input \ctl_rf_c4_rf_chdad_reg[18]/NET0131  ;
  input \ctl_rf_c4_rf_chdad_reg[19]/NET0131  ;
  input \ctl_rf_c4_rf_chdad_reg[1]/NET0131  ;
  input \ctl_rf_c4_rf_chdad_reg[20]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[21]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[22]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[23]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[24]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[25]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[26]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[27]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[28]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[29]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[2]/NET0131  ;
  input \ctl_rf_c4_rf_chdad_reg[30]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[31]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[3]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[4]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[5]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[6]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[7]/P0002  ;
  input \ctl_rf_c4_rf_chdad_reg[8]/NET0131  ;
  input \ctl_rf_c4_rf_chdad_reg[9]/P0002  ;
  input \ctl_rf_c4_rf_chllp_cnt_reg[0]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_cnt_reg[1]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_cnt_reg[2]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_cnt_reg[3]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_on_reg/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[0]/P0002  ;
  input \ctl_rf_c4_rf_chllp_reg[10]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[11]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[12]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[13]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[14]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[15]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[16]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[17]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[18]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[19]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[1]/P0002  ;
  input \ctl_rf_c4_rf_chllp_reg[20]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[21]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[22]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[23]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[24]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[25]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[26]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[27]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[28]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[29]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[2]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[30]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[31]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[3]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[4]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[5]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[6]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[7]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[8]/NET0131  ;
  input \ctl_rf_c4_rf_chllp_reg[9]/NET0131  ;
  input \ctl_rf_c4_rf_chllpen_reg/NET0131  ;
  input \ctl_rf_c4_rf_chpri_reg[0]/NET0131  ;
  input \ctl_rf_c4_rf_chpri_reg[1]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[0]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[10]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[11]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[12]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[13]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[14]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[15]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[16]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[17]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[18]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[19]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[1]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[20]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[21]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[22]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[23]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[24]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[25]/P0002  ;
  input \ctl_rf_c4_rf_chsad_reg[26]/P0002  ;
  input \ctl_rf_c4_rf_chsad_reg[27]/P0002  ;
  input \ctl_rf_c4_rf_chsad_reg[28]/P0002  ;
  input \ctl_rf_c4_rf_chsad_reg[29]/P0002  ;
  input \ctl_rf_c4_rf_chsad_reg[2]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[30]/P0002  ;
  input \ctl_rf_c4_rf_chsad_reg[31]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[3]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[4]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[5]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[6]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[7]/NET0131  ;
  input \ctl_rf_c4_rf_chsad_reg[8]/P0002  ;
  input \ctl_rf_c4_rf_chsad_reg[9]/NET0131  ;
  input \ctl_rf_c4_rf_chtsz_reg[0]/P0002  ;
  input \ctl_rf_c4_rf_chtsz_reg[10]/P0002  ;
  input \ctl_rf_c4_rf_chtsz_reg[11]/P0002  ;
  input \ctl_rf_c4_rf_chtsz_reg[1]/P0002  ;
  input \ctl_rf_c4_rf_chtsz_reg[2]/P0002  ;
  input \ctl_rf_c4_rf_chtsz_reg[3]/P0002  ;
  input \ctl_rf_c4_rf_chtsz_reg[4]/NET0131  ;
  input \ctl_rf_c4_rf_chtsz_reg[5]/NET0131  ;
  input \ctl_rf_c4_rf_chtsz_reg[6]/NET0131  ;
  input \ctl_rf_c4_rf_chtsz_reg[7]/NET0131  ;
  input \ctl_rf_c4_rf_chtsz_reg[8]/P0002  ;
  input \ctl_rf_c4_rf_chtsz_reg[9]/P0002  ;
  input \ctl_rf_c4_rf_dad_ctl0_reg/NET0131  ;
  input \ctl_rf_c4_rf_dad_ctl1_reg/NET0131  ;
  input \ctl_rf_c4_rf_dreqmode_reg/NET0131  ;
  input \ctl_rf_c4_rf_dst_sel_reg/NET0131  ;
  input \ctl_rf_c4_rf_dwidth_reg[0]/NET0131  ;
  input \ctl_rf_c4_rf_dwidth_reg[1]/NET0131  ;
  input \ctl_rf_c4_rf_dwidth_reg[2]/NET0131  ;
  input \ctl_rf_c4_rf_int_abt_msk_reg/NET0131  ;
  input \ctl_rf_c4_rf_int_err_msk_reg/NET0131  ;
  input \ctl_rf_c4_rf_int_tc1_msk_reg/NET0131  ;
  input \ctl_rf_c4_rf_int_tc_msk_reg/NET0131  ;
  input \ctl_rf_c4_rf_mode_reg/NET0131  ;
  input \ctl_rf_c4_rf_prot1_reg/NET0131  ;
  input \ctl_rf_c4_rf_prot2_reg/NET0131  ;
  input \ctl_rf_c4_rf_prot3_reg/NET0131  ;
  input \ctl_rf_c4_rf_sad_ctl0_reg/NET0131  ;
  input \ctl_rf_c4_rf_sad_ctl1_reg/NET0131  ;
  input \ctl_rf_c4_rf_src_sel_reg/NET0131  ;
  input \ctl_rf_c4_rf_src_sz_reg[0]/NET0131  ;
  input \ctl_rf_c4_rf_src_sz_reg[1]/NET0131  ;
  input \ctl_rf_c4_rf_src_sz_reg[2]/NET0131  ;
  input \ctl_rf_c4_rf_swidth_reg[0]/NET0131  ;
  input \ctl_rf_c4_rf_swidth_reg[1]/NET0131  ;
  input \ctl_rf_c4_rf_swidth_reg[2]/NET0131  ;
  input \ctl_rf_c4brbs_reg[16]/NET0131  ;
  input \ctl_rf_c4brbs_reg[17]/NET0131  ;
  input \ctl_rf_c4brbs_reg[18]/NET0131  ;
  input \ctl_rf_c4brbs_reg[19]/NET0131  ;
  input \ctl_rf_c4brbs_reg[20]/NET0131  ;
  input \ctl_rf_c4brbs_reg[21]/NET0131  ;
  input \ctl_rf_c4brbs_reg[22]/NET0131  ;
  input \ctl_rf_c4brbs_reg[23]/NET0131  ;
  input \ctl_rf_c4brbs_reg[24]/NET0131  ;
  input \ctl_rf_c4brbs_reg[25]/NET0131  ;
  input \ctl_rf_c4brbs_reg[26]/NET0131  ;
  input \ctl_rf_c4brbs_reg[27]/NET0131  ;
  input \ctl_rf_c4brbs_reg[28]/NET0131  ;
  input \ctl_rf_c4brbs_reg[29]/NET0131  ;
  input \ctl_rf_c4brbs_reg[30]/NET0131  ;
  input \ctl_rf_c4brbs_reg[31]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[16]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[17]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[18]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[19]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[20]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[21]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[22]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[23]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[24]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[25]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[26]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[27]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[28]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[29]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[30]/NET0131  ;
  input \ctl_rf_c4dmabs_reg[31]/NET0131  ;
  input \ctl_rf_c5_rf_autold_reg/NET0131  ;
  input \ctl_rf_c5_rf_ch_en_reg/NET0131  ;
  input \ctl_rf_c5_rf_chabt_reg/NET0131  ;
  input \ctl_rf_c5_rf_chdad_reg[0]/NET0131  ;
  input \ctl_rf_c5_rf_chdad_reg[10]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[11]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[12]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[13]/NET0131  ;
  input \ctl_rf_c5_rf_chdad_reg[14]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[15]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[16]/NET0131  ;
  input \ctl_rf_c5_rf_chdad_reg[17]/NET0131  ;
  input \ctl_rf_c5_rf_chdad_reg[18]/NET0131  ;
  input \ctl_rf_c5_rf_chdad_reg[19]/NET0131  ;
  input \ctl_rf_c5_rf_chdad_reg[1]/NET0131  ;
  input \ctl_rf_c5_rf_chdad_reg[20]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[21]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[22]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[23]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[24]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[25]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[26]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[27]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[28]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[29]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[2]/NET0131  ;
  input \ctl_rf_c5_rf_chdad_reg[30]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[31]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[3]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[4]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[5]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[6]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[7]/P0002  ;
  input \ctl_rf_c5_rf_chdad_reg[8]/NET0131  ;
  input \ctl_rf_c5_rf_chdad_reg[9]/P0002  ;
  input \ctl_rf_c5_rf_chllp_cnt_reg[0]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_cnt_reg[1]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_cnt_reg[2]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_cnt_reg[3]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_on_reg/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[0]/P0002  ;
  input \ctl_rf_c5_rf_chllp_reg[10]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[11]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[12]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[13]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[14]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[15]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[16]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[17]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[18]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[19]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[1]/P0002  ;
  input \ctl_rf_c5_rf_chllp_reg[20]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[21]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[22]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[23]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[24]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[25]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[26]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[27]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[28]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[29]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[2]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[30]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[31]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[3]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[4]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[5]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[6]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[7]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[8]/NET0131  ;
  input \ctl_rf_c5_rf_chllp_reg[9]/NET0131  ;
  input \ctl_rf_c5_rf_chllpen_reg/NET0131  ;
  input \ctl_rf_c5_rf_chpri_reg[0]/NET0131  ;
  input \ctl_rf_c5_rf_chpri_reg[1]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[0]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[10]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[11]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[12]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[13]/P0002  ;
  input \ctl_rf_c5_rf_chsad_reg[14]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[15]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[16]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[17]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[18]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[19]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[1]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[20]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[21]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[22]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[23]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[24]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[25]/P0002  ;
  input \ctl_rf_c5_rf_chsad_reg[26]/P0002  ;
  input \ctl_rf_c5_rf_chsad_reg[27]/P0002  ;
  input \ctl_rf_c5_rf_chsad_reg[28]/P0002  ;
  input \ctl_rf_c5_rf_chsad_reg[29]/P0002  ;
  input \ctl_rf_c5_rf_chsad_reg[2]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[30]/P0002  ;
  input \ctl_rf_c5_rf_chsad_reg[31]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[3]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[4]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[5]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[6]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[7]/NET0131  ;
  input \ctl_rf_c5_rf_chsad_reg[8]/P0002  ;
  input \ctl_rf_c5_rf_chsad_reg[9]/NET0131  ;
  input \ctl_rf_c5_rf_chtsz_reg[0]/P0002  ;
  input \ctl_rf_c5_rf_chtsz_reg[10]/P0002  ;
  input \ctl_rf_c5_rf_chtsz_reg[11]/P0002  ;
  input \ctl_rf_c5_rf_chtsz_reg[1]/P0002  ;
  input \ctl_rf_c5_rf_chtsz_reg[2]/P0002  ;
  input \ctl_rf_c5_rf_chtsz_reg[3]/P0002  ;
  input \ctl_rf_c5_rf_chtsz_reg[4]/NET0131  ;
  input \ctl_rf_c5_rf_chtsz_reg[5]/NET0131  ;
  input \ctl_rf_c5_rf_chtsz_reg[6]/NET0131  ;
  input \ctl_rf_c5_rf_chtsz_reg[7]/NET0131  ;
  input \ctl_rf_c5_rf_chtsz_reg[8]/P0002  ;
  input \ctl_rf_c5_rf_chtsz_reg[9]/P0002  ;
  input \ctl_rf_c5_rf_dad_ctl0_reg/NET0131  ;
  input \ctl_rf_c5_rf_dad_ctl1_reg/NET0131  ;
  input \ctl_rf_c5_rf_dreqmode_reg/NET0131  ;
  input \ctl_rf_c5_rf_dst_sel_reg/NET0131  ;
  input \ctl_rf_c5_rf_dwidth_reg[0]/NET0131  ;
  input \ctl_rf_c5_rf_dwidth_reg[1]/NET0131  ;
  input \ctl_rf_c5_rf_dwidth_reg[2]/NET0131  ;
  input \ctl_rf_c5_rf_int_abt_msk_reg/NET0131  ;
  input \ctl_rf_c5_rf_int_err_msk_reg/NET0131  ;
  input \ctl_rf_c5_rf_int_tc1_msk_reg/NET0131  ;
  input \ctl_rf_c5_rf_int_tc_msk_reg/NET0131  ;
  input \ctl_rf_c5_rf_mode_reg/NET0131  ;
  input \ctl_rf_c5_rf_prot1_reg/NET0131  ;
  input \ctl_rf_c5_rf_prot2_reg/NET0131  ;
  input \ctl_rf_c5_rf_prot3_reg/NET0131  ;
  input \ctl_rf_c5_rf_sad_ctl0_reg/NET0131  ;
  input \ctl_rf_c5_rf_sad_ctl1_reg/NET0131  ;
  input \ctl_rf_c5_rf_src_sel_reg/NET0131  ;
  input \ctl_rf_c5_rf_src_sz_reg[0]/NET0131  ;
  input \ctl_rf_c5_rf_src_sz_reg[1]/NET0131  ;
  input \ctl_rf_c5_rf_src_sz_reg[2]/NET0131  ;
  input \ctl_rf_c5_rf_swidth_reg[0]/NET0131  ;
  input \ctl_rf_c5_rf_swidth_reg[1]/NET0131  ;
  input \ctl_rf_c5_rf_swidth_reg[2]/NET0131  ;
  input \ctl_rf_c5brbs_reg[16]/NET0131  ;
  input \ctl_rf_c5brbs_reg[17]/NET0131  ;
  input \ctl_rf_c5brbs_reg[18]/NET0131  ;
  input \ctl_rf_c5brbs_reg[19]/NET0131  ;
  input \ctl_rf_c5brbs_reg[20]/NET0131  ;
  input \ctl_rf_c5brbs_reg[21]/NET0131  ;
  input \ctl_rf_c5brbs_reg[22]/NET0131  ;
  input \ctl_rf_c5brbs_reg[23]/NET0131  ;
  input \ctl_rf_c5brbs_reg[24]/NET0131  ;
  input \ctl_rf_c5brbs_reg[25]/NET0131  ;
  input \ctl_rf_c5brbs_reg[26]/NET0131  ;
  input \ctl_rf_c5brbs_reg[27]/NET0131  ;
  input \ctl_rf_c5brbs_reg[28]/NET0131  ;
  input \ctl_rf_c5brbs_reg[29]/NET0131  ;
  input \ctl_rf_c5brbs_reg[30]/NET0131  ;
  input \ctl_rf_c5brbs_reg[31]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[16]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[17]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[18]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[19]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[20]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[21]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[22]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[23]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[24]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[25]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[26]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[27]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[28]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[29]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[30]/NET0131  ;
  input \ctl_rf_c5dmabs_reg[31]/NET0131  ;
  input \ctl_rf_c6_rf_autold_reg/NET0131  ;
  input \ctl_rf_c6_rf_ch_en_reg/NET0131  ;
  input \ctl_rf_c6_rf_chabt_reg/NET0131  ;
  input \ctl_rf_c6_rf_chdad_reg[0]/NET0131  ;
  input \ctl_rf_c6_rf_chdad_reg[10]/NET0131  ;
  input \ctl_rf_c6_rf_chdad_reg[11]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[12]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[13]/NET0131  ;
  input \ctl_rf_c6_rf_chdad_reg[14]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[15]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[16]/NET0131  ;
  input \ctl_rf_c6_rf_chdad_reg[17]/NET0131  ;
  input \ctl_rf_c6_rf_chdad_reg[18]/NET0131  ;
  input \ctl_rf_c6_rf_chdad_reg[19]/NET0131  ;
  input \ctl_rf_c6_rf_chdad_reg[1]/NET0131  ;
  input \ctl_rf_c6_rf_chdad_reg[20]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[21]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[22]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[23]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[24]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[25]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[26]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[27]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[28]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[29]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[2]/NET0131  ;
  input \ctl_rf_c6_rf_chdad_reg[30]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[31]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[3]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[4]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[5]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[6]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[7]/P0002  ;
  input \ctl_rf_c6_rf_chdad_reg[8]/NET0131  ;
  input \ctl_rf_c6_rf_chdad_reg[9]/P0002  ;
  input \ctl_rf_c6_rf_chllp_cnt_reg[0]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_cnt_reg[1]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_cnt_reg[2]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_cnt_reg[3]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_on_reg/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[0]/P0002  ;
  input \ctl_rf_c6_rf_chllp_reg[10]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[11]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[12]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[13]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[14]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[15]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[16]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[17]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[18]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[19]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[1]/P0002  ;
  input \ctl_rf_c6_rf_chllp_reg[20]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[21]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[22]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[23]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[24]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[25]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[26]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[27]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[28]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[29]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[2]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[30]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[31]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[3]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[4]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[5]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[6]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[7]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[8]/NET0131  ;
  input \ctl_rf_c6_rf_chllp_reg[9]/NET0131  ;
  input \ctl_rf_c6_rf_chllpen_reg/NET0131  ;
  input \ctl_rf_c6_rf_chpri_reg[0]/NET0131  ;
  input \ctl_rf_c6_rf_chpri_reg[1]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[0]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[10]/P0002  ;
  input \ctl_rf_c6_rf_chsad_reg[11]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[12]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[13]/P0002  ;
  input \ctl_rf_c6_rf_chsad_reg[14]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[15]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[16]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[17]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[18]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[19]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[1]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[20]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[21]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[22]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[23]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[24]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[25]/P0002  ;
  input \ctl_rf_c6_rf_chsad_reg[26]/P0002  ;
  input \ctl_rf_c6_rf_chsad_reg[27]/P0002  ;
  input \ctl_rf_c6_rf_chsad_reg[28]/P0002  ;
  input \ctl_rf_c6_rf_chsad_reg[29]/P0002  ;
  input \ctl_rf_c6_rf_chsad_reg[2]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[30]/P0002  ;
  input \ctl_rf_c6_rf_chsad_reg[31]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[3]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[4]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[5]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[6]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[7]/NET0131  ;
  input \ctl_rf_c6_rf_chsad_reg[8]/P0002  ;
  input \ctl_rf_c6_rf_chsad_reg[9]/NET0131  ;
  input \ctl_rf_c6_rf_chtsz_reg[0]/P0002  ;
  input \ctl_rf_c6_rf_chtsz_reg[10]/P0002  ;
  input \ctl_rf_c6_rf_chtsz_reg[11]/P0002  ;
  input \ctl_rf_c6_rf_chtsz_reg[1]/P0002  ;
  input \ctl_rf_c6_rf_chtsz_reg[2]/P0002  ;
  input \ctl_rf_c6_rf_chtsz_reg[3]/P0002  ;
  input \ctl_rf_c6_rf_chtsz_reg[4]/NET0131  ;
  input \ctl_rf_c6_rf_chtsz_reg[5]/NET0131  ;
  input \ctl_rf_c6_rf_chtsz_reg[6]/NET0131  ;
  input \ctl_rf_c6_rf_chtsz_reg[7]/NET0131  ;
  input \ctl_rf_c6_rf_chtsz_reg[8]/P0002  ;
  input \ctl_rf_c6_rf_chtsz_reg[9]/P0002  ;
  input \ctl_rf_c6_rf_dad_ctl0_reg/NET0131  ;
  input \ctl_rf_c6_rf_dad_ctl1_reg/NET0131  ;
  input \ctl_rf_c6_rf_dreqmode_reg/NET0131  ;
  input \ctl_rf_c6_rf_dst_sel_reg/NET0131  ;
  input \ctl_rf_c6_rf_dwidth_reg[0]/NET0131  ;
  input \ctl_rf_c6_rf_dwidth_reg[1]/NET0131  ;
  input \ctl_rf_c6_rf_dwidth_reg[2]/NET0131  ;
  input \ctl_rf_c6_rf_int_abt_msk_reg/NET0131  ;
  input \ctl_rf_c6_rf_int_err_msk_reg/NET0131  ;
  input \ctl_rf_c6_rf_int_tc1_msk_reg/NET0131  ;
  input \ctl_rf_c6_rf_int_tc_msk_reg/NET0131  ;
  input \ctl_rf_c6_rf_mode_reg/NET0131  ;
  input \ctl_rf_c6_rf_prot1_reg/NET0131  ;
  input \ctl_rf_c6_rf_prot2_reg/NET0131  ;
  input \ctl_rf_c6_rf_prot3_reg/NET0131  ;
  input \ctl_rf_c6_rf_sad_ctl0_reg/NET0131  ;
  input \ctl_rf_c6_rf_sad_ctl1_reg/NET0131  ;
  input \ctl_rf_c6_rf_src_sel_reg/NET0131  ;
  input \ctl_rf_c6_rf_src_sz_reg[0]/NET0131  ;
  input \ctl_rf_c6_rf_src_sz_reg[1]/NET0131  ;
  input \ctl_rf_c6_rf_src_sz_reg[2]/NET0131  ;
  input \ctl_rf_c6_rf_swidth_reg[0]/NET0131  ;
  input \ctl_rf_c6_rf_swidth_reg[1]/NET0131  ;
  input \ctl_rf_c6_rf_swidth_reg[2]/NET0131  ;
  input \ctl_rf_c6brbs_reg[16]/NET0131  ;
  input \ctl_rf_c6brbs_reg[17]/NET0131  ;
  input \ctl_rf_c6brbs_reg[18]/NET0131  ;
  input \ctl_rf_c6brbs_reg[19]/NET0131  ;
  input \ctl_rf_c6brbs_reg[20]/NET0131  ;
  input \ctl_rf_c6brbs_reg[21]/NET0131  ;
  input \ctl_rf_c6brbs_reg[22]/NET0131  ;
  input \ctl_rf_c6brbs_reg[23]/NET0131  ;
  input \ctl_rf_c6brbs_reg[24]/NET0131  ;
  input \ctl_rf_c6brbs_reg[25]/NET0131  ;
  input \ctl_rf_c6brbs_reg[26]/NET0131  ;
  input \ctl_rf_c6brbs_reg[27]/NET0131  ;
  input \ctl_rf_c6brbs_reg[28]/NET0131  ;
  input \ctl_rf_c6brbs_reg[29]/NET0131  ;
  input \ctl_rf_c6brbs_reg[30]/NET0131  ;
  input \ctl_rf_c6brbs_reg[31]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[16]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[17]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[18]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[19]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[20]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[21]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[22]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[23]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[24]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[25]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[26]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[27]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[28]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[29]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[30]/NET0131  ;
  input \ctl_rf_c6dmabs_reg[31]/NET0131  ;
  input \ctl_rf_c7_rf_autold_reg/NET0131  ;
  input \ctl_rf_c7_rf_ch_en_reg/NET0131  ;
  input \ctl_rf_c7_rf_chabt_reg/NET0131  ;
  input \ctl_rf_c7_rf_chdad_reg[0]/NET0131  ;
  input \ctl_rf_c7_rf_chdad_reg[10]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[11]/NET0131  ;
  input \ctl_rf_c7_rf_chdad_reg[12]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[13]/NET0131  ;
  input \ctl_rf_c7_rf_chdad_reg[14]/NET0131  ;
  input \ctl_rf_c7_rf_chdad_reg[15]/NET0131  ;
  input \ctl_rf_c7_rf_chdad_reg[16]/NET0131  ;
  input \ctl_rf_c7_rf_chdad_reg[17]/NET0131  ;
  input \ctl_rf_c7_rf_chdad_reg[18]/NET0131  ;
  input \ctl_rf_c7_rf_chdad_reg[19]/NET0131  ;
  input \ctl_rf_c7_rf_chdad_reg[1]/NET0131  ;
  input \ctl_rf_c7_rf_chdad_reg[20]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[21]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[22]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[23]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[24]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[25]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[26]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[27]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[28]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[29]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[2]/NET0131  ;
  input \ctl_rf_c7_rf_chdad_reg[30]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[31]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[3]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[4]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[5]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[6]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[7]/P0002  ;
  input \ctl_rf_c7_rf_chdad_reg[8]/NET0131  ;
  input \ctl_rf_c7_rf_chdad_reg[9]/P0002  ;
  input \ctl_rf_c7_rf_chllp_cnt_reg[0]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_cnt_reg[1]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_cnt_reg[2]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_cnt_reg[3]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_on_reg/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[0]/P0002  ;
  input \ctl_rf_c7_rf_chllp_reg[10]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[11]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[12]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[13]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[14]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[15]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[16]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[17]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[18]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[19]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[1]/P0002  ;
  input \ctl_rf_c7_rf_chllp_reg[20]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[21]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[22]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[23]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[24]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[25]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[26]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[27]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[28]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[29]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[2]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[30]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[31]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[3]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[4]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[5]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[6]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[7]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[8]/NET0131  ;
  input \ctl_rf_c7_rf_chllp_reg[9]/NET0131  ;
  input \ctl_rf_c7_rf_chllpen_reg/NET0131  ;
  input \ctl_rf_c7_rf_chpri_reg[0]/NET0131  ;
  input \ctl_rf_c7_rf_chpri_reg[1]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[0]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[10]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[11]/P0002  ;
  input \ctl_rf_c7_rf_chsad_reg[12]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[13]/P0002  ;
  input \ctl_rf_c7_rf_chsad_reg[14]/P0002  ;
  input \ctl_rf_c7_rf_chsad_reg[15]/P0002  ;
  input \ctl_rf_c7_rf_chsad_reg[16]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[17]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[18]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[19]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[1]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[20]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[21]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[22]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[23]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[24]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[25]/P0002  ;
  input \ctl_rf_c7_rf_chsad_reg[26]/P0002  ;
  input \ctl_rf_c7_rf_chsad_reg[27]/P0002  ;
  input \ctl_rf_c7_rf_chsad_reg[28]/P0002  ;
  input \ctl_rf_c7_rf_chsad_reg[29]/P0002  ;
  input \ctl_rf_c7_rf_chsad_reg[2]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[30]/P0002  ;
  input \ctl_rf_c7_rf_chsad_reg[31]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[3]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[4]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[5]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[6]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[7]/NET0131  ;
  input \ctl_rf_c7_rf_chsad_reg[8]/P0002  ;
  input \ctl_rf_c7_rf_chsad_reg[9]/NET0131  ;
  input \ctl_rf_c7_rf_chtsz_reg[0]/P0002  ;
  input \ctl_rf_c7_rf_chtsz_reg[10]/P0002  ;
  input \ctl_rf_c7_rf_chtsz_reg[11]/P0002  ;
  input \ctl_rf_c7_rf_chtsz_reg[1]/P0002  ;
  input \ctl_rf_c7_rf_chtsz_reg[2]/P0002  ;
  input \ctl_rf_c7_rf_chtsz_reg[3]/P0002  ;
  input \ctl_rf_c7_rf_chtsz_reg[4]/NET0131  ;
  input \ctl_rf_c7_rf_chtsz_reg[5]/NET0131  ;
  input \ctl_rf_c7_rf_chtsz_reg[6]/NET0131  ;
  input \ctl_rf_c7_rf_chtsz_reg[7]/NET0131  ;
  input \ctl_rf_c7_rf_chtsz_reg[8]/P0002  ;
  input \ctl_rf_c7_rf_chtsz_reg[9]/P0002  ;
  input \ctl_rf_c7_rf_dad_ctl0_reg/NET0131  ;
  input \ctl_rf_c7_rf_dad_ctl1_reg/NET0131  ;
  input \ctl_rf_c7_rf_dreqmode_reg/NET0131  ;
  input \ctl_rf_c7_rf_dst_sel_reg/NET0131  ;
  input \ctl_rf_c7_rf_dwidth_reg[0]/NET0131  ;
  input \ctl_rf_c7_rf_dwidth_reg[1]/NET0131  ;
  input \ctl_rf_c7_rf_dwidth_reg[2]/NET0131  ;
  input \ctl_rf_c7_rf_int_abt_msk_reg/NET0131  ;
  input \ctl_rf_c7_rf_int_err_msk_reg/NET0131  ;
  input \ctl_rf_c7_rf_int_tc1_msk_reg/NET0131  ;
  input \ctl_rf_c7_rf_int_tc_msk_reg/NET0131  ;
  input \ctl_rf_c7_rf_mode_reg/NET0131  ;
  input \ctl_rf_c7_rf_prot1_reg/NET0131  ;
  input \ctl_rf_c7_rf_prot2_reg/NET0131  ;
  input \ctl_rf_c7_rf_prot3_reg/NET0131  ;
  input \ctl_rf_c7_rf_sad_ctl0_reg/NET0131  ;
  input \ctl_rf_c7_rf_sad_ctl1_reg/NET0131  ;
  input \ctl_rf_c7_rf_src_sel_reg/NET0131  ;
  input \ctl_rf_c7_rf_src_sz_reg[0]/NET0131  ;
  input \ctl_rf_c7_rf_src_sz_reg[1]/NET0131  ;
  input \ctl_rf_c7_rf_src_sz_reg[2]/NET0131  ;
  input \ctl_rf_c7_rf_swidth_reg[0]/NET0131  ;
  input \ctl_rf_c7_rf_swidth_reg[1]/NET0131  ;
  input \ctl_rf_c7_rf_swidth_reg[2]/NET0131  ;
  input \ctl_rf_c7brbs_reg[16]/NET0131  ;
  input \ctl_rf_c7brbs_reg[17]/NET0131  ;
  input \ctl_rf_c7brbs_reg[18]/NET0131  ;
  input \ctl_rf_c7brbs_reg[19]/NET0131  ;
  input \ctl_rf_c7brbs_reg[20]/NET0131  ;
  input \ctl_rf_c7brbs_reg[21]/NET0131  ;
  input \ctl_rf_c7brbs_reg[22]/NET0131  ;
  input \ctl_rf_c7brbs_reg[23]/NET0131  ;
  input \ctl_rf_c7brbs_reg[24]/NET0131  ;
  input \ctl_rf_c7brbs_reg[25]/NET0131  ;
  input \ctl_rf_c7brbs_reg[26]/NET0131  ;
  input \ctl_rf_c7brbs_reg[27]/NET0131  ;
  input \ctl_rf_c7brbs_reg[28]/NET0131  ;
  input \ctl_rf_c7brbs_reg[29]/NET0131  ;
  input \ctl_rf_c7brbs_reg[30]/NET0131  ;
  input \ctl_rf_c7brbs_reg[31]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[16]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[17]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[18]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[19]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[20]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[21]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[22]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[23]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[24]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[25]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[26]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[27]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[28]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[29]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[30]/NET0131  ;
  input \ctl_rf_c7dmabs_reg[31]/NET0131  ;
  input \ctl_rf_dmacen_reg/NET0131  ;
  input \ctl_rf_m0end_reg/NET0131  ;
  input \ctl_rf_m1end_reg/NET0131  ;
  input \ctl_rf_rf_sel_d1_reg/NET0131  ;
  input \ctl_rf_sync_reg[0]/NET0131  ;
  input \ctl_rf_sync_reg[1]/NET0131  ;
  input \ctl_rf_sync_reg[2]/NET0131  ;
  input \ctl_rf_sync_reg[3]/NET0131  ;
  input \ctl_rf_sync_reg[4]/NET0131  ;
  input \ctl_rf_sync_reg[5]/NET0131  ;
  input \ctl_rf_sync_reg[6]/NET0131  ;
  input \ctl_rf_sync_reg[7]/NET0131  ;
  input \ctl_rf_tc_reg[0]/NET0131  ;
  input \ctl_rf_tc_reg[1]/NET0131  ;
  input \ctl_rf_tc_reg[2]/NET0131  ;
  input \ctl_rf_tc_reg[3]/NET0131  ;
  input \ctl_rf_tc_reg[4]/NET0131  ;
  input \ctl_rf_tc_reg[5]/NET0131  ;
  input \ctl_rf_tc_reg[6]/NET0131  ;
  input \ctl_rf_tc_reg[7]/NET0131  ;
  input \de_bst_cnt_reg[0]/NET0131  ;
  input \de_bst_cnt_reg[2]/NET0131  ;
  input \de_bst_cnt_reg[3]/NET0131  ;
  input \de_bst_cnt_reg[4]/NET0131  ;
  input \de_bst_cnt_reg[5]/NET0131  ;
  input \de_bst_cnt_reg[6]/NET0131  ;
  input \de_bst_cnt_reg[7]/NET0131  ;
  input \de_bst_cnt_reg[8]/NET0131  ;
  input \de_de_st_reg[0]/NET0131  ;
  input \de_de_st_reg[1]/NET0131  ;
  input \de_de_st_reg[2]/NET0131  ;
  input \de_de_st_reg[5]/NET0131  ;
  input \de_de_st_reg[6]/NET0131  ;
  input \de_m0_arb_st_reg/NET0131  ;
  input \de_m0_is_llp_reg/NET0131  ;
  input \de_m1_arb_st_reg[0]/NET0131  ;
  input \de_m1_arb_st_reg[1]/NET0131  ;
  input \de_m1_is_llp_reg/NET0131  ;
  input \de_st_rd_msk_reg/NET0131  ;
  input \de_tsz_cnt_reg[0]/NET0131  ;
  input \de_tsz_cnt_reg[10]/NET0131  ;
  input \de_tsz_cnt_reg[11]/NET0131  ;
  input \de_tsz_cnt_reg[1]/NET0131  ;
  input \de_tsz_cnt_reg[2]/NET0131  ;
  input \de_tsz_cnt_reg[3]/NET0131  ;
  input \de_tsz_cnt_reg[4]/NET0131  ;
  input \de_tsz_cnt_reg[5]/NET0131  ;
  input \de_tsz_cnt_reg[6]/NET0131  ;
  input \de_tsz_cnt_reg[7]/NET0131  ;
  input \de_tsz_cnt_reg[8]/NET0131  ;
  input \de_tsz_cnt_reg[9]/NET0131  ;
  input \dma_ack[0]_pad  ;
  input \dma_ack[1]_pad  ;
  input \dma_ack[2]_pad  ;
  input \dma_ack[3]_pad  ;
  input \dma_ack[4]_pad  ;
  input \dma_ack[5]_pad  ;
  input \dma_ack[6]_pad  ;
  input \dma_ack[7]_pad  ;
  input \dma_tc[0]_pad  ;
  input \dma_tc[1]_pad  ;
  input \dma_tc[2]_pad  ;
  input \dma_tc[3]_pad  ;
  input \dma_tc[4]_pad  ;
  input \dma_tc[5]_pad  ;
  input \dma_tc[6]_pad  ;
  input \dma_tc[7]_pad  ;
  input \h0burst[0]_pad  ;
  input \h0grant_pad  ;
  input \h0readyin_pad  ;
  input \h0req_pad  ;
  input \h0resp[0]_pad  ;
  input \h0resp[1]_pad  ;
  input \h0write_pad  ;
  input \h1burst[0]_pad  ;
  input \h1prot[0]_pad  ;
  input \h1rdt0_br[0]_pad  ;
  input \h1rdt0_br[10]_pad  ;
  input \h1rdt0_br[11]_pad  ;
  input \h1rdt0_br[12]_pad  ;
  input \h1rdt0_br[13]_pad  ;
  input \h1rdt0_br[14]_pad  ;
  input \h1rdt0_br[15]_pad  ;
  input \h1rdt0_br[16]_pad  ;
  input \h1rdt0_br[17]_pad  ;
  input \h1rdt0_br[18]_pad  ;
  input \h1rdt0_br[19]_pad  ;
  input \h1rdt0_br[1]_pad  ;
  input \h1rdt0_br[20]_pad  ;
  input \h1rdt0_br[21]_pad  ;
  input \h1rdt0_br[22]_pad  ;
  input \h1rdt0_br[23]_pad  ;
  input \h1rdt0_br[24]_pad  ;
  input \h1rdt0_br[25]_pad  ;
  input \h1rdt0_br[26]_pad  ;
  input \h1rdt0_br[27]_pad  ;
  input \h1rdt0_br[28]_pad  ;
  input \h1rdt0_br[29]_pad  ;
  input \h1rdt0_br[2]_pad  ;
  input \h1rdt0_br[30]_pad  ;
  input \h1rdt0_br[31]_pad  ;
  input \h1rdt0_br[3]_pad  ;
  input \h1rdt0_br[4]_pad  ;
  input \h1rdt0_br[5]_pad  ;
  input \h1rdt0_br[6]_pad  ;
  input \h1rdt0_br[7]_pad  ;
  input \h1rdt0_br[8]_pad  ;
  input \h1rdt0_br[9]_pad  ;
  input \h1rdt0_dma[0]_pad  ;
  input \h1rdt0_dma[10]_pad  ;
  input \h1rdt0_dma[11]_pad  ;
  input \h1rdt0_dma[12]_pad  ;
  input \h1rdt0_dma[13]_pad  ;
  input \h1rdt0_dma[14]_pad  ;
  input \h1rdt0_dma[15]_pad  ;
  input \h1rdt0_dma[16]_pad  ;
  input \h1rdt0_dma[17]_pad  ;
  input \h1rdt0_dma[18]_pad  ;
  input \h1rdt0_dma[19]_pad  ;
  input \h1rdt0_dma[1]_pad  ;
  input \h1rdt0_dma[20]_pad  ;
  input \h1rdt0_dma[21]_pad  ;
  input \h1rdt0_dma[22]_pad  ;
  input \h1rdt0_dma[23]_pad  ;
  input \h1rdt0_dma[24]_pad  ;
  input \h1rdt0_dma[25]_pad  ;
  input \h1rdt0_dma[26]_pad  ;
  input \h1rdt0_dma[27]_pad  ;
  input \h1rdt0_dma[28]_pad  ;
  input \h1rdt0_dma[29]_pad  ;
  input \h1rdt0_dma[2]_pad  ;
  input \h1rdt0_dma[30]_pad  ;
  input \h1rdt0_dma[31]_pad  ;
  input \h1rdt0_dma[3]_pad  ;
  input \h1rdt0_dma[4]_pad  ;
  input \h1rdt0_dma[5]_pad  ;
  input \h1rdt0_dma[6]_pad  ;
  input \h1rdt0_dma[7]_pad  ;
  input \h1rdt0_dma[8]_pad  ;
  input \h1rdt0_dma[9]_pad  ;
  input \h1rdt1_br[0]_pad  ;
  input \h1rdt1_br[10]_pad  ;
  input \h1rdt1_br[11]_pad  ;
  input \h1rdt1_br[12]_pad  ;
  input \h1rdt1_br[13]_pad  ;
  input \h1rdt1_br[14]_pad  ;
  input \h1rdt1_br[15]_pad  ;
  input \h1rdt1_br[16]_pad  ;
  input \h1rdt1_br[17]_pad  ;
  input \h1rdt1_br[18]_pad  ;
  input \h1rdt1_br[19]_pad  ;
  input \h1rdt1_br[1]_pad  ;
  input \h1rdt1_br[20]_pad  ;
  input \h1rdt1_br[21]_pad  ;
  input \h1rdt1_br[22]_pad  ;
  input \h1rdt1_br[23]_pad  ;
  input \h1rdt1_br[24]_pad  ;
  input \h1rdt1_br[25]_pad  ;
  input \h1rdt1_br[26]_pad  ;
  input \h1rdt1_br[27]_pad  ;
  input \h1rdt1_br[28]_pad  ;
  input \h1rdt1_br[29]_pad  ;
  input \h1rdt1_br[2]_pad  ;
  input \h1rdt1_br[30]_pad  ;
  input \h1rdt1_br[31]_pad  ;
  input \h1rdt1_br[3]_pad  ;
  input \h1rdt1_br[4]_pad  ;
  input \h1rdt1_br[5]_pad  ;
  input \h1rdt1_br[6]_pad  ;
  input \h1rdt1_br[7]_pad  ;
  input \h1rdt1_br[8]_pad  ;
  input \h1rdt1_br[9]_pad  ;
  input \h1rdt1_dma[0]_pad  ;
  input \h1rdt1_dma[10]_pad  ;
  input \h1rdt1_dma[11]_pad  ;
  input \h1rdt1_dma[12]_pad  ;
  input \h1rdt1_dma[13]_pad  ;
  input \h1rdt1_dma[14]_pad  ;
  input \h1rdt1_dma[15]_pad  ;
  input \h1rdt1_dma[16]_pad  ;
  input \h1rdt1_dma[17]_pad  ;
  input \h1rdt1_dma[18]_pad  ;
  input \h1rdt1_dma[19]_pad  ;
  input \h1rdt1_dma[1]_pad  ;
  input \h1rdt1_dma[20]_pad  ;
  input \h1rdt1_dma[21]_pad  ;
  input \h1rdt1_dma[22]_pad  ;
  input \h1rdt1_dma[23]_pad  ;
  input \h1rdt1_dma[24]_pad  ;
  input \h1rdt1_dma[25]_pad  ;
  input \h1rdt1_dma[26]_pad  ;
  input \h1rdt1_dma[27]_pad  ;
  input \h1rdt1_dma[28]_pad  ;
  input \h1rdt1_dma[29]_pad  ;
  input \h1rdt1_dma[2]_pad  ;
  input \h1rdt1_dma[30]_pad  ;
  input \h1rdt1_dma[31]_pad  ;
  input \h1rdt1_dma[3]_pad  ;
  input \h1rdt1_dma[4]_pad  ;
  input \h1rdt1_dma[5]_pad  ;
  input \h1rdt1_dma[6]_pad  ;
  input \h1rdt1_dma[7]_pad  ;
  input \h1rdt1_dma[8]_pad  ;
  input \h1rdt1_dma[9]_pad  ;
  input \h1rdt2_br[0]_pad  ;
  input \h1rdt2_br[10]_pad  ;
  input \h1rdt2_br[11]_pad  ;
  input \h1rdt2_br[12]_pad  ;
  input \h1rdt2_br[13]_pad  ;
  input \h1rdt2_br[14]_pad  ;
  input \h1rdt2_br[15]_pad  ;
  input \h1rdt2_br[16]_pad  ;
  input \h1rdt2_br[17]_pad  ;
  input \h1rdt2_br[18]_pad  ;
  input \h1rdt2_br[19]_pad  ;
  input \h1rdt2_br[1]_pad  ;
  input \h1rdt2_br[20]_pad  ;
  input \h1rdt2_br[21]_pad  ;
  input \h1rdt2_br[22]_pad  ;
  input \h1rdt2_br[23]_pad  ;
  input \h1rdt2_br[24]_pad  ;
  input \h1rdt2_br[25]_pad  ;
  input \h1rdt2_br[26]_pad  ;
  input \h1rdt2_br[27]_pad  ;
  input \h1rdt2_br[28]_pad  ;
  input \h1rdt2_br[29]_pad  ;
  input \h1rdt2_br[2]_pad  ;
  input \h1rdt2_br[30]_pad  ;
  input \h1rdt2_br[31]_pad  ;
  input \h1rdt2_br[3]_pad  ;
  input \h1rdt2_br[4]_pad  ;
  input \h1rdt2_br[5]_pad  ;
  input \h1rdt2_br[6]_pad  ;
  input \h1rdt2_br[7]_pad  ;
  input \h1rdt2_br[8]_pad  ;
  input \h1rdt2_br[9]_pad  ;
  input \h1rdt2_dma[0]_pad  ;
  input \h1rdt2_dma[10]_pad  ;
  input \h1rdt2_dma[11]_pad  ;
  input \h1rdt2_dma[12]_pad  ;
  input \h1rdt2_dma[13]_pad  ;
  input \h1rdt2_dma[14]_pad  ;
  input \h1rdt2_dma[15]_pad  ;
  input \h1rdt2_dma[16]_pad  ;
  input \h1rdt2_dma[17]_pad  ;
  input \h1rdt2_dma[18]_pad  ;
  input \h1rdt2_dma[19]_pad  ;
  input \h1rdt2_dma[1]_pad  ;
  input \h1rdt2_dma[20]_pad  ;
  input \h1rdt2_dma[21]_pad  ;
  input \h1rdt2_dma[22]_pad  ;
  input \h1rdt2_dma[23]_pad  ;
  input \h1rdt2_dma[24]_pad  ;
  input \h1rdt2_dma[25]_pad  ;
  input \h1rdt2_dma[26]_pad  ;
  input \h1rdt2_dma[27]_pad  ;
  input \h1rdt2_dma[28]_pad  ;
  input \h1rdt2_dma[29]_pad  ;
  input \h1rdt2_dma[2]_pad  ;
  input \h1rdt2_dma[30]_pad  ;
  input \h1rdt2_dma[31]_pad  ;
  input \h1rdt2_dma[3]_pad  ;
  input \h1rdt2_dma[4]_pad  ;
  input \h1rdt2_dma[5]_pad  ;
  input \h1rdt2_dma[6]_pad  ;
  input \h1rdt2_dma[7]_pad  ;
  input \h1rdt2_dma[8]_pad  ;
  input \h1rdt2_dma[9]_pad  ;
  input \h1rdt3_br[0]_pad  ;
  input \h1rdt3_br[10]_pad  ;
  input \h1rdt3_br[11]_pad  ;
  input \h1rdt3_br[12]_pad  ;
  input \h1rdt3_br[13]_pad  ;
  input \h1rdt3_br[14]_pad  ;
  input \h1rdt3_br[15]_pad  ;
  input \h1rdt3_br[16]_pad  ;
  input \h1rdt3_br[17]_pad  ;
  input \h1rdt3_br[18]_pad  ;
  input \h1rdt3_br[19]_pad  ;
  input \h1rdt3_br[1]_pad  ;
  input \h1rdt3_br[20]_pad  ;
  input \h1rdt3_br[21]_pad  ;
  input \h1rdt3_br[22]_pad  ;
  input \h1rdt3_br[23]_pad  ;
  input \h1rdt3_br[24]_pad  ;
  input \h1rdt3_br[25]_pad  ;
  input \h1rdt3_br[26]_pad  ;
  input \h1rdt3_br[27]_pad  ;
  input \h1rdt3_br[28]_pad  ;
  input \h1rdt3_br[29]_pad  ;
  input \h1rdt3_br[2]_pad  ;
  input \h1rdt3_br[30]_pad  ;
  input \h1rdt3_br[31]_pad  ;
  input \h1rdt3_br[3]_pad  ;
  input \h1rdt3_br[4]_pad  ;
  input \h1rdt3_br[5]_pad  ;
  input \h1rdt3_br[6]_pad  ;
  input \h1rdt3_br[7]_pad  ;
  input \h1rdt3_br[8]_pad  ;
  input \h1rdt3_br[9]_pad  ;
  input \h1rdt3_dma[0]_pad  ;
  input \h1rdt3_dma[10]_pad  ;
  input \h1rdt3_dma[11]_pad  ;
  input \h1rdt3_dma[12]_pad  ;
  input \h1rdt3_dma[13]_pad  ;
  input \h1rdt3_dma[14]_pad  ;
  input \h1rdt3_dma[15]_pad  ;
  input \h1rdt3_dma[16]_pad  ;
  input \h1rdt3_dma[17]_pad  ;
  input \h1rdt3_dma[18]_pad  ;
  input \h1rdt3_dma[19]_pad  ;
  input \h1rdt3_dma[1]_pad  ;
  input \h1rdt3_dma[20]_pad  ;
  input \h1rdt3_dma[21]_pad  ;
  input \h1rdt3_dma[22]_pad  ;
  input \h1rdt3_dma[23]_pad  ;
  input \h1rdt3_dma[24]_pad  ;
  input \h1rdt3_dma[25]_pad  ;
  input \h1rdt3_dma[26]_pad  ;
  input \h1rdt3_dma[27]_pad  ;
  input \h1rdt3_dma[28]_pad  ;
  input \h1rdt3_dma[29]_pad  ;
  input \h1rdt3_dma[2]_pad  ;
  input \h1rdt3_dma[30]_pad  ;
  input \h1rdt3_dma[31]_pad  ;
  input \h1rdt3_dma[3]_pad  ;
  input \h1rdt3_dma[4]_pad  ;
  input \h1rdt3_dma[5]_pad  ;
  input \h1rdt3_dma[6]_pad  ;
  input \h1rdt3_dma[7]_pad  ;
  input \h1rdt3_dma[8]_pad  ;
  input \h1rdt3_dma[9]_pad  ;
  input \h1rdt4_br[0]_pad  ;
  input \h1rdt4_br[10]_pad  ;
  input \h1rdt4_br[11]_pad  ;
  input \h1rdt4_br[12]_pad  ;
  input \h1rdt4_br[13]_pad  ;
  input \h1rdt4_br[14]_pad  ;
  input \h1rdt4_br[15]_pad  ;
  input \h1rdt4_br[16]_pad  ;
  input \h1rdt4_br[17]_pad  ;
  input \h1rdt4_br[18]_pad  ;
  input \h1rdt4_br[19]_pad  ;
  input \h1rdt4_br[1]_pad  ;
  input \h1rdt4_br[20]_pad  ;
  input \h1rdt4_br[21]_pad  ;
  input \h1rdt4_br[22]_pad  ;
  input \h1rdt4_br[23]_pad  ;
  input \h1rdt4_br[24]_pad  ;
  input \h1rdt4_br[25]_pad  ;
  input \h1rdt4_br[26]_pad  ;
  input \h1rdt4_br[27]_pad  ;
  input \h1rdt4_br[28]_pad  ;
  input \h1rdt4_br[29]_pad  ;
  input \h1rdt4_br[2]_pad  ;
  input \h1rdt4_br[30]_pad  ;
  input \h1rdt4_br[31]_pad  ;
  input \h1rdt4_br[3]_pad  ;
  input \h1rdt4_br[4]_pad  ;
  input \h1rdt4_br[5]_pad  ;
  input \h1rdt4_br[6]_pad  ;
  input \h1rdt4_br[7]_pad  ;
  input \h1rdt4_br[8]_pad  ;
  input \h1rdt4_br[9]_pad  ;
  input \h1rdt4_dma[0]_pad  ;
  input \h1rdt4_dma[10]_pad  ;
  input \h1rdt4_dma[11]_pad  ;
  input \h1rdt4_dma[12]_pad  ;
  input \h1rdt4_dma[13]_pad  ;
  input \h1rdt4_dma[14]_pad  ;
  input \h1rdt4_dma[15]_pad  ;
  input \h1rdt4_dma[16]_pad  ;
  input \h1rdt4_dma[17]_pad  ;
  input \h1rdt4_dma[18]_pad  ;
  input \h1rdt4_dma[19]_pad  ;
  input \h1rdt4_dma[1]_pad  ;
  input \h1rdt4_dma[20]_pad  ;
  input \h1rdt4_dma[21]_pad  ;
  input \h1rdt4_dma[22]_pad  ;
  input \h1rdt4_dma[23]_pad  ;
  input \h1rdt4_dma[24]_pad  ;
  input \h1rdt4_dma[25]_pad  ;
  input \h1rdt4_dma[26]_pad  ;
  input \h1rdt4_dma[27]_pad  ;
  input \h1rdt4_dma[28]_pad  ;
  input \h1rdt4_dma[29]_pad  ;
  input \h1rdt4_dma[2]_pad  ;
  input \h1rdt4_dma[30]_pad  ;
  input \h1rdt4_dma[31]_pad  ;
  input \h1rdt4_dma[3]_pad  ;
  input \h1rdt4_dma[4]_pad  ;
  input \h1rdt4_dma[5]_pad  ;
  input \h1rdt4_dma[6]_pad  ;
  input \h1rdt4_dma[7]_pad  ;
  input \h1rdt4_dma[8]_pad  ;
  input \h1rdt4_dma[9]_pad  ;
  input \h1rdt5_br[0]_pad  ;
  input \h1rdt5_br[10]_pad  ;
  input \h1rdt5_br[11]_pad  ;
  input \h1rdt5_br[12]_pad  ;
  input \h1rdt5_br[13]_pad  ;
  input \h1rdt5_br[14]_pad  ;
  input \h1rdt5_br[15]_pad  ;
  input \h1rdt5_br[16]_pad  ;
  input \h1rdt5_br[17]_pad  ;
  input \h1rdt5_br[18]_pad  ;
  input \h1rdt5_br[19]_pad  ;
  input \h1rdt5_br[1]_pad  ;
  input \h1rdt5_br[20]_pad  ;
  input \h1rdt5_br[21]_pad  ;
  input \h1rdt5_br[22]_pad  ;
  input \h1rdt5_br[23]_pad  ;
  input \h1rdt5_br[24]_pad  ;
  input \h1rdt5_br[25]_pad  ;
  input \h1rdt5_br[26]_pad  ;
  input \h1rdt5_br[27]_pad  ;
  input \h1rdt5_br[28]_pad  ;
  input \h1rdt5_br[29]_pad  ;
  input \h1rdt5_br[2]_pad  ;
  input \h1rdt5_br[30]_pad  ;
  input \h1rdt5_br[31]_pad  ;
  input \h1rdt5_br[3]_pad  ;
  input \h1rdt5_br[4]_pad  ;
  input \h1rdt5_br[5]_pad  ;
  input \h1rdt5_br[6]_pad  ;
  input \h1rdt5_br[7]_pad  ;
  input \h1rdt5_br[8]_pad  ;
  input \h1rdt5_br[9]_pad  ;
  input \h1rdt5_dma[0]_pad  ;
  input \h1rdt5_dma[10]_pad  ;
  input \h1rdt5_dma[11]_pad  ;
  input \h1rdt5_dma[12]_pad  ;
  input \h1rdt5_dma[13]_pad  ;
  input \h1rdt5_dma[14]_pad  ;
  input \h1rdt5_dma[15]_pad  ;
  input \h1rdt5_dma[16]_pad  ;
  input \h1rdt5_dma[17]_pad  ;
  input \h1rdt5_dma[18]_pad  ;
  input \h1rdt5_dma[19]_pad  ;
  input \h1rdt5_dma[1]_pad  ;
  input \h1rdt5_dma[20]_pad  ;
  input \h1rdt5_dma[21]_pad  ;
  input \h1rdt5_dma[22]_pad  ;
  input \h1rdt5_dma[23]_pad  ;
  input \h1rdt5_dma[24]_pad  ;
  input \h1rdt5_dma[25]_pad  ;
  input \h1rdt5_dma[26]_pad  ;
  input \h1rdt5_dma[27]_pad  ;
  input \h1rdt5_dma[28]_pad  ;
  input \h1rdt5_dma[29]_pad  ;
  input \h1rdt5_dma[2]_pad  ;
  input \h1rdt5_dma[30]_pad  ;
  input \h1rdt5_dma[31]_pad  ;
  input \h1rdt5_dma[3]_pad  ;
  input \h1rdt5_dma[4]_pad  ;
  input \h1rdt5_dma[5]_pad  ;
  input \h1rdt5_dma[6]_pad  ;
  input \h1rdt5_dma[7]_pad  ;
  input \h1rdt5_dma[8]_pad  ;
  input \h1rdt5_dma[9]_pad  ;
  input \h1rdt6_br[0]_pad  ;
  input \h1rdt6_br[10]_pad  ;
  input \h1rdt6_br[11]_pad  ;
  input \h1rdt6_br[12]_pad  ;
  input \h1rdt6_br[13]_pad  ;
  input \h1rdt6_br[14]_pad  ;
  input \h1rdt6_br[15]_pad  ;
  input \h1rdt6_br[16]_pad  ;
  input \h1rdt6_br[17]_pad  ;
  input \h1rdt6_br[18]_pad  ;
  input \h1rdt6_br[19]_pad  ;
  input \h1rdt6_br[1]_pad  ;
  input \h1rdt6_br[20]_pad  ;
  input \h1rdt6_br[21]_pad  ;
  input \h1rdt6_br[22]_pad  ;
  input \h1rdt6_br[23]_pad  ;
  input \h1rdt6_br[24]_pad  ;
  input \h1rdt6_br[25]_pad  ;
  input \h1rdt6_br[26]_pad  ;
  input \h1rdt6_br[27]_pad  ;
  input \h1rdt6_br[28]_pad  ;
  input \h1rdt6_br[29]_pad  ;
  input \h1rdt6_br[2]_pad  ;
  input \h1rdt6_br[30]_pad  ;
  input \h1rdt6_br[31]_pad  ;
  input \h1rdt6_br[3]_pad  ;
  input \h1rdt6_br[4]_pad  ;
  input \h1rdt6_br[5]_pad  ;
  input \h1rdt6_br[6]_pad  ;
  input \h1rdt6_br[7]_pad  ;
  input \h1rdt6_br[8]_pad  ;
  input \h1rdt6_br[9]_pad  ;
  input \h1rdt6_dma[0]_pad  ;
  input \h1rdt6_dma[10]_pad  ;
  input \h1rdt6_dma[11]_pad  ;
  input \h1rdt6_dma[12]_pad  ;
  input \h1rdt6_dma[13]_pad  ;
  input \h1rdt6_dma[14]_pad  ;
  input \h1rdt6_dma[15]_pad  ;
  input \h1rdt6_dma[16]_pad  ;
  input \h1rdt6_dma[17]_pad  ;
  input \h1rdt6_dma[18]_pad  ;
  input \h1rdt6_dma[19]_pad  ;
  input \h1rdt6_dma[1]_pad  ;
  input \h1rdt6_dma[20]_pad  ;
  input \h1rdt6_dma[21]_pad  ;
  input \h1rdt6_dma[22]_pad  ;
  input \h1rdt6_dma[23]_pad  ;
  input \h1rdt6_dma[24]_pad  ;
  input \h1rdt6_dma[25]_pad  ;
  input \h1rdt6_dma[26]_pad  ;
  input \h1rdt6_dma[27]_pad  ;
  input \h1rdt6_dma[28]_pad  ;
  input \h1rdt6_dma[29]_pad  ;
  input \h1rdt6_dma[2]_pad  ;
  input \h1rdt6_dma[30]_pad  ;
  input \h1rdt6_dma[31]_pad  ;
  input \h1rdt6_dma[3]_pad  ;
  input \h1rdt6_dma[4]_pad  ;
  input \h1rdt6_dma[5]_pad  ;
  input \h1rdt6_dma[6]_pad  ;
  input \h1rdt6_dma[7]_pad  ;
  input \h1rdt6_dma[8]_pad  ;
  input \h1rdt6_dma[9]_pad  ;
  input \h1rdt7_br[0]_pad  ;
  input \h1rdt7_br[10]_pad  ;
  input \h1rdt7_br[11]_pad  ;
  input \h1rdt7_br[12]_pad  ;
  input \h1rdt7_br[13]_pad  ;
  input \h1rdt7_br[14]_pad  ;
  input \h1rdt7_br[15]_pad  ;
  input \h1rdt7_br[16]_pad  ;
  input \h1rdt7_br[17]_pad  ;
  input \h1rdt7_br[18]_pad  ;
  input \h1rdt7_br[19]_pad  ;
  input \h1rdt7_br[1]_pad  ;
  input \h1rdt7_br[20]_pad  ;
  input \h1rdt7_br[21]_pad  ;
  input \h1rdt7_br[22]_pad  ;
  input \h1rdt7_br[23]_pad  ;
  input \h1rdt7_br[24]_pad  ;
  input \h1rdt7_br[25]_pad  ;
  input \h1rdt7_br[26]_pad  ;
  input \h1rdt7_br[27]_pad  ;
  input \h1rdt7_br[28]_pad  ;
  input \h1rdt7_br[29]_pad  ;
  input \h1rdt7_br[2]_pad  ;
  input \h1rdt7_br[30]_pad  ;
  input \h1rdt7_br[31]_pad  ;
  input \h1rdt7_br[3]_pad  ;
  input \h1rdt7_br[4]_pad  ;
  input \h1rdt7_br[5]_pad  ;
  input \h1rdt7_br[6]_pad  ;
  input \h1rdt7_br[7]_pad  ;
  input \h1rdt7_br[8]_pad  ;
  input \h1rdt7_br[9]_pad  ;
  input \h1rdt7_dma[0]_pad  ;
  input \h1rdt7_dma[10]_pad  ;
  input \h1rdt7_dma[11]_pad  ;
  input \h1rdt7_dma[12]_pad  ;
  input \h1rdt7_dma[13]_pad  ;
  input \h1rdt7_dma[14]_pad  ;
  input \h1rdt7_dma[15]_pad  ;
  input \h1rdt7_dma[16]_pad  ;
  input \h1rdt7_dma[17]_pad  ;
  input \h1rdt7_dma[18]_pad  ;
  input \h1rdt7_dma[19]_pad  ;
  input \h1rdt7_dma[1]_pad  ;
  input \h1rdt7_dma[20]_pad  ;
  input \h1rdt7_dma[21]_pad  ;
  input \h1rdt7_dma[22]_pad  ;
  input \h1rdt7_dma[23]_pad  ;
  input \h1rdt7_dma[24]_pad  ;
  input \h1rdt7_dma[25]_pad  ;
  input \h1rdt7_dma[26]_pad  ;
  input \h1rdt7_dma[27]_pad  ;
  input \h1rdt7_dma[28]_pad  ;
  input \h1rdt7_dma[29]_pad  ;
  input \h1rdt7_dma[2]_pad  ;
  input \h1rdt7_dma[30]_pad  ;
  input \h1rdt7_dma[31]_pad  ;
  input \h1rdt7_dma[3]_pad  ;
  input \h1rdt7_dma[4]_pad  ;
  input \h1rdt7_dma[5]_pad  ;
  input \h1rdt7_dma[6]_pad  ;
  input \h1rdt7_dma[7]_pad  ;
  input \h1rdt7_dma[8]_pad  ;
  input \h1rdt7_dma[9]_pad  ;
  input \h1rdy0_br_pad  ;
  input \h1rdy0_dma_pad  ;
  input \h1rdy1_br_pad  ;
  input \h1rdy1_dma_pad  ;
  input \h1rdy2_br_pad  ;
  input \h1rdy2_dma_pad  ;
  input \h1rdy3_br_pad  ;
  input \h1rdy3_dma_pad  ;
  input \h1rdy4_br_pad  ;
  input \h1rdy4_dma_pad  ;
  input \h1rdy5_br_pad  ;
  input \h1rdy5_dma_pad  ;
  input \h1rdy6_br_pad  ;
  input \h1rdy6_dma_pad  ;
  input \h1rdy7_br_pad  ;
  input \h1rdy7_dma_pad  ;
  input \h1rp0_br[0]_pad  ;
  input \h1rp0_br[1]_pad  ;
  input \h1rp0_dma[0]_pad  ;
  input \h1rp0_dma[1]_pad  ;
  input \h1rp1_br[0]_pad  ;
  input \h1rp1_br[1]_pad  ;
  input \h1rp1_dma[0]_pad  ;
  input \h1rp1_dma[1]_pad  ;
  input \h1rp2_br[0]_pad  ;
  input \h1rp2_br[1]_pad  ;
  input \h1rp2_dma[0]_pad  ;
  input \h1rp2_dma[1]_pad  ;
  input \h1rp3_br[0]_pad  ;
  input \h1rp3_br[1]_pad  ;
  input \h1rp3_dma[0]_pad  ;
  input \h1rp3_dma[1]_pad  ;
  input \h1rp4_br[0]_pad  ;
  input \h1rp4_br[1]_pad  ;
  input \h1rp4_dma[0]_pad  ;
  input \h1rp4_dma[1]_pad  ;
  input \h1rp5_br[0]_pad  ;
  input \h1rp5_br[1]_pad  ;
  input \h1rp5_dma[0]_pad  ;
  input \h1rp5_dma[1]_pad  ;
  input \h1rp6_br[0]_pad  ;
  input \h1rp6_br[1]_pad  ;
  input \h1rp6_dma[0]_pad  ;
  input \h1rp6_dma[1]_pad  ;
  input \h1rp7_br[0]_pad  ;
  input \h1rp7_br[1]_pad  ;
  input \h1rp7_dma[0]_pad  ;
  input \h1rp7_dma[1]_pad  ;
  input \h1size[0]_pad  ;
  input \h1size[1]_pad  ;
  input \h1size[2]_pad  ;
  input \h1write_pad  ;
  input \haddr[0]_pad  ;
  input \haddr[1]_pad  ;
  input \haddr[2]_pad  ;
  input \haddr[3]_pad  ;
  input \haddr[4]_pad  ;
  input \haddr[5]_pad  ;
  input \haddr[6]_pad  ;
  input \haddr[7]_pad  ;
  input \haddr[8]_pad  ;
  input \hrdata_reg[0]_pad  ;
  input \hrdata_reg[10]_pad  ;
  input \hrdata_reg[11]_pad  ;
  input \hrdata_reg[12]_pad  ;
  input \hrdata_reg[13]_pad  ;
  input \hrdata_reg[14]_pad  ;
  input \hrdata_reg[15]_pad  ;
  input \hrdata_reg[16]_pad  ;
  input \hrdata_reg[17]_pad  ;
  input \hrdata_reg[18]_pad  ;
  input \hrdata_reg[19]_pad  ;
  input \hrdata_reg[1]_pad  ;
  input \hrdata_reg[20]_pad  ;
  input \hrdata_reg[21]_pad  ;
  input \hrdata_reg[22]_pad  ;
  input \hrdata_reg[23]_pad  ;
  input \hrdata_reg[24]_pad  ;
  input \hrdata_reg[25]_pad  ;
  input \hrdata_reg[26]_pad  ;
  input \hrdata_reg[27]_pad  ;
  input \hrdata_reg[28]_pad  ;
  input \hrdata_reg[29]_pad  ;
  input \hrdata_reg[2]_pad  ;
  input \hrdata_reg[30]_pad  ;
  input \hrdata_reg[31]_pad  ;
  input \hrdata_reg[3]_pad  ;
  input \hrdata_reg[4]_pad  ;
  input \hrdata_reg[5]_pad  ;
  input \hrdata_reg[6]_pad  ;
  input \hrdata_reg[7]_pad  ;
  input \hrdata_reg[8]_pad  ;
  input \hrdata_reg[9]_pad  ;
  input hreadyin_pad ;
  input hreadyout_br_pad ;
  input \hresp_br[0]_pad  ;
  input \hresp_br[1]_pad  ;
  input hsel_br_pad ;
  input hsel_reg_pad ;
  input \hsize[0]_pad  ;
  input \hsize[1]_pad  ;
  input \hsize[2]_pad  ;
  input \htrans[0]_pad  ;
  input \htrans[1]_pad  ;
  input \hwdata[0]_pad  ;
  input \hwdata[10]_pad  ;
  input \hwdata[11]_pad  ;
  input \hwdata[12]_pad  ;
  input \hwdata[13]_pad  ;
  input \hwdata[14]_pad  ;
  input \hwdata[15]_pad  ;
  input \hwdata[16]_pad  ;
  input \hwdata[17]_pad  ;
  input \hwdata[18]_pad  ;
  input \hwdata[19]_pad  ;
  input \hwdata[1]_pad  ;
  input \hwdata[20]_pad  ;
  input \hwdata[21]_pad  ;
  input \hwdata[22]_pad  ;
  input \hwdata[23]_pad  ;
  input \hwdata[24]_pad  ;
  input \hwdata[25]_pad  ;
  input \hwdata[26]_pad  ;
  input \hwdata[27]_pad  ;
  input \hwdata[28]_pad  ;
  input \hwdata[29]_pad  ;
  input \hwdata[2]_pad  ;
  input \hwdata[30]_pad  ;
  input \hwdata[31]_pad  ;
  input \hwdata[3]_pad  ;
  input \hwdata[4]_pad  ;
  input \hwdata[5]_pad  ;
  input \hwdata[6]_pad  ;
  input \hwdata[7]_pad  ;
  input \hwdata[8]_pad  ;
  input \hwdata[9]_pad  ;
  input hwrite_pad ;
  input \m1_mux_hrdy_df_reg/NET0131  ;
  input \m1_mux_hrmxnof_reg/NET0131  ;
  input \m1_mux_hrp_df_reg[0]/NET0131  ;
  input \m1_mux_mux_no_reg[0]/NET0131  ;
  input \m1_mux_mux_no_reg[1]/NET0131  ;
  input \m1_mux_mux_no_reg[2]/NET0131  ;
  input \m1_mux_mux_no_reg[3]/NET0131  ;
  output \_al_n1  ;
  output \g16/_0_  ;
  output \g58487/_0_  ;
  output \g58489/_0_  ;
  output \g58491/_0_  ;
  output \g58493/_0_  ;
  output \g58495/_0_  ;
  output \g58497/_0_  ;
  output \g58499/_0_  ;
  output \g58500/_0_  ;
  output \g58501/_0_  ;
  output \g58502/_0_  ;
  output \g58504/_0_  ;
  output \g58505/_0_  ;
  output \g58507/_0_  ;
  output \g58508/_0_  ;
  output \g58509/_0_  ;
  output \g58510/_0_  ;
  output \g58556/_0_  ;
  output \g58557/_0_  ;
  output \g58558/_0_  ;
  output \g58559/_0_  ;
  output \g58560/_0_  ;
  output \g58561/_0_  ;
  output \g58562/_0_  ;
  output \g58563/_0_  ;
  output \g58566/_0_  ;
  output \g58567/_0_  ;
  output \g58568/_0_  ;
  output \g58569/_0_  ;
  output \g58570/_0_  ;
  output \g58571/_0_  ;
  output \g58572/_0_  ;
  output \g58573/_0_  ;
  output \g58574/_0_  ;
  output \g58575/_0_  ;
  output \g58576/_0_  ;
  output \g58577/_0_  ;
  output \g58578/_0_  ;
  output \g58579/_0_  ;
  output \g58580/_0_  ;
  output \g58581/_0_  ;
  output \g58584/_0_  ;
  output \g58585/_0_  ;
  output \g58586/_0_  ;
  output \g58587/_0_  ;
  output \g58588/_0_  ;
  output \g58589/_0_  ;
  output \g58590/_0_  ;
  output \g58591/_0_  ;
  output \g58592/_0_  ;
  output \g58593/_0_  ;
  output \g58594/_0_  ;
  output \g58595/_0_  ;
  output \g58596/_0_  ;
  output \g58597/_0_  ;
  output \g58598/_0_  ;
  output \g58599/_0_  ;
  output \g58600/_0_  ;
  output \g58601/_0_  ;
  output \g58602/_0_  ;
  output \g58603/_0_  ;
  output \g58604/_0_  ;
  output \g58605/_0_  ;
  output \g58606/_0_  ;
  output \g58607/_0_  ;
  output \g58608/_0_  ;
  output \g58609/_0_  ;
  output \g58610/_0_  ;
  output \g58611/_0_  ;
  output \g58612/_0_  ;
  output \g58613/_0_  ;
  output \g58614/_0_  ;
  output \g58615/_0_  ;
  output \g58616/_0_  ;
  output \g58617/_0_  ;
  output \g58618/_0_  ;
  output \g58619/_0_  ;
  output \g58620/_0_  ;
  output \g58621/_0_  ;
  output \g58622/_0_  ;
  output \g58623/_0_  ;
  output \g58624/_0_  ;
  output \g58625/_0_  ;
  output \g58626/_0_  ;
  output \g58627/_0_  ;
  output \g58723/_0_  ;
  output \g58734/_0_  ;
  output \g58737/_0_  ;
  output \g58741/_0_  ;
  output \g58749/_0_  ;
  output \g58754/_0_  ;
  output \g58762/_0_  ;
  output \g58763/_0_  ;
  output \g58764/_0_  ;
  output \g58765/_0_  ;
  output \g58766/_0_  ;
  output \g58767/_0_  ;
  output \g58768/_0_  ;
  output \g58769/_0_  ;
  output \g58770/_0_  ;
  output \g58771/_0_  ;
  output \g59788/_0_  ;
  output \g59832/_0_  ;
  output \g59873/_0_  ;
  output \g59874/_0_  ;
  output \g59893/_0_  ;
  output \g59894/_0_  ;
  output \g59895/_0_  ;
  output \g59896/_0_  ;
  output \g59923/_0_  ;
  output \g60031/_0_  ;
  output \g60032/_0_  ;
  output \g60033/_0_  ;
  output \g60036/_0_  ;
  output \g60037/_0_  ;
  output \g60038/_0_  ;
  output \g60165/_0_  ;
  output \g60186/_2__syn_2  ;
  output \g60187/_0_  ;
  output \g60188/_0_  ;
  output \g60258/_0_  ;
  output \g60259/_0_  ;
  output \g60260/_0_  ;
  output \g60261/_0_  ;
  output \g60263/_0_  ;
  output \g60264/_0_  ;
  output \g60265/_0_  ;
  output \g60266/_0_  ;
  output \g60267/_0_  ;
  output \g60303/_3_  ;
  output \g60360/_0_  ;
  output \g60361/_0_  ;
  output \g60401/_00_  ;
  output \g60428/_0_  ;
  output \g60429/_0_  ;
  output \g60448/_0_  ;
  output \g60449/_0_  ;
  output \g60974/_0_  ;
  output \g61072/_0_  ;
  output \g61073/_0_  ;
  output \g61074/_0_  ;
  output \g61075/_0_  ;
  output \g61076/_0_  ;
  output \g61077/_0_  ;
  output \g61078/_0_  ;
  output \g61079/_0_  ;
  output \g61486/_0_  ;
  output \g61502/_3_  ;
  output \g61879/_0_  ;
  output \g62077/_0_  ;
  output \g62078/_0_  ;
  output \g62079/_0_  ;
  output \g62080/_0_  ;
  output \g62081/_0_  ;
  output \g62082/_0_  ;
  output \g62083/_0_  ;
  output \g62084/_0_  ;
  output \g62085/_0_  ;
  output \g62086/_0_  ;
  output \g62087/_0_  ;
  output \g62088/_0_  ;
  output \g62089/_0_  ;
  output \g62090/_0_  ;
  output \g62091/_0_  ;
  output \g62629/_0_  ;
  output \g62630/_0_  ;
  output \g62631/_0_  ;
  output \g62632/_0_  ;
  output \g62633/_0_  ;
  output \g62634/_0_  ;
  output \g62635/_0_  ;
  output \g62637/_0_  ;
  output \g62638/_0_  ;
  output \g62639/_0_  ;
  output \g62641/_0_  ;
  output \g62643/_0_  ;
  output \g62645/_0_  ;
  output \g62646/_0_  ;
  output \g62647/_0_  ;
  output \g62648/_0_  ;
  output \g62649/_0_  ;
  output \g62650/_0_  ;
  output \g62651/_0_  ;
  output \g62652/_0_  ;
  output \g62655/_0_  ;
  output \g62656/_0_  ;
  output \g62657/_0_  ;
  output \g62658/_0_  ;
  output \g62659/_0_  ;
  output \g62660/_0_  ;
  output \g62661/_0_  ;
  output \g62662/_0_  ;
  output \g62663/_0_  ;
  output \g62664/_0_  ;
  output \g62665/_0_  ;
  output \g62667/_0_  ;
  output \g62668/_0_  ;
  output \g62669/_0_  ;
  output \g62670/_0_  ;
  output \g62671/_0_  ;
  output \g62672/_0_  ;
  output \g62673/_0_  ;
  output \g62674/_0_  ;
  output \g62675/_0_  ;
  output \g62676/_0_  ;
  output \g62677/_0_  ;
  output \g62678/_0_  ;
  output \g62679/_0_  ;
  output \g62680/_0_  ;
  output \g62681/_0_  ;
  output \g62682/_0_  ;
  output \g62683/_0_  ;
  output \g62684/_0_  ;
  output \g62685/_0_  ;
  output \g62686/_0_  ;
  output \g62687/_0_  ;
  output \g62688/_0_  ;
  output \g62689/_0_  ;
  output \g62690/_0_  ;
  output \g62691/_0_  ;
  output \g62692/_0_  ;
  output \g62693/_0_  ;
  output \g62694/_0_  ;
  output \g62695/_0_  ;
  output \g62696/_0_  ;
  output \g62697/_0_  ;
  output \g62698/_0_  ;
  output \g62699/_0_  ;
  output \g62700/_0_  ;
  output \g62701/_0_  ;
  output \g62702/_0_  ;
  output \g62703/_0_  ;
  output \g62704/_0_  ;
  output \g62705/_0_  ;
  output \g62706/_0_  ;
  output \g62707/_0_  ;
  output \g62708/_0_  ;
  output \g62709/_0_  ;
  output \g62710/_0_  ;
  output \g62711/_0_  ;
  output \g62712/_0_  ;
  output \g62713/_0_  ;
  output \g62714/_0_  ;
  output \g62715/_0_  ;
  output \g62716/_0_  ;
  output \g62721/_0_  ;
  output \g62722/_0_  ;
  output \g62723/_0_  ;
  output \g62725/_0_  ;
  output \g62726/_0_  ;
  output \g62727/_0_  ;
  output \g62728/_0_  ;
  output \g62729/_0_  ;
  output \g62730/_0_  ;
  output \g62731/_0_  ;
  output \g62732/_0_  ;
  output \g62733/_0_  ;
  output \g62734/_0_  ;
  output \g62735/_0_  ;
  output \g62736/_0_  ;
  output \g62737/_0_  ;
  output \g62738/_0_  ;
  output \g62739/_0_  ;
  output \g62740/_0_  ;
  output \g62741/_0_  ;
  output \g62742/_0_  ;
  output \g62743/_0_  ;
  output \g62744/_0_  ;
  output \g62745/_0_  ;
  output \g62746/_0_  ;
  output \g62747/_0_  ;
  output \g62748/_0_  ;
  output \g62749/_0_  ;
  output \g62750/_0_  ;
  output \g62751/_0_  ;
  output \g62752/_0_  ;
  output \g62753/_0_  ;
  output \g62754/_0_  ;
  output \g62755/_0_  ;
  output \g62756/_0_  ;
  output \g62757/_0_  ;
  output \g62758/_0_  ;
  output \g62759/_0_  ;
  output \g62760/_0_  ;
  output \g62761/_0_  ;
  output \g62762/_0_  ;
  output \g62763/_0_  ;
  output \g62764/_0_  ;
  output \g62765/_0_  ;
  output \g62766/_0_  ;
  output \g62767/_0_  ;
  output \g62768/_0_  ;
  output \g62769/_0_  ;
  output \g62770/_0_  ;
  output \g62771/_0_  ;
  output \g62772/_0_  ;
  output \g62773/_0_  ;
  output \g62774/_0_  ;
  output \g62775/_0_  ;
  output \g62776/_0_  ;
  output \g62777/_0_  ;
  output \g62778/_0_  ;
  output \g62779/_0_  ;
  output \g62780/_0_  ;
  output \g62781/_0_  ;
  output \g62783/_0_  ;
  output \g62784/_0_  ;
  output \g62785/_0_  ;
  output \g62786/_0_  ;
  output \g62787/_0_  ;
  output \g62788/_0_  ;
  output \g62789/_0_  ;
  output \g62790/_0_  ;
  output \g62791/_0_  ;
  output \g62792/_0_  ;
  output \g62793/_0_  ;
  output \g62794/_0_  ;
  output \g62795/_0_  ;
  output \g62797/_0_  ;
  output \g62798/_0_  ;
  output \g62799/_0_  ;
  output \g62800/_0_  ;
  output \g62801/_0_  ;
  output \g62802/_0_  ;
  output \g62803/_0_  ;
  output \g62804/_0_  ;
  output \g62805/_0_  ;
  output \g62806/_0_  ;
  output \g62807/_0_  ;
  output \g62808/_0_  ;
  output \g62809/_0_  ;
  output \g62810/_0_  ;
  output \g62811/_0_  ;
  output \g62812/_0_  ;
  output \g62813/_0_  ;
  output \g62814/_0_  ;
  output \g62815/_0_  ;
  output \g62816/_0_  ;
  output \g62817/_0_  ;
  output \g62818/_0_  ;
  output \g63108/_0_  ;
  output \g63117/_0_  ;
  output \g63125/_0_  ;
  output \g63126/_0_  ;
  output \g63127/_0_  ;
  output \g63128/_0_  ;
  output \g63129/_0_  ;
  output \g63130/_0_  ;
  output \g63131/_0_  ;
  output \g63132/_0_  ;
  output \g63133/_0_  ;
  output \g63134/_0_  ;
  output \g63135/_0_  ;
  output \g63136/_0_  ;
  output \g63137/_0_  ;
  output \g63138/_0_  ;
  output \g63139/_0_  ;
  output \g63140/_0_  ;
  output \g63141/_0_  ;
  output \g63142/_0_  ;
  output \g63143/_0_  ;
  output \g63144/_0_  ;
  output \g63145/_0_  ;
  output \g63146/_0_  ;
  output \g63147/_0_  ;
  output \g63148/_0_  ;
  output \g63149/_0_  ;
  output \g63150/_0_  ;
  output \g63151/_0_  ;
  output \g63152/_0_  ;
  output \g63153/_0_  ;
  output \g63154/_0_  ;
  output \g63155/_0_  ;
  output \g63156/_0_  ;
  output \g63157/_0_  ;
  output \g63159/_0_  ;
  output \g63160/_0_  ;
  output \g63161/_0_  ;
  output \g63162/_0_  ;
  output \g63163/_0_  ;
  output \g63164/_0_  ;
  output \g63165/_0_  ;
  output \g63166/_0_  ;
  output \g63167/_0_  ;
  output \g63168/_0_  ;
  output \g63169/_0_  ;
  output \g63170/_0_  ;
  output \g63171/_0_  ;
  output \g63172/_0_  ;
  output \g63173/_0_  ;
  output \g63174/_0_  ;
  output \g63175/_0_  ;
  output \g63176/_0_  ;
  output \g63177/_0_  ;
  output \g63178/_0_  ;
  output \g63179/_0_  ;
  output \g63180/_0_  ;
  output \g63181/_0_  ;
  output \g63182/_0_  ;
  output \g63183/_0_  ;
  output \g63184/_0_  ;
  output \g63185/_0_  ;
  output \g63186/_0_  ;
  output \g63187/_0_  ;
  output \g63188/_0_  ;
  output \g63189/_0_  ;
  output \g63190/_0_  ;
  output \g63191/_0_  ;
  output \g63192/_0_  ;
  output \g63193/_0_  ;
  output \g63194/_0_  ;
  output \g63195/_0_  ;
  output \g63196/_0_  ;
  output \g63197/_0_  ;
  output \g63198/_0_  ;
  output \g63199/_0_  ;
  output \g63200/_0_  ;
  output \g63201/_0_  ;
  output \g63202/_0_  ;
  output \g63203/_0_  ;
  output \g63204/_0_  ;
  output \g63205/_0_  ;
  output \g63206/_0_  ;
  output \g63207/_0_  ;
  output \g63208/_0_  ;
  output \g63209/_0_  ;
  output \g63210/_0_  ;
  output \g63211/_0_  ;
  output \g63212/_0_  ;
  output \g63213/_0_  ;
  output \g63214/_0_  ;
  output \g63215/_0_  ;
  output \g63216/_0_  ;
  output \g63217/_0_  ;
  output \g63218/_0_  ;
  output \g63219/_0_  ;
  output \g63220/_0_  ;
  output \g63221/_0_  ;
  output \g63222/_0_  ;
  output \g63223/_0_  ;
  output \g63224/_0_  ;
  output \g63225/_0_  ;
  output \g63226/_0_  ;
  output \g63228/_0_  ;
  output \g63229/_0_  ;
  output \g63231/_0_  ;
  output \g63232/_0_  ;
  output \g63233/_0_  ;
  output \g63234/_0_  ;
  output \g63235/_0_  ;
  output \g63236/_0_  ;
  output \g63237/_0_  ;
  output \g63238/_0_  ;
  output \g63239/_0_  ;
  output \g63240/_0_  ;
  output \g63241/_0_  ;
  output \g63242/_0_  ;
  output \g63244/_0_  ;
  output \g63246/_0_  ;
  output \g63247/_0_  ;
  output \g63248/_0_  ;
  output \g63249/_0_  ;
  output \g63250/_0_  ;
  output \g63251/_0_  ;
  output \g63252/_0_  ;
  output \g63253/_0_  ;
  output \g63254/_0_  ;
  output \g63255/_0_  ;
  output \g63256/_0_  ;
  output \g63257/_0_  ;
  output \g63258/_0_  ;
  output \g63259/_0_  ;
  output \g63260/_0_  ;
  output \g63261/_0_  ;
  output \g63262/_0_  ;
  output \g63263/_0_  ;
  output \g63264/_0_  ;
  output \g63265/_0_  ;
  output \g63266/_0_  ;
  output \g63267/_0_  ;
  output \g63268/_0_  ;
  output \g63269/_0_  ;
  output \g63270/_0_  ;
  output \g63272/_0_  ;
  output \g63291/_0_  ;
  output \g63292/_0_  ;
  output \g63293/_0_  ;
  output \g63294/_0_  ;
  output \g63295/_0_  ;
  output \g63298/_0_  ;
  output \g63299/_0_  ;
  output \g63300/_0_  ;
  output \g63301/_0_  ;
  output \g63302/_0_  ;
  output \g63303/_0_  ;
  output \g63304/_0_  ;
  output \g63305/_0_  ;
  output \g63306/_0_  ;
  output \g63307/_0_  ;
  output \g63308/_0_  ;
  output \g63309/_0_  ;
  output \g63310/_0_  ;
  output \g63311/_0_  ;
  output \g63312/_0_  ;
  output \g63313/_0_  ;
  output \g63314/_0_  ;
  output \g63315/_0_  ;
  output \g63316/_0_  ;
  output \g63317/_0_  ;
  output \g63318/_0_  ;
  output \g63320/_0_  ;
  output \g63322/_0_  ;
  output \g63323/_0_  ;
  output \g63324/_0_  ;
  output \g63325/_0_  ;
  output \g63326/_0_  ;
  output \g63327/_0_  ;
  output \g63328/_0_  ;
  output \g63329/_0_  ;
  output \g63330/_0_  ;
  output \g63331/_0_  ;
  output \g63332/_0_  ;
  output \g63333/_0_  ;
  output \g63334/_0_  ;
  output \g63335/_0_  ;
  output \g63336/_0_  ;
  output \g63337/_0_  ;
  output \g63338/_0_  ;
  output \g63339/_0_  ;
  output \g63340/_0_  ;
  output \g63341/_0_  ;
  output \g63342/_0_  ;
  output \g63343/_0_  ;
  output \g63344/_0_  ;
  output \g63345/_0_  ;
  output \g63346/_0_  ;
  output \g63347/_0_  ;
  output \g63348/_0_  ;
  output \g63349/_0_  ;
  output \g63350/_0_  ;
  output \g63351/_0_  ;
  output \g63352/_0_  ;
  output \g63353/_0_  ;
  output \g63354/_0_  ;
  output \g63355/_0_  ;
  output \g63356/_0_  ;
  output \g63357/_0_  ;
  output \g63358/_0_  ;
  output \g63359/_0_  ;
  output \g63360/_0_  ;
  output \g63361/_0_  ;
  output \g63362/_0_  ;
  output \g63363/_0_  ;
  output \g63364/_0_  ;
  output \g63365/_0_  ;
  output \g63366/_0_  ;
  output \g63367/_0_  ;
  output \g63368/_0_  ;
  output \g63369/_0_  ;
  output \g63370/_0_  ;
  output \g63371/_0_  ;
  output \g63372/_0_  ;
  output \g63373/_0_  ;
  output \g63374/_0_  ;
  output \g63375/_0_  ;
  output \g63376/_0_  ;
  output \g63377/_0_  ;
  output \g63378/_0_  ;
  output \g63379/_0_  ;
  output \g63380/_0_  ;
  output \g63383/_3_  ;
  output \g63386/_0_  ;
  output \g63387/_0_  ;
  output \g63388/_0_  ;
  output \g63389/_0_  ;
  output \g63390/_0_  ;
  output \g63391/_0_  ;
  output \g63392/_0_  ;
  output \g63419/_0_  ;
  output \g63421/_0_  ;
  output \g63422/_0_  ;
  output \g63423/_0_  ;
  output \g63424/_0_  ;
  output \g63425/_0_  ;
  output \g63536/_3_  ;
  output \g63625/_0_  ;
  output \g63628/_0_  ;
  output \g63871/_0_  ;
  output \g63874/_0_  ;
  output \g63889/_0_  ;
  output \g63933/_0_  ;
  output \g63945/_0_  ;
  output \g63959/_0_  ;
  output \g63962/_0_  ;
  output \g63974/_0_  ;
  output \g63977/_0_  ;
  output \g64035/_0_  ;
  output \g64435/_3_  ;
  output \g64939/_0_  ;
  output \g65149/_0_  ;
  output \g65632/_3_  ;
  output \g65633/_0_  ;
  output \g65634/_0_  ;
  output \g65635/_0_  ;
  output \g65636/_0_  ;
  output \g65638/_3_  ;
  output \g65640/_3_  ;
  output \g65999/_0_  ;
  output \g66912/_0_  ;
  output \g66914/_0_  ;
  output \g67555/_3_  ;
  output \g67564/_3_  ;
  output \g67567/_3_  ;
  output \g67735/_0_  ;
  output \g67736/_0_  ;
  output \g67737/_0_  ;
  output \g67738/_0_  ;
  output \g67758/_0_  ;
  output \g67760/_0_  ;
  output \g67761/_0_  ;
  output \g67763/_0_  ;
  output \g67766/_0_  ;
  output \g67810/_0_  ;
  output \g67816/_0_  ;
  output \g67902/_0_  ;
  output \g67927/_0_  ;
  output \g67936/_0_  ;
  output \g68067/_0_  ;
  output \g68068/_0_  ;
  output \g68069/_0_  ;
  output \g68070/_0_  ;
  output \g68071/_0_  ;
  output \g68072/_0_  ;
  output \g68073/_0_  ;
  output \g68074/_0_  ;
  output \g68075/_0_  ;
  output \g68076/_0_  ;
  output \g68077/_0_  ;
  output \g68078/_0_  ;
  output \g68079/_0_  ;
  output \g68080/_0_  ;
  output \g68081/_0_  ;
  output \g68082/_0_  ;
  output \g68083/_0_  ;
  output \g68084/_0_  ;
  output \g68085/_0_  ;
  output \g68086/_0_  ;
  output \g68087/_0_  ;
  output \g68088/_0_  ;
  output \g68089/_0_  ;
  output \g68090/_0_  ;
  output \g68091/_0_  ;
  output \g68096/_0_  ;
  output \g68160/_0_  ;
  output \g68218/_0_  ;
  output \g68219/_0_  ;
  output \g68220/_0_  ;
  output \g68221/_0_  ;
  output \g68222/_0_  ;
  output \g68226/_0_  ;
  output \g68247/_0_  ;
  output \g68252/_0_  ;
  output \g68632/_0_  ;
  output \g68633/_0_  ;
  output \g68635/_0_  ;
  output \g68640/_0_  ;
  output \g68642/_0_  ;
  output \g68643/_0_  ;
  output \g68644/_0_  ;
  output \g68645/_0_  ;
  output \g68649/_0_  ;
  output \g68668/_2_  ;
  output \g68670/_0_  ;
  output \g68681/_3_  ;
  output \g68689/_0_  ;
  output \g68690/_0_  ;
  output \g68691/_0_  ;
  output \g68692/_0_  ;
  output \g68693/_0_  ;
  output \g68694/_0_  ;
  output \g68695/_0_  ;
  output \g68737/_0_  ;
  output \g68742/_0_  ;
  output \g68745/_0_  ;
  output \g68750/_0_  ;
  output \g68759/_0_  ;
  output \g68761/_0_  ;
  output \g68774/_0_  ;
  output \g68775/_0_  ;
  output \g68776/_0_  ;
  output \g68777/_0_  ;
  output \g68778/_0_  ;
  output \g68780/_0_  ;
  output \g68781/_0_  ;
  output \g68782/_0_  ;
  output \g68783/_0_  ;
  output \g68784/_0_  ;
  output \g68785/_0_  ;
  output \g68786/_0_  ;
  output \g68787/_0_  ;
  output \g68790/_0_  ;
  output \g68791/_0_  ;
  output \g68793/_0_  ;
  output \g68794/_0_  ;
  output \g68795/_0_  ;
  output \g68796/_0_  ;
  output \g68797/_0_  ;
  output \g68804/_0_  ;
  output \g68805/_0_  ;
  output \g68807/_0_  ;
  output \g68809/_0_  ;
  output \g68864/_3_  ;
  output \g68865/_3_  ;
  output \g68866/_3_  ;
  output \g68867/_3_  ;
  output \g68868/_3_  ;
  output \g68869/_3_  ;
  output \g68870/_3_  ;
  output \g68871/_3_  ;
  output \g68872/_3_  ;
  output \g68873/_3_  ;
  output \g68874/_3_  ;
  output \g68875/_3_  ;
  output \g68876/_3_  ;
  output \g68877/_3_  ;
  output \g68878/_3_  ;
  output \g68879/_3_  ;
  output \g68880/_3_  ;
  output \g68881/_3_  ;
  output \g68882/_3_  ;
  output \g68883/_3_  ;
  output \g68884/_3_  ;
  output \g68885/_3_  ;
  output \g68886/_3_  ;
  output \g68887/_3_  ;
  output \g68888/_3_  ;
  output \g68889/_3_  ;
  output \g68890/_3_  ;
  output \g68891/_3_  ;
  output \g68892/_3_  ;
  output \g68893/_3_  ;
  output \g68894/_3_  ;
  output \g68895/_3_  ;
  output \g69037/_1__syn_2  ;
  output \g69077/_0_  ;
  output \g69081/_0_  ;
  output \g69084/_0_  ;
  output \g69085/_0_  ;
  output \g69086/_0_  ;
  output \g69088/_0_  ;
  output \g69094/_0_  ;
  output \g69095/_0_  ;
  output \g69097/_0_  ;
  output \g69114/_3_  ;
  output \g69116/_3_  ;
  output \g69118/_3_  ;
  output \g69120/_3_  ;
  output \g69122/_3_  ;
  output \g69124/_3_  ;
  output \g69126/_3_  ;
  output \g69128/_3_  ;
  output \g69581/_3_  ;
  output \g70303/_1__syn_2  ;
  output \g70304/_1__syn_2  ;
  output \g70305/_1__syn_2  ;
  output \g70306/_1__syn_2  ;
  output \g70353/_1__syn_2  ;
  output \g70359/_2_  ;
  output \g70364/_1__syn_2  ;
  output \g70375/_1__syn_2  ;
  output \g70380/_2_  ;
  output \g70383/_1__syn_2  ;
  output \g70394/_2_  ;
  output \g70395/_2_  ;
  output \g70396/_1__syn_2  ;
  output \g70398/_1__syn_2  ;
  output \g70407/_1_  ;
  output \g70416/_1__syn_2  ;
  output \g70418/_1__syn_2  ;
  output \g70419/_2_  ;
  output \g70424/_1_  ;
  output \g70465/_2_  ;
  output \g70511/_1_  ;
  output \g70512/_1_  ;
  output \g70513/_2_  ;
  output \g70514/_2_  ;
  output \g70516/_2_  ;
  output \g70518/_2_  ;
  output \g70519/_2_  ;
  output \g70520/_2_  ;
  output \g70530/_2_  ;
  output \g70534/_3_  ;
  output \g70536/_3_  ;
  output \g70540/_3_  ;
  output \g70541/_2_  ;
  output \g70545/_3_  ;
  output \g70546/_2_  ;
  output \g70547/_2_  ;
  output \g70550/_3_  ;
  output \g70551/_2_  ;
  output \g70552/_2_  ;
  output \g70558/_3_  ;
  output \g70559/_2_  ;
  output \g70560/_2_  ;
  output \g70562/_3_  ;
  output \g70564/_3_  ;
  output \g70567/_3_  ;
  output \g70568/_2_  ;
  output \g70571/_3_  ;
  output \g70577/_0_  ;
  output \g70578/_2_  ;
  output \g70585/_3_  ;
  output \g70586/_2_  ;
  output \g70587/_2_  ;
  output \g70588/_3_  ;
  output \g70602/_3_  ;
  output \g70841/_0_  ;
  output \g70842/_0_  ;
  output \g70843/_0_  ;
  output \g70844/_0_  ;
  output \g70845/_0_  ;
  output \g70846/_0_  ;
  output \g70847/_0_  ;
  output \g70848/_0_  ;
  output \g70849/_0_  ;
  output \g70850/_0_  ;
  output \g70851/_0_  ;
  output \g70852/_0_  ;
  output \g70853/_0_  ;
  output \g70854/_0_  ;
  output \g70855/_0_  ;
  output \g70856/_0_  ;
  output \g70857/_0_  ;
  output \g70858/_0_  ;
  output \g70859/_0_  ;
  output \g70860/_0_  ;
  output \g70861/_0_  ;
  output \g70862/_0_  ;
  output \g70863/_0_  ;
  output \g70864/_0_  ;
  output \g70865/_0_  ;
  output \g70866/_0_  ;
  output \g70867/_0_  ;
  output \g70868/_0_  ;
  output \g70869/_0_  ;
  output \g70870/_0_  ;
  output \g70871/_0_  ;
  output \g70872/_0_  ;
  output \g70944/_1__syn_2  ;
  output \g71042/_1__syn_2  ;
  output \g71064/_1__syn_2  ;
  output \g71065/_1__syn_2  ;
  output \g71076/_1__syn_2  ;
  output \g71077/_1__syn_2  ;
  output \g71202/_1__syn_2  ;
  output \g71204/_1__syn_2  ;
  output \g71236/_0_  ;
  output \g71237/_0_  ;
  output \g71241/_0_  ;
  output \g71242/_0_  ;
  output \g71245/_0_  ;
  output \g71246/_0_  ;
  output \g71306/_0_  ;
  output \g71308/_0_  ;
  output \g71309/_0_  ;
  output \g71310/_0_  ;
  output \g71355/_0_  ;
  output \g71416/_0_  ;
  output \g71417/_0_  ;
  output \g71420/_0_  ;
  output \g71432/_0_  ;
  output \g71434/_0_  ;
  output \g71435/_0_  ;
  output \g71436/_0_  ;
  output \g71446/_0_  ;
  output \g71449/_0_  ;
  output \g71451/_0_  ;
  output \g71452/_0_  ;
  output \g71485/_0_  ;
  output \g71494/_0_  ;
  output \g71499/_0_  ;
  output \g71500/_0_  ;
  output \g71501/_0_  ;
  output \g71502/_0_  ;
  output \g71503/_0_  ;
  output \g71504/_0_  ;
  output \g71505/_0_  ;
  output \g71506/_0_  ;
  output \g71815/_0_  ;
  output \g71823/_0_  ;
  output \g71832/_0_  ;
  output \g71833/_0__syn_2  ;
  output \g71837/_0_  ;
  output \g71838/_0_  ;
  output \g71846/_1__syn_2  ;
  output \g71847/_1__syn_2  ;
  output \g71849/_0_  ;
  output \g71854/_0_  ;
  output \g71858/_1__syn_2  ;
  output \g71859/_1__syn_2  ;
  output \g71863/_0_  ;
  output \g71867/_0_  ;
  output \g71869/_0_  ;
  output \g71872/_1_  ;
  output \g71873/_1__syn_2  ;
  output \g71874/_1__syn_2  ;
  output \g71875/_0_  ;
  output \g71877/_1__syn_2  ;
  output \g71881/_0_  ;
  output \g71906/_0_  ;
  output \g71907/_1__syn_2  ;
  output \g71910/_0_  ;
  output \g71911/_0_  ;
  output \g71912/_1__syn_2  ;
  output \g71913/_1__syn_2  ;
  output \g71914/_1__syn_2  ;
  output \g71918/_0_  ;
  output \g71921/_0_  ;
  output \g71922/_0_  ;
  output \g71929/_1__syn_2  ;
  output \g71931/_1__syn_2  ;
  output \g71938/_1__syn_2  ;
  output \g71942/_0_  ;
  output \g71946/_1__syn_2  ;
  output \g71947/_0_  ;
  output \g71951/_0_  ;
  output \g71958/_1__syn_2  ;
  output \g71965/_0_  ;
  output \g71970/_1__syn_2  ;
  output \g71972/_1__syn_2  ;
  output \g71973/_1__syn_2  ;
  output \g71986/_1__syn_2  ;
  output \g71987/_1__syn_2  ;
  output \g71990/_1__syn_2  ;
  output \g71991/_1__syn_2  ;
  output \g71992/_1__syn_2  ;
  output \g71994/_1__syn_2  ;
  output \g71997/_1__syn_2  ;
  output \g72001/_1__syn_2  ;
  output \g72013/_1__syn_2  ;
  output \g72021/_1__syn_2  ;
  output \g72030/_0_  ;
  output \g72031/_0__syn_2  ;
  output \g72036/_1__syn_2  ;
  output \g72038/_0_  ;
  output \g72042/_1__syn_2  ;
  output \g72047/_1__syn_2  ;
  output \g72048/_1__syn_2  ;
  output \g72049/_1__syn_2  ;
  output \g72056/_0_  ;
  output \g72064/_1__syn_2  ;
  output \g72073/_1__syn_2  ;
  output \g72075/_0_  ;
  output \g72078/_0_  ;
  output \g72081/_0_  ;
  output \g72091/_0_  ;
  output \g72096/_0_  ;
  output \g72100/_1__syn_2  ;
  output \g72113/_0_  ;
  output \g72118/_0_  ;
  output \g72121/_1__syn_2  ;
  output \g72122/_1__syn_2  ;
  output \g72125/_1__syn_2  ;
  output \g72128/_0_  ;
  output \g72140/_0_  ;
  output \g72144/_1__syn_2  ;
  output \g72154/_1__syn_2  ;
  output \g72159/_0_  ;
  output \g72164/_1__syn_2  ;
  output \g72165/_1__syn_2  ;
  output \g72167/_1__syn_2  ;
  output \g72170/_1__syn_2  ;
  output \g72172/_1__syn_2  ;
  output \g72173/_0_  ;
  output \g72177/_1__syn_2  ;
  output \g72189/_0_  ;
  output \g72194/_0_  ;
  output \g72196/_0_  ;
  output \g72198/_0_  ;
  output \g72206/_1__syn_2  ;
  output \g72209/_1__syn_2  ;
  output \g72210/_1__syn_2  ;
  output \g72211/_0_  ;
  output \g72215/_0_  ;
  output \g72227/_1__syn_2  ;
  output \g72229/_1__syn_2  ;
  output \g72230/_0_  ;
  output \g72239/_0_  ;
  output \g72250/_3_  ;
  output \g72251/_3_  ;
  output \g72252/_3_  ;
  output \g72253/_3_  ;
  output \g72254/_3_  ;
  output \g72255/_3_  ;
  output \g72256/_3_  ;
  output \g72257/_3_  ;
  output \g72259/_3_  ;
  output \g72260/_3_  ;
  output \g72261/_3_  ;
  output \g72262/_3_  ;
  output \g72263/_3_  ;
  output \g72264/_3_  ;
  output \g72265/_3_  ;
  output \g72266/_3_  ;
  output \g72267/_3_  ;
  output \g72273/_3_  ;
  output \g72275/_3_  ;
  output \g72282/_3_  ;
  output \g72285/_3_  ;
  output \g72293/_3_  ;
  output \g72304/_3_  ;
  output \g72305/_3_  ;
  output \g72306/_3_  ;
  output \g72307/_3_  ;
  output \g72309/_3_  ;
  output \g72310/_3_  ;
  output \g72324/_3_  ;
  output \g72325/_3_  ;
  output \g72326/_3_  ;
  output \g72327/_3_  ;
  output \g72711/_0_  ;
  output \g72763/_0_  ;
  output \g72966/_0_  ;
  output \g72967/_0_  ;
  output \g73018/_0_  ;
  output \g73058/_0_  ;
  output \g73062/_0_  ;
  output \g73067/_0_  ;
  output \g73068/_0_  ;
  output \g73207/_0_  ;
  output \g75007/_1__syn_2  ;
  output \g75568/_1_  ;
  output \g75792/_0_  ;
  output \g75836/_0_  ;
  output \g76027/_0_  ;
  output \g76034/_0_  ;
  output \g76108/_0_  ;
  output \g76130/_0_  ;
  output \g76266/_0_  ;
  output \g76315/_0_  ;
  output \g76569/_0_  ;
  output \g76714/_0_  ;
  output \g77122/_1__syn_2  ;
  output \g77709/_1_  ;
  output \g81909/_0_  ;
  output \g81922/_0_  ;
  output \g81926/_1__syn_2  ;
  output \g82197/_1_  ;
  output \g82272/_0_  ;
  output \g82291/_0_  ;
  output \g82716/_0_  ;
  output \g82718/_0_  ;
  output \g82738/_0_  ;
  output \g82769/_0_  ;
  output \g82775/_0_  ;
  output \g82779/_1__syn_2  ;
  output \g82804/_0_  ;
  output \g82810/_0_  ;
  output \g82817/_0_  ;
  output \g82823/_0_  ;
  output \g82835/_0_  ;
  output \g82841/_0_  ;
  output \g82847/_0_  ;
  output \g82853/_0_  ;
  output \g82859/_0_  ;
  output \g82862/_1__syn_2  ;
  output \g82956/_0_  ;
  output \g82959/_1_  ;
  output \g83020/_0_  ;
  output \g83025/_0_  ;
  output \g83078/_0_  ;
  output \g83083/_0_  ;
  output \g83121/_0_  ;
  output \g83135/_0_  ;
  output \g83205/_0_  ;
  output \g83240/_0_  ;
  output \g83509/_1__syn_2  ;
  output \g83769/_0_  ;
  output \h0lock_pad  ;
  output \h1sel_br[7]_pad  ;
  output \h1sel_dma[0]_pad  ;
  output \h1sel_dma[4]_pad  ;
  output \h1sel_dma[7]_pad  ;
  wire n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 ;
  assign n2228 = ~\ahb_slv_slv_ad_d1o_reg[6]/NET0131  & ~\ahb_slv_slv_ad_d1o_reg[7]/NET0131  ;
  assign n2229 = \ahb_slv_slv_wr_d1o_reg/NET0131  & n2228 ;
  assign n2230 = ~\ahb_slv_slv_ad_d1o_reg[2]/NET0131  & \ahb_slv_slv_ad_d1o_reg[8]/NET0131  ;
  assign n2231 = n2229 & n2230 ;
  assign n2232 = \ahb_slv_slv_ad_d1o_reg[5]/NET0131  & \ctl_rf_rf_sel_d1_reg/NET0131  ;
  assign n2233 = \ahb_slv_slv_ad_d1o_reg[3]/NET0131  & ~\ahb_slv_slv_ad_d1o_reg[4]/NET0131  ;
  assign n2234 = n2232 & n2233 ;
  assign n2235 = \ctl_rf_be_d1_reg[0]/P0001  & n2234 ;
  assign n2236 = n2231 & n2235 ;
  assign n2237 = ~\ctl_rf_c1_rf_chsad_reg[7]/NET0131  & ~n2236 ;
  assign n2238 = \ahb_slv_slv_sz_d1o_reg[0]/NET0131  & ~\ahb_slv_slv_sz_d1o_reg[1]/NET0131  ;
  assign n2239 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \ctl_rf_m0end_reg/NET0131  ;
  assign n2240 = n2238 & n2239 ;
  assign n2241 = ~\ahb_slv_slv_sz_d1o_reg[0]/NET0131  & ~\ahb_slv_slv_sz_d1o_reg[1]/NET0131  ;
  assign n2242 = n2239 & n2241 ;
  assign n2243 = \hwdata[7]_pad  & ~n2242 ;
  assign n2244 = \hwdata[31]_pad  & n2242 ;
  assign n2245 = ~n2243 & ~n2244 ;
  assign n2246 = ~n2240 & ~n2245 ;
  assign n2247 = \hwdata[23]_pad  & n2240 ;
  assign n2248 = n2236 & ~n2247 ;
  assign n2249 = ~n2246 & n2248 ;
  assign n2250 = ~n2237 & ~n2249 ;
  assign n2251 = \ahb_slv_slv_ad_d1o_reg[2]/NET0131  & \ahb_slv_slv_ad_d1o_reg[8]/NET0131  ;
  assign n2252 = n2229 & n2251 ;
  assign n2253 = \ctl_rf_be_d1_reg[2]/P0001  & n2234 ;
  assign n2254 = n2252 & n2253 ;
  assign n2255 = ~\ctl_rf_c1_rf_chdad_reg[17]/NET0131  & ~n2254 ;
  assign n2256 = \hwdata[17]_pad  & ~n2242 ;
  assign n2257 = \hwdata[9]_pad  & n2242 ;
  assign n2258 = ~n2256 & ~n2257 ;
  assign n2259 = ~n2240 & ~n2258 ;
  assign n2260 = \hwdata[1]_pad  & n2240 ;
  assign n2261 = n2254 & ~n2260 ;
  assign n2262 = ~n2259 & n2261 ;
  assign n2263 = ~n2255 & ~n2262 ;
  assign n2264 = \ahb_slv_slv_ad_d1o_reg[6]/NET0131  & \ahb_slv_slv_wr_d1o_reg/NET0131  ;
  assign n2265 = ~\ahb_slv_slv_ad_d1o_reg[7]/NET0131  & n2264 ;
  assign n2266 = n2251 & n2265 ;
  assign n2267 = n2253 & n2266 ;
  assign n2268 = ~\ctl_rf_c3_rf_chdad_reg[17]/NET0131  & ~n2267 ;
  assign n2269 = ~n2260 & n2267 ;
  assign n2270 = ~n2259 & n2269 ;
  assign n2271 = ~n2268 & ~n2270 ;
  assign n2272 = ~\ahb_slv_slv_ad_d1o_reg[6]/NET0131  & \ahb_slv_slv_ad_d1o_reg[7]/NET0131  ;
  assign n2273 = \ahb_slv_slv_wr_d1o_reg/NET0131  & n2272 ;
  assign n2274 = n2251 & n2273 ;
  assign n2275 = ~\ahb_slv_slv_ad_d1o_reg[5]/NET0131  & \ctl_rf_rf_sel_d1_reg/NET0131  ;
  assign n2276 = n2233 & n2275 ;
  assign n2277 = \ctl_rf_be_d1_reg[2]/P0001  & n2276 ;
  assign n2278 = n2274 & n2277 ;
  assign n2279 = ~\ctl_rf_c4_rf_chdad_reg[17]/NET0131  & ~n2278 ;
  assign n2280 = ~n2260 & n2278 ;
  assign n2281 = ~n2259 & n2280 ;
  assign n2282 = ~n2279 & ~n2281 ;
  assign n2283 = n2253 & n2274 ;
  assign n2284 = ~\ctl_rf_c5_rf_chdad_reg[17]/NET0131  & ~n2283 ;
  assign n2285 = ~n2260 & n2283 ;
  assign n2286 = ~n2259 & n2285 ;
  assign n2287 = ~n2284 & ~n2286 ;
  assign n2288 = \ahb_slv_slv_ad_d1o_reg[7]/NET0131  & n2264 ;
  assign n2289 = n2251 & n2288 ;
  assign n2290 = n2277 & n2289 ;
  assign n2291 = ~\ctl_rf_c6_rf_chdad_reg[17]/NET0131  & ~n2290 ;
  assign n2292 = ~n2260 & n2290 ;
  assign n2293 = ~n2259 & n2292 ;
  assign n2294 = ~n2291 & ~n2293 ;
  assign n2295 = n2253 & n2289 ;
  assign n2296 = ~\ctl_rf_c7_rf_chdad_reg[17]/NET0131  & ~n2295 ;
  assign n2297 = ~n2260 & n2295 ;
  assign n2298 = ~n2259 & n2297 ;
  assign n2299 = ~n2296 & ~n2298 ;
  assign n2300 = \ctl_rf_be_d1_reg[3]/P0001  & n2234 ;
  assign n2301 = n2231 & n2300 ;
  assign n2302 = ~\ctl_rf_c1_rf_chsad_reg[31]/NET0131  & ~n2301 ;
  assign n2303 = \hwdata[31]_pad  & ~n2242 ;
  assign n2304 = \hwdata[7]_pad  & n2242 ;
  assign n2305 = ~n2303 & ~n2304 ;
  assign n2306 = ~n2240 & ~n2305 ;
  assign n2307 = \hwdata[15]_pad  & n2240 ;
  assign n2308 = n2301 & ~n2307 ;
  assign n2309 = ~n2306 & n2308 ;
  assign n2310 = ~n2302 & ~n2309 ;
  assign n2311 = n2230 & n2265 ;
  assign n2312 = n2300 & n2311 ;
  assign n2313 = ~\ctl_rf_c3_rf_chsad_reg[31]/NET0131  & ~n2312 ;
  assign n2314 = ~n2307 & n2312 ;
  assign n2315 = ~n2306 & n2314 ;
  assign n2316 = ~n2313 & ~n2315 ;
  assign n2317 = n2230 & n2273 ;
  assign n2318 = \ctl_rf_be_d1_reg[3]/P0001  & n2276 ;
  assign n2319 = n2317 & n2318 ;
  assign n2320 = ~\ctl_rf_c4_rf_chsad_reg[31]/NET0131  & ~n2319 ;
  assign n2321 = ~n2307 & n2319 ;
  assign n2322 = ~n2306 & n2321 ;
  assign n2323 = ~n2320 & ~n2322 ;
  assign n2324 = n2230 & n2288 ;
  assign n2325 = n2318 & n2324 ;
  assign n2326 = ~\ctl_rf_c6_rf_chsad_reg[31]/NET0131  & ~n2325 ;
  assign n2327 = ~n2307 & n2325 ;
  assign n2328 = ~n2306 & n2327 ;
  assign n2329 = ~n2326 & ~n2328 ;
  assign n2330 = n2231 & n2318 ;
  assign n2331 = ~\ctl_rf_c0_rf_chsad_reg[31]/NET0131  & ~n2330 ;
  assign n2332 = ~n2307 & n2330 ;
  assign n2333 = ~n2306 & n2332 ;
  assign n2334 = ~n2331 & ~n2333 ;
  assign n2335 = n2266 & n2277 ;
  assign n2336 = ~\ctl_rf_c2_rf_chdad_reg[17]/NET0131  & ~n2335 ;
  assign n2337 = ~n2260 & n2335 ;
  assign n2338 = ~n2259 & n2337 ;
  assign n2339 = ~n2336 & ~n2338 ;
  assign n2340 = n2311 & n2318 ;
  assign n2341 = ~\ctl_rf_c2_rf_chsad_reg[31]/NET0131  & ~n2340 ;
  assign n2342 = ~n2307 & n2340 ;
  assign n2343 = ~n2306 & n2342 ;
  assign n2344 = ~n2341 & ~n2343 ;
  assign n2345 = n2300 & n2317 ;
  assign n2346 = ~\ctl_rf_c5_rf_chsad_reg[31]/NET0131  & ~n2345 ;
  assign n2347 = ~n2307 & n2345 ;
  assign n2348 = ~n2306 & n2347 ;
  assign n2349 = ~n2346 & ~n2348 ;
  assign n2350 = n2300 & n2324 ;
  assign n2351 = ~\ctl_rf_c7_rf_chsad_reg[31]/NET0131  & ~n2350 ;
  assign n2352 = ~n2307 & n2350 ;
  assign n2353 = ~n2306 & n2352 ;
  assign n2354 = ~n2351 & ~n2353 ;
  assign n2355 = n2252 & n2277 ;
  assign n2356 = ~\ctl_rf_c0_rf_chdad_reg[17]/NET0131  & ~n2355 ;
  assign n2357 = ~n2260 & n2355 ;
  assign n2358 = ~n2259 & n2357 ;
  assign n2359 = ~n2356 & ~n2358 ;
  assign n2360 = n2231 & n2253 ;
  assign n2361 = ~\ctl_rf_c1_rf_chsad_reg[21]/NET0131  & ~n2360 ;
  assign n2362 = \hwdata[21]_pad  & ~n2242 ;
  assign n2363 = \hwdata[13]_pad  & n2242 ;
  assign n2364 = ~n2362 & ~n2363 ;
  assign n2365 = ~n2240 & ~n2364 ;
  assign n2366 = \hwdata[5]_pad  & n2240 ;
  assign n2367 = n2360 & ~n2366 ;
  assign n2368 = ~n2365 & n2367 ;
  assign n2369 = ~n2361 & ~n2368 ;
  assign n2370 = n2253 & n2311 ;
  assign n2371 = ~\ctl_rf_c3_rf_chsad_reg[21]/NET0131  & ~n2370 ;
  assign n2372 = ~n2366 & n2370 ;
  assign n2373 = ~n2365 & n2372 ;
  assign n2374 = ~n2371 & ~n2373 ;
  assign n2375 = n2277 & n2317 ;
  assign n2376 = ~\ctl_rf_c4_rf_chsad_reg[21]/NET0131  & ~n2375 ;
  assign n2377 = ~n2366 & n2375 ;
  assign n2378 = ~n2365 & n2377 ;
  assign n2379 = ~n2376 & ~n2378 ;
  assign n2380 = n2253 & n2317 ;
  assign n2381 = ~\ctl_rf_c5_rf_chsad_reg[21]/NET0131  & ~n2380 ;
  assign n2382 = ~n2366 & n2380 ;
  assign n2383 = ~n2365 & n2382 ;
  assign n2384 = ~n2381 & ~n2383 ;
  assign n2385 = n2277 & n2324 ;
  assign n2386 = ~\ctl_rf_c6_rf_chsad_reg[21]/NET0131  & ~n2385 ;
  assign n2387 = ~n2366 & n2385 ;
  assign n2388 = ~n2365 & n2387 ;
  assign n2389 = ~n2386 & ~n2388 ;
  assign n2390 = n2253 & n2324 ;
  assign n2391 = ~\ctl_rf_c7_rf_chsad_reg[21]/NET0131  & ~n2390 ;
  assign n2392 = ~n2366 & n2390 ;
  assign n2393 = ~n2365 & n2392 ;
  assign n2394 = ~n2391 & ~n2393 ;
  assign n2395 = ~\ctl_rf_c1_rf_chdad_reg[18]/NET0131  & ~n2254 ;
  assign n2396 = \hwdata[18]_pad  & ~n2242 ;
  assign n2397 = \hwdata[10]_pad  & n2242 ;
  assign n2398 = ~n2396 & ~n2397 ;
  assign n2399 = ~n2240 & ~n2398 ;
  assign n2400 = \hwdata[2]_pad  & n2240 ;
  assign n2401 = n2254 & ~n2400 ;
  assign n2402 = ~n2399 & n2401 ;
  assign n2403 = ~n2395 & ~n2402 ;
  assign n2404 = ~\ctl_rf_c1_rf_chdad_reg[19]/NET0131  & ~n2254 ;
  assign n2405 = \hwdata[19]_pad  & ~n2242 ;
  assign n2406 = \hwdata[11]_pad  & n2242 ;
  assign n2407 = ~n2405 & ~n2406 ;
  assign n2408 = ~n2240 & ~n2407 ;
  assign n2409 = \hwdata[3]_pad  & n2240 ;
  assign n2410 = n2254 & ~n2409 ;
  assign n2411 = ~n2408 & n2410 ;
  assign n2412 = ~n2404 & ~n2411 ;
  assign n2413 = ~\ctl_rf_c3_rf_chdad_reg[18]/NET0131  & ~n2267 ;
  assign n2414 = n2267 & ~n2400 ;
  assign n2415 = ~n2399 & n2414 ;
  assign n2416 = ~n2413 & ~n2415 ;
  assign n2417 = ~\ctl_rf_c3_rf_chdad_reg[19]/NET0131  & ~n2267 ;
  assign n2418 = n2267 & ~n2409 ;
  assign n2419 = ~n2408 & n2418 ;
  assign n2420 = ~n2417 & ~n2419 ;
  assign n2421 = ~\ctl_rf_c3_rf_chsad_reg[18]/NET0131  & ~n2370 ;
  assign n2422 = n2370 & ~n2400 ;
  assign n2423 = ~n2399 & n2422 ;
  assign n2424 = ~n2421 & ~n2423 ;
  assign n2425 = ~\ctl_rf_c3_rf_chsad_reg[19]/NET0131  & ~n2370 ;
  assign n2426 = n2370 & ~n2409 ;
  assign n2427 = ~n2408 & n2426 ;
  assign n2428 = ~n2425 & ~n2427 ;
  assign n2429 = ~\ctl_rf_c4_rf_chdad_reg[19]/NET0131  & ~n2278 ;
  assign n2430 = n2278 & ~n2409 ;
  assign n2431 = ~n2408 & n2430 ;
  assign n2432 = ~n2429 & ~n2431 ;
  assign n2433 = ~\ctl_rf_c4_rf_chdad_reg[18]/NET0131  & ~n2278 ;
  assign n2434 = n2278 & ~n2400 ;
  assign n2435 = ~n2399 & n2434 ;
  assign n2436 = ~n2433 & ~n2435 ;
  assign n2437 = ~\ctl_rf_c4_rf_chsad_reg[18]/NET0131  & ~n2375 ;
  assign n2438 = n2375 & ~n2400 ;
  assign n2439 = ~n2399 & n2438 ;
  assign n2440 = ~n2437 & ~n2439 ;
  assign n2441 = ~\ctl_rf_c4_rf_chsad_reg[19]/NET0131  & ~n2375 ;
  assign n2442 = n2375 & ~n2409 ;
  assign n2443 = ~n2408 & n2442 ;
  assign n2444 = ~n2441 & ~n2443 ;
  assign n2445 = ~\ctl_rf_c5_rf_chdad_reg[18]/NET0131  & ~n2283 ;
  assign n2446 = n2283 & ~n2400 ;
  assign n2447 = ~n2399 & n2446 ;
  assign n2448 = ~n2445 & ~n2447 ;
  assign n2449 = ~\ctl_rf_c5_rf_chdad_reg[19]/NET0131  & ~n2283 ;
  assign n2450 = n2283 & ~n2409 ;
  assign n2451 = ~n2408 & n2450 ;
  assign n2452 = ~n2449 & ~n2451 ;
  assign n2453 = ~\ctl_rf_c5_rf_chsad_reg[18]/NET0131  & ~n2380 ;
  assign n2454 = n2380 & ~n2400 ;
  assign n2455 = ~n2399 & n2454 ;
  assign n2456 = ~n2453 & ~n2455 ;
  assign n2457 = ~\ctl_rf_c5_rf_chsad_reg[19]/NET0131  & ~n2380 ;
  assign n2458 = n2380 & ~n2409 ;
  assign n2459 = ~n2408 & n2458 ;
  assign n2460 = ~n2457 & ~n2459 ;
  assign n2461 = ~\ctl_rf_c6_rf_chdad_reg[18]/NET0131  & ~n2290 ;
  assign n2462 = n2290 & ~n2400 ;
  assign n2463 = ~n2399 & n2462 ;
  assign n2464 = ~n2461 & ~n2463 ;
  assign n2465 = ~\ctl_rf_c6_rf_chdad_reg[19]/NET0131  & ~n2290 ;
  assign n2466 = n2290 & ~n2409 ;
  assign n2467 = ~n2408 & n2466 ;
  assign n2468 = ~n2465 & ~n2467 ;
  assign n2469 = ~\ctl_rf_c6_rf_chsad_reg[18]/NET0131  & ~n2385 ;
  assign n2470 = n2385 & ~n2400 ;
  assign n2471 = ~n2399 & n2470 ;
  assign n2472 = ~n2469 & ~n2471 ;
  assign n2473 = ~\ctl_rf_c6_rf_chsad_reg[19]/NET0131  & ~n2385 ;
  assign n2474 = n2385 & ~n2409 ;
  assign n2475 = ~n2408 & n2474 ;
  assign n2476 = ~n2473 & ~n2475 ;
  assign n2477 = ~\ctl_rf_c7_rf_chsad_reg[18]/NET0131  & ~n2390 ;
  assign n2478 = n2390 & ~n2400 ;
  assign n2479 = ~n2399 & n2478 ;
  assign n2480 = ~n2477 & ~n2479 ;
  assign n2481 = ~\ctl_rf_c7_rf_chsad_reg[19]/NET0131  & ~n2390 ;
  assign n2482 = n2390 & ~n2409 ;
  assign n2483 = ~n2408 & n2482 ;
  assign n2484 = ~n2481 & ~n2483 ;
  assign n2485 = n2231 & n2277 ;
  assign n2486 = ~\ctl_rf_c0_rf_chsad_reg[21]/NET0131  & ~n2485 ;
  assign n2487 = ~n2366 & n2485 ;
  assign n2488 = ~n2365 & n2487 ;
  assign n2489 = ~n2486 & ~n2488 ;
  assign n2490 = n2277 & n2311 ;
  assign n2491 = ~\ctl_rf_c2_rf_chsad_reg[21]/NET0131  & ~n2490 ;
  assign n2492 = ~n2366 & n2490 ;
  assign n2493 = ~n2365 & n2492 ;
  assign n2494 = ~n2491 & ~n2493 ;
  assign n2495 = ~\ctl_rf_c1_rf_chsad_reg[22]/NET0131  & ~n2360 ;
  assign n2496 = \hwdata[22]_pad  & ~n2242 ;
  assign n2497 = \hwdata[14]_pad  & n2242 ;
  assign n2498 = ~n2496 & ~n2497 ;
  assign n2499 = ~n2240 & ~n2498 ;
  assign n2500 = \hwdata[6]_pad  & n2240 ;
  assign n2501 = n2360 & ~n2500 ;
  assign n2502 = ~n2499 & n2501 ;
  assign n2503 = ~n2495 & ~n2502 ;
  assign n2504 = ~\ctl_rf_c3_rf_chsad_reg[22]/NET0131  & ~n2370 ;
  assign n2505 = n2370 & ~n2500 ;
  assign n2506 = ~n2499 & n2505 ;
  assign n2507 = ~n2504 & ~n2506 ;
  assign n2508 = ~\ctl_rf_c4_rf_chsad_reg[22]/NET0131  & ~n2375 ;
  assign n2509 = n2375 & ~n2500 ;
  assign n2510 = ~n2499 & n2509 ;
  assign n2511 = ~n2508 & ~n2510 ;
  assign n2512 = ~\ctl_rf_c5_rf_chsad_reg[22]/NET0131  & ~n2380 ;
  assign n2513 = n2380 & ~n2500 ;
  assign n2514 = ~n2499 & n2513 ;
  assign n2515 = ~n2512 & ~n2514 ;
  assign n2516 = ~\ctl_rf_c6_rf_chsad_reg[22]/NET0131  & ~n2385 ;
  assign n2517 = n2385 & ~n2500 ;
  assign n2518 = ~n2499 & n2517 ;
  assign n2519 = ~n2516 & ~n2518 ;
  assign n2520 = ~\ctl_rf_c7_rf_chsad_reg[22]/NET0131  & ~n2390 ;
  assign n2521 = n2390 & ~n2500 ;
  assign n2522 = ~n2499 & n2521 ;
  assign n2523 = ~n2520 & ~n2522 ;
  assign n2524 = ~\ctl_rf_c1_rf_chsad_reg[23]/NET0131  & ~n2360 ;
  assign n2525 = \hwdata[23]_pad  & ~n2242 ;
  assign n2526 = \hwdata[15]_pad  & n2242 ;
  assign n2527 = ~n2525 & ~n2526 ;
  assign n2528 = ~n2240 & ~n2527 ;
  assign n2529 = \hwdata[7]_pad  & n2240 ;
  assign n2530 = n2360 & ~n2529 ;
  assign n2531 = ~n2528 & n2530 ;
  assign n2532 = ~n2524 & ~n2531 ;
  assign n2533 = ~\ctl_rf_c3_rf_chsad_reg[23]/NET0131  & ~n2370 ;
  assign n2534 = n2370 & ~n2529 ;
  assign n2535 = ~n2528 & n2534 ;
  assign n2536 = ~n2533 & ~n2535 ;
  assign n2537 = ~\ctl_rf_c4_rf_chsad_reg[23]/NET0131  & ~n2375 ;
  assign n2538 = n2375 & ~n2529 ;
  assign n2539 = ~n2528 & n2538 ;
  assign n2540 = ~n2537 & ~n2539 ;
  assign n2541 = ~\ctl_rf_c5_rf_chsad_reg[23]/NET0131  & ~n2380 ;
  assign n2542 = n2380 & ~n2529 ;
  assign n2543 = ~n2528 & n2542 ;
  assign n2544 = ~n2541 & ~n2543 ;
  assign n2545 = ~\ctl_rf_c6_rf_chsad_reg[23]/NET0131  & ~n2385 ;
  assign n2546 = n2385 & ~n2529 ;
  assign n2547 = ~n2528 & n2546 ;
  assign n2548 = ~n2545 & ~n2547 ;
  assign n2549 = ~\ctl_rf_c7_rf_chsad_reg[23]/NET0131  & ~n2390 ;
  assign n2550 = n2390 & ~n2529 ;
  assign n2551 = ~n2528 & n2550 ;
  assign n2552 = ~n2549 & ~n2551 ;
  assign n2553 = ~\ctl_rf_c0_rf_chsad_reg[18]/NET0131  & ~n2485 ;
  assign n2554 = ~n2400 & n2485 ;
  assign n2555 = ~n2399 & n2554 ;
  assign n2556 = ~n2553 & ~n2555 ;
  assign n2557 = ~\ctl_rf_c0_rf_chsad_reg[19]/NET0131  & ~n2485 ;
  assign n2558 = ~n2409 & n2485 ;
  assign n2559 = ~n2408 & n2558 ;
  assign n2560 = ~n2557 & ~n2559 ;
  assign n2561 = ~\ctl_rf_c1_rf_chsad_reg[20]/NET0131  & ~n2360 ;
  assign n2562 = \hwdata[20]_pad  & ~n2242 ;
  assign n2563 = \hwdata[12]_pad  & n2242 ;
  assign n2564 = ~n2562 & ~n2563 ;
  assign n2565 = ~n2240 & ~n2564 ;
  assign n2566 = \hwdata[4]_pad  & n2240 ;
  assign n2567 = n2360 & ~n2566 ;
  assign n2568 = ~n2565 & n2567 ;
  assign n2569 = ~n2561 & ~n2568 ;
  assign n2570 = ~\ctl_rf_c1_rf_chsad_reg[24]/NET0131  & ~n2301 ;
  assign n2571 = \hwdata[24]_pad  & ~n2242 ;
  assign n2572 = \hwdata[0]_pad  & n2242 ;
  assign n2573 = ~n2571 & ~n2572 ;
  assign n2574 = ~n2240 & ~n2573 ;
  assign n2575 = \hwdata[8]_pad  & n2240 ;
  assign n2576 = n2301 & ~n2575 ;
  assign n2577 = ~n2574 & n2576 ;
  assign n2578 = ~n2570 & ~n2577 ;
  assign n2579 = ~\ctl_rf_c2_rf_chdad_reg[18]/NET0131  & ~n2335 ;
  assign n2580 = n2335 & ~n2400 ;
  assign n2581 = ~n2399 & n2580 ;
  assign n2582 = ~n2579 & ~n2581 ;
  assign n2583 = ~\ctl_rf_c2_rf_chdad_reg[19]/NET0131  & ~n2335 ;
  assign n2584 = n2335 & ~n2409 ;
  assign n2585 = ~n2408 & n2584 ;
  assign n2586 = ~n2583 & ~n2585 ;
  assign n2587 = ~\ctl_rf_c2_rf_chsad_reg[19]/NET0131  & ~n2490 ;
  assign n2588 = ~n2409 & n2490 ;
  assign n2589 = ~n2408 & n2588 ;
  assign n2590 = ~n2587 & ~n2589 ;
  assign n2591 = ~\ctl_rf_c2_rf_chsad_reg[18]/NET0131  & ~n2490 ;
  assign n2592 = ~n2400 & n2490 ;
  assign n2593 = ~n2399 & n2592 ;
  assign n2594 = ~n2591 & ~n2593 ;
  assign n2595 = ~\ctl_rf_c3_rf_chsad_reg[20]/NET0131  & ~n2370 ;
  assign n2596 = n2370 & ~n2566 ;
  assign n2597 = ~n2565 & n2596 ;
  assign n2598 = ~n2595 & ~n2597 ;
  assign n2599 = ~\ctl_rf_c3_rf_chsad_reg[24]/NET0131  & ~n2312 ;
  assign n2600 = n2312 & ~n2575 ;
  assign n2601 = ~n2574 & n2600 ;
  assign n2602 = ~n2599 & ~n2601 ;
  assign n2603 = ~\ctl_rf_c4_rf_chsad_reg[20]/NET0131  & ~n2375 ;
  assign n2604 = n2375 & ~n2566 ;
  assign n2605 = ~n2565 & n2604 ;
  assign n2606 = ~n2603 & ~n2605 ;
  assign n2607 = ~\ctl_rf_c4_rf_chsad_reg[24]/NET0131  & ~n2319 ;
  assign n2608 = n2319 & ~n2575 ;
  assign n2609 = ~n2574 & n2608 ;
  assign n2610 = ~n2607 & ~n2609 ;
  assign n2611 = ~\ctl_rf_c6_rf_chsad_reg[20]/NET0131  & ~n2385 ;
  assign n2612 = n2385 & ~n2566 ;
  assign n2613 = ~n2565 & n2612 ;
  assign n2614 = ~n2611 & ~n2613 ;
  assign n2615 = ~\ctl_rf_c6_rf_chsad_reg[24]/NET0131  & ~n2325 ;
  assign n2616 = n2325 & ~n2575 ;
  assign n2617 = ~n2574 & n2616 ;
  assign n2618 = ~n2615 & ~n2617 ;
  assign n2619 = ~\ctl_rf_c0_rf_chdad_reg[18]/NET0131  & ~n2355 ;
  assign n2620 = n2355 & ~n2400 ;
  assign n2621 = ~n2399 & n2620 ;
  assign n2622 = ~n2619 & ~n2621 ;
  assign n2623 = ~\ctl_rf_c0_rf_chdad_reg[19]/NET0131  & ~n2355 ;
  assign n2624 = n2355 & ~n2409 ;
  assign n2625 = ~n2408 & n2624 ;
  assign n2626 = ~n2623 & ~n2625 ;
  assign n2627 = ~\ctl_rf_c0_rf_chsad_reg[20]/NET0131  & ~n2485 ;
  assign n2628 = n2485 & ~n2566 ;
  assign n2629 = ~n2565 & n2628 ;
  assign n2630 = ~n2627 & ~n2629 ;
  assign n2631 = ~\ctl_rf_c0_rf_chsad_reg[22]/NET0131  & ~n2485 ;
  assign n2632 = n2485 & ~n2500 ;
  assign n2633 = ~n2499 & n2632 ;
  assign n2634 = ~n2631 & ~n2633 ;
  assign n2635 = ~\ctl_rf_c0_rf_chsad_reg[23]/NET0131  & ~n2485 ;
  assign n2636 = n2485 & ~n2529 ;
  assign n2637 = ~n2528 & n2636 ;
  assign n2638 = ~n2635 & ~n2637 ;
  assign n2639 = ~\ctl_rf_c0_rf_chsad_reg[24]/NET0131  & ~n2330 ;
  assign n2640 = n2330 & ~n2575 ;
  assign n2641 = ~n2574 & n2640 ;
  assign n2642 = ~n2639 & ~n2641 ;
  assign n2643 = ~\ctl_rf_c2_rf_chsad_reg[20]/NET0131  & ~n2490 ;
  assign n2644 = n2490 & ~n2566 ;
  assign n2645 = ~n2565 & n2644 ;
  assign n2646 = ~n2643 & ~n2645 ;
  assign n2647 = ~\ctl_rf_c2_rf_chsad_reg[22]/NET0131  & ~n2490 ;
  assign n2648 = n2490 & ~n2500 ;
  assign n2649 = ~n2499 & n2648 ;
  assign n2650 = ~n2647 & ~n2649 ;
  assign n2651 = ~\ctl_rf_c2_rf_chsad_reg[23]/NET0131  & ~n2490 ;
  assign n2652 = n2490 & ~n2529 ;
  assign n2653 = ~n2528 & n2652 ;
  assign n2654 = ~n2651 & ~n2653 ;
  assign n2655 = ~\ctl_rf_c2_rf_chsad_reg[24]/NET0131  & ~n2340 ;
  assign n2656 = n2340 & ~n2575 ;
  assign n2657 = ~n2574 & n2656 ;
  assign n2658 = ~n2655 & ~n2657 ;
  assign n2659 = ~\ctl_rf_c5_rf_chsad_reg[20]/NET0131  & ~n2380 ;
  assign n2660 = n2380 & ~n2566 ;
  assign n2661 = ~n2565 & n2660 ;
  assign n2662 = ~n2659 & ~n2661 ;
  assign n2663 = ~\ctl_rf_c5_rf_chsad_reg[24]/NET0131  & ~n2345 ;
  assign n2664 = n2345 & ~n2575 ;
  assign n2665 = ~n2574 & n2664 ;
  assign n2666 = ~n2663 & ~n2665 ;
  assign n2667 = ~\ctl_rf_c7_rf_chsad_reg[20]/NET0131  & ~n2390 ;
  assign n2668 = n2390 & ~n2566 ;
  assign n2669 = ~n2565 & n2668 ;
  assign n2670 = ~n2667 & ~n2669 ;
  assign n2671 = ~\ctl_rf_c7_rf_chsad_reg[24]/NET0131  & ~n2350 ;
  assign n2672 = n2350 & ~n2575 ;
  assign n2673 = ~n2574 & n2672 ;
  assign n2674 = ~n2671 & ~n2673 ;
  assign n2675 = ~\ctl_rf_c1_rf_chsad_reg[16]/NET0131  & ~n2360 ;
  assign n2676 = \hwdata[16]_pad  & ~n2242 ;
  assign n2677 = \hwdata[8]_pad  & n2242 ;
  assign n2678 = ~n2676 & ~n2677 ;
  assign n2679 = ~n2240 & ~n2678 ;
  assign n2680 = \hwdata[0]_pad  & n2240 ;
  assign n2681 = n2360 & ~n2680 ;
  assign n2682 = ~n2679 & n2681 ;
  assign n2683 = ~n2675 & ~n2682 ;
  assign n2684 = ~\ctl_rf_c3_rf_chsad_reg[16]/NET0131  & ~n2370 ;
  assign n2685 = n2370 & ~n2680 ;
  assign n2686 = ~n2679 & n2685 ;
  assign n2687 = ~n2684 & ~n2686 ;
  assign n2688 = ~\ctl_rf_c4_rf_chdad_reg[16]/NET0131  & ~n2278 ;
  assign n2689 = n2278 & ~n2680 ;
  assign n2690 = ~n2679 & n2689 ;
  assign n2691 = ~n2688 & ~n2690 ;
  assign n2692 = ~\ctl_rf_c4_rf_chsad_reg[16]/NET0131  & ~n2375 ;
  assign n2693 = n2375 & ~n2680 ;
  assign n2694 = ~n2679 & n2693 ;
  assign n2695 = ~n2692 & ~n2694 ;
  assign n2696 = ~\ctl_rf_c6_rf_chdad_reg[16]/NET0131  & ~n2290 ;
  assign n2697 = n2290 & ~n2680 ;
  assign n2698 = ~n2679 & n2697 ;
  assign n2699 = ~n2696 & ~n2698 ;
  assign n2700 = ~\ctl_rf_c6_rf_chsad_reg[16]/NET0131  & ~n2385 ;
  assign n2701 = n2385 & ~n2680 ;
  assign n2702 = ~n2679 & n2701 ;
  assign n2703 = ~n2700 & ~n2702 ;
  assign n2704 = ~\ctl_rf_c0_rf_chsad_reg[16]/NET0131  & ~n2485 ;
  assign n2705 = n2485 & ~n2680 ;
  assign n2706 = ~n2679 & n2705 ;
  assign n2707 = ~n2704 & ~n2706 ;
  assign n2708 = ~\ctl_rf_c1_rf_chdad_reg[16]/NET0131  & ~n2254 ;
  assign n2709 = n2254 & ~n2680 ;
  assign n2710 = ~n2679 & n2709 ;
  assign n2711 = ~n2708 & ~n2710 ;
  assign n2712 = ~\ctl_rf_c2_rf_chdad_reg[16]/NET0131  & ~n2335 ;
  assign n2713 = n2335 & ~n2680 ;
  assign n2714 = ~n2679 & n2713 ;
  assign n2715 = ~n2712 & ~n2714 ;
  assign n2716 = ~\ctl_rf_c2_rf_chsad_reg[16]/NET0131  & ~n2490 ;
  assign n2717 = n2490 & ~n2680 ;
  assign n2718 = ~n2679 & n2717 ;
  assign n2719 = ~n2716 & ~n2718 ;
  assign n2720 = ~\ctl_rf_c3_rf_chdad_reg[16]/NET0131  & ~n2267 ;
  assign n2721 = n2267 & ~n2680 ;
  assign n2722 = ~n2679 & n2721 ;
  assign n2723 = ~n2720 & ~n2722 ;
  assign n2724 = ~\ctl_rf_c5_rf_chdad_reg[16]/NET0131  & ~n2283 ;
  assign n2725 = n2283 & ~n2680 ;
  assign n2726 = ~n2679 & n2725 ;
  assign n2727 = ~n2724 & ~n2726 ;
  assign n2728 = ~\ctl_rf_c5_rf_chsad_reg[16]/NET0131  & ~n2380 ;
  assign n2729 = n2380 & ~n2680 ;
  assign n2730 = ~n2679 & n2729 ;
  assign n2731 = ~n2728 & ~n2730 ;
  assign n2732 = ~\ctl_rf_c7_rf_chdad_reg[16]/NET0131  & ~n2295 ;
  assign n2733 = n2295 & ~n2680 ;
  assign n2734 = ~n2679 & n2733 ;
  assign n2735 = ~n2732 & ~n2734 ;
  assign n2736 = ~\ctl_rf_c7_rf_chsad_reg[16]/NET0131  & ~n2390 ;
  assign n2737 = n2390 & ~n2680 ;
  assign n2738 = ~n2679 & n2737 ;
  assign n2739 = ~n2736 & ~n2738 ;
  assign n2740 = ~\ctl_rf_c0_rf_chdad_reg[16]/NET0131  & ~n2355 ;
  assign n2741 = n2355 & ~n2680 ;
  assign n2742 = ~n2679 & n2741 ;
  assign n2743 = ~n2740 & ~n2742 ;
  assign n2744 = ~\m1_mux_mux_no_reg[2]/NET0131  & \m1_mux_mux_no_reg[3]/NET0131  ;
  assign n2745 = ~\m1_mux_mux_no_reg[0]/NET0131  & \m1_mux_mux_no_reg[1]/NET0131  ;
  assign n2746 = n2744 & n2745 ;
  assign n2747 = \h1rdy2_br_pad  & n2746 ;
  assign n2748 = ~\m1_mux_hrmxnof_reg/NET0131  & ~n2747 ;
  assign n2749 = \m1_mux_mux_no_reg[0]/NET0131  & \m1_mux_mux_no_reg[1]/NET0131  ;
  assign n2750 = \m1_mux_mux_no_reg[2]/NET0131  & \m1_mux_mux_no_reg[3]/NET0131  ;
  assign n2751 = n2749 & n2750 ;
  assign n2752 = \h1rdy7_br_pad  & n2751 ;
  assign n2753 = n2745 & n2750 ;
  assign n2754 = \h1rdy6_br_pad  & n2753 ;
  assign n2755 = ~n2752 & ~n2754 ;
  assign n2756 = ~\m1_mux_mux_no_reg[2]/NET0131  & ~\m1_mux_mux_no_reg[3]/NET0131  ;
  assign n2757 = n2749 & n2756 ;
  assign n2758 = \h1rdy3_dma_pad  & n2757 ;
  assign n2759 = \m1_mux_mux_no_reg[0]/NET0131  & ~\m1_mux_mux_no_reg[1]/NET0131  ;
  assign n2760 = n2756 & n2759 ;
  assign n2761 = \h1rdy1_dma_pad  & n2760 ;
  assign n2762 = ~n2758 & ~n2761 ;
  assign n2763 = n2755 & n2762 ;
  assign n2764 = n2748 & n2763 ;
  assign n2765 = n2744 & n2749 ;
  assign n2766 = \h1rdy3_br_pad  & n2765 ;
  assign n2767 = n2744 & n2759 ;
  assign n2768 = \h1rdy1_br_pad  & n2767 ;
  assign n2769 = \m1_mux_mux_no_reg[2]/NET0131  & ~\m1_mux_mux_no_reg[3]/NET0131  ;
  assign n2770 = n2759 & n2769 ;
  assign n2771 = \h1rdy5_dma_pad  & n2770 ;
  assign n2772 = ~n2768 & ~n2771 ;
  assign n2773 = ~n2766 & n2772 ;
  assign n2774 = n2749 & n2769 ;
  assign n2775 = \h1rdy7_dma_pad  & n2774 ;
  assign n2776 = ~\m1_mux_mux_no_reg[0]/NET0131  & ~\m1_mux_mux_no_reg[1]/NET0131  ;
  assign n2777 = n2750 & n2776 ;
  assign n2778 = \h1rdy4_br_pad  & n2777 ;
  assign n2779 = ~n2775 & ~n2778 ;
  assign n2780 = n2744 & n2776 ;
  assign n2781 = \h1rdy0_br_pad  & n2780 ;
  assign n2782 = n2750 & n2759 ;
  assign n2783 = \h1rdy5_br_pad  & n2782 ;
  assign n2784 = ~n2781 & ~n2783 ;
  assign n2785 = n2779 & n2784 ;
  assign n2786 = n2745 & n2756 ;
  assign n2787 = \h1rdy2_dma_pad  & n2786 ;
  assign n2788 = n2769 & n2776 ;
  assign n2789 = \h1rdy4_dma_pad  & n2788 ;
  assign n2790 = ~n2787 & ~n2789 ;
  assign n2791 = n2745 & n2769 ;
  assign n2792 = \h1rdy6_dma_pad  & n2791 ;
  assign n2793 = n2756 & n2776 ;
  assign n2794 = \h1rdy0_dma_pad  & n2793 ;
  assign n2795 = ~n2792 & ~n2794 ;
  assign n2796 = n2790 & n2795 ;
  assign n2797 = n2785 & n2796 ;
  assign n2798 = n2773 & n2797 ;
  assign n2799 = n2764 & n2798 ;
  assign n2800 = ~\ahb_mst1_mx_cmd_st_reg[1]/NET0131  & ~\ahb_mst1_mx_dtp_reg/NET0131  ;
  assign n2801 = \ahb_slv_slv_br_req_reg/NET0131  & n2800 ;
  assign n2802 = \ahb_slv_slv_br_req_reg/NET0131  & \de_m1_arb_st_reg[1]/NET0131  ;
  assign n2803 = n2801 & ~n2802 ;
  assign n2804 = ~\de_tsz_cnt_reg[10]/NET0131  & ~\de_tsz_cnt_reg[11]/NET0131  ;
  assign n2805 = ~\de_tsz_cnt_reg[2]/NET0131  & ~\de_tsz_cnt_reg[3]/NET0131  ;
  assign n2806 = ~\de_tsz_cnt_reg[4]/NET0131  & ~\de_tsz_cnt_reg[5]/NET0131  ;
  assign n2807 = n2805 & n2806 ;
  assign n2808 = n2804 & n2807 ;
  assign n2809 = ~\de_tsz_cnt_reg[6]/NET0131  & ~\de_tsz_cnt_reg[7]/NET0131  ;
  assign n2810 = ~\de_tsz_cnt_reg[8]/NET0131  & ~\de_tsz_cnt_reg[9]/NET0131  ;
  assign n2811 = n2809 & n2810 ;
  assign n2812 = ~\de_tsz_cnt_reg[0]/NET0131  & ~\de_tsz_cnt_reg[1]/NET0131  ;
  assign n2813 = n2811 & n2812 ;
  assign n2814 = n2808 & n2813 ;
  assign n2815 = ~\de_de_st_reg[1]/NET0131  & ~\de_de_st_reg[2]/NET0131  ;
  assign n2816 = \ch_sel_arb_chcsr_reg_reg[2]/NET0131  & ~n2815 ;
  assign n2817 = ~\de_bst_cnt_reg[5]/NET0131  & ~\de_bst_cnt_reg[6]/NET0131  ;
  assign n2818 = ~\de_bst_cnt_reg[7]/NET0131  & ~\de_bst_cnt_reg[8]/NET0131  ;
  assign n2819 = n2817 & n2818 ;
  assign n2820 = ~\de_bst_cnt_reg[2]/NET0131  & ~\de_bst_cnt_reg[3]/NET0131  ;
  assign n2821 = ~\de_bst_cnt_reg[0]/NET0131  & ~\de_bst_cnt_reg[4]/NET0131  ;
  assign n2822 = n2820 & n2821 ;
  assign n2823 = n2819 & n2822 ;
  assign n2824 = n2816 & ~n2823 ;
  assign n2825 = ~n2814 & n2824 ;
  assign n2826 = \de_de_st_reg[6]/NET0131  & \de_m1_is_llp_reg/NET0131  ;
  assign n2827 = ~n2802 & ~n2826 ;
  assign n2828 = ~n2825 & n2827 ;
  assign n2829 = ~n2803 & ~n2828 ;
  assign n2830 = ~\m1_mux_hrdy_df_reg/NET0131  & \m1_mux_hrmxnof_reg/NET0131  ;
  assign n2831 = ~\de_de_st_reg[5]/NET0131  & n2800 ;
  assign n2832 = ~n2830 & n2831 ;
  assign n2833 = n2829 & n2832 ;
  assign n2834 = ~n2799 & n2833 ;
  assign n2835 = ~\ch_sel_arb_chcsr_reg_reg[3]/NET0131  & ~\ch_sel_arb_chcsr_reg_reg[4]/NET0131  ;
  assign n2836 = ~\de_de_st_reg[6]/NET0131  & \de_m1_arb_st_reg[0]/NET0131  ;
  assign n2837 = ~n2835 & n2836 ;
  assign n2838 = ~\ch_sel_arb_chcsr_reg_reg[5]/NET0131  & ~\ch_sel_arb_chcsr_reg_reg[6]/NET0131  ;
  assign n2839 = ~\de_de_st_reg[6]/NET0131  & ~\de_m1_arb_st_reg[0]/NET0131  ;
  assign n2840 = ~n2838 & n2839 ;
  assign n2841 = ~n2837 & ~n2840 ;
  assign n2842 = ~\de_m1_arb_st_reg[1]/NET0131  & n2841 ;
  assign n2843 = n2834 & ~n2842 ;
  assign n2844 = ~\h1burst[0]_pad  & ~n2834 ;
  assign n2845 = ~n2843 & ~n2844 ;
  assign n2846 = ~\ahb_mst1_mx_cmd_st_reg[0]/NET0131  & ~\ahb_mst1_mx_cmd_st_reg[1]/NET0131  ;
  assign n2847 = n2834 & n2846 ;
  assign n2848 = \m1_mux_hrmxnof_reg/NET0131  & ~\m1_mux_hrp_df_reg[0]/NET0131  ;
  assign n2849 = \h1rp0_br[0]_pad  & n2780 ;
  assign n2850 = ~\m1_mux_hrmxnof_reg/NET0131  & ~n2849 ;
  assign n2851 = \h1rp0_dma[0]_pad  & n2793 ;
  assign n2852 = \h1rp4_dma[0]_pad  & n2788 ;
  assign n2853 = ~n2851 & ~n2852 ;
  assign n2854 = \h1rp2_br[0]_pad  & n2746 ;
  assign n2855 = \h1rp2_dma[0]_pad  & n2786 ;
  assign n2856 = ~n2854 & ~n2855 ;
  assign n2857 = n2853 & n2856 ;
  assign n2858 = n2850 & n2857 ;
  assign n2859 = \h1rp4_br[0]_pad  & n2777 ;
  assign n2860 = \h1rp3_br[0]_pad  & n2765 ;
  assign n2861 = \h1rp1_br[0]_pad  & n2767 ;
  assign n2862 = ~n2860 & ~n2861 ;
  assign n2863 = ~n2859 & n2862 ;
  assign n2864 = \h1rp3_dma[0]_pad  & n2757 ;
  assign n2865 = \h1rp1_dma[0]_pad  & n2760 ;
  assign n2866 = ~n2864 & ~n2865 ;
  assign n2867 = \h1rp5_dma[0]_pad  & n2770 ;
  assign n2868 = \h1rp6_br[0]_pad  & n2753 ;
  assign n2869 = ~n2867 & ~n2868 ;
  assign n2870 = n2866 & n2869 ;
  assign n2871 = \h1rp5_br[0]_pad  & n2782 ;
  assign n2872 = \h1rp7_br[0]_pad  & n2751 ;
  assign n2873 = ~n2871 & ~n2872 ;
  assign n2874 = \h1rp6_dma[0]_pad  & n2791 ;
  assign n2875 = \h1rp7_dma[0]_pad  & n2774 ;
  assign n2876 = ~n2874 & ~n2875 ;
  assign n2877 = n2873 & n2876 ;
  assign n2878 = n2870 & n2877 ;
  assign n2879 = n2863 & n2878 ;
  assign n2880 = n2858 & n2879 ;
  assign n2881 = ~n2848 & ~n2880 ;
  assign n2882 = \h1rp0_dma[1]_pad  & n2793 ;
  assign n2883 = \h1rp5_dma[1]_pad  & n2770 ;
  assign n2884 = ~n2882 & ~n2883 ;
  assign n2885 = \h1rp6_dma[1]_pad  & n2791 ;
  assign n2886 = \h1rp6_br[1]_pad  & n2753 ;
  assign n2887 = ~n2885 & ~n2886 ;
  assign n2888 = n2884 & n2887 ;
  assign n2889 = \h1rp0_br[1]_pad  & n2780 ;
  assign n2890 = \h1rp1_dma[1]_pad  & n2760 ;
  assign n2891 = ~n2889 & ~n2890 ;
  assign n2892 = \h1rp7_dma[1]_pad  & n2774 ;
  assign n2893 = \h1rp5_br[1]_pad  & n2782 ;
  assign n2894 = ~n2892 & ~n2893 ;
  assign n2895 = n2891 & n2894 ;
  assign n2896 = n2888 & n2895 ;
  assign n2897 = \h1rp1_br[1]_pad  & n2767 ;
  assign n2898 = \h1rp7_br[1]_pad  & n2751 ;
  assign n2899 = ~n2897 & ~n2898 ;
  assign n2900 = \h1rp4_dma[1]_pad  & n2788 ;
  assign n2901 = \h1rp4_br[1]_pad  & n2777 ;
  assign n2902 = ~n2900 & ~n2901 ;
  assign n2903 = n2899 & n2902 ;
  assign n2904 = \h1rp3_dma[1]_pad  & n2757 ;
  assign n2905 = \h1rp3_br[1]_pad  & n2765 ;
  assign n2906 = ~n2904 & ~n2905 ;
  assign n2907 = \h1rp2_br[1]_pad  & n2746 ;
  assign n2908 = \h1rp2_dma[1]_pad  & n2786 ;
  assign n2909 = ~n2907 & ~n2908 ;
  assign n2910 = n2906 & n2909 ;
  assign n2911 = n2903 & n2910 ;
  assign n2912 = n2896 & n2911 ;
  assign n2913 = ~\m1_mux_hrmxnof_reg/NET0131  & ~n2912 ;
  assign n2914 = ~\de_m1_arb_st_reg[0]/NET0131  & ~\de_m1_arb_st_reg[1]/NET0131  ;
  assign n2915 = \ch_sel_arb_chcsr_reg_reg[2]/NET0131  & n2914 ;
  assign n2916 = ~\ahb_mst1_mx_cmd_st_reg[0]/NET0131  & ~n2838 ;
  assign n2917 = ~\de_tsz_cnt_reg[0]/NET0131  & \de_tsz_cnt_reg[1]/NET0131  ;
  assign n2918 = n2811 & n2917 ;
  assign n2919 = n2808 & n2918 ;
  assign n2920 = ~n2916 & ~n2919 ;
  assign n2921 = n2915 & ~n2920 ;
  assign n2922 = \de_m1_arb_st_reg[0]/NET0131  & ~\de_m1_arb_st_reg[1]/NET0131  ;
  assign n2923 = ~\ahb_mst1_mx_cmd_st_reg[0]/NET0131  & \ch_sel_arb_chcsr_reg_reg[1]/NET0131  ;
  assign n2924 = ~n2835 & n2923 ;
  assign n2925 = n2922 & n2924 ;
  assign n2926 = \ahb_mst1_mx_cmd_st_reg[1]/NET0131  & ~\ahb_slv_slv_br_req_reg/NET0131  ;
  assign n2927 = ~n2925 & n2926 ;
  assign n2928 = ~n2921 & n2927 ;
  assign n2929 = ~n2913 & n2928 ;
  assign n2930 = ~n2881 & n2929 ;
  assign n2931 = ~n2847 & ~n2930 ;
  assign n2932 = ~\ahb_mst0_mx_cmd_st_reg[1]/NET0131  & ~\ahb_mst0_mx_dtp_reg/NET0131  ;
  assign n2933 = ~\de_de_st_reg[5]/NET0131  & \h0grant_pad  ;
  assign n2934 = \h0readyin_pad  & n2933 ;
  assign n2935 = n2932 & n2934 ;
  assign n2936 = ~\h0burst[0]_pad  & ~n2935 ;
  assign n2937 = ~\ch_sel_arb_chcsr_reg_reg[2]/NET0131  & ~n2815 ;
  assign n2938 = ~n2823 & n2937 ;
  assign n2939 = ~n2814 & n2938 ;
  assign n2940 = \de_de_st_reg[6]/NET0131  & \de_m0_is_llp_reg/NET0131  ;
  assign n2941 = ~\h0burst[0]_pad  & ~n2940 ;
  assign n2942 = ~n2939 & n2941 ;
  assign n2943 = ~n2936 & ~n2942 ;
  assign n2944 = ~n2939 & ~n2940 ;
  assign n2945 = ~\de_de_st_reg[6]/NET0131  & \de_m0_arb_st_reg/NET0131  ;
  assign n2946 = ~n2835 & n2945 ;
  assign n2947 = ~\de_de_st_reg[6]/NET0131  & ~\de_m0_arb_st_reg/NET0131  ;
  assign n2948 = ~n2838 & n2947 ;
  assign n2949 = ~n2946 & ~n2948 ;
  assign n2950 = n2935 & ~n2949 ;
  assign n2951 = ~n2944 & n2950 ;
  assign n2952 = n2943 & ~n2951 ;
  assign n2953 = \ahb_mst0_mx_cmd_st_reg[0]/NET0131  & \ahb_mst0_mx_cmd_st_reg[1]/NET0131  ;
  assign n2954 = ~n2838 & ~n2953 ;
  assign n2955 = ~n2919 & ~n2954 ;
  assign n2956 = ~\ch_sel_arb_chcsr_reg_reg[2]/NET0131  & ~\de_m0_arb_st_reg/NET0131  ;
  assign n2957 = ~n2955 & n2956 ;
  assign n2958 = \de_m0_arb_st_reg/NET0131  & ~n2835 ;
  assign n2959 = ~\ahb_mst0_mx_cmd_st_reg[0]/NET0131  & ~\ch_sel_arb_chcsr_reg_reg[1]/NET0131  ;
  assign n2960 = n2958 & n2959 ;
  assign n2961 = \ahb_mst0_mx_cmd_st_reg[1]/NET0131  & \h0grant_pad  ;
  assign n2962 = ~\h0resp[0]_pad  & ~\h0resp[1]_pad  ;
  assign n2963 = n2961 & n2962 ;
  assign n2964 = ~n2960 & n2963 ;
  assign n2965 = ~n2957 & n2964 ;
  assign n2966 = ~\ahb_mst0_mx_cmd_st_reg[0]/NET0131  & n2935 ;
  assign n2967 = ~n2944 & n2966 ;
  assign n2968 = ~n2965 & ~n2967 ;
  assign n2969 = \ch_sel_dma_rrarb1_state_reg[0]/NET0131  & \ch_sel_dma_rrarb1_state_reg[2]/NET0131  ;
  assign n2970 = \ctl_rf_c4_rf_ch_en_reg/NET0131  & ~\ctl_rf_c4_rf_chabt_reg/NET0131  ;
  assign n2971 = \ctl_rf_dmacen_reg/NET0131  & n2970 ;
  assign n2972 = ~\ctl_rf_c4_rf_mode_reg/NET0131  & n2971 ;
  assign n2973 = \ch_sel_fix_pri_sel_reg[0]/NET0131  & ~\ch_sel_fix_pri_sel_reg[1]/NET0131  ;
  assign n2974 = \ch_sel_dma_rrarb1_state_reg[0]/NET0131  & n2973 ;
  assign n2975 = ~\ch_sel_fix_pri_sel_reg[0]/NET0131  & \ch_sel_fix_pri_sel_reg[1]/NET0131  ;
  assign n2976 = \ch_sel_dma_rrarb2_state_reg[0]/NET0131  & n2975 ;
  assign n2977 = ~n2974 & ~n2976 ;
  assign n2978 = ~\ch_sel_fix_pri_sel_reg[0]/NET0131  & ~\ch_sel_fix_pri_sel_reg[1]/NET0131  ;
  assign n2979 = \ch_sel_dma_rrarb0_state_reg[0]/NET0131  & n2978 ;
  assign n2980 = \ch_sel_fix_pri_sel_reg[0]/NET0131  & \ch_sel_fix_pri_sel_reg[1]/NET0131  ;
  assign n2981 = \ch_sel_dma_rrarb3_state_reg[0]/NET0131  & n2980 ;
  assign n2982 = ~n2979 & ~n2981 ;
  assign n2983 = n2977 & n2982 ;
  assign n2984 = \de_de_st_reg[5]/NET0131  & n2983 ;
  assign n2985 = \ch_sel_dma_rrarb2_state_reg[1]/NET0131  & n2975 ;
  assign n2986 = \ch_sel_dma_rrarb3_state_reg[1]/NET0131  & n2980 ;
  assign n2987 = ~n2985 & ~n2986 ;
  assign n2988 = \ch_sel_dma_rrarb0_state_reg[1]/NET0131  & n2978 ;
  assign n2989 = \ch_sel_dma_rrarb1_state_reg[1]/NET0131  & n2973 ;
  assign n2990 = ~n2988 & ~n2989 ;
  assign n2991 = n2987 & n2990 ;
  assign n2992 = \ch_sel_dma_rrarb2_state_reg[2]/NET0131  & n2975 ;
  assign n2993 = \ch_sel_dma_rrarb3_state_reg[2]/NET0131  & n2980 ;
  assign n2994 = ~n2992 & ~n2993 ;
  assign n2995 = \ch_sel_dma_rrarb0_state_reg[2]/NET0131  & n2978 ;
  assign n2996 = \ch_sel_dma_rrarb1_state_reg[2]/NET0131  & n2973 ;
  assign n2997 = ~n2995 & ~n2996 ;
  assign n2998 = n2994 & n2997 ;
  assign n2999 = n2991 & ~n2998 ;
  assign n3000 = n2984 & n2999 ;
  assign n3001 = ~\ch_sel_dma_reqd1_reg[4]/NET0131  & ~\ctl_rf_sync_reg[4]/NET0131  ;
  assign n3002 = ~\ch_sel_dma_reqd2_reg[4]/NET0131  & \ctl_rf_sync_reg[4]/NET0131  ;
  assign n3003 = ~n3001 & ~n3002 ;
  assign n3004 = ~\dma_ack[4]_pad  & n3003 ;
  assign n3005 = n2971 & n3004 ;
  assign n3006 = ~n3000 & n3005 ;
  assign n3007 = ~n2972 & ~n3006 ;
  assign n3008 = \ctl_rf_c6_rf_ch_en_reg/NET0131  & ~\ctl_rf_c6_rf_chabt_reg/NET0131  ;
  assign n3009 = \ctl_rf_dmacen_reg/NET0131  & n3008 ;
  assign n3010 = ~\ctl_rf_c6_rf_mode_reg/NET0131  & n3009 ;
  assign n3011 = ~n2991 & ~n2998 ;
  assign n3012 = n2984 & n3011 ;
  assign n3013 = ~\ch_sel_dma_reqd1_reg[6]/NET0131  & ~\ctl_rf_sync_reg[6]/NET0131  ;
  assign n3014 = ~\ch_sel_dma_reqd2_reg[6]/NET0131  & \ctl_rf_sync_reg[6]/NET0131  ;
  assign n3015 = ~n3013 & ~n3014 ;
  assign n3016 = ~\dma_ack[6]_pad  & n3015 ;
  assign n3017 = n3009 & n3016 ;
  assign n3018 = ~n3012 & n3017 ;
  assign n3019 = ~n3010 & ~n3018 ;
  assign n3020 = n3007 & n3019 ;
  assign n3021 = \ctl_rf_c3_rf_ch_en_reg/NET0131  & ~\ctl_rf_c3_rf_chabt_reg/NET0131  ;
  assign n3022 = \ctl_rf_dmacen_reg/NET0131  & n3021 ;
  assign n3023 = ~\ctl_rf_c3_rf_mode_reg/NET0131  & n3022 ;
  assign n3024 = ~n2991 & n2998 ;
  assign n3025 = \de_de_st_reg[5]/NET0131  & ~n2983 ;
  assign n3026 = n3024 & n3025 ;
  assign n3027 = ~\ch_sel_dma_reqd1_reg[3]/NET0131  & ~\ctl_rf_sync_reg[3]/NET0131  ;
  assign n3028 = ~\ch_sel_dma_reqd2_reg[3]/P0001  & \ctl_rf_sync_reg[3]/NET0131  ;
  assign n3029 = ~n3027 & ~n3028 ;
  assign n3030 = ~\dma_ack[3]_pad  & n3029 ;
  assign n3031 = n3022 & n3030 ;
  assign n3032 = ~n3026 & n3031 ;
  assign n3033 = ~n3023 & ~n3032 ;
  assign n3034 = \ctl_rf_c5_rf_ch_en_reg/NET0131  & ~\ctl_rf_c5_rf_chabt_reg/NET0131  ;
  assign n3035 = \ctl_rf_dmacen_reg/NET0131  & n3034 ;
  assign n3036 = ~\ctl_rf_c5_rf_mode_reg/NET0131  & n3035 ;
  assign n3037 = n2999 & n3025 ;
  assign n3038 = ~\ch_sel_dma_reqd1_reg[5]/NET0131  & ~\ctl_rf_sync_reg[5]/NET0131  ;
  assign n3039 = ~\ch_sel_dma_reqd2_reg[5]/NET0131  & \ctl_rf_sync_reg[5]/NET0131  ;
  assign n3040 = ~n3038 & ~n3039 ;
  assign n3041 = ~\dma_ack[5]_pad  & n3040 ;
  assign n3042 = n3035 & n3041 ;
  assign n3043 = ~n3037 & n3042 ;
  assign n3044 = ~n3036 & ~n3043 ;
  assign n3045 = n3033 & n3044 ;
  assign n3046 = n3020 & n3045 ;
  assign n3047 = \ctl_rf_c0_rf_ch_en_reg/NET0131  & ~\ctl_rf_c0_rf_chabt_reg/NET0131  ;
  assign n3048 = \ctl_rf_dmacen_reg/NET0131  & n3047 ;
  assign n3049 = ~\ctl_rf_c0_rf_mode_reg/NET0131  & n3048 ;
  assign n3050 = n2991 & n2998 ;
  assign n3051 = n2984 & n3050 ;
  assign n3052 = ~\ch_sel_dma_reqd1_reg[0]/NET0131  & ~\ctl_rf_sync_reg[0]/NET0131  ;
  assign n3053 = ~\ch_sel_dma_reqd2_reg[0]/NET0131  & \ctl_rf_sync_reg[0]/NET0131  ;
  assign n3054 = ~n3052 & ~n3053 ;
  assign n3055 = ~\dma_ack[0]_pad  & n3054 ;
  assign n3056 = n3048 & n3055 ;
  assign n3057 = ~n3051 & n3056 ;
  assign n3058 = ~n3049 & ~n3057 ;
  assign n3059 = \ctl_rf_c2_rf_ch_en_reg/NET0131  & ~\ctl_rf_c2_rf_chabt_reg/NET0131  ;
  assign n3060 = \ctl_rf_dmacen_reg/NET0131  & n3059 ;
  assign n3061 = ~\ctl_rf_c2_rf_mode_reg/NET0131  & n3060 ;
  assign n3062 = n2984 & n3024 ;
  assign n3063 = ~\ch_sel_dma_reqd1_reg[2]/NET0131  & ~\ctl_rf_sync_reg[2]/NET0131  ;
  assign n3064 = ~\ch_sel_dma_reqd2_reg[2]/P0001  & \ctl_rf_sync_reg[2]/NET0131  ;
  assign n3065 = ~n3063 & ~n3064 ;
  assign n3066 = ~\dma_ack[2]_pad  & n3065 ;
  assign n3067 = n3060 & n3066 ;
  assign n3068 = ~n3062 & n3067 ;
  assign n3069 = ~n3061 & ~n3068 ;
  assign n3070 = n3058 & n3069 ;
  assign n3071 = \ctl_rf_c1_rf_ch_en_reg/NET0131  & ~\ctl_rf_c1_rf_chabt_reg/NET0131  ;
  assign n3072 = \ctl_rf_dmacen_reg/NET0131  & n3071 ;
  assign n3073 = ~\ctl_rf_c1_rf_mode_reg/NET0131  & n3072 ;
  assign n3074 = n3025 & n3050 ;
  assign n3075 = ~\ch_sel_dma_reqd1_reg[1]/NET0131  & ~\ctl_rf_sync_reg[1]/NET0131  ;
  assign n3076 = ~\ch_sel_dma_reqd2_reg[1]/P0001  & \ctl_rf_sync_reg[1]/NET0131  ;
  assign n3077 = ~n3075 & ~n3076 ;
  assign n3078 = ~\dma_ack[1]_pad  & n3077 ;
  assign n3079 = n3072 & n3078 ;
  assign n3080 = ~n3074 & n3079 ;
  assign n3081 = ~n3073 & ~n3080 ;
  assign n3082 = \ctl_rf_c7_rf_ch_en_reg/NET0131  & ~\ctl_rf_c7_rf_chabt_reg/NET0131  ;
  assign n3083 = \ctl_rf_dmacen_reg/NET0131  & n3082 ;
  assign n3084 = ~\ctl_rf_c7_rf_mode_reg/NET0131  & n3083 ;
  assign n3085 = n3011 & n3025 ;
  assign n3086 = ~\ch_sel_dma_reqd1_reg[7]/NET0131  & ~\ctl_rf_sync_reg[7]/NET0131  ;
  assign n3087 = ~\ch_sel_dma_reqd2_reg[7]/NET0131  & \ctl_rf_sync_reg[7]/NET0131  ;
  assign n3088 = ~n3086 & ~n3087 ;
  assign n3089 = ~\dma_ack[7]_pad  & n3088 ;
  assign n3090 = n3083 & n3089 ;
  assign n3091 = ~n3085 & n3090 ;
  assign n3092 = ~n3084 & ~n3091 ;
  assign n3093 = n3081 & n3092 ;
  assign n3094 = n3070 & n3093 ;
  assign n3095 = n3046 & n3094 ;
  assign n3096 = ~\ch_sel_vld_req_any_d1_reg/NET0131  & \de_de_st_reg[0]/NET0131  ;
  assign n3097 = ~n3095 & n3096 ;
  assign n3098 = ~\ctl_rf_c4_rf_chabt_reg/NET0131  & ~\ctl_rf_c5_rf_chabt_reg/NET0131  ;
  assign n3099 = ~\ctl_rf_c6_rf_chabt_reg/NET0131  & ~\ctl_rf_c7_rf_chabt_reg/NET0131  ;
  assign n3100 = n3098 & n3099 ;
  assign n3101 = ~\ctl_rf_c0_rf_chabt_reg/NET0131  & ~\ctl_rf_c1_rf_chabt_reg/NET0131  ;
  assign n3102 = ~\ctl_rf_c2_rf_chabt_reg/NET0131  & ~\ctl_rf_c3_rf_chabt_reg/NET0131  ;
  assign n3103 = n3101 & n3102 ;
  assign n3104 = n3100 & n3103 ;
  assign n3105 = \de_de_st_reg[0]/NET0131  & ~n3104 ;
  assign n3106 = ~\ch_sel_de_stup_d1_reg/NET0131  & ~n3105 ;
  assign n3107 = ~n3097 & n3106 ;
  assign n3108 = n2969 & n3107 ;
  assign n3109 = \ctl_rf_c1_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c1_rf_chpri_reg[1]/NET0131  ;
  assign n3110 = ~n3081 & n3109 ;
  assign n3111 = \ctl_rf_c0_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c0_rf_chpri_reg[1]/NET0131  ;
  assign n3112 = ~n3058 & n3111 ;
  assign n3113 = n3110 & ~n3112 ;
  assign n3114 = \ctl_rf_c7_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c7_rf_chpri_reg[1]/NET0131  ;
  assign n3115 = ~n3092 & n3114 ;
  assign n3116 = ~n3113 & ~n3115 ;
  assign n3117 = \ctl_rf_c3_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c3_rf_chpri_reg[1]/NET0131  ;
  assign n3118 = ~n3033 & n3117 ;
  assign n3119 = \ctl_rf_c2_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c2_rf_chpri_reg[1]/NET0131  ;
  assign n3120 = ~n3069 & n3119 ;
  assign n3121 = ~n3112 & ~n3120 ;
  assign n3122 = n3118 & n3121 ;
  assign n3123 = n3116 & ~n3122 ;
  assign n3124 = \ctl_rf_c4_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c4_rf_chpri_reg[1]/NET0131  ;
  assign n3125 = ~n3007 & n3124 ;
  assign n3126 = n3121 & ~n3125 ;
  assign n3127 = n3123 & ~n3126 ;
  assign n3128 = \ctl_rf_c6_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c6_rf_chpri_reg[1]/NET0131  ;
  assign n3129 = ~n3019 & n3128 ;
  assign n3130 = ~\ch_sel_dma_rrarb1_state_reg[1]/NET0131  & ~n3129 ;
  assign n3131 = n2969 & n3130 ;
  assign n3132 = ~n3127 & n3131 ;
  assign n3133 = ~n3108 & ~n3132 ;
  assign n3134 = ~\ch_sel_dma_rrarb1_state_reg[0]/NET0131  & ~\ch_sel_dma_rrarb1_state_reg[2]/NET0131  ;
  assign n3135 = \ch_sel_dma_rrarb1_state_reg[1]/NET0131  & n3134 ;
  assign n3136 = ~n3106 & n3135 ;
  assign n3137 = n3096 & n3135 ;
  assign n3138 = ~n3095 & n3137 ;
  assign n3139 = ~n3136 & ~n3138 ;
  assign n3140 = \ctl_rf_c5_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c5_rf_chpri_reg[1]/NET0131  ;
  assign n3141 = ~n3044 & n3140 ;
  assign n3142 = ~n3118 & ~n3141 ;
  assign n3143 = n3116 & n3142 ;
  assign n3144 = n3129 & ~n3141 ;
  assign n3145 = ~n3125 & ~n3144 ;
  assign n3146 = ~n3118 & ~n3145 ;
  assign n3147 = ~n3143 & ~n3146 ;
  assign n3148 = ~n3139 & n3147 ;
  assign n3149 = ~n3125 & n3141 ;
  assign n3150 = ~n3118 & ~n3149 ;
  assign n3151 = ~n3120 & ~n3150 ;
  assign n3152 = ~n3112 & ~n3129 ;
  assign n3153 = n3115 & ~n3129 ;
  assign n3154 = ~n3152 & ~n3153 ;
  assign n3155 = ~n3120 & ~n3125 ;
  assign n3156 = ~n3154 & n3155 ;
  assign n3157 = ~n3151 & ~n3156 ;
  assign n3158 = ~n3107 & n3157 ;
  assign n3159 = \ch_sel_dma_rrarb1_state_reg[0]/NET0131  & ~\ch_sel_dma_rrarb1_state_reg[2]/NET0131  ;
  assign n3160 = ~\ch_sel_dma_rrarb1_state_reg[1]/NET0131  & n3159 ;
  assign n3161 = ~n3158 & n3160 ;
  assign n3162 = ~n3148 & ~n3161 ;
  assign n3163 = n3133 & n3162 ;
  assign n3164 = n3121 & ~n3150 ;
  assign n3165 = n3116 & ~n3164 ;
  assign n3166 = \ch_sel_dma_rrarb1_state_reg[1]/NET0131  & ~n3165 ;
  assign n3167 = ~n3115 & ~n3141 ;
  assign n3168 = ~n3113 & n3167 ;
  assign n3169 = ~n3122 & n3168 ;
  assign n3170 = ~\ch_sel_dma_rrarb1_state_reg[1]/NET0131  & ~n3144 ;
  assign n3171 = ~n3169 & n3170 ;
  assign n3172 = ~n3166 & ~n3171 ;
  assign n3173 = ~\ch_sel_dma_rrarb1_state_reg[0]/NET0131  & \ch_sel_dma_rrarb1_state_reg[2]/NET0131  ;
  assign n3174 = ~n3106 & n3173 ;
  assign n3175 = n3096 & n3173 ;
  assign n3176 = ~n3095 & n3175 ;
  assign n3177 = ~n3174 & ~n3176 ;
  assign n3178 = ~n3172 & ~n3177 ;
  assign n3179 = \ch_sel_dma_rrarb1_state_reg[1]/NET0131  & n3159 ;
  assign n3180 = ~n3110 & n3120 ;
  assign n3181 = ~n3125 & n3152 ;
  assign n3182 = ~n3180 & n3181 ;
  assign n3183 = ~n3125 & n3153 ;
  assign n3184 = ~n3149 & ~n3183 ;
  assign n3185 = ~n3182 & n3184 ;
  assign n3186 = ~n3107 & n3185 ;
  assign n3187 = n3179 & ~n3186 ;
  assign n3188 = ~\ch_sel_dma_rrarb1_state_reg[1]/NET0131  & ~n3106 ;
  assign n3189 = ~\ch_sel_dma_rrarb1_state_reg[1]/NET0131  & n3096 ;
  assign n3190 = ~n3095 & n3189 ;
  assign n3191 = ~n3188 & ~n3190 ;
  assign n3192 = ~n3110 & ~n3118 ;
  assign n3193 = ~n3149 & n3192 ;
  assign n3194 = ~n3183 & n3193 ;
  assign n3195 = n3134 & ~n3180 ;
  assign n3196 = ~n3194 & n3195 ;
  assign n3197 = ~n3191 & n3196 ;
  assign n3198 = ~n3113 & ~n3121 ;
  assign n3199 = ~n3113 & ~n3118 ;
  assign n3200 = ~n3145 & n3199 ;
  assign n3201 = ~n3198 & ~n3200 ;
  assign n3202 = \ch_sel_dma_rrarb1_state_reg[1]/NET0131  & n2969 ;
  assign n3203 = n3201 & n3202 ;
  assign n3204 = ~n3197 & ~n3203 ;
  assign n3205 = ~n3187 & n3204 ;
  assign n3206 = ~n3178 & n3205 ;
  assign n3207 = n3163 & n3206 ;
  assign n3208 = ~\ch_sel_dma_rrarb3_state_reg[1]/NET0131  & ~n3106 ;
  assign n3209 = ~\ch_sel_dma_rrarb3_state_reg[1]/NET0131  & n3096 ;
  assign n3210 = ~n3095 & n3209 ;
  assign n3211 = ~n3208 & ~n3210 ;
  assign n3212 = ~\ch_sel_dma_rrarb3_state_reg[0]/NET0131  & \ch_sel_dma_rrarb3_state_reg[2]/NET0131  ;
  assign n3213 = ~n3211 & n3212 ;
  assign n3214 = \ctl_rf_c5_rf_chpri_reg[0]/NET0131  & \ctl_rf_c5_rf_chpri_reg[1]/NET0131  ;
  assign n3215 = ~n3044 & n3214 ;
  assign n3216 = \ctl_rf_c6_rf_chpri_reg[0]/NET0131  & \ctl_rf_c6_rf_chpri_reg[1]/NET0131  ;
  assign n3217 = ~n3019 & n3216 ;
  assign n3218 = \ctl_rf_c7_rf_chpri_reg[0]/NET0131  & \ctl_rf_c7_rf_chpri_reg[1]/NET0131  ;
  assign n3219 = ~n3092 & n3218 ;
  assign n3220 = ~n3217 & n3219 ;
  assign n3221 = ~n3215 & ~n3220 ;
  assign n3222 = \ctl_rf_c1_rf_chpri_reg[0]/NET0131  & \ctl_rf_c1_rf_chpri_reg[1]/NET0131  ;
  assign n3223 = ~n3081 & n3222 ;
  assign n3224 = \ctl_rf_c3_rf_chpri_reg[0]/NET0131  & \ctl_rf_c3_rf_chpri_reg[1]/NET0131  ;
  assign n3225 = ~n3033 & n3224 ;
  assign n3226 = ~n3223 & ~n3225 ;
  assign n3227 = \ctl_rf_c2_rf_chpri_reg[0]/NET0131  & \ctl_rf_c2_rf_chpri_reg[1]/NET0131  ;
  assign n3228 = ~n3069 & n3227 ;
  assign n3229 = ~n3223 & n3228 ;
  assign n3230 = \ctl_rf_c0_rf_chpri_reg[0]/NET0131  & \ctl_rf_c0_rf_chpri_reg[1]/NET0131  ;
  assign n3231 = ~n3058 & n3230 ;
  assign n3232 = ~n3217 & ~n3231 ;
  assign n3233 = ~n3229 & n3232 ;
  assign n3234 = ~n3226 & n3233 ;
  assign n3235 = n3221 & ~n3234 ;
  assign n3236 = n3213 & ~n3235 ;
  assign n3237 = \ch_sel_dma_rrarb3_state_reg[0]/NET0131  & \ch_sel_dma_rrarb3_state_reg[2]/NET0131  ;
  assign n3238 = n3106 & n3237 ;
  assign n3239 = ~n3097 & n3238 ;
  assign n3240 = ~n3236 & ~n3239 ;
  assign n3241 = \ctl_rf_c4_rf_chpri_reg[0]/NET0131  & \ctl_rf_c4_rf_chpri_reg[1]/NET0131  ;
  assign n3242 = ~n3007 & n3241 ;
  assign n3243 = n3215 & ~n3242 ;
  assign n3244 = ~n3225 & ~n3243 ;
  assign n3245 = ~n3228 & ~n3244 ;
  assign n3246 = ~n3228 & ~n3242 ;
  assign n3247 = ~n3220 & ~n3232 ;
  assign n3248 = n3246 & ~n3247 ;
  assign n3249 = ~n3245 & ~n3248 ;
  assign n3250 = ~n3107 & n3249 ;
  assign n3251 = \ch_sel_dma_rrarb3_state_reg[0]/NET0131  & ~\ch_sel_dma_rrarb3_state_reg[2]/NET0131  ;
  assign n3252 = ~\ch_sel_dma_rrarb3_state_reg[1]/NET0131  & n3251 ;
  assign n3253 = ~n3250 & n3252 ;
  assign n3254 = \ch_sel_dma_rrarb3_state_reg[1]/NET0131  & n3251 ;
  assign n3255 = ~n3221 & ~n3242 ;
  assign n3256 = n3233 & ~n3242 ;
  assign n3257 = ~n3255 & ~n3256 ;
  assign n3258 = ~n3107 & n3257 ;
  assign n3259 = n3254 & ~n3258 ;
  assign n3260 = ~n3253 & ~n3259 ;
  assign n3261 = n3240 & n3260 ;
  assign n3262 = ~\ch_sel_dma_rrarb3_state_reg[0]/NET0131  & ~\ch_sel_dma_rrarb3_state_reg[2]/NET0131  ;
  assign n3263 = ~n3226 & ~n3229 ;
  assign n3264 = ~n3221 & n3246 ;
  assign n3265 = ~n3263 & ~n3264 ;
  assign n3266 = ~n3211 & ~n3265 ;
  assign n3267 = n3262 & n3266 ;
  assign n3268 = ~n3220 & ~n3223 ;
  assign n3269 = ~n3242 & ~n3268 ;
  assign n3270 = ~n3247 & n3269 ;
  assign n3271 = n3244 & ~n3270 ;
  assign n3272 = \ch_sel_dma_rrarb3_state_reg[1]/NET0131  & ~n3106 ;
  assign n3273 = \ch_sel_dma_rrarb3_state_reg[1]/NET0131  & n3096 ;
  assign n3274 = ~n3095 & n3273 ;
  assign n3275 = ~n3272 & ~n3274 ;
  assign n3276 = n3262 & ~n3275 ;
  assign n3277 = ~n3271 & n3276 ;
  assign n3278 = ~n3267 & ~n3277 ;
  assign n3279 = \ch_sel_dma_rrarb3_state_reg[1]/NET0131  & \ctl_rf_c5_rf_chpri_reg[1]/NET0131  ;
  assign n3280 = \ctl_rf_c5_rf_chpri_reg[0]/NET0131  & n3279 ;
  assign n3281 = ~n3044 & n3280 ;
  assign n3282 = n3217 & ~n3281 ;
  assign n3283 = n3246 & ~n3282 ;
  assign n3284 = ~n3231 & n3283 ;
  assign n3285 = ~\ch_sel_dma_rrarb3_state_reg[1]/NET0131  & \ctl_rf_c6_rf_chpri_reg[1]/NET0131  ;
  assign n3286 = \ctl_rf_c6_rf_chpri_reg[0]/NET0131  & n3285 ;
  assign n3287 = ~n3019 & n3286 ;
  assign n3288 = ~n3231 & ~n3287 ;
  assign n3289 = n3263 & n3288 ;
  assign n3290 = ~n3284 & ~n3289 ;
  assign n3291 = ~\ch_sel_dma_rrarb3_state_reg[1]/NET0131  & n3220 ;
  assign n3292 = n3290 & ~n3291 ;
  assign n3293 = n3237 & ~n3292 ;
  assign n3294 = n3226 & ~n3243 ;
  assign n3295 = ~n3229 & ~n3294 ;
  assign n3296 = ~n3231 & n3295 ;
  assign n3297 = ~n3219 & ~n3296 ;
  assign n3298 = n3212 & ~n3275 ;
  assign n3299 = ~n3297 & n3298 ;
  assign n3300 = ~n3293 & ~n3299 ;
  assign n3301 = n3278 & n3300 ;
  assign n3302 = n3261 & n3301 ;
  assign n3303 = ~\ch_sel_dma_rrarb0_state_reg[0]/NET0131  & ~\ch_sel_dma_rrarb0_state_reg[2]/NET0131  ;
  assign n3304 = ~\ch_sel_dma_rrarb0_state_reg[1]/NET0131  & n3303 ;
  assign n3305 = ~\ctl_rf_c1_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c1_rf_chpri_reg[1]/NET0131  ;
  assign n3306 = ~n3081 & n3305 ;
  assign n3307 = n3304 & n3306 ;
  assign n3308 = ~\ctl_rf_c3_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c3_rf_chpri_reg[1]/NET0131  ;
  assign n3309 = ~n3033 & n3308 ;
  assign n3310 = ~\ctl_rf_c4_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c4_rf_chpri_reg[1]/NET0131  ;
  assign n3311 = ~n3007 & n3310 ;
  assign n3312 = ~n3309 & n3311 ;
  assign n3313 = ~\ctl_rf_c6_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c6_rf_chpri_reg[1]/NET0131  ;
  assign n3314 = ~n3019 & n3313 ;
  assign n3315 = ~\ctl_rf_c7_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c7_rf_chpri_reg[1]/NET0131  ;
  assign n3316 = ~n3092 & n3315 ;
  assign n3317 = ~n3314 & n3316 ;
  assign n3318 = ~\ctl_rf_c5_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c5_rf_chpri_reg[1]/NET0131  ;
  assign n3319 = ~n3044 & n3318 ;
  assign n3320 = ~n3309 & ~n3319 ;
  assign n3321 = ~n3317 & n3320 ;
  assign n3322 = ~n3312 & ~n3321 ;
  assign n3323 = ~\ctl_rf_c2_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c2_rf_chpri_reg[1]/NET0131  ;
  assign n3324 = ~n3069 & n3323 ;
  assign n3325 = n3304 & ~n3324 ;
  assign n3326 = n3322 & n3325 ;
  assign n3327 = ~n3307 & ~n3326 ;
  assign n3328 = ~n3312 & ~n3320 ;
  assign n3329 = ~\ctl_rf_c0_rf_chpri_reg[0]/NET0131  & ~\ctl_rf_c0_rf_chpri_reg[1]/NET0131  ;
  assign n3330 = ~n3058 & n3329 ;
  assign n3331 = ~n3324 & ~n3330 ;
  assign n3332 = \ch_sel_dma_rrarb0_state_reg[2]/NET0131  & ~n3331 ;
  assign n3333 = n3328 & ~n3332 ;
  assign n3334 = ~n3311 & ~n3314 ;
  assign n3335 = ~\ch_sel_dma_rrarb0_state_reg[2]/NET0131  & ~n3334 ;
  assign n3336 = n3306 & ~n3330 ;
  assign n3337 = ~n3316 & ~n3336 ;
  assign n3338 = ~n3335 & ~n3337 ;
  assign n3339 = ~n3333 & ~n3338 ;
  assign n3340 = ~\ch_sel_dma_rrarb0_state_reg[0]/NET0131  & \ch_sel_dma_rrarb0_state_reg[1]/NET0131  ;
  assign n3341 = ~n3339 & n3340 ;
  assign n3342 = n3327 & ~n3341 ;
  assign n3343 = ~n3107 & ~n3342 ;
  assign n3344 = \ch_sel_dma_rrarb0_state_reg[0]/NET0131  & ~\ch_sel_dma_rrarb0_state_reg[2]/NET0131  ;
  assign n3345 = ~\ch_sel_dma_rrarb0_state_reg[1]/NET0131  & n3344 ;
  assign n3346 = ~n3316 & n3330 ;
  assign n3347 = n3334 & ~n3346 ;
  assign n3348 = ~n3328 & ~n3347 ;
  assign n3349 = ~n3324 & ~n3348 ;
  assign n3350 = ~n3107 & ~n3349 ;
  assign n3351 = n3345 & ~n3350 ;
  assign n3352 = \ch_sel_dma_rrarb0_state_reg[1]/NET0131  & n3344 ;
  assign n3353 = ~n3317 & ~n3319 ;
  assign n3354 = ~n3311 & ~n3353 ;
  assign n3355 = ~n3331 & ~n3336 ;
  assign n3356 = n3334 & ~n3355 ;
  assign n3357 = ~n3354 & ~n3356 ;
  assign n3358 = ~n3107 & n3357 ;
  assign n3359 = n3352 & ~n3358 ;
  assign n3360 = ~n3351 & ~n3359 ;
  assign n3361 = ~n3314 & n3336 ;
  assign n3362 = n3309 & ~n3314 ;
  assign n3363 = n3331 & n3362 ;
  assign n3364 = ~n3361 & ~n3363 ;
  assign n3365 = n3353 & n3364 ;
  assign n3366 = ~\ch_sel_dma_rrarb0_state_reg[1]/NET0131  & \ch_sel_dma_rrarb0_state_reg[2]/NET0131  ;
  assign n3367 = ~\ch_sel_dma_rrarb0_state_reg[0]/NET0131  & n3366 ;
  assign n3368 = ~n3106 & n3367 ;
  assign n3369 = n3096 & n3367 ;
  assign n3370 = ~n3095 & n3369 ;
  assign n3371 = ~n3368 & ~n3370 ;
  assign n3372 = ~n3365 & ~n3371 ;
  assign n3373 = \ch_sel_dma_rrarb0_state_reg[0]/NET0131  & \ch_sel_dma_rrarb0_state_reg[2]/NET0131  ;
  assign n3374 = n3107 & n3373 ;
  assign n3375 = n3320 & ~n3336 ;
  assign n3376 = \ch_sel_dma_rrarb0_state_reg[1]/NET0131  & ~n3375 ;
  assign n3377 = n3314 & ~n3376 ;
  assign n3378 = ~n3312 & n3331 ;
  assign n3379 = ~\ch_sel_dma_rrarb0_state_reg[1]/NET0131  & ~\ctl_rf_c7_rf_chpri_reg[1]/NET0131  ;
  assign n3380 = ~\ctl_rf_c7_rf_chpri_reg[0]/NET0131  & n3379 ;
  assign n3381 = ~n3092 & n3380 ;
  assign n3382 = ~n3336 & ~n3381 ;
  assign n3383 = ~n3378 & n3382 ;
  assign n3384 = n3373 & ~n3383 ;
  assign n3385 = ~n3377 & n3384 ;
  assign n3386 = ~n3374 & ~n3385 ;
  assign n3387 = ~n3372 & n3386 ;
  assign n3388 = n3360 & n3387 ;
  assign n3389 = ~n3343 & n3388 ;
  assign n3390 = ~\ctl_rf_c3_rf_chpri_reg[0]/NET0131  & \ctl_rf_c3_rf_chpri_reg[1]/NET0131  ;
  assign n3391 = ~n3033 & n3390 ;
  assign n3392 = ~\ctl_rf_c1_rf_chpri_reg[0]/NET0131  & \ctl_rf_c1_rf_chpri_reg[1]/NET0131  ;
  assign n3393 = ~n3081 & n3392 ;
  assign n3394 = ~\ctl_rf_c0_rf_chpri_reg[0]/NET0131  & \ctl_rf_c0_rf_chpri_reg[1]/NET0131  ;
  assign n3395 = ~n3058 & n3394 ;
  assign n3396 = n3393 & ~n3395 ;
  assign n3397 = ~\ctl_rf_c5_rf_chpri_reg[0]/NET0131  & \ctl_rf_c5_rf_chpri_reg[1]/NET0131  ;
  assign n3398 = ~n3044 & n3397 ;
  assign n3399 = ~\ctl_rf_c7_rf_chpri_reg[0]/NET0131  & \ctl_rf_c7_rf_chpri_reg[1]/NET0131  ;
  assign n3400 = ~n3092 & n3399 ;
  assign n3401 = ~n3398 & ~n3400 ;
  assign n3402 = ~n3396 & n3401 ;
  assign n3403 = ~\ctl_rf_c4_rf_chpri_reg[0]/NET0131  & \ctl_rf_c4_rf_chpri_reg[1]/NET0131  ;
  assign n3404 = ~n3007 & n3403 ;
  assign n3405 = ~\ctl_rf_c6_rf_chpri_reg[0]/NET0131  & \ctl_rf_c6_rf_chpri_reg[1]/NET0131  ;
  assign n3406 = ~n3019 & n3405 ;
  assign n3407 = ~n3398 & n3406 ;
  assign n3408 = ~n3404 & ~n3407 ;
  assign n3409 = ~n3402 & n3408 ;
  assign n3410 = ~n3391 & ~n3409 ;
  assign n3411 = ~\ch_sel_dma_rrarb2_state_reg[0]/NET0131  & \ch_sel_dma_rrarb2_state_reg[1]/NET0131  ;
  assign n3412 = ~\ch_sel_dma_rrarb2_state_reg[2]/NET0131  & n3411 ;
  assign n3413 = ~n3106 & n3412 ;
  assign n3414 = n3096 & n3412 ;
  assign n3415 = ~n3095 & n3414 ;
  assign n3416 = ~n3413 & ~n3415 ;
  assign n3417 = ~n3410 & ~n3416 ;
  assign n3418 = ~\ch_sel_dma_rrarb2_state_reg[1]/NET0131  & ~\ch_sel_dma_rrarb2_state_reg[2]/NET0131  ;
  assign n3419 = \ch_sel_dma_rrarb2_state_reg[0]/NET0131  & ~n3418 ;
  assign n3420 = n3106 & n3419 ;
  assign n3421 = ~n3097 & n3420 ;
  assign n3422 = ~n3417 & ~n3421 ;
  assign n3423 = \ch_sel_dma_rrarb2_state_reg[0]/NET0131  & ~\ch_sel_dma_rrarb2_state_reg[2]/NET0131  ;
  assign n3424 = \ch_sel_dma_rrarb2_state_reg[1]/NET0131  & n3423 ;
  assign n3425 = n3398 & ~n3404 ;
  assign n3426 = ~n3404 & ~n3406 ;
  assign n3427 = n3400 & n3426 ;
  assign n3428 = ~n3425 & ~n3427 ;
  assign n3429 = ~\ctl_rf_c2_rf_chpri_reg[0]/NET0131  & \ctl_rf_c2_rf_chpri_reg[1]/NET0131  ;
  assign n3430 = ~n3069 & n3429 ;
  assign n3431 = ~n3395 & ~n3430 ;
  assign n3432 = ~n3396 & ~n3431 ;
  assign n3433 = n3426 & ~n3432 ;
  assign n3434 = n3428 & ~n3433 ;
  assign n3435 = n3424 & ~n3434 ;
  assign n3436 = ~n3391 & ~n3393 ;
  assign n3437 = ~n3432 & ~n3436 ;
  assign n3438 = ~n3404 & n3431 ;
  assign n3439 = ~n3407 & n3438 ;
  assign n3440 = ~n3437 & ~n3439 ;
  assign n3441 = \ch_sel_dma_rrarb2_state_reg[1]/NET0131  & \ch_sel_dma_rrarb2_state_reg[2]/NET0131  ;
  assign n3442 = \ch_sel_dma_rrarb2_state_reg[0]/NET0131  & n3441 ;
  assign n3443 = ~n3440 & n3442 ;
  assign n3444 = ~n3435 & ~n3443 ;
  assign n3445 = n3422 & n3444 ;
  assign n3446 = ~n3400 & n3432 ;
  assign n3447 = ~n3400 & ~n3425 ;
  assign n3448 = n3436 & n3447 ;
  assign n3449 = ~n3446 & ~n3448 ;
  assign n3450 = \ch_sel_dma_rrarb2_state_reg[2]/NET0131  & n3411 ;
  assign n3451 = ~n3106 & n3450 ;
  assign n3452 = n3096 & n3450 ;
  assign n3453 = ~n3095 & n3452 ;
  assign n3454 = ~n3451 & ~n3453 ;
  assign n3455 = n3449 & ~n3454 ;
  assign n3456 = ~n3400 & ~n3438 ;
  assign n3457 = ~n3437 & n3456 ;
  assign n3458 = ~\ch_sel_dma_rrarb2_state_reg[1]/NET0131  & \ch_sel_dma_rrarb2_state_reg[2]/NET0131  ;
  assign n3459 = \ch_sel_dma_rrarb2_state_reg[0]/NET0131  & n3458 ;
  assign n3460 = ~n3406 & n3459 ;
  assign n3461 = ~n3457 & n3460 ;
  assign n3462 = ~n3455 & ~n3461 ;
  assign n3463 = n3445 & n3462 ;
  assign n3464 = ~\ch_sel_dma_rrarb2_state_reg[0]/NET0131  & n3418 ;
  assign n3465 = n3393 & n3464 ;
  assign n3466 = ~n3391 & ~n3425 ;
  assign n3467 = ~n3427 & n3466 ;
  assign n3468 = ~n3430 & n3464 ;
  assign n3469 = ~n3467 & n3468 ;
  assign n3470 = ~n3465 & ~n3469 ;
  assign n3471 = n3401 & ~n3437 ;
  assign n3472 = ~\ch_sel_dma_rrarb2_state_reg[0]/NET0131  & n3458 ;
  assign n3473 = ~n3407 & n3472 ;
  assign n3474 = ~n3471 & n3473 ;
  assign n3475 = n3470 & ~n3474 ;
  assign n3476 = ~n3107 & ~n3475 ;
  assign n3477 = ~n3430 & ~n3467 ;
  assign n3478 = n3426 & n3431 ;
  assign n3479 = ~n3107 & ~n3478 ;
  assign n3480 = ~n3477 & n3479 ;
  assign n3481 = \ch_sel_dma_rrarb2_state_reg[0]/NET0131  & n3418 ;
  assign n3482 = ~n3480 & n3481 ;
  assign n3483 = ~n3476 & ~n3482 ;
  assign n3484 = n3463 & n3483 ;
  assign n3485 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \de_m1_arb_st_reg[1]/NET0131  ;
  assign n3486 = \ahb_mst0_m0_m1_diff_tx_reg/NET0131  & \ch_sel_arb_chcsr_reg_reg[1]/NET0131  ;
  assign n3487 = ~\de_m1_is_llp_reg/NET0131  & ~n3486 ;
  assign n3488 = n2816 & n3487 ;
  assign n3489 = \de_m1_is_llp_reg/NET0131  & ~n3486 ;
  assign n3490 = ~n2816 & n3489 ;
  assign n3491 = ~n3488 & ~n3490 ;
  assign n3492 = ~\de_m1_is_llp_reg/NET0131  & n3486 ;
  assign n3493 = ~n2816 & n3492 ;
  assign n3494 = \h1size[2]_pad  & ~n3493 ;
  assign n3495 = n3491 & n3494 ;
  assign n3496 = \ch_sel_arb_chcsr_reg_reg[10]/NET0131  & ~\de_m1_is_llp_reg/NET0131  ;
  assign n3497 = n3486 & n3496 ;
  assign n3498 = ~n2816 & n3497 ;
  assign n3499 = \ch_sel_arb_chcsr_reg_reg[13]/NET0131  & \ch_sel_arb_chcsr_reg_reg[2]/NET0131  ;
  assign n3500 = ~n2815 & n3499 ;
  assign n3501 = n3487 & n3500 ;
  assign n3502 = ~\de_m1_arb_st_reg[1]/NET0131  & ~n3501 ;
  assign n3503 = ~n3498 & n3502 ;
  assign n3504 = ~n3495 & n3503 ;
  assign n3505 = ~n3485 & ~n3504 ;
  assign n3506 = n2834 & ~n3505 ;
  assign n3507 = ~\h1size[2]_pad  & ~n2834 ;
  assign n3508 = ~n3506 & ~n3507 ;
  assign n3509 = n3118 & n3134 ;
  assign n3510 = ~n3110 & ~n3112 ;
  assign n3511 = ~n3115 & ~n3129 ;
  assign n3512 = ~n3510 & n3511 ;
  assign n3513 = ~n3125 & ~n3141 ;
  assign n3514 = n3134 & n3513 ;
  assign n3515 = ~n3512 & n3514 ;
  assign n3516 = ~n3509 & ~n3515 ;
  assign n3517 = ~n3107 & n3516 ;
  assign n3518 = \ch_sel_dma_rrarb1_state_reg[1]/NET0131  & ~n3517 ;
  assign n3519 = ~\ch_sel_dma_rrarb1_state_reg[0]/NET0131  & ~\ctl_rf_c7_rf_chpri_reg[1]/NET0131  ;
  assign n3520 = \ctl_rf_c7_rf_chpri_reg[0]/NET0131  & n3519 ;
  assign n3521 = ~n3092 & n3520 ;
  assign n3522 = \ch_sel_dma_rrarb1_state_reg[1]/NET0131  & n3521 ;
  assign n3523 = ~n3118 & ~n3120 ;
  assign n3524 = ~n3513 & n3523 ;
  assign n3525 = \ch_sel_dma_rrarb1_state_reg[1]/NET0131  & n3510 ;
  assign n3526 = ~n3524 & n3525 ;
  assign n3527 = ~n3522 & ~n3526 ;
  assign n3528 = n3510 & ~n3523 ;
  assign n3529 = n3511 & ~n3528 ;
  assign n3530 = ~\ch_sel_dma_rrarb1_state_reg[0]/NET0131  & ~n3141 ;
  assign n3531 = ~n3529 & n3530 ;
  assign n3532 = ~n3191 & n3531 ;
  assign n3533 = n3527 & ~n3532 ;
  assign n3534 = \ch_sel_dma_rrarb1_state_reg[2]/NET0131  & ~n3533 ;
  assign n3535 = n3179 & n3513 ;
  assign n3536 = ~n3512 & n3535 ;
  assign n3537 = ~n3511 & n3513 ;
  assign n3538 = n3523 & ~n3537 ;
  assign n3539 = ~\ch_sel_dma_rrarb1_state_reg[0]/NET0131  & ~\ctl_rf_c1_rf_chpri_reg[1]/NET0131  ;
  assign n3540 = \ctl_rf_c1_rf_chpri_reg[0]/NET0131  & n3539 ;
  assign n3541 = ~n3081 & n3540 ;
  assign n3542 = ~\ch_sel_dma_rrarb1_state_reg[2]/NET0131  & ~n3541 ;
  assign n3543 = ~n3538 & n3542 ;
  assign n3544 = n2969 & ~n3529 ;
  assign n3545 = ~n3543 & ~n3544 ;
  assign n3546 = ~n3191 & ~n3545 ;
  assign n3547 = ~n3536 & ~n3546 ;
  assign n3548 = ~n3534 & n3547 ;
  assign n3549 = ~n3518 & n3548 ;
  assign n3550 = ~n3391 & ~n3430 ;
  assign n3551 = ~n3398 & ~n3404 ;
  assign n3552 = ~n3400 & ~n3406 ;
  assign n3553 = n3551 & ~n3552 ;
  assign n3554 = n3550 & ~n3553 ;
  assign n3555 = ~\ch_sel_dma_rrarb2_state_reg[0]/NET0131  & \ctl_rf_c1_rf_chpri_reg[1]/NET0131  ;
  assign n3556 = ~\ctl_rf_c1_rf_chpri_reg[0]/NET0131  & n3555 ;
  assign n3557 = ~n3081 & n3556 ;
  assign n3558 = n3418 & ~n3557 ;
  assign n3559 = ~n3554 & n3558 ;
  assign n3560 = ~n3393 & ~n3395 ;
  assign n3561 = ~n3550 & n3560 ;
  assign n3562 = n3552 & ~n3561 ;
  assign n3563 = ~\ch_sel_dma_rrarb2_state_reg[0]/NET0131  & \ctl_rf_c5_rf_chpri_reg[1]/NET0131  ;
  assign n3564 = ~\ctl_rf_c5_rf_chpri_reg[0]/NET0131  & n3563 ;
  assign n3565 = ~n3044 & n3564 ;
  assign n3566 = n3458 & ~n3565 ;
  assign n3567 = ~n3562 & n3566 ;
  assign n3568 = ~n3559 & ~n3567 ;
  assign n3569 = ~n3107 & ~n3568 ;
  assign n3570 = n3552 & ~n3560 ;
  assign n3571 = n3423 & n3551 ;
  assign n3572 = ~n3570 & n3571 ;
  assign n3573 = \ch_sel_dma_rrarb2_state_reg[1]/NET0131  & n3572 ;
  assign n3574 = \ch_sel_dma_rrarb2_state_reg[1]/NET0131  & n3106 ;
  assign n3575 = ~n3097 & n3574 ;
  assign n3576 = ~n3573 & ~n3575 ;
  assign n3577 = n3391 & n3412 ;
  assign n3578 = n3412 & n3551 ;
  assign n3579 = ~n3570 & n3578 ;
  assign n3580 = ~n3577 & ~n3579 ;
  assign n3581 = n3550 & ~n3551 ;
  assign n3582 = n3441 & n3560 ;
  assign n3583 = ~n3581 & n3582 ;
  assign n3584 = n3399 & n3450 ;
  assign n3585 = ~n3092 & n3584 ;
  assign n3586 = ~n3583 & ~n3585 ;
  assign n3587 = n3580 & n3586 ;
  assign n3588 = n3576 & n3587 ;
  assign n3589 = ~n3569 & n3588 ;
  assign n3590 = ~\ch_sel_dma_rrarb3_state_reg[0]/NET0131  & \ctl_rf_c7_rf_chpri_reg[1]/NET0131  ;
  assign n3591 = \ctl_rf_c7_rf_chpri_reg[0]/NET0131  & n3590 ;
  assign n3592 = ~n3092 & n3591 ;
  assign n3593 = \ch_sel_dma_rrarb3_state_reg[1]/NET0131  & \ch_sel_dma_rrarb3_state_reg[2]/NET0131  ;
  assign n3594 = n3592 & n3593 ;
  assign n3595 = ~n3215 & ~n3242 ;
  assign n3596 = ~n3225 & ~n3228 ;
  assign n3597 = ~n3595 & n3596 ;
  assign n3598 = ~n3223 & ~n3231 ;
  assign n3599 = n3593 & n3598 ;
  assign n3600 = ~n3597 & n3599 ;
  assign n3601 = ~n3594 & ~n3600 ;
  assign n3602 = ~n3217 & ~n3219 ;
  assign n3603 = ~n3598 & n3602 ;
  assign n3604 = n3254 & n3595 ;
  assign n3605 = ~n3603 & n3604 ;
  assign n3606 = \ch_sel_dma_rrarb3_state_reg[1]/NET0131  & ~n3262 ;
  assign n3607 = n3106 & n3606 ;
  assign n3608 = ~n3097 & n3607 ;
  assign n3609 = ~n3605 & ~n3608 ;
  assign n3610 = n3601 & n3609 ;
  assign n3611 = n3595 & ~n3602 ;
  assign n3612 = n3596 & ~n3611 ;
  assign n3613 = ~\ch_sel_dma_rrarb3_state_reg[0]/NET0131  & \ctl_rf_c1_rf_chpri_reg[1]/NET0131  ;
  assign n3614 = \ctl_rf_c1_rf_chpri_reg[0]/NET0131  & n3613 ;
  assign n3615 = ~n3081 & n3614 ;
  assign n3616 = ~\ch_sel_dma_rrarb3_state_reg[1]/NET0131  & ~\ch_sel_dma_rrarb3_state_reg[2]/NET0131  ;
  assign n3617 = ~n3615 & n3616 ;
  assign n3618 = ~n3106 & n3617 ;
  assign n3619 = n3096 & n3617 ;
  assign n3620 = ~n3095 & n3619 ;
  assign n3621 = ~n3618 & ~n3620 ;
  assign n3622 = ~n3612 & ~n3621 ;
  assign n3623 = ~n3596 & n3598 ;
  assign n3624 = n3602 & ~n3623 ;
  assign n3625 = n3237 & ~n3624 ;
  assign n3626 = ~n3211 & n3625 ;
  assign n3627 = ~n3622 & ~n3626 ;
  assign n3628 = n3610 & n3627 ;
  assign n3629 = \ch_sel_dma_rrarb3_state_reg[1]/NET0131  & n3262 ;
  assign n3630 = n3595 & ~n3603 ;
  assign n3631 = ~n3106 & ~n3225 ;
  assign n3632 = n3096 & ~n3225 ;
  assign n3633 = ~n3095 & n3632 ;
  assign n3634 = ~n3631 & ~n3633 ;
  assign n3635 = ~n3630 & ~n3634 ;
  assign n3636 = n3629 & ~n3635 ;
  assign n3637 = n3212 & ~n3215 ;
  assign n3638 = ~n3624 & n3637 ;
  assign n3639 = ~n3211 & n3638 ;
  assign n3640 = ~n3636 & ~n3639 ;
  assign n3641 = n3628 & n3640 ;
  assign n3642 = \ch_sel_dma_rrarb1_state_reg[1]/NET0131  & ~n3521 ;
  assign n3643 = ~\ch_sel_dma_rrarb1_state_reg[0]/NET0131  & ~\ctl_rf_c5_rf_chpri_reg[1]/NET0131  ;
  assign n3644 = \ctl_rf_c5_rf_chpri_reg[0]/NET0131  & n3643 ;
  assign n3645 = ~n3044 & n3644 ;
  assign n3646 = n3511 & ~n3645 ;
  assign n3647 = ~n3642 & ~n3646 ;
  assign n3648 = n3510 & n3523 ;
  assign n3649 = ~n3647 & ~n3648 ;
  assign n3650 = ~n3107 & n3649 ;
  assign n3651 = \ch_sel_dma_rrarb1_state_reg[2]/NET0131  & ~n3650 ;
  assign n3652 = ~\ch_sel_dma_rrarb1_state_reg[1]/NET0131  & ~\ch_sel_dma_rrarb1_state_reg[2]/NET0131  ;
  assign n3653 = ~n3541 & n3652 ;
  assign n3654 = n3523 & n3653 ;
  assign n3655 = ~n3118 & n3135 ;
  assign n3656 = ~n3179 & ~n3655 ;
  assign n3657 = ~n3654 & n3656 ;
  assign n3658 = n3511 & n3513 ;
  assign n3659 = ~n3657 & ~n3658 ;
  assign n3660 = ~n3107 & n3659 ;
  assign n3661 = ~n3651 & ~n3660 ;
  assign n3662 = ~n3391 & n3412 ;
  assign n3663 = n3550 & n3558 ;
  assign n3664 = ~n3662 & ~n3663 ;
  assign n3665 = ~n3424 & n3664 ;
  assign n3666 = n3551 & n3552 ;
  assign n3667 = ~n3107 & ~n3666 ;
  assign n3668 = ~n3665 & n3667 ;
  assign n3669 = n3431 & n3436 ;
  assign n3670 = \ch_sel_dma_rrarb2_state_reg[2]/NET0131  & n3669 ;
  assign n3671 = \ch_sel_dma_rrarb2_state_reg[2]/NET0131  & n3106 ;
  assign n3672 = ~n3097 & n3671 ;
  assign n3673 = ~n3670 & ~n3672 ;
  assign n3674 = ~n3458 & ~n3585 ;
  assign n3675 = ~n3565 & ~n3585 ;
  assign n3676 = n3552 & n3675 ;
  assign n3677 = ~n3674 & ~n3676 ;
  assign n3678 = n3673 & ~n3677 ;
  assign n3679 = ~n3668 & n3678 ;
  assign n3680 = \ch_sel_dma_rrarb3_state_reg[1]/NET0131  & ~n3592 ;
  assign n3681 = ~\ch_sel_dma_rrarb3_state_reg[0]/NET0131  & \ctl_rf_c5_rf_chpri_reg[1]/NET0131  ;
  assign n3682 = \ctl_rf_c5_rf_chpri_reg[0]/NET0131  & n3681 ;
  assign n3683 = ~n3044 & n3682 ;
  assign n3684 = n3602 & ~n3683 ;
  assign n3685 = ~n3680 & ~n3684 ;
  assign n3686 = n3596 & n3598 ;
  assign n3687 = ~n3685 & ~n3686 ;
  assign n3688 = ~n3107 & n3687 ;
  assign n3689 = \ch_sel_dma_rrarb3_state_reg[2]/NET0131  & ~n3688 ;
  assign n3690 = n3595 & n3602 ;
  assign n3691 = n3596 & n3617 ;
  assign n3692 = ~n3225 & n3629 ;
  assign n3693 = ~n3254 & ~n3692 ;
  assign n3694 = ~n3691 & n3693 ;
  assign n3695 = ~n3690 & ~n3694 ;
  assign n3696 = ~n3107 & n3695 ;
  assign n3697 = ~n3689 & ~n3696 ;
  assign n3698 = n3304 & ~n3306 ;
  assign n3699 = ~n3345 & ~n3698 ;
  assign n3700 = ~n3309 & ~n3324 ;
  assign n3701 = ~n3311 & ~n3319 ;
  assign n3702 = ~n3314 & ~n3316 ;
  assign n3703 = n3701 & ~n3702 ;
  assign n3704 = n3700 & ~n3703 ;
  assign n3705 = ~n3699 & ~n3704 ;
  assign n3706 = ~n3306 & ~n3330 ;
  assign n3707 = ~n3700 & n3706 ;
  assign n3708 = n3702 & ~n3707 ;
  assign n3709 = ~\ch_sel_dma_rrarb0_state_reg[0]/NET0131  & ~\ctl_rf_c5_rf_chpri_reg[1]/NET0131  ;
  assign n3710 = ~\ctl_rf_c5_rf_chpri_reg[0]/NET0131  & n3709 ;
  assign n3711 = ~n3044 & n3710 ;
  assign n3712 = n3366 & ~n3711 ;
  assign n3713 = ~n3708 & n3712 ;
  assign n3714 = ~n3705 & ~n3713 ;
  assign n3715 = ~n3107 & ~n3714 ;
  assign n3716 = \ch_sel_dma_rrarb0_state_reg[1]/NET0131  & n3303 ;
  assign n3717 = n3308 & n3716 ;
  assign n3718 = ~n3033 & n3717 ;
  assign n3719 = ~\ch_sel_dma_rrarb0_state_reg[0]/NET0131  & ~\ctl_rf_c7_rf_chpri_reg[1]/NET0131  ;
  assign n3720 = ~\ctl_rf_c7_rf_chpri_reg[0]/NET0131  & n3719 ;
  assign n3721 = ~n3092 & n3720 ;
  assign n3722 = \ch_sel_dma_rrarb0_state_reg[1]/NET0131  & \ch_sel_dma_rrarb0_state_reg[2]/NET0131  ;
  assign n3723 = n3721 & n3722 ;
  assign n3724 = ~n3718 & ~n3723 ;
  assign n3725 = ~\ch_sel_dma_rrarb0_state_reg[1]/NET0131  & n3724 ;
  assign n3726 = ~\ch_sel_dma_rrarb0_state_reg[2]/NET0131  & n3703 ;
  assign n3727 = ~n3107 & ~n3726 ;
  assign n3728 = \ch_sel_dma_rrarb0_state_reg[2]/NET0131  & ~n3700 ;
  assign n3729 = ~n3701 & ~n3728 ;
  assign n3730 = n3706 & ~n3729 ;
  assign n3731 = n3724 & ~n3730 ;
  assign n3732 = n3727 & n3731 ;
  assign n3733 = ~n3725 & ~n3732 ;
  assign n3734 = ~n3715 & ~n3733 ;
  assign n3735 = n2935 & ~n2944 ;
  assign n3736 = \ch_sel_dma_rrarb0_state_reg[1]/NET0131  & ~n3721 ;
  assign n3737 = n3702 & ~n3711 ;
  assign n3738 = ~n3736 & ~n3737 ;
  assign n3739 = n3700 & n3706 ;
  assign n3740 = ~n3738 & ~n3739 ;
  assign n3741 = ~n3107 & n3740 ;
  assign n3742 = \ch_sel_dma_rrarb0_state_reg[2]/NET0131  & ~n3741 ;
  assign n3743 = n3324 & ~n3716 ;
  assign n3744 = ~n3345 & ~n3716 ;
  assign n3745 = ~n3698 & n3744 ;
  assign n3746 = ~n3743 & ~n3745 ;
  assign n3747 = ~n3309 & n3746 ;
  assign n3748 = ~n3352 & ~n3747 ;
  assign n3749 = n3701 & n3702 ;
  assign n3750 = ~n3107 & ~n3749 ;
  assign n3751 = ~n3748 & n3750 ;
  assign n3752 = ~n3742 & ~n3751 ;
  assign n3753 = \ahb_mst1_mx_cmd_st_reg[0]/NET0131  & ~\ahb_mst1_mx_cmd_st_reg[1]/NET0131  ;
  assign n3754 = ~n2930 & ~n3753 ;
  assign n3755 = ~\ahb_slv_slv_ad_d1o_reg[3]/NET0131  & ~\ahb_slv_slv_ad_d1o_reg[4]/NET0131  ;
  assign n3756 = n2275 & n3755 ;
  assign n3757 = n2317 & n3756 ;
  assign n3758 = ~\ctl_rf_be_d1_reg[2]/P0001  & n3757 ;
  assign n3759 = \hwdata[15]_pad  & ~n2242 ;
  assign n3760 = \hwdata[23]_pad  & n2242 ;
  assign n3761 = ~n3759 & ~n3760 ;
  assign n3762 = ~n2240 & ~n3761 ;
  assign n3763 = \hwdata[31]_pad  & n2240 ;
  assign n3764 = n3757 & ~n3763 ;
  assign n3765 = ~n3762 & n3764 ;
  assign n3766 = ~n3758 & ~n3765 ;
  assign n3767 = \hwdata[0]_pad  & ~n2242 ;
  assign n3768 = \hwdata[24]_pad  & n2242 ;
  assign n3769 = ~n3767 & ~n3768 ;
  assign n3770 = ~n2240 & ~n3769 ;
  assign n3771 = \hwdata[16]_pad  & n2240 ;
  assign n3772 = ~n3770 & ~n3771 ;
  assign n3773 = \ctl_rf_be_d1_reg[0]/P0001  & ~n3772 ;
  assign n3774 = ~n3766 & n3773 ;
  assign n3775 = \ctl_rf_c1_rf_chabt_reg/NET0131  & ~n2983 ;
  assign n3776 = n3050 & n3775 ;
  assign n3777 = \ctl_rf_c4_rf_chabt_reg/NET0131  & n2983 ;
  assign n3778 = n2999 & n3777 ;
  assign n3779 = ~n3776 & ~n3778 ;
  assign n3780 = \ctl_rf_c7_rf_chabt_reg/NET0131  & ~n2983 ;
  assign n3781 = n3011 & n3780 ;
  assign n3782 = \ctl_rf_c0_rf_chabt_reg/NET0131  & n2983 ;
  assign n3783 = n3050 & n3782 ;
  assign n3784 = ~n3781 & ~n3783 ;
  assign n3785 = n3779 & n3784 ;
  assign n3786 = \ctl_rf_c5_rf_chabt_reg/NET0131  & ~n2983 ;
  assign n3787 = n2999 & n3786 ;
  assign n3788 = \ctl_rf_c6_rf_chabt_reg/NET0131  & n2983 ;
  assign n3789 = n3011 & n3788 ;
  assign n3790 = ~n3787 & ~n3789 ;
  assign n3791 = \ctl_rf_c2_rf_chabt_reg/NET0131  & n2983 ;
  assign n3792 = n3024 & n3791 ;
  assign n3793 = \ctl_rf_c3_rf_chabt_reg/NET0131  & ~n2983 ;
  assign n3794 = n3024 & n3793 ;
  assign n3795 = ~n3792 & ~n3794 ;
  assign n3796 = n3790 & n3795 ;
  assign n3797 = n3785 & n3796 ;
  assign n3798 = n3000 & ~n3797 ;
  assign n3799 = n2983 & n3024 ;
  assign n3800 = ~\ctl_rf_c2_rf_chllp_reg[28]/NET0131  & ~\ctl_rf_c2_rf_chllp_reg[29]/NET0131  ;
  assign n3801 = ~\ctl_rf_c2_rf_chllp_reg[2]/NET0131  & ~\ctl_rf_c2_rf_chllp_reg[30]/NET0131  ;
  assign n3802 = n3800 & n3801 ;
  assign n3803 = ~\ctl_rf_c2_rf_chllp_reg[24]/NET0131  & ~\ctl_rf_c2_rf_chllp_reg[25]/NET0131  ;
  assign n3804 = ~\ctl_rf_c2_rf_chllp_reg[26]/NET0131  & ~\ctl_rf_c2_rf_chllp_reg[27]/NET0131  ;
  assign n3805 = n3803 & n3804 ;
  assign n3806 = n3802 & n3805 ;
  assign n3807 = ~\ctl_rf_c2_rf_chllp_reg[6]/NET0131  & ~\ctl_rf_c2_rf_chllp_reg[7]/NET0131  ;
  assign n3808 = ~\ctl_rf_c2_rf_chllp_reg[8]/NET0131  & ~\ctl_rf_c2_rf_chllp_reg[9]/NET0131  ;
  assign n3809 = n3807 & n3808 ;
  assign n3810 = ~\ctl_rf_c2_rf_chllp_reg[31]/NET0131  & ~\ctl_rf_c2_rf_chllp_reg[3]/NET0131  ;
  assign n3811 = ~\ctl_rf_c2_rf_chllp_reg[4]/NET0131  & ~\ctl_rf_c2_rf_chllp_reg[5]/NET0131  ;
  assign n3812 = n3810 & n3811 ;
  assign n3813 = n3809 & n3812 ;
  assign n3814 = n3806 & n3813 ;
  assign n3815 = ~\ctl_rf_c2_rf_chllp_reg[10]/NET0131  & ~\ctl_rf_c2_rf_chllp_reg[11]/NET0131  ;
  assign n3816 = ~\ctl_rf_c2_rf_chllp_reg[12]/NET0131  & ~\ctl_rf_c2_rf_chllp_reg[13]/NET0131  ;
  assign n3817 = ~\ctl_rf_c2_rf_chllp_reg[14]/NET0131  & ~\ctl_rf_c2_rf_chllp_reg[15]/NET0131  ;
  assign n3818 = n3816 & n3817 ;
  assign n3819 = n3815 & n3818 ;
  assign n3820 = ~\ctl_rf_c2_rf_chllp_reg[20]/NET0131  & ~\ctl_rf_c2_rf_chllp_reg[21]/NET0131  ;
  assign n3821 = ~\ctl_rf_c2_rf_chllp_reg[22]/NET0131  & ~\ctl_rf_c2_rf_chllp_reg[23]/NET0131  ;
  assign n3822 = n3820 & n3821 ;
  assign n3823 = ~\ctl_rf_c2_rf_chllp_reg[16]/NET0131  & ~\ctl_rf_c2_rf_chllp_reg[17]/NET0131  ;
  assign n3824 = ~\ctl_rf_c2_rf_chllp_reg[18]/NET0131  & ~\ctl_rf_c2_rf_chllp_reg[19]/NET0131  ;
  assign n3825 = n3823 & n3824 ;
  assign n3826 = n3822 & n3825 ;
  assign n3827 = n3819 & n3826 ;
  assign n3828 = n3814 & n3827 ;
  assign n3829 = n3799 & ~n3828 ;
  assign n3830 = n2983 & n2999 ;
  assign n3831 = ~\ctl_rf_c4_rf_chllp_reg[28]/NET0131  & ~\ctl_rf_c4_rf_chllp_reg[29]/NET0131  ;
  assign n3832 = ~\ctl_rf_c4_rf_chllp_reg[2]/NET0131  & ~\ctl_rf_c4_rf_chllp_reg[30]/NET0131  ;
  assign n3833 = n3831 & n3832 ;
  assign n3834 = ~\ctl_rf_c4_rf_chllp_reg[24]/NET0131  & ~\ctl_rf_c4_rf_chllp_reg[25]/NET0131  ;
  assign n3835 = ~\ctl_rf_c4_rf_chllp_reg[26]/NET0131  & ~\ctl_rf_c4_rf_chllp_reg[27]/NET0131  ;
  assign n3836 = n3834 & n3835 ;
  assign n3837 = n3833 & n3836 ;
  assign n3838 = ~\ctl_rf_c4_rf_chllp_reg[6]/NET0131  & ~\ctl_rf_c4_rf_chllp_reg[7]/NET0131  ;
  assign n3839 = ~\ctl_rf_c4_rf_chllp_reg[8]/NET0131  & ~\ctl_rf_c4_rf_chllp_reg[9]/NET0131  ;
  assign n3840 = n3838 & n3839 ;
  assign n3841 = ~\ctl_rf_c4_rf_chllp_reg[31]/NET0131  & ~\ctl_rf_c4_rf_chllp_reg[3]/NET0131  ;
  assign n3842 = ~\ctl_rf_c4_rf_chllp_reg[4]/NET0131  & ~\ctl_rf_c4_rf_chllp_reg[5]/NET0131  ;
  assign n3843 = n3841 & n3842 ;
  assign n3844 = n3840 & n3843 ;
  assign n3845 = n3837 & n3844 ;
  assign n3846 = ~\ctl_rf_c4_rf_chllp_reg[10]/NET0131  & ~\ctl_rf_c4_rf_chllp_reg[11]/NET0131  ;
  assign n3847 = ~\ctl_rf_c4_rf_chllp_reg[12]/NET0131  & ~\ctl_rf_c4_rf_chllp_reg[13]/NET0131  ;
  assign n3848 = ~\ctl_rf_c4_rf_chllp_reg[14]/NET0131  & ~\ctl_rf_c4_rf_chllp_reg[15]/NET0131  ;
  assign n3849 = n3847 & n3848 ;
  assign n3850 = n3846 & n3849 ;
  assign n3851 = ~\ctl_rf_c4_rf_chllp_reg[20]/NET0131  & ~\ctl_rf_c4_rf_chllp_reg[21]/NET0131  ;
  assign n3852 = ~\ctl_rf_c4_rf_chllp_reg[22]/NET0131  & ~\ctl_rf_c4_rf_chllp_reg[23]/NET0131  ;
  assign n3853 = n3851 & n3852 ;
  assign n3854 = ~\ctl_rf_c4_rf_chllp_reg[16]/NET0131  & ~\ctl_rf_c4_rf_chllp_reg[17]/NET0131  ;
  assign n3855 = ~\ctl_rf_c4_rf_chllp_reg[18]/NET0131  & ~\ctl_rf_c4_rf_chllp_reg[19]/NET0131  ;
  assign n3856 = n3854 & n3855 ;
  assign n3857 = n3853 & n3856 ;
  assign n3858 = n3850 & n3857 ;
  assign n3859 = n3845 & n3858 ;
  assign n3860 = n3830 & ~n3859 ;
  assign n3861 = ~n3829 & ~n3860 ;
  assign n3862 = ~n2983 & n3050 ;
  assign n3863 = ~\ctl_rf_c1_rf_chllp_reg[28]/NET0131  & ~\ctl_rf_c1_rf_chllp_reg[29]/NET0131  ;
  assign n3864 = ~\ctl_rf_c1_rf_chllp_reg[2]/NET0131  & ~\ctl_rf_c1_rf_chllp_reg[30]/NET0131  ;
  assign n3865 = n3863 & n3864 ;
  assign n3866 = ~\ctl_rf_c1_rf_chllp_reg[24]/NET0131  & ~\ctl_rf_c1_rf_chllp_reg[25]/NET0131  ;
  assign n3867 = ~\ctl_rf_c1_rf_chllp_reg[26]/NET0131  & ~\ctl_rf_c1_rf_chllp_reg[27]/NET0131  ;
  assign n3868 = n3866 & n3867 ;
  assign n3869 = n3865 & n3868 ;
  assign n3870 = ~\ctl_rf_c1_rf_chllp_reg[6]/NET0131  & ~\ctl_rf_c1_rf_chllp_reg[7]/NET0131  ;
  assign n3871 = ~\ctl_rf_c1_rf_chllp_reg[8]/NET0131  & ~\ctl_rf_c1_rf_chllp_reg[9]/NET0131  ;
  assign n3872 = n3870 & n3871 ;
  assign n3873 = ~\ctl_rf_c1_rf_chllp_reg[31]/NET0131  & ~\ctl_rf_c1_rf_chllp_reg[3]/NET0131  ;
  assign n3874 = ~\ctl_rf_c1_rf_chllp_reg[4]/NET0131  & ~\ctl_rf_c1_rf_chllp_reg[5]/NET0131  ;
  assign n3875 = n3873 & n3874 ;
  assign n3876 = n3872 & n3875 ;
  assign n3877 = n3869 & n3876 ;
  assign n3878 = ~\ctl_rf_c1_rf_chllp_reg[10]/NET0131  & ~\ctl_rf_c1_rf_chllp_reg[11]/NET0131  ;
  assign n3879 = ~\ctl_rf_c1_rf_chllp_reg[12]/NET0131  & ~\ctl_rf_c1_rf_chllp_reg[13]/NET0131  ;
  assign n3880 = ~\ctl_rf_c1_rf_chllp_reg[14]/NET0131  & ~\ctl_rf_c1_rf_chllp_reg[15]/NET0131  ;
  assign n3881 = n3879 & n3880 ;
  assign n3882 = n3878 & n3881 ;
  assign n3883 = ~\ctl_rf_c1_rf_chllp_reg[20]/NET0131  & ~\ctl_rf_c1_rf_chllp_reg[21]/NET0131  ;
  assign n3884 = ~\ctl_rf_c1_rf_chllp_reg[22]/NET0131  & ~\ctl_rf_c1_rf_chllp_reg[23]/NET0131  ;
  assign n3885 = n3883 & n3884 ;
  assign n3886 = ~\ctl_rf_c1_rf_chllp_reg[16]/NET0131  & ~\ctl_rf_c1_rf_chllp_reg[17]/NET0131  ;
  assign n3887 = ~\ctl_rf_c1_rf_chllp_reg[18]/NET0131  & ~\ctl_rf_c1_rf_chllp_reg[19]/NET0131  ;
  assign n3888 = n3886 & n3887 ;
  assign n3889 = n3885 & n3888 ;
  assign n3890 = n3882 & n3889 ;
  assign n3891 = n3877 & n3890 ;
  assign n3892 = n3862 & ~n3891 ;
  assign n3893 = ~n2983 & n3024 ;
  assign n3894 = ~\ctl_rf_c3_rf_chllp_reg[28]/NET0131  & ~\ctl_rf_c3_rf_chllp_reg[29]/NET0131  ;
  assign n3895 = ~\ctl_rf_c3_rf_chllp_reg[2]/NET0131  & ~\ctl_rf_c3_rf_chllp_reg[30]/NET0131  ;
  assign n3896 = n3894 & n3895 ;
  assign n3897 = ~\ctl_rf_c3_rf_chllp_reg[24]/NET0131  & ~\ctl_rf_c3_rf_chllp_reg[25]/NET0131  ;
  assign n3898 = ~\ctl_rf_c3_rf_chllp_reg[26]/NET0131  & ~\ctl_rf_c3_rf_chllp_reg[27]/NET0131  ;
  assign n3899 = n3897 & n3898 ;
  assign n3900 = n3896 & n3899 ;
  assign n3901 = ~\ctl_rf_c3_rf_chllp_reg[6]/NET0131  & ~\ctl_rf_c3_rf_chllp_reg[7]/NET0131  ;
  assign n3902 = ~\ctl_rf_c3_rf_chllp_reg[8]/NET0131  & ~\ctl_rf_c3_rf_chllp_reg[9]/NET0131  ;
  assign n3903 = n3901 & n3902 ;
  assign n3904 = ~\ctl_rf_c3_rf_chllp_reg[31]/NET0131  & ~\ctl_rf_c3_rf_chllp_reg[3]/NET0131  ;
  assign n3905 = ~\ctl_rf_c3_rf_chllp_reg[4]/NET0131  & ~\ctl_rf_c3_rf_chllp_reg[5]/NET0131  ;
  assign n3906 = n3904 & n3905 ;
  assign n3907 = n3903 & n3906 ;
  assign n3908 = n3900 & n3907 ;
  assign n3909 = ~\ctl_rf_c3_rf_chllp_reg[10]/NET0131  & ~\ctl_rf_c3_rf_chllp_reg[11]/NET0131  ;
  assign n3910 = ~\ctl_rf_c3_rf_chllp_reg[12]/NET0131  & ~\ctl_rf_c3_rf_chllp_reg[13]/NET0131  ;
  assign n3911 = ~\ctl_rf_c3_rf_chllp_reg[14]/NET0131  & ~\ctl_rf_c3_rf_chllp_reg[15]/NET0131  ;
  assign n3912 = n3910 & n3911 ;
  assign n3913 = n3909 & n3912 ;
  assign n3914 = ~\ctl_rf_c3_rf_chllp_reg[20]/NET0131  & ~\ctl_rf_c3_rf_chllp_reg[21]/NET0131  ;
  assign n3915 = ~\ctl_rf_c3_rf_chllp_reg[22]/NET0131  & ~\ctl_rf_c3_rf_chllp_reg[23]/NET0131  ;
  assign n3916 = n3914 & n3915 ;
  assign n3917 = ~\ctl_rf_c3_rf_chllp_reg[16]/NET0131  & ~\ctl_rf_c3_rf_chllp_reg[17]/NET0131  ;
  assign n3918 = ~\ctl_rf_c3_rf_chllp_reg[18]/NET0131  & ~\ctl_rf_c3_rf_chllp_reg[19]/NET0131  ;
  assign n3919 = n3917 & n3918 ;
  assign n3920 = n3916 & n3919 ;
  assign n3921 = n3913 & n3920 ;
  assign n3922 = n3908 & n3921 ;
  assign n3923 = n3893 & ~n3922 ;
  assign n3924 = ~n3892 & ~n3923 ;
  assign n3925 = n3861 & n3924 ;
  assign n3926 = ~n2983 & n3011 ;
  assign n3927 = ~\ctl_rf_c7_rf_chllp_reg[28]/NET0131  & ~\ctl_rf_c7_rf_chllp_reg[29]/NET0131  ;
  assign n3928 = ~\ctl_rf_c7_rf_chllp_reg[2]/NET0131  & ~\ctl_rf_c7_rf_chllp_reg[30]/NET0131  ;
  assign n3929 = n3927 & n3928 ;
  assign n3930 = ~\ctl_rf_c7_rf_chllp_reg[24]/NET0131  & ~\ctl_rf_c7_rf_chllp_reg[25]/NET0131  ;
  assign n3931 = ~\ctl_rf_c7_rf_chllp_reg[26]/NET0131  & ~\ctl_rf_c7_rf_chllp_reg[27]/NET0131  ;
  assign n3932 = n3930 & n3931 ;
  assign n3933 = n3929 & n3932 ;
  assign n3934 = ~\ctl_rf_c7_rf_chllp_reg[6]/NET0131  & ~\ctl_rf_c7_rf_chllp_reg[7]/NET0131  ;
  assign n3935 = ~\ctl_rf_c7_rf_chllp_reg[8]/NET0131  & ~\ctl_rf_c7_rf_chllp_reg[9]/NET0131  ;
  assign n3936 = n3934 & n3935 ;
  assign n3937 = ~\ctl_rf_c7_rf_chllp_reg[31]/NET0131  & ~\ctl_rf_c7_rf_chllp_reg[3]/NET0131  ;
  assign n3938 = ~\ctl_rf_c7_rf_chllp_reg[4]/NET0131  & ~\ctl_rf_c7_rf_chllp_reg[5]/NET0131  ;
  assign n3939 = n3937 & n3938 ;
  assign n3940 = n3936 & n3939 ;
  assign n3941 = n3933 & n3940 ;
  assign n3942 = ~\ctl_rf_c7_rf_chllp_reg[10]/NET0131  & ~\ctl_rf_c7_rf_chllp_reg[11]/NET0131  ;
  assign n3943 = ~\ctl_rf_c7_rf_chllp_reg[12]/NET0131  & ~\ctl_rf_c7_rf_chllp_reg[13]/NET0131  ;
  assign n3944 = ~\ctl_rf_c7_rf_chllp_reg[14]/NET0131  & ~\ctl_rf_c7_rf_chllp_reg[15]/NET0131  ;
  assign n3945 = n3943 & n3944 ;
  assign n3946 = n3942 & n3945 ;
  assign n3947 = ~\ctl_rf_c7_rf_chllp_reg[20]/NET0131  & ~\ctl_rf_c7_rf_chllp_reg[21]/NET0131  ;
  assign n3948 = ~\ctl_rf_c7_rf_chllp_reg[22]/NET0131  & ~\ctl_rf_c7_rf_chllp_reg[23]/NET0131  ;
  assign n3949 = n3947 & n3948 ;
  assign n3950 = ~\ctl_rf_c7_rf_chllp_reg[16]/NET0131  & ~\ctl_rf_c7_rf_chllp_reg[17]/NET0131  ;
  assign n3951 = ~\ctl_rf_c7_rf_chllp_reg[18]/NET0131  & ~\ctl_rf_c7_rf_chllp_reg[19]/NET0131  ;
  assign n3952 = n3950 & n3951 ;
  assign n3953 = n3949 & n3952 ;
  assign n3954 = n3946 & n3953 ;
  assign n3955 = n3941 & n3954 ;
  assign n3956 = n3926 & ~n3955 ;
  assign n3957 = ~n2983 & n2999 ;
  assign n3958 = ~\ctl_rf_c5_rf_chllp_reg[28]/NET0131  & ~\ctl_rf_c5_rf_chllp_reg[29]/NET0131  ;
  assign n3959 = ~\ctl_rf_c5_rf_chllp_reg[2]/NET0131  & ~\ctl_rf_c5_rf_chllp_reg[30]/NET0131  ;
  assign n3960 = n3958 & n3959 ;
  assign n3961 = ~\ctl_rf_c5_rf_chllp_reg[24]/NET0131  & ~\ctl_rf_c5_rf_chllp_reg[25]/NET0131  ;
  assign n3962 = ~\ctl_rf_c5_rf_chllp_reg[26]/NET0131  & ~\ctl_rf_c5_rf_chllp_reg[27]/NET0131  ;
  assign n3963 = n3961 & n3962 ;
  assign n3964 = n3960 & n3963 ;
  assign n3965 = ~\ctl_rf_c5_rf_chllp_reg[6]/NET0131  & ~\ctl_rf_c5_rf_chllp_reg[7]/NET0131  ;
  assign n3966 = ~\ctl_rf_c5_rf_chllp_reg[8]/NET0131  & ~\ctl_rf_c5_rf_chllp_reg[9]/NET0131  ;
  assign n3967 = n3965 & n3966 ;
  assign n3968 = ~\ctl_rf_c5_rf_chllp_reg[31]/NET0131  & ~\ctl_rf_c5_rf_chllp_reg[3]/NET0131  ;
  assign n3969 = ~\ctl_rf_c5_rf_chllp_reg[4]/NET0131  & ~\ctl_rf_c5_rf_chllp_reg[5]/NET0131  ;
  assign n3970 = n3968 & n3969 ;
  assign n3971 = n3967 & n3970 ;
  assign n3972 = n3964 & n3971 ;
  assign n3973 = ~\ctl_rf_c5_rf_chllp_reg[10]/NET0131  & ~\ctl_rf_c5_rf_chllp_reg[11]/NET0131  ;
  assign n3974 = ~\ctl_rf_c5_rf_chllp_reg[12]/NET0131  & ~\ctl_rf_c5_rf_chllp_reg[13]/NET0131  ;
  assign n3975 = ~\ctl_rf_c5_rf_chllp_reg[14]/NET0131  & ~\ctl_rf_c5_rf_chllp_reg[15]/NET0131  ;
  assign n3976 = n3974 & n3975 ;
  assign n3977 = n3973 & n3976 ;
  assign n3978 = ~\ctl_rf_c5_rf_chllp_reg[20]/NET0131  & ~\ctl_rf_c5_rf_chllp_reg[21]/NET0131  ;
  assign n3979 = ~\ctl_rf_c5_rf_chllp_reg[22]/NET0131  & ~\ctl_rf_c5_rf_chllp_reg[23]/NET0131  ;
  assign n3980 = n3978 & n3979 ;
  assign n3981 = ~\ctl_rf_c5_rf_chllp_reg[16]/NET0131  & ~\ctl_rf_c5_rf_chllp_reg[17]/NET0131  ;
  assign n3982 = ~\ctl_rf_c5_rf_chllp_reg[18]/NET0131  & ~\ctl_rf_c5_rf_chllp_reg[19]/NET0131  ;
  assign n3983 = n3981 & n3982 ;
  assign n3984 = n3980 & n3983 ;
  assign n3985 = n3977 & n3984 ;
  assign n3986 = n3972 & n3985 ;
  assign n3987 = n3957 & ~n3986 ;
  assign n3988 = ~n3956 & ~n3987 ;
  assign n3989 = n2983 & n3050 ;
  assign n3990 = ~\ctl_rf_c0_rf_chllp_reg[28]/NET0131  & ~\ctl_rf_c0_rf_chllp_reg[29]/NET0131  ;
  assign n3991 = ~\ctl_rf_c0_rf_chllp_reg[2]/NET0131  & ~\ctl_rf_c0_rf_chllp_reg[30]/NET0131  ;
  assign n3992 = n3990 & n3991 ;
  assign n3993 = ~\ctl_rf_c0_rf_chllp_reg[24]/NET0131  & ~\ctl_rf_c0_rf_chllp_reg[25]/NET0131  ;
  assign n3994 = ~\ctl_rf_c0_rf_chllp_reg[26]/NET0131  & ~\ctl_rf_c0_rf_chllp_reg[27]/NET0131  ;
  assign n3995 = n3993 & n3994 ;
  assign n3996 = n3992 & n3995 ;
  assign n3997 = ~\ctl_rf_c0_rf_chllp_reg[6]/NET0131  & ~\ctl_rf_c0_rf_chllp_reg[7]/NET0131  ;
  assign n3998 = ~\ctl_rf_c0_rf_chllp_reg[8]/NET0131  & ~\ctl_rf_c0_rf_chllp_reg[9]/NET0131  ;
  assign n3999 = n3997 & n3998 ;
  assign n4000 = ~\ctl_rf_c0_rf_chllp_reg[31]/NET0131  & ~\ctl_rf_c0_rf_chllp_reg[3]/NET0131  ;
  assign n4001 = ~\ctl_rf_c0_rf_chllp_reg[4]/NET0131  & ~\ctl_rf_c0_rf_chllp_reg[5]/NET0131  ;
  assign n4002 = n4000 & n4001 ;
  assign n4003 = n3999 & n4002 ;
  assign n4004 = n3996 & n4003 ;
  assign n4005 = ~\ctl_rf_c0_rf_chllp_reg[10]/NET0131  & ~\ctl_rf_c0_rf_chllp_reg[11]/NET0131  ;
  assign n4006 = ~\ctl_rf_c0_rf_chllp_reg[12]/NET0131  & ~\ctl_rf_c0_rf_chllp_reg[13]/NET0131  ;
  assign n4007 = ~\ctl_rf_c0_rf_chllp_reg[14]/NET0131  & ~\ctl_rf_c0_rf_chllp_reg[15]/NET0131  ;
  assign n4008 = n4006 & n4007 ;
  assign n4009 = n4005 & n4008 ;
  assign n4010 = ~\ctl_rf_c0_rf_chllp_reg[20]/NET0131  & ~\ctl_rf_c0_rf_chllp_reg[21]/NET0131  ;
  assign n4011 = ~\ctl_rf_c0_rf_chllp_reg[22]/NET0131  & ~\ctl_rf_c0_rf_chllp_reg[23]/NET0131  ;
  assign n4012 = n4010 & n4011 ;
  assign n4013 = ~\ctl_rf_c0_rf_chllp_reg[16]/NET0131  & ~\ctl_rf_c0_rf_chllp_reg[17]/NET0131  ;
  assign n4014 = ~\ctl_rf_c0_rf_chllp_reg[18]/NET0131  & ~\ctl_rf_c0_rf_chllp_reg[19]/NET0131  ;
  assign n4015 = n4013 & n4014 ;
  assign n4016 = n4012 & n4015 ;
  assign n4017 = n4009 & n4016 ;
  assign n4018 = n4004 & n4017 ;
  assign n4019 = n3989 & ~n4018 ;
  assign n4020 = n2983 & n3011 ;
  assign n4021 = ~\ctl_rf_c6_rf_chllp_reg[28]/NET0131  & ~\ctl_rf_c6_rf_chllp_reg[29]/NET0131  ;
  assign n4022 = ~\ctl_rf_c6_rf_chllp_reg[2]/NET0131  & ~\ctl_rf_c6_rf_chllp_reg[30]/NET0131  ;
  assign n4023 = n4021 & n4022 ;
  assign n4024 = ~\ctl_rf_c6_rf_chllp_reg[24]/NET0131  & ~\ctl_rf_c6_rf_chllp_reg[25]/NET0131  ;
  assign n4025 = ~\ctl_rf_c6_rf_chllp_reg[26]/NET0131  & ~\ctl_rf_c6_rf_chllp_reg[27]/NET0131  ;
  assign n4026 = n4024 & n4025 ;
  assign n4027 = n4023 & n4026 ;
  assign n4028 = ~\ctl_rf_c6_rf_chllp_reg[6]/NET0131  & ~\ctl_rf_c6_rf_chllp_reg[7]/NET0131  ;
  assign n4029 = ~\ctl_rf_c6_rf_chllp_reg[8]/NET0131  & ~\ctl_rf_c6_rf_chllp_reg[9]/NET0131  ;
  assign n4030 = n4028 & n4029 ;
  assign n4031 = ~\ctl_rf_c6_rf_chllp_reg[31]/NET0131  & ~\ctl_rf_c6_rf_chllp_reg[3]/NET0131  ;
  assign n4032 = ~\ctl_rf_c6_rf_chllp_reg[4]/NET0131  & ~\ctl_rf_c6_rf_chllp_reg[5]/NET0131  ;
  assign n4033 = n4031 & n4032 ;
  assign n4034 = n4030 & n4033 ;
  assign n4035 = n4027 & n4034 ;
  assign n4036 = ~\ctl_rf_c6_rf_chllp_reg[10]/NET0131  & ~\ctl_rf_c6_rf_chllp_reg[11]/NET0131  ;
  assign n4037 = ~\ctl_rf_c6_rf_chllp_reg[12]/NET0131  & ~\ctl_rf_c6_rf_chllp_reg[13]/NET0131  ;
  assign n4038 = ~\ctl_rf_c6_rf_chllp_reg[14]/NET0131  & ~\ctl_rf_c6_rf_chllp_reg[15]/NET0131  ;
  assign n4039 = n4037 & n4038 ;
  assign n4040 = n4036 & n4039 ;
  assign n4041 = ~\ctl_rf_c6_rf_chllp_reg[20]/NET0131  & ~\ctl_rf_c6_rf_chllp_reg[21]/NET0131  ;
  assign n4042 = ~\ctl_rf_c6_rf_chllp_reg[22]/NET0131  & ~\ctl_rf_c6_rf_chllp_reg[23]/NET0131  ;
  assign n4043 = n4041 & n4042 ;
  assign n4044 = ~\ctl_rf_c6_rf_chllp_reg[16]/NET0131  & ~\ctl_rf_c6_rf_chllp_reg[17]/NET0131  ;
  assign n4045 = ~\ctl_rf_c6_rf_chllp_reg[18]/NET0131  & ~\ctl_rf_c6_rf_chllp_reg[19]/NET0131  ;
  assign n4046 = n4044 & n4045 ;
  assign n4047 = n4043 & n4046 ;
  assign n4048 = n4040 & n4047 ;
  assign n4049 = n4035 & n4048 ;
  assign n4050 = n4020 & ~n4049 ;
  assign n4051 = ~n4019 & ~n4050 ;
  assign n4052 = n3988 & n4051 ;
  assign n4053 = n3925 & n4052 ;
  assign n4054 = n2814 & n3000 ;
  assign n4055 = n4053 & n4054 ;
  assign n4056 = ~n3798 & ~n4055 ;
  assign n4057 = \ctl_rf_be_d1_reg[0]/P0001  & ~n3766 ;
  assign n4058 = ~\de_de_st_reg[0]/NET0131  & n2983 ;
  assign n4059 = n2999 & n4058 ;
  assign n4060 = \ctl_rf_c4_rf_chabt_reg/NET0131  & ~n4059 ;
  assign n4061 = \ctl_rf_c4_rf_ch_en_reg/NET0131  & ~n4060 ;
  assign n4062 = ~n4057 & n4061 ;
  assign n4063 = n4056 & n4062 ;
  assign n4064 = ~n3774 & ~n4063 ;
  assign n4065 = n2232 & n3755 ;
  assign n4066 = n2317 & n4065 ;
  assign n4067 = ~\ctl_rf_be_d1_reg[2]/P0001  & n4066 ;
  assign n4068 = ~n3763 & n4066 ;
  assign n4069 = ~n3762 & n4068 ;
  assign n4070 = ~n4067 & ~n4069 ;
  assign n4071 = n3773 & ~n4070 ;
  assign n4072 = n3037 & ~n3797 ;
  assign n4073 = n2814 & n3037 ;
  assign n4074 = n4053 & n4073 ;
  assign n4075 = ~n4072 & ~n4074 ;
  assign n4076 = \ctl_rf_be_d1_reg[0]/P0001  & ~n4070 ;
  assign n4077 = ~\de_de_st_reg[0]/NET0131  & ~n2983 ;
  assign n4078 = n2999 & n4077 ;
  assign n4079 = \ctl_rf_c5_rf_chabt_reg/NET0131  & ~n4078 ;
  assign n4080 = \ctl_rf_c5_rf_ch_en_reg/NET0131  & ~n4079 ;
  assign n4081 = ~n4076 & n4080 ;
  assign n4082 = n4075 & n4081 ;
  assign n4083 = ~n4071 & ~n4082 ;
  assign n4084 = n2324 & n3756 ;
  assign n4085 = ~\ctl_rf_be_d1_reg[2]/P0001  & n4084 ;
  assign n4086 = ~n3763 & n4084 ;
  assign n4087 = ~n3762 & n4086 ;
  assign n4088 = ~n4085 & ~n4087 ;
  assign n4089 = n3773 & ~n4088 ;
  assign n4090 = n3012 & ~n3797 ;
  assign n4091 = n2814 & n3012 ;
  assign n4092 = n4053 & n4091 ;
  assign n4093 = ~n4090 & ~n4092 ;
  assign n4094 = \ctl_rf_be_d1_reg[0]/P0001  & ~n4088 ;
  assign n4095 = n3011 & n4058 ;
  assign n4096 = \ctl_rf_c6_rf_chabt_reg/NET0131  & ~n4095 ;
  assign n4097 = \ctl_rf_c6_rf_ch_en_reg/NET0131  & ~n4096 ;
  assign n4098 = ~n4094 & n4097 ;
  assign n4099 = n4093 & n4098 ;
  assign n4100 = ~n4089 & ~n4099 ;
  assign n4101 = n2324 & n4065 ;
  assign n4102 = ~\ctl_rf_be_d1_reg[2]/P0001  & n4101 ;
  assign n4103 = ~n3763 & n4101 ;
  assign n4104 = ~n3762 & n4103 ;
  assign n4105 = ~n4102 & ~n4104 ;
  assign n4106 = n3773 & ~n4105 ;
  assign n4107 = n3085 & ~n3797 ;
  assign n4108 = n2814 & n3085 ;
  assign n4109 = n4053 & n4108 ;
  assign n4110 = ~n4107 & ~n4109 ;
  assign n4111 = \ctl_rf_be_d1_reg[0]/P0001  & ~n4105 ;
  assign n4112 = n3011 & n4077 ;
  assign n4113 = \ctl_rf_c7_rf_chabt_reg/NET0131  & ~n4112 ;
  assign n4114 = \ctl_rf_c7_rf_ch_en_reg/NET0131  & ~n4113 ;
  assign n4115 = ~n4111 & n4114 ;
  assign n4116 = n4110 & n4115 ;
  assign n4117 = ~n4106 & ~n4116 ;
  assign n4118 = n2231 & n4065 ;
  assign n4119 = ~\ctl_rf_be_d1_reg[2]/P0001  & n4118 ;
  assign n4120 = ~n3763 & n4118 ;
  assign n4121 = ~n3762 & n4120 ;
  assign n4122 = ~n4119 & ~n4121 ;
  assign n4123 = n3773 & ~n4122 ;
  assign n4124 = n3074 & ~n3797 ;
  assign n4125 = n2814 & n3074 ;
  assign n4126 = n4053 & n4125 ;
  assign n4127 = ~n4124 & ~n4126 ;
  assign n4128 = \ctl_rf_be_d1_reg[0]/P0001  & ~n4122 ;
  assign n4129 = n3050 & n4077 ;
  assign n4130 = \ctl_rf_c1_rf_chabt_reg/NET0131  & ~n4129 ;
  assign n4131 = \ctl_rf_c1_rf_ch_en_reg/NET0131  & ~n4130 ;
  assign n4132 = ~n4128 & n4131 ;
  assign n4133 = n4127 & n4132 ;
  assign n4134 = ~n4123 & ~n4133 ;
  assign n4135 = n2311 & n3756 ;
  assign n4136 = ~\ctl_rf_be_d1_reg[2]/P0001  & n4135 ;
  assign n4137 = ~n3763 & n4135 ;
  assign n4138 = ~n3762 & n4137 ;
  assign n4139 = ~n4136 & ~n4138 ;
  assign n4140 = n3773 & ~n4139 ;
  assign n4141 = n3062 & ~n3797 ;
  assign n4142 = n2814 & n3062 ;
  assign n4143 = n4053 & n4142 ;
  assign n4144 = ~n4141 & ~n4143 ;
  assign n4145 = \ctl_rf_be_d1_reg[0]/P0001  & ~n4139 ;
  assign n4146 = n3024 & n4058 ;
  assign n4147 = \ctl_rf_c2_rf_chabt_reg/NET0131  & ~n4146 ;
  assign n4148 = \ctl_rf_c2_rf_ch_en_reg/NET0131  & ~n4147 ;
  assign n4149 = ~n4145 & n4148 ;
  assign n4150 = n4144 & n4149 ;
  assign n4151 = ~n4140 & ~n4150 ;
  assign n4152 = n2311 & n4065 ;
  assign n4153 = ~\ctl_rf_be_d1_reg[2]/P0001  & n4152 ;
  assign n4154 = ~n3763 & n4152 ;
  assign n4155 = ~n3762 & n4154 ;
  assign n4156 = ~n4153 & ~n4155 ;
  assign n4157 = n3773 & ~n4156 ;
  assign n4158 = n3026 & ~n3797 ;
  assign n4159 = n2814 & n3026 ;
  assign n4160 = n4053 & n4159 ;
  assign n4161 = ~n4158 & ~n4160 ;
  assign n4162 = \ctl_rf_be_d1_reg[0]/P0001  & ~n4156 ;
  assign n4163 = n3024 & n4077 ;
  assign n4164 = \ctl_rf_c3_rf_chabt_reg/NET0131  & ~n4163 ;
  assign n4165 = \ctl_rf_c3_rf_ch_en_reg/NET0131  & ~n4164 ;
  assign n4166 = ~n4162 & n4165 ;
  assign n4167 = n4161 & n4166 ;
  assign n4168 = ~n4157 & ~n4167 ;
  assign n4169 = n2231 & n3756 ;
  assign n4170 = ~\ctl_rf_be_d1_reg[2]/P0001  & n4169 ;
  assign n4171 = ~n3763 & n4169 ;
  assign n4172 = ~n3762 & n4171 ;
  assign n4173 = ~n4170 & ~n4172 ;
  assign n4174 = n3773 & ~n4173 ;
  assign n4175 = n3051 & ~n3797 ;
  assign n4176 = n2814 & n3051 ;
  assign n4177 = n4053 & n4176 ;
  assign n4178 = ~n4175 & ~n4177 ;
  assign n4179 = \ctl_rf_be_d1_reg[0]/P0001  & ~n4173 ;
  assign n4180 = n3050 & n4058 ;
  assign n4181 = \ctl_rf_c0_rf_chabt_reg/NET0131  & ~n4180 ;
  assign n4182 = \ctl_rf_c0_rf_ch_en_reg/NET0131  & ~n4181 ;
  assign n4183 = ~n4179 & n4182 ;
  assign n4184 = n4178 & n4183 ;
  assign n4185 = ~n4174 & ~n4184 ;
  assign n4186 = \ctl_rf_c1_rf_chtsz_reg[2]/P0002  & ~n2983 ;
  assign n4187 = n3050 & n4186 ;
  assign n4188 = \ctl_rf_c2_rf_chtsz_reg[2]/P0002  & n2983 ;
  assign n4189 = n3024 & n4188 ;
  assign n4190 = ~n4187 & ~n4189 ;
  assign n4191 = \ctl_rf_c7_rf_chtsz_reg[2]/P0002  & ~n2983 ;
  assign n4192 = n3011 & n4191 ;
  assign n4193 = \ctl_rf_c0_rf_chtsz_reg[2]/P0002  & n2983 ;
  assign n4194 = n3050 & n4193 ;
  assign n4195 = ~n4192 & ~n4194 ;
  assign n4196 = n4190 & n4195 ;
  assign n4197 = \ctl_rf_c3_rf_chtsz_reg[2]/P0002  & ~n2983 ;
  assign n4198 = n3024 & n4197 ;
  assign n4199 = \ctl_rf_c6_rf_chtsz_reg[2]/P0002  & n2983 ;
  assign n4200 = n3011 & n4199 ;
  assign n4201 = ~n4198 & ~n4200 ;
  assign n4202 = \ctl_rf_c4_rf_chtsz_reg[2]/P0002  & n2983 ;
  assign n4203 = n2999 & n4202 ;
  assign n4204 = \ctl_rf_c5_rf_chtsz_reg[2]/P0002  & ~n2983 ;
  assign n4205 = n2999 & n4204 ;
  assign n4206 = ~n4203 & ~n4205 ;
  assign n4207 = n4201 & n4206 ;
  assign n4208 = n4196 & n4207 ;
  assign n4209 = \ctl_rf_c1_rf_chtsz_reg[4]/NET0131  & ~n2983 ;
  assign n4210 = n3050 & n4209 ;
  assign n4211 = \ctl_rf_c2_rf_chtsz_reg[4]/NET0131  & n2983 ;
  assign n4212 = n3024 & n4211 ;
  assign n4213 = ~n4210 & ~n4212 ;
  assign n4214 = \ctl_rf_c7_rf_chtsz_reg[4]/NET0131  & ~n2983 ;
  assign n4215 = n3011 & n4214 ;
  assign n4216 = \ctl_rf_c0_rf_chtsz_reg[4]/NET0131  & n2983 ;
  assign n4217 = n3050 & n4216 ;
  assign n4218 = ~n4215 & ~n4217 ;
  assign n4219 = n4213 & n4218 ;
  assign n4220 = \ctl_rf_c3_rf_chtsz_reg[4]/NET0131  & ~n2983 ;
  assign n4221 = n3024 & n4220 ;
  assign n4222 = \ctl_rf_c6_rf_chtsz_reg[4]/NET0131  & n2983 ;
  assign n4223 = n3011 & n4222 ;
  assign n4224 = ~n4221 & ~n4223 ;
  assign n4225 = \ctl_rf_c4_rf_chtsz_reg[4]/NET0131  & n2983 ;
  assign n4226 = n2999 & n4225 ;
  assign n4227 = \ctl_rf_c5_rf_chtsz_reg[4]/NET0131  & ~n2983 ;
  assign n4228 = n2999 & n4227 ;
  assign n4229 = ~n4226 & ~n4228 ;
  assign n4230 = n4224 & n4229 ;
  assign n4231 = n4219 & n4230 ;
  assign n4232 = n4208 & n4231 ;
  assign n4233 = \ctl_rf_c1_rf_chtsz_reg[1]/P0002  & ~n2983 ;
  assign n4234 = n3050 & n4233 ;
  assign n4235 = \ctl_rf_c2_rf_chtsz_reg[1]/P0002  & n2983 ;
  assign n4236 = n3024 & n4235 ;
  assign n4237 = ~n4234 & ~n4236 ;
  assign n4238 = \ctl_rf_c7_rf_chtsz_reg[1]/P0002  & ~n2983 ;
  assign n4239 = n3011 & n4238 ;
  assign n4240 = \ctl_rf_c0_rf_chtsz_reg[1]/P0002  & n2983 ;
  assign n4241 = n3050 & n4240 ;
  assign n4242 = ~n4239 & ~n4241 ;
  assign n4243 = n4237 & n4242 ;
  assign n4244 = \ctl_rf_c3_rf_chtsz_reg[1]/P0002  & ~n2983 ;
  assign n4245 = n3024 & n4244 ;
  assign n4246 = \ctl_rf_c6_rf_chtsz_reg[1]/P0002  & n2983 ;
  assign n4247 = n3011 & n4246 ;
  assign n4248 = ~n4245 & ~n4247 ;
  assign n4249 = \ctl_rf_c4_rf_chtsz_reg[1]/P0002  & n2983 ;
  assign n4250 = n2999 & n4249 ;
  assign n4251 = \ctl_rf_c5_rf_chtsz_reg[1]/P0002  & ~n2983 ;
  assign n4252 = n2999 & n4251 ;
  assign n4253 = ~n4250 & ~n4252 ;
  assign n4254 = n4248 & n4253 ;
  assign n4255 = n4243 & n4254 ;
  assign n4256 = \ctl_rf_c1_rf_chtsz_reg[11]/P0002  & ~n2983 ;
  assign n4257 = n3050 & n4256 ;
  assign n4258 = \ctl_rf_c2_rf_chtsz_reg[11]/P0002  & n2983 ;
  assign n4259 = n3024 & n4258 ;
  assign n4260 = ~n4257 & ~n4259 ;
  assign n4261 = \ctl_rf_c7_rf_chtsz_reg[11]/P0002  & ~n2983 ;
  assign n4262 = n3011 & n4261 ;
  assign n4263 = \ctl_rf_c0_rf_chtsz_reg[11]/P0002  & n2983 ;
  assign n4264 = n3050 & n4263 ;
  assign n4265 = ~n4262 & ~n4264 ;
  assign n4266 = n4260 & n4265 ;
  assign n4267 = \ctl_rf_c3_rf_chtsz_reg[11]/P0002  & ~n2983 ;
  assign n4268 = n3024 & n4267 ;
  assign n4269 = \ctl_rf_c6_rf_chtsz_reg[11]/P0002  & n2983 ;
  assign n4270 = n3011 & n4269 ;
  assign n4271 = ~n4268 & ~n4270 ;
  assign n4272 = \ctl_rf_c4_rf_chtsz_reg[11]/P0002  & n2983 ;
  assign n4273 = n2999 & n4272 ;
  assign n4274 = \ctl_rf_c5_rf_chtsz_reg[11]/P0002  & ~n2983 ;
  assign n4275 = n2999 & n4274 ;
  assign n4276 = ~n4273 & ~n4275 ;
  assign n4277 = n4271 & n4276 ;
  assign n4278 = n4266 & n4277 ;
  assign n4279 = n4255 & n4278 ;
  assign n4280 = n4232 & n4279 ;
  assign n4281 = \ctl_rf_c1_rf_chtsz_reg[5]/NET0131  & ~n2983 ;
  assign n4282 = n3050 & n4281 ;
  assign n4283 = \ctl_rf_c2_rf_chtsz_reg[5]/NET0131  & n2983 ;
  assign n4284 = n3024 & n4283 ;
  assign n4285 = ~n4282 & ~n4284 ;
  assign n4286 = \ctl_rf_c7_rf_chtsz_reg[5]/NET0131  & ~n2983 ;
  assign n4287 = n3011 & n4286 ;
  assign n4288 = \ctl_rf_c0_rf_chtsz_reg[5]/NET0131  & n2983 ;
  assign n4289 = n3050 & n4288 ;
  assign n4290 = ~n4287 & ~n4289 ;
  assign n4291 = n4285 & n4290 ;
  assign n4292 = \ctl_rf_c3_rf_chtsz_reg[5]/NET0131  & ~n2983 ;
  assign n4293 = n3024 & n4292 ;
  assign n4294 = \ctl_rf_c6_rf_chtsz_reg[5]/NET0131  & n2983 ;
  assign n4295 = n3011 & n4294 ;
  assign n4296 = ~n4293 & ~n4295 ;
  assign n4297 = \ctl_rf_c4_rf_chtsz_reg[5]/NET0131  & n2983 ;
  assign n4298 = n2999 & n4297 ;
  assign n4299 = \ctl_rf_c5_rf_chtsz_reg[5]/NET0131  & ~n2983 ;
  assign n4300 = n2999 & n4299 ;
  assign n4301 = ~n4298 & ~n4300 ;
  assign n4302 = n4296 & n4301 ;
  assign n4303 = n4291 & n4302 ;
  assign n4304 = \ctl_rf_c7_rf_chllpen_reg/NET0131  & ~n2983 ;
  assign n4305 = n3011 & n4304 ;
  assign n4306 = \ctl_rf_c3_rf_chllpen_reg/NET0131  & ~n2983 ;
  assign n4307 = n3024 & n4306 ;
  assign n4308 = ~n4305 & ~n4307 ;
  assign n4309 = \ctl_rf_c1_rf_chllpen_reg/NET0131  & ~n2983 ;
  assign n4310 = n3050 & n4309 ;
  assign n4311 = \ctl_rf_c0_rf_chllpen_reg/NET0131  & n2983 ;
  assign n4312 = n3050 & n4311 ;
  assign n4313 = ~n4310 & ~n4312 ;
  assign n4314 = n4308 & n4313 ;
  assign n4315 = \ctl_rf_c2_rf_chllpen_reg/NET0131  & n2983 ;
  assign n4316 = n3024 & n4315 ;
  assign n4317 = \ctl_rf_c6_rf_chllpen_reg/NET0131  & n2983 ;
  assign n4318 = n3011 & n4317 ;
  assign n4319 = ~n4316 & ~n4318 ;
  assign n4320 = \ctl_rf_c4_rf_chllpen_reg/NET0131  & n2983 ;
  assign n4321 = n2999 & n4320 ;
  assign n4322 = \ctl_rf_c5_rf_chllpen_reg/NET0131  & ~n2983 ;
  assign n4323 = n2999 & n4322 ;
  assign n4324 = ~n4321 & ~n4323 ;
  assign n4325 = n4319 & n4324 ;
  assign n4326 = n4314 & n4325 ;
  assign n4327 = n4303 & n4326 ;
  assign n4328 = \ctl_rf_c1_rf_chtsz_reg[3]/P0002  & ~n2983 ;
  assign n4329 = n3050 & n4328 ;
  assign n4330 = \ctl_rf_c2_rf_chtsz_reg[3]/P0002  & n2983 ;
  assign n4331 = n3024 & n4330 ;
  assign n4332 = ~n4329 & ~n4331 ;
  assign n4333 = \ctl_rf_c7_rf_chtsz_reg[3]/P0002  & ~n2983 ;
  assign n4334 = n3011 & n4333 ;
  assign n4335 = \ctl_rf_c0_rf_chtsz_reg[3]/P0002  & n2983 ;
  assign n4336 = n3050 & n4335 ;
  assign n4337 = ~n4334 & ~n4336 ;
  assign n4338 = n4332 & n4337 ;
  assign n4339 = \ctl_rf_c3_rf_chtsz_reg[3]/P0002  & ~n2983 ;
  assign n4340 = n3024 & n4339 ;
  assign n4341 = \ctl_rf_c6_rf_chtsz_reg[3]/P0002  & n2983 ;
  assign n4342 = n3011 & n4341 ;
  assign n4343 = ~n4340 & ~n4342 ;
  assign n4344 = \ctl_rf_c4_rf_chtsz_reg[3]/P0002  & n2983 ;
  assign n4345 = n2999 & n4344 ;
  assign n4346 = \ctl_rf_c5_rf_chtsz_reg[3]/P0002  & ~n2983 ;
  assign n4347 = n2999 & n4346 ;
  assign n4348 = ~n4345 & ~n4347 ;
  assign n4349 = n4343 & n4348 ;
  assign n4350 = n4338 & n4349 ;
  assign n4351 = \ctl_rf_c1_rf_chtsz_reg[8]/P0002  & ~n2983 ;
  assign n4352 = n3050 & n4351 ;
  assign n4353 = \ctl_rf_c2_rf_chtsz_reg[8]/P0002  & n2983 ;
  assign n4354 = n3024 & n4353 ;
  assign n4355 = ~n4352 & ~n4354 ;
  assign n4356 = \ctl_rf_c7_rf_chtsz_reg[8]/P0002  & ~n2983 ;
  assign n4357 = n3011 & n4356 ;
  assign n4358 = \ctl_rf_c0_rf_chtsz_reg[8]/P0002  & n2983 ;
  assign n4359 = n3050 & n4358 ;
  assign n4360 = ~n4357 & ~n4359 ;
  assign n4361 = n4355 & n4360 ;
  assign n4362 = \ctl_rf_c3_rf_chtsz_reg[8]/P0002  & ~n2983 ;
  assign n4363 = n3024 & n4362 ;
  assign n4364 = \ctl_rf_c6_rf_chtsz_reg[8]/P0002  & n2983 ;
  assign n4365 = n3011 & n4364 ;
  assign n4366 = ~n4363 & ~n4365 ;
  assign n4367 = \ctl_rf_c4_rf_chtsz_reg[8]/P0002  & n2983 ;
  assign n4368 = n2999 & n4367 ;
  assign n4369 = \ctl_rf_c5_rf_chtsz_reg[8]/P0002  & ~n2983 ;
  assign n4370 = n2999 & n4369 ;
  assign n4371 = ~n4368 & ~n4370 ;
  assign n4372 = n4366 & n4371 ;
  assign n4373 = n4361 & n4372 ;
  assign n4374 = n4350 & n4373 ;
  assign n4375 = n4327 & n4374 ;
  assign n4376 = n4280 & n4375 ;
  assign n4377 = \ctl_rf_c1_rf_chtsz_reg[7]/NET0131  & ~n2983 ;
  assign n4378 = n3050 & n4377 ;
  assign n4379 = \ctl_rf_c2_rf_chtsz_reg[7]/NET0131  & n2983 ;
  assign n4380 = n3024 & n4379 ;
  assign n4381 = ~n4378 & ~n4380 ;
  assign n4382 = \ctl_rf_c7_rf_chtsz_reg[7]/NET0131  & ~n2983 ;
  assign n4383 = n3011 & n4382 ;
  assign n4384 = \ctl_rf_c0_rf_chtsz_reg[7]/NET0131  & n2983 ;
  assign n4385 = n3050 & n4384 ;
  assign n4386 = ~n4383 & ~n4385 ;
  assign n4387 = n4381 & n4386 ;
  assign n4388 = \ctl_rf_c3_rf_chtsz_reg[7]/NET0131  & ~n2983 ;
  assign n4389 = n3024 & n4388 ;
  assign n4390 = \ctl_rf_c6_rf_chtsz_reg[7]/NET0131  & n2983 ;
  assign n4391 = n3011 & n4390 ;
  assign n4392 = ~n4389 & ~n4391 ;
  assign n4393 = \ctl_rf_c4_rf_chtsz_reg[7]/NET0131  & n2983 ;
  assign n4394 = n2999 & n4393 ;
  assign n4395 = \ctl_rf_c5_rf_chtsz_reg[7]/NET0131  & ~n2983 ;
  assign n4396 = n2999 & n4395 ;
  assign n4397 = ~n4394 & ~n4396 ;
  assign n4398 = n4392 & n4397 ;
  assign n4399 = n4387 & n4398 ;
  assign n4400 = \ctl_rf_c1_rf_chtsz_reg[9]/P0002  & ~n2983 ;
  assign n4401 = n3050 & n4400 ;
  assign n4402 = \ctl_rf_c2_rf_chtsz_reg[9]/P0002  & n2983 ;
  assign n4403 = n3024 & n4402 ;
  assign n4404 = ~n4401 & ~n4403 ;
  assign n4405 = \ctl_rf_c7_rf_chtsz_reg[9]/P0002  & ~n2983 ;
  assign n4406 = n3011 & n4405 ;
  assign n4407 = \ctl_rf_c0_rf_chtsz_reg[9]/P0002  & n2983 ;
  assign n4408 = n3050 & n4407 ;
  assign n4409 = ~n4406 & ~n4408 ;
  assign n4410 = n4404 & n4409 ;
  assign n4411 = \ctl_rf_c3_rf_chtsz_reg[9]/P0002  & ~n2983 ;
  assign n4412 = n3024 & n4411 ;
  assign n4413 = \ctl_rf_c6_rf_chtsz_reg[9]/P0002  & n2983 ;
  assign n4414 = n3011 & n4413 ;
  assign n4415 = ~n4412 & ~n4414 ;
  assign n4416 = \ctl_rf_c4_rf_chtsz_reg[9]/P0002  & n2983 ;
  assign n4417 = n2999 & n4416 ;
  assign n4418 = \ctl_rf_c5_rf_chtsz_reg[9]/P0002  & ~n2983 ;
  assign n4419 = n2999 & n4418 ;
  assign n4420 = ~n4417 & ~n4419 ;
  assign n4421 = n4415 & n4420 ;
  assign n4422 = n4410 & n4421 ;
  assign n4423 = n4399 & n4422 ;
  assign n4424 = \ctl_rf_c1_rf_chtsz_reg[10]/P0002  & ~n2983 ;
  assign n4425 = n3050 & n4424 ;
  assign n4426 = \ctl_rf_c2_rf_chtsz_reg[10]/P0002  & n2983 ;
  assign n4427 = n3024 & n4426 ;
  assign n4428 = ~n4425 & ~n4427 ;
  assign n4429 = \ctl_rf_c7_rf_chtsz_reg[10]/P0002  & ~n2983 ;
  assign n4430 = n3011 & n4429 ;
  assign n4431 = \ctl_rf_c0_rf_chtsz_reg[10]/P0002  & n2983 ;
  assign n4432 = n3050 & n4431 ;
  assign n4433 = ~n4430 & ~n4432 ;
  assign n4434 = n4428 & n4433 ;
  assign n4435 = \ctl_rf_c3_rf_chtsz_reg[10]/P0002  & ~n2983 ;
  assign n4436 = n3024 & n4435 ;
  assign n4437 = \ctl_rf_c6_rf_chtsz_reg[10]/P0002  & n2983 ;
  assign n4438 = n3011 & n4437 ;
  assign n4439 = ~n4436 & ~n4438 ;
  assign n4440 = \ctl_rf_c4_rf_chtsz_reg[10]/P0002  & n2983 ;
  assign n4441 = n2999 & n4440 ;
  assign n4442 = \ctl_rf_c5_rf_chtsz_reg[10]/P0002  & ~n2983 ;
  assign n4443 = n2999 & n4442 ;
  assign n4444 = ~n4441 & ~n4443 ;
  assign n4445 = n4439 & n4444 ;
  assign n4446 = n4434 & n4445 ;
  assign n4447 = \ctl_rf_c1_rf_chtsz_reg[6]/NET0131  & ~n2983 ;
  assign n4448 = n3050 & n4447 ;
  assign n4449 = \ctl_rf_c2_rf_chtsz_reg[6]/NET0131  & n2983 ;
  assign n4450 = n3024 & n4449 ;
  assign n4451 = ~n4448 & ~n4450 ;
  assign n4452 = \ctl_rf_c7_rf_chtsz_reg[6]/NET0131  & ~n2983 ;
  assign n4453 = n3011 & n4452 ;
  assign n4454 = \ctl_rf_c0_rf_chtsz_reg[6]/NET0131  & n2983 ;
  assign n4455 = n3050 & n4454 ;
  assign n4456 = ~n4453 & ~n4455 ;
  assign n4457 = n4451 & n4456 ;
  assign n4458 = \ctl_rf_c3_rf_chtsz_reg[6]/NET0131  & ~n2983 ;
  assign n4459 = n3024 & n4458 ;
  assign n4460 = \ctl_rf_c6_rf_chtsz_reg[6]/NET0131  & n2983 ;
  assign n4461 = n3011 & n4460 ;
  assign n4462 = ~n4459 & ~n4461 ;
  assign n4463 = \ctl_rf_c4_rf_chtsz_reg[6]/NET0131  & n2983 ;
  assign n4464 = n2999 & n4463 ;
  assign n4465 = \ctl_rf_c5_rf_chtsz_reg[6]/NET0131  & ~n2983 ;
  assign n4466 = n2999 & n4465 ;
  assign n4467 = ~n4464 & ~n4466 ;
  assign n4468 = n4462 & n4467 ;
  assign n4469 = n4457 & n4468 ;
  assign n4470 = n4446 & n4469 ;
  assign n4471 = n4423 & n4470 ;
  assign n4472 = ~\de_de_st_reg[5]/NET0131  & ~\de_de_st_reg[6]/NET0131  ;
  assign n4473 = ~\de_de_st_reg[2]/NET0131  & n4472 ;
  assign n4474 = \de_de_st_reg[0]/NET0131  & ~\de_de_st_reg[1]/NET0131  ;
  assign n4475 = n4473 & n4474 ;
  assign n4476 = \ctl_rf_c1_rf_chtsz_reg[0]/P0002  & ~n2983 ;
  assign n4477 = n3050 & n4476 ;
  assign n4478 = \ctl_rf_c2_rf_chtsz_reg[0]/P0002  & n2983 ;
  assign n4479 = n3024 & n4478 ;
  assign n4480 = ~n4477 & ~n4479 ;
  assign n4481 = \ctl_rf_c7_rf_chtsz_reg[0]/P0002  & ~n2983 ;
  assign n4482 = n3011 & n4481 ;
  assign n4483 = \ctl_rf_c0_rf_chtsz_reg[0]/P0002  & n2983 ;
  assign n4484 = n3050 & n4483 ;
  assign n4485 = ~n4482 & ~n4484 ;
  assign n4486 = n4480 & n4485 ;
  assign n4487 = \ctl_rf_c3_rf_chtsz_reg[0]/P0002  & ~n2983 ;
  assign n4488 = n3024 & n4487 ;
  assign n4489 = \ctl_rf_c6_rf_chtsz_reg[0]/P0002  & n2983 ;
  assign n4490 = n3011 & n4489 ;
  assign n4491 = ~n4488 & ~n4490 ;
  assign n4492 = \ctl_rf_c4_rf_chtsz_reg[0]/P0002  & n2983 ;
  assign n4493 = n2999 & n4492 ;
  assign n4494 = \ctl_rf_c5_rf_chtsz_reg[0]/P0002  & ~n2983 ;
  assign n4495 = n2999 & n4494 ;
  assign n4496 = ~n4493 & ~n4495 ;
  assign n4497 = n4491 & n4496 ;
  assign n4498 = n4486 & n4497 ;
  assign n4499 = \ch_sel_arb_req_reg/NET0131  & ~n3105 ;
  assign n4500 = n4498 & n4499 ;
  assign n4501 = n4475 & n4500 ;
  assign n4502 = n4471 & n4501 ;
  assign n4503 = n4376 & n4502 ;
  assign n4504 = ~\ch_sel_arb_chcsr_reg_reg[1]/NET0131  & ~\ch_sel_arb_chcsr_reg_reg[2]/NET0131  ;
  assign n4505 = \ch_sel_arb_chcsr_reg_reg[1]/NET0131  & \ch_sel_arb_chcsr_reg_reg[2]/NET0131  ;
  assign n4506 = ~n4504 & ~n4505 ;
  assign n4507 = \de_tsz_cnt_reg[0]/NET0131  & ~\de_tsz_cnt_reg[1]/NET0131  ;
  assign n4508 = n2811 & n4507 ;
  assign n4509 = n2808 & n4508 ;
  assign n4510 = \de_bst_cnt_reg[0]/NET0131  & ~\de_bst_cnt_reg[4]/NET0131  ;
  assign n4511 = n2820 & n4510 ;
  assign n4512 = n2819 & n4511 ;
  assign n4513 = ~n4509 & ~n4512 ;
  assign n4514 = ~n4506 & ~n4513 ;
  assign n4515 = ~\de_de_st_reg[0]/NET0131  & \de_de_st_reg[1]/NET0131  ;
  assign n4516 = n4473 & n4515 ;
  assign n4517 = ~n4514 & n4516 ;
  assign n4518 = \ahb_mst1_mx_cmd_st_reg[1]/NET0131  & ~n2830 ;
  assign n4519 = n2915 & n4518 ;
  assign n4520 = ~n2799 & n4519 ;
  assign n4521 = \ahb_mst0_mx_cmd_st_reg[1]/NET0131  & \h0readyin_pad  ;
  assign n4522 = n2956 & n4521 ;
  assign n4523 = n4516 & ~n4522 ;
  assign n4524 = ~n4520 & n4523 ;
  assign n4525 = ~n4517 & ~n4524 ;
  assign n4526 = n4471 & n4500 ;
  assign n4527 = n4376 & n4526 ;
  assign n4528 = \ch_sel_arb_req_reg/NET0131  & n4475 ;
  assign n4529 = ~n3105 & n4528 ;
  assign n4530 = n4326 & n4529 ;
  assign n4531 = ~n4527 & n4530 ;
  assign n4532 = n4525 & ~n4531 ;
  assign n4533 = \ahb_mst0_mx_cmd_st_reg[0]/NET0131  & ~\ahb_mst0_mx_cmd_st_reg[1]/NET0131  ;
  assign n4534 = ~n2964 & ~n4533 ;
  assign n4535 = n2956 & ~n4533 ;
  assign n4536 = ~n2955 & n4535 ;
  assign n4537 = ~n4534 & ~n4536 ;
  assign n4538 = ~\h0req_pad  & ~n2944 ;
  assign n4539 = ~\ch_sel_arb_chcsr_reg_reg[2]/NET0131  & \de_de_st_reg[1]/NET0131  ;
  assign n4540 = \ch_sel_arb_chcsr_reg_reg[1]/NET0131  & n4539 ;
  assign n4541 = ~\de_de_st_reg[5]/NET0131  & \h0req_pad  ;
  assign n4542 = ~n4540 & n4541 ;
  assign n4543 = ~n2823 & n4541 ;
  assign n4544 = ~n2814 & n4543 ;
  assign n4545 = ~n4542 & ~n4544 ;
  assign n4546 = ~n4538 & n4545 ;
  assign n4547 = ~\de_de_st_reg[0]/NET0131  & ~\de_de_st_reg[1]/NET0131  ;
  assign n4548 = \de_de_st_reg[2]/NET0131  & n4472 ;
  assign n4549 = n4547 & n4548 ;
  assign n4550 = ~n4520 & ~n4522 ;
  assign n4551 = n4514 & n4516 ;
  assign n4552 = ~n4550 & n4551 ;
  assign n4553 = ~n4549 & ~n4552 ;
  assign n4554 = n3686 & n3690 ;
  assign n4555 = ~n3107 & ~n4554 ;
  assign n4556 = n3648 & n3658 ;
  assign n4557 = n3666 & n3669 ;
  assign n4558 = ~n4556 & n4557 ;
  assign n4559 = ~n3107 & n4558 ;
  assign n4560 = \ch_sel_fix_pri_sel_reg[0]/NET0131  & n3106 ;
  assign n4561 = ~n3097 & n4560 ;
  assign n4562 = ~n4559 & ~n4561 ;
  assign n4563 = ~n4555 & n4562 ;
  assign n4564 = ~\ch_sel_fix_pri_sel_reg[1]/NET0131  & n3106 ;
  assign n4565 = ~n3097 & n4564 ;
  assign n4566 = ~n3107 & n4557 ;
  assign n4567 = ~n4555 & n4566 ;
  assign n4568 = ~n4565 & ~n4567 ;
  assign n4569 = hsel_reg_pad & \htrans[1]_pad  ;
  assign n4570 = \hrdata_reg[16]_pad  & ~n4569 ;
  assign n4571 = ~\hsize[1]_pad  & ~\hsize[2]_pad  ;
  assign n4572 = \ctl_rf_m0end_reg/NET0131  & \hsize[0]_pad  ;
  assign n4573 = n4571 & n4572 ;
  assign n4574 = ~\haddr[4]_pad  & ~\haddr[5]_pad  ;
  assign n4575 = ~\haddr[6]_pad  & \haddr[7]_pad  ;
  assign n4576 = n4574 & n4575 ;
  assign n4577 = ~\haddr[2]_pad  & ~\haddr[3]_pad  ;
  assign n4578 = \ctl_rf_c4_rf_ch_en_reg/NET0131  & n4577 ;
  assign n4579 = \haddr[2]_pad  & ~\haddr[3]_pad  ;
  assign n4580 = \ctl_rf_c4_rf_int_tc1_msk_reg/NET0131  & n4579 ;
  assign n4581 = ~n4578 & ~n4580 ;
  assign n4582 = \haddr[2]_pad  & \haddr[3]_pad  ;
  assign n4583 = \ctl_rf_c4_rf_chdad_reg[0]/NET0131  & n4582 ;
  assign n4584 = ~\haddr[2]_pad  & \haddr[3]_pad  ;
  assign n4585 = \ctl_rf_c4_rf_chsad_reg[0]/NET0131  & n4584 ;
  assign n4586 = ~n4583 & ~n4585 ;
  assign n4587 = n4581 & n4586 ;
  assign n4588 = n4576 & ~n4587 ;
  assign n4589 = \haddr[6]_pad  & ~\haddr[7]_pad  ;
  assign n4590 = n4574 & n4589 ;
  assign n4591 = \ctl_rf_c2_rf_int_tc1_msk_reg/NET0131  & n4579 ;
  assign n4592 = \ctl_rf_c2_rf_chsad_reg[0]/NET0131  & n4584 ;
  assign n4593 = ~n4591 & ~n4592 ;
  assign n4594 = \ctl_rf_c2_rf_ch_en_reg/NET0131  & n4577 ;
  assign n4595 = \ctl_rf_c2_rf_chdad_reg[0]/NET0131  & n4582 ;
  assign n4596 = ~n4594 & ~n4595 ;
  assign n4597 = n4593 & n4596 ;
  assign n4598 = n4590 & ~n4597 ;
  assign n4599 = ~n4588 & ~n4598 ;
  assign n4600 = ~\haddr[4]_pad  & \haddr[5]_pad  ;
  assign n4601 = n4575 & n4600 ;
  assign n4602 = \ctl_rf_c5_rf_int_tc1_msk_reg/NET0131  & n4579 ;
  assign n4603 = \ctl_rf_c5_rf_chdad_reg[0]/NET0131  & n4582 ;
  assign n4604 = ~n4602 & ~n4603 ;
  assign n4605 = \ctl_rf_c5_rf_chsad_reg[0]/NET0131  & n4584 ;
  assign n4606 = \ctl_rf_c5_rf_ch_en_reg/NET0131  & n4577 ;
  assign n4607 = ~n4605 & ~n4606 ;
  assign n4608 = n4604 & n4607 ;
  assign n4609 = n4601 & ~n4608 ;
  assign n4610 = \haddr[6]_pad  & \haddr[7]_pad  ;
  assign n4611 = n4574 & n4610 ;
  assign n4612 = \ctl_rf_c6_rf_int_tc1_msk_reg/NET0131  & n4579 ;
  assign n4613 = \ctl_rf_c6_rf_chdad_reg[0]/NET0131  & n4582 ;
  assign n4614 = ~n4612 & ~n4613 ;
  assign n4615 = \ctl_rf_c6_rf_chsad_reg[0]/NET0131  & n4584 ;
  assign n4616 = \ctl_rf_c6_rf_ch_en_reg/NET0131  & n4577 ;
  assign n4617 = ~n4615 & ~n4616 ;
  assign n4618 = n4614 & n4617 ;
  assign n4619 = n4611 & ~n4618 ;
  assign n4620 = ~n4609 & ~n4619 ;
  assign n4621 = n4599 & n4620 ;
  assign n4622 = ~\haddr[6]_pad  & ~\haddr[7]_pad  ;
  assign n4623 = n4574 & n4622 ;
  assign n4624 = \ctl_rf_c0_rf_int_tc1_msk_reg/NET0131  & n4579 ;
  assign n4625 = \ctl_rf_c0_rf_chdad_reg[0]/NET0131  & n4582 ;
  assign n4626 = ~n4624 & ~n4625 ;
  assign n4627 = \ctl_rf_c0_rf_chsad_reg[0]/NET0131  & n4584 ;
  assign n4628 = \ctl_rf_c0_rf_ch_en_reg/NET0131  & n4577 ;
  assign n4629 = ~n4627 & ~n4628 ;
  assign n4630 = n4626 & n4629 ;
  assign n4631 = n4623 & ~n4630 ;
  assign n4632 = n4600 & n4622 ;
  assign n4633 = \ctl_rf_c1_rf_int_tc1_msk_reg/NET0131  & n4579 ;
  assign n4634 = \ctl_rf_c1_rf_chdad_reg[0]/NET0131  & n4582 ;
  assign n4635 = ~n4633 & ~n4634 ;
  assign n4636 = \ctl_rf_c1_rf_chsad_reg[0]/NET0131  & n4584 ;
  assign n4637 = \ctl_rf_c1_rf_ch_en_reg/NET0131  & n4577 ;
  assign n4638 = ~n4636 & ~n4637 ;
  assign n4639 = n4635 & n4638 ;
  assign n4640 = n4632 & ~n4639 ;
  assign n4641 = ~n4631 & ~n4640 ;
  assign n4642 = n4600 & n4610 ;
  assign n4643 = \ctl_rf_c7_rf_ch_en_reg/NET0131  & n4577 ;
  assign n4644 = \ctl_rf_c7_rf_int_tc1_msk_reg/NET0131  & n4579 ;
  assign n4645 = ~n4643 & ~n4644 ;
  assign n4646 = \ctl_rf_c7_rf_chdad_reg[0]/NET0131  & n4582 ;
  assign n4647 = \ctl_rf_c7_rf_chsad_reg[0]/NET0131  & n4584 ;
  assign n4648 = ~n4646 & ~n4647 ;
  assign n4649 = n4645 & n4648 ;
  assign n4650 = n4642 & ~n4649 ;
  assign n4651 = n4589 & n4600 ;
  assign n4652 = \ctl_rf_c3_rf_int_tc1_msk_reg/NET0131  & n4579 ;
  assign n4653 = \ctl_rf_c3_rf_chsad_reg[0]/NET0131  & n4584 ;
  assign n4654 = ~n4652 & ~n4653 ;
  assign n4655 = \ctl_rf_c3_rf_ch_en_reg/NET0131  & n4577 ;
  assign n4656 = \ctl_rf_c3_rf_chdad_reg[0]/NET0131  & n4582 ;
  assign n4657 = ~n4655 & ~n4656 ;
  assign n4658 = n4654 & n4657 ;
  assign n4659 = n4651 & ~n4658 ;
  assign n4660 = ~n4650 & ~n4659 ;
  assign n4661 = n4641 & n4660 ;
  assign n4662 = \haddr[4]_pad  & ~\haddr[5]_pad  ;
  assign n4663 = n4589 & n4662 ;
  assign n4664 = \ctl_rf_c2_rf_chllp_reg[0]/P0002  & n4577 ;
  assign n4665 = \ctl_rf_c2_rf_chtsz_reg[0]/P0002  & n4579 ;
  assign n4666 = ~n4664 & ~n4665 ;
  assign n4667 = n4663 & ~n4666 ;
  assign n4668 = \haddr[4]_pad  & \haddr[5]_pad  ;
  assign n4669 = n4610 & n4668 ;
  assign n4670 = \ctl_rf_c7_rf_chllp_reg[0]/P0002  & n4577 ;
  assign n4671 = \ctl_rf_c7_rf_chtsz_reg[0]/P0002  & n4579 ;
  assign n4672 = ~n4670 & ~n4671 ;
  assign n4673 = n4669 & ~n4672 ;
  assign n4674 = ~n4667 & ~n4673 ;
  assign n4675 = n4622 & n4662 ;
  assign n4676 = \ctl_rf_c0_rf_chllp_reg[0]/P0002  & n4577 ;
  assign n4677 = \ctl_rf_c0_rf_chtsz_reg[0]/P0002  & n4579 ;
  assign n4678 = ~n4676 & ~n4677 ;
  assign n4679 = n4675 & ~n4678 ;
  assign n4680 = n4575 & n4668 ;
  assign n4681 = \ctl_rf_c5_rf_chllp_reg[0]/P0002  & n4577 ;
  assign n4682 = \ctl_rf_c5_rf_chtsz_reg[0]/P0002  & n4579 ;
  assign n4683 = ~n4681 & ~n4682 ;
  assign n4684 = n4680 & ~n4683 ;
  assign n4685 = ~n4679 & ~n4684 ;
  assign n4686 = n4674 & n4685 ;
  assign n4687 = n4575 & n4662 ;
  assign n4688 = \ctl_rf_c4_rf_chllp_reg[0]/P0002  & n4577 ;
  assign n4689 = \ctl_rf_c4_rf_chtsz_reg[0]/P0002  & n4579 ;
  assign n4690 = ~n4688 & ~n4689 ;
  assign n4691 = n4687 & ~n4690 ;
  assign n4692 = n4622 & n4668 ;
  assign n4693 = \ctl_rf_c1_rf_chllp_reg[0]/P0002  & n4577 ;
  assign n4694 = \ctl_rf_c1_rf_chtsz_reg[0]/P0002  & n4579 ;
  assign n4695 = ~n4693 & ~n4694 ;
  assign n4696 = n4692 & ~n4695 ;
  assign n4697 = ~n4691 & ~n4696 ;
  assign n4698 = n4589 & n4668 ;
  assign n4699 = \ctl_rf_c3_rf_chllp_reg[0]/P0002  & n4577 ;
  assign n4700 = \ctl_rf_c3_rf_chtsz_reg[0]/P0002  & n4579 ;
  assign n4701 = ~n4699 & ~n4700 ;
  assign n4702 = n4698 & ~n4701 ;
  assign n4703 = n4610 & n4662 ;
  assign n4704 = \ctl_rf_c6_rf_chllp_reg[0]/P0002  & n4577 ;
  assign n4705 = \ctl_rf_c6_rf_chtsz_reg[0]/P0002  & n4579 ;
  assign n4706 = ~n4704 & ~n4705 ;
  assign n4707 = n4703 & ~n4706 ;
  assign n4708 = ~n4702 & ~n4707 ;
  assign n4709 = n4697 & n4708 ;
  assign n4710 = n4686 & n4709 ;
  assign n4711 = n4661 & n4710 ;
  assign n4712 = n4621 & n4711 ;
  assign n4713 = \haddr[8]_pad  & ~n4712 ;
  assign n4714 = ~\haddr[8]_pad  & n4622 ;
  assign n4715 = n4577 & n4600 ;
  assign n4716 = ~\de_de_st_reg[0]/NET0131  & n4715 ;
  assign n4717 = n2983 & n4716 ;
  assign n4718 = n3050 & n4717 ;
  assign n4719 = n4579 & n4662 ;
  assign n4720 = \ctl_rf_tc_reg[0]/NET0131  & n4719 ;
  assign n4721 = ~\haddr[3]_pad  & n4574 ;
  assign n4722 = ~\ctl_rf_c0_rf_int_tc1_msk_reg/NET0131  & \ctl_rf_tc_reg[0]/NET0131  ;
  assign n4723 = n4721 & n4722 ;
  assign n4724 = ~n4720 & ~n4723 ;
  assign n4725 = n4584 & n4600 ;
  assign n4726 = \ctl_rf_sync_reg[0]/NET0131  & n4725 ;
  assign n4727 = n4582 & n4662 ;
  assign n4728 = \ctl_rf_c0_rf_ch_en_reg/NET0131  & n4727 ;
  assign n4729 = ~n4726 & ~n4728 ;
  assign n4730 = n4579 & n4600 ;
  assign n4731 = \ctl_rf_dmacen_reg/NET0131  & n4730 ;
  assign n4732 = \ctl_rf_abt_reg[0]/NET0131  & ~\ctl_rf_c0_rf_int_abt_msk_reg/NET0131  ;
  assign n4733 = n4574 & n4577 ;
  assign n4734 = n4732 & n4733 ;
  assign n4735 = ~n4731 & ~n4734 ;
  assign n4736 = n4729 & n4735 ;
  assign n4737 = n4724 & n4736 ;
  assign n4738 = ~n4718 & n4737 ;
  assign n4739 = n4714 & ~n4738 ;
  assign n4740 = n4573 & ~n4739 ;
  assign n4741 = ~n4713 & n4740 ;
  assign n4742 = n4569 & ~n4741 ;
  assign n4743 = n4573 & n4742 ;
  assign n4744 = \ctl_rf_m0end_reg/NET0131  & ~\hsize[0]_pad  ;
  assign n4745 = n4571 & n4744 ;
  assign n4746 = ~\haddr[8]_pad  & n4745 ;
  assign n4747 = ~\de_de_st_reg[0]/NET0131  & n4579 ;
  assign n4748 = ~n2983 & n4747 ;
  assign n4749 = n3011 & n4748 ;
  assign n4750 = \ctl_rf_c7_rf_chsad_reg[8]/P0002  & n4584 ;
  assign n4751 = \ctl_rf_c7_rf_dwidth_reg[0]/NET0131  & n4577 ;
  assign n4752 = \ctl_rf_c7_rf_chdad_reg[8]/NET0131  & n4582 ;
  assign n4753 = ~n4751 & ~n4752 ;
  assign n4754 = ~n4750 & n4753 ;
  assign n4755 = ~n4749 & n4754 ;
  assign n4756 = n4642 & ~n4755 ;
  assign n4757 = \ctl_rf_c6_rf_chllp_reg[8]/NET0131  & n4577 ;
  assign n4758 = \ctl_rf_c6_rf_chtsz_reg[8]/P0002  & n4579 ;
  assign n4759 = ~n4757 & ~n4758 ;
  assign n4760 = n4703 & ~n4759 ;
  assign n4761 = \ctl_rf_c3_rf_chllp_reg[8]/NET0131  & n4577 ;
  assign n4762 = \ctl_rf_c3_rf_chtsz_reg[8]/P0002  & n4579 ;
  assign n4763 = ~n4761 & ~n4762 ;
  assign n4764 = n4698 & ~n4763 ;
  assign n4765 = ~n4760 & ~n4764 ;
  assign n4766 = \ctl_rf_c7_rf_chllp_reg[8]/NET0131  & n4577 ;
  assign n4767 = \ctl_rf_c7_rf_chtsz_reg[8]/P0002  & n4579 ;
  assign n4768 = ~n4766 & ~n4767 ;
  assign n4769 = n4669 & ~n4768 ;
  assign n4770 = \ctl_rf_c4_rf_chllp_reg[8]/NET0131  & n4577 ;
  assign n4771 = \ctl_rf_c4_rf_chtsz_reg[8]/P0002  & n4579 ;
  assign n4772 = ~n4770 & ~n4771 ;
  assign n4773 = n4687 & ~n4772 ;
  assign n4774 = ~n4769 & ~n4773 ;
  assign n4775 = n4765 & n4774 ;
  assign n4776 = \ctl_rf_c2_rf_chllp_reg[8]/NET0131  & n4577 ;
  assign n4777 = \ctl_rf_c2_rf_chtsz_reg[8]/P0002  & n4579 ;
  assign n4778 = ~n4776 & ~n4777 ;
  assign n4779 = n4663 & ~n4778 ;
  assign n4780 = \ctl_rf_c0_rf_chllp_reg[8]/NET0131  & n4577 ;
  assign n4781 = \ctl_rf_c0_rf_chtsz_reg[8]/P0002  & n4579 ;
  assign n4782 = ~n4780 & ~n4781 ;
  assign n4783 = n4675 & ~n4782 ;
  assign n4784 = ~n4779 & ~n4783 ;
  assign n4785 = \ctl_rf_c1_rf_chllp_reg[8]/NET0131  & n4577 ;
  assign n4786 = \ctl_rf_c1_rf_chtsz_reg[8]/P0002  & n4579 ;
  assign n4787 = ~n4785 & ~n4786 ;
  assign n4788 = n4692 & ~n4787 ;
  assign n4789 = \ctl_rf_c5_rf_chllp_reg[8]/NET0131  & n4577 ;
  assign n4790 = \ctl_rf_c5_rf_chtsz_reg[8]/P0002  & n4579 ;
  assign n4791 = ~n4789 & ~n4790 ;
  assign n4792 = n4680 & ~n4791 ;
  assign n4793 = ~n4788 & ~n4792 ;
  assign n4794 = n4784 & n4793 ;
  assign n4795 = n4775 & n4794 ;
  assign n4796 = ~n4756 & n4795 ;
  assign n4797 = n2983 & n4747 ;
  assign n4798 = n3011 & n4797 ;
  assign n4799 = \ctl_rf_c6_rf_chsad_reg[8]/P0002  & n4584 ;
  assign n4800 = \ctl_rf_c6_rf_dwidth_reg[0]/NET0131  & n4577 ;
  assign n4801 = \ctl_rf_c6_rf_chdad_reg[8]/NET0131  & n4582 ;
  assign n4802 = ~n4800 & ~n4801 ;
  assign n4803 = ~n4799 & n4802 ;
  assign n4804 = ~n4798 & n4803 ;
  assign n4805 = n4611 & ~n4804 ;
  assign n4806 = n3050 & n4748 ;
  assign n4807 = \ctl_rf_c1_rf_chsad_reg[8]/P0002  & n4584 ;
  assign n4808 = \ctl_rf_c1_rf_chdad_reg[8]/NET0131  & n4582 ;
  assign n4809 = \ctl_rf_c1_rf_dwidth_reg[0]/NET0131  & n4577 ;
  assign n4810 = ~n4808 & ~n4809 ;
  assign n4811 = ~n4807 & n4810 ;
  assign n4812 = ~n4806 & n4811 ;
  assign n4813 = n4632 & ~n4812 ;
  assign n4814 = ~n4805 & ~n4813 ;
  assign n4815 = n2999 & n4748 ;
  assign n4816 = \ctl_rf_c5_rf_chsad_reg[8]/P0002  & n4584 ;
  assign n4817 = \ctl_rf_c5_rf_chdad_reg[8]/NET0131  & n4582 ;
  assign n4818 = \ctl_rf_c5_rf_dwidth_reg[0]/NET0131  & n4577 ;
  assign n4819 = ~n4817 & ~n4818 ;
  assign n4820 = ~n4816 & n4819 ;
  assign n4821 = ~n4815 & n4820 ;
  assign n4822 = n4601 & ~n4821 ;
  assign n4823 = n3024 & n4797 ;
  assign n4824 = \ctl_rf_c2_rf_chsad_reg[8]/P0002  & n4584 ;
  assign n4825 = \ctl_rf_c2_rf_dwidth_reg[0]/NET0131  & n4577 ;
  assign n4826 = \ctl_rf_c2_rf_chdad_reg[8]/NET0131  & n4582 ;
  assign n4827 = ~n4825 & ~n4826 ;
  assign n4828 = ~n4824 & n4827 ;
  assign n4829 = ~n4823 & n4828 ;
  assign n4830 = n4590 & ~n4829 ;
  assign n4831 = ~n4822 & ~n4830 ;
  assign n4832 = n4814 & n4831 ;
  assign n4833 = n4796 & n4832 ;
  assign n4834 = n3050 & n4797 ;
  assign n4835 = \ctl_rf_c0_rf_chsad_reg[8]/P0002  & n4584 ;
  assign n4836 = \ctl_rf_c0_rf_chdad_reg[8]/NET0131  & n4582 ;
  assign n4837 = \ctl_rf_c0_rf_dwidth_reg[0]/NET0131  & n4577 ;
  assign n4838 = ~n4836 & ~n4837 ;
  assign n4839 = ~n4835 & n4838 ;
  assign n4840 = ~n4834 & n4839 ;
  assign n4841 = n4623 & ~n4840 ;
  assign n4842 = n3024 & n4748 ;
  assign n4843 = \ctl_rf_c3_rf_chsad_reg[8]/P0002  & n4584 ;
  assign n4844 = \ctl_rf_c3_rf_dwidth_reg[0]/NET0131  & n4577 ;
  assign n4845 = \ctl_rf_c3_rf_chdad_reg[8]/NET0131  & n4582 ;
  assign n4846 = ~n4844 & ~n4845 ;
  assign n4847 = ~n4843 & n4846 ;
  assign n4848 = ~n4842 & n4847 ;
  assign n4849 = n4651 & ~n4848 ;
  assign n4850 = n2999 & n4797 ;
  assign n4851 = \ctl_rf_c4_rf_chsad_reg[8]/P0002  & n4584 ;
  assign n4852 = \ctl_rf_c4_rf_chdad_reg[8]/NET0131  & n4582 ;
  assign n4853 = \ctl_rf_c4_rf_dwidth_reg[0]/NET0131  & n4577 ;
  assign n4854 = ~n4852 & ~n4853 ;
  assign n4855 = ~n4851 & n4854 ;
  assign n4856 = ~n4850 & n4855 ;
  assign n4857 = n4576 & ~n4856 ;
  assign n4858 = ~n4849 & ~n4857 ;
  assign n4859 = ~n4841 & n4858 ;
  assign n4860 = n4745 & n4859 ;
  assign n4861 = n4833 & n4860 ;
  assign n4862 = ~n4746 & ~n4861 ;
  assign n4863 = \ctl_rf_c0_rf_src_sz_reg[0]/NET0131  & n4577 ;
  assign n4864 = \ctl_rf_c0_rf_chllp_cnt_reg[0]/NET0131  & n4579 ;
  assign n4865 = ~n4863 & ~n4864 ;
  assign n4866 = \ctl_rf_c0_rf_chsad_reg[16]/NET0131  & n4584 ;
  assign n4867 = \ctl_rf_c0_rf_chdad_reg[16]/NET0131  & n4582 ;
  assign n4868 = ~n4866 & ~n4867 ;
  assign n4869 = n4865 & n4868 ;
  assign n4870 = n4623 & ~n4869 ;
  assign n4871 = \haddr[8]_pad  & ~n4870 ;
  assign n4872 = \ctl_rf_c2_rf_chllp_cnt_reg[0]/NET0131  & n4579 ;
  assign n4873 = \ctl_rf_c2_rf_chdad_reg[16]/NET0131  & n4582 ;
  assign n4874 = ~n4872 & ~n4873 ;
  assign n4875 = \ctl_rf_c2_rf_chsad_reg[16]/NET0131  & n4584 ;
  assign n4876 = \ctl_rf_c2_rf_src_sz_reg[0]/NET0131  & n4577 ;
  assign n4877 = ~n4875 & ~n4876 ;
  assign n4878 = n4874 & n4877 ;
  assign n4879 = n4590 & ~n4878 ;
  assign n4880 = \ctl_rf_c6_rf_chllp_cnt_reg[0]/NET0131  & n4579 ;
  assign n4881 = \ctl_rf_c6_rf_chsad_reg[16]/NET0131  & n4584 ;
  assign n4882 = ~n4880 & ~n4881 ;
  assign n4883 = \ctl_rf_c6_rf_src_sz_reg[0]/NET0131  & n4577 ;
  assign n4884 = \ctl_rf_c6_rf_chdad_reg[16]/NET0131  & n4582 ;
  assign n4885 = ~n4883 & ~n4884 ;
  assign n4886 = n4882 & n4885 ;
  assign n4887 = n4611 & ~n4886 ;
  assign n4888 = ~n4879 & ~n4887 ;
  assign n4889 = \ctl_rf_c1_rf_src_sz_reg[0]/NET0131  & n4577 ;
  assign n4890 = \ctl_rf_c1_rf_chllp_cnt_reg[0]/NET0131  & n4579 ;
  assign n4891 = ~n4889 & ~n4890 ;
  assign n4892 = \ctl_rf_c1_rf_chdad_reg[16]/NET0131  & n4582 ;
  assign n4893 = \ctl_rf_c1_rf_chsad_reg[16]/NET0131  & n4584 ;
  assign n4894 = ~n4892 & ~n4893 ;
  assign n4895 = n4891 & n4894 ;
  assign n4896 = n4632 & ~n4895 ;
  assign n4897 = \ctl_rf_c7_rf_chllp_cnt_reg[0]/NET0131  & n4579 ;
  assign n4898 = \ctl_rf_c7_rf_chdad_reg[16]/NET0131  & n4582 ;
  assign n4899 = ~n4897 & ~n4898 ;
  assign n4900 = \ctl_rf_c7_rf_chsad_reg[16]/NET0131  & n4584 ;
  assign n4901 = \ctl_rf_c7_rf_src_sz_reg[0]/NET0131  & n4577 ;
  assign n4902 = ~n4900 & ~n4901 ;
  assign n4903 = n4899 & n4902 ;
  assign n4904 = n4642 & ~n4903 ;
  assign n4905 = ~n4896 & ~n4904 ;
  assign n4906 = n4888 & n4905 ;
  assign n4907 = n4871 & n4906 ;
  assign n4908 = \ctl_rf_c1_rf_chllp_reg[16]/NET0131  & n4692 ;
  assign n4909 = \ctl_rf_c3_rf_chllp_reg[16]/NET0131  & n4698 ;
  assign n4910 = ~n4908 & ~n4909 ;
  assign n4911 = \ctl_rf_c0_rf_chllp_reg[16]/NET0131  & n4675 ;
  assign n4912 = \ctl_rf_c4_rf_chllp_reg[16]/NET0131  & n4687 ;
  assign n4913 = ~n4911 & ~n4912 ;
  assign n4914 = n4910 & n4913 ;
  assign n4915 = \ctl_rf_c6_rf_chllp_reg[16]/NET0131  & n4703 ;
  assign n4916 = \ctl_rf_c5_rf_chllp_reg[16]/NET0131  & n4680 ;
  assign n4917 = ~n4915 & ~n4916 ;
  assign n4918 = \ctl_rf_c2_rf_chllp_reg[16]/NET0131  & n4663 ;
  assign n4919 = \ctl_rf_c7_rf_chllp_reg[16]/NET0131  & n4669 ;
  assign n4920 = ~n4918 & ~n4919 ;
  assign n4921 = n4917 & n4920 ;
  assign n4922 = n4914 & n4921 ;
  assign n4923 = n4577 & ~n4922 ;
  assign n4924 = \ctl_rf_c4_rf_src_sz_reg[0]/NET0131  & n4577 ;
  assign n4925 = \ctl_rf_c4_rf_chsad_reg[16]/NET0131  & n4584 ;
  assign n4926 = ~n4924 & ~n4925 ;
  assign n4927 = \ctl_rf_c4_rf_chllp_cnt_reg[0]/NET0131  & n4579 ;
  assign n4928 = \ctl_rf_c4_rf_chdad_reg[16]/NET0131  & n4582 ;
  assign n4929 = ~n4927 & ~n4928 ;
  assign n4930 = n4926 & n4929 ;
  assign n4931 = n4576 & ~n4930 ;
  assign n4932 = \ctl_rf_c5_rf_chllp_cnt_reg[0]/NET0131  & n4579 ;
  assign n4933 = \ctl_rf_c5_rf_chdad_reg[16]/NET0131  & n4582 ;
  assign n4934 = ~n4932 & ~n4933 ;
  assign n4935 = \ctl_rf_c5_rf_chsad_reg[16]/NET0131  & n4584 ;
  assign n4936 = \ctl_rf_c5_rf_src_sz_reg[0]/NET0131  & n4577 ;
  assign n4937 = ~n4935 & ~n4936 ;
  assign n4938 = n4934 & n4937 ;
  assign n4939 = n4601 & ~n4938 ;
  assign n4940 = \ctl_rf_c3_rf_chllp_cnt_reg[0]/NET0131  & n4579 ;
  assign n4941 = \ctl_rf_c3_rf_chsad_reg[16]/NET0131  & n4584 ;
  assign n4942 = ~n4940 & ~n4941 ;
  assign n4943 = \ctl_rf_c3_rf_src_sz_reg[0]/NET0131  & n4577 ;
  assign n4944 = \ctl_rf_c3_rf_chdad_reg[16]/NET0131  & n4582 ;
  assign n4945 = ~n4943 & ~n4944 ;
  assign n4946 = n4942 & n4945 ;
  assign n4947 = n4651 & ~n4946 ;
  assign n4948 = ~n4939 & ~n4947 ;
  assign n4949 = ~n4931 & n4948 ;
  assign n4950 = ~n4923 & n4949 ;
  assign n4951 = n4907 & n4950 ;
  assign n4952 = \ctl_rf_c4dmabs_reg[16]/NET0131  & \haddr[4]_pad  ;
  assign n4953 = n4577 & n4952 ;
  assign n4954 = \ctl_rf_c5dmabs_reg[16]/NET0131  & \haddr[4]_pad  ;
  assign n4955 = n4579 & n4954 ;
  assign n4956 = ~n4953 & ~n4955 ;
  assign n4957 = \ctl_rf_c0dmabs_reg[16]/NET0131  & ~\haddr[4]_pad  ;
  assign n4958 = n4577 & n4957 ;
  assign n4959 = \ctl_rf_c6dmabs_reg[16]/NET0131  & \haddr[4]_pad  ;
  assign n4960 = n4584 & n4959 ;
  assign n4961 = ~n4958 & ~n4960 ;
  assign n4962 = n4956 & n4961 ;
  assign n4963 = \ctl_rf_c7dmabs_reg[16]/NET0131  & \haddr[4]_pad  ;
  assign n4964 = n4582 & n4963 ;
  assign n4965 = \ctl_rf_c2dmabs_reg[16]/NET0131  & ~\haddr[4]_pad  ;
  assign n4966 = n4584 & n4965 ;
  assign n4967 = ~n4964 & ~n4966 ;
  assign n4968 = \ctl_rf_c1dmabs_reg[16]/NET0131  & ~\haddr[4]_pad  ;
  assign n4969 = n4579 & n4968 ;
  assign n4970 = \ctl_rf_c3dmabs_reg[16]/NET0131  & ~\haddr[4]_pad  ;
  assign n4971 = n4582 & n4970 ;
  assign n4972 = ~n4969 & ~n4971 ;
  assign n4973 = n4967 & n4972 ;
  assign n4974 = n4962 & n4973 ;
  assign n4975 = n4589 & ~n4974 ;
  assign n4976 = \ctl_rf_c1brbs_reg[16]/NET0131  & ~\haddr[4]_pad  ;
  assign n4977 = n4579 & n4976 ;
  assign n4978 = \ctl_rf_c5brbs_reg[16]/NET0131  & \haddr[4]_pad  ;
  assign n4979 = n4579 & n4978 ;
  assign n4980 = ~n4977 & ~n4979 ;
  assign n4981 = \ctl_rf_c0brbs_reg[16]/NET0131  & ~\haddr[4]_pad  ;
  assign n4982 = n4577 & n4981 ;
  assign n4983 = \ctl_rf_c7brbs_reg[16]/NET0131  & \haddr[4]_pad  ;
  assign n4984 = n4582 & n4983 ;
  assign n4985 = ~n4982 & ~n4984 ;
  assign n4986 = n4980 & n4985 ;
  assign n4987 = \ctl_rf_c6brbs_reg[16]/NET0131  & \haddr[4]_pad  ;
  assign n4988 = n4584 & n4987 ;
  assign n4989 = \ctl_rf_c2brbs_reg[16]/NET0131  & ~\haddr[4]_pad  ;
  assign n4990 = n4584 & n4989 ;
  assign n4991 = ~n4988 & ~n4990 ;
  assign n4992 = \ctl_rf_c4brbs_reg[16]/NET0131  & \haddr[4]_pad  ;
  assign n4993 = n4577 & n4992 ;
  assign n4994 = \ctl_rf_c3brbs_reg[16]/NET0131  & ~\haddr[4]_pad  ;
  assign n4995 = n4582 & n4994 ;
  assign n4996 = ~n4993 & ~n4995 ;
  assign n4997 = n4991 & n4996 ;
  assign n4998 = n4986 & n4997 ;
  assign n4999 = n4575 & ~n4998 ;
  assign n5000 = \ctl_rf_abt_reg[0]/NET0131  & n4622 ;
  assign n5001 = ~\haddr[8]_pad  & ~n5000 ;
  assign n5002 = n4574 & n4582 ;
  assign n5003 = ~\ctl_rf_c0_rf_int_abt_msk_reg/NET0131  & n5002 ;
  assign n5004 = n4584 & n4662 ;
  assign n5005 = ~\haddr[8]_pad  & ~n5004 ;
  assign n5006 = ~n5003 & n5005 ;
  assign n5007 = ~n5001 & ~n5006 ;
  assign n5008 = ~n4999 & ~n5007 ;
  assign n5009 = ~n4975 & n5008 ;
  assign n5010 = ~n4951 & ~n5009 ;
  assign n5011 = ~n4745 & ~n5010 ;
  assign n5012 = n4742 & ~n5011 ;
  assign n5013 = n4862 & n5012 ;
  assign n5014 = ~n4743 & ~n5013 ;
  assign n5015 = ~n4570 & n5014 ;
  assign n5016 = \hrdata_reg[8]_pad  & ~n4569 ;
  assign n5017 = n4569 & ~n4573 ;
  assign n5018 = \ctl_rf_c3_rf_chllp_reg[24]/NET0131  & n4698 ;
  assign n5019 = \ctl_rf_c5_rf_chllp_reg[24]/NET0131  & n4680 ;
  assign n5020 = \ctl_rf_c2_rf_chllp_reg[24]/NET0131  & n4663 ;
  assign n5021 = ~n5019 & ~n5020 ;
  assign n5022 = ~n5018 & n5021 ;
  assign n5023 = \ctl_rf_c0_rf_chllp_reg[24]/NET0131  & n4675 ;
  assign n5024 = \ctl_rf_c1_rf_chllp_reg[24]/NET0131  & n4692 ;
  assign n5025 = ~n5023 & ~n5024 ;
  assign n5026 = \ctl_rf_c4_rf_chllp_reg[24]/NET0131  & n4687 ;
  assign n5027 = \ctl_rf_c7_rf_chllp_reg[24]/NET0131  & n4669 ;
  assign n5028 = ~n5026 & ~n5027 ;
  assign n5029 = \ctl_rf_c1_rf_dreqmode_reg/NET0131  & n4632 ;
  assign n5030 = \ctl_rf_c6_rf_chllp_reg[24]/NET0131  & n4703 ;
  assign n5031 = ~n5029 & ~n5030 ;
  assign n5032 = n5028 & n5031 ;
  assign n5033 = n5025 & n5032 ;
  assign n5034 = n5022 & n5033 ;
  assign n5035 = n4577 & ~n5034 ;
  assign n5036 = \ctl_rf_c6_rf_chdad_reg[24]/P0002  & n4582 ;
  assign n5037 = \ctl_rf_c6_rf_chsad_reg[24]/NET0131  & n4584 ;
  assign n5038 = \ctl_rf_c6_rf_dreqmode_reg/NET0131  & n4577 ;
  assign n5039 = ~n5037 & ~n5038 ;
  assign n5040 = ~n5036 & n5039 ;
  assign n5041 = n4611 & ~n5040 ;
  assign n5042 = \ctl_rf_c7_rf_chdad_reg[24]/P0002  & n4582 ;
  assign n5043 = \ctl_rf_c7_rf_chsad_reg[24]/NET0131  & n4584 ;
  assign n5044 = \ctl_rf_c7_rf_dreqmode_reg/NET0131  & n4577 ;
  assign n5045 = ~n5043 & ~n5044 ;
  assign n5046 = ~n5042 & n5045 ;
  assign n5047 = n4642 & ~n5046 ;
  assign n5048 = ~n5041 & ~n5047 ;
  assign n5049 = \ctl_rf_c0_rf_dreqmode_reg/NET0131  & n4577 ;
  assign n5050 = \ctl_rf_c0_rf_chsad_reg[24]/NET0131  & n4584 ;
  assign n5051 = \ctl_rf_c0_rf_chdad_reg[24]/P0002  & n4582 ;
  assign n5052 = ~n5050 & ~n5051 ;
  assign n5053 = ~n5049 & n5052 ;
  assign n5054 = n4623 & ~n5053 ;
  assign n5055 = \ctl_rf_c5_rf_chdad_reg[24]/P0002  & n4582 ;
  assign n5056 = \ctl_rf_c5_rf_chsad_reg[24]/NET0131  & n4584 ;
  assign n5057 = \ctl_rf_c5_rf_dreqmode_reg/NET0131  & n4577 ;
  assign n5058 = ~n5056 & ~n5057 ;
  assign n5059 = ~n5055 & n5058 ;
  assign n5060 = n4601 & ~n5059 ;
  assign n5061 = ~n5054 & ~n5060 ;
  assign n5062 = n5048 & n5061 ;
  assign n5063 = \ctl_rf_c3_rf_chdad_reg[24]/P0002  & n4582 ;
  assign n5064 = \ctl_rf_c3_rf_chsad_reg[24]/NET0131  & n4584 ;
  assign n5065 = \ctl_rf_c3_rf_dreqmode_reg/NET0131  & n4577 ;
  assign n5066 = ~n5064 & ~n5065 ;
  assign n5067 = ~n5063 & n5066 ;
  assign n5068 = n4651 & ~n5067 ;
  assign n5069 = \ctl_rf_c1_rf_chdad_reg[24]/P0002  & n4582 ;
  assign n5070 = \ctl_rf_c1_rf_chsad_reg[24]/NET0131  & n4584 ;
  assign n5071 = ~n5069 & ~n5070 ;
  assign n5072 = n4632 & ~n5071 ;
  assign n5073 = \haddr[8]_pad  & ~n5072 ;
  assign n5074 = ~n5068 & n5073 ;
  assign n5075 = \ctl_rf_c4_rf_dreqmode_reg/NET0131  & n4577 ;
  assign n5076 = \ctl_rf_c4_rf_chdad_reg[24]/P0002  & n4582 ;
  assign n5077 = \ctl_rf_c4_rf_chsad_reg[24]/NET0131  & n4584 ;
  assign n5078 = ~n5076 & ~n5077 ;
  assign n5079 = ~n5075 & n5078 ;
  assign n5080 = n4576 & ~n5079 ;
  assign n5081 = \ctl_rf_c2_rf_dreqmode_reg/NET0131  & n4577 ;
  assign n5082 = \ctl_rf_c2_rf_chsad_reg[24]/NET0131  & n4584 ;
  assign n5083 = \ctl_rf_c2_rf_chdad_reg[24]/P0002  & n4582 ;
  assign n5084 = ~n5082 & ~n5083 ;
  assign n5085 = ~n5081 & n5084 ;
  assign n5086 = n4590 & ~n5085 ;
  assign n5087 = ~n5080 & ~n5086 ;
  assign n5088 = n5074 & n5087 ;
  assign n5089 = n5062 & n5088 ;
  assign n5090 = ~n5035 & n5089 ;
  assign n5091 = \ctl_rf_c5brbs_reg[24]/NET0131  & \haddr[4]_pad  ;
  assign n5092 = n4579 & n5091 ;
  assign n5093 = \ctl_rf_c6brbs_reg[24]/NET0131  & \haddr[4]_pad  ;
  assign n5094 = n4584 & n5093 ;
  assign n5095 = ~n5092 & ~n5094 ;
  assign n5096 = \ctl_rf_c2brbs_reg[24]/NET0131  & ~\haddr[4]_pad  ;
  assign n5097 = n4584 & n5096 ;
  assign n5098 = \ctl_rf_c4brbs_reg[24]/NET0131  & \haddr[4]_pad  ;
  assign n5099 = n4577 & n5098 ;
  assign n5100 = ~n5097 & ~n5099 ;
  assign n5101 = n5095 & n5100 ;
  assign n5102 = \ctl_rf_c3brbs_reg[24]/NET0131  & ~\haddr[4]_pad  ;
  assign n5103 = n4582 & n5102 ;
  assign n5104 = \ctl_rf_c1brbs_reg[24]/NET0131  & ~\haddr[4]_pad  ;
  assign n5105 = n4579 & n5104 ;
  assign n5106 = ~n5103 & ~n5105 ;
  assign n5107 = \ctl_rf_c0brbs_reg[24]/NET0131  & ~\haddr[4]_pad  ;
  assign n5108 = n4577 & n5107 ;
  assign n5109 = \ctl_rf_c7brbs_reg[24]/NET0131  & \haddr[4]_pad  ;
  assign n5110 = n4582 & n5109 ;
  assign n5111 = ~n5108 & ~n5110 ;
  assign n5112 = n5106 & n5111 ;
  assign n5113 = n5101 & n5112 ;
  assign n5114 = n4575 & ~n5113 ;
  assign n5115 = \ctl_rf_c2dmabs_reg[24]/NET0131  & ~\haddr[4]_pad  ;
  assign n5116 = n4584 & n5115 ;
  assign n5117 = \ctl_rf_c6dmabs_reg[24]/NET0131  & \haddr[4]_pad  ;
  assign n5118 = n4584 & n5117 ;
  assign n5119 = ~n5116 & ~n5118 ;
  assign n5120 = \ctl_rf_c1dmabs_reg[24]/NET0131  & ~\haddr[4]_pad  ;
  assign n5121 = n4579 & n5120 ;
  assign n5122 = \ctl_rf_c3dmabs_reg[24]/NET0131  & ~\haddr[4]_pad  ;
  assign n5123 = n4582 & n5122 ;
  assign n5124 = ~n5121 & ~n5123 ;
  assign n5125 = n5119 & n5124 ;
  assign n5126 = \ctl_rf_c4dmabs_reg[24]/NET0131  & \haddr[4]_pad  ;
  assign n5127 = n4577 & n5126 ;
  assign n5128 = \ctl_rf_c0dmabs_reg[24]/NET0131  & ~\haddr[4]_pad  ;
  assign n5129 = n4577 & n5128 ;
  assign n5130 = ~n5127 & ~n5129 ;
  assign n5131 = \ctl_rf_c5dmabs_reg[24]/NET0131  & \haddr[4]_pad  ;
  assign n5132 = n4579 & n5131 ;
  assign n5133 = \ctl_rf_c7dmabs_reg[24]/NET0131  & \haddr[4]_pad  ;
  assign n5134 = n4582 & n5133 ;
  assign n5135 = ~n5132 & ~n5134 ;
  assign n5136 = n5130 & n5135 ;
  assign n5137 = n5125 & n5136 ;
  assign n5138 = n4589 & ~n5137 ;
  assign n5139 = ~\haddr[8]_pad  & ~n5138 ;
  assign n5140 = ~n5114 & n5139 ;
  assign n5141 = n4569 & ~n5140 ;
  assign n5142 = ~n5090 & n5141 ;
  assign n5143 = ~n5017 & ~n5142 ;
  assign n5144 = n4573 & ~n5143 ;
  assign n5145 = ~\haddr[8]_pad  & ~n4745 ;
  assign n5146 = ~n4745 & n4859 ;
  assign n5147 = n4833 & n5146 ;
  assign n5148 = ~n5145 & ~n5147 ;
  assign n5149 = n4745 & ~n5010 ;
  assign n5150 = ~n5143 & ~n5149 ;
  assign n5151 = n5148 & n5150 ;
  assign n5152 = ~n5144 & ~n5151 ;
  assign n5153 = ~n5016 & n5152 ;
  assign n5154 = \hrdata_reg[24]_pad  & ~n4569 ;
  assign n5155 = ~\haddr[8]_pad  & n4573 ;
  assign n5156 = n4573 & n4859 ;
  assign n5157 = n4833 & n5156 ;
  assign n5158 = ~n5155 & ~n5157 ;
  assign n5159 = ~n5090 & ~n5140 ;
  assign n5160 = ~n4745 & ~n5159 ;
  assign n5161 = ~n4739 & n4745 ;
  assign n5162 = ~n4713 & n5161 ;
  assign n5163 = ~n5160 & ~n5162 ;
  assign n5164 = ~n4573 & ~n5163 ;
  assign n5165 = n4569 & ~n5164 ;
  assign n5166 = n5158 & n5165 ;
  assign n5167 = ~n5154 & ~n5166 ;
  assign n5168 = \de_de_st_reg[5]/NET0131  & n3047 ;
  assign n5169 = n2983 & n5168 ;
  assign n5170 = n3050 & n5169 ;
  assign n5171 = n2814 & n5170 ;
  assign n5172 = ~n4053 & n5171 ;
  assign n5173 = ~\de_de_st_reg[0]/NET0131  & ~\de_de_st_reg[5]/NET0131  ;
  assign n5174 = n2983 & n5173 ;
  assign n5175 = n3050 & n5174 ;
  assign n5176 = \ctl_rf_c0_rf_chabt_reg/NET0131  & ~n5175 ;
  assign n5177 = \ctl_rf_c0_rf_chllpen_reg/NET0131  & ~n5170 ;
  assign n5178 = ~n5176 & n5177 ;
  assign n5179 = ~n5172 & ~n5178 ;
  assign n5180 = \de_de_st_reg[5]/NET0131  & n3071 ;
  assign n5181 = ~n2983 & n5180 ;
  assign n5182 = n3050 & n5181 ;
  assign n5183 = n2814 & n5182 ;
  assign n5184 = ~n4053 & n5183 ;
  assign n5185 = ~n2983 & n5173 ;
  assign n5186 = n3050 & n5185 ;
  assign n5187 = \ctl_rf_c1_rf_chabt_reg/NET0131  & ~n5186 ;
  assign n5188 = \ctl_rf_c1_rf_chllpen_reg/NET0131  & ~n5182 ;
  assign n5189 = ~n5187 & n5188 ;
  assign n5190 = ~n5184 & ~n5189 ;
  assign n5191 = \de_de_st_reg[5]/NET0131  & n3059 ;
  assign n5192 = n2983 & n5191 ;
  assign n5193 = n3024 & n5192 ;
  assign n5194 = n2814 & n5193 ;
  assign n5195 = ~n4053 & n5194 ;
  assign n5196 = n3024 & n5174 ;
  assign n5197 = \ctl_rf_c2_rf_chabt_reg/NET0131  & ~n5196 ;
  assign n5198 = \ctl_rf_c2_rf_chllpen_reg/NET0131  & ~n5193 ;
  assign n5199 = ~n5197 & n5198 ;
  assign n5200 = ~n5195 & ~n5199 ;
  assign n5201 = \de_de_st_reg[5]/NET0131  & n3021 ;
  assign n5202 = ~n2983 & n5201 ;
  assign n5203 = n3024 & n5202 ;
  assign n5204 = n2814 & n5203 ;
  assign n5205 = ~n4053 & n5204 ;
  assign n5206 = n3024 & n5185 ;
  assign n5207 = \ctl_rf_c3_rf_chabt_reg/NET0131  & ~n5206 ;
  assign n5208 = \ctl_rf_c3_rf_chllpen_reg/NET0131  & ~n5203 ;
  assign n5209 = ~n5207 & n5208 ;
  assign n5210 = ~n5205 & ~n5209 ;
  assign n5211 = \de_de_st_reg[5]/NET0131  & n2970 ;
  assign n5212 = n2983 & n5211 ;
  assign n5213 = n2999 & n5212 ;
  assign n5214 = n2814 & n5213 ;
  assign n5215 = ~n4053 & n5214 ;
  assign n5216 = n2999 & n5174 ;
  assign n5217 = \ctl_rf_c4_rf_chabt_reg/NET0131  & ~n5216 ;
  assign n5218 = \ctl_rf_c4_rf_chllpen_reg/NET0131  & ~n5213 ;
  assign n5219 = ~n5217 & n5218 ;
  assign n5220 = ~n5215 & ~n5219 ;
  assign n5221 = \de_de_st_reg[5]/NET0131  & n3034 ;
  assign n5222 = ~n2983 & n5221 ;
  assign n5223 = n2999 & n5222 ;
  assign n5224 = n2814 & n5223 ;
  assign n5225 = ~n4053 & n5224 ;
  assign n5226 = n2999 & n5185 ;
  assign n5227 = \ctl_rf_c5_rf_chabt_reg/NET0131  & ~n5226 ;
  assign n5228 = \ctl_rf_c5_rf_chllpen_reg/NET0131  & ~n5223 ;
  assign n5229 = ~n5227 & n5228 ;
  assign n5230 = ~n5225 & ~n5229 ;
  assign n5231 = \de_de_st_reg[5]/NET0131  & n3008 ;
  assign n5232 = n2983 & n5231 ;
  assign n5233 = n3011 & n5232 ;
  assign n5234 = n2814 & n5233 ;
  assign n5235 = ~n4053 & n5234 ;
  assign n5236 = n3011 & n5174 ;
  assign n5237 = \ctl_rf_c6_rf_chabt_reg/NET0131  & ~n5236 ;
  assign n5238 = \ctl_rf_c6_rf_chllpen_reg/NET0131  & ~n5233 ;
  assign n5239 = ~n5237 & n5238 ;
  assign n5240 = ~n5235 & ~n5239 ;
  assign n5241 = \de_de_st_reg[5]/NET0131  & n3082 ;
  assign n5242 = ~n2983 & n5241 ;
  assign n5243 = n3011 & n5242 ;
  assign n5244 = n2814 & n5243 ;
  assign n5245 = ~n4053 & n5244 ;
  assign n5246 = n3011 & n5185 ;
  assign n5247 = \ctl_rf_c7_rf_chabt_reg/NET0131  & ~n5246 ;
  assign n5248 = \ctl_rf_c7_rf_chllpen_reg/NET0131  & ~n5243 ;
  assign n5249 = ~n5247 & n5248 ;
  assign n5250 = ~n5245 & ~n5249 ;
  assign n5251 = ~n4326 & n4529 ;
  assign n5252 = ~\de_de_st_reg[2]/NET0131  & ~\de_de_st_reg[5]/NET0131  ;
  assign n5253 = \de_de_st_reg[6]/NET0131  & n5252 ;
  assign n5254 = n4547 & n5253 ;
  assign n5255 = ~n5251 & ~n5254 ;
  assign n5256 = \de_de_st_reg[1]/NET0131  & \de_de_st_reg[2]/NET0131  ;
  assign n5257 = ~\de_de_st_reg[0]/NET0131  & ~n5256 ;
  assign n5258 = ~n2815 & n4472 ;
  assign n5259 = n5257 & n5258 ;
  assign n5260 = ~n5254 & ~n5259 ;
  assign n5261 = ~n4475 & ~n5260 ;
  assign n5262 = ~n4529 & ~n5261 ;
  assign n5263 = \ch_sel_arb_req_reg/NET0131  & ~\de_de_st_reg[5]/NET0131  ;
  assign n5264 = ~n3105 & n5263 ;
  assign n5265 = ~\ch_sel_arb_req_reg/NET0131  & ~\ch_sel_de_stup_d1_reg/NET0131  ;
  assign n5266 = ~n3105 & n5265 ;
  assign n5267 = ~n3095 & n5266 ;
  assign n5268 = ~n5264 & ~n5267 ;
  assign n5269 = \hrdata_reg[0]_pad  & ~n4569 ;
  assign n5270 = n4569 & ~n5009 ;
  assign n5271 = ~n4951 & n5270 ;
  assign n5272 = ~n5017 & ~n5271 ;
  assign n5273 = ~n5269 & n5272 ;
  assign n5274 = n4745 & ~n5159 ;
  assign n5275 = ~n4739 & ~n4745 ;
  assign n5276 = ~n4713 & n5275 ;
  assign n5277 = ~n5274 & ~n5276 ;
  assign n5278 = ~n4573 & ~n5269 ;
  assign n5279 = ~n5277 & n5278 ;
  assign n5280 = ~n5273 & ~n5279 ;
  assign n5281 = \hrdata_reg[1]_pad  & ~n4569 ;
  assign n5282 = \ctl_rf_c0_rf_src_sz_reg[1]/NET0131  & n4577 ;
  assign n5283 = \ctl_rf_c0_rf_chllp_cnt_reg[1]/NET0131  & n4579 ;
  assign n5284 = ~n5282 & ~n5283 ;
  assign n5285 = \ctl_rf_c0_rf_chdad_reg[17]/NET0131  & n4582 ;
  assign n5286 = \ctl_rf_c0_rf_chsad_reg[17]/NET0131  & n4584 ;
  assign n5287 = ~n5285 & ~n5286 ;
  assign n5288 = n5284 & n5287 ;
  assign n5289 = n4623 & ~n5288 ;
  assign n5290 = \haddr[8]_pad  & ~n5289 ;
  assign n5291 = \ctl_rf_c2_rf_chllp_cnt_reg[1]/NET0131  & n4579 ;
  assign n5292 = \ctl_rf_c2_rf_chdad_reg[17]/NET0131  & n4582 ;
  assign n5293 = ~n5291 & ~n5292 ;
  assign n5294 = \ctl_rf_c2_rf_chsad_reg[17]/NET0131  & n4584 ;
  assign n5295 = \ctl_rf_c2_rf_src_sz_reg[1]/NET0131  & n4577 ;
  assign n5296 = ~n5294 & ~n5295 ;
  assign n5297 = n5293 & n5296 ;
  assign n5298 = n4590 & ~n5297 ;
  assign n5299 = \ctl_rf_c4_rf_chllp_cnt_reg[1]/NET0131  & n4579 ;
  assign n5300 = \ctl_rf_c4_rf_chdad_reg[17]/NET0131  & n4582 ;
  assign n5301 = ~n5299 & ~n5300 ;
  assign n5302 = \ctl_rf_c4_rf_chsad_reg[17]/NET0131  & n4584 ;
  assign n5303 = \ctl_rf_c4_rf_src_sz_reg[1]/NET0131  & n4577 ;
  assign n5304 = ~n5302 & ~n5303 ;
  assign n5305 = n5301 & n5304 ;
  assign n5306 = n4576 & ~n5305 ;
  assign n5307 = ~n5298 & ~n5306 ;
  assign n5308 = \ctl_rf_c7_rf_chllp_cnt_reg[1]/NET0131  & n4579 ;
  assign n5309 = \ctl_rf_c7_rf_chdad_reg[17]/NET0131  & n4582 ;
  assign n5310 = ~n5308 & ~n5309 ;
  assign n5311 = \ctl_rf_c7_rf_chsad_reg[17]/NET0131  & n4584 ;
  assign n5312 = \ctl_rf_c7_rf_src_sz_reg[1]/NET0131  & n4577 ;
  assign n5313 = ~n5311 & ~n5312 ;
  assign n5314 = n5310 & n5313 ;
  assign n5315 = n4642 & ~n5314 ;
  assign n5316 = \ctl_rf_c1_rf_src_sz_reg[1]/NET0131  & n4577 ;
  assign n5317 = \ctl_rf_c1_rf_chllp_cnt_reg[1]/NET0131  & n4579 ;
  assign n5318 = ~n5316 & ~n5317 ;
  assign n5319 = \ctl_rf_c1_rf_chdad_reg[17]/NET0131  & n4582 ;
  assign n5320 = \ctl_rf_c1_rf_chsad_reg[17]/NET0131  & n4584 ;
  assign n5321 = ~n5319 & ~n5320 ;
  assign n5322 = n5318 & n5321 ;
  assign n5323 = n4632 & ~n5322 ;
  assign n5324 = ~n5315 & ~n5323 ;
  assign n5325 = n5307 & n5324 ;
  assign n5326 = n5290 & n5325 ;
  assign n5327 = \ctl_rf_c5_rf_chllp_reg[17]/NET0131  & n4680 ;
  assign n5328 = \ctl_rf_c3_rf_chllp_reg[17]/NET0131  & n4698 ;
  assign n5329 = ~n5327 & ~n5328 ;
  assign n5330 = \ctl_rf_c0_rf_chllp_reg[17]/NET0131  & n4675 ;
  assign n5331 = \ctl_rf_c4_rf_chllp_reg[17]/NET0131  & n4687 ;
  assign n5332 = ~n5330 & ~n5331 ;
  assign n5333 = n5329 & n5332 ;
  assign n5334 = \ctl_rf_c6_rf_chllp_reg[17]/NET0131  & n4703 ;
  assign n5335 = \ctl_rf_c2_rf_chllp_reg[17]/NET0131  & n4663 ;
  assign n5336 = ~n5334 & ~n5335 ;
  assign n5337 = \ctl_rf_c1_rf_chllp_reg[17]/NET0131  & n4692 ;
  assign n5338 = \ctl_rf_c7_rf_chllp_reg[17]/NET0131  & n4669 ;
  assign n5339 = ~n5337 & ~n5338 ;
  assign n5340 = n5336 & n5339 ;
  assign n5341 = n5333 & n5340 ;
  assign n5342 = n4577 & ~n5341 ;
  assign n5343 = \ctl_rf_c6_rf_chdad_reg[17]/NET0131  & n4582 ;
  assign n5344 = \ctl_rf_c6_rf_src_sz_reg[1]/NET0131  & n4577 ;
  assign n5345 = ~n5343 & ~n5344 ;
  assign n5346 = \ctl_rf_c6_rf_chllp_cnt_reg[1]/NET0131  & n4579 ;
  assign n5347 = \ctl_rf_c6_rf_chsad_reg[17]/NET0131  & n4584 ;
  assign n5348 = ~n5346 & ~n5347 ;
  assign n5349 = n5345 & n5348 ;
  assign n5350 = n4611 & ~n5349 ;
  assign n5351 = \ctl_rf_c5_rf_chllp_cnt_reg[1]/NET0131  & n4579 ;
  assign n5352 = \ctl_rf_c5_rf_chdad_reg[17]/NET0131  & n4582 ;
  assign n5353 = ~n5351 & ~n5352 ;
  assign n5354 = \ctl_rf_c5_rf_chsad_reg[17]/NET0131  & n4584 ;
  assign n5355 = \ctl_rf_c5_rf_src_sz_reg[1]/NET0131  & n4577 ;
  assign n5356 = ~n5354 & ~n5355 ;
  assign n5357 = n5353 & n5356 ;
  assign n5358 = n4601 & ~n5357 ;
  assign n5359 = \ctl_rf_c3_rf_chllp_cnt_reg[1]/NET0131  & n4579 ;
  assign n5360 = \ctl_rf_c3_rf_chsad_reg[17]/NET0131  & n4584 ;
  assign n5361 = ~n5359 & ~n5360 ;
  assign n5362 = \ctl_rf_c3_rf_src_sz_reg[1]/NET0131  & n4577 ;
  assign n5363 = \ctl_rf_c3_rf_chdad_reg[17]/NET0131  & n4582 ;
  assign n5364 = ~n5362 & ~n5363 ;
  assign n5365 = n5361 & n5364 ;
  assign n5366 = n4651 & ~n5365 ;
  assign n5367 = ~n5358 & ~n5366 ;
  assign n5368 = ~n5350 & n5367 ;
  assign n5369 = ~n5342 & n5368 ;
  assign n5370 = n5326 & n5369 ;
  assign n5371 = \ctl_rf_c1brbs_reg[17]/NET0131  & ~\haddr[4]_pad  ;
  assign n5372 = n4579 & n5371 ;
  assign n5373 = \ctl_rf_c3brbs_reg[17]/NET0131  & ~\haddr[4]_pad  ;
  assign n5374 = n4582 & n5373 ;
  assign n5375 = ~n5372 & ~n5374 ;
  assign n5376 = \ctl_rf_c0brbs_reg[17]/NET0131  & ~\haddr[4]_pad  ;
  assign n5377 = n4577 & n5376 ;
  assign n5378 = \ctl_rf_c7brbs_reg[17]/NET0131  & \haddr[4]_pad  ;
  assign n5379 = n4582 & n5378 ;
  assign n5380 = ~n5377 & ~n5379 ;
  assign n5381 = n5375 & n5380 ;
  assign n5382 = \ctl_rf_c6brbs_reg[17]/NET0131  & \haddr[4]_pad  ;
  assign n5383 = n4584 & n5382 ;
  assign n5384 = \ctl_rf_c4brbs_reg[17]/NET0131  & \haddr[4]_pad  ;
  assign n5385 = n4577 & n5384 ;
  assign n5386 = ~n5383 & ~n5385 ;
  assign n5387 = \ctl_rf_c2brbs_reg[17]/NET0131  & ~\haddr[4]_pad  ;
  assign n5388 = n4584 & n5387 ;
  assign n5389 = \ctl_rf_c5brbs_reg[17]/NET0131  & \haddr[4]_pad  ;
  assign n5390 = n4579 & n5389 ;
  assign n5391 = ~n5388 & ~n5390 ;
  assign n5392 = n5386 & n5391 ;
  assign n5393 = n5381 & n5392 ;
  assign n5394 = n4575 & ~n5393 ;
  assign n5395 = \ctl_rf_c2dmabs_reg[17]/NET0131  & ~\haddr[4]_pad  ;
  assign n5396 = n4584 & n5395 ;
  assign n5397 = \ctl_rf_c3dmabs_reg[17]/NET0131  & ~\haddr[4]_pad  ;
  assign n5398 = n4582 & n5397 ;
  assign n5399 = ~n5396 & ~n5398 ;
  assign n5400 = \ctl_rf_c0dmabs_reg[17]/NET0131  & ~\haddr[4]_pad  ;
  assign n5401 = n4577 & n5400 ;
  assign n5402 = \ctl_rf_c6dmabs_reg[17]/NET0131  & \haddr[4]_pad  ;
  assign n5403 = n4584 & n5402 ;
  assign n5404 = ~n5401 & ~n5403 ;
  assign n5405 = n5399 & n5404 ;
  assign n5406 = \ctl_rf_c7dmabs_reg[17]/NET0131  & \haddr[4]_pad  ;
  assign n5407 = n4582 & n5406 ;
  assign n5408 = \ctl_rf_c4dmabs_reg[17]/NET0131  & \haddr[4]_pad  ;
  assign n5409 = n4577 & n5408 ;
  assign n5410 = ~n5407 & ~n5409 ;
  assign n5411 = \ctl_rf_c1dmabs_reg[17]/NET0131  & ~\haddr[4]_pad  ;
  assign n5412 = n4579 & n5411 ;
  assign n5413 = \ctl_rf_c5dmabs_reg[17]/NET0131  & \haddr[4]_pad  ;
  assign n5414 = n4579 & n5413 ;
  assign n5415 = ~n5412 & ~n5414 ;
  assign n5416 = n5410 & n5415 ;
  assign n5417 = n5405 & n5416 ;
  assign n5418 = n4589 & ~n5417 ;
  assign n5419 = \ctl_rf_abt_reg[1]/NET0131  & n4622 ;
  assign n5420 = ~\haddr[8]_pad  & ~n5419 ;
  assign n5421 = ~\ctl_rf_c1_rf_int_abt_msk_reg/NET0131  & n5002 ;
  assign n5422 = n5005 & ~n5421 ;
  assign n5423 = ~n5420 & ~n5422 ;
  assign n5424 = ~n5418 & ~n5423 ;
  assign n5425 = ~n5394 & n5424 ;
  assign n5426 = n4569 & ~n5425 ;
  assign n5427 = ~n5370 & n5426 ;
  assign n5428 = ~n5017 & ~n5427 ;
  assign n5429 = ~n5281 & n5428 ;
  assign n5430 = \ctl_rf_c5dmabs_reg[25]/NET0131  & \haddr[4]_pad  ;
  assign n5431 = n4579 & n5430 ;
  assign n5432 = \ctl_rf_c6dmabs_reg[25]/NET0131  & \haddr[4]_pad  ;
  assign n5433 = n4584 & n5432 ;
  assign n5434 = ~n5431 & ~n5433 ;
  assign n5435 = \ctl_rf_c2dmabs_reg[25]/NET0131  & ~\haddr[4]_pad  ;
  assign n5436 = n4584 & n5435 ;
  assign n5437 = \ctl_rf_c4dmabs_reg[25]/NET0131  & \haddr[4]_pad  ;
  assign n5438 = n4577 & n5437 ;
  assign n5439 = ~n5436 & ~n5438 ;
  assign n5440 = n5434 & n5439 ;
  assign n5441 = \ctl_rf_c3dmabs_reg[25]/NET0131  & ~\haddr[4]_pad  ;
  assign n5442 = n4582 & n5441 ;
  assign n5443 = \ctl_rf_c1dmabs_reg[25]/NET0131  & ~\haddr[4]_pad  ;
  assign n5444 = n4579 & n5443 ;
  assign n5445 = ~n5442 & ~n5444 ;
  assign n5446 = \ctl_rf_c0dmabs_reg[25]/NET0131  & ~\haddr[4]_pad  ;
  assign n5447 = n4577 & n5446 ;
  assign n5448 = \ctl_rf_c7dmabs_reg[25]/NET0131  & \haddr[4]_pad  ;
  assign n5449 = n4582 & n5448 ;
  assign n5450 = ~n5447 & ~n5449 ;
  assign n5451 = n5445 & n5450 ;
  assign n5452 = n5440 & n5451 ;
  assign n5453 = n4589 & ~n5452 ;
  assign n5454 = \ctl_rf_c2brbs_reg[25]/NET0131  & ~\haddr[4]_pad  ;
  assign n5455 = n4584 & n5454 ;
  assign n5456 = \ctl_rf_c6brbs_reg[25]/NET0131  & \haddr[4]_pad  ;
  assign n5457 = n4584 & n5456 ;
  assign n5458 = ~n5455 & ~n5457 ;
  assign n5459 = \ctl_rf_c1brbs_reg[25]/NET0131  & ~\haddr[4]_pad  ;
  assign n5460 = n4579 & n5459 ;
  assign n5461 = \ctl_rf_c3brbs_reg[25]/NET0131  & ~\haddr[4]_pad  ;
  assign n5462 = n4582 & n5461 ;
  assign n5463 = ~n5460 & ~n5462 ;
  assign n5464 = n5458 & n5463 ;
  assign n5465 = \ctl_rf_c4brbs_reg[25]/NET0131  & \haddr[4]_pad  ;
  assign n5466 = n4577 & n5465 ;
  assign n5467 = \ctl_rf_c0brbs_reg[25]/NET0131  & ~\haddr[4]_pad  ;
  assign n5468 = n4577 & n5467 ;
  assign n5469 = ~n5466 & ~n5468 ;
  assign n5470 = \ctl_rf_c5brbs_reg[25]/NET0131  & \haddr[4]_pad  ;
  assign n5471 = n4579 & n5470 ;
  assign n5472 = \ctl_rf_c7brbs_reg[25]/NET0131  & \haddr[4]_pad  ;
  assign n5473 = n4582 & n5472 ;
  assign n5474 = ~n5471 & ~n5473 ;
  assign n5475 = n5469 & n5474 ;
  assign n5476 = n5464 & n5475 ;
  assign n5477 = n4575 & ~n5476 ;
  assign n5478 = ~\haddr[8]_pad  & ~n5477 ;
  assign n5479 = ~n5453 & n5478 ;
  assign n5480 = n4745 & n5479 ;
  assign n5481 = \ctl_rf_c4_rf_chdad_reg[25]/P0002  & n4582 ;
  assign n5482 = \ctl_rf_c4_rf_chsad_reg[25]/P0002  & n4584 ;
  assign n5483 = ~n5481 & ~n5482 ;
  assign n5484 = n4576 & ~n5483 ;
  assign n5485 = \ctl_rf_c1_rf_chdad_reg[25]/P0002  & n4582 ;
  assign n5486 = \ctl_rf_c1_rf_chsad_reg[25]/P0002  & n4584 ;
  assign n5487 = ~n5485 & ~n5486 ;
  assign n5488 = n4632 & ~n5487 ;
  assign n5489 = \ctl_rf_c3_rf_chdad_reg[25]/P0002  & n4582 ;
  assign n5490 = \ctl_rf_c3_rf_chsad_reg[25]/P0002  & n4584 ;
  assign n5491 = ~n5489 & ~n5490 ;
  assign n5492 = n4651 & ~n5491 ;
  assign n5493 = ~n5488 & ~n5492 ;
  assign n5494 = ~n5484 & n5493 ;
  assign n5495 = \ctl_rf_c7_rf_chdad_reg[25]/P0002  & n4582 ;
  assign n5496 = \ctl_rf_c7_rf_chsad_reg[25]/P0002  & n4584 ;
  assign n5497 = ~n5495 & ~n5496 ;
  assign n5498 = n4642 & ~n5497 ;
  assign n5499 = \haddr[8]_pad  & ~n5498 ;
  assign n5500 = \ctl_rf_c6_rf_chdad_reg[25]/P0002  & n4582 ;
  assign n5501 = \ctl_rf_c6_rf_chsad_reg[25]/P0002  & n4584 ;
  assign n5502 = ~n5500 & ~n5501 ;
  assign n5503 = n4611 & ~n5502 ;
  assign n5504 = \ctl_rf_c2_rf_chdad_reg[25]/P0002  & n4582 ;
  assign n5505 = \ctl_rf_c2_rf_chsad_reg[25]/P0002  & n4584 ;
  assign n5506 = ~n5504 & ~n5505 ;
  assign n5507 = n4590 & ~n5506 ;
  assign n5508 = ~n5503 & ~n5507 ;
  assign n5509 = \ctl_rf_c5_rf_chdad_reg[25]/P0002  & n4582 ;
  assign n5510 = \ctl_rf_c5_rf_chsad_reg[25]/P0002  & n4584 ;
  assign n5511 = ~n5509 & ~n5510 ;
  assign n5512 = n4601 & ~n5511 ;
  assign n5513 = \ctl_rf_c0_rf_chdad_reg[25]/P0002  & n4582 ;
  assign n5514 = \ctl_rf_c0_rf_chsad_reg[25]/P0002  & n4584 ;
  assign n5515 = ~n5513 & ~n5514 ;
  assign n5516 = n4623 & ~n5515 ;
  assign n5517 = ~n5512 & ~n5516 ;
  assign n5518 = n5508 & n5517 ;
  assign n5519 = n5499 & n5518 ;
  assign n5520 = n5494 & n5519 ;
  assign n5521 = \ctl_rf_c1_rf_chllp_reg[25]/NET0131  & n4692 ;
  assign n5522 = \ctl_rf_c3_rf_chllp_reg[25]/NET0131  & n4698 ;
  assign n5523 = ~n5521 & ~n5522 ;
  assign n5524 = \ctl_rf_c0_rf_chllp_reg[25]/NET0131  & n4675 ;
  assign n5525 = \ctl_rf_c4_rf_chllp_reg[25]/NET0131  & n4687 ;
  assign n5526 = ~n5524 & ~n5525 ;
  assign n5527 = n5523 & n5526 ;
  assign n5528 = \ctl_rf_c6_rf_chllp_reg[25]/NET0131  & n4703 ;
  assign n5529 = \ctl_rf_c5_rf_chllp_reg[25]/NET0131  & n4680 ;
  assign n5530 = ~n5528 & ~n5529 ;
  assign n5531 = \ctl_rf_c2_rf_chllp_reg[25]/NET0131  & n4663 ;
  assign n5532 = \ctl_rf_c7_rf_chllp_reg[25]/NET0131  & n4669 ;
  assign n5533 = ~n5531 & ~n5532 ;
  assign n5534 = n5530 & n5533 ;
  assign n5535 = n5527 & n5534 ;
  assign n5536 = n4577 & ~n5535 ;
  assign n5537 = n4745 & ~n5536 ;
  assign n5538 = n5520 & n5537 ;
  assign n5539 = ~n5480 & ~n5538 ;
  assign n5540 = \ctl_rf_c7_rf_chsad_reg[1]/NET0131  & n4584 ;
  assign n5541 = \ctl_rf_c7_rf_chdad_reg[1]/NET0131  & n4582 ;
  assign n5542 = ~n5540 & ~n5541 ;
  assign n5543 = \ctl_rf_c7_rf_dst_sel_reg/NET0131  & n4577 ;
  assign n5544 = \ctl_rf_c7_rf_int_err_msk_reg/NET0131  & n4579 ;
  assign n5545 = ~n5543 & ~n5544 ;
  assign n5546 = n5542 & n5545 ;
  assign n5547 = n4642 & ~n5546 ;
  assign n5548 = \ctl_rf_c3_rf_dst_sel_reg/NET0131  & n4577 ;
  assign n5549 = \ctl_rf_c3_rf_chsad_reg[1]/NET0131  & n4584 ;
  assign n5550 = ~n5548 & ~n5549 ;
  assign n5551 = \ctl_rf_c3_rf_chdad_reg[1]/NET0131  & n4582 ;
  assign n5552 = \ctl_rf_c3_rf_int_err_msk_reg/NET0131  & n4579 ;
  assign n5553 = ~n5551 & ~n5552 ;
  assign n5554 = n5550 & n5553 ;
  assign n5555 = n4651 & ~n5554 ;
  assign n5556 = ~n5547 & ~n5555 ;
  assign n5557 = \ctl_rf_c0_rf_chsad_reg[1]/NET0131  & n4584 ;
  assign n5558 = \ctl_rf_c0_rf_dst_sel_reg/NET0131  & n4577 ;
  assign n5559 = ~n5557 & ~n5558 ;
  assign n5560 = \ctl_rf_c0_rf_chdad_reg[1]/NET0131  & n4582 ;
  assign n5561 = \ctl_rf_c0_rf_int_err_msk_reg/NET0131  & n4579 ;
  assign n5562 = ~n5560 & ~n5561 ;
  assign n5563 = n5559 & n5562 ;
  assign n5564 = n4623 & ~n5563 ;
  assign n5565 = \ctl_rf_c1_rf_chsad_reg[1]/NET0131  & n4584 ;
  assign n5566 = \ctl_rf_c1_rf_chdad_reg[1]/NET0131  & n4582 ;
  assign n5567 = ~n5565 & ~n5566 ;
  assign n5568 = \ctl_rf_c1_rf_dst_sel_reg/NET0131  & n4577 ;
  assign n5569 = \ctl_rf_c1_rf_int_err_msk_reg/NET0131  & n4579 ;
  assign n5570 = ~n5568 & ~n5569 ;
  assign n5571 = n5567 & n5570 ;
  assign n5572 = n4632 & ~n5571 ;
  assign n5573 = ~n5564 & ~n5572 ;
  assign n5574 = n5556 & n5573 ;
  assign n5575 = \ctl_rf_c5_rf_chsad_reg[1]/NET0131  & n4584 ;
  assign n5576 = \ctl_rf_c5_rf_chdad_reg[1]/NET0131  & n4582 ;
  assign n5577 = ~n5575 & ~n5576 ;
  assign n5578 = \ctl_rf_c5_rf_dst_sel_reg/NET0131  & n4577 ;
  assign n5579 = \ctl_rf_c5_rf_int_err_msk_reg/NET0131  & n4579 ;
  assign n5580 = ~n5578 & ~n5579 ;
  assign n5581 = n5577 & n5580 ;
  assign n5582 = n4601 & ~n5581 ;
  assign n5583 = \ctl_rf_c6_rf_dst_sel_reg/NET0131  & n4577 ;
  assign n5584 = \ctl_rf_c6_rf_chsad_reg[1]/NET0131  & n4584 ;
  assign n5585 = ~n5583 & ~n5584 ;
  assign n5586 = \ctl_rf_c6_rf_chdad_reg[1]/NET0131  & n4582 ;
  assign n5587 = \ctl_rf_c6_rf_int_err_msk_reg/NET0131  & n4579 ;
  assign n5588 = ~n5586 & ~n5587 ;
  assign n5589 = n5585 & n5588 ;
  assign n5590 = n4611 & ~n5589 ;
  assign n5591 = ~n5582 & ~n5590 ;
  assign n5592 = \ctl_rf_c4_rf_chsad_reg[1]/NET0131  & n4584 ;
  assign n5593 = \ctl_rf_c4_rf_dst_sel_reg/NET0131  & n4577 ;
  assign n5594 = ~n5592 & ~n5593 ;
  assign n5595 = \ctl_rf_c4_rf_chdad_reg[1]/NET0131  & n4582 ;
  assign n5596 = \ctl_rf_c4_rf_int_err_msk_reg/NET0131  & n4579 ;
  assign n5597 = ~n5595 & ~n5596 ;
  assign n5598 = n5594 & n5597 ;
  assign n5599 = n4576 & ~n5598 ;
  assign n5600 = \ctl_rf_c2_rf_chsad_reg[1]/NET0131  & n4584 ;
  assign n5601 = \ctl_rf_c2_rf_chdad_reg[1]/NET0131  & n4582 ;
  assign n5602 = ~n5600 & ~n5601 ;
  assign n5603 = \ctl_rf_c2_rf_dst_sel_reg/NET0131  & n4577 ;
  assign n5604 = \ctl_rf_c2_rf_int_err_msk_reg/NET0131  & n4579 ;
  assign n5605 = ~n5603 & ~n5604 ;
  assign n5606 = n5602 & n5605 ;
  assign n5607 = n4590 & ~n5606 ;
  assign n5608 = ~n5599 & ~n5607 ;
  assign n5609 = n5591 & n5608 ;
  assign n5610 = \ctl_rf_c0_rf_chllp_reg[1]/P0002  & n4577 ;
  assign n5611 = \ctl_rf_c0_rf_chtsz_reg[1]/P0002  & n4579 ;
  assign n5612 = ~n5610 & ~n5611 ;
  assign n5613 = n4675 & ~n5612 ;
  assign n5614 = \ctl_rf_c3_rf_chllp_reg[1]/P0002  & n4577 ;
  assign n5615 = \ctl_rf_c3_rf_chtsz_reg[1]/P0002  & n4579 ;
  assign n5616 = ~n5614 & ~n5615 ;
  assign n5617 = n4698 & ~n5616 ;
  assign n5618 = ~n5613 & ~n5617 ;
  assign n5619 = \ctl_rf_c1_rf_chllp_reg[1]/P0002  & n4577 ;
  assign n5620 = \ctl_rf_c1_rf_chtsz_reg[1]/P0002  & n4579 ;
  assign n5621 = ~n5619 & ~n5620 ;
  assign n5622 = n4692 & ~n5621 ;
  assign n5623 = \ctl_rf_c2_rf_chllp_reg[1]/P0002  & n4577 ;
  assign n5624 = \ctl_rf_c2_rf_chtsz_reg[1]/P0002  & n4579 ;
  assign n5625 = ~n5623 & ~n5624 ;
  assign n5626 = n4663 & ~n5625 ;
  assign n5627 = ~n5622 & ~n5626 ;
  assign n5628 = n5618 & n5627 ;
  assign n5629 = \ctl_rf_c7_rf_chllp_reg[1]/P0002  & n4577 ;
  assign n5630 = \ctl_rf_c7_rf_chtsz_reg[1]/P0002  & n4579 ;
  assign n5631 = ~n5629 & ~n5630 ;
  assign n5632 = n4669 & ~n5631 ;
  assign n5633 = \ctl_rf_c5_rf_chllp_reg[1]/P0002  & n4577 ;
  assign n5634 = \ctl_rf_c5_rf_chtsz_reg[1]/P0002  & n4579 ;
  assign n5635 = ~n5633 & ~n5634 ;
  assign n5636 = n4680 & ~n5635 ;
  assign n5637 = ~n5632 & ~n5636 ;
  assign n5638 = \ctl_rf_c6_rf_chllp_reg[1]/P0002  & n4577 ;
  assign n5639 = \ctl_rf_c6_rf_chtsz_reg[1]/P0002  & n4579 ;
  assign n5640 = ~n5638 & ~n5639 ;
  assign n5641 = n4703 & ~n5640 ;
  assign n5642 = \ctl_rf_c4_rf_chllp_reg[1]/P0002  & n4577 ;
  assign n5643 = \ctl_rf_c4_rf_chtsz_reg[1]/P0002  & n4579 ;
  assign n5644 = ~n5642 & ~n5643 ;
  assign n5645 = n4687 & ~n5644 ;
  assign n5646 = ~n5641 & ~n5645 ;
  assign n5647 = n5637 & n5646 ;
  assign n5648 = n5628 & n5647 ;
  assign n5649 = n5609 & n5648 ;
  assign n5650 = n5574 & n5649 ;
  assign n5651 = \haddr[8]_pad  & ~n5650 ;
  assign n5652 = ~n2983 & n4716 ;
  assign n5653 = n3050 & n5652 ;
  assign n5654 = \ctl_rf_c1_rf_int_tc1_msk_reg/NET0131  & ~\haddr[4]_pad  ;
  assign n5655 = ~\haddr[5]_pad  & n4579 ;
  assign n5656 = ~n5654 & n5655 ;
  assign n5657 = \ctl_rf_tc_reg[1]/NET0131  & n5656 ;
  assign n5658 = \ctl_rf_m0end_reg/NET0131  & n4730 ;
  assign n5659 = \ctl_rf_c1_rf_ch_en_reg/NET0131  & n4727 ;
  assign n5660 = ~n5658 & ~n5659 ;
  assign n5661 = ~\ctl_rf_c1_rf_int_tc1_msk_reg/NET0131  & \ctl_rf_tc_reg[1]/NET0131  ;
  assign n5662 = \ctl_rf_abt_reg[1]/NET0131  & ~\ctl_rf_c1_rf_int_abt_msk_reg/NET0131  ;
  assign n5663 = ~n5661 & ~n5662 ;
  assign n5664 = n4733 & ~n5663 ;
  assign n5665 = \ctl_rf_sync_reg[1]/NET0131  & n4725 ;
  assign n5666 = ~n5664 & ~n5665 ;
  assign n5667 = n5660 & n5666 ;
  assign n5668 = ~n5657 & n5667 ;
  assign n5669 = ~n5653 & n5668 ;
  assign n5670 = n4714 & ~n5669 ;
  assign n5671 = ~n4745 & ~n5670 ;
  assign n5672 = ~n5651 & n5671 ;
  assign n5673 = n5539 & ~n5672 ;
  assign n5674 = ~n4573 & ~n5281 ;
  assign n5675 = ~n5673 & n5674 ;
  assign n5676 = ~n5429 & ~n5675 ;
  assign n5677 = \hrdata_reg[25]_pad  & ~n4569 ;
  assign n5678 = \ctl_rf_c2_rf_chsad_reg[9]/NET0131  & n4584 ;
  assign n5679 = \ctl_rf_c2_rf_dwidth_reg[1]/NET0131  & n4577 ;
  assign n5680 = \ctl_rf_c2_rf_chdad_reg[9]/P0002  & n4582 ;
  assign n5681 = ~n5679 & ~n5680 ;
  assign n5682 = ~n5678 & n5681 ;
  assign n5683 = n4590 & ~n5682 ;
  assign n5684 = \ctl_rf_c0_rf_chsad_reg[9]/NET0131  & n4584 ;
  assign n5685 = \ctl_rf_c0_rf_dwidth_reg[1]/NET0131  & n4577 ;
  assign n5686 = \ctl_rf_c0_rf_chdad_reg[9]/P0002  & n4582 ;
  assign n5687 = ~n5685 & ~n5686 ;
  assign n5688 = ~n5684 & n5687 ;
  assign n5689 = n4623 & ~n5688 ;
  assign n5690 = ~n5683 & ~n5689 ;
  assign n5691 = \ctl_rf_c3_rf_chsad_reg[9]/NET0131  & n4584 ;
  assign n5692 = \ctl_rf_c3_rf_dwidth_reg[1]/NET0131  & n4577 ;
  assign n5693 = \ctl_rf_c3_rf_chdad_reg[9]/P0002  & n4582 ;
  assign n5694 = ~n5692 & ~n5693 ;
  assign n5695 = ~n5691 & n5694 ;
  assign n5696 = n4651 & ~n5695 ;
  assign n5697 = \ctl_rf_c5_rf_chsad_reg[9]/NET0131  & n4584 ;
  assign n5698 = \ctl_rf_c5_rf_dwidth_reg[1]/NET0131  & n4577 ;
  assign n5699 = \ctl_rf_c5_rf_chdad_reg[9]/P0002  & n4582 ;
  assign n5700 = ~n5698 & ~n5699 ;
  assign n5701 = ~n5697 & n5700 ;
  assign n5702 = n4601 & ~n5701 ;
  assign n5703 = ~n5696 & ~n5702 ;
  assign n5704 = n5690 & n5703 ;
  assign n5705 = \ctl_rf_c3_rf_chllp_reg[9]/NET0131  & n4577 ;
  assign n5706 = \ctl_rf_c3_rf_chtsz_reg[9]/P0002  & n4579 ;
  assign n5707 = ~n5705 & ~n5706 ;
  assign n5708 = n4698 & ~n5707 ;
  assign n5709 = \ctl_rf_c2_rf_chllp_reg[9]/NET0131  & n4577 ;
  assign n5710 = \ctl_rf_c2_rf_chtsz_reg[9]/P0002  & n4579 ;
  assign n5711 = ~n5709 & ~n5710 ;
  assign n5712 = n4663 & ~n5711 ;
  assign n5713 = ~n5708 & ~n5712 ;
  assign n5714 = \ctl_rf_c1_rf_chllp_reg[9]/NET0131  & n4577 ;
  assign n5715 = \ctl_rf_c1_rf_chtsz_reg[9]/P0002  & n4579 ;
  assign n5716 = ~n5714 & ~n5715 ;
  assign n5717 = n4692 & ~n5716 ;
  assign n5718 = \ctl_rf_c0_rf_chllp_reg[9]/NET0131  & n4577 ;
  assign n5719 = \ctl_rf_c0_rf_chtsz_reg[9]/P0002  & n4579 ;
  assign n5720 = ~n5718 & ~n5719 ;
  assign n5721 = n4675 & ~n5720 ;
  assign n5722 = ~n5717 & ~n5721 ;
  assign n5723 = n5713 & n5722 ;
  assign n5724 = \ctl_rf_c5_rf_chllp_reg[9]/NET0131  & n4577 ;
  assign n5725 = \ctl_rf_c5_rf_chtsz_reg[9]/P0002  & n4579 ;
  assign n5726 = ~n5724 & ~n5725 ;
  assign n5727 = n4680 & ~n5726 ;
  assign n5728 = \ctl_rf_c4_rf_chllp_reg[9]/NET0131  & n4577 ;
  assign n5729 = \ctl_rf_c4_rf_chtsz_reg[9]/P0002  & n4579 ;
  assign n5730 = ~n5728 & ~n5729 ;
  assign n5731 = n4687 & ~n5730 ;
  assign n5732 = ~n5727 & ~n5731 ;
  assign n5733 = \ctl_rf_c6_rf_chllp_reg[9]/NET0131  & n4577 ;
  assign n5734 = \ctl_rf_c6_rf_chtsz_reg[9]/P0002  & n4579 ;
  assign n5735 = ~n5733 & ~n5734 ;
  assign n5736 = n4703 & ~n5735 ;
  assign n5737 = \ctl_rf_c7_rf_chllp_reg[9]/NET0131  & n4577 ;
  assign n5738 = \ctl_rf_c7_rf_chtsz_reg[9]/P0002  & n4579 ;
  assign n5739 = ~n5737 & ~n5738 ;
  assign n5740 = n4669 & ~n5739 ;
  assign n5741 = ~n5736 & ~n5740 ;
  assign n5742 = n5732 & n5741 ;
  assign n5743 = n5723 & n5742 ;
  assign n5744 = n5704 & n5743 ;
  assign n5745 = \ctl_rf_c1_rf_chsad_reg[9]/NET0131  & n4584 ;
  assign n5746 = \ctl_rf_c1_rf_dwidth_reg[1]/NET0131  & n4577 ;
  assign n5747 = \ctl_rf_c1_rf_chdad_reg[9]/P0002  & n4582 ;
  assign n5748 = ~n5746 & ~n5747 ;
  assign n5749 = ~n5745 & n5748 ;
  assign n5750 = n4632 & ~n5749 ;
  assign n5751 = \ctl_rf_c4_rf_chsad_reg[9]/NET0131  & n4584 ;
  assign n5752 = \ctl_rf_c4_rf_dwidth_reg[1]/NET0131  & n4577 ;
  assign n5753 = \ctl_rf_c4_rf_chdad_reg[9]/P0002  & n4582 ;
  assign n5754 = ~n5752 & ~n5753 ;
  assign n5755 = ~n5751 & n5754 ;
  assign n5756 = n4576 & ~n5755 ;
  assign n5757 = ~n5750 & ~n5756 ;
  assign n5758 = \ctl_rf_c6_rf_chsad_reg[9]/NET0131  & n4584 ;
  assign n5759 = \ctl_rf_c6_rf_dwidth_reg[1]/NET0131  & n4577 ;
  assign n5760 = \ctl_rf_c6_rf_chdad_reg[9]/P0002  & n4582 ;
  assign n5761 = ~n5759 & ~n5760 ;
  assign n5762 = ~n5758 & n5761 ;
  assign n5763 = n4611 & ~n5762 ;
  assign n5764 = \ctl_rf_c7_rf_chsad_reg[9]/NET0131  & n4584 ;
  assign n5765 = \ctl_rf_c7_rf_dwidth_reg[1]/NET0131  & n4577 ;
  assign n5766 = \ctl_rf_c7_rf_chdad_reg[9]/P0002  & n4582 ;
  assign n5767 = ~n5765 & ~n5766 ;
  assign n5768 = ~n5764 & n5767 ;
  assign n5769 = n4642 & ~n5768 ;
  assign n5770 = ~n5763 & ~n5769 ;
  assign n5771 = n5757 & n5770 ;
  assign n5772 = n4573 & n5771 ;
  assign n5773 = n5744 & n5772 ;
  assign n5774 = ~n5155 & ~n5773 ;
  assign n5775 = n4569 & n5774 ;
  assign n5776 = ~n5677 & ~n5775 ;
  assign n5777 = ~n4745 & n5479 ;
  assign n5778 = ~n4745 & ~n5536 ;
  assign n5779 = n5520 & n5778 ;
  assign n5780 = ~n5777 & ~n5779 ;
  assign n5781 = n4745 & ~n5670 ;
  assign n5782 = ~n5651 & n5781 ;
  assign n5783 = n5780 & ~n5782 ;
  assign n5784 = ~n4573 & ~n5677 ;
  assign n5785 = ~n5783 & n5784 ;
  assign n5786 = ~n5776 & ~n5785 ;
  assign n5787 = \hrdata_reg[26]_pad  & ~n4569 ;
  assign n5788 = \ctl_rf_c2_rf_chsad_reg[10]/NET0131  & n4584 ;
  assign n5789 = \ctl_rf_c2_rf_dwidth_reg[2]/NET0131  & n4577 ;
  assign n5790 = \ctl_rf_c2_rf_chdad_reg[10]/P0002  & n4582 ;
  assign n5791 = ~n5789 & ~n5790 ;
  assign n5792 = ~n5788 & n5791 ;
  assign n5793 = n4590 & ~n5792 ;
  assign n5794 = \ctl_rf_c0_rf_chsad_reg[10]/NET0131  & n4584 ;
  assign n5795 = \ctl_rf_c0_rf_dwidth_reg[2]/NET0131  & n4577 ;
  assign n5796 = \ctl_rf_c0_rf_chdad_reg[10]/P0002  & n4582 ;
  assign n5797 = ~n5795 & ~n5796 ;
  assign n5798 = ~n5794 & n5797 ;
  assign n5799 = n4623 & ~n5798 ;
  assign n5800 = ~n5793 & ~n5799 ;
  assign n5801 = \ctl_rf_c5_rf_chsad_reg[10]/NET0131  & n4584 ;
  assign n5802 = \ctl_rf_c5_rf_dwidth_reg[2]/NET0131  & n4577 ;
  assign n5803 = \ctl_rf_c5_rf_chdad_reg[10]/P0002  & n4582 ;
  assign n5804 = ~n5802 & ~n5803 ;
  assign n5805 = ~n5801 & n5804 ;
  assign n5806 = n4601 & ~n5805 ;
  assign n5807 = \ctl_rf_c3_rf_chdad_reg[10]/NET0131  & n4582 ;
  assign n5808 = \ctl_rf_c3_rf_dwidth_reg[2]/NET0131  & n4577 ;
  assign n5809 = \ctl_rf_c3_rf_chsad_reg[10]/P0002  & n4584 ;
  assign n5810 = ~n5808 & ~n5809 ;
  assign n5811 = ~n5807 & n5810 ;
  assign n5812 = n4651 & ~n5811 ;
  assign n5813 = ~n5806 & ~n5812 ;
  assign n5814 = n5800 & n5813 ;
  assign n5815 = \ctl_rf_c3_rf_chllp_reg[10]/NET0131  & n4577 ;
  assign n5816 = \ctl_rf_c3_rf_chtsz_reg[10]/P0002  & n4579 ;
  assign n5817 = ~n5815 & ~n5816 ;
  assign n5818 = n4698 & ~n5817 ;
  assign n5819 = \ctl_rf_c5_rf_chllp_reg[10]/NET0131  & n4577 ;
  assign n5820 = \ctl_rf_c5_rf_chtsz_reg[10]/P0002  & n4579 ;
  assign n5821 = ~n5819 & ~n5820 ;
  assign n5822 = n4680 & ~n5821 ;
  assign n5823 = ~n5818 & ~n5822 ;
  assign n5824 = \ctl_rf_c0_rf_chllp_reg[10]/NET0131  & n4577 ;
  assign n5825 = \ctl_rf_c0_rf_chtsz_reg[10]/P0002  & n4579 ;
  assign n5826 = ~n5824 & ~n5825 ;
  assign n5827 = n4675 & ~n5826 ;
  assign n5828 = \ctl_rf_c1_rf_chllp_reg[10]/NET0131  & n4577 ;
  assign n5829 = \ctl_rf_c1_rf_chtsz_reg[10]/P0002  & n4579 ;
  assign n5830 = ~n5828 & ~n5829 ;
  assign n5831 = n4692 & ~n5830 ;
  assign n5832 = ~n5827 & ~n5831 ;
  assign n5833 = n5823 & n5832 ;
  assign n5834 = \ctl_rf_c2_rf_chllp_reg[10]/NET0131  & n4577 ;
  assign n5835 = \ctl_rf_c2_rf_chtsz_reg[10]/P0002  & n4579 ;
  assign n5836 = ~n5834 & ~n5835 ;
  assign n5837 = n4663 & ~n5836 ;
  assign n5838 = \ctl_rf_c4_rf_chllp_reg[10]/NET0131  & n4577 ;
  assign n5839 = \ctl_rf_c4_rf_chtsz_reg[10]/P0002  & n4579 ;
  assign n5840 = ~n5838 & ~n5839 ;
  assign n5841 = n4687 & ~n5840 ;
  assign n5842 = ~n5837 & ~n5841 ;
  assign n5843 = \ctl_rf_c6_rf_chllp_reg[10]/NET0131  & n4577 ;
  assign n5844 = \ctl_rf_c6_rf_chtsz_reg[10]/P0002  & n4579 ;
  assign n5845 = ~n5843 & ~n5844 ;
  assign n5846 = n4703 & ~n5845 ;
  assign n5847 = \ctl_rf_c7_rf_chllp_reg[10]/NET0131  & n4577 ;
  assign n5848 = \ctl_rf_c7_rf_chtsz_reg[10]/P0002  & n4579 ;
  assign n5849 = ~n5847 & ~n5848 ;
  assign n5850 = n4669 & ~n5849 ;
  assign n5851 = ~n5846 & ~n5850 ;
  assign n5852 = n5842 & n5851 ;
  assign n5853 = n5833 & n5852 ;
  assign n5854 = n5814 & n5853 ;
  assign n5855 = \ctl_rf_c1_rf_chdad_reg[10]/NET0131  & n4582 ;
  assign n5856 = \ctl_rf_c1_rf_dwidth_reg[2]/NET0131  & n4577 ;
  assign n5857 = \ctl_rf_c1_rf_chsad_reg[10]/P0002  & n4584 ;
  assign n5858 = ~n5856 & ~n5857 ;
  assign n5859 = ~n5855 & n5858 ;
  assign n5860 = n4632 & ~n5859 ;
  assign n5861 = \ctl_rf_c4_rf_chsad_reg[10]/NET0131  & n4584 ;
  assign n5862 = \ctl_rf_c4_rf_dwidth_reg[2]/NET0131  & n4577 ;
  assign n5863 = \ctl_rf_c4_rf_chdad_reg[10]/P0002  & n4582 ;
  assign n5864 = ~n5862 & ~n5863 ;
  assign n5865 = ~n5861 & n5864 ;
  assign n5866 = n4576 & ~n5865 ;
  assign n5867 = ~n5860 & ~n5866 ;
  assign n5868 = \ctl_rf_c7_rf_chsad_reg[10]/NET0131  & n4584 ;
  assign n5869 = \ctl_rf_c7_rf_dwidth_reg[2]/NET0131  & n4577 ;
  assign n5870 = \ctl_rf_c7_rf_chdad_reg[10]/P0002  & n4582 ;
  assign n5871 = ~n5869 & ~n5870 ;
  assign n5872 = ~n5868 & n5871 ;
  assign n5873 = n4642 & ~n5872 ;
  assign n5874 = \ctl_rf_c6_rf_chdad_reg[10]/NET0131  & n4582 ;
  assign n5875 = \ctl_rf_c6_rf_dwidth_reg[2]/NET0131  & n4577 ;
  assign n5876 = \ctl_rf_c6_rf_chsad_reg[10]/P0002  & n4584 ;
  assign n5877 = ~n5875 & ~n5876 ;
  assign n5878 = ~n5874 & n5877 ;
  assign n5879 = n4611 & ~n5878 ;
  assign n5880 = ~n5873 & ~n5879 ;
  assign n5881 = n5867 & n5880 ;
  assign n5882 = n4573 & n5881 ;
  assign n5883 = n5854 & n5882 ;
  assign n5884 = ~n5155 & ~n5883 ;
  assign n5885 = n4569 & n5884 ;
  assign n5886 = ~n5787 & ~n5885 ;
  assign n5887 = \ctl_rf_c5brbs_reg[26]/NET0131  & \haddr[4]_pad  ;
  assign n5888 = n4579 & n5887 ;
  assign n5889 = \ctl_rf_c6brbs_reg[26]/NET0131  & \haddr[4]_pad  ;
  assign n5890 = n4584 & n5889 ;
  assign n5891 = ~n5888 & ~n5890 ;
  assign n5892 = \ctl_rf_c1brbs_reg[26]/NET0131  & ~\haddr[4]_pad  ;
  assign n5893 = n4579 & n5892 ;
  assign n5894 = \ctl_rf_c2brbs_reg[26]/NET0131  & ~\haddr[4]_pad  ;
  assign n5895 = n4584 & n5894 ;
  assign n5896 = ~n5893 & ~n5895 ;
  assign n5897 = n5891 & n5896 ;
  assign n5898 = \ctl_rf_c3brbs_reg[26]/NET0131  & ~\haddr[4]_pad  ;
  assign n5899 = n4582 & n5898 ;
  assign n5900 = \ctl_rf_c4brbs_reg[26]/NET0131  & \haddr[4]_pad  ;
  assign n5901 = n4577 & n5900 ;
  assign n5902 = ~n5899 & ~n5901 ;
  assign n5903 = \ctl_rf_c0brbs_reg[26]/NET0131  & ~\haddr[4]_pad  ;
  assign n5904 = n4577 & n5903 ;
  assign n5905 = \ctl_rf_c7brbs_reg[26]/NET0131  & \haddr[4]_pad  ;
  assign n5906 = n4582 & n5905 ;
  assign n5907 = ~n5904 & ~n5906 ;
  assign n5908 = n5902 & n5907 ;
  assign n5909 = n5897 & n5908 ;
  assign n5910 = n4575 & ~n5909 ;
  assign n5911 = \ctl_rf_c1dmabs_reg[26]/NET0131  & ~\haddr[4]_pad  ;
  assign n5912 = n4579 & n5911 ;
  assign n5913 = \ctl_rf_c6dmabs_reg[26]/NET0131  & \haddr[4]_pad  ;
  assign n5914 = n4584 & n5913 ;
  assign n5915 = ~n5912 & ~n5914 ;
  assign n5916 = \ctl_rf_c4dmabs_reg[26]/NET0131  & \haddr[4]_pad  ;
  assign n5917 = n4577 & n5916 ;
  assign n5918 = \ctl_rf_c3dmabs_reg[26]/NET0131  & ~\haddr[4]_pad  ;
  assign n5919 = n4582 & n5918 ;
  assign n5920 = ~n5917 & ~n5919 ;
  assign n5921 = n5915 & n5920 ;
  assign n5922 = \ctl_rf_c2dmabs_reg[26]/NET0131  & ~\haddr[4]_pad  ;
  assign n5923 = n4584 & n5922 ;
  assign n5924 = \ctl_rf_c0dmabs_reg[26]/NET0131  & ~\haddr[4]_pad  ;
  assign n5925 = n4577 & n5924 ;
  assign n5926 = ~n5923 & ~n5925 ;
  assign n5927 = \ctl_rf_c5dmabs_reg[26]/NET0131  & \haddr[4]_pad  ;
  assign n5928 = n4579 & n5927 ;
  assign n5929 = \ctl_rf_c7dmabs_reg[26]/NET0131  & \haddr[4]_pad  ;
  assign n5930 = n4582 & n5929 ;
  assign n5931 = ~n5928 & ~n5930 ;
  assign n5932 = n5926 & n5931 ;
  assign n5933 = n5921 & n5932 ;
  assign n5934 = n4589 & ~n5933 ;
  assign n5935 = ~\haddr[8]_pad  & ~n5934 ;
  assign n5936 = ~n5910 & n5935 ;
  assign n5937 = ~n4745 & n5936 ;
  assign n5938 = \ctl_rf_c3_rf_chdad_reg[26]/P0002  & n4582 ;
  assign n5939 = \ctl_rf_c3_rf_chsad_reg[26]/P0002  & n4584 ;
  assign n5940 = ~n5938 & ~n5939 ;
  assign n5941 = n4651 & ~n5940 ;
  assign n5942 = \ctl_rf_c5_rf_chdad_reg[26]/P0002  & n4582 ;
  assign n5943 = \ctl_rf_c5_rf_chsad_reg[26]/P0002  & n4584 ;
  assign n5944 = ~n5942 & ~n5943 ;
  assign n5945 = n4601 & ~n5944 ;
  assign n5946 = \ctl_rf_c7_rf_chdad_reg[26]/P0002  & n4582 ;
  assign n5947 = \ctl_rf_c7_rf_chsad_reg[26]/P0002  & n4584 ;
  assign n5948 = ~n5946 & ~n5947 ;
  assign n5949 = n4642 & ~n5948 ;
  assign n5950 = ~n5945 & ~n5949 ;
  assign n5951 = ~n5941 & n5950 ;
  assign n5952 = \ctl_rf_c2_rf_chdad_reg[26]/P0002  & n4582 ;
  assign n5953 = \ctl_rf_c2_rf_chsad_reg[26]/P0002  & n4584 ;
  assign n5954 = ~n5952 & ~n5953 ;
  assign n5955 = n4590 & ~n5954 ;
  assign n5956 = \haddr[8]_pad  & ~n5955 ;
  assign n5957 = \ctl_rf_c0_rf_chdad_reg[26]/P0002  & n4582 ;
  assign n5958 = \ctl_rf_c0_rf_chsad_reg[26]/P0002  & n4584 ;
  assign n5959 = ~n5957 & ~n5958 ;
  assign n5960 = n4623 & ~n5959 ;
  assign n5961 = \ctl_rf_c6_rf_chdad_reg[26]/P0002  & n4582 ;
  assign n5962 = \ctl_rf_c6_rf_chsad_reg[26]/P0002  & n4584 ;
  assign n5963 = ~n5961 & ~n5962 ;
  assign n5964 = n4611 & ~n5963 ;
  assign n5965 = ~n5960 & ~n5964 ;
  assign n5966 = \ctl_rf_c1_rf_chdad_reg[26]/P0002  & n4582 ;
  assign n5967 = \ctl_rf_c1_rf_chsad_reg[26]/P0002  & n4584 ;
  assign n5968 = ~n5966 & ~n5967 ;
  assign n5969 = n4632 & ~n5968 ;
  assign n5970 = \ctl_rf_c4_rf_chdad_reg[26]/P0002  & n4582 ;
  assign n5971 = \ctl_rf_c4_rf_chsad_reg[26]/P0002  & n4584 ;
  assign n5972 = ~n5970 & ~n5971 ;
  assign n5973 = n4576 & ~n5972 ;
  assign n5974 = ~n5969 & ~n5973 ;
  assign n5975 = n5965 & n5974 ;
  assign n5976 = n5956 & n5975 ;
  assign n5977 = n5951 & n5976 ;
  assign n5978 = \ctl_rf_c4_rf_chllp_reg[26]/NET0131  & n4687 ;
  assign n5979 = \ctl_rf_c0_rf_chllp_reg[26]/NET0131  & n4675 ;
  assign n5980 = ~n5978 & ~n5979 ;
  assign n5981 = \ctl_rf_c3_rf_chllp_reg[26]/NET0131  & n4698 ;
  assign n5982 = \ctl_rf_c1_rf_chllp_reg[26]/NET0131  & n4692 ;
  assign n5983 = ~n5981 & ~n5982 ;
  assign n5984 = n5980 & n5983 ;
  assign n5985 = \ctl_rf_c5_rf_chllp_reg[26]/NET0131  & n4680 ;
  assign n5986 = \ctl_rf_c6_rf_chllp_reg[26]/NET0131  & n4703 ;
  assign n5987 = ~n5985 & ~n5986 ;
  assign n5988 = \ctl_rf_c7_rf_chllp_reg[26]/NET0131  & n4669 ;
  assign n5989 = \ctl_rf_c2_rf_chllp_reg[26]/NET0131  & n4663 ;
  assign n5990 = ~n5988 & ~n5989 ;
  assign n5991 = n5987 & n5990 ;
  assign n5992 = n5984 & n5991 ;
  assign n5993 = n4577 & ~n5992 ;
  assign n5994 = ~n4745 & ~n5993 ;
  assign n5995 = n5977 & n5994 ;
  assign n5996 = ~n5937 & ~n5995 ;
  assign n5997 = \ctl_rf_c7_rf_int_abt_msk_reg/NET0131  & n4579 ;
  assign n5998 = \ctl_rf_c7_rf_chdad_reg[2]/NET0131  & n4582 ;
  assign n5999 = ~n5997 & ~n5998 ;
  assign n6000 = \ctl_rf_c7_rf_chsad_reg[2]/NET0131  & n4584 ;
  assign n6001 = \ctl_rf_c7_rf_src_sel_reg/NET0131  & n4577 ;
  assign n6002 = ~n6000 & ~n6001 ;
  assign n6003 = n5999 & n6002 ;
  assign n6004 = n4642 & ~n6003 ;
  assign n6005 = \ctl_rf_c2_rf_int_abt_msk_reg/NET0131  & n4579 ;
  assign n6006 = \ctl_rf_c2_rf_chdad_reg[2]/NET0131  & n4582 ;
  assign n6007 = ~n6005 & ~n6006 ;
  assign n6008 = \ctl_rf_c2_rf_src_sel_reg/NET0131  & n4577 ;
  assign n6009 = \ctl_rf_c2_rf_chsad_reg[2]/NET0131  & n4584 ;
  assign n6010 = ~n6008 & ~n6009 ;
  assign n6011 = n6007 & n6010 ;
  assign n6012 = n4590 & ~n6011 ;
  assign n6013 = ~n6004 & ~n6012 ;
  assign n6014 = \ctl_rf_c5_rf_src_sel_reg/NET0131  & n4577 ;
  assign n6015 = \ctl_rf_c5_rf_int_abt_msk_reg/NET0131  & n4579 ;
  assign n6016 = ~n6014 & ~n6015 ;
  assign n6017 = \ctl_rf_c5_rf_chdad_reg[2]/NET0131  & n4582 ;
  assign n6018 = \ctl_rf_c5_rf_chsad_reg[2]/NET0131  & n4584 ;
  assign n6019 = ~n6017 & ~n6018 ;
  assign n6020 = n6016 & n6019 ;
  assign n6021 = n4601 & ~n6020 ;
  assign n6022 = \ctl_rf_c1_rf_int_abt_msk_reg/NET0131  & n4579 ;
  assign n6023 = \ctl_rf_c1_rf_chsad_reg[2]/NET0131  & n4584 ;
  assign n6024 = ~n6022 & ~n6023 ;
  assign n6025 = \ctl_rf_c1_rf_chdad_reg[2]/NET0131  & n4582 ;
  assign n6026 = \ctl_rf_c1_rf_src_sel_reg/NET0131  & n4577 ;
  assign n6027 = ~n6025 & ~n6026 ;
  assign n6028 = n6024 & n6027 ;
  assign n6029 = n4632 & ~n6028 ;
  assign n6030 = ~n6021 & ~n6029 ;
  assign n6031 = n6013 & n6030 ;
  assign n6032 = \ctl_rf_c0_rf_int_abt_msk_reg/NET0131  & n4579 ;
  assign n6033 = \ctl_rf_c0_rf_chdad_reg[2]/NET0131  & n4582 ;
  assign n6034 = ~n6032 & ~n6033 ;
  assign n6035 = \ctl_rf_c0_rf_chsad_reg[2]/NET0131  & n4584 ;
  assign n6036 = \ctl_rf_c0_rf_src_sel_reg/NET0131  & n4577 ;
  assign n6037 = ~n6035 & ~n6036 ;
  assign n6038 = n6034 & n6037 ;
  assign n6039 = n4623 & ~n6038 ;
  assign n6040 = \ctl_rf_c6_rf_int_abt_msk_reg/NET0131  & n4579 ;
  assign n6041 = \ctl_rf_c6_rf_chsad_reg[2]/NET0131  & n4584 ;
  assign n6042 = ~n6040 & ~n6041 ;
  assign n6043 = \ctl_rf_c6_rf_src_sel_reg/NET0131  & n4577 ;
  assign n6044 = \ctl_rf_c6_rf_chdad_reg[2]/NET0131  & n4582 ;
  assign n6045 = ~n6043 & ~n6044 ;
  assign n6046 = n6042 & n6045 ;
  assign n6047 = n4611 & ~n6046 ;
  assign n6048 = ~n6039 & ~n6047 ;
  assign n6049 = \ctl_rf_c4_rf_src_sel_reg/NET0131  & n4577 ;
  assign n6050 = \ctl_rf_c4_rf_int_abt_msk_reg/NET0131  & n4579 ;
  assign n6051 = ~n6049 & ~n6050 ;
  assign n6052 = \ctl_rf_c4_rf_chdad_reg[2]/NET0131  & n4582 ;
  assign n6053 = \ctl_rf_c4_rf_chsad_reg[2]/NET0131  & n4584 ;
  assign n6054 = ~n6052 & ~n6053 ;
  assign n6055 = n6051 & n6054 ;
  assign n6056 = n4576 & ~n6055 ;
  assign n6057 = \ctl_rf_c3_rf_int_abt_msk_reg/NET0131  & n4579 ;
  assign n6058 = \ctl_rf_c3_rf_chdad_reg[2]/NET0131  & n4582 ;
  assign n6059 = ~n6057 & ~n6058 ;
  assign n6060 = \ctl_rf_c3_rf_chsad_reg[2]/NET0131  & n4584 ;
  assign n6061 = \ctl_rf_c3_rf_src_sel_reg/NET0131  & n4577 ;
  assign n6062 = ~n6060 & ~n6061 ;
  assign n6063 = n6059 & n6062 ;
  assign n6064 = n4651 & ~n6063 ;
  assign n6065 = ~n6056 & ~n6064 ;
  assign n6066 = n6048 & n6065 ;
  assign n6067 = \ctl_rf_c0_rf_chllp_reg[2]/NET0131  & n4577 ;
  assign n6068 = \ctl_rf_c0_rf_chtsz_reg[2]/P0002  & n4579 ;
  assign n6069 = ~n6067 & ~n6068 ;
  assign n6070 = n4675 & ~n6069 ;
  assign n6071 = \ctl_rf_c4_rf_chllp_reg[2]/NET0131  & n4577 ;
  assign n6072 = \ctl_rf_c4_rf_chtsz_reg[2]/P0002  & n4579 ;
  assign n6073 = ~n6071 & ~n6072 ;
  assign n6074 = n4687 & ~n6073 ;
  assign n6075 = ~n6070 & ~n6074 ;
  assign n6076 = \ctl_rf_c1_rf_chllp_reg[2]/NET0131  & n4577 ;
  assign n6077 = \ctl_rf_c1_rf_chtsz_reg[2]/P0002  & n4579 ;
  assign n6078 = ~n6076 & ~n6077 ;
  assign n6079 = n4692 & ~n6078 ;
  assign n6080 = \ctl_rf_c2_rf_chllp_reg[2]/NET0131  & n4577 ;
  assign n6081 = \ctl_rf_c2_rf_chtsz_reg[2]/P0002  & n4579 ;
  assign n6082 = ~n6080 & ~n6081 ;
  assign n6083 = n4663 & ~n6082 ;
  assign n6084 = ~n6079 & ~n6083 ;
  assign n6085 = n6075 & n6084 ;
  assign n6086 = \ctl_rf_c7_rf_chllp_reg[2]/NET0131  & n4577 ;
  assign n6087 = \ctl_rf_c7_rf_chtsz_reg[2]/P0002  & n4579 ;
  assign n6088 = ~n6086 & ~n6087 ;
  assign n6089 = n4669 & ~n6088 ;
  assign n6090 = \ctl_rf_c5_rf_chllp_reg[2]/NET0131  & n4577 ;
  assign n6091 = \ctl_rf_c5_rf_chtsz_reg[2]/P0002  & n4579 ;
  assign n6092 = ~n6090 & ~n6091 ;
  assign n6093 = n4680 & ~n6092 ;
  assign n6094 = ~n6089 & ~n6093 ;
  assign n6095 = \ctl_rf_c3_rf_chllp_reg[2]/NET0131  & n4577 ;
  assign n6096 = \ctl_rf_c3_rf_chtsz_reg[2]/P0002  & n4579 ;
  assign n6097 = ~n6095 & ~n6096 ;
  assign n6098 = n4698 & ~n6097 ;
  assign n6099 = \ctl_rf_c6_rf_chllp_reg[2]/NET0131  & n4577 ;
  assign n6100 = \ctl_rf_c6_rf_chtsz_reg[2]/P0002  & n4579 ;
  assign n6101 = ~n6099 & ~n6100 ;
  assign n6102 = n4703 & ~n6101 ;
  assign n6103 = ~n6098 & ~n6102 ;
  assign n6104 = n6094 & n6103 ;
  assign n6105 = n6085 & n6104 ;
  assign n6106 = n6066 & n6105 ;
  assign n6107 = n6031 & n6106 ;
  assign n6108 = \haddr[8]_pad  & ~n6107 ;
  assign n6109 = n3024 & n4717 ;
  assign n6110 = \ctl_rf_c2_rf_int_tc1_msk_reg/NET0131  & ~\haddr[4]_pad  ;
  assign n6111 = n5655 & ~n6110 ;
  assign n6112 = \ctl_rf_tc_reg[2]/NET0131  & n6111 ;
  assign n6113 = \ctl_rf_m1end_reg/NET0131  & n4730 ;
  assign n6114 = \ctl_rf_c2_rf_ch_en_reg/NET0131  & n4727 ;
  assign n6115 = ~n6113 & ~n6114 ;
  assign n6116 = ~\ctl_rf_c2_rf_int_tc1_msk_reg/NET0131  & \ctl_rf_tc_reg[2]/NET0131  ;
  assign n6117 = \ctl_rf_abt_reg[2]/NET0131  & ~\ctl_rf_c2_rf_int_abt_msk_reg/NET0131  ;
  assign n6118 = ~n6116 & ~n6117 ;
  assign n6119 = n4733 & ~n6118 ;
  assign n6120 = \ctl_rf_sync_reg[2]/NET0131  & n4725 ;
  assign n6121 = ~n6119 & ~n6120 ;
  assign n6122 = n6115 & n6121 ;
  assign n6123 = ~n6112 & n6122 ;
  assign n6124 = ~n6109 & n6123 ;
  assign n6125 = n4714 & ~n6124 ;
  assign n6126 = n4745 & ~n6125 ;
  assign n6127 = ~n6108 & n6126 ;
  assign n6128 = n5996 & ~n6127 ;
  assign n6129 = ~n4573 & ~n5787 ;
  assign n6130 = ~n6128 & n6129 ;
  assign n6131 = ~n5886 & ~n6130 ;
  assign n6132 = \hrdata_reg[27]_pad  & ~n4569 ;
  assign n6133 = \ctl_rf_c5_rf_chsad_reg[11]/NET0131  & n4584 ;
  assign n6134 = \ctl_rf_c5_rf_swidth_reg[0]/NET0131  & n4577 ;
  assign n6135 = \ctl_rf_c5_rf_chdad_reg[11]/P0002  & n4582 ;
  assign n6136 = ~n6134 & ~n6135 ;
  assign n6137 = ~n6133 & n6136 ;
  assign n6138 = n4601 & ~n6137 ;
  assign n6139 = \ctl_rf_c0_rf_chdad_reg[11]/NET0131  & n4582 ;
  assign n6140 = \ctl_rf_c0_rf_swidth_reg[0]/NET0131  & n4577 ;
  assign n6141 = \ctl_rf_c0_rf_chsad_reg[11]/P0002  & n4584 ;
  assign n6142 = ~n6140 & ~n6141 ;
  assign n6143 = ~n6139 & n6142 ;
  assign n6144 = n4623 & ~n6143 ;
  assign n6145 = ~n6138 & ~n6144 ;
  assign n6146 = \ctl_rf_c3_rf_chdad_reg[11]/NET0131  & n4582 ;
  assign n6147 = \ctl_rf_c3_rf_swidth_reg[0]/NET0131  & n4577 ;
  assign n6148 = \ctl_rf_c3_rf_chsad_reg[11]/P0002  & n4584 ;
  assign n6149 = ~n6147 & ~n6148 ;
  assign n6150 = ~n6146 & n6149 ;
  assign n6151 = n4651 & ~n6150 ;
  assign n6152 = \ctl_rf_c2_rf_chsad_reg[11]/NET0131  & n4584 ;
  assign n6153 = \ctl_rf_c2_rf_swidth_reg[0]/NET0131  & n4577 ;
  assign n6154 = \ctl_rf_c2_rf_chdad_reg[11]/P0002  & n4582 ;
  assign n6155 = ~n6153 & ~n6154 ;
  assign n6156 = ~n6152 & n6155 ;
  assign n6157 = n4590 & ~n6156 ;
  assign n6158 = ~n6151 & ~n6157 ;
  assign n6159 = n6145 & n6158 ;
  assign n6160 = \ctl_rf_c3_rf_chllp_reg[11]/NET0131  & n4577 ;
  assign n6161 = \ctl_rf_c3_rf_chtsz_reg[11]/P0002  & n4579 ;
  assign n6162 = ~n6160 & ~n6161 ;
  assign n6163 = n4698 & ~n6162 ;
  assign n6164 = \ctl_rf_c2_rf_chllp_reg[11]/NET0131  & n4577 ;
  assign n6165 = \ctl_rf_c2_rf_chtsz_reg[11]/P0002  & n4579 ;
  assign n6166 = ~n6164 & ~n6165 ;
  assign n6167 = n4663 & ~n6166 ;
  assign n6168 = ~n6163 & ~n6167 ;
  assign n6169 = \ctl_rf_c1_rf_chllp_reg[11]/NET0131  & n4577 ;
  assign n6170 = \ctl_rf_c1_rf_chtsz_reg[11]/P0002  & n4579 ;
  assign n6171 = ~n6169 & ~n6170 ;
  assign n6172 = n4692 & ~n6171 ;
  assign n6173 = \ctl_rf_c0_rf_chllp_reg[11]/NET0131  & n4577 ;
  assign n6174 = \ctl_rf_c0_rf_chtsz_reg[11]/P0002  & n4579 ;
  assign n6175 = ~n6173 & ~n6174 ;
  assign n6176 = n4675 & ~n6175 ;
  assign n6177 = ~n6172 & ~n6176 ;
  assign n6178 = n6168 & n6177 ;
  assign n6179 = \ctl_rf_c5_rf_chllp_reg[11]/NET0131  & n4577 ;
  assign n6180 = \ctl_rf_c5_rf_chtsz_reg[11]/P0002  & n4579 ;
  assign n6181 = ~n6179 & ~n6180 ;
  assign n6182 = n4680 & ~n6181 ;
  assign n6183 = \ctl_rf_c4_rf_chllp_reg[11]/NET0131  & n4577 ;
  assign n6184 = \ctl_rf_c4_rf_chtsz_reg[11]/P0002  & n4579 ;
  assign n6185 = ~n6183 & ~n6184 ;
  assign n6186 = n4687 & ~n6185 ;
  assign n6187 = ~n6182 & ~n6186 ;
  assign n6188 = \ctl_rf_c6_rf_chllp_reg[11]/NET0131  & n4577 ;
  assign n6189 = \ctl_rf_c6_rf_chtsz_reg[11]/P0002  & n4579 ;
  assign n6190 = ~n6188 & ~n6189 ;
  assign n6191 = n4703 & ~n6190 ;
  assign n6192 = \ctl_rf_c7_rf_chllp_reg[11]/NET0131  & n4577 ;
  assign n6193 = \ctl_rf_c7_rf_chtsz_reg[11]/P0002  & n4579 ;
  assign n6194 = ~n6192 & ~n6193 ;
  assign n6195 = n4669 & ~n6194 ;
  assign n6196 = ~n6191 & ~n6195 ;
  assign n6197 = n6187 & n6196 ;
  assign n6198 = n6178 & n6197 ;
  assign n6199 = n6159 & n6198 ;
  assign n6200 = \ctl_rf_c1_rf_chsad_reg[11]/NET0131  & n4584 ;
  assign n6201 = \ctl_rf_c1_rf_swidth_reg[0]/NET0131  & n4577 ;
  assign n6202 = \ctl_rf_c1_rf_chdad_reg[11]/P0002  & n4582 ;
  assign n6203 = ~n6201 & ~n6202 ;
  assign n6204 = ~n6200 & n6203 ;
  assign n6205 = n4632 & ~n6204 ;
  assign n6206 = \ctl_rf_c4_rf_chsad_reg[11]/NET0131  & n4584 ;
  assign n6207 = \ctl_rf_c4_rf_swidth_reg[0]/NET0131  & n4577 ;
  assign n6208 = \ctl_rf_c4_rf_chdad_reg[11]/P0002  & n4582 ;
  assign n6209 = ~n6207 & ~n6208 ;
  assign n6210 = ~n6206 & n6209 ;
  assign n6211 = n4576 & ~n6210 ;
  assign n6212 = ~n6205 & ~n6211 ;
  assign n6213 = \ctl_rf_c6_rf_chsad_reg[11]/NET0131  & n4584 ;
  assign n6214 = \ctl_rf_c6_rf_swidth_reg[0]/NET0131  & n4577 ;
  assign n6215 = \ctl_rf_c6_rf_chdad_reg[11]/P0002  & n4582 ;
  assign n6216 = ~n6214 & ~n6215 ;
  assign n6217 = ~n6213 & n6216 ;
  assign n6218 = n4611 & ~n6217 ;
  assign n6219 = \ctl_rf_c7_rf_chdad_reg[11]/NET0131  & n4582 ;
  assign n6220 = \ctl_rf_c7_rf_swidth_reg[0]/NET0131  & n4577 ;
  assign n6221 = \ctl_rf_c7_rf_chsad_reg[11]/P0002  & n4584 ;
  assign n6222 = ~n6220 & ~n6221 ;
  assign n6223 = ~n6219 & n6222 ;
  assign n6224 = n4642 & ~n6223 ;
  assign n6225 = ~n6218 & ~n6224 ;
  assign n6226 = n6212 & n6225 ;
  assign n6227 = n4573 & n6226 ;
  assign n6228 = n6199 & n6227 ;
  assign n6229 = ~n5155 & ~n6228 ;
  assign n6230 = n4569 & n6229 ;
  assign n6231 = ~n6132 & ~n6230 ;
  assign n6232 = \ctl_rf_c5dmabs_reg[27]/NET0131  & \haddr[4]_pad  ;
  assign n6233 = n4579 & n6232 ;
  assign n6234 = \ctl_rf_c6dmabs_reg[27]/NET0131  & \haddr[4]_pad  ;
  assign n6235 = n4584 & n6234 ;
  assign n6236 = ~n6233 & ~n6235 ;
  assign n6237 = \ctl_rf_c1dmabs_reg[27]/NET0131  & ~\haddr[4]_pad  ;
  assign n6238 = n4579 & n6237 ;
  assign n6239 = \ctl_rf_c2dmabs_reg[27]/NET0131  & ~\haddr[4]_pad  ;
  assign n6240 = n4584 & n6239 ;
  assign n6241 = ~n6238 & ~n6240 ;
  assign n6242 = n6236 & n6241 ;
  assign n6243 = \ctl_rf_c3dmabs_reg[27]/NET0131  & ~\haddr[4]_pad  ;
  assign n6244 = n4582 & n6243 ;
  assign n6245 = \ctl_rf_c4dmabs_reg[27]/NET0131  & \haddr[4]_pad  ;
  assign n6246 = n4577 & n6245 ;
  assign n6247 = ~n6244 & ~n6246 ;
  assign n6248 = \ctl_rf_c0dmabs_reg[27]/NET0131  & ~\haddr[4]_pad  ;
  assign n6249 = n4577 & n6248 ;
  assign n6250 = \ctl_rf_c7dmabs_reg[27]/NET0131  & \haddr[4]_pad  ;
  assign n6251 = n4582 & n6250 ;
  assign n6252 = ~n6249 & ~n6251 ;
  assign n6253 = n6247 & n6252 ;
  assign n6254 = n6242 & n6253 ;
  assign n6255 = n4589 & ~n6254 ;
  assign n6256 = \ctl_rf_c1brbs_reg[27]/NET0131  & ~\haddr[4]_pad  ;
  assign n6257 = n4579 & n6256 ;
  assign n6258 = \ctl_rf_c6brbs_reg[27]/NET0131  & \haddr[4]_pad  ;
  assign n6259 = n4584 & n6258 ;
  assign n6260 = ~n6257 & ~n6259 ;
  assign n6261 = \ctl_rf_c4brbs_reg[27]/NET0131  & \haddr[4]_pad  ;
  assign n6262 = n4577 & n6261 ;
  assign n6263 = \ctl_rf_c3brbs_reg[27]/NET0131  & ~\haddr[4]_pad  ;
  assign n6264 = n4582 & n6263 ;
  assign n6265 = ~n6262 & ~n6264 ;
  assign n6266 = n6260 & n6265 ;
  assign n6267 = \ctl_rf_c2brbs_reg[27]/NET0131  & ~\haddr[4]_pad  ;
  assign n6268 = n4584 & n6267 ;
  assign n6269 = \ctl_rf_c0brbs_reg[27]/NET0131  & ~\haddr[4]_pad  ;
  assign n6270 = n4577 & n6269 ;
  assign n6271 = ~n6268 & ~n6270 ;
  assign n6272 = \ctl_rf_c5brbs_reg[27]/NET0131  & \haddr[4]_pad  ;
  assign n6273 = n4579 & n6272 ;
  assign n6274 = \ctl_rf_c7brbs_reg[27]/NET0131  & \haddr[4]_pad  ;
  assign n6275 = n4582 & n6274 ;
  assign n6276 = ~n6273 & ~n6275 ;
  assign n6277 = n6271 & n6276 ;
  assign n6278 = n6266 & n6277 ;
  assign n6279 = n4575 & ~n6278 ;
  assign n6280 = ~\haddr[8]_pad  & ~n6279 ;
  assign n6281 = ~n6255 & n6280 ;
  assign n6282 = ~n4745 & n6281 ;
  assign n6283 = \ctl_rf_c3_rf_chdad_reg[27]/P0002  & n4582 ;
  assign n6284 = \ctl_rf_c3_rf_chsad_reg[27]/P0002  & n4584 ;
  assign n6285 = ~n6283 & ~n6284 ;
  assign n6286 = n4651 & ~n6285 ;
  assign n6287 = \ctl_rf_c5_rf_chdad_reg[27]/P0002  & n4582 ;
  assign n6288 = \ctl_rf_c5_rf_chsad_reg[27]/P0002  & n4584 ;
  assign n6289 = ~n6287 & ~n6288 ;
  assign n6290 = n4601 & ~n6289 ;
  assign n6291 = \ctl_rf_c6_rf_chdad_reg[27]/P0002  & n4582 ;
  assign n6292 = \ctl_rf_c6_rf_chsad_reg[27]/P0002  & n4584 ;
  assign n6293 = ~n6291 & ~n6292 ;
  assign n6294 = n4611 & ~n6293 ;
  assign n6295 = ~n6290 & ~n6294 ;
  assign n6296 = ~n6286 & n6295 ;
  assign n6297 = \ctl_rf_c2_rf_chdad_reg[27]/P0002  & n4582 ;
  assign n6298 = \ctl_rf_c2_rf_chsad_reg[27]/P0002  & n4584 ;
  assign n6299 = ~n6297 & ~n6298 ;
  assign n6300 = n4590 & ~n6299 ;
  assign n6301 = \haddr[8]_pad  & ~n6300 ;
  assign n6302 = \ctl_rf_c0_rf_chdad_reg[27]/P0002  & n4582 ;
  assign n6303 = \ctl_rf_c0_rf_chsad_reg[27]/P0002  & n4584 ;
  assign n6304 = ~n6302 & ~n6303 ;
  assign n6305 = n4623 & ~n6304 ;
  assign n6306 = \ctl_rf_c1_rf_chdad_reg[27]/P0002  & n4582 ;
  assign n6307 = \ctl_rf_c1_rf_chsad_reg[27]/P0002  & n4584 ;
  assign n6308 = ~n6306 & ~n6307 ;
  assign n6309 = n4632 & ~n6308 ;
  assign n6310 = ~n6305 & ~n6309 ;
  assign n6311 = \ctl_rf_c4_rf_chdad_reg[27]/P0002  & n4582 ;
  assign n6312 = \ctl_rf_c4_rf_chsad_reg[27]/P0002  & n4584 ;
  assign n6313 = ~n6311 & ~n6312 ;
  assign n6314 = n4576 & ~n6313 ;
  assign n6315 = \ctl_rf_c7_rf_chdad_reg[27]/P0002  & n4582 ;
  assign n6316 = \ctl_rf_c7_rf_chsad_reg[27]/P0002  & n4584 ;
  assign n6317 = ~n6315 & ~n6316 ;
  assign n6318 = n4642 & ~n6317 ;
  assign n6319 = ~n6314 & ~n6318 ;
  assign n6320 = n6310 & n6319 ;
  assign n6321 = n6301 & n6320 ;
  assign n6322 = n6296 & n6321 ;
  assign n6323 = \ctl_rf_c4_rf_chllp_reg[27]/NET0131  & n4687 ;
  assign n6324 = \ctl_rf_c0_rf_chllp_reg[27]/NET0131  & n4675 ;
  assign n6325 = ~n6323 & ~n6324 ;
  assign n6326 = \ctl_rf_c3_rf_chllp_reg[27]/NET0131  & n4698 ;
  assign n6327 = \ctl_rf_c1_rf_chllp_reg[27]/NET0131  & n4692 ;
  assign n6328 = ~n6326 & ~n6327 ;
  assign n6329 = n6325 & n6328 ;
  assign n6330 = \ctl_rf_c5_rf_chllp_reg[27]/NET0131  & n4680 ;
  assign n6331 = \ctl_rf_c6_rf_chllp_reg[27]/NET0131  & n4703 ;
  assign n6332 = ~n6330 & ~n6331 ;
  assign n6333 = \ctl_rf_c7_rf_chllp_reg[27]/NET0131  & n4669 ;
  assign n6334 = \ctl_rf_c2_rf_chllp_reg[27]/NET0131  & n4663 ;
  assign n6335 = ~n6333 & ~n6334 ;
  assign n6336 = n6332 & n6335 ;
  assign n6337 = n6329 & n6336 ;
  assign n6338 = n4577 & ~n6337 ;
  assign n6339 = ~n4745 & ~n6338 ;
  assign n6340 = n6322 & n6339 ;
  assign n6341 = ~n6282 & ~n6340 ;
  assign n6342 = \ctl_rf_c5_rf_chsad_reg[3]/NET0131  & n4584 ;
  assign n6343 = \ctl_rf_c5_rf_dad_ctl0_reg/NET0131  & n4577 ;
  assign n6344 = \ctl_rf_c5_rf_chdad_reg[3]/P0002  & n4582 ;
  assign n6345 = ~n6343 & ~n6344 ;
  assign n6346 = ~n6342 & n6345 ;
  assign n6347 = n4601 & ~n6346 ;
  assign n6348 = \ctl_rf_c3_rf_chsad_reg[3]/NET0131  & n4584 ;
  assign n6349 = \ctl_rf_c3_rf_dad_ctl0_reg/NET0131  & n4577 ;
  assign n6350 = \ctl_rf_c3_rf_chdad_reg[3]/P0002  & n4582 ;
  assign n6351 = ~n6349 & ~n6350 ;
  assign n6352 = ~n6348 & n6351 ;
  assign n6353 = n4651 & ~n6352 ;
  assign n6354 = ~n6347 & ~n6353 ;
  assign n6355 = \ctl_rf_c0_rf_chsad_reg[3]/NET0131  & n4584 ;
  assign n6356 = \ctl_rf_c0_rf_dad_ctl0_reg/NET0131  & n4577 ;
  assign n6357 = \ctl_rf_c0_rf_chdad_reg[3]/P0002  & n4582 ;
  assign n6358 = ~n6356 & ~n6357 ;
  assign n6359 = ~n6355 & n6358 ;
  assign n6360 = n4623 & ~n6359 ;
  assign n6361 = \ctl_rf_c2_rf_chsad_reg[3]/NET0131  & n4584 ;
  assign n6362 = \ctl_rf_c2_rf_dad_ctl0_reg/NET0131  & n4577 ;
  assign n6363 = \ctl_rf_c2_rf_chdad_reg[3]/P0002  & n4582 ;
  assign n6364 = ~n6362 & ~n6363 ;
  assign n6365 = ~n6361 & n6364 ;
  assign n6366 = n4590 & ~n6365 ;
  assign n6367 = ~n6360 & ~n6366 ;
  assign n6368 = n6354 & n6367 ;
  assign n6369 = \ctl_rf_c7_rf_chsad_reg[3]/NET0131  & n4584 ;
  assign n6370 = \ctl_rf_c7_rf_dad_ctl0_reg/NET0131  & n4577 ;
  assign n6371 = \ctl_rf_c7_rf_chdad_reg[3]/P0002  & n4582 ;
  assign n6372 = ~n6370 & ~n6371 ;
  assign n6373 = ~n6369 & n6372 ;
  assign n6374 = n4642 & ~n6373 ;
  assign n6375 = \ctl_rf_c6_rf_chsad_reg[3]/NET0131  & n4584 ;
  assign n6376 = \ctl_rf_c6_rf_dad_ctl0_reg/NET0131  & n4577 ;
  assign n6377 = \ctl_rf_c6_rf_chdad_reg[3]/P0002  & n4582 ;
  assign n6378 = ~n6376 & ~n6377 ;
  assign n6379 = ~n6375 & n6378 ;
  assign n6380 = n4611 & ~n6379 ;
  assign n6381 = ~n6374 & ~n6380 ;
  assign n6382 = \ctl_rf_c1_rf_chsad_reg[3]/NET0131  & n4584 ;
  assign n6383 = \ctl_rf_c1_rf_dad_ctl0_reg/NET0131  & n4577 ;
  assign n6384 = \ctl_rf_c1_rf_chdad_reg[3]/P0002  & n4582 ;
  assign n6385 = ~n6383 & ~n6384 ;
  assign n6386 = ~n6382 & n6385 ;
  assign n6387 = n4632 & ~n6386 ;
  assign n6388 = \ctl_rf_c4_rf_chsad_reg[3]/NET0131  & n4584 ;
  assign n6389 = \ctl_rf_c4_rf_dad_ctl0_reg/NET0131  & n4577 ;
  assign n6390 = \ctl_rf_c4_rf_chdad_reg[3]/P0002  & n4582 ;
  assign n6391 = ~n6389 & ~n6390 ;
  assign n6392 = ~n6388 & n6391 ;
  assign n6393 = n4576 & ~n6392 ;
  assign n6394 = ~n6387 & ~n6393 ;
  assign n6395 = n6381 & n6394 ;
  assign n6396 = \ctl_rf_c2_rf_chllp_reg[3]/NET0131  & n4577 ;
  assign n6397 = \ctl_rf_c2_rf_chtsz_reg[3]/P0002  & n4579 ;
  assign n6398 = ~n6396 & ~n6397 ;
  assign n6399 = n4663 & ~n6398 ;
  assign n6400 = \ctl_rf_c7_rf_chllp_reg[3]/NET0131  & n4577 ;
  assign n6401 = \ctl_rf_c7_rf_chtsz_reg[3]/P0002  & n4579 ;
  assign n6402 = ~n6400 & ~n6401 ;
  assign n6403 = n4669 & ~n6402 ;
  assign n6404 = ~n6399 & ~n6403 ;
  assign n6405 = \ctl_rf_c4_rf_chllp_reg[3]/NET0131  & n4577 ;
  assign n6406 = \ctl_rf_c4_rf_chtsz_reg[3]/P0002  & n4579 ;
  assign n6407 = ~n6405 & ~n6406 ;
  assign n6408 = n4687 & ~n6407 ;
  assign n6409 = \ctl_rf_c3_rf_chllp_reg[3]/NET0131  & n4577 ;
  assign n6410 = \ctl_rf_c3_rf_chtsz_reg[3]/P0002  & n4579 ;
  assign n6411 = ~n6409 & ~n6410 ;
  assign n6412 = n4698 & ~n6411 ;
  assign n6413 = ~n6408 & ~n6412 ;
  assign n6414 = n6404 & n6413 ;
  assign n6415 = \ctl_rf_c6_rf_chllp_reg[3]/NET0131  & n4577 ;
  assign n6416 = \ctl_rf_c6_rf_chtsz_reg[3]/P0002  & n4579 ;
  assign n6417 = ~n6415 & ~n6416 ;
  assign n6418 = n4703 & ~n6417 ;
  assign n6419 = \ctl_rf_c5_rf_chllp_reg[3]/NET0131  & n4577 ;
  assign n6420 = \ctl_rf_c5_rf_chtsz_reg[3]/P0002  & n4579 ;
  assign n6421 = ~n6419 & ~n6420 ;
  assign n6422 = n4680 & ~n6421 ;
  assign n6423 = ~n6418 & ~n6422 ;
  assign n6424 = \ctl_rf_c0_rf_chllp_reg[3]/NET0131  & n4577 ;
  assign n6425 = \ctl_rf_c0_rf_chtsz_reg[3]/P0002  & n4579 ;
  assign n6426 = ~n6424 & ~n6425 ;
  assign n6427 = n4675 & ~n6426 ;
  assign n6428 = \ctl_rf_c1_rf_chllp_reg[3]/NET0131  & n4577 ;
  assign n6429 = \ctl_rf_c1_rf_chtsz_reg[3]/P0002  & n4579 ;
  assign n6430 = ~n6428 & ~n6429 ;
  assign n6431 = n4692 & ~n6430 ;
  assign n6432 = ~n6427 & ~n6431 ;
  assign n6433 = n6423 & n6432 ;
  assign n6434 = n6414 & n6433 ;
  assign n6435 = n6395 & n6434 ;
  assign n6436 = n6368 & n6435 ;
  assign n6437 = \haddr[8]_pad  & ~n6436 ;
  assign n6438 = n3024 & n5652 ;
  assign n6439 = \ctl_rf_tc_reg[3]/NET0131  & n4719 ;
  assign n6440 = ~\ctl_rf_c3_rf_int_tc1_msk_reg/NET0131  & \ctl_rf_tc_reg[3]/NET0131  ;
  assign n6441 = n4721 & n6440 ;
  assign n6442 = ~n6439 & ~n6441 ;
  assign n6443 = \ctl_rf_abt_reg[3]/NET0131  & ~\ctl_rf_c3_rf_int_abt_msk_reg/NET0131  ;
  assign n6444 = n4733 & n6443 ;
  assign n6445 = \ctl_rf_sync_reg[3]/NET0131  & n4725 ;
  assign n6446 = \ctl_rf_c3_rf_ch_en_reg/NET0131  & n4727 ;
  assign n6447 = ~n6445 & ~n6446 ;
  assign n6448 = ~n6444 & n6447 ;
  assign n6449 = n6442 & n6448 ;
  assign n6450 = ~n6438 & n6449 ;
  assign n6451 = n4714 & ~n6450 ;
  assign n6452 = n4745 & ~n6451 ;
  assign n6453 = ~n6437 & n6452 ;
  assign n6454 = n6341 & ~n6453 ;
  assign n6455 = ~n4573 & ~n6132 ;
  assign n6456 = ~n6454 & n6455 ;
  assign n6457 = ~n6231 & ~n6456 ;
  assign n6458 = \hrdata_reg[28]_pad  & ~n4569 ;
  assign n6459 = \ctl_rf_c0_rf_chdad_reg[12]/NET0131  & n4582 ;
  assign n6460 = \ctl_rf_c0_rf_swidth_reg[1]/NET0131  & n4577 ;
  assign n6461 = \ctl_rf_c0_rf_chsad_reg[12]/P0002  & n4584 ;
  assign n6462 = ~n6460 & ~n6461 ;
  assign n6463 = ~n6459 & n6462 ;
  assign n6464 = n4623 & ~n6463 ;
  assign n6465 = \ctl_rf_c7_rf_chsad_reg[12]/NET0131  & n4584 ;
  assign n6466 = \ctl_rf_c7_rf_swidth_reg[1]/NET0131  & n4577 ;
  assign n6467 = \ctl_rf_c7_rf_chdad_reg[12]/P0002  & n4582 ;
  assign n6468 = ~n6466 & ~n6467 ;
  assign n6469 = ~n6465 & n6468 ;
  assign n6470 = n4642 & ~n6469 ;
  assign n6471 = ~n6464 & ~n6470 ;
  assign n6472 = \ctl_rf_c6_rf_chsad_reg[12]/NET0131  & n4584 ;
  assign n6473 = \ctl_rf_c6_rf_swidth_reg[1]/NET0131  & n4577 ;
  assign n6474 = \ctl_rf_c6_rf_chdad_reg[12]/P0002  & n4582 ;
  assign n6475 = ~n6473 & ~n6474 ;
  assign n6476 = ~n6472 & n6475 ;
  assign n6477 = n4611 & ~n6476 ;
  assign n6478 = \ctl_rf_c1_rf_chdad_reg[12]/NET0131  & n4582 ;
  assign n6479 = \ctl_rf_c1_rf_swidth_reg[1]/NET0131  & n4577 ;
  assign n6480 = \ctl_rf_c1_rf_chsad_reg[12]/P0002  & n4584 ;
  assign n6481 = ~n6479 & ~n6480 ;
  assign n6482 = ~n6478 & n6481 ;
  assign n6483 = n4632 & ~n6482 ;
  assign n6484 = ~n6477 & ~n6483 ;
  assign n6485 = n6471 & n6484 ;
  assign n6486 = \ctl_rf_c5_rf_chsad_reg[12]/NET0131  & n4584 ;
  assign n6487 = \ctl_rf_c5_rf_swidth_reg[1]/NET0131  & n4577 ;
  assign n6488 = \ctl_rf_c5_rf_chdad_reg[12]/P0002  & n4582 ;
  assign n6489 = ~n6487 & ~n6488 ;
  assign n6490 = ~n6486 & n6489 ;
  assign n6491 = n4601 & ~n6490 ;
  assign n6492 = \ctl_rf_c2_rf_chsad_reg[12]/NET0131  & n4584 ;
  assign n6493 = \ctl_rf_c2_rf_swidth_reg[1]/NET0131  & n4577 ;
  assign n6494 = \ctl_rf_c2_rf_chdad_reg[12]/P0002  & n4582 ;
  assign n6495 = ~n6493 & ~n6494 ;
  assign n6496 = ~n6492 & n6495 ;
  assign n6497 = n4590 & ~n6496 ;
  assign n6498 = ~n6491 & ~n6497 ;
  assign n6499 = \ctl_rf_c4_rf_chsad_reg[12]/NET0131  & n4584 ;
  assign n6500 = \ctl_rf_c4_rf_swidth_reg[1]/NET0131  & n4577 ;
  assign n6501 = \ctl_rf_c4_rf_chdad_reg[12]/P0002  & n4582 ;
  assign n6502 = ~n6500 & ~n6501 ;
  assign n6503 = ~n6499 & n6502 ;
  assign n6504 = n4576 & ~n6503 ;
  assign n6505 = \ctl_rf_c3_rf_chdad_reg[12]/NET0131  & n4582 ;
  assign n6506 = \ctl_rf_c3_rf_swidth_reg[1]/NET0131  & n4577 ;
  assign n6507 = \ctl_rf_c3_rf_chsad_reg[12]/P0002  & n4584 ;
  assign n6508 = ~n6506 & ~n6507 ;
  assign n6509 = ~n6505 & n6508 ;
  assign n6510 = n4651 & ~n6509 ;
  assign n6511 = ~n6504 & ~n6510 ;
  assign n6512 = n6498 & n6511 ;
  assign n6513 = n6485 & n6512 ;
  assign n6514 = \ctl_rf_c5_rf_chllp_reg[12]/NET0131  & n4680 ;
  assign n6515 = \ctl_rf_c6_rf_chllp_reg[12]/NET0131  & n4703 ;
  assign n6516 = ~n6514 & ~n6515 ;
  assign n6517 = \ctl_rf_c1_rf_chllp_reg[12]/NET0131  & n4692 ;
  assign n6518 = \ctl_rf_c3_rf_chllp_reg[12]/NET0131  & n4698 ;
  assign n6519 = ~n6517 & ~n6518 ;
  assign n6520 = n6516 & n6519 ;
  assign n6521 = \ctl_rf_c0_rf_chllp_reg[12]/NET0131  & n4675 ;
  assign n6522 = \ctl_rf_c7_rf_chllp_reg[12]/NET0131  & n4669 ;
  assign n6523 = ~n6521 & ~n6522 ;
  assign n6524 = \ctl_rf_c2_rf_chllp_reg[12]/NET0131  & n4663 ;
  assign n6525 = \ctl_rf_c4_rf_chllp_reg[12]/NET0131  & n4687 ;
  assign n6526 = ~n6524 & ~n6525 ;
  assign n6527 = n6523 & n6526 ;
  assign n6528 = n6520 & n6527 ;
  assign n6529 = n4577 & ~n6528 ;
  assign n6530 = n4573 & ~n6529 ;
  assign n6531 = n6513 & n6530 ;
  assign n6532 = ~n5155 & ~n6531 ;
  assign n6533 = n4569 & n6532 ;
  assign n6534 = ~n6458 & ~n6533 ;
  assign n6535 = \ctl_rf_c5dmabs_reg[28]/NET0131  & \haddr[4]_pad  ;
  assign n6536 = n4579 & n6535 ;
  assign n6537 = \ctl_rf_c6dmabs_reg[28]/NET0131  & \haddr[4]_pad  ;
  assign n6538 = n4584 & n6537 ;
  assign n6539 = ~n6536 & ~n6538 ;
  assign n6540 = \ctl_rf_c1dmabs_reg[28]/NET0131  & ~\haddr[4]_pad  ;
  assign n6541 = n4579 & n6540 ;
  assign n6542 = \ctl_rf_c2dmabs_reg[28]/NET0131  & ~\haddr[4]_pad  ;
  assign n6543 = n4584 & n6542 ;
  assign n6544 = ~n6541 & ~n6543 ;
  assign n6545 = n6539 & n6544 ;
  assign n6546 = \ctl_rf_c3dmabs_reg[28]/NET0131  & ~\haddr[4]_pad  ;
  assign n6547 = n4582 & n6546 ;
  assign n6548 = \ctl_rf_c4dmabs_reg[28]/NET0131  & \haddr[4]_pad  ;
  assign n6549 = n4577 & n6548 ;
  assign n6550 = ~n6547 & ~n6549 ;
  assign n6551 = \ctl_rf_c0dmabs_reg[28]/NET0131  & ~\haddr[4]_pad  ;
  assign n6552 = n4577 & n6551 ;
  assign n6553 = \ctl_rf_c7dmabs_reg[28]/NET0131  & \haddr[4]_pad  ;
  assign n6554 = n4582 & n6553 ;
  assign n6555 = ~n6552 & ~n6554 ;
  assign n6556 = n6550 & n6555 ;
  assign n6557 = n6545 & n6556 ;
  assign n6558 = n4589 & ~n6557 ;
  assign n6559 = \ctl_rf_c1brbs_reg[28]/NET0131  & ~\haddr[4]_pad  ;
  assign n6560 = n4579 & n6559 ;
  assign n6561 = \ctl_rf_c6brbs_reg[28]/NET0131  & \haddr[4]_pad  ;
  assign n6562 = n4584 & n6561 ;
  assign n6563 = ~n6560 & ~n6562 ;
  assign n6564 = \ctl_rf_c4brbs_reg[28]/NET0131  & \haddr[4]_pad  ;
  assign n6565 = n4577 & n6564 ;
  assign n6566 = \ctl_rf_c3brbs_reg[28]/NET0131  & ~\haddr[4]_pad  ;
  assign n6567 = n4582 & n6566 ;
  assign n6568 = ~n6565 & ~n6567 ;
  assign n6569 = n6563 & n6568 ;
  assign n6570 = \ctl_rf_c2brbs_reg[28]/NET0131  & ~\haddr[4]_pad  ;
  assign n6571 = n4584 & n6570 ;
  assign n6572 = \ctl_rf_c0brbs_reg[28]/NET0131  & ~\haddr[4]_pad  ;
  assign n6573 = n4577 & n6572 ;
  assign n6574 = ~n6571 & ~n6573 ;
  assign n6575 = \ctl_rf_c5brbs_reg[28]/NET0131  & \haddr[4]_pad  ;
  assign n6576 = n4579 & n6575 ;
  assign n6577 = \ctl_rf_c7brbs_reg[28]/NET0131  & \haddr[4]_pad  ;
  assign n6578 = n4582 & n6577 ;
  assign n6579 = ~n6576 & ~n6578 ;
  assign n6580 = n6574 & n6579 ;
  assign n6581 = n6569 & n6580 ;
  assign n6582 = n4575 & ~n6581 ;
  assign n6583 = ~\haddr[8]_pad  & ~n6582 ;
  assign n6584 = ~n6558 & n6583 ;
  assign n6585 = ~n4745 & n6584 ;
  assign n6586 = \ctl_rf_c3_rf_chdad_reg[28]/P0002  & n4582 ;
  assign n6587 = \ctl_rf_c3_rf_chsad_reg[28]/P0002  & n4584 ;
  assign n6588 = ~n6586 & ~n6587 ;
  assign n6589 = n4651 & ~n6588 ;
  assign n6590 = \ctl_rf_c5_rf_chdad_reg[28]/P0002  & n4582 ;
  assign n6591 = \ctl_rf_c5_rf_chsad_reg[28]/P0002  & n4584 ;
  assign n6592 = ~n6590 & ~n6591 ;
  assign n6593 = n4601 & ~n6592 ;
  assign n6594 = \ctl_rf_c6_rf_chdad_reg[28]/P0002  & n4582 ;
  assign n6595 = \ctl_rf_c6_rf_chsad_reg[28]/P0002  & n4584 ;
  assign n6596 = ~n6594 & ~n6595 ;
  assign n6597 = n4611 & ~n6596 ;
  assign n6598 = ~n6593 & ~n6597 ;
  assign n6599 = ~n6589 & n6598 ;
  assign n6600 = \ctl_rf_c0_rf_chdad_reg[28]/P0002  & n4582 ;
  assign n6601 = \ctl_rf_c0_rf_chsad_reg[28]/P0002  & n4584 ;
  assign n6602 = ~n6600 & ~n6601 ;
  assign n6603 = n4623 & ~n6602 ;
  assign n6604 = \haddr[8]_pad  & ~n6603 ;
  assign n6605 = \ctl_rf_c2_rf_chdad_reg[28]/P0002  & n4582 ;
  assign n6606 = \ctl_rf_c2_rf_chsad_reg[28]/P0002  & n4584 ;
  assign n6607 = ~n6605 & ~n6606 ;
  assign n6608 = n4590 & ~n6607 ;
  assign n6609 = \ctl_rf_c4_rf_chdad_reg[28]/P0002  & n4582 ;
  assign n6610 = \ctl_rf_c4_rf_chsad_reg[28]/P0002  & n4584 ;
  assign n6611 = ~n6609 & ~n6610 ;
  assign n6612 = n4576 & ~n6611 ;
  assign n6613 = ~n6608 & ~n6612 ;
  assign n6614 = \ctl_rf_c1_rf_chdad_reg[28]/P0002  & n4582 ;
  assign n6615 = \ctl_rf_c1_rf_chsad_reg[28]/P0002  & n4584 ;
  assign n6616 = ~n6614 & ~n6615 ;
  assign n6617 = n4632 & ~n6616 ;
  assign n6618 = \ctl_rf_c7_rf_chdad_reg[28]/P0002  & n4582 ;
  assign n6619 = \ctl_rf_c7_rf_chsad_reg[28]/P0002  & n4584 ;
  assign n6620 = ~n6618 & ~n6619 ;
  assign n6621 = n4642 & ~n6620 ;
  assign n6622 = ~n6617 & ~n6621 ;
  assign n6623 = n6613 & n6622 ;
  assign n6624 = n6604 & n6623 ;
  assign n6625 = n6599 & n6624 ;
  assign n6626 = \ctl_rf_c4_rf_chllp_reg[28]/NET0131  & n4687 ;
  assign n6627 = \ctl_rf_c0_rf_chllp_reg[28]/NET0131  & n4675 ;
  assign n6628 = ~n6626 & ~n6627 ;
  assign n6629 = \ctl_rf_c3_rf_chllp_reg[28]/NET0131  & n4698 ;
  assign n6630 = \ctl_rf_c1_rf_chllp_reg[28]/NET0131  & n4692 ;
  assign n6631 = ~n6629 & ~n6630 ;
  assign n6632 = n6628 & n6631 ;
  assign n6633 = \ctl_rf_c5_rf_chllp_reg[28]/NET0131  & n4680 ;
  assign n6634 = \ctl_rf_c6_rf_chllp_reg[28]/NET0131  & n4703 ;
  assign n6635 = ~n6633 & ~n6634 ;
  assign n6636 = \ctl_rf_c7_rf_chllp_reg[28]/NET0131  & n4669 ;
  assign n6637 = \ctl_rf_c2_rf_chllp_reg[28]/NET0131  & n4663 ;
  assign n6638 = ~n6636 & ~n6637 ;
  assign n6639 = n6635 & n6638 ;
  assign n6640 = n6632 & n6639 ;
  assign n6641 = n4577 & ~n6640 ;
  assign n6642 = ~n4745 & ~n6641 ;
  assign n6643 = n6625 & n6642 ;
  assign n6644 = ~n6585 & ~n6643 ;
  assign n6645 = \ctl_rf_c4_rf_chsad_reg[4]/NET0131  & n4584 ;
  assign n6646 = \ctl_rf_c4_rf_dad_ctl1_reg/NET0131  & n4577 ;
  assign n6647 = \ctl_rf_c4_rf_chdad_reg[4]/P0002  & n4582 ;
  assign n6648 = ~n6646 & ~n6647 ;
  assign n6649 = ~n6645 & n6648 ;
  assign n6650 = n4576 & ~n6649 ;
  assign n6651 = \ctl_rf_c6_rf_chsad_reg[4]/NET0131  & n4584 ;
  assign n6652 = \ctl_rf_c6_rf_dad_ctl1_reg/NET0131  & n4577 ;
  assign n6653 = \ctl_rf_c6_rf_chdad_reg[4]/P0002  & n4582 ;
  assign n6654 = ~n6652 & ~n6653 ;
  assign n6655 = ~n6651 & n6654 ;
  assign n6656 = n4611 & ~n6655 ;
  assign n6657 = ~n6650 & ~n6656 ;
  assign n6658 = \ctl_rf_c7_rf_chsad_reg[4]/NET0131  & n4584 ;
  assign n6659 = \ctl_rf_c7_rf_dad_ctl1_reg/NET0131  & n4577 ;
  assign n6660 = \ctl_rf_c7_rf_chdad_reg[4]/P0002  & n4582 ;
  assign n6661 = ~n6659 & ~n6660 ;
  assign n6662 = ~n6658 & n6661 ;
  assign n6663 = n4642 & ~n6662 ;
  assign n6664 = \ctl_rf_c1_rf_chsad_reg[4]/NET0131  & n4584 ;
  assign n6665 = \ctl_rf_c1_rf_dad_ctl1_reg/NET0131  & n4577 ;
  assign n6666 = \ctl_rf_c1_rf_chdad_reg[4]/P0002  & n4582 ;
  assign n6667 = ~n6665 & ~n6666 ;
  assign n6668 = ~n6664 & n6667 ;
  assign n6669 = n4632 & ~n6668 ;
  assign n6670 = ~n6663 & ~n6669 ;
  assign n6671 = n6657 & n6670 ;
  assign n6672 = \ctl_rf_c0_rf_chsad_reg[4]/NET0131  & n4584 ;
  assign n6673 = \ctl_rf_c0_rf_dad_ctl1_reg/NET0131  & n4577 ;
  assign n6674 = \ctl_rf_c0_rf_chdad_reg[4]/P0002  & n4582 ;
  assign n6675 = ~n6673 & ~n6674 ;
  assign n6676 = ~n6672 & n6675 ;
  assign n6677 = n4623 & ~n6676 ;
  assign n6678 = \ctl_rf_c5_rf_chsad_reg[4]/NET0131  & n4584 ;
  assign n6679 = \ctl_rf_c5_rf_dad_ctl1_reg/NET0131  & n4577 ;
  assign n6680 = \ctl_rf_c5_rf_chdad_reg[4]/P0002  & n4582 ;
  assign n6681 = ~n6679 & ~n6680 ;
  assign n6682 = ~n6678 & n6681 ;
  assign n6683 = n4601 & ~n6682 ;
  assign n6684 = ~n6677 & ~n6683 ;
  assign n6685 = \ctl_rf_c3_rf_chsad_reg[4]/NET0131  & n4584 ;
  assign n6686 = \ctl_rf_c3_rf_dad_ctl1_reg/NET0131  & n4577 ;
  assign n6687 = \ctl_rf_c3_rf_chdad_reg[4]/P0002  & n4582 ;
  assign n6688 = ~n6686 & ~n6687 ;
  assign n6689 = ~n6685 & n6688 ;
  assign n6690 = n4651 & ~n6689 ;
  assign n6691 = \ctl_rf_c2_rf_chsad_reg[4]/NET0131  & n4584 ;
  assign n6692 = \ctl_rf_c2_rf_dad_ctl1_reg/NET0131  & n4577 ;
  assign n6693 = \ctl_rf_c2_rf_chdad_reg[4]/P0002  & n4582 ;
  assign n6694 = ~n6692 & ~n6693 ;
  assign n6695 = ~n6691 & n6694 ;
  assign n6696 = n4590 & ~n6695 ;
  assign n6697 = ~n6690 & ~n6696 ;
  assign n6698 = n6684 & n6697 ;
  assign n6699 = \ctl_rf_c7_rf_chllp_reg[4]/NET0131  & n4577 ;
  assign n6700 = \ctl_rf_c7_rf_chtsz_reg[4]/NET0131  & n4579 ;
  assign n6701 = ~n6699 & ~n6700 ;
  assign n6702 = n4669 & ~n6701 ;
  assign n6703 = \ctl_rf_c2_rf_chllp_reg[4]/NET0131  & n4577 ;
  assign n6704 = \ctl_rf_c2_rf_chtsz_reg[4]/NET0131  & n4579 ;
  assign n6705 = ~n6703 & ~n6704 ;
  assign n6706 = n4663 & ~n6705 ;
  assign n6707 = ~n6702 & ~n6706 ;
  assign n6708 = \ctl_rf_c1_rf_chllp_reg[4]/NET0131  & n4577 ;
  assign n6709 = \ctl_rf_c1_rf_chtsz_reg[4]/NET0131  & n4579 ;
  assign n6710 = ~n6708 & ~n6709 ;
  assign n6711 = n4692 & ~n6710 ;
  assign n6712 = \ctl_rf_c0_rf_chllp_reg[4]/NET0131  & n4577 ;
  assign n6713 = \ctl_rf_c0_rf_chtsz_reg[4]/NET0131  & n4579 ;
  assign n6714 = ~n6712 & ~n6713 ;
  assign n6715 = n4675 & ~n6714 ;
  assign n6716 = ~n6711 & ~n6715 ;
  assign n6717 = n6707 & n6716 ;
  assign n6718 = \ctl_rf_c5_rf_chllp_reg[4]/NET0131  & n4577 ;
  assign n6719 = \ctl_rf_c5_rf_chtsz_reg[4]/NET0131  & n4579 ;
  assign n6720 = ~n6718 & ~n6719 ;
  assign n6721 = n4680 & ~n6720 ;
  assign n6722 = \ctl_rf_c6_rf_chllp_reg[4]/NET0131  & n4577 ;
  assign n6723 = \ctl_rf_c6_rf_chtsz_reg[4]/NET0131  & n4579 ;
  assign n6724 = ~n6722 & ~n6723 ;
  assign n6725 = n4703 & ~n6724 ;
  assign n6726 = ~n6721 & ~n6725 ;
  assign n6727 = \ctl_rf_c3_rf_chllp_reg[4]/NET0131  & n4577 ;
  assign n6728 = \ctl_rf_c3_rf_chtsz_reg[4]/NET0131  & n4579 ;
  assign n6729 = ~n6727 & ~n6728 ;
  assign n6730 = n4698 & ~n6729 ;
  assign n6731 = \ctl_rf_c4_rf_chllp_reg[4]/NET0131  & n4577 ;
  assign n6732 = \ctl_rf_c4_rf_chtsz_reg[4]/NET0131  & n4579 ;
  assign n6733 = ~n6731 & ~n6732 ;
  assign n6734 = n4687 & ~n6733 ;
  assign n6735 = ~n6730 & ~n6734 ;
  assign n6736 = n6726 & n6735 ;
  assign n6737 = n6717 & n6736 ;
  assign n6738 = n6698 & n6737 ;
  assign n6739 = n6671 & n6738 ;
  assign n6740 = \haddr[8]_pad  & ~n6739 ;
  assign n6741 = n2999 & n4717 ;
  assign n6742 = \ctl_rf_tc_reg[4]/NET0131  & n4719 ;
  assign n6743 = ~\ctl_rf_c4_rf_int_tc1_msk_reg/NET0131  & \ctl_rf_tc_reg[4]/NET0131  ;
  assign n6744 = n4721 & n6743 ;
  assign n6745 = ~n6742 & ~n6744 ;
  assign n6746 = \ctl_rf_abt_reg[4]/NET0131  & ~\ctl_rf_c4_rf_int_abt_msk_reg/NET0131  ;
  assign n6747 = n4733 & n6746 ;
  assign n6748 = \ctl_rf_sync_reg[4]/NET0131  & n4725 ;
  assign n6749 = \ctl_rf_c4_rf_ch_en_reg/NET0131  & n4727 ;
  assign n6750 = ~n6748 & ~n6749 ;
  assign n6751 = ~n6747 & n6750 ;
  assign n6752 = n6745 & n6751 ;
  assign n6753 = ~n6741 & n6752 ;
  assign n6754 = n4714 & ~n6753 ;
  assign n6755 = n4745 & ~n6754 ;
  assign n6756 = ~n6740 & n6755 ;
  assign n6757 = n6644 & ~n6756 ;
  assign n6758 = ~n4573 & ~n6458 ;
  assign n6759 = ~n6757 & n6758 ;
  assign n6760 = ~n6534 & ~n6759 ;
  assign n6761 = \hrdata_reg[29]_pad  & ~n4569 ;
  assign n6762 = \ctl_rf_c7_rf_chdad_reg[13]/NET0131  & n4582 ;
  assign n6763 = \ctl_rf_c7_rf_swidth_reg[2]/NET0131  & n4577 ;
  assign n6764 = \ctl_rf_c7_rf_chsad_reg[13]/P0002  & n4584 ;
  assign n6765 = ~n6763 & ~n6764 ;
  assign n6766 = ~n6762 & n6765 ;
  assign n6767 = n4642 & ~n6766 ;
  assign n6768 = \ctl_rf_c0_rf_chsad_reg[13]/NET0131  & n4584 ;
  assign n6769 = \ctl_rf_c0_rf_swidth_reg[2]/NET0131  & n4577 ;
  assign n6770 = \ctl_rf_c0_rf_chdad_reg[13]/P0002  & n4582 ;
  assign n6771 = ~n6769 & ~n6770 ;
  assign n6772 = ~n6768 & n6771 ;
  assign n6773 = n4623 & ~n6772 ;
  assign n6774 = ~n6767 & ~n6773 ;
  assign n6775 = \ctl_rf_c3_rf_chsad_reg[13]/NET0131  & n4584 ;
  assign n6776 = \ctl_rf_c3_rf_swidth_reg[2]/NET0131  & n4577 ;
  assign n6777 = \ctl_rf_c3_rf_chdad_reg[13]/P0002  & n4582 ;
  assign n6778 = ~n6776 & ~n6777 ;
  assign n6779 = ~n6775 & n6778 ;
  assign n6780 = n4651 & ~n6779 ;
  assign n6781 = \ctl_rf_c5_rf_chdad_reg[13]/NET0131  & n4582 ;
  assign n6782 = \ctl_rf_c5_rf_swidth_reg[2]/NET0131  & n4577 ;
  assign n6783 = \ctl_rf_c5_rf_chsad_reg[13]/P0002  & n4584 ;
  assign n6784 = ~n6782 & ~n6783 ;
  assign n6785 = ~n6781 & n6784 ;
  assign n6786 = n4601 & ~n6785 ;
  assign n6787 = ~n6780 & ~n6786 ;
  assign n6788 = n6774 & n6787 ;
  assign n6789 = \ctl_rf_c6_rf_chdad_reg[13]/NET0131  & n4582 ;
  assign n6790 = \ctl_rf_c6_rf_swidth_reg[2]/NET0131  & n4577 ;
  assign n6791 = \ctl_rf_c6_rf_chsad_reg[13]/P0002  & n4584 ;
  assign n6792 = ~n6790 & ~n6791 ;
  assign n6793 = ~n6789 & n6792 ;
  assign n6794 = n4611 & ~n6793 ;
  assign n6795 = \ctl_rf_c4_rf_chsad_reg[13]/NET0131  & n4584 ;
  assign n6796 = \ctl_rf_c4_rf_swidth_reg[2]/NET0131  & n4577 ;
  assign n6797 = \ctl_rf_c4_rf_chdad_reg[13]/P0002  & n4582 ;
  assign n6798 = ~n6796 & ~n6797 ;
  assign n6799 = ~n6795 & n6798 ;
  assign n6800 = n4576 & ~n6799 ;
  assign n6801 = ~n6794 & ~n6800 ;
  assign n6802 = \ctl_rf_c2_rf_chsad_reg[13]/NET0131  & n4584 ;
  assign n6803 = \ctl_rf_c2_rf_swidth_reg[2]/NET0131  & n4577 ;
  assign n6804 = \ctl_rf_c2_rf_chdad_reg[13]/P0002  & n4582 ;
  assign n6805 = ~n6803 & ~n6804 ;
  assign n6806 = ~n6802 & n6805 ;
  assign n6807 = n4590 & ~n6806 ;
  assign n6808 = \ctl_rf_c1_rf_chdad_reg[13]/NET0131  & n4582 ;
  assign n6809 = \ctl_rf_c1_rf_swidth_reg[2]/NET0131  & n4577 ;
  assign n6810 = \ctl_rf_c1_rf_chsad_reg[13]/P0002  & n4584 ;
  assign n6811 = ~n6809 & ~n6810 ;
  assign n6812 = ~n6808 & n6811 ;
  assign n6813 = n4632 & ~n6812 ;
  assign n6814 = ~n6807 & ~n6813 ;
  assign n6815 = n6801 & n6814 ;
  assign n6816 = n6788 & n6815 ;
  assign n6817 = \ctl_rf_c4_rf_chllp_reg[13]/NET0131  & n4687 ;
  assign n6818 = \ctl_rf_c1_rf_chllp_reg[13]/NET0131  & n4692 ;
  assign n6819 = ~n6817 & ~n6818 ;
  assign n6820 = \ctl_rf_c6_rf_chllp_reg[13]/NET0131  & n4703 ;
  assign n6821 = \ctl_rf_c2_rf_chllp_reg[13]/NET0131  & n4663 ;
  assign n6822 = ~n6820 & ~n6821 ;
  assign n6823 = n6819 & n6822 ;
  assign n6824 = \ctl_rf_c7_rf_chllp_reg[13]/NET0131  & n4669 ;
  assign n6825 = \ctl_rf_c0_rf_chllp_reg[13]/NET0131  & n4675 ;
  assign n6826 = ~n6824 & ~n6825 ;
  assign n6827 = \ctl_rf_c3_rf_chllp_reg[13]/NET0131  & n4698 ;
  assign n6828 = \ctl_rf_c5_rf_chllp_reg[13]/NET0131  & n4680 ;
  assign n6829 = ~n6827 & ~n6828 ;
  assign n6830 = n6826 & n6829 ;
  assign n6831 = n6823 & n6830 ;
  assign n6832 = n4577 & ~n6831 ;
  assign n6833 = n4573 & ~n6832 ;
  assign n6834 = n6816 & n6833 ;
  assign n6835 = ~n5155 & ~n6834 ;
  assign n6836 = n4569 & n6835 ;
  assign n6837 = ~n6761 & ~n6836 ;
  assign n6838 = \ctl_rf_c5dmabs_reg[29]/NET0131  & \haddr[4]_pad  ;
  assign n6839 = n4579 & n6838 ;
  assign n6840 = \ctl_rf_c6dmabs_reg[29]/NET0131  & \haddr[4]_pad  ;
  assign n6841 = n4584 & n6840 ;
  assign n6842 = ~n6839 & ~n6841 ;
  assign n6843 = \ctl_rf_c1dmabs_reg[29]/NET0131  & ~\haddr[4]_pad  ;
  assign n6844 = n4579 & n6843 ;
  assign n6845 = \ctl_rf_c2dmabs_reg[29]/NET0131  & ~\haddr[4]_pad  ;
  assign n6846 = n4584 & n6845 ;
  assign n6847 = ~n6844 & ~n6846 ;
  assign n6848 = n6842 & n6847 ;
  assign n6849 = \ctl_rf_c3dmabs_reg[29]/NET0131  & ~\haddr[4]_pad  ;
  assign n6850 = n4582 & n6849 ;
  assign n6851 = \ctl_rf_c4dmabs_reg[29]/NET0131  & \haddr[4]_pad  ;
  assign n6852 = n4577 & n6851 ;
  assign n6853 = ~n6850 & ~n6852 ;
  assign n6854 = \ctl_rf_c0dmabs_reg[29]/NET0131  & ~\haddr[4]_pad  ;
  assign n6855 = n4577 & n6854 ;
  assign n6856 = \ctl_rf_c7dmabs_reg[29]/NET0131  & \haddr[4]_pad  ;
  assign n6857 = n4582 & n6856 ;
  assign n6858 = ~n6855 & ~n6857 ;
  assign n6859 = n6853 & n6858 ;
  assign n6860 = n6848 & n6859 ;
  assign n6861 = n4589 & ~n6860 ;
  assign n6862 = \ctl_rf_c1brbs_reg[29]/NET0131  & ~\haddr[4]_pad  ;
  assign n6863 = n4579 & n6862 ;
  assign n6864 = \ctl_rf_c6brbs_reg[29]/NET0131  & \haddr[4]_pad  ;
  assign n6865 = n4584 & n6864 ;
  assign n6866 = ~n6863 & ~n6865 ;
  assign n6867 = \ctl_rf_c4brbs_reg[29]/NET0131  & \haddr[4]_pad  ;
  assign n6868 = n4577 & n6867 ;
  assign n6869 = \ctl_rf_c3brbs_reg[29]/NET0131  & ~\haddr[4]_pad  ;
  assign n6870 = n4582 & n6869 ;
  assign n6871 = ~n6868 & ~n6870 ;
  assign n6872 = n6866 & n6871 ;
  assign n6873 = \ctl_rf_c2brbs_reg[29]/NET0131  & ~\haddr[4]_pad  ;
  assign n6874 = n4584 & n6873 ;
  assign n6875 = \ctl_rf_c0brbs_reg[29]/NET0131  & ~\haddr[4]_pad  ;
  assign n6876 = n4577 & n6875 ;
  assign n6877 = ~n6874 & ~n6876 ;
  assign n6878 = \ctl_rf_c5brbs_reg[29]/NET0131  & \haddr[4]_pad  ;
  assign n6879 = n4579 & n6878 ;
  assign n6880 = \ctl_rf_c7brbs_reg[29]/NET0131  & \haddr[4]_pad  ;
  assign n6881 = n4582 & n6880 ;
  assign n6882 = ~n6879 & ~n6881 ;
  assign n6883 = n6877 & n6882 ;
  assign n6884 = n6872 & n6883 ;
  assign n6885 = n4575 & ~n6884 ;
  assign n6886 = ~\haddr[8]_pad  & ~n6885 ;
  assign n6887 = ~n6861 & n6886 ;
  assign n6888 = ~n4745 & n6887 ;
  assign n6889 = \ctl_rf_c6_rf_chdad_reg[29]/P0002  & n4582 ;
  assign n6890 = \ctl_rf_c6_rf_chsad_reg[29]/P0002  & n4584 ;
  assign n6891 = ~n6889 & ~n6890 ;
  assign n6892 = n4611 & ~n6891 ;
  assign n6893 = \ctl_rf_c7_rf_chdad_reg[29]/P0002  & n4582 ;
  assign n6894 = \ctl_rf_c7_rf_chsad_reg[29]/P0002  & n4584 ;
  assign n6895 = ~n6893 & ~n6894 ;
  assign n6896 = n4642 & ~n6895 ;
  assign n6897 = \ctl_rf_c3_rf_chdad_reg[29]/P0002  & n4582 ;
  assign n6898 = \ctl_rf_c3_rf_chsad_reg[29]/P0002  & n4584 ;
  assign n6899 = ~n6897 & ~n6898 ;
  assign n6900 = n4651 & ~n6899 ;
  assign n6901 = ~n6896 & ~n6900 ;
  assign n6902 = ~n6892 & n6901 ;
  assign n6903 = \ctl_rf_c1_rf_chdad_reg[29]/P0002  & n4582 ;
  assign n6904 = \ctl_rf_c1_rf_chsad_reg[29]/P0002  & n4584 ;
  assign n6905 = ~n6903 & ~n6904 ;
  assign n6906 = n4632 & ~n6905 ;
  assign n6907 = \haddr[8]_pad  & ~n6906 ;
  assign n6908 = \ctl_rf_c4_rf_chdad_reg[29]/P0002  & n4582 ;
  assign n6909 = \ctl_rf_c4_rf_chsad_reg[29]/P0002  & n4584 ;
  assign n6910 = ~n6908 & ~n6909 ;
  assign n6911 = n4576 & ~n6910 ;
  assign n6912 = \ctl_rf_c2_rf_chdad_reg[29]/P0002  & n4582 ;
  assign n6913 = \ctl_rf_c2_rf_chsad_reg[29]/P0002  & n4584 ;
  assign n6914 = ~n6912 & ~n6913 ;
  assign n6915 = n4590 & ~n6914 ;
  assign n6916 = ~n6911 & ~n6915 ;
  assign n6917 = \ctl_rf_c0_rf_chdad_reg[29]/P0002  & n4582 ;
  assign n6918 = \ctl_rf_c0_rf_chsad_reg[29]/P0002  & n4584 ;
  assign n6919 = ~n6917 & ~n6918 ;
  assign n6920 = n4623 & ~n6919 ;
  assign n6921 = \ctl_rf_c5_rf_chdad_reg[29]/P0002  & n4582 ;
  assign n6922 = \ctl_rf_c5_rf_chsad_reg[29]/P0002  & n4584 ;
  assign n6923 = ~n6921 & ~n6922 ;
  assign n6924 = n4601 & ~n6923 ;
  assign n6925 = ~n6920 & ~n6924 ;
  assign n6926 = n6916 & n6925 ;
  assign n6927 = n6907 & n6926 ;
  assign n6928 = n6902 & n6927 ;
  assign n6929 = \ctl_rf_c1_rf_chllp_reg[29]/NET0131  & n4692 ;
  assign n6930 = \ctl_rf_c3_rf_chllp_reg[29]/NET0131  & n4698 ;
  assign n6931 = ~n6929 & ~n6930 ;
  assign n6932 = \ctl_rf_c0_rf_chllp_reg[29]/NET0131  & n4675 ;
  assign n6933 = \ctl_rf_c4_rf_chllp_reg[29]/NET0131  & n4687 ;
  assign n6934 = ~n6932 & ~n6933 ;
  assign n6935 = n6931 & n6934 ;
  assign n6936 = \ctl_rf_c6_rf_chllp_reg[29]/NET0131  & n4703 ;
  assign n6937 = \ctl_rf_c5_rf_chllp_reg[29]/NET0131  & n4680 ;
  assign n6938 = ~n6936 & ~n6937 ;
  assign n6939 = \ctl_rf_c2_rf_chllp_reg[29]/NET0131  & n4663 ;
  assign n6940 = \ctl_rf_c7_rf_chllp_reg[29]/NET0131  & n4669 ;
  assign n6941 = ~n6939 & ~n6940 ;
  assign n6942 = n6938 & n6941 ;
  assign n6943 = n6935 & n6942 ;
  assign n6944 = n4577 & ~n6943 ;
  assign n6945 = ~n4745 & ~n6944 ;
  assign n6946 = n6928 & n6945 ;
  assign n6947 = ~n6888 & ~n6946 ;
  assign n6948 = \ctl_rf_c2_rf_chsad_reg[5]/NET0131  & n4584 ;
  assign n6949 = \ctl_rf_c2_rf_sad_ctl0_reg/NET0131  & n4577 ;
  assign n6950 = \ctl_rf_c2_rf_chdad_reg[5]/P0002  & n4582 ;
  assign n6951 = ~n6949 & ~n6950 ;
  assign n6952 = ~n6948 & n6951 ;
  assign n6953 = n4590 & ~n6952 ;
  assign n6954 = \ctl_rf_c3_rf_chsad_reg[5]/NET0131  & n4584 ;
  assign n6955 = \ctl_rf_c3_rf_sad_ctl0_reg/NET0131  & n4577 ;
  assign n6956 = \ctl_rf_c3_rf_chdad_reg[5]/P0002  & n4582 ;
  assign n6957 = ~n6955 & ~n6956 ;
  assign n6958 = ~n6954 & n6957 ;
  assign n6959 = n4651 & ~n6958 ;
  assign n6960 = ~n6953 & ~n6959 ;
  assign n6961 = \ctl_rf_c0_rf_chsad_reg[5]/NET0131  & n4584 ;
  assign n6962 = \ctl_rf_c0_rf_sad_ctl0_reg/NET0131  & n4577 ;
  assign n6963 = \ctl_rf_c0_rf_chdad_reg[5]/P0002  & n4582 ;
  assign n6964 = ~n6962 & ~n6963 ;
  assign n6965 = ~n6961 & n6964 ;
  assign n6966 = n4623 & ~n6965 ;
  assign n6967 = \ctl_rf_c5_rf_chsad_reg[5]/NET0131  & n4584 ;
  assign n6968 = \ctl_rf_c5_rf_sad_ctl0_reg/NET0131  & n4577 ;
  assign n6969 = \ctl_rf_c5_rf_chdad_reg[5]/P0002  & n4582 ;
  assign n6970 = ~n6968 & ~n6969 ;
  assign n6971 = ~n6967 & n6970 ;
  assign n6972 = n4601 & ~n6971 ;
  assign n6973 = ~n6966 & ~n6972 ;
  assign n6974 = n6960 & n6973 ;
  assign n6975 = \ctl_rf_c4_rf_chsad_reg[5]/NET0131  & n4584 ;
  assign n6976 = \ctl_rf_c4_rf_sad_ctl0_reg/NET0131  & n4577 ;
  assign n6977 = \ctl_rf_c4_rf_chdad_reg[5]/P0002  & n4582 ;
  assign n6978 = ~n6976 & ~n6977 ;
  assign n6979 = ~n6975 & n6978 ;
  assign n6980 = n4576 & ~n6979 ;
  assign n6981 = \ctl_rf_c6_rf_chsad_reg[5]/NET0131  & n4584 ;
  assign n6982 = \ctl_rf_c6_rf_sad_ctl0_reg/NET0131  & n4577 ;
  assign n6983 = \ctl_rf_c6_rf_chdad_reg[5]/P0002  & n4582 ;
  assign n6984 = ~n6982 & ~n6983 ;
  assign n6985 = ~n6981 & n6984 ;
  assign n6986 = n4611 & ~n6985 ;
  assign n6987 = ~n6980 & ~n6986 ;
  assign n6988 = \ctl_rf_c7_rf_chsad_reg[5]/NET0131  & n4584 ;
  assign n6989 = \ctl_rf_c7_rf_sad_ctl0_reg/NET0131  & n4577 ;
  assign n6990 = \ctl_rf_c7_rf_chdad_reg[5]/P0002  & n4582 ;
  assign n6991 = ~n6989 & ~n6990 ;
  assign n6992 = ~n6988 & n6991 ;
  assign n6993 = n4642 & ~n6992 ;
  assign n6994 = \ctl_rf_c1_rf_chsad_reg[5]/NET0131  & n4584 ;
  assign n6995 = \ctl_rf_c1_rf_sad_ctl0_reg/NET0131  & n4577 ;
  assign n6996 = \ctl_rf_c1_rf_chdad_reg[5]/P0002  & n4582 ;
  assign n6997 = ~n6995 & ~n6996 ;
  assign n6998 = ~n6994 & n6997 ;
  assign n6999 = n4632 & ~n6998 ;
  assign n7000 = ~n6993 & ~n6999 ;
  assign n7001 = n6987 & n7000 ;
  assign n7002 = \ctl_rf_c0_rf_chllp_reg[5]/NET0131  & n4577 ;
  assign n7003 = \ctl_rf_c0_rf_chtsz_reg[5]/NET0131  & n4579 ;
  assign n7004 = ~n7002 & ~n7003 ;
  assign n7005 = n4675 & ~n7004 ;
  assign n7006 = \ctl_rf_c7_rf_chllp_reg[5]/NET0131  & n4577 ;
  assign n7007 = \ctl_rf_c7_rf_chtsz_reg[5]/NET0131  & n4579 ;
  assign n7008 = ~n7006 & ~n7007 ;
  assign n7009 = n4669 & ~n7008 ;
  assign n7010 = ~n7005 & ~n7009 ;
  assign n7011 = \ctl_rf_c4_rf_chllp_reg[5]/NET0131  & n4577 ;
  assign n7012 = \ctl_rf_c4_rf_chtsz_reg[5]/NET0131  & n4579 ;
  assign n7013 = ~n7011 & ~n7012 ;
  assign n7014 = n4687 & ~n7013 ;
  assign n7015 = \ctl_rf_c3_rf_chllp_reg[5]/NET0131  & n4577 ;
  assign n7016 = \ctl_rf_c3_rf_chtsz_reg[5]/NET0131  & n4579 ;
  assign n7017 = ~n7015 & ~n7016 ;
  assign n7018 = n4698 & ~n7017 ;
  assign n7019 = ~n7014 & ~n7018 ;
  assign n7020 = n7010 & n7019 ;
  assign n7021 = \ctl_rf_c6_rf_chllp_reg[5]/NET0131  & n4577 ;
  assign n7022 = \ctl_rf_c6_rf_chtsz_reg[5]/NET0131  & n4579 ;
  assign n7023 = ~n7021 & ~n7022 ;
  assign n7024 = n4703 & ~n7023 ;
  assign n7025 = \ctl_rf_c2_rf_chllp_reg[5]/NET0131  & n4577 ;
  assign n7026 = \ctl_rf_c2_rf_chtsz_reg[5]/NET0131  & n4579 ;
  assign n7027 = ~n7025 & ~n7026 ;
  assign n7028 = n4663 & ~n7027 ;
  assign n7029 = ~n7024 & ~n7028 ;
  assign n7030 = \ctl_rf_c1_rf_chllp_reg[5]/NET0131  & n4577 ;
  assign n7031 = \ctl_rf_c1_rf_chtsz_reg[5]/NET0131  & n4579 ;
  assign n7032 = ~n7030 & ~n7031 ;
  assign n7033 = n4692 & ~n7032 ;
  assign n7034 = \ctl_rf_c5_rf_chllp_reg[5]/NET0131  & n4577 ;
  assign n7035 = \ctl_rf_c5_rf_chtsz_reg[5]/NET0131  & n4579 ;
  assign n7036 = ~n7034 & ~n7035 ;
  assign n7037 = n4680 & ~n7036 ;
  assign n7038 = ~n7033 & ~n7037 ;
  assign n7039 = n7029 & n7038 ;
  assign n7040 = n7020 & n7039 ;
  assign n7041 = n7001 & n7040 ;
  assign n7042 = n6974 & n7041 ;
  assign n7043 = \haddr[8]_pad  & ~n7042 ;
  assign n7044 = n2999 & n5652 ;
  assign n7045 = \ctl_rf_tc_reg[5]/NET0131  & n4719 ;
  assign n7046 = ~\ctl_rf_c5_rf_int_tc1_msk_reg/NET0131  & \ctl_rf_tc_reg[5]/NET0131  ;
  assign n7047 = n4721 & n7046 ;
  assign n7048 = ~n7045 & ~n7047 ;
  assign n7049 = \ctl_rf_abt_reg[5]/NET0131  & ~\ctl_rf_c5_rf_int_abt_msk_reg/NET0131  ;
  assign n7050 = n4733 & n7049 ;
  assign n7051 = \ctl_rf_sync_reg[5]/NET0131  & n4725 ;
  assign n7052 = \ctl_rf_c5_rf_ch_en_reg/NET0131  & n4727 ;
  assign n7053 = ~n7051 & ~n7052 ;
  assign n7054 = ~n7050 & n7053 ;
  assign n7055 = n7048 & n7054 ;
  assign n7056 = ~n7044 & n7055 ;
  assign n7057 = n4714 & ~n7056 ;
  assign n7058 = n4745 & ~n7057 ;
  assign n7059 = ~n7043 & n7058 ;
  assign n7060 = n6947 & ~n7059 ;
  assign n7061 = ~n4573 & ~n6761 ;
  assign n7062 = ~n7060 & n7061 ;
  assign n7063 = ~n6837 & ~n7062 ;
  assign n7064 = \hrdata_reg[2]_pad  & ~n4569 ;
  assign n7065 = n4569 & ~n4573 ;
  assign n7066 = \ctl_rf_c0_rf_chllp_cnt_reg[2]/NET0131  & n4579 ;
  assign n7067 = \ctl_rf_c0_rf_chdad_reg[18]/NET0131  & n4582 ;
  assign n7068 = ~n7066 & ~n7067 ;
  assign n7069 = \ctl_rf_c0_rf_chsad_reg[18]/NET0131  & n4584 ;
  assign n7070 = \ctl_rf_c0_rf_src_sz_reg[2]/NET0131  & n4577 ;
  assign n7071 = ~n7069 & ~n7070 ;
  assign n7072 = n7068 & n7071 ;
  assign n7073 = n4623 & ~n7072 ;
  assign n7074 = \haddr[8]_pad  & ~n7073 ;
  assign n7075 = \ctl_rf_c2_rf_chllp_cnt_reg[2]/NET0131  & n4579 ;
  assign n7076 = \ctl_rf_c2_rf_chsad_reg[18]/NET0131  & n4584 ;
  assign n7077 = ~n7075 & ~n7076 ;
  assign n7078 = \ctl_rf_c2_rf_src_sz_reg[2]/NET0131  & n4577 ;
  assign n7079 = \ctl_rf_c2_rf_chdad_reg[18]/NET0131  & n4582 ;
  assign n7080 = ~n7078 & ~n7079 ;
  assign n7081 = n7077 & n7080 ;
  assign n7082 = n4590 & ~n7081 ;
  assign n7083 = \ctl_rf_c6_rf_chllp_cnt_reg[2]/NET0131  & n4579 ;
  assign n7084 = \ctl_rf_c6_rf_chdad_reg[18]/NET0131  & n4582 ;
  assign n7085 = ~n7083 & ~n7084 ;
  assign n7086 = \ctl_rf_c6_rf_chsad_reg[18]/NET0131  & n4584 ;
  assign n7087 = \ctl_rf_c6_rf_src_sz_reg[2]/NET0131  & n4577 ;
  assign n7088 = ~n7086 & ~n7087 ;
  assign n7089 = n7085 & n7088 ;
  assign n7090 = n4611 & ~n7089 ;
  assign n7091 = ~n7082 & ~n7090 ;
  assign n7092 = \ctl_rf_c1_rf_src_sz_reg[2]/NET0131  & n4577 ;
  assign n7093 = \ctl_rf_c1_rf_chllp_cnt_reg[2]/NET0131  & n4579 ;
  assign n7094 = ~n7092 & ~n7093 ;
  assign n7095 = \ctl_rf_c1_rf_chdad_reg[18]/NET0131  & n4582 ;
  assign n7096 = \ctl_rf_c1_rf_chsad_reg[18]/NET0131  & n4584 ;
  assign n7097 = ~n7095 & ~n7096 ;
  assign n7098 = n7094 & n7097 ;
  assign n7099 = n4632 & ~n7098 ;
  assign n7100 = \ctl_rf_c7_rf_src_sz_reg[2]/NET0131  & n4577 ;
  assign n7101 = \ctl_rf_c7_rf_chllp_cnt_reg[2]/NET0131  & n4579 ;
  assign n7102 = ~n7100 & ~n7101 ;
  assign n7103 = \ctl_rf_c7_rf_chdad_reg[18]/NET0131  & n4582 ;
  assign n7104 = \ctl_rf_c7_rf_chsad_reg[18]/NET0131  & n4584 ;
  assign n7105 = ~n7103 & ~n7104 ;
  assign n7106 = n7102 & n7105 ;
  assign n7107 = n4642 & ~n7106 ;
  assign n7108 = ~n7099 & ~n7107 ;
  assign n7109 = n7091 & n7108 ;
  assign n7110 = n7074 & n7109 ;
  assign n7111 = \ctl_rf_c5_rf_chllp_reg[18]/NET0131  & n4680 ;
  assign n7112 = \ctl_rf_c3_rf_chllp_reg[18]/NET0131  & n4698 ;
  assign n7113 = ~n7111 & ~n7112 ;
  assign n7114 = \ctl_rf_c0_rf_chllp_reg[18]/NET0131  & n4675 ;
  assign n7115 = \ctl_rf_c4_rf_chllp_reg[18]/NET0131  & n4687 ;
  assign n7116 = ~n7114 & ~n7115 ;
  assign n7117 = n7113 & n7116 ;
  assign n7118 = \ctl_rf_c6_rf_chllp_reg[18]/NET0131  & n4703 ;
  assign n7119 = \ctl_rf_c2_rf_chllp_reg[18]/NET0131  & n4663 ;
  assign n7120 = ~n7118 & ~n7119 ;
  assign n7121 = \ctl_rf_c1_rf_chllp_reg[18]/NET0131  & n4692 ;
  assign n7122 = \ctl_rf_c7_rf_chllp_reg[18]/NET0131  & n4669 ;
  assign n7123 = ~n7121 & ~n7122 ;
  assign n7124 = n7120 & n7123 ;
  assign n7125 = n7117 & n7124 ;
  assign n7126 = n4577 & ~n7125 ;
  assign n7127 = \ctl_rf_c4_rf_src_sz_reg[2]/NET0131  & n4577 ;
  assign n7128 = \ctl_rf_c4_rf_chsad_reg[18]/NET0131  & n4584 ;
  assign n7129 = ~n7127 & ~n7128 ;
  assign n7130 = \ctl_rf_c4_rf_chllp_cnt_reg[2]/NET0131  & n4579 ;
  assign n7131 = \ctl_rf_c4_rf_chdad_reg[18]/NET0131  & n4582 ;
  assign n7132 = ~n7130 & ~n7131 ;
  assign n7133 = n7129 & n7132 ;
  assign n7134 = n4576 & ~n7133 ;
  assign n7135 = \ctl_rf_c5_rf_src_sz_reg[2]/NET0131  & n4577 ;
  assign n7136 = \ctl_rf_c5_rf_chllp_cnt_reg[2]/NET0131  & n4579 ;
  assign n7137 = ~n7135 & ~n7136 ;
  assign n7138 = \ctl_rf_c5_rf_chdad_reg[18]/NET0131  & n4582 ;
  assign n7139 = \ctl_rf_c5_rf_chsad_reg[18]/NET0131  & n4584 ;
  assign n7140 = ~n7138 & ~n7139 ;
  assign n7141 = n7137 & n7140 ;
  assign n7142 = n4601 & ~n7141 ;
  assign n7143 = \ctl_rf_c3_rf_chllp_cnt_reg[2]/NET0131  & n4579 ;
  assign n7144 = \ctl_rf_c3_rf_chdad_reg[18]/NET0131  & n4582 ;
  assign n7145 = ~n7143 & ~n7144 ;
  assign n7146 = \ctl_rf_c3_rf_chsad_reg[18]/NET0131  & n4584 ;
  assign n7147 = \ctl_rf_c3_rf_src_sz_reg[2]/NET0131  & n4577 ;
  assign n7148 = ~n7146 & ~n7147 ;
  assign n7149 = n7145 & n7148 ;
  assign n7150 = n4651 & ~n7149 ;
  assign n7151 = ~n7142 & ~n7150 ;
  assign n7152 = ~n7134 & n7151 ;
  assign n7153 = ~n7126 & n7152 ;
  assign n7154 = n7110 & n7153 ;
  assign n7155 = \ctl_rf_c1brbs_reg[18]/NET0131  & ~\haddr[4]_pad  ;
  assign n7156 = n4579 & n7155 ;
  assign n7157 = \ctl_rf_c3brbs_reg[18]/NET0131  & ~\haddr[4]_pad  ;
  assign n7158 = n4582 & n7157 ;
  assign n7159 = ~n7156 & ~n7158 ;
  assign n7160 = \ctl_rf_c0brbs_reg[18]/NET0131  & ~\haddr[4]_pad  ;
  assign n7161 = n4577 & n7160 ;
  assign n7162 = \ctl_rf_c7brbs_reg[18]/NET0131  & \haddr[4]_pad  ;
  assign n7163 = n4582 & n7162 ;
  assign n7164 = ~n7161 & ~n7163 ;
  assign n7165 = n7159 & n7164 ;
  assign n7166 = \ctl_rf_c6brbs_reg[18]/NET0131  & \haddr[4]_pad  ;
  assign n7167 = n4584 & n7166 ;
  assign n7168 = \ctl_rf_c4brbs_reg[18]/NET0131  & \haddr[4]_pad  ;
  assign n7169 = n4577 & n7168 ;
  assign n7170 = ~n7167 & ~n7169 ;
  assign n7171 = \ctl_rf_c2brbs_reg[18]/NET0131  & ~\haddr[4]_pad  ;
  assign n7172 = n4584 & n7171 ;
  assign n7173 = \ctl_rf_c5brbs_reg[18]/NET0131  & \haddr[4]_pad  ;
  assign n7174 = n4579 & n7173 ;
  assign n7175 = ~n7172 & ~n7174 ;
  assign n7176 = n7170 & n7175 ;
  assign n7177 = n7165 & n7176 ;
  assign n7178 = n4575 & ~n7177 ;
  assign n7179 = \ctl_rf_c2dmabs_reg[18]/NET0131  & ~\haddr[4]_pad  ;
  assign n7180 = n4584 & n7179 ;
  assign n7181 = \ctl_rf_c3dmabs_reg[18]/NET0131  & ~\haddr[4]_pad  ;
  assign n7182 = n4582 & n7181 ;
  assign n7183 = ~n7180 & ~n7182 ;
  assign n7184 = \ctl_rf_c0dmabs_reg[18]/NET0131  & ~\haddr[4]_pad  ;
  assign n7185 = n4577 & n7184 ;
  assign n7186 = \ctl_rf_c6dmabs_reg[18]/NET0131  & \haddr[4]_pad  ;
  assign n7187 = n4584 & n7186 ;
  assign n7188 = ~n7185 & ~n7187 ;
  assign n7189 = n7183 & n7188 ;
  assign n7190 = \ctl_rf_c7dmabs_reg[18]/NET0131  & \haddr[4]_pad  ;
  assign n7191 = n4582 & n7190 ;
  assign n7192 = \ctl_rf_c4dmabs_reg[18]/NET0131  & \haddr[4]_pad  ;
  assign n7193 = n4577 & n7192 ;
  assign n7194 = ~n7191 & ~n7193 ;
  assign n7195 = \ctl_rf_c1dmabs_reg[18]/NET0131  & ~\haddr[4]_pad  ;
  assign n7196 = n4579 & n7195 ;
  assign n7197 = \ctl_rf_c5dmabs_reg[18]/NET0131  & \haddr[4]_pad  ;
  assign n7198 = n4579 & n7197 ;
  assign n7199 = ~n7196 & ~n7198 ;
  assign n7200 = n7194 & n7199 ;
  assign n7201 = n7189 & n7200 ;
  assign n7202 = n4589 & ~n7201 ;
  assign n7203 = \ctl_rf_abt_reg[2]/NET0131  & n4622 ;
  assign n7204 = ~\haddr[8]_pad  & ~n7203 ;
  assign n7205 = ~\ctl_rf_c2_rf_int_abt_msk_reg/NET0131  & n5002 ;
  assign n7206 = n5005 & ~n7205 ;
  assign n7207 = ~n7204 & ~n7206 ;
  assign n7208 = ~n7202 & ~n7207 ;
  assign n7209 = ~n7178 & n7208 ;
  assign n7210 = n4569 & ~n7209 ;
  assign n7211 = ~n7154 & n7210 ;
  assign n7212 = ~n7065 & ~n7211 ;
  assign n7213 = ~n7064 & n7212 ;
  assign n7214 = n4745 & n5936 ;
  assign n7215 = n4745 & ~n5993 ;
  assign n7216 = n5977 & n7215 ;
  assign n7217 = ~n7214 & ~n7216 ;
  assign n7218 = ~n4745 & ~n6125 ;
  assign n7219 = ~n6108 & n7218 ;
  assign n7220 = n7217 & ~n7219 ;
  assign n7221 = ~n4573 & ~n7064 ;
  assign n7222 = ~n7220 & n7221 ;
  assign n7223 = ~n7213 & ~n7222 ;
  assign n7224 = \hrdata_reg[30]_pad  & ~n4569 ;
  assign n7225 = \ctl_rf_c0_rf_autold_reg/NET0131  & n4577 ;
  assign n7226 = \ctl_rf_c0_rf_chdad_reg[14]/NET0131  & n4582 ;
  assign n7227 = \ctl_rf_c0_rf_chsad_reg[14]/P0002  & n4584 ;
  assign n7228 = ~n7226 & ~n7227 ;
  assign n7229 = ~n7225 & n7228 ;
  assign n7230 = n4623 & ~n7229 ;
  assign n7231 = \ctl_rf_c7_rf_autold_reg/NET0131  & n4577 ;
  assign n7232 = \ctl_rf_c7_rf_chdad_reg[14]/NET0131  & n4582 ;
  assign n7233 = \ctl_rf_c7_rf_chsad_reg[14]/P0002  & n4584 ;
  assign n7234 = ~n7232 & ~n7233 ;
  assign n7235 = ~n7231 & n7234 ;
  assign n7236 = n4642 & ~n7235 ;
  assign n7237 = ~n7230 & ~n7236 ;
  assign n7238 = \ctl_rf_c6_rf_autold_reg/NET0131  & n4577 ;
  assign n7239 = \ctl_rf_c6_rf_chsad_reg[14]/NET0131  & n4584 ;
  assign n7240 = \ctl_rf_c6_rf_chdad_reg[14]/P0002  & n4582 ;
  assign n7241 = ~n7239 & ~n7240 ;
  assign n7242 = ~n7238 & n7241 ;
  assign n7243 = n4611 & ~n7242 ;
  assign n7244 = \ctl_rf_c1_rf_autold_reg/NET0131  & n4577 ;
  assign n7245 = \ctl_rf_c1_rf_chdad_reg[14]/NET0131  & n4582 ;
  assign n7246 = \ctl_rf_c1_rf_chsad_reg[14]/P0002  & n4584 ;
  assign n7247 = ~n7245 & ~n7246 ;
  assign n7248 = ~n7244 & n7247 ;
  assign n7249 = n4632 & ~n7248 ;
  assign n7250 = ~n7243 & ~n7249 ;
  assign n7251 = n7237 & n7250 ;
  assign n7252 = \ctl_rf_c3_rf_autold_reg/NET0131  & n4577 ;
  assign n7253 = \ctl_rf_c3_rf_chsad_reg[14]/NET0131  & n4584 ;
  assign n7254 = \ctl_rf_c3_rf_chdad_reg[14]/P0002  & n4582 ;
  assign n7255 = ~n7253 & ~n7254 ;
  assign n7256 = ~n7252 & n7255 ;
  assign n7257 = n4651 & ~n7256 ;
  assign n7258 = \ctl_rf_c2_rf_autold_reg/NET0131  & n4577 ;
  assign n7259 = \ctl_rf_c2_rf_chsad_reg[14]/NET0131  & n4584 ;
  assign n7260 = \ctl_rf_c2_rf_chdad_reg[14]/P0002  & n4582 ;
  assign n7261 = ~n7259 & ~n7260 ;
  assign n7262 = ~n7258 & n7261 ;
  assign n7263 = n4590 & ~n7262 ;
  assign n7264 = ~n7257 & ~n7263 ;
  assign n7265 = \ctl_rf_c4_rf_autold_reg/NET0131  & n4577 ;
  assign n7266 = \ctl_rf_c4_rf_chsad_reg[14]/NET0131  & n4584 ;
  assign n7267 = \ctl_rf_c4_rf_chdad_reg[14]/P0002  & n4582 ;
  assign n7268 = ~n7266 & ~n7267 ;
  assign n7269 = ~n7265 & n7268 ;
  assign n7270 = n4576 & ~n7269 ;
  assign n7271 = \ctl_rf_c5_rf_autold_reg/NET0131  & n4577 ;
  assign n7272 = \ctl_rf_c5_rf_chsad_reg[14]/NET0131  & n4584 ;
  assign n7273 = \ctl_rf_c5_rf_chdad_reg[14]/P0002  & n4582 ;
  assign n7274 = ~n7272 & ~n7273 ;
  assign n7275 = ~n7271 & n7274 ;
  assign n7276 = n4601 & ~n7275 ;
  assign n7277 = ~n7270 & ~n7276 ;
  assign n7278 = n7264 & n7277 ;
  assign n7279 = n7251 & n7278 ;
  assign n7280 = \ctl_rf_c5_rf_chllp_reg[14]/NET0131  & n4680 ;
  assign n7281 = \ctl_rf_c6_rf_chllp_reg[14]/NET0131  & n4703 ;
  assign n7282 = ~n7280 & ~n7281 ;
  assign n7283 = \ctl_rf_c1_rf_chllp_reg[14]/NET0131  & n4692 ;
  assign n7284 = \ctl_rf_c3_rf_chllp_reg[14]/NET0131  & n4698 ;
  assign n7285 = ~n7283 & ~n7284 ;
  assign n7286 = n7282 & n7285 ;
  assign n7287 = \ctl_rf_c0_rf_chllp_reg[14]/NET0131  & n4675 ;
  assign n7288 = \ctl_rf_c7_rf_chllp_reg[14]/NET0131  & n4669 ;
  assign n7289 = ~n7287 & ~n7288 ;
  assign n7290 = \ctl_rf_c2_rf_chllp_reg[14]/NET0131  & n4663 ;
  assign n7291 = \ctl_rf_c4_rf_chllp_reg[14]/NET0131  & n4687 ;
  assign n7292 = ~n7290 & ~n7291 ;
  assign n7293 = n7289 & n7292 ;
  assign n7294 = n7286 & n7293 ;
  assign n7295 = n4577 & ~n7294 ;
  assign n7296 = n4573 & ~n7295 ;
  assign n7297 = n7279 & n7296 ;
  assign n7298 = ~n5155 & ~n7297 ;
  assign n7299 = n4569 & n7298 ;
  assign n7300 = ~n7224 & ~n7299 ;
  assign n7301 = \ctl_rf_c5dmabs_reg[30]/NET0131  & \haddr[4]_pad  ;
  assign n7302 = n4579 & n7301 ;
  assign n7303 = \ctl_rf_c6dmabs_reg[30]/NET0131  & \haddr[4]_pad  ;
  assign n7304 = n4584 & n7303 ;
  assign n7305 = ~n7302 & ~n7304 ;
  assign n7306 = \ctl_rf_c1dmabs_reg[30]/NET0131  & ~\haddr[4]_pad  ;
  assign n7307 = n4579 & n7306 ;
  assign n7308 = \ctl_rf_c2dmabs_reg[30]/NET0131  & ~\haddr[4]_pad  ;
  assign n7309 = n4584 & n7308 ;
  assign n7310 = ~n7307 & ~n7309 ;
  assign n7311 = n7305 & n7310 ;
  assign n7312 = \ctl_rf_c3dmabs_reg[30]/NET0131  & ~\haddr[4]_pad  ;
  assign n7313 = n4582 & n7312 ;
  assign n7314 = \ctl_rf_c4dmabs_reg[30]/NET0131  & \haddr[4]_pad  ;
  assign n7315 = n4577 & n7314 ;
  assign n7316 = ~n7313 & ~n7315 ;
  assign n7317 = \ctl_rf_c0dmabs_reg[30]/NET0131  & ~\haddr[4]_pad  ;
  assign n7318 = n4577 & n7317 ;
  assign n7319 = \ctl_rf_c7dmabs_reg[30]/NET0131  & \haddr[4]_pad  ;
  assign n7320 = n4582 & n7319 ;
  assign n7321 = ~n7318 & ~n7320 ;
  assign n7322 = n7316 & n7321 ;
  assign n7323 = n7311 & n7322 ;
  assign n7324 = n4589 & ~n7323 ;
  assign n7325 = \ctl_rf_c1brbs_reg[30]/NET0131  & ~\haddr[4]_pad  ;
  assign n7326 = n4579 & n7325 ;
  assign n7327 = \ctl_rf_c7brbs_reg[30]/NET0131  & \haddr[4]_pad  ;
  assign n7328 = n4582 & n7327 ;
  assign n7329 = ~n7326 & ~n7328 ;
  assign n7330 = \ctl_rf_c4brbs_reg[30]/NET0131  & \haddr[4]_pad  ;
  assign n7331 = n4577 & n7330 ;
  assign n7332 = \ctl_rf_c5brbs_reg[30]/NET0131  & \haddr[4]_pad  ;
  assign n7333 = n4579 & n7332 ;
  assign n7334 = ~n7331 & ~n7333 ;
  assign n7335 = n7329 & n7334 ;
  assign n7336 = \ctl_rf_c2brbs_reg[30]/NET0131  & ~\haddr[4]_pad  ;
  assign n7337 = n4584 & n7336 ;
  assign n7338 = \ctl_rf_c0brbs_reg[30]/NET0131  & ~\haddr[4]_pad  ;
  assign n7339 = n4577 & n7338 ;
  assign n7340 = ~n7337 & ~n7339 ;
  assign n7341 = \ctl_rf_c3brbs_reg[30]/NET0131  & ~\haddr[4]_pad  ;
  assign n7342 = n4582 & n7341 ;
  assign n7343 = \ctl_rf_c6brbs_reg[30]/NET0131  & \haddr[4]_pad  ;
  assign n7344 = n4584 & n7343 ;
  assign n7345 = ~n7342 & ~n7344 ;
  assign n7346 = n7340 & n7345 ;
  assign n7347 = n7335 & n7346 ;
  assign n7348 = n4575 & ~n7347 ;
  assign n7349 = ~\haddr[8]_pad  & ~n7348 ;
  assign n7350 = ~n7324 & n7349 ;
  assign n7351 = ~n4745 & n7350 ;
  assign n7352 = \ctl_rf_c6_rf_chdad_reg[30]/P0002  & n4582 ;
  assign n7353 = \ctl_rf_c6_rf_chsad_reg[30]/P0002  & n4584 ;
  assign n7354 = ~n7352 & ~n7353 ;
  assign n7355 = n4611 & ~n7354 ;
  assign n7356 = \ctl_rf_c7_rf_chdad_reg[30]/P0002  & n4582 ;
  assign n7357 = \ctl_rf_c7_rf_chsad_reg[30]/P0002  & n4584 ;
  assign n7358 = ~n7356 & ~n7357 ;
  assign n7359 = n4642 & ~n7358 ;
  assign n7360 = \ctl_rf_c3_rf_chdad_reg[30]/P0002  & n4582 ;
  assign n7361 = \ctl_rf_c3_rf_chsad_reg[30]/P0002  & n4584 ;
  assign n7362 = ~n7360 & ~n7361 ;
  assign n7363 = n4651 & ~n7362 ;
  assign n7364 = ~n7359 & ~n7363 ;
  assign n7365 = ~n7355 & n7364 ;
  assign n7366 = \ctl_rf_c1_rf_chdad_reg[30]/P0002  & n4582 ;
  assign n7367 = \ctl_rf_c1_rf_chsad_reg[30]/P0002  & n4584 ;
  assign n7368 = ~n7366 & ~n7367 ;
  assign n7369 = n4632 & ~n7368 ;
  assign n7370 = \haddr[8]_pad  & ~n7369 ;
  assign n7371 = \ctl_rf_c4_rf_chdad_reg[30]/P0002  & n4582 ;
  assign n7372 = \ctl_rf_c4_rf_chsad_reg[30]/P0002  & n4584 ;
  assign n7373 = ~n7371 & ~n7372 ;
  assign n7374 = n4576 & ~n7373 ;
  assign n7375 = \ctl_rf_c2_rf_chdad_reg[30]/P0002  & n4582 ;
  assign n7376 = \ctl_rf_c2_rf_chsad_reg[30]/P0002  & n4584 ;
  assign n7377 = ~n7375 & ~n7376 ;
  assign n7378 = n4590 & ~n7377 ;
  assign n7379 = ~n7374 & ~n7378 ;
  assign n7380 = \ctl_rf_c0_rf_chdad_reg[30]/P0002  & n4582 ;
  assign n7381 = \ctl_rf_c0_rf_chsad_reg[30]/P0002  & n4584 ;
  assign n7382 = ~n7380 & ~n7381 ;
  assign n7383 = n4623 & ~n7382 ;
  assign n7384 = \ctl_rf_c5_rf_chdad_reg[30]/P0002  & n4582 ;
  assign n7385 = \ctl_rf_c5_rf_chsad_reg[30]/P0002  & n4584 ;
  assign n7386 = ~n7384 & ~n7385 ;
  assign n7387 = n4601 & ~n7386 ;
  assign n7388 = ~n7383 & ~n7387 ;
  assign n7389 = n7379 & n7388 ;
  assign n7390 = n7370 & n7389 ;
  assign n7391 = n7365 & n7390 ;
  assign n7392 = \ctl_rf_c1_rf_chllp_reg[30]/NET0131  & n4692 ;
  assign n7393 = \ctl_rf_c3_rf_chllp_reg[30]/NET0131  & n4698 ;
  assign n7394 = ~n7392 & ~n7393 ;
  assign n7395 = \ctl_rf_c0_rf_chllp_reg[30]/NET0131  & n4675 ;
  assign n7396 = \ctl_rf_c4_rf_chllp_reg[30]/NET0131  & n4687 ;
  assign n7397 = ~n7395 & ~n7396 ;
  assign n7398 = n7394 & n7397 ;
  assign n7399 = \ctl_rf_c6_rf_chllp_reg[30]/NET0131  & n4703 ;
  assign n7400 = \ctl_rf_c5_rf_chllp_reg[30]/NET0131  & n4680 ;
  assign n7401 = ~n7399 & ~n7400 ;
  assign n7402 = \ctl_rf_c2_rf_chllp_reg[30]/NET0131  & n4663 ;
  assign n7403 = \ctl_rf_c7_rf_chllp_reg[30]/NET0131  & n4669 ;
  assign n7404 = ~n7402 & ~n7403 ;
  assign n7405 = n7401 & n7404 ;
  assign n7406 = n7398 & n7405 ;
  assign n7407 = n4577 & ~n7406 ;
  assign n7408 = ~n4745 & ~n7407 ;
  assign n7409 = n7391 & n7408 ;
  assign n7410 = ~n7351 & ~n7409 ;
  assign n7411 = \ctl_rf_c5_rf_chsad_reg[6]/NET0131  & n4584 ;
  assign n7412 = \ctl_rf_c5_rf_sad_ctl1_reg/NET0131  & n4577 ;
  assign n7413 = \ctl_rf_c5_rf_chdad_reg[6]/P0002  & n4582 ;
  assign n7414 = ~n7412 & ~n7413 ;
  assign n7415 = ~n7411 & n7414 ;
  assign n7416 = n4601 & ~n7415 ;
  assign n7417 = \ctl_rf_c2_rf_chsad_reg[6]/NET0131  & n4584 ;
  assign n7418 = \ctl_rf_c2_rf_sad_ctl1_reg/NET0131  & n4577 ;
  assign n7419 = \ctl_rf_c2_rf_chdad_reg[6]/P0002  & n4582 ;
  assign n7420 = ~n7418 & ~n7419 ;
  assign n7421 = ~n7417 & n7420 ;
  assign n7422 = n4590 & ~n7421 ;
  assign n7423 = ~n7416 & ~n7422 ;
  assign n7424 = \ctl_rf_c0_rf_chsad_reg[6]/NET0131  & n4584 ;
  assign n7425 = \ctl_rf_c0_rf_sad_ctl1_reg/NET0131  & n4577 ;
  assign n7426 = \ctl_rf_c0_rf_chdad_reg[6]/P0002  & n4582 ;
  assign n7427 = ~n7425 & ~n7426 ;
  assign n7428 = ~n7424 & n7427 ;
  assign n7429 = n4623 & ~n7428 ;
  assign n7430 = \ctl_rf_c3_rf_chsad_reg[6]/NET0131  & n4584 ;
  assign n7431 = \ctl_rf_c3_rf_sad_ctl1_reg/NET0131  & n4577 ;
  assign n7432 = \ctl_rf_c3_rf_chdad_reg[6]/P0002  & n4582 ;
  assign n7433 = ~n7431 & ~n7432 ;
  assign n7434 = ~n7430 & n7433 ;
  assign n7435 = n4651 & ~n7434 ;
  assign n7436 = ~n7429 & ~n7435 ;
  assign n7437 = n7423 & n7436 ;
  assign n7438 = \ctl_rf_c7_rf_chsad_reg[6]/NET0131  & n4584 ;
  assign n7439 = \ctl_rf_c7_rf_sad_ctl1_reg/NET0131  & n4577 ;
  assign n7440 = \ctl_rf_c7_rf_chdad_reg[6]/P0002  & n4582 ;
  assign n7441 = ~n7439 & ~n7440 ;
  assign n7442 = ~n7438 & n7441 ;
  assign n7443 = n4642 & ~n7442 ;
  assign n7444 = \ctl_rf_c4_rf_chsad_reg[6]/NET0131  & n4584 ;
  assign n7445 = \ctl_rf_c4_rf_sad_ctl1_reg/NET0131  & n4577 ;
  assign n7446 = \ctl_rf_c4_rf_chdad_reg[6]/P0002  & n4582 ;
  assign n7447 = ~n7445 & ~n7446 ;
  assign n7448 = ~n7444 & n7447 ;
  assign n7449 = n4576 & ~n7448 ;
  assign n7450 = ~n7443 & ~n7449 ;
  assign n7451 = \ctl_rf_c1_rf_chsad_reg[6]/NET0131  & n4584 ;
  assign n7452 = \ctl_rf_c1_rf_sad_ctl1_reg/NET0131  & n4577 ;
  assign n7453 = \ctl_rf_c1_rf_chdad_reg[6]/P0002  & n4582 ;
  assign n7454 = ~n7452 & ~n7453 ;
  assign n7455 = ~n7451 & n7454 ;
  assign n7456 = n4632 & ~n7455 ;
  assign n7457 = \ctl_rf_c6_rf_chsad_reg[6]/NET0131  & n4584 ;
  assign n7458 = \ctl_rf_c6_rf_sad_ctl1_reg/NET0131  & n4577 ;
  assign n7459 = \ctl_rf_c6_rf_chdad_reg[6]/P0002  & n4582 ;
  assign n7460 = ~n7458 & ~n7459 ;
  assign n7461 = ~n7457 & n7460 ;
  assign n7462 = n4611 & ~n7461 ;
  assign n7463 = ~n7456 & ~n7462 ;
  assign n7464 = n7450 & n7463 ;
  assign n7465 = \ctl_rf_c2_rf_chllp_reg[6]/NET0131  & n4577 ;
  assign n7466 = \ctl_rf_c2_rf_chtsz_reg[6]/NET0131  & n4579 ;
  assign n7467 = ~n7465 & ~n7466 ;
  assign n7468 = n4663 & ~n7467 ;
  assign n7469 = \ctl_rf_c3_rf_chllp_reg[6]/NET0131  & n4577 ;
  assign n7470 = \ctl_rf_c3_rf_chtsz_reg[6]/NET0131  & n4579 ;
  assign n7471 = ~n7469 & ~n7470 ;
  assign n7472 = n4698 & ~n7471 ;
  assign n7473 = ~n7468 & ~n7472 ;
  assign n7474 = \ctl_rf_c7_rf_chllp_reg[6]/NET0131  & n4577 ;
  assign n7475 = \ctl_rf_c7_rf_chtsz_reg[6]/NET0131  & n4579 ;
  assign n7476 = ~n7474 & ~n7475 ;
  assign n7477 = n4669 & ~n7476 ;
  assign n7478 = \ctl_rf_c4_rf_chllp_reg[6]/NET0131  & n4577 ;
  assign n7479 = \ctl_rf_c4_rf_chtsz_reg[6]/NET0131  & n4579 ;
  assign n7480 = ~n7478 & ~n7479 ;
  assign n7481 = n4687 & ~n7480 ;
  assign n7482 = ~n7477 & ~n7481 ;
  assign n7483 = n7473 & n7482 ;
  assign n7484 = \ctl_rf_c6_rf_chllp_reg[6]/NET0131  & n4577 ;
  assign n7485 = \ctl_rf_c6_rf_chtsz_reg[6]/NET0131  & n4579 ;
  assign n7486 = ~n7484 & ~n7485 ;
  assign n7487 = n4703 & ~n7486 ;
  assign n7488 = \ctl_rf_c5_rf_chllp_reg[6]/NET0131  & n4577 ;
  assign n7489 = \ctl_rf_c5_rf_chtsz_reg[6]/NET0131  & n4579 ;
  assign n7490 = ~n7488 & ~n7489 ;
  assign n7491 = n4680 & ~n7490 ;
  assign n7492 = ~n7487 & ~n7491 ;
  assign n7493 = \ctl_rf_c0_rf_chllp_reg[6]/NET0131  & n4577 ;
  assign n7494 = \ctl_rf_c0_rf_chtsz_reg[6]/NET0131  & n4579 ;
  assign n7495 = ~n7493 & ~n7494 ;
  assign n7496 = n4675 & ~n7495 ;
  assign n7497 = \ctl_rf_c1_rf_chllp_reg[6]/NET0131  & n4577 ;
  assign n7498 = \ctl_rf_c1_rf_chtsz_reg[6]/NET0131  & n4579 ;
  assign n7499 = ~n7497 & ~n7498 ;
  assign n7500 = n4692 & ~n7499 ;
  assign n7501 = ~n7496 & ~n7500 ;
  assign n7502 = n7492 & n7501 ;
  assign n7503 = n7483 & n7502 ;
  assign n7504 = n7464 & n7503 ;
  assign n7505 = n7437 & n7504 ;
  assign n7506 = \haddr[8]_pad  & ~n7505 ;
  assign n7507 = n3011 & n4717 ;
  assign n7508 = \ctl_rf_tc_reg[6]/NET0131  & n4719 ;
  assign n7509 = ~\ctl_rf_c6_rf_int_tc1_msk_reg/NET0131  & \ctl_rf_tc_reg[6]/NET0131  ;
  assign n7510 = n4721 & n7509 ;
  assign n7511 = ~n7508 & ~n7510 ;
  assign n7512 = \ctl_rf_abt_reg[6]/NET0131  & ~\ctl_rf_c6_rf_int_abt_msk_reg/NET0131  ;
  assign n7513 = n4733 & n7512 ;
  assign n7514 = \ctl_rf_sync_reg[6]/NET0131  & n4725 ;
  assign n7515 = \ctl_rf_c6_rf_ch_en_reg/NET0131  & n4727 ;
  assign n7516 = ~n7514 & ~n7515 ;
  assign n7517 = ~n7513 & n7516 ;
  assign n7518 = n7511 & n7517 ;
  assign n7519 = ~n7507 & n7518 ;
  assign n7520 = n4714 & ~n7519 ;
  assign n7521 = n4745 & ~n7520 ;
  assign n7522 = ~n7506 & n7521 ;
  assign n7523 = n7410 & ~n7522 ;
  assign n7524 = ~n4573 & ~n7224 ;
  assign n7525 = ~n7523 & n7524 ;
  assign n7526 = ~n7300 & ~n7525 ;
  assign n7527 = \hrdata_reg[31]_pad  & ~n4569 ;
  assign n7528 = \ctl_rf_c0_rf_chdad_reg[15]/NET0131  & n4582 ;
  assign n7529 = \ctl_rf_c0_rf_chabt_reg/NET0131  & n4577 ;
  assign n7530 = \ctl_rf_c0_rf_chsad_reg[15]/P0002  & n4584 ;
  assign n7531 = ~n7529 & ~n7530 ;
  assign n7532 = ~n7528 & n7531 ;
  assign n7533 = n4623 & ~n7532 ;
  assign n7534 = \ctl_rf_c6_rf_chsad_reg[15]/NET0131  & n4584 ;
  assign n7535 = \ctl_rf_c6_rf_chabt_reg/NET0131  & n4577 ;
  assign n7536 = \ctl_rf_c6_rf_chdad_reg[15]/P0002  & n4582 ;
  assign n7537 = ~n7535 & ~n7536 ;
  assign n7538 = ~n7534 & n7537 ;
  assign n7539 = n4611 & ~n7538 ;
  assign n7540 = ~n7533 & ~n7539 ;
  assign n7541 = \ctl_rf_c7_rf_chdad_reg[15]/NET0131  & n4582 ;
  assign n7542 = \ctl_rf_c7_rf_chabt_reg/NET0131  & n4577 ;
  assign n7543 = \ctl_rf_c7_rf_chsad_reg[15]/P0002  & n4584 ;
  assign n7544 = ~n7542 & ~n7543 ;
  assign n7545 = ~n7541 & n7544 ;
  assign n7546 = n4642 & ~n7545 ;
  assign n7547 = \ctl_rf_c1_rf_chdad_reg[15]/NET0131  & n4582 ;
  assign n7548 = \ctl_rf_c1_rf_chabt_reg/NET0131  & n4577 ;
  assign n7549 = \ctl_rf_c1_rf_chsad_reg[15]/P0002  & n4584 ;
  assign n7550 = ~n7548 & ~n7549 ;
  assign n7551 = ~n7547 & n7550 ;
  assign n7552 = n4632 & ~n7551 ;
  assign n7553 = ~n7546 & ~n7552 ;
  assign n7554 = n7540 & n7553 ;
  assign n7555 = \ctl_rf_c3_rf_chdad_reg[15]/NET0131  & n4582 ;
  assign n7556 = \ctl_rf_c3_rf_chabt_reg/NET0131  & n4577 ;
  assign n7557 = \ctl_rf_c3_rf_chsad_reg[15]/P0002  & n4584 ;
  assign n7558 = ~n7556 & ~n7557 ;
  assign n7559 = ~n7555 & n7558 ;
  assign n7560 = n4651 & ~n7559 ;
  assign n7561 = \ctl_rf_c2_rf_chsad_reg[15]/NET0131  & n4584 ;
  assign n7562 = \ctl_rf_c2_rf_chabt_reg/NET0131  & n4577 ;
  assign n7563 = \ctl_rf_c2_rf_chdad_reg[15]/P0002  & n4582 ;
  assign n7564 = ~n7562 & ~n7563 ;
  assign n7565 = ~n7561 & n7564 ;
  assign n7566 = n4590 & ~n7565 ;
  assign n7567 = ~n7560 & ~n7566 ;
  assign n7568 = \ctl_rf_c4_rf_chsad_reg[15]/NET0131  & n4584 ;
  assign n7569 = \ctl_rf_c4_rf_chabt_reg/NET0131  & n4577 ;
  assign n7570 = \ctl_rf_c4_rf_chdad_reg[15]/P0002  & n4582 ;
  assign n7571 = ~n7569 & ~n7570 ;
  assign n7572 = ~n7568 & n7571 ;
  assign n7573 = n4576 & ~n7572 ;
  assign n7574 = \ctl_rf_c5_rf_chsad_reg[15]/NET0131  & n4584 ;
  assign n7575 = \ctl_rf_c5_rf_chabt_reg/NET0131  & n4577 ;
  assign n7576 = \ctl_rf_c5_rf_chdad_reg[15]/P0002  & n4582 ;
  assign n7577 = ~n7575 & ~n7576 ;
  assign n7578 = ~n7574 & n7577 ;
  assign n7579 = n4601 & ~n7578 ;
  assign n7580 = ~n7573 & ~n7579 ;
  assign n7581 = n7567 & n7580 ;
  assign n7582 = n7554 & n7581 ;
  assign n7583 = \ctl_rf_c5_rf_chllp_reg[15]/NET0131  & n4680 ;
  assign n7584 = \ctl_rf_c6_rf_chllp_reg[15]/NET0131  & n4703 ;
  assign n7585 = ~n7583 & ~n7584 ;
  assign n7586 = \ctl_rf_c0_rf_chllp_reg[15]/NET0131  & n4675 ;
  assign n7587 = \ctl_rf_c3_rf_chllp_reg[15]/NET0131  & n4698 ;
  assign n7588 = ~n7586 & ~n7587 ;
  assign n7589 = n7585 & n7588 ;
  assign n7590 = \ctl_rf_c1_rf_chllp_reg[15]/NET0131  & n4692 ;
  assign n7591 = \ctl_rf_c7_rf_chllp_reg[15]/NET0131  & n4669 ;
  assign n7592 = ~n7590 & ~n7591 ;
  assign n7593 = \ctl_rf_c2_rf_chllp_reg[15]/NET0131  & n4663 ;
  assign n7594 = \ctl_rf_c4_rf_chllp_reg[15]/NET0131  & n4687 ;
  assign n7595 = ~n7593 & ~n7594 ;
  assign n7596 = n7592 & n7595 ;
  assign n7597 = n7589 & n7596 ;
  assign n7598 = n4577 & ~n7597 ;
  assign n7599 = n4573 & ~n7598 ;
  assign n7600 = n7582 & n7599 ;
  assign n7601 = ~n5155 & ~n7600 ;
  assign n7602 = n4569 & n7601 ;
  assign n7603 = ~n7527 & ~n7602 ;
  assign n7604 = \haddr[8]_pad  & ~n4632 ;
  assign n7605 = \ctl_rf_c1_rf_int_tc_msk_reg/NET0131  & n4577 ;
  assign n7606 = \ctl_rf_c1_rf_chdad_reg[31]/P0002  & n4582 ;
  assign n7607 = ~n7605 & ~n7606 ;
  assign n7608 = \ctl_rf_c1_rf_chsad_reg[31]/NET0131  & n4584 ;
  assign n7609 = \haddr[8]_pad  & ~n7608 ;
  assign n7610 = n7607 & n7609 ;
  assign n7611 = ~n7604 & ~n7610 ;
  assign n7612 = \ctl_rf_c7_rf_chsad_reg[31]/NET0131  & n4584 ;
  assign n7613 = \ctl_rf_c7_rf_int_tc_msk_reg/NET0131  & n4577 ;
  assign n7614 = \ctl_rf_c7_rf_chdad_reg[31]/P0002  & n4582 ;
  assign n7615 = ~n7613 & ~n7614 ;
  assign n7616 = ~n7612 & n7615 ;
  assign n7617 = n4642 & ~n7616 ;
  assign n7618 = \ctl_rf_c0_rf_chdad_reg[31]/P0002  & n4582 ;
  assign n7619 = \ctl_rf_c0_rf_chsad_reg[31]/NET0131  & n4584 ;
  assign n7620 = \ctl_rf_c0_rf_int_tc_msk_reg/NET0131  & n4577 ;
  assign n7621 = ~n7619 & ~n7620 ;
  assign n7622 = ~n7618 & n7621 ;
  assign n7623 = n4623 & ~n7622 ;
  assign n7624 = ~n7617 & ~n7623 ;
  assign n7625 = \ctl_rf_c5_rf_chsad_reg[31]/NET0131  & n4584 ;
  assign n7626 = \ctl_rf_c5_rf_int_tc_msk_reg/NET0131  & n4577 ;
  assign n7627 = \ctl_rf_c5_rf_chdad_reg[31]/P0002  & n4582 ;
  assign n7628 = ~n7626 & ~n7627 ;
  assign n7629 = ~n7625 & n7628 ;
  assign n7630 = n4601 & ~n7629 ;
  assign n7631 = \ctl_rf_c2_rf_chsad_reg[31]/NET0131  & n4584 ;
  assign n7632 = \ctl_rf_c2_rf_int_tc_msk_reg/NET0131  & n4577 ;
  assign n7633 = \ctl_rf_c2_rf_chdad_reg[31]/P0002  & n4582 ;
  assign n7634 = ~n7632 & ~n7633 ;
  assign n7635 = ~n7631 & n7634 ;
  assign n7636 = n4590 & ~n7635 ;
  assign n7637 = ~n7630 & ~n7636 ;
  assign n7638 = n7624 & n7637 ;
  assign n7639 = ~n7611 & n7638 ;
  assign n7640 = \ctl_rf_c5_rf_chllp_reg[31]/NET0131  & n4680 ;
  assign n7641 = \ctl_rf_c0_rf_chllp_reg[31]/NET0131  & n4675 ;
  assign n7642 = ~n7640 & ~n7641 ;
  assign n7643 = \ctl_rf_c2_rf_chllp_reg[31]/NET0131  & n4663 ;
  assign n7644 = \ctl_rf_c6_rf_chllp_reg[31]/NET0131  & n4703 ;
  assign n7645 = ~n7643 & ~n7644 ;
  assign n7646 = n7642 & n7645 ;
  assign n7647 = \ctl_rf_c1_rf_chllp_reg[31]/NET0131  & n4692 ;
  assign n7648 = \ctl_rf_c3_rf_chllp_reg[31]/NET0131  & n4698 ;
  assign n7649 = ~n7647 & ~n7648 ;
  assign n7650 = \ctl_rf_c4_rf_chllp_reg[31]/NET0131  & n4687 ;
  assign n7651 = \ctl_rf_c7_rf_chllp_reg[31]/NET0131  & n4669 ;
  assign n7652 = ~n7650 & ~n7651 ;
  assign n7653 = n7649 & n7652 ;
  assign n7654 = n7646 & n7653 ;
  assign n7655 = n4577 & ~n7654 ;
  assign n7656 = \ctl_rf_c3_rf_chdad_reg[31]/P0002  & n4582 ;
  assign n7657 = \ctl_rf_c3_rf_chsad_reg[31]/NET0131  & n4584 ;
  assign n7658 = \ctl_rf_c3_rf_int_tc_msk_reg/NET0131  & n4577 ;
  assign n7659 = ~n7657 & ~n7658 ;
  assign n7660 = ~n7656 & n7659 ;
  assign n7661 = n4651 & ~n7660 ;
  assign n7662 = \ctl_rf_c4_rf_chsad_reg[31]/NET0131  & n4584 ;
  assign n7663 = \ctl_rf_c4_rf_int_tc_msk_reg/NET0131  & n4577 ;
  assign n7664 = \ctl_rf_c4_rf_chdad_reg[31]/P0002  & n4582 ;
  assign n7665 = ~n7663 & ~n7664 ;
  assign n7666 = ~n7662 & n7665 ;
  assign n7667 = n4576 & ~n7666 ;
  assign n7668 = \ctl_rf_c6_rf_chsad_reg[31]/NET0131  & n4584 ;
  assign n7669 = \ctl_rf_c6_rf_int_tc_msk_reg/NET0131  & n4577 ;
  assign n7670 = \ctl_rf_c6_rf_chdad_reg[31]/P0002  & n4582 ;
  assign n7671 = ~n7669 & ~n7670 ;
  assign n7672 = ~n7668 & n7671 ;
  assign n7673 = n4611 & ~n7672 ;
  assign n7674 = ~n7667 & ~n7673 ;
  assign n7675 = ~n7661 & n7674 ;
  assign n7676 = ~n7655 & n7675 ;
  assign n7677 = n7639 & n7676 ;
  assign n7678 = \ctl_rf_c5brbs_reg[31]/NET0131  & \haddr[4]_pad  ;
  assign n7679 = n4579 & n7678 ;
  assign n7680 = \ctl_rf_c6brbs_reg[31]/NET0131  & \haddr[4]_pad  ;
  assign n7681 = n4584 & n7680 ;
  assign n7682 = ~n7679 & ~n7681 ;
  assign n7683 = \ctl_rf_c1brbs_reg[31]/NET0131  & ~\haddr[4]_pad  ;
  assign n7684 = n4579 & n7683 ;
  assign n7685 = \ctl_rf_c2brbs_reg[31]/NET0131  & ~\haddr[4]_pad  ;
  assign n7686 = n4584 & n7685 ;
  assign n7687 = ~n7684 & ~n7686 ;
  assign n7688 = n7682 & n7687 ;
  assign n7689 = \ctl_rf_c3brbs_reg[31]/NET0131  & ~\haddr[4]_pad  ;
  assign n7690 = n4582 & n7689 ;
  assign n7691 = \ctl_rf_c4brbs_reg[31]/NET0131  & \haddr[4]_pad  ;
  assign n7692 = n4577 & n7691 ;
  assign n7693 = ~n7690 & ~n7692 ;
  assign n7694 = \ctl_rf_c0brbs_reg[31]/NET0131  & ~\haddr[4]_pad  ;
  assign n7695 = n4577 & n7694 ;
  assign n7696 = \ctl_rf_c7brbs_reg[31]/NET0131  & \haddr[4]_pad  ;
  assign n7697 = n4582 & n7696 ;
  assign n7698 = ~n7695 & ~n7697 ;
  assign n7699 = n7693 & n7698 ;
  assign n7700 = n7688 & n7699 ;
  assign n7701 = n4575 & ~n7700 ;
  assign n7702 = \ctl_rf_c1dmabs_reg[31]/NET0131  & ~\haddr[4]_pad  ;
  assign n7703 = n4579 & n7702 ;
  assign n7704 = \ctl_rf_c6dmabs_reg[31]/NET0131  & \haddr[4]_pad  ;
  assign n7705 = n4584 & n7704 ;
  assign n7706 = ~n7703 & ~n7705 ;
  assign n7707 = \ctl_rf_c4dmabs_reg[31]/NET0131  & \haddr[4]_pad  ;
  assign n7708 = n4577 & n7707 ;
  assign n7709 = \ctl_rf_c3dmabs_reg[31]/NET0131  & ~\haddr[4]_pad  ;
  assign n7710 = n4582 & n7709 ;
  assign n7711 = ~n7708 & ~n7710 ;
  assign n7712 = n7706 & n7711 ;
  assign n7713 = \ctl_rf_c2dmabs_reg[31]/NET0131  & ~\haddr[4]_pad  ;
  assign n7714 = n4584 & n7713 ;
  assign n7715 = \ctl_rf_c0dmabs_reg[31]/NET0131  & ~\haddr[4]_pad  ;
  assign n7716 = n4577 & n7715 ;
  assign n7717 = ~n7714 & ~n7716 ;
  assign n7718 = \ctl_rf_c5dmabs_reg[31]/NET0131  & \haddr[4]_pad  ;
  assign n7719 = n4579 & n7718 ;
  assign n7720 = \ctl_rf_c7dmabs_reg[31]/NET0131  & \haddr[4]_pad  ;
  assign n7721 = n4582 & n7720 ;
  assign n7722 = ~n7719 & ~n7721 ;
  assign n7723 = n7717 & n7722 ;
  assign n7724 = n7712 & n7723 ;
  assign n7725 = n4589 & ~n7724 ;
  assign n7726 = ~\haddr[8]_pad  & ~n7725 ;
  assign n7727 = ~n7701 & n7726 ;
  assign n7728 = ~n7677 & ~n7727 ;
  assign n7729 = ~n4745 & ~n7728 ;
  assign n7730 = \ctl_rf_c4_rf_chsad_reg[7]/NET0131  & n4584 ;
  assign n7731 = \ctl_rf_c4_rf_mode_reg/NET0131  & n4577 ;
  assign n7732 = \ctl_rf_c4_rf_chdad_reg[7]/P0002  & n4582 ;
  assign n7733 = ~n7731 & ~n7732 ;
  assign n7734 = ~n7730 & n7733 ;
  assign n7735 = n4576 & ~n7734 ;
  assign n7736 = \ctl_rf_c6_rf_chsad_reg[7]/NET0131  & n4584 ;
  assign n7737 = \ctl_rf_c6_rf_mode_reg/NET0131  & n4577 ;
  assign n7738 = \ctl_rf_c6_rf_chdad_reg[7]/P0002  & n4582 ;
  assign n7739 = ~n7737 & ~n7738 ;
  assign n7740 = ~n7736 & n7739 ;
  assign n7741 = n4611 & ~n7740 ;
  assign n7742 = ~n7735 & ~n7741 ;
  assign n7743 = \ctl_rf_c7_rf_chsad_reg[7]/NET0131  & n4584 ;
  assign n7744 = \ctl_rf_c7_rf_mode_reg/NET0131  & n4577 ;
  assign n7745 = \ctl_rf_c7_rf_chdad_reg[7]/P0002  & n4582 ;
  assign n7746 = ~n7744 & ~n7745 ;
  assign n7747 = ~n7743 & n7746 ;
  assign n7748 = n4642 & ~n7747 ;
  assign n7749 = \ctl_rf_c1_rf_chsad_reg[7]/NET0131  & n4584 ;
  assign n7750 = \ctl_rf_c1_rf_mode_reg/NET0131  & n4577 ;
  assign n7751 = \ctl_rf_c1_rf_chdad_reg[7]/P0002  & n4582 ;
  assign n7752 = ~n7750 & ~n7751 ;
  assign n7753 = ~n7749 & n7752 ;
  assign n7754 = n4632 & ~n7753 ;
  assign n7755 = ~n7748 & ~n7754 ;
  assign n7756 = n7742 & n7755 ;
  assign n7757 = \ctl_rf_c0_rf_chsad_reg[7]/NET0131  & n4584 ;
  assign n7758 = \ctl_rf_c0_rf_mode_reg/NET0131  & n4577 ;
  assign n7759 = \ctl_rf_c0_rf_chdad_reg[7]/P0002  & n4582 ;
  assign n7760 = ~n7758 & ~n7759 ;
  assign n7761 = ~n7757 & n7760 ;
  assign n7762 = n4623 & ~n7761 ;
  assign n7763 = \ctl_rf_c5_rf_chsad_reg[7]/NET0131  & n4584 ;
  assign n7764 = \ctl_rf_c5_rf_mode_reg/NET0131  & n4577 ;
  assign n7765 = \ctl_rf_c5_rf_chdad_reg[7]/P0002  & n4582 ;
  assign n7766 = ~n7764 & ~n7765 ;
  assign n7767 = ~n7763 & n7766 ;
  assign n7768 = n4601 & ~n7767 ;
  assign n7769 = ~n7762 & ~n7768 ;
  assign n7770 = \ctl_rf_c3_rf_chsad_reg[7]/NET0131  & n4584 ;
  assign n7771 = \ctl_rf_c3_rf_mode_reg/NET0131  & n4577 ;
  assign n7772 = \ctl_rf_c3_rf_chdad_reg[7]/P0002  & n4582 ;
  assign n7773 = ~n7771 & ~n7772 ;
  assign n7774 = ~n7770 & n7773 ;
  assign n7775 = n4651 & ~n7774 ;
  assign n7776 = \ctl_rf_c2_rf_chsad_reg[7]/NET0131  & n4584 ;
  assign n7777 = \ctl_rf_c2_rf_mode_reg/NET0131  & n4577 ;
  assign n7778 = \ctl_rf_c2_rf_chdad_reg[7]/P0002  & n4582 ;
  assign n7779 = ~n7777 & ~n7778 ;
  assign n7780 = ~n7776 & n7779 ;
  assign n7781 = n4590 & ~n7780 ;
  assign n7782 = ~n7775 & ~n7781 ;
  assign n7783 = n7769 & n7782 ;
  assign n7784 = \ctl_rf_c3_rf_chllp_reg[7]/NET0131  & n4577 ;
  assign n7785 = \ctl_rf_c3_rf_chtsz_reg[7]/NET0131  & n4579 ;
  assign n7786 = ~n7784 & ~n7785 ;
  assign n7787 = n4698 & ~n7786 ;
  assign n7788 = \ctl_rf_c0_rf_chllp_reg[7]/NET0131  & n4577 ;
  assign n7789 = \ctl_rf_c0_rf_chtsz_reg[7]/NET0131  & n4579 ;
  assign n7790 = ~n7788 & ~n7789 ;
  assign n7791 = n4675 & ~n7790 ;
  assign n7792 = ~n7787 & ~n7791 ;
  assign n7793 = \ctl_rf_c5_rf_chllp_reg[7]/NET0131  & n4577 ;
  assign n7794 = \ctl_rf_c5_rf_chtsz_reg[7]/NET0131  & n4579 ;
  assign n7795 = ~n7793 & ~n7794 ;
  assign n7796 = n4680 & ~n7795 ;
  assign n7797 = \ctl_rf_c1_rf_chllp_reg[7]/NET0131  & n4577 ;
  assign n7798 = \ctl_rf_c1_rf_chtsz_reg[7]/NET0131  & n4579 ;
  assign n7799 = ~n7797 & ~n7798 ;
  assign n7800 = n4692 & ~n7799 ;
  assign n7801 = ~n7796 & ~n7800 ;
  assign n7802 = n7792 & n7801 ;
  assign n7803 = \ctl_rf_c2_rf_chllp_reg[7]/NET0131  & n4577 ;
  assign n7804 = \ctl_rf_c2_rf_chtsz_reg[7]/NET0131  & n4579 ;
  assign n7805 = ~n7803 & ~n7804 ;
  assign n7806 = n4663 & ~n7805 ;
  assign n7807 = \ctl_rf_c7_rf_chllp_reg[7]/NET0131  & n4577 ;
  assign n7808 = \ctl_rf_c7_rf_chtsz_reg[7]/NET0131  & n4579 ;
  assign n7809 = ~n7807 & ~n7808 ;
  assign n7810 = n4669 & ~n7809 ;
  assign n7811 = ~n7806 & ~n7810 ;
  assign n7812 = \ctl_rf_c4_rf_chllp_reg[7]/NET0131  & n4577 ;
  assign n7813 = \ctl_rf_c4_rf_chtsz_reg[7]/NET0131  & n4579 ;
  assign n7814 = ~n7812 & ~n7813 ;
  assign n7815 = n4687 & ~n7814 ;
  assign n7816 = \ctl_rf_c6_rf_chllp_reg[7]/NET0131  & n4577 ;
  assign n7817 = \ctl_rf_c6_rf_chtsz_reg[7]/NET0131  & n4579 ;
  assign n7818 = ~n7816 & ~n7817 ;
  assign n7819 = n4703 & ~n7818 ;
  assign n7820 = ~n7815 & ~n7819 ;
  assign n7821 = n7811 & n7820 ;
  assign n7822 = n7802 & n7821 ;
  assign n7823 = n7783 & n7822 ;
  assign n7824 = n7756 & n7823 ;
  assign n7825 = \haddr[8]_pad  & ~n7824 ;
  assign n7826 = n3011 & n5652 ;
  assign n7827 = \ctl_rf_tc_reg[7]/NET0131  & n4719 ;
  assign n7828 = ~\ctl_rf_c7_rf_int_tc1_msk_reg/NET0131  & \ctl_rf_tc_reg[7]/NET0131  ;
  assign n7829 = n4721 & n7828 ;
  assign n7830 = ~n7827 & ~n7829 ;
  assign n7831 = \ctl_rf_abt_reg[7]/NET0131  & ~\ctl_rf_c7_rf_int_abt_msk_reg/NET0131  ;
  assign n7832 = n4733 & n7831 ;
  assign n7833 = \ctl_rf_sync_reg[7]/NET0131  & n4725 ;
  assign n7834 = \ctl_rf_c7_rf_ch_en_reg/NET0131  & n4727 ;
  assign n7835 = ~n7833 & ~n7834 ;
  assign n7836 = ~n7832 & n7835 ;
  assign n7837 = n7830 & n7836 ;
  assign n7838 = ~n7826 & n7837 ;
  assign n7839 = n4714 & ~n7838 ;
  assign n7840 = n4745 & ~n7839 ;
  assign n7841 = ~n7825 & n7840 ;
  assign n7842 = ~n7729 & ~n7841 ;
  assign n7843 = ~n4573 & ~n7527 ;
  assign n7844 = ~n7842 & n7843 ;
  assign n7845 = ~n7603 & ~n7844 ;
  assign n7846 = \hrdata_reg[3]_pad  & ~n4569 ;
  assign n7847 = \ctl_rf_c0_rf_chllp_cnt_reg[3]/NET0131  & n4579 ;
  assign n7848 = \ctl_rf_c0_rf_chdad_reg[19]/NET0131  & n4582 ;
  assign n7849 = ~n7847 & ~n7848 ;
  assign n7850 = \ctl_rf_c0_rf_chsad_reg[19]/NET0131  & n4584 ;
  assign n7851 = \ctl_rf_c0_rf_prot1_reg/NET0131  & n4577 ;
  assign n7852 = ~n7850 & ~n7851 ;
  assign n7853 = n7849 & n7852 ;
  assign n7854 = n4623 & ~n7853 ;
  assign n7855 = \haddr[8]_pad  & ~n7854 ;
  assign n7856 = \ctl_rf_c2_rf_chllp_cnt_reg[3]/NET0131  & n4579 ;
  assign n7857 = \ctl_rf_c2_rf_chsad_reg[19]/NET0131  & n4584 ;
  assign n7858 = ~n7856 & ~n7857 ;
  assign n7859 = \ctl_rf_c2_rf_prot1_reg/NET0131  & n4577 ;
  assign n7860 = \ctl_rf_c2_rf_chdad_reg[19]/NET0131  & n4582 ;
  assign n7861 = ~n7859 & ~n7860 ;
  assign n7862 = n7858 & n7861 ;
  assign n7863 = n4590 & ~n7862 ;
  assign n7864 = \ctl_rf_c4_rf_chllp_cnt_reg[3]/NET0131  & n4579 ;
  assign n7865 = \ctl_rf_c4_rf_chdad_reg[19]/NET0131  & n4582 ;
  assign n7866 = ~n7864 & ~n7865 ;
  assign n7867 = \ctl_rf_c4_rf_chsad_reg[19]/NET0131  & n4584 ;
  assign n7868 = \ctl_rf_c4_rf_prot1_reg/NET0131  & n4577 ;
  assign n7869 = ~n7867 & ~n7868 ;
  assign n7870 = n7866 & n7869 ;
  assign n7871 = n4576 & ~n7870 ;
  assign n7872 = ~n7863 & ~n7871 ;
  assign n7873 = \ctl_rf_c7_rf_prot1_reg/NET0131  & n4577 ;
  assign n7874 = \ctl_rf_c7_rf_chllp_cnt_reg[3]/NET0131  & n4579 ;
  assign n7875 = ~n7873 & ~n7874 ;
  assign n7876 = \ctl_rf_c7_rf_chdad_reg[19]/NET0131  & n4582 ;
  assign n7877 = \ctl_rf_c7_rf_chsad_reg[19]/NET0131  & n4584 ;
  assign n7878 = ~n7876 & ~n7877 ;
  assign n7879 = n7875 & n7878 ;
  assign n7880 = n4642 & ~n7879 ;
  assign n7881 = \ctl_rf_c1_rf_prot1_reg/NET0131  & n4577 ;
  assign n7882 = \ctl_rf_c1_rf_chllp_cnt_reg[3]/NET0131  & n4579 ;
  assign n7883 = ~n7881 & ~n7882 ;
  assign n7884 = \ctl_rf_c1_rf_chdad_reg[19]/NET0131  & n4582 ;
  assign n7885 = \ctl_rf_c1_rf_chsad_reg[19]/NET0131  & n4584 ;
  assign n7886 = ~n7884 & ~n7885 ;
  assign n7887 = n7883 & n7886 ;
  assign n7888 = n4632 & ~n7887 ;
  assign n7889 = ~n7880 & ~n7888 ;
  assign n7890 = n7872 & n7889 ;
  assign n7891 = n7855 & n7890 ;
  assign n7892 = \ctl_rf_c1_rf_chllp_reg[19]/NET0131  & n4692 ;
  assign n7893 = \ctl_rf_c3_rf_chllp_reg[19]/NET0131  & n4698 ;
  assign n7894 = ~n7892 & ~n7893 ;
  assign n7895 = \ctl_rf_c0_rf_chllp_reg[19]/NET0131  & n4675 ;
  assign n7896 = \ctl_rf_c4_rf_chllp_reg[19]/NET0131  & n4687 ;
  assign n7897 = ~n7895 & ~n7896 ;
  assign n7898 = n7894 & n7897 ;
  assign n7899 = \ctl_rf_c6_rf_chllp_reg[19]/NET0131  & n4703 ;
  assign n7900 = \ctl_rf_c5_rf_chllp_reg[19]/NET0131  & n4680 ;
  assign n7901 = ~n7899 & ~n7900 ;
  assign n7902 = \ctl_rf_c2_rf_chllp_reg[19]/NET0131  & n4663 ;
  assign n7903 = \ctl_rf_c7_rf_chllp_reg[19]/NET0131  & n4669 ;
  assign n7904 = ~n7902 & ~n7903 ;
  assign n7905 = n7901 & n7904 ;
  assign n7906 = n7898 & n7905 ;
  assign n7907 = n4577 & ~n7906 ;
  assign n7908 = \ctl_rf_c6_rf_prot1_reg/NET0131  & n4577 ;
  assign n7909 = \ctl_rf_c6_rf_chsad_reg[19]/NET0131  & n4584 ;
  assign n7910 = ~n7908 & ~n7909 ;
  assign n7911 = \ctl_rf_c6_rf_chllp_cnt_reg[3]/NET0131  & n4579 ;
  assign n7912 = \ctl_rf_c6_rf_chdad_reg[19]/NET0131  & n4582 ;
  assign n7913 = ~n7911 & ~n7912 ;
  assign n7914 = n7910 & n7913 ;
  assign n7915 = n4611 & ~n7914 ;
  assign n7916 = \ctl_rf_c5_rf_prot1_reg/NET0131  & n4577 ;
  assign n7917 = \ctl_rf_c5_rf_chllp_cnt_reg[3]/NET0131  & n4579 ;
  assign n7918 = ~n7916 & ~n7917 ;
  assign n7919 = \ctl_rf_c5_rf_chdad_reg[19]/NET0131  & n4582 ;
  assign n7920 = \ctl_rf_c5_rf_chsad_reg[19]/NET0131  & n4584 ;
  assign n7921 = ~n7919 & ~n7920 ;
  assign n7922 = n7918 & n7921 ;
  assign n7923 = n4601 & ~n7922 ;
  assign n7924 = \ctl_rf_c3_rf_chllp_cnt_reg[3]/NET0131  & n4579 ;
  assign n7925 = \ctl_rf_c3_rf_chdad_reg[19]/NET0131  & n4582 ;
  assign n7926 = ~n7924 & ~n7925 ;
  assign n7927 = \ctl_rf_c3_rf_chsad_reg[19]/NET0131  & n4584 ;
  assign n7928 = \ctl_rf_c3_rf_prot1_reg/NET0131  & n4577 ;
  assign n7929 = ~n7927 & ~n7928 ;
  assign n7930 = n7926 & n7929 ;
  assign n7931 = n4651 & ~n7930 ;
  assign n7932 = ~n7923 & ~n7931 ;
  assign n7933 = ~n7915 & n7932 ;
  assign n7934 = ~n7907 & n7933 ;
  assign n7935 = n7891 & n7934 ;
  assign n7936 = \ctl_rf_c1dmabs_reg[19]/NET0131  & ~\haddr[4]_pad  ;
  assign n7937 = n4579 & n7936 ;
  assign n7938 = \ctl_rf_c3dmabs_reg[19]/NET0131  & ~\haddr[4]_pad  ;
  assign n7939 = n4582 & n7938 ;
  assign n7940 = ~n7937 & ~n7939 ;
  assign n7941 = \ctl_rf_c0dmabs_reg[19]/NET0131  & ~\haddr[4]_pad  ;
  assign n7942 = n4577 & n7941 ;
  assign n7943 = \ctl_rf_c7dmabs_reg[19]/NET0131  & \haddr[4]_pad  ;
  assign n7944 = n4582 & n7943 ;
  assign n7945 = ~n7942 & ~n7944 ;
  assign n7946 = n7940 & n7945 ;
  assign n7947 = \ctl_rf_c6dmabs_reg[19]/NET0131  & \haddr[4]_pad  ;
  assign n7948 = n4584 & n7947 ;
  assign n7949 = \ctl_rf_c4dmabs_reg[19]/NET0131  & \haddr[4]_pad  ;
  assign n7950 = n4577 & n7949 ;
  assign n7951 = ~n7948 & ~n7950 ;
  assign n7952 = \ctl_rf_c2dmabs_reg[19]/NET0131  & ~\haddr[4]_pad  ;
  assign n7953 = n4584 & n7952 ;
  assign n7954 = \ctl_rf_c5dmabs_reg[19]/NET0131  & \haddr[4]_pad  ;
  assign n7955 = n4579 & n7954 ;
  assign n7956 = ~n7953 & ~n7955 ;
  assign n7957 = n7951 & n7956 ;
  assign n7958 = n7946 & n7957 ;
  assign n7959 = n4589 & ~n7958 ;
  assign n7960 = \ctl_rf_c2brbs_reg[19]/NET0131  & ~\haddr[4]_pad  ;
  assign n7961 = n4584 & n7960 ;
  assign n7962 = \ctl_rf_c3brbs_reg[19]/NET0131  & ~\haddr[4]_pad  ;
  assign n7963 = n4582 & n7962 ;
  assign n7964 = ~n7961 & ~n7963 ;
  assign n7965 = \ctl_rf_c0brbs_reg[19]/NET0131  & ~\haddr[4]_pad  ;
  assign n7966 = n4577 & n7965 ;
  assign n7967 = \ctl_rf_c6brbs_reg[19]/NET0131  & \haddr[4]_pad  ;
  assign n7968 = n4584 & n7967 ;
  assign n7969 = ~n7966 & ~n7968 ;
  assign n7970 = n7964 & n7969 ;
  assign n7971 = \ctl_rf_c7brbs_reg[19]/NET0131  & \haddr[4]_pad  ;
  assign n7972 = n4582 & n7971 ;
  assign n7973 = \ctl_rf_c4brbs_reg[19]/NET0131  & \haddr[4]_pad  ;
  assign n7974 = n4577 & n7973 ;
  assign n7975 = ~n7972 & ~n7974 ;
  assign n7976 = \ctl_rf_c1brbs_reg[19]/NET0131  & ~\haddr[4]_pad  ;
  assign n7977 = n4579 & n7976 ;
  assign n7978 = \ctl_rf_c5brbs_reg[19]/NET0131  & \haddr[4]_pad  ;
  assign n7979 = n4579 & n7978 ;
  assign n7980 = ~n7977 & ~n7979 ;
  assign n7981 = n7975 & n7980 ;
  assign n7982 = n7970 & n7981 ;
  assign n7983 = n4575 & ~n7982 ;
  assign n7984 = \ctl_rf_abt_reg[3]/NET0131  & n4622 ;
  assign n7985 = ~\haddr[8]_pad  & ~n7984 ;
  assign n7986 = ~\ctl_rf_c3_rf_int_abt_msk_reg/NET0131  & n5002 ;
  assign n7987 = n5005 & ~n7986 ;
  assign n7988 = ~n7985 & ~n7987 ;
  assign n7989 = ~n7983 & ~n7988 ;
  assign n7990 = ~n7959 & n7989 ;
  assign n7991 = n4569 & ~n7990 ;
  assign n7992 = ~n7935 & n7991 ;
  assign n7993 = ~n7065 & ~n7992 ;
  assign n7994 = ~n7846 & n7993 ;
  assign n7995 = n4745 & n6281 ;
  assign n7996 = n4745 & ~n6338 ;
  assign n7997 = n6322 & n7996 ;
  assign n7998 = ~n7995 & ~n7997 ;
  assign n7999 = ~n4745 & ~n6451 ;
  assign n8000 = ~n6437 & n7999 ;
  assign n8001 = n7998 & ~n8000 ;
  assign n8002 = ~n4573 & ~n7846 ;
  assign n8003 = ~n8001 & n8002 ;
  assign n8004 = ~n7994 & ~n8003 ;
  assign n8005 = \hrdata_reg[4]_pad  & ~n4569 ;
  assign n8006 = \haddr[8]_pad  & ~n4576 ;
  assign n8007 = \ctl_rf_c4_rf_prot2_reg/NET0131  & n4577 ;
  assign n8008 = \ctl_rf_c4_rf_chdad_reg[20]/P0002  & n4582 ;
  assign n8009 = ~n8007 & ~n8008 ;
  assign n8010 = \ctl_rf_c4_rf_chsad_reg[20]/NET0131  & n4584 ;
  assign n8011 = \haddr[8]_pad  & ~n8010 ;
  assign n8012 = n8009 & n8011 ;
  assign n8013 = ~n8006 & ~n8012 ;
  assign n8014 = \ctl_rf_c6_rf_chsad_reg[20]/NET0131  & n4584 ;
  assign n8015 = \ctl_rf_c6_rf_prot2_reg/NET0131  & n4577 ;
  assign n8016 = \ctl_rf_c6_rf_chdad_reg[20]/P0002  & n4582 ;
  assign n8017 = ~n8015 & ~n8016 ;
  assign n8018 = ~n8014 & n8017 ;
  assign n8019 = n4611 & ~n8018 ;
  assign n8020 = \ctl_rf_c7_rf_chdad_reg[20]/P0002  & n4582 ;
  assign n8021 = \ctl_rf_c7_rf_chsad_reg[20]/NET0131  & n4584 ;
  assign n8022 = \ctl_rf_c7_rf_prot2_reg/NET0131  & n4577 ;
  assign n8023 = ~n8021 & ~n8022 ;
  assign n8024 = ~n8020 & n8023 ;
  assign n8025 = n4642 & ~n8024 ;
  assign n8026 = ~n8019 & ~n8025 ;
  assign n8027 = \ctl_rf_c5_rf_chsad_reg[20]/NET0131  & n4584 ;
  assign n8028 = \ctl_rf_c5_rf_prot2_reg/NET0131  & n4577 ;
  assign n8029 = \ctl_rf_c5_rf_chdad_reg[20]/P0002  & n4582 ;
  assign n8030 = ~n8028 & ~n8029 ;
  assign n8031 = ~n8027 & n8030 ;
  assign n8032 = n4601 & ~n8031 ;
  assign n8033 = \ctl_rf_c2_rf_chsad_reg[20]/NET0131  & n4584 ;
  assign n8034 = \ctl_rf_c2_rf_prot2_reg/NET0131  & n4577 ;
  assign n8035 = \ctl_rf_c2_rf_chdad_reg[20]/P0002  & n4582 ;
  assign n8036 = ~n8034 & ~n8035 ;
  assign n8037 = ~n8033 & n8036 ;
  assign n8038 = n4590 & ~n8037 ;
  assign n8039 = ~n8032 & ~n8038 ;
  assign n8040 = n8026 & n8039 ;
  assign n8041 = ~n8013 & n8040 ;
  assign n8042 = \ctl_rf_c1_rf_chllp_reg[20]/NET0131  & n4692 ;
  assign n8043 = \ctl_rf_c3_rf_chllp_reg[20]/NET0131  & n4698 ;
  assign n8044 = ~n8042 & ~n8043 ;
  assign n8045 = \ctl_rf_c0_rf_chllp_reg[20]/NET0131  & n4675 ;
  assign n8046 = \ctl_rf_c6_rf_chllp_reg[20]/NET0131  & n4703 ;
  assign n8047 = ~n8045 & ~n8046 ;
  assign n8048 = n8044 & n8047 ;
  assign n8049 = \ctl_rf_c4_rf_chllp_reg[20]/NET0131  & n4687 ;
  assign n8050 = \ctl_rf_c2_rf_chllp_reg[20]/NET0131  & n4663 ;
  assign n8051 = ~n8049 & ~n8050 ;
  assign n8052 = \ctl_rf_c5_rf_chllp_reg[20]/NET0131  & n4680 ;
  assign n8053 = \ctl_rf_c7_rf_chllp_reg[20]/NET0131  & n4669 ;
  assign n8054 = ~n8052 & ~n8053 ;
  assign n8055 = n8051 & n8054 ;
  assign n8056 = n8048 & n8055 ;
  assign n8057 = n4577 & ~n8056 ;
  assign n8058 = \ctl_rf_c0_rf_chdad_reg[20]/P0002  & n4582 ;
  assign n8059 = \ctl_rf_c0_rf_chsad_reg[20]/NET0131  & n4584 ;
  assign n8060 = \ctl_rf_c0_rf_prot2_reg/NET0131  & n4577 ;
  assign n8061 = ~n8059 & ~n8060 ;
  assign n8062 = ~n8058 & n8061 ;
  assign n8063 = n4623 & ~n8062 ;
  assign n8064 = \ctl_rf_c3_rf_chsad_reg[20]/NET0131  & n4584 ;
  assign n8065 = \ctl_rf_c3_rf_prot2_reg/NET0131  & n4577 ;
  assign n8066 = \ctl_rf_c3_rf_chdad_reg[20]/P0002  & n4582 ;
  assign n8067 = ~n8065 & ~n8066 ;
  assign n8068 = ~n8064 & n8067 ;
  assign n8069 = n4651 & ~n8068 ;
  assign n8070 = \ctl_rf_c1_rf_chsad_reg[20]/NET0131  & n4584 ;
  assign n8071 = \ctl_rf_c1_rf_prot2_reg/NET0131  & n4577 ;
  assign n8072 = \ctl_rf_c1_rf_chdad_reg[20]/P0002  & n4582 ;
  assign n8073 = ~n8071 & ~n8072 ;
  assign n8074 = ~n8070 & n8073 ;
  assign n8075 = n4632 & ~n8074 ;
  assign n8076 = ~n8069 & ~n8075 ;
  assign n8077 = ~n8063 & n8076 ;
  assign n8078 = ~n8057 & n8077 ;
  assign n8079 = n8041 & n8078 ;
  assign n8080 = \ctl_rf_c1dmabs_reg[20]/NET0131  & ~\haddr[4]_pad  ;
  assign n8081 = n4579 & n8080 ;
  assign n8082 = \ctl_rf_c3dmabs_reg[20]/NET0131  & ~\haddr[4]_pad  ;
  assign n8083 = n4582 & n8082 ;
  assign n8084 = ~n8081 & ~n8083 ;
  assign n8085 = \ctl_rf_c0dmabs_reg[20]/NET0131  & ~\haddr[4]_pad  ;
  assign n8086 = n4577 & n8085 ;
  assign n8087 = \ctl_rf_c7dmabs_reg[20]/NET0131  & \haddr[4]_pad  ;
  assign n8088 = n4582 & n8087 ;
  assign n8089 = ~n8086 & ~n8088 ;
  assign n8090 = n8084 & n8089 ;
  assign n8091 = \ctl_rf_c6dmabs_reg[20]/NET0131  & \haddr[4]_pad  ;
  assign n8092 = n4584 & n8091 ;
  assign n8093 = \ctl_rf_c4dmabs_reg[20]/NET0131  & \haddr[4]_pad  ;
  assign n8094 = n4577 & n8093 ;
  assign n8095 = ~n8092 & ~n8094 ;
  assign n8096 = \ctl_rf_c2dmabs_reg[20]/NET0131  & ~\haddr[4]_pad  ;
  assign n8097 = n4584 & n8096 ;
  assign n8098 = \ctl_rf_c5dmabs_reg[20]/NET0131  & \haddr[4]_pad  ;
  assign n8099 = n4579 & n8098 ;
  assign n8100 = ~n8097 & ~n8099 ;
  assign n8101 = n8095 & n8100 ;
  assign n8102 = n8090 & n8101 ;
  assign n8103 = n4589 & ~n8102 ;
  assign n8104 = \ctl_rf_c2brbs_reg[20]/NET0131  & ~\haddr[4]_pad  ;
  assign n8105 = n4584 & n8104 ;
  assign n8106 = \ctl_rf_c3brbs_reg[20]/NET0131  & ~\haddr[4]_pad  ;
  assign n8107 = n4582 & n8106 ;
  assign n8108 = ~n8105 & ~n8107 ;
  assign n8109 = \ctl_rf_c0brbs_reg[20]/NET0131  & ~\haddr[4]_pad  ;
  assign n8110 = n4577 & n8109 ;
  assign n8111 = \ctl_rf_c6brbs_reg[20]/NET0131  & \haddr[4]_pad  ;
  assign n8112 = n4584 & n8111 ;
  assign n8113 = ~n8110 & ~n8112 ;
  assign n8114 = n8108 & n8113 ;
  assign n8115 = \ctl_rf_c7brbs_reg[20]/NET0131  & \haddr[4]_pad  ;
  assign n8116 = n4582 & n8115 ;
  assign n8117 = \ctl_rf_c4brbs_reg[20]/NET0131  & \haddr[4]_pad  ;
  assign n8118 = n4577 & n8117 ;
  assign n8119 = ~n8116 & ~n8118 ;
  assign n8120 = \ctl_rf_c1brbs_reg[20]/NET0131  & ~\haddr[4]_pad  ;
  assign n8121 = n4579 & n8120 ;
  assign n8122 = \ctl_rf_c5brbs_reg[20]/NET0131  & \haddr[4]_pad  ;
  assign n8123 = n4579 & n8122 ;
  assign n8124 = ~n8121 & ~n8123 ;
  assign n8125 = n8119 & n8124 ;
  assign n8126 = n8114 & n8125 ;
  assign n8127 = n4575 & ~n8126 ;
  assign n8128 = \ctl_rf_abt_reg[4]/NET0131  & n4622 ;
  assign n8129 = ~\haddr[8]_pad  & ~n8128 ;
  assign n8130 = ~\ctl_rf_c4_rf_int_abt_msk_reg/NET0131  & n5002 ;
  assign n8131 = n5005 & ~n8130 ;
  assign n8132 = ~n8129 & ~n8131 ;
  assign n8133 = ~n8127 & ~n8132 ;
  assign n8134 = ~n8103 & n8133 ;
  assign n8135 = n4569 & ~n8134 ;
  assign n8136 = ~n8079 & n8135 ;
  assign n8137 = ~n7065 & ~n8136 ;
  assign n8138 = ~n8005 & n8137 ;
  assign n8139 = n4745 & n6584 ;
  assign n8140 = n4745 & ~n6641 ;
  assign n8141 = n6625 & n8140 ;
  assign n8142 = ~n8139 & ~n8141 ;
  assign n8143 = ~n4745 & ~n6754 ;
  assign n8144 = ~n6740 & n8143 ;
  assign n8145 = n8142 & ~n8144 ;
  assign n8146 = ~n4573 & ~n8005 ;
  assign n8147 = ~n8145 & n8146 ;
  assign n8148 = ~n8138 & ~n8147 ;
  assign n8149 = \hrdata_reg[5]_pad  & ~n4569 ;
  assign n8150 = \haddr[8]_pad  & ~n4623 ;
  assign n8151 = \ctl_rf_c0_rf_prot3_reg/NET0131  & n4577 ;
  assign n8152 = \ctl_rf_c0_rf_chdad_reg[21]/P0002  & n4582 ;
  assign n8153 = ~n8151 & ~n8152 ;
  assign n8154 = \ctl_rf_c0_rf_chsad_reg[21]/NET0131  & n4584 ;
  assign n8155 = \haddr[8]_pad  & ~n8154 ;
  assign n8156 = n8153 & n8155 ;
  assign n8157 = ~n8150 & ~n8156 ;
  assign n8158 = \ctl_rf_c3_rf_chsad_reg[21]/NET0131  & n4584 ;
  assign n8159 = \ctl_rf_c3_rf_prot3_reg/NET0131  & n4577 ;
  assign n8160 = \ctl_rf_c3_rf_chdad_reg[21]/P0002  & n4582 ;
  assign n8161 = ~n8159 & ~n8160 ;
  assign n8162 = ~n8158 & n8161 ;
  assign n8163 = n4651 & ~n8162 ;
  assign n8164 = \ctl_rf_c5_rf_chdad_reg[21]/P0002  & n4582 ;
  assign n8165 = \ctl_rf_c5_rf_chsad_reg[21]/NET0131  & n4584 ;
  assign n8166 = \ctl_rf_c5_rf_prot3_reg/NET0131  & n4577 ;
  assign n8167 = ~n8165 & ~n8166 ;
  assign n8168 = ~n8164 & n8167 ;
  assign n8169 = n4601 & ~n8168 ;
  assign n8170 = ~n8163 & ~n8169 ;
  assign n8171 = \ctl_rf_c1_rf_chsad_reg[21]/NET0131  & n4584 ;
  assign n8172 = \ctl_rf_c1_rf_prot3_reg/NET0131  & n4577 ;
  assign n8173 = \ctl_rf_c1_rf_chdad_reg[21]/P0002  & n4582 ;
  assign n8174 = ~n8172 & ~n8173 ;
  assign n8175 = ~n8171 & n8174 ;
  assign n8176 = n4632 & ~n8175 ;
  assign n8177 = \ctl_rf_c4_rf_chsad_reg[21]/NET0131  & n4584 ;
  assign n8178 = \ctl_rf_c4_rf_prot3_reg/NET0131  & n4577 ;
  assign n8179 = \ctl_rf_c4_rf_chdad_reg[21]/P0002  & n4582 ;
  assign n8180 = ~n8178 & ~n8179 ;
  assign n8181 = ~n8177 & n8180 ;
  assign n8182 = n4576 & ~n8181 ;
  assign n8183 = ~n8176 & ~n8182 ;
  assign n8184 = n8170 & n8183 ;
  assign n8185 = ~n8157 & n8184 ;
  assign n8186 = \ctl_rf_c4_rf_chllp_reg[21]/NET0131  & n4687 ;
  assign n8187 = \ctl_rf_c2_rf_chllp_reg[21]/NET0131  & n4663 ;
  assign n8188 = ~n8186 & ~n8187 ;
  assign n8189 = \ctl_rf_c3_rf_chllp_reg[21]/NET0131  & n4698 ;
  assign n8190 = \ctl_rf_c1_rf_chllp_reg[21]/NET0131  & n4692 ;
  assign n8191 = ~n8189 & ~n8190 ;
  assign n8192 = n8188 & n8191 ;
  assign n8193 = \ctl_rf_c5_rf_chllp_reg[21]/NET0131  & n4680 ;
  assign n8194 = \ctl_rf_c7_rf_chllp_reg[21]/NET0131  & n4669 ;
  assign n8195 = ~n8193 & ~n8194 ;
  assign n8196 = \ctl_rf_c6_rf_chllp_reg[21]/NET0131  & n4703 ;
  assign n8197 = \ctl_rf_c0_rf_chllp_reg[21]/NET0131  & n4675 ;
  assign n8198 = ~n8196 & ~n8197 ;
  assign n8199 = n8195 & n8198 ;
  assign n8200 = n8192 & n8199 ;
  assign n8201 = n4577 & ~n8200 ;
  assign n8202 = \ctl_rf_c7_rf_chdad_reg[21]/P0002  & n4582 ;
  assign n8203 = \ctl_rf_c7_rf_chsad_reg[21]/NET0131  & n4584 ;
  assign n8204 = \ctl_rf_c7_rf_prot3_reg/NET0131  & n4577 ;
  assign n8205 = ~n8203 & ~n8204 ;
  assign n8206 = ~n8202 & n8205 ;
  assign n8207 = n4642 & ~n8206 ;
  assign n8208 = \ctl_rf_c6_rf_chsad_reg[21]/NET0131  & n4584 ;
  assign n8209 = \ctl_rf_c6_rf_prot3_reg/NET0131  & n4577 ;
  assign n8210 = \ctl_rf_c6_rf_chdad_reg[21]/P0002  & n4582 ;
  assign n8211 = ~n8209 & ~n8210 ;
  assign n8212 = ~n8208 & n8211 ;
  assign n8213 = n4611 & ~n8212 ;
  assign n8214 = \ctl_rf_c2_rf_chsad_reg[21]/NET0131  & n4584 ;
  assign n8215 = \ctl_rf_c2_rf_prot3_reg/NET0131  & n4577 ;
  assign n8216 = \ctl_rf_c2_rf_chdad_reg[21]/P0002  & n4582 ;
  assign n8217 = ~n8215 & ~n8216 ;
  assign n8218 = ~n8214 & n8217 ;
  assign n8219 = n4590 & ~n8218 ;
  assign n8220 = ~n8213 & ~n8219 ;
  assign n8221 = ~n8207 & n8220 ;
  assign n8222 = ~n8201 & n8221 ;
  assign n8223 = n8185 & n8222 ;
  assign n8224 = \ctl_rf_c1brbs_reg[21]/NET0131  & ~\haddr[4]_pad  ;
  assign n8225 = n4579 & n8224 ;
  assign n8226 = \ctl_rf_c3brbs_reg[21]/NET0131  & ~\haddr[4]_pad  ;
  assign n8227 = n4582 & n8226 ;
  assign n8228 = ~n8225 & ~n8227 ;
  assign n8229 = \ctl_rf_c0brbs_reg[21]/NET0131  & ~\haddr[4]_pad  ;
  assign n8230 = n4577 & n8229 ;
  assign n8231 = \ctl_rf_c7brbs_reg[21]/NET0131  & \haddr[4]_pad  ;
  assign n8232 = n4582 & n8231 ;
  assign n8233 = ~n8230 & ~n8232 ;
  assign n8234 = n8228 & n8233 ;
  assign n8235 = \ctl_rf_c6brbs_reg[21]/NET0131  & \haddr[4]_pad  ;
  assign n8236 = n4584 & n8235 ;
  assign n8237 = \ctl_rf_c4brbs_reg[21]/NET0131  & \haddr[4]_pad  ;
  assign n8238 = n4577 & n8237 ;
  assign n8239 = ~n8236 & ~n8238 ;
  assign n8240 = \ctl_rf_c2brbs_reg[21]/NET0131  & ~\haddr[4]_pad  ;
  assign n8241 = n4584 & n8240 ;
  assign n8242 = \ctl_rf_c5brbs_reg[21]/NET0131  & \haddr[4]_pad  ;
  assign n8243 = n4579 & n8242 ;
  assign n8244 = ~n8241 & ~n8243 ;
  assign n8245 = n8239 & n8244 ;
  assign n8246 = n8234 & n8245 ;
  assign n8247 = n4575 & ~n8246 ;
  assign n8248 = \ctl_rf_c2dmabs_reg[21]/NET0131  & ~\haddr[4]_pad  ;
  assign n8249 = n4584 & n8248 ;
  assign n8250 = \ctl_rf_c3dmabs_reg[21]/NET0131  & ~\haddr[4]_pad  ;
  assign n8251 = n4582 & n8250 ;
  assign n8252 = ~n8249 & ~n8251 ;
  assign n8253 = \ctl_rf_c0dmabs_reg[21]/NET0131  & ~\haddr[4]_pad  ;
  assign n8254 = n4577 & n8253 ;
  assign n8255 = \ctl_rf_c6dmabs_reg[21]/NET0131  & \haddr[4]_pad  ;
  assign n8256 = n4584 & n8255 ;
  assign n8257 = ~n8254 & ~n8256 ;
  assign n8258 = n8252 & n8257 ;
  assign n8259 = \ctl_rf_c7dmabs_reg[21]/NET0131  & \haddr[4]_pad  ;
  assign n8260 = n4582 & n8259 ;
  assign n8261 = \ctl_rf_c4dmabs_reg[21]/NET0131  & \haddr[4]_pad  ;
  assign n8262 = n4577 & n8261 ;
  assign n8263 = ~n8260 & ~n8262 ;
  assign n8264 = \ctl_rf_c1dmabs_reg[21]/NET0131  & ~\haddr[4]_pad  ;
  assign n8265 = n4579 & n8264 ;
  assign n8266 = \ctl_rf_c5dmabs_reg[21]/NET0131  & \haddr[4]_pad  ;
  assign n8267 = n4579 & n8266 ;
  assign n8268 = ~n8265 & ~n8267 ;
  assign n8269 = n8263 & n8268 ;
  assign n8270 = n8258 & n8269 ;
  assign n8271 = n4589 & ~n8270 ;
  assign n8272 = \ctl_rf_abt_reg[5]/NET0131  & n4622 ;
  assign n8273 = ~\haddr[8]_pad  & ~n8272 ;
  assign n8274 = ~\ctl_rf_c5_rf_int_abt_msk_reg/NET0131  & n5002 ;
  assign n8275 = n5005 & ~n8274 ;
  assign n8276 = ~n8273 & ~n8275 ;
  assign n8277 = ~n8271 & ~n8276 ;
  assign n8278 = ~n8247 & n8277 ;
  assign n8279 = n4569 & ~n8278 ;
  assign n8280 = ~n8223 & n8279 ;
  assign n8281 = ~n7065 & ~n8280 ;
  assign n8282 = ~n8149 & n8281 ;
  assign n8283 = n4745 & n6887 ;
  assign n8284 = n4745 & ~n6944 ;
  assign n8285 = n6928 & n8284 ;
  assign n8286 = ~n8283 & ~n8285 ;
  assign n8287 = ~n4745 & ~n7057 ;
  assign n8288 = ~n7043 & n8287 ;
  assign n8289 = n8286 & ~n8288 ;
  assign n8290 = ~n4573 & ~n8149 ;
  assign n8291 = ~n8289 & n8290 ;
  assign n8292 = ~n8282 & ~n8291 ;
  assign n8293 = \hrdata_reg[6]_pad  & ~n4569 ;
  assign n8294 = \haddr[8]_pad  & ~n4642 ;
  assign n8295 = \ctl_rf_c7_rf_chpri_reg[0]/NET0131  & n4577 ;
  assign n8296 = \ctl_rf_c7_rf_chdad_reg[22]/P0002  & n4582 ;
  assign n8297 = ~n8295 & ~n8296 ;
  assign n8298 = \ctl_rf_c7_rf_chsad_reg[22]/NET0131  & n4584 ;
  assign n8299 = \haddr[8]_pad  & ~n8298 ;
  assign n8300 = n8297 & n8299 ;
  assign n8301 = ~n8294 & ~n8300 ;
  assign n8302 = \ctl_rf_c6_rf_chsad_reg[22]/NET0131  & n4584 ;
  assign n8303 = \ctl_rf_c6_rf_chpri_reg[0]/NET0131  & n4577 ;
  assign n8304 = \ctl_rf_c6_rf_chdad_reg[22]/P0002  & n4582 ;
  assign n8305 = ~n8303 & ~n8304 ;
  assign n8306 = ~n8302 & n8305 ;
  assign n8307 = n4611 & ~n8306 ;
  assign n8308 = \ctl_rf_c4_rf_chdad_reg[22]/P0002  & n4582 ;
  assign n8309 = \ctl_rf_c4_rf_chsad_reg[22]/NET0131  & n4584 ;
  assign n8310 = \ctl_rf_c4_rf_chpri_reg[0]/NET0131  & n4577 ;
  assign n8311 = ~n8309 & ~n8310 ;
  assign n8312 = ~n8308 & n8311 ;
  assign n8313 = n4576 & ~n8312 ;
  assign n8314 = ~n8307 & ~n8313 ;
  assign n8315 = \ctl_rf_c0_rf_chsad_reg[22]/NET0131  & n4584 ;
  assign n8316 = \ctl_rf_c0_rf_chpri_reg[0]/NET0131  & n4577 ;
  assign n8317 = \ctl_rf_c0_rf_chdad_reg[22]/P0002  & n4582 ;
  assign n8318 = ~n8316 & ~n8317 ;
  assign n8319 = ~n8315 & n8318 ;
  assign n8320 = n4623 & ~n8319 ;
  assign n8321 = \ctl_rf_c3_rf_chsad_reg[22]/NET0131  & n4584 ;
  assign n8322 = \ctl_rf_c3_rf_chpri_reg[0]/NET0131  & n4577 ;
  assign n8323 = \ctl_rf_c3_rf_chdad_reg[22]/P0002  & n4582 ;
  assign n8324 = ~n8322 & ~n8323 ;
  assign n8325 = ~n8321 & n8324 ;
  assign n8326 = n4651 & ~n8325 ;
  assign n8327 = ~n8320 & ~n8326 ;
  assign n8328 = n8314 & n8327 ;
  assign n8329 = ~n8301 & n8328 ;
  assign n8330 = \ctl_rf_c1_rf_chllp_reg[22]/NET0131  & n4692 ;
  assign n8331 = \ctl_rf_c3_rf_chllp_reg[22]/NET0131  & n4698 ;
  assign n8332 = ~n8330 & ~n8331 ;
  assign n8333 = \ctl_rf_c0_rf_chllp_reg[22]/NET0131  & n4675 ;
  assign n8334 = \ctl_rf_c6_rf_chllp_reg[22]/NET0131  & n4703 ;
  assign n8335 = ~n8333 & ~n8334 ;
  assign n8336 = n8332 & n8335 ;
  assign n8337 = \ctl_rf_c4_rf_chllp_reg[22]/NET0131  & n4687 ;
  assign n8338 = \ctl_rf_c2_rf_chllp_reg[22]/NET0131  & n4663 ;
  assign n8339 = ~n8337 & ~n8338 ;
  assign n8340 = \ctl_rf_c5_rf_chllp_reg[22]/NET0131  & n4680 ;
  assign n8341 = \ctl_rf_c7_rf_chllp_reg[22]/NET0131  & n4669 ;
  assign n8342 = ~n8340 & ~n8341 ;
  assign n8343 = n8339 & n8342 ;
  assign n8344 = n8336 & n8343 ;
  assign n8345 = n4577 & ~n8344 ;
  assign n8346 = \ctl_rf_c5_rf_chdad_reg[22]/P0002  & n4582 ;
  assign n8347 = \ctl_rf_c5_rf_chsad_reg[22]/NET0131  & n4584 ;
  assign n8348 = \ctl_rf_c5_rf_chpri_reg[0]/NET0131  & n4577 ;
  assign n8349 = ~n8347 & ~n8348 ;
  assign n8350 = ~n8346 & n8349 ;
  assign n8351 = n4601 & ~n8350 ;
  assign n8352 = \ctl_rf_c2_rf_chsad_reg[22]/NET0131  & n4584 ;
  assign n8353 = \ctl_rf_c2_rf_chpri_reg[0]/NET0131  & n4577 ;
  assign n8354 = \ctl_rf_c2_rf_chdad_reg[22]/P0002  & n4582 ;
  assign n8355 = ~n8353 & ~n8354 ;
  assign n8356 = ~n8352 & n8355 ;
  assign n8357 = n4590 & ~n8356 ;
  assign n8358 = \ctl_rf_c1_rf_chsad_reg[22]/NET0131  & n4584 ;
  assign n8359 = \ctl_rf_c1_rf_chpri_reg[0]/NET0131  & n4577 ;
  assign n8360 = \ctl_rf_c1_rf_chdad_reg[22]/P0002  & n4582 ;
  assign n8361 = ~n8359 & ~n8360 ;
  assign n8362 = ~n8358 & n8361 ;
  assign n8363 = n4632 & ~n8362 ;
  assign n8364 = ~n8357 & ~n8363 ;
  assign n8365 = ~n8351 & n8364 ;
  assign n8366 = ~n8345 & n8365 ;
  assign n8367 = n8329 & n8366 ;
  assign n8368 = \ctl_rf_c1brbs_reg[22]/NET0131  & ~\haddr[4]_pad  ;
  assign n8369 = n4579 & n8368 ;
  assign n8370 = \ctl_rf_c3brbs_reg[22]/NET0131  & ~\haddr[4]_pad  ;
  assign n8371 = n4582 & n8370 ;
  assign n8372 = ~n8369 & ~n8371 ;
  assign n8373 = \ctl_rf_c0brbs_reg[22]/NET0131  & ~\haddr[4]_pad  ;
  assign n8374 = n4577 & n8373 ;
  assign n8375 = \ctl_rf_c7brbs_reg[22]/NET0131  & \haddr[4]_pad  ;
  assign n8376 = n4582 & n8375 ;
  assign n8377 = ~n8374 & ~n8376 ;
  assign n8378 = n8372 & n8377 ;
  assign n8379 = \ctl_rf_c6brbs_reg[22]/NET0131  & \haddr[4]_pad  ;
  assign n8380 = n4584 & n8379 ;
  assign n8381 = \ctl_rf_c4brbs_reg[22]/NET0131  & \haddr[4]_pad  ;
  assign n8382 = n4577 & n8381 ;
  assign n8383 = ~n8380 & ~n8382 ;
  assign n8384 = \ctl_rf_c2brbs_reg[22]/NET0131  & ~\haddr[4]_pad  ;
  assign n8385 = n4584 & n8384 ;
  assign n8386 = \ctl_rf_c5brbs_reg[22]/NET0131  & \haddr[4]_pad  ;
  assign n8387 = n4579 & n8386 ;
  assign n8388 = ~n8385 & ~n8387 ;
  assign n8389 = n8383 & n8388 ;
  assign n8390 = n8378 & n8389 ;
  assign n8391 = n4575 & ~n8390 ;
  assign n8392 = \ctl_rf_c2dmabs_reg[22]/NET0131  & ~\haddr[4]_pad  ;
  assign n8393 = n4584 & n8392 ;
  assign n8394 = \ctl_rf_c3dmabs_reg[22]/NET0131  & ~\haddr[4]_pad  ;
  assign n8395 = n4582 & n8394 ;
  assign n8396 = ~n8393 & ~n8395 ;
  assign n8397 = \ctl_rf_c0dmabs_reg[22]/NET0131  & ~\haddr[4]_pad  ;
  assign n8398 = n4577 & n8397 ;
  assign n8399 = \ctl_rf_c6dmabs_reg[22]/NET0131  & \haddr[4]_pad  ;
  assign n8400 = n4584 & n8399 ;
  assign n8401 = ~n8398 & ~n8400 ;
  assign n8402 = n8396 & n8401 ;
  assign n8403 = \ctl_rf_c7dmabs_reg[22]/NET0131  & \haddr[4]_pad  ;
  assign n8404 = n4582 & n8403 ;
  assign n8405 = \ctl_rf_c4dmabs_reg[22]/NET0131  & \haddr[4]_pad  ;
  assign n8406 = n4577 & n8405 ;
  assign n8407 = ~n8404 & ~n8406 ;
  assign n8408 = \ctl_rf_c1dmabs_reg[22]/NET0131  & ~\haddr[4]_pad  ;
  assign n8409 = n4579 & n8408 ;
  assign n8410 = \ctl_rf_c5dmabs_reg[22]/NET0131  & \haddr[4]_pad  ;
  assign n8411 = n4579 & n8410 ;
  assign n8412 = ~n8409 & ~n8411 ;
  assign n8413 = n8407 & n8412 ;
  assign n8414 = n8402 & n8413 ;
  assign n8415 = n4589 & ~n8414 ;
  assign n8416 = \ctl_rf_abt_reg[6]/NET0131  & n4622 ;
  assign n8417 = ~\haddr[8]_pad  & ~n8416 ;
  assign n8418 = ~\ctl_rf_c6_rf_int_abt_msk_reg/NET0131  & n5002 ;
  assign n8419 = n5005 & ~n8418 ;
  assign n8420 = ~n8417 & ~n8419 ;
  assign n8421 = ~n8415 & ~n8420 ;
  assign n8422 = ~n8391 & n8421 ;
  assign n8423 = n4569 & ~n8422 ;
  assign n8424 = ~n8367 & n8423 ;
  assign n8425 = ~n7065 & ~n8424 ;
  assign n8426 = ~n8293 & n8425 ;
  assign n8427 = n4745 & n7350 ;
  assign n8428 = n4745 & ~n7407 ;
  assign n8429 = n7391 & n8428 ;
  assign n8430 = ~n8427 & ~n8429 ;
  assign n8431 = ~n4745 & ~n7520 ;
  assign n8432 = ~n7506 & n8431 ;
  assign n8433 = n8430 & ~n8432 ;
  assign n8434 = ~n4573 & ~n8293 ;
  assign n8435 = ~n8433 & n8434 ;
  assign n8436 = ~n8426 & ~n8435 ;
  assign n8437 = \hrdata_reg[7]_pad  & ~n4569 ;
  assign n8438 = \ctl_rf_c4_rf_chpri_reg[1]/NET0131  & n4577 ;
  assign n8439 = \ctl_rf_c4_rf_chdad_reg[23]/P0002  & n4582 ;
  assign n8440 = ~n8438 & ~n8439 ;
  assign n8441 = \ctl_rf_c4_rf_chsad_reg[23]/NET0131  & n4584 ;
  assign n8442 = \haddr[8]_pad  & ~n8441 ;
  assign n8443 = n8440 & n8442 ;
  assign n8444 = ~n8006 & ~n8443 ;
  assign n8445 = \ctl_rf_c1_rf_chsad_reg[23]/NET0131  & n4584 ;
  assign n8446 = \ctl_rf_c1_rf_chpri_reg[1]/NET0131  & n4577 ;
  assign n8447 = \ctl_rf_c1_rf_chdad_reg[23]/P0002  & n4582 ;
  assign n8448 = ~n8446 & ~n8447 ;
  assign n8449 = ~n8445 & n8448 ;
  assign n8450 = n4632 & ~n8449 ;
  assign n8451 = \ctl_rf_c6_rf_chdad_reg[23]/P0002  & n4582 ;
  assign n8452 = \ctl_rf_c6_rf_chsad_reg[23]/NET0131  & n4584 ;
  assign n8453 = \ctl_rf_c6_rf_chpri_reg[1]/NET0131  & n4577 ;
  assign n8454 = ~n8452 & ~n8453 ;
  assign n8455 = ~n8451 & n8454 ;
  assign n8456 = n4611 & ~n8455 ;
  assign n8457 = ~n8450 & ~n8456 ;
  assign n8458 = \ctl_rf_c0_rf_chsad_reg[23]/NET0131  & n4584 ;
  assign n8459 = \ctl_rf_c0_rf_chpri_reg[1]/NET0131  & n4577 ;
  assign n8460 = \ctl_rf_c0_rf_chdad_reg[23]/P0002  & n4582 ;
  assign n8461 = ~n8459 & ~n8460 ;
  assign n8462 = ~n8458 & n8461 ;
  assign n8463 = n4623 & ~n8462 ;
  assign n8464 = \ctl_rf_c2_rf_chsad_reg[23]/NET0131  & n4584 ;
  assign n8465 = \ctl_rf_c2_rf_chpri_reg[1]/NET0131  & n4577 ;
  assign n8466 = \ctl_rf_c2_rf_chdad_reg[23]/P0002  & n4582 ;
  assign n8467 = ~n8465 & ~n8466 ;
  assign n8468 = ~n8464 & n8467 ;
  assign n8469 = n4590 & ~n8468 ;
  assign n8470 = ~n8463 & ~n8469 ;
  assign n8471 = n8457 & n8470 ;
  assign n8472 = ~n8444 & n8471 ;
  assign n8473 = \ctl_rf_c5_rf_chllp_reg[23]/NET0131  & n4680 ;
  assign n8474 = \ctl_rf_c0_rf_chllp_reg[23]/NET0131  & n4675 ;
  assign n8475 = ~n8473 & ~n8474 ;
  assign n8476 = \ctl_rf_c2_rf_chllp_reg[23]/NET0131  & n4663 ;
  assign n8477 = \ctl_rf_c6_rf_chllp_reg[23]/NET0131  & n4703 ;
  assign n8478 = ~n8476 & ~n8477 ;
  assign n8479 = n8475 & n8478 ;
  assign n8480 = \ctl_rf_c1_rf_chllp_reg[23]/NET0131  & n4692 ;
  assign n8481 = \ctl_rf_c3_rf_chllp_reg[23]/NET0131  & n4698 ;
  assign n8482 = ~n8480 & ~n8481 ;
  assign n8483 = \ctl_rf_c4_rf_chllp_reg[23]/NET0131  & n4687 ;
  assign n8484 = \ctl_rf_c7_rf_chllp_reg[23]/NET0131  & n4669 ;
  assign n8485 = ~n8483 & ~n8484 ;
  assign n8486 = n8482 & n8485 ;
  assign n8487 = n8479 & n8486 ;
  assign n8488 = n4577 & ~n8487 ;
  assign n8489 = \ctl_rf_c5_rf_chdad_reg[23]/P0002  & n4582 ;
  assign n8490 = \ctl_rf_c5_rf_chsad_reg[23]/NET0131  & n4584 ;
  assign n8491 = \ctl_rf_c5_rf_chpri_reg[1]/NET0131  & n4577 ;
  assign n8492 = ~n8490 & ~n8491 ;
  assign n8493 = ~n8489 & n8492 ;
  assign n8494 = n4601 & ~n8493 ;
  assign n8495 = \ctl_rf_c3_rf_chsad_reg[23]/NET0131  & n4584 ;
  assign n8496 = \ctl_rf_c3_rf_chpri_reg[1]/NET0131  & n4577 ;
  assign n8497 = \ctl_rf_c3_rf_chdad_reg[23]/P0002  & n4582 ;
  assign n8498 = ~n8496 & ~n8497 ;
  assign n8499 = ~n8495 & n8498 ;
  assign n8500 = n4651 & ~n8499 ;
  assign n8501 = \ctl_rf_c7_rf_chsad_reg[23]/NET0131  & n4584 ;
  assign n8502 = \ctl_rf_c7_rf_chpri_reg[1]/NET0131  & n4577 ;
  assign n8503 = \ctl_rf_c7_rf_chdad_reg[23]/P0002  & n4582 ;
  assign n8504 = ~n8502 & ~n8503 ;
  assign n8505 = ~n8501 & n8504 ;
  assign n8506 = n4642 & ~n8505 ;
  assign n8507 = ~n8500 & ~n8506 ;
  assign n8508 = ~n8494 & n8507 ;
  assign n8509 = ~n8488 & n8508 ;
  assign n8510 = n8472 & n8509 ;
  assign n8511 = \ctl_rf_c1brbs_reg[23]/NET0131  & ~\haddr[4]_pad  ;
  assign n8512 = n4579 & n8511 ;
  assign n8513 = \ctl_rf_c3brbs_reg[23]/NET0131  & ~\haddr[4]_pad  ;
  assign n8514 = n4582 & n8513 ;
  assign n8515 = ~n8512 & ~n8514 ;
  assign n8516 = \ctl_rf_c0brbs_reg[23]/NET0131  & ~\haddr[4]_pad  ;
  assign n8517 = n4577 & n8516 ;
  assign n8518 = \ctl_rf_c7brbs_reg[23]/NET0131  & \haddr[4]_pad  ;
  assign n8519 = n4582 & n8518 ;
  assign n8520 = ~n8517 & ~n8519 ;
  assign n8521 = n8515 & n8520 ;
  assign n8522 = \ctl_rf_c6brbs_reg[23]/NET0131  & \haddr[4]_pad  ;
  assign n8523 = n4584 & n8522 ;
  assign n8524 = \ctl_rf_c4brbs_reg[23]/NET0131  & \haddr[4]_pad  ;
  assign n8525 = n4577 & n8524 ;
  assign n8526 = ~n8523 & ~n8525 ;
  assign n8527 = \ctl_rf_c2brbs_reg[23]/NET0131  & ~\haddr[4]_pad  ;
  assign n8528 = n4584 & n8527 ;
  assign n8529 = \ctl_rf_c5brbs_reg[23]/NET0131  & \haddr[4]_pad  ;
  assign n8530 = n4579 & n8529 ;
  assign n8531 = ~n8528 & ~n8530 ;
  assign n8532 = n8526 & n8531 ;
  assign n8533 = n8521 & n8532 ;
  assign n8534 = n4575 & ~n8533 ;
  assign n8535 = \ctl_rf_c2dmabs_reg[23]/NET0131  & ~\haddr[4]_pad  ;
  assign n8536 = n4584 & n8535 ;
  assign n8537 = \ctl_rf_c3dmabs_reg[23]/NET0131  & ~\haddr[4]_pad  ;
  assign n8538 = n4582 & n8537 ;
  assign n8539 = ~n8536 & ~n8538 ;
  assign n8540 = \ctl_rf_c0dmabs_reg[23]/NET0131  & ~\haddr[4]_pad  ;
  assign n8541 = n4577 & n8540 ;
  assign n8542 = \ctl_rf_c6dmabs_reg[23]/NET0131  & \haddr[4]_pad  ;
  assign n8543 = n4584 & n8542 ;
  assign n8544 = ~n8541 & ~n8543 ;
  assign n8545 = n8539 & n8544 ;
  assign n8546 = \ctl_rf_c7dmabs_reg[23]/NET0131  & \haddr[4]_pad  ;
  assign n8547 = n4582 & n8546 ;
  assign n8548 = \ctl_rf_c4dmabs_reg[23]/NET0131  & \haddr[4]_pad  ;
  assign n8549 = n4577 & n8548 ;
  assign n8550 = ~n8547 & ~n8549 ;
  assign n8551 = \ctl_rf_c1dmabs_reg[23]/NET0131  & ~\haddr[4]_pad  ;
  assign n8552 = n4579 & n8551 ;
  assign n8553 = \ctl_rf_c5dmabs_reg[23]/NET0131  & \haddr[4]_pad  ;
  assign n8554 = n4579 & n8553 ;
  assign n8555 = ~n8552 & ~n8554 ;
  assign n8556 = n8550 & n8555 ;
  assign n8557 = n8545 & n8556 ;
  assign n8558 = n4589 & ~n8557 ;
  assign n8559 = \ctl_rf_abt_reg[7]/NET0131  & n4622 ;
  assign n8560 = ~\haddr[8]_pad  & ~n8559 ;
  assign n8561 = ~\ctl_rf_c7_rf_int_abt_msk_reg/NET0131  & n5002 ;
  assign n8562 = n5005 & ~n8561 ;
  assign n8563 = ~n8560 & ~n8562 ;
  assign n8564 = ~n8558 & ~n8563 ;
  assign n8565 = ~n8534 & n8564 ;
  assign n8566 = n4569 & ~n8565 ;
  assign n8567 = ~n8510 & n8566 ;
  assign n8568 = ~n7065 & ~n8567 ;
  assign n8569 = ~n8437 & n8568 ;
  assign n8570 = n4745 & ~n7728 ;
  assign n8571 = ~n4745 & ~n7839 ;
  assign n8572 = ~n7825 & n8571 ;
  assign n8573 = ~n8570 & ~n8572 ;
  assign n8574 = ~n4573 & ~n8437 ;
  assign n8575 = ~n8573 & n8574 ;
  assign n8576 = ~n8569 & ~n8575 ;
  assign n8577 = ~\ahb_slv_slv_ad_d1o_reg[3]/NET0131  & \ahb_slv_slv_ad_d1o_reg[4]/NET0131  ;
  assign n8578 = n2229 & n8577 ;
  assign n8579 = n2232 & n2251 ;
  assign n8580 = \ctl_rf_be_d1_reg[0]/P0001  & n8579 ;
  assign n8581 = n8578 & n8580 ;
  assign n8582 = ~\ctl_rf_c1_rf_chtsz_reg[5]/NET0131  & ~n8581 ;
  assign n8583 = \hwdata[5]_pad  & ~n2242 ;
  assign n8584 = \hwdata[29]_pad  & n2242 ;
  assign n8585 = ~n8583 & ~n8584 ;
  assign n8586 = ~n2240 & ~n8585 ;
  assign n8587 = \hwdata[21]_pad  & n2240 ;
  assign n8588 = n8581 & ~n8587 ;
  assign n8589 = ~n8586 & n8588 ;
  assign n8590 = ~n8582 & ~n8589 ;
  assign n8591 = ~\ctl_rf_c1_rf_chtsz_reg[6]/NET0131  & ~n8581 ;
  assign n8592 = \hwdata[6]_pad  & ~n2242 ;
  assign n8593 = \hwdata[30]_pad  & n2242 ;
  assign n8594 = ~n8592 & ~n8593 ;
  assign n8595 = ~n2240 & ~n8594 ;
  assign n8596 = \hwdata[22]_pad  & n2240 ;
  assign n8597 = n8581 & ~n8596 ;
  assign n8598 = ~n8595 & n8597 ;
  assign n8599 = ~n8591 & ~n8598 ;
  assign n8600 = ~\ctl_rf_c1_rf_chtsz_reg[7]/NET0131  & ~n8581 ;
  assign n8601 = ~n2247 & n8581 ;
  assign n8602 = ~n2246 & n8601 ;
  assign n8603 = ~n8600 & ~n8602 ;
  assign n8604 = n2235 & n2311 ;
  assign n8605 = ~\ctl_rf_c3_rf_chsad_reg[7]/NET0131  & ~n8604 ;
  assign n8606 = ~n2247 & n8604 ;
  assign n8607 = ~n2246 & n8606 ;
  assign n8608 = ~n8605 & ~n8607 ;
  assign n8609 = n2265 & n8577 ;
  assign n8610 = n8580 & n8609 ;
  assign n8611 = ~\ctl_rf_c3_rf_chtsz_reg[5]/NET0131  & ~n8610 ;
  assign n8612 = ~n8587 & n8610 ;
  assign n8613 = ~n8586 & n8612 ;
  assign n8614 = ~n8611 & ~n8613 ;
  assign n8615 = ~\ctl_rf_c3_rf_chtsz_reg[6]/NET0131  & ~n8610 ;
  assign n8616 = ~n8596 & n8610 ;
  assign n8617 = ~n8595 & n8616 ;
  assign n8618 = ~n8615 & ~n8617 ;
  assign n8619 = ~\ctl_rf_c3_rf_chtsz_reg[7]/NET0131  & ~n8610 ;
  assign n8620 = ~n2247 & n8610 ;
  assign n8621 = ~n2246 & n8620 ;
  assign n8622 = ~n8619 & ~n8621 ;
  assign n8623 = \ctl_rf_be_d1_reg[0]/P0001  & n2276 ;
  assign n8624 = n2317 & n8623 ;
  assign n8625 = ~\ctl_rf_c4_rf_chsad_reg[7]/NET0131  & ~n8624 ;
  assign n8626 = ~n2247 & n8624 ;
  assign n8627 = ~n2246 & n8626 ;
  assign n8628 = ~n8625 & ~n8627 ;
  assign n8629 = n2273 & n8577 ;
  assign n8630 = n2251 & n2275 ;
  assign n8631 = \ctl_rf_be_d1_reg[0]/P0001  & n8630 ;
  assign n8632 = n8629 & n8631 ;
  assign n8633 = ~\ctl_rf_c4_rf_chtsz_reg[5]/NET0131  & ~n8632 ;
  assign n8634 = ~n8587 & n8632 ;
  assign n8635 = ~n8586 & n8634 ;
  assign n8636 = ~n8633 & ~n8635 ;
  assign n8637 = ~\ctl_rf_c4_rf_chtsz_reg[6]/NET0131  & ~n8632 ;
  assign n8638 = ~n8596 & n8632 ;
  assign n8639 = ~n8595 & n8638 ;
  assign n8640 = ~n8637 & ~n8639 ;
  assign n8641 = n2235 & n2317 ;
  assign n8642 = ~\ctl_rf_c5_rf_chsad_reg[7]/NET0131  & ~n8641 ;
  assign n8643 = ~n2247 & n8641 ;
  assign n8644 = ~n2246 & n8643 ;
  assign n8645 = ~n8642 & ~n8644 ;
  assign n8646 = n8580 & n8629 ;
  assign n8647 = ~\ctl_rf_c5_rf_chtsz_reg[6]/NET0131  & ~n8646 ;
  assign n8648 = ~n8596 & n8646 ;
  assign n8649 = ~n8595 & n8648 ;
  assign n8650 = ~n8647 & ~n8649 ;
  assign n8651 = n2324 & n8623 ;
  assign n8652 = ~\ctl_rf_c6_rf_chsad_reg[7]/NET0131  & ~n8651 ;
  assign n8653 = ~n2247 & n8651 ;
  assign n8654 = ~n2246 & n8653 ;
  assign n8655 = ~n8652 & ~n8654 ;
  assign n8656 = n2275 & n2288 ;
  assign n8657 = n2251 & n8577 ;
  assign n8658 = \ctl_rf_be_d1_reg[0]/P0001  & n8657 ;
  assign n8659 = n8656 & n8658 ;
  assign n8660 = ~\ctl_rf_c6_rf_chtsz_reg[5]/NET0131  & ~n8659 ;
  assign n8661 = ~n8587 & n8659 ;
  assign n8662 = ~n8586 & n8661 ;
  assign n8663 = ~n8660 & ~n8662 ;
  assign n8664 = ~\ctl_rf_c6_rf_chtsz_reg[6]/NET0131  & ~n8659 ;
  assign n8665 = ~n8596 & n8659 ;
  assign n8666 = ~n8595 & n8665 ;
  assign n8667 = ~n8664 & ~n8666 ;
  assign n8668 = ~\ctl_rf_c6_rf_chtsz_reg[7]/NET0131  & ~n8659 ;
  assign n8669 = ~n2247 & n8659 ;
  assign n8670 = ~n2246 & n8669 ;
  assign n8671 = ~n8668 & ~n8670 ;
  assign n8672 = n2235 & n2324 ;
  assign n8673 = ~\ctl_rf_c7_rf_chsad_reg[7]/NET0131  & ~n8672 ;
  assign n8674 = ~n2247 & n8672 ;
  assign n8675 = ~n2246 & n8674 ;
  assign n8676 = ~n8673 & ~n8675 ;
  assign n8677 = n2232 & n2288 ;
  assign n8678 = n8658 & n8677 ;
  assign n8679 = ~\ctl_rf_c7_rf_chtsz_reg[5]/NET0131  & ~n8678 ;
  assign n8680 = ~n8587 & n8678 ;
  assign n8681 = ~n8586 & n8680 ;
  assign n8682 = ~n8679 & ~n8681 ;
  assign n8683 = ~\ctl_rf_c7_rf_chtsz_reg[6]/NET0131  & ~n8678 ;
  assign n8684 = ~n8596 & n8678 ;
  assign n8685 = ~n8595 & n8684 ;
  assign n8686 = ~n8683 & ~n8685 ;
  assign n8687 = ~\ctl_rf_c7_rf_chtsz_reg[7]/NET0131  & ~n8678 ;
  assign n8688 = ~n2247 & n8678 ;
  assign n8689 = ~n2246 & n8688 ;
  assign n8690 = ~n8687 & ~n8689 ;
  assign n8691 = n2231 & n8623 ;
  assign n8692 = ~\ctl_rf_c0_rf_chsad_reg[7]/NET0131  & ~n8691 ;
  assign n8693 = ~n2247 & n8691 ;
  assign n8694 = ~n2246 & n8693 ;
  assign n8695 = ~n8692 & ~n8694 ;
  assign n8696 = n8578 & n8631 ;
  assign n8697 = ~\ctl_rf_c0_rf_chtsz_reg[5]/NET0131  & ~n8696 ;
  assign n8698 = ~n8587 & n8696 ;
  assign n8699 = ~n8586 & n8698 ;
  assign n8700 = ~n8697 & ~n8699 ;
  assign n8701 = ~\ctl_rf_c0_rf_chtsz_reg[6]/NET0131  & ~n8696 ;
  assign n8702 = ~n8596 & n8696 ;
  assign n8703 = ~n8595 & n8702 ;
  assign n8704 = ~n8701 & ~n8703 ;
  assign n8705 = ~\ctl_rf_c0_rf_chtsz_reg[7]/NET0131  & ~n8696 ;
  assign n8706 = ~n2247 & n8696 ;
  assign n8707 = ~n2246 & n8706 ;
  assign n8708 = ~n8705 & ~n8707 ;
  assign n8709 = ~\ctl_rf_c1_rf_chtsz_reg[4]/NET0131  & ~n8581 ;
  assign n8710 = \hwdata[4]_pad  & ~n2242 ;
  assign n8711 = \hwdata[28]_pad  & n2242 ;
  assign n8712 = ~n8710 & ~n8711 ;
  assign n8713 = ~n2240 & ~n8712 ;
  assign n8714 = \hwdata[20]_pad  & n2240 ;
  assign n8715 = n8581 & ~n8714 ;
  assign n8716 = ~n8713 & n8715 ;
  assign n8717 = ~n8709 & ~n8716 ;
  assign n8718 = n2311 & n8623 ;
  assign n8719 = ~\ctl_rf_c2_rf_chsad_reg[7]/NET0131  & ~n8718 ;
  assign n8720 = ~n2247 & n8718 ;
  assign n8721 = ~n2246 & n8720 ;
  assign n8722 = ~n8719 & ~n8721 ;
  assign n8723 = n8609 & n8631 ;
  assign n8724 = ~\ctl_rf_c2_rf_chtsz_reg[5]/NET0131  & ~n8723 ;
  assign n8725 = ~n8587 & n8723 ;
  assign n8726 = ~n8586 & n8725 ;
  assign n8727 = ~n8724 & ~n8726 ;
  assign n8728 = ~\ctl_rf_c2_rf_chtsz_reg[6]/NET0131  & ~n8723 ;
  assign n8729 = ~n8596 & n8723 ;
  assign n8730 = ~n8595 & n8729 ;
  assign n8731 = ~n8728 & ~n8730 ;
  assign n8732 = ~\ctl_rf_c2_rf_chtsz_reg[7]/NET0131  & ~n8723 ;
  assign n8733 = ~n2247 & n8723 ;
  assign n8734 = ~n2246 & n8733 ;
  assign n8735 = ~n8732 & ~n8734 ;
  assign n8736 = ~\ctl_rf_c3_rf_chtsz_reg[4]/NET0131  & ~n8610 ;
  assign n8737 = n8610 & ~n8714 ;
  assign n8738 = ~n8713 & n8737 ;
  assign n8739 = ~n8736 & ~n8738 ;
  assign n8740 = ~\ctl_rf_c4_rf_chtsz_reg[4]/NET0131  & ~n8632 ;
  assign n8741 = n8632 & ~n8714 ;
  assign n8742 = ~n8713 & n8741 ;
  assign n8743 = ~n8740 & ~n8742 ;
  assign n8744 = ~\ctl_rf_c6_rf_chtsz_reg[4]/NET0131  & ~n8659 ;
  assign n8745 = n8659 & ~n8714 ;
  assign n8746 = ~n8713 & n8745 ;
  assign n8747 = ~n8744 & ~n8746 ;
  assign n8748 = ~\ctl_rf_c7_rf_chtsz_reg[4]/NET0131  & ~n8678 ;
  assign n8749 = n8678 & ~n8714 ;
  assign n8750 = ~n8713 & n8749 ;
  assign n8751 = ~n8748 & ~n8750 ;
  assign n8752 = \ctl_rf_be_d1_reg[1]/P0001  & n2234 ;
  assign n8753 = n2252 & n8752 ;
  assign n8754 = ~\ctl_rf_c1_rf_chdad_reg[10]/NET0131  & ~n8753 ;
  assign n8755 = \hwdata[10]_pad  & ~n2242 ;
  assign n8756 = \hwdata[18]_pad  & n2242 ;
  assign n8757 = ~n8755 & ~n8756 ;
  assign n8758 = ~n2240 & ~n8757 ;
  assign n8759 = \hwdata[26]_pad  & n2240 ;
  assign n8760 = n8753 & ~n8759 ;
  assign n8761 = ~n8758 & n8760 ;
  assign n8762 = ~n8754 & ~n8761 ;
  assign n8763 = ~\ctl_rf_c1_rf_chdad_reg[12]/NET0131  & ~n8753 ;
  assign n8764 = \hwdata[12]_pad  & ~n2242 ;
  assign n8765 = \hwdata[20]_pad  & n2242 ;
  assign n8766 = ~n8764 & ~n8765 ;
  assign n8767 = ~n2240 & ~n8766 ;
  assign n8768 = \hwdata[28]_pad  & n2240 ;
  assign n8769 = n8753 & ~n8768 ;
  assign n8770 = ~n8767 & n8769 ;
  assign n8771 = ~n8763 & ~n8770 ;
  assign n8772 = ~\ctl_rf_c1_rf_chdad_reg[15]/NET0131  & ~n8753 ;
  assign n8773 = ~n3763 & n8753 ;
  assign n8774 = ~n3762 & n8773 ;
  assign n8775 = ~n8772 & ~n8774 ;
  assign n8776 = ~\ctl_rf_c1_rf_chdad_reg[8]/NET0131  & ~n8753 ;
  assign n8777 = \hwdata[8]_pad  & ~n2242 ;
  assign n8778 = \hwdata[16]_pad  & n2242 ;
  assign n8779 = ~n8777 & ~n8778 ;
  assign n8780 = ~n2240 & ~n8779 ;
  assign n8781 = \hwdata[24]_pad  & n2240 ;
  assign n8782 = n8753 & ~n8781 ;
  assign n8783 = ~n8780 & n8782 ;
  assign n8784 = ~n8776 & ~n8783 ;
  assign n8785 = n2231 & n8752 ;
  assign n8786 = ~\ctl_rf_c1_rf_chsad_reg[11]/NET0131  & ~n8785 ;
  assign n8787 = \hwdata[11]_pad  & ~n2242 ;
  assign n8788 = \hwdata[19]_pad  & n2242 ;
  assign n8789 = ~n8787 & ~n8788 ;
  assign n8790 = ~n2240 & ~n8789 ;
  assign n8791 = \hwdata[27]_pad  & n2240 ;
  assign n8792 = n8785 & ~n8791 ;
  assign n8793 = ~n8790 & n8792 ;
  assign n8794 = ~n8786 & ~n8793 ;
  assign n8795 = ~\ctl_rf_c1_rf_chsad_reg[5]/NET0131  & ~n2236 ;
  assign n8796 = n2236 & ~n8587 ;
  assign n8797 = ~n8586 & n8796 ;
  assign n8798 = ~n8795 & ~n8797 ;
  assign n8799 = ~\ctl_rf_c1_rf_chsad_reg[6]/NET0131  & ~n2236 ;
  assign n8800 = n2236 & ~n8596 ;
  assign n8801 = ~n8595 & n8800 ;
  assign n8802 = ~n8799 & ~n8801 ;
  assign n8803 = ~\ctl_rf_c1_rf_chsad_reg[9]/NET0131  & ~n8785 ;
  assign n8804 = \hwdata[9]_pad  & ~n2242 ;
  assign n8805 = \hwdata[17]_pad  & n2242 ;
  assign n8806 = ~n8804 & ~n8805 ;
  assign n8807 = ~n2240 & ~n8806 ;
  assign n8808 = \hwdata[25]_pad  & n2240 ;
  assign n8809 = n8785 & ~n8808 ;
  assign n8810 = ~n8807 & n8809 ;
  assign n8811 = ~n8803 & ~n8810 ;
  assign n8812 = n2266 & n8752 ;
  assign n8813 = ~\ctl_rf_c3_rf_chdad_reg[10]/NET0131  & ~n8812 ;
  assign n8814 = ~n8759 & n8812 ;
  assign n8815 = ~n8758 & n8814 ;
  assign n8816 = ~n8813 & ~n8815 ;
  assign n8817 = ~\ctl_rf_c3_rf_chdad_reg[11]/NET0131  & ~n8812 ;
  assign n8818 = ~n8791 & n8812 ;
  assign n8819 = ~n8790 & n8818 ;
  assign n8820 = ~n8817 & ~n8819 ;
  assign n8821 = ~\ctl_rf_c3_rf_chdad_reg[12]/NET0131  & ~n8812 ;
  assign n8822 = ~n8768 & n8812 ;
  assign n8823 = ~n8767 & n8822 ;
  assign n8824 = ~n8821 & ~n8823 ;
  assign n8825 = ~\ctl_rf_c3_rf_chdad_reg[15]/NET0131  & ~n8812 ;
  assign n8826 = ~n3763 & n8812 ;
  assign n8827 = ~n3762 & n8826 ;
  assign n8828 = ~n8825 & ~n8827 ;
  assign n8829 = ~\ctl_rf_c3_rf_chdad_reg[8]/NET0131  & ~n8812 ;
  assign n8830 = ~n8781 & n8812 ;
  assign n8831 = ~n8780 & n8830 ;
  assign n8832 = ~n8829 & ~n8831 ;
  assign n8833 = ~\ctl_rf_c3_rf_chsad_reg[5]/NET0131  & ~n8604 ;
  assign n8834 = ~n8587 & n8604 ;
  assign n8835 = ~n8586 & n8834 ;
  assign n8836 = ~n8833 & ~n8835 ;
  assign n8837 = ~\ctl_rf_c3_rf_chsad_reg[6]/NET0131  & ~n8604 ;
  assign n8838 = ~n8596 & n8604 ;
  assign n8839 = ~n8595 & n8838 ;
  assign n8840 = ~n8837 & ~n8839 ;
  assign n8841 = n2311 & n8752 ;
  assign n8842 = ~\ctl_rf_c3_rf_chsad_reg[9]/NET0131  & ~n8841 ;
  assign n8843 = ~n8808 & n8841 ;
  assign n8844 = ~n8807 & n8843 ;
  assign n8845 = ~n8842 & ~n8844 ;
  assign n8846 = \ctl_rf_be_d1_reg[1]/P0001  & n2276 ;
  assign n8847 = n2274 & n8846 ;
  assign n8848 = ~\ctl_rf_c4_rf_chdad_reg[8]/NET0131  & ~n8847 ;
  assign n8849 = ~n8781 & n8847 ;
  assign n8850 = ~n8780 & n8849 ;
  assign n8851 = ~n8848 & ~n8850 ;
  assign n8852 = n2317 & n8846 ;
  assign n8853 = ~\ctl_rf_c4_rf_chsad_reg[10]/NET0131  & ~n8852 ;
  assign n8854 = ~n8759 & n8852 ;
  assign n8855 = ~n8758 & n8854 ;
  assign n8856 = ~n8853 & ~n8855 ;
  assign n8857 = ~\ctl_rf_c4_rf_chsad_reg[11]/NET0131  & ~n8852 ;
  assign n8858 = ~n8791 & n8852 ;
  assign n8859 = ~n8790 & n8858 ;
  assign n8860 = ~n8857 & ~n8859 ;
  assign n8861 = ~\ctl_rf_c4_rf_chsad_reg[12]/NET0131  & ~n8852 ;
  assign n8862 = ~n8768 & n8852 ;
  assign n8863 = ~n8767 & n8862 ;
  assign n8864 = ~n8861 & ~n8863 ;
  assign n8865 = ~\ctl_rf_c4_rf_chsad_reg[15]/NET0131  & ~n8852 ;
  assign n8866 = ~n3763 & n8852 ;
  assign n8867 = ~n3762 & n8866 ;
  assign n8868 = ~n8865 & ~n8867 ;
  assign n8869 = ~\ctl_rf_c4_rf_chsad_reg[5]/NET0131  & ~n8624 ;
  assign n8870 = ~n8587 & n8624 ;
  assign n8871 = ~n8586 & n8870 ;
  assign n8872 = ~n8869 & ~n8871 ;
  assign n8873 = ~\ctl_rf_c4_rf_chsad_reg[6]/NET0131  & ~n8624 ;
  assign n8874 = ~n8596 & n8624 ;
  assign n8875 = ~n8595 & n8874 ;
  assign n8876 = ~n8873 & ~n8875 ;
  assign n8877 = ~\ctl_rf_c4_rf_chsad_reg[9]/NET0131  & ~n8852 ;
  assign n8878 = ~n8808 & n8852 ;
  assign n8879 = ~n8807 & n8878 ;
  assign n8880 = ~n8877 & ~n8879 ;
  assign n8881 = n2274 & n8752 ;
  assign n8882 = ~\ctl_rf_c5_rf_chdad_reg[8]/NET0131  & ~n8881 ;
  assign n8883 = ~n8781 & n8881 ;
  assign n8884 = ~n8780 & n8883 ;
  assign n8885 = ~n8882 & ~n8884 ;
  assign n8886 = n2317 & n8752 ;
  assign n8887 = ~\ctl_rf_c5_rf_chsad_reg[10]/NET0131  & ~n8886 ;
  assign n8888 = ~n8759 & n8886 ;
  assign n8889 = ~n8758 & n8888 ;
  assign n8890 = ~n8887 & ~n8889 ;
  assign n8891 = ~\ctl_rf_c5_rf_chsad_reg[11]/NET0131  & ~n8886 ;
  assign n8892 = ~n8791 & n8886 ;
  assign n8893 = ~n8790 & n8892 ;
  assign n8894 = ~n8891 & ~n8893 ;
  assign n8895 = ~\ctl_rf_c5_rf_chsad_reg[12]/NET0131  & ~n8886 ;
  assign n8896 = ~n8768 & n8886 ;
  assign n8897 = ~n8767 & n8896 ;
  assign n8898 = ~n8895 & ~n8897 ;
  assign n8899 = ~\ctl_rf_c5_rf_chsad_reg[15]/NET0131  & ~n8886 ;
  assign n8900 = ~n3763 & n8886 ;
  assign n8901 = ~n3762 & n8900 ;
  assign n8902 = ~n8899 & ~n8901 ;
  assign n8903 = ~\ctl_rf_c5_rf_chsad_reg[5]/NET0131  & ~n8641 ;
  assign n8904 = ~n8587 & n8641 ;
  assign n8905 = ~n8586 & n8904 ;
  assign n8906 = ~n8903 & ~n8905 ;
  assign n8907 = ~\ctl_rf_c5_rf_chsad_reg[6]/NET0131  & ~n8641 ;
  assign n8908 = ~n8596 & n8641 ;
  assign n8909 = ~n8595 & n8908 ;
  assign n8910 = ~n8907 & ~n8909 ;
  assign n8911 = ~\ctl_rf_c5_rf_chsad_reg[9]/NET0131  & ~n8886 ;
  assign n8912 = ~n8808 & n8886 ;
  assign n8913 = ~n8807 & n8912 ;
  assign n8914 = ~n8911 & ~n8913 ;
  assign n8915 = n2289 & n8846 ;
  assign n8916 = ~\ctl_rf_c6_rf_chdad_reg[10]/NET0131  & ~n8915 ;
  assign n8917 = ~n8759 & n8915 ;
  assign n8918 = ~n8758 & n8917 ;
  assign n8919 = ~n8916 & ~n8918 ;
  assign n8920 = ~\ctl_rf_c6_rf_chdad_reg[8]/NET0131  & ~n8915 ;
  assign n8921 = ~n8781 & n8915 ;
  assign n8922 = ~n8780 & n8921 ;
  assign n8923 = ~n8920 & ~n8922 ;
  assign n8924 = n2324 & n8846 ;
  assign n8925 = ~\ctl_rf_c6_rf_chsad_reg[11]/NET0131  & ~n8924 ;
  assign n8926 = ~n8791 & n8924 ;
  assign n8927 = ~n8790 & n8926 ;
  assign n8928 = ~n8925 & ~n8927 ;
  assign n8929 = ~\ctl_rf_c6_rf_chsad_reg[12]/NET0131  & ~n8924 ;
  assign n8930 = ~n8768 & n8924 ;
  assign n8931 = ~n8767 & n8930 ;
  assign n8932 = ~n8929 & ~n8931 ;
  assign n8933 = ~\ctl_rf_c6_rf_chsad_reg[15]/NET0131  & ~n8924 ;
  assign n8934 = ~n3763 & n8924 ;
  assign n8935 = ~n3762 & n8934 ;
  assign n8936 = ~n8933 & ~n8935 ;
  assign n8937 = ~\ctl_rf_c6_rf_chsad_reg[5]/NET0131  & ~n8651 ;
  assign n8938 = ~n8587 & n8651 ;
  assign n8939 = ~n8586 & n8938 ;
  assign n8940 = ~n8937 & ~n8939 ;
  assign n8941 = ~\ctl_rf_c6_rf_chsad_reg[6]/NET0131  & ~n8651 ;
  assign n8942 = ~n8596 & n8651 ;
  assign n8943 = ~n8595 & n8942 ;
  assign n8944 = ~n8941 & ~n8943 ;
  assign n8945 = ~\ctl_rf_c6_rf_chsad_reg[9]/NET0131  & ~n8924 ;
  assign n8946 = ~n8808 & n8924 ;
  assign n8947 = ~n8807 & n8946 ;
  assign n8948 = ~n8945 & ~n8947 ;
  assign n8949 = n2289 & n8752 ;
  assign n8950 = ~\ctl_rf_c7_rf_chdad_reg[11]/NET0131  & ~n8949 ;
  assign n8951 = ~n8791 & n8949 ;
  assign n8952 = ~n8790 & n8951 ;
  assign n8953 = ~n8950 & ~n8952 ;
  assign n8954 = ~\ctl_rf_c7_rf_chdad_reg[15]/NET0131  & ~n8949 ;
  assign n8955 = ~n3763 & n8949 ;
  assign n8956 = ~n3762 & n8955 ;
  assign n8957 = ~n8954 & ~n8956 ;
  assign n8958 = ~\ctl_rf_c7_rf_chdad_reg[8]/NET0131  & ~n8949 ;
  assign n8959 = ~n8781 & n8949 ;
  assign n8960 = ~n8780 & n8959 ;
  assign n8961 = ~n8958 & ~n8960 ;
  assign n8962 = n2324 & n8752 ;
  assign n8963 = ~\ctl_rf_c7_rf_chsad_reg[10]/NET0131  & ~n8962 ;
  assign n8964 = ~n8759 & n8962 ;
  assign n8965 = ~n8758 & n8964 ;
  assign n8966 = ~n8963 & ~n8965 ;
  assign n8967 = ~\ctl_rf_c7_rf_chsad_reg[12]/NET0131  & ~n8962 ;
  assign n8968 = ~n8768 & n8962 ;
  assign n8969 = ~n8767 & n8968 ;
  assign n8970 = ~n8967 & ~n8969 ;
  assign n8971 = ~\ctl_rf_c7_rf_chsad_reg[5]/NET0131  & ~n8672 ;
  assign n8972 = ~n8587 & n8672 ;
  assign n8973 = ~n8586 & n8972 ;
  assign n8974 = ~n8971 & ~n8973 ;
  assign n8975 = ~\ctl_rf_c7_rf_chsad_reg[6]/NET0131  & ~n8672 ;
  assign n8976 = ~n8596 & n8672 ;
  assign n8977 = ~n8595 & n8976 ;
  assign n8978 = ~n8975 & ~n8977 ;
  assign n8979 = ~\ctl_rf_c7_rf_chsad_reg[9]/NET0131  & ~n8962 ;
  assign n8980 = ~n8808 & n8962 ;
  assign n8981 = ~n8807 & n8980 ;
  assign n8982 = ~n8979 & ~n8981 ;
  assign n8983 = ~\ctl_rf_c1_rf_chsad_reg[0]/NET0131  & ~n2236 ;
  assign n8984 = n2236 & ~n3771 ;
  assign n8985 = ~n3770 & n8984 ;
  assign n8986 = ~n8983 & ~n8985 ;
  assign n8987 = ~\ctl_rf_c1_rf_chsad_reg[1]/NET0131  & ~n2236 ;
  assign n8988 = \hwdata[1]_pad  & ~n2242 ;
  assign n8989 = \hwdata[25]_pad  & n2242 ;
  assign n8990 = ~n8988 & ~n8989 ;
  assign n8991 = ~n2240 & ~n8990 ;
  assign n8992 = \hwdata[17]_pad  & n2240 ;
  assign n8993 = n2236 & ~n8992 ;
  assign n8994 = ~n8991 & n8993 ;
  assign n8995 = ~n8987 & ~n8994 ;
  assign n8996 = ~\ctl_rf_c1_rf_chsad_reg[2]/NET0131  & ~n2236 ;
  assign n8997 = \hwdata[2]_pad  & ~n2242 ;
  assign n8998 = \hwdata[26]_pad  & n2242 ;
  assign n8999 = ~n8997 & ~n8998 ;
  assign n9000 = ~n2240 & ~n8999 ;
  assign n9001 = \hwdata[18]_pad  & n2240 ;
  assign n9002 = n2236 & ~n9001 ;
  assign n9003 = ~n9000 & n9002 ;
  assign n9004 = ~n8996 & ~n9003 ;
  assign n9005 = ~\ctl_rf_c1_rf_chsad_reg[4]/NET0131  & ~n2236 ;
  assign n9006 = n2236 & ~n8714 ;
  assign n9007 = ~n8713 & n9006 ;
  assign n9008 = ~n9005 & ~n9007 ;
  assign n9009 = ~\ctl_rf_c3_rf_chsad_reg[0]/NET0131  & ~n8604 ;
  assign n9010 = ~n3771 & n8604 ;
  assign n9011 = ~n3770 & n9010 ;
  assign n9012 = ~n9009 & ~n9011 ;
  assign n9013 = ~\ctl_rf_c3_rf_chsad_reg[13]/NET0131  & ~n8841 ;
  assign n9014 = \hwdata[13]_pad  & ~n2242 ;
  assign n9015 = \hwdata[21]_pad  & n2242 ;
  assign n9016 = ~n9014 & ~n9015 ;
  assign n9017 = ~n2240 & ~n9016 ;
  assign n9018 = \hwdata[29]_pad  & n2240 ;
  assign n9019 = n8841 & ~n9018 ;
  assign n9020 = ~n9017 & n9019 ;
  assign n9021 = ~n9013 & ~n9020 ;
  assign n9022 = ~\ctl_rf_c3_rf_chsad_reg[14]/NET0131  & ~n8841 ;
  assign n9023 = \hwdata[14]_pad  & ~n2242 ;
  assign n9024 = \hwdata[22]_pad  & n2242 ;
  assign n9025 = ~n9023 & ~n9024 ;
  assign n9026 = ~n2240 & ~n9025 ;
  assign n9027 = \hwdata[30]_pad  & n2240 ;
  assign n9028 = n8841 & ~n9027 ;
  assign n9029 = ~n9026 & n9028 ;
  assign n9030 = ~n9022 & ~n9029 ;
  assign n9031 = ~\ctl_rf_c3_rf_chsad_reg[1]/NET0131  & ~n8604 ;
  assign n9032 = n8604 & ~n8992 ;
  assign n9033 = ~n8991 & n9032 ;
  assign n9034 = ~n9031 & ~n9033 ;
  assign n9035 = ~\ctl_rf_c3_rf_chsad_reg[2]/NET0131  & ~n8604 ;
  assign n9036 = n8604 & ~n9001 ;
  assign n9037 = ~n9000 & n9036 ;
  assign n9038 = ~n9035 & ~n9037 ;
  assign n9039 = ~\ctl_rf_c3_rf_chsad_reg[3]/NET0131  & ~n8604 ;
  assign n9040 = \hwdata[3]_pad  & ~n2242 ;
  assign n9041 = \hwdata[27]_pad  & n2242 ;
  assign n9042 = ~n9040 & ~n9041 ;
  assign n9043 = ~n2240 & ~n9042 ;
  assign n9044 = \hwdata[19]_pad  & n2240 ;
  assign n9045 = n8604 & ~n9044 ;
  assign n9046 = ~n9043 & n9045 ;
  assign n9047 = ~n9039 & ~n9046 ;
  assign n9048 = ~\ctl_rf_c3_rf_chsad_reg[4]/NET0131  & ~n8604 ;
  assign n9049 = n8604 & ~n8714 ;
  assign n9050 = ~n8713 & n9049 ;
  assign n9051 = ~n9048 & ~n9050 ;
  assign n9052 = n2274 & n8623 ;
  assign n9053 = ~\ctl_rf_c4_rf_chdad_reg[0]/NET0131  & ~n9052 ;
  assign n9054 = ~n3771 & n9052 ;
  assign n9055 = ~n3770 & n9054 ;
  assign n9056 = ~n9053 & ~n9055 ;
  assign n9057 = ~\ctl_rf_c4_rf_chdad_reg[1]/NET0131  & ~n9052 ;
  assign n9058 = ~n8992 & n9052 ;
  assign n9059 = ~n8991 & n9058 ;
  assign n9060 = ~n9057 & ~n9059 ;
  assign n9061 = ~\ctl_rf_c4_rf_chdad_reg[2]/NET0131  & ~n9052 ;
  assign n9062 = ~n9001 & n9052 ;
  assign n9063 = ~n9000 & n9062 ;
  assign n9064 = ~n9061 & ~n9063 ;
  assign n9065 = ~\ctl_rf_c4_rf_chsad_reg[0]/NET0131  & ~n8624 ;
  assign n9066 = ~n3771 & n8624 ;
  assign n9067 = ~n3770 & n9066 ;
  assign n9068 = ~n9065 & ~n9067 ;
  assign n9069 = ~\ctl_rf_c4_rf_chsad_reg[13]/NET0131  & ~n8852 ;
  assign n9070 = n8852 & ~n9018 ;
  assign n9071 = ~n9017 & n9070 ;
  assign n9072 = ~n9069 & ~n9071 ;
  assign n9073 = ~\ctl_rf_c4_rf_chsad_reg[14]/NET0131  & ~n8852 ;
  assign n9074 = n8852 & ~n9027 ;
  assign n9075 = ~n9026 & n9074 ;
  assign n9076 = ~n9073 & ~n9075 ;
  assign n9077 = ~\ctl_rf_c4_rf_chsad_reg[1]/NET0131  & ~n8624 ;
  assign n9078 = n8624 & ~n8992 ;
  assign n9079 = ~n8991 & n9078 ;
  assign n9080 = ~n9077 & ~n9079 ;
  assign n9081 = ~\ctl_rf_c4_rf_chsad_reg[2]/NET0131  & ~n8624 ;
  assign n9082 = n8624 & ~n9001 ;
  assign n9083 = ~n9000 & n9082 ;
  assign n9084 = ~n9081 & ~n9083 ;
  assign n9085 = ~\ctl_rf_c4_rf_chsad_reg[3]/NET0131  & ~n8624 ;
  assign n9086 = n8624 & ~n9044 ;
  assign n9087 = ~n9043 & n9086 ;
  assign n9088 = ~n9085 & ~n9087 ;
  assign n9089 = ~\ctl_rf_c4_rf_chsad_reg[4]/NET0131  & ~n8624 ;
  assign n9090 = n8624 & ~n8714 ;
  assign n9091 = ~n8713 & n9090 ;
  assign n9092 = ~n9089 & ~n9091 ;
  assign n9093 = n2289 & n8623 ;
  assign n9094 = ~\ctl_rf_c6_rf_chdad_reg[0]/NET0131  & ~n9093 ;
  assign n9095 = ~n3771 & n9093 ;
  assign n9096 = ~n3770 & n9095 ;
  assign n9097 = ~n9094 & ~n9096 ;
  assign n9098 = ~\ctl_rf_c6_rf_chdad_reg[13]/NET0131  & ~n8915 ;
  assign n9099 = n8915 & ~n9018 ;
  assign n9100 = ~n9017 & n9099 ;
  assign n9101 = ~n9098 & ~n9100 ;
  assign n9102 = ~\ctl_rf_c6_rf_chdad_reg[1]/NET0131  & ~n9093 ;
  assign n9103 = ~n8992 & n9093 ;
  assign n9104 = ~n8991 & n9103 ;
  assign n9105 = ~n9102 & ~n9104 ;
  assign n9106 = ~\ctl_rf_c6_rf_chdad_reg[2]/NET0131  & ~n9093 ;
  assign n9107 = ~n9001 & n9093 ;
  assign n9108 = ~n9000 & n9107 ;
  assign n9109 = ~n9106 & ~n9108 ;
  assign n9110 = ~\ctl_rf_c6_rf_chsad_reg[0]/NET0131  & ~n8651 ;
  assign n9111 = ~n3771 & n8651 ;
  assign n9112 = ~n3770 & n9111 ;
  assign n9113 = ~n9110 & ~n9112 ;
  assign n9114 = ~\ctl_rf_c6_rf_chsad_reg[14]/NET0131  & ~n8924 ;
  assign n9115 = n8924 & ~n9027 ;
  assign n9116 = ~n9026 & n9115 ;
  assign n9117 = ~n9114 & ~n9116 ;
  assign n9118 = ~\ctl_rf_c6_rf_chsad_reg[1]/NET0131  & ~n8651 ;
  assign n9119 = n8651 & ~n8992 ;
  assign n9120 = ~n8991 & n9119 ;
  assign n9121 = ~n9118 & ~n9120 ;
  assign n9122 = ~\ctl_rf_c6_rf_chsad_reg[2]/NET0131  & ~n8651 ;
  assign n9123 = n8651 & ~n9001 ;
  assign n9124 = ~n9000 & n9123 ;
  assign n9125 = ~n9122 & ~n9124 ;
  assign n9126 = ~\ctl_rf_c6_rf_chsad_reg[3]/NET0131  & ~n8651 ;
  assign n9127 = n8651 & ~n9044 ;
  assign n9128 = ~n9043 & n9127 ;
  assign n9129 = ~n9126 & ~n9128 ;
  assign n9130 = ~\ctl_rf_c6_rf_chsad_reg[4]/NET0131  & ~n8651 ;
  assign n9131 = n8651 & ~n8714 ;
  assign n9132 = ~n8713 & n9131 ;
  assign n9133 = ~n9130 & ~n9132 ;
  assign n9134 = n2252 & n8623 ;
  assign n9135 = ~\ctl_rf_c0_rf_chdad_reg[1]/NET0131  & ~n9134 ;
  assign n9136 = ~n8992 & n9134 ;
  assign n9137 = ~n8991 & n9136 ;
  assign n9138 = ~n9135 & ~n9137 ;
  assign n9139 = ~\ctl_rf_c0_rf_chdad_reg[2]/NET0131  & ~n9134 ;
  assign n9140 = ~n9001 & n9134 ;
  assign n9141 = ~n9000 & n9140 ;
  assign n9142 = ~n9139 & ~n9141 ;
  assign n9143 = n2252 & n8846 ;
  assign n9144 = ~\ctl_rf_c0_rf_chdad_reg[8]/NET0131  & ~n9143 ;
  assign n9145 = ~n8781 & n9143 ;
  assign n9146 = ~n8780 & n9145 ;
  assign n9147 = ~n9144 & ~n9146 ;
  assign n9148 = ~\ctl_rf_c0_rf_chsad_reg[0]/NET0131  & ~n8691 ;
  assign n9149 = ~n3771 & n8691 ;
  assign n9150 = ~n3770 & n9149 ;
  assign n9151 = ~n9148 & ~n9150 ;
  assign n9152 = n2231 & n8846 ;
  assign n9153 = ~\ctl_rf_c0_rf_chsad_reg[10]/NET0131  & ~n9152 ;
  assign n9154 = ~n8759 & n9152 ;
  assign n9155 = ~n8758 & n9154 ;
  assign n9156 = ~n9153 & ~n9155 ;
  assign n9157 = ~\ctl_rf_c0_rf_chsad_reg[13]/NET0131  & ~n9152 ;
  assign n9158 = ~n9018 & n9152 ;
  assign n9159 = ~n9017 & n9158 ;
  assign n9160 = ~n9157 & ~n9159 ;
  assign n9161 = ~\ctl_rf_c0_rf_chsad_reg[1]/NET0131  & ~n8691 ;
  assign n9162 = n8691 & ~n8992 ;
  assign n9163 = ~n8991 & n9162 ;
  assign n9164 = ~n9161 & ~n9163 ;
  assign n9165 = ~\ctl_rf_c0_rf_chsad_reg[2]/NET0131  & ~n8691 ;
  assign n9166 = n8691 & ~n9001 ;
  assign n9167 = ~n9000 & n9166 ;
  assign n9168 = ~n9165 & ~n9167 ;
  assign n9169 = ~\ctl_rf_c0_rf_chsad_reg[3]/NET0131  & ~n8691 ;
  assign n9170 = n8691 & ~n9044 ;
  assign n9171 = ~n9043 & n9170 ;
  assign n9172 = ~n9169 & ~n9171 ;
  assign n9173 = ~\ctl_rf_c0_rf_chsad_reg[4]/NET0131  & ~n8691 ;
  assign n9174 = n8691 & ~n8714 ;
  assign n9175 = ~n8713 & n9174 ;
  assign n9176 = ~n9173 & ~n9175 ;
  assign n9177 = ~\ctl_rf_c0_rf_chsad_reg[5]/NET0131  & ~n8691 ;
  assign n9178 = ~n8587 & n8691 ;
  assign n9179 = ~n8586 & n9178 ;
  assign n9180 = ~n9177 & ~n9179 ;
  assign n9181 = ~\ctl_rf_c0_rf_chsad_reg[6]/NET0131  & ~n8691 ;
  assign n9182 = ~n8596 & n8691 ;
  assign n9183 = ~n8595 & n9182 ;
  assign n9184 = ~n9181 & ~n9183 ;
  assign n9185 = ~\ctl_rf_c0_rf_chsad_reg[9]/NET0131  & ~n9152 ;
  assign n9186 = ~n8808 & n9152 ;
  assign n9187 = ~n8807 & n9186 ;
  assign n9188 = ~n9185 & ~n9187 ;
  assign n9189 = ~\ctl_rf_c0_rf_chtsz_reg[4]/NET0131  & ~n8696 ;
  assign n9190 = n8696 & ~n8714 ;
  assign n9191 = ~n8713 & n9190 ;
  assign n9192 = ~n9189 & ~n9191 ;
  assign n9193 = n2235 & n2252 ;
  assign n9194 = ~\ctl_rf_c1_rf_chdad_reg[0]/NET0131  & ~n9193 ;
  assign n9195 = ~n3771 & n9193 ;
  assign n9196 = ~n3770 & n9195 ;
  assign n9197 = ~n9194 & ~n9196 ;
  assign n9198 = ~\ctl_rf_c1_rf_chdad_reg[13]/NET0131  & ~n8753 ;
  assign n9199 = n8753 & ~n9018 ;
  assign n9200 = ~n9017 & n9199 ;
  assign n9201 = ~n9198 & ~n9200 ;
  assign n9202 = ~\ctl_rf_c1_rf_chdad_reg[14]/NET0131  & ~n8753 ;
  assign n9203 = n8753 & ~n9027 ;
  assign n9204 = ~n9026 & n9203 ;
  assign n9205 = ~n9202 & ~n9204 ;
  assign n9206 = ~\ctl_rf_c1_rf_chdad_reg[1]/NET0131  & ~n9193 ;
  assign n9207 = ~n8992 & n9193 ;
  assign n9208 = ~n8991 & n9207 ;
  assign n9209 = ~n9206 & ~n9208 ;
  assign n9210 = ~\ctl_rf_c1_rf_chdad_reg[2]/NET0131  & ~n9193 ;
  assign n9211 = ~n9001 & n9193 ;
  assign n9212 = ~n9000 & n9211 ;
  assign n9213 = ~n9210 & ~n9212 ;
  assign n9214 = n2266 & n8623 ;
  assign n9215 = ~\ctl_rf_c2_rf_chdad_reg[0]/NET0131  & ~n9214 ;
  assign n9216 = ~n3771 & n9214 ;
  assign n9217 = ~n3770 & n9216 ;
  assign n9218 = ~n9215 & ~n9217 ;
  assign n9219 = ~\ctl_rf_c2_rf_chdad_reg[1]/NET0131  & ~n9214 ;
  assign n9220 = ~n8992 & n9214 ;
  assign n9221 = ~n8991 & n9220 ;
  assign n9222 = ~n9219 & ~n9221 ;
  assign n9223 = ~\ctl_rf_c2_rf_chdad_reg[2]/NET0131  & ~n9214 ;
  assign n9224 = ~n9001 & n9214 ;
  assign n9225 = ~n9000 & n9224 ;
  assign n9226 = ~n9223 & ~n9225 ;
  assign n9227 = n2266 & n8846 ;
  assign n9228 = ~\ctl_rf_c2_rf_chdad_reg[8]/NET0131  & ~n9227 ;
  assign n9229 = ~n8781 & n9227 ;
  assign n9230 = ~n8780 & n9229 ;
  assign n9231 = ~n9228 & ~n9230 ;
  assign n9232 = n2311 & n8846 ;
  assign n9233 = ~\ctl_rf_c2_rf_chsad_reg[10]/NET0131  & ~n9232 ;
  assign n9234 = ~n8759 & n9232 ;
  assign n9235 = ~n8758 & n9234 ;
  assign n9236 = ~n9233 & ~n9235 ;
  assign n9237 = ~\ctl_rf_c2_rf_chsad_reg[0]/NET0131  & ~n8718 ;
  assign n9238 = ~n3771 & n8718 ;
  assign n9239 = ~n3770 & n9238 ;
  assign n9240 = ~n9237 & ~n9239 ;
  assign n9241 = ~\ctl_rf_c2_rf_chsad_reg[11]/NET0131  & ~n9232 ;
  assign n9242 = ~n8791 & n9232 ;
  assign n9243 = ~n8790 & n9242 ;
  assign n9244 = ~n9241 & ~n9243 ;
  assign n9245 = ~\ctl_rf_c2_rf_chsad_reg[12]/NET0131  & ~n9232 ;
  assign n9246 = ~n8768 & n9232 ;
  assign n9247 = ~n8767 & n9246 ;
  assign n9248 = ~n9245 & ~n9247 ;
  assign n9249 = ~\ctl_rf_c2_rf_chsad_reg[13]/NET0131  & ~n9232 ;
  assign n9250 = ~n9018 & n9232 ;
  assign n9251 = ~n9017 & n9250 ;
  assign n9252 = ~n9249 & ~n9251 ;
  assign n9253 = ~\ctl_rf_c2_rf_chsad_reg[14]/NET0131  & ~n9232 ;
  assign n9254 = ~n9027 & n9232 ;
  assign n9255 = ~n9026 & n9254 ;
  assign n9256 = ~n9253 & ~n9255 ;
  assign n9257 = ~\ctl_rf_c2_rf_chsad_reg[1]/NET0131  & ~n8718 ;
  assign n9258 = n8718 & ~n8992 ;
  assign n9259 = ~n8991 & n9258 ;
  assign n9260 = ~n9257 & ~n9259 ;
  assign n9261 = ~\ctl_rf_c2_rf_chsad_reg[2]/NET0131  & ~n8718 ;
  assign n9262 = n8718 & ~n9001 ;
  assign n9263 = ~n9000 & n9262 ;
  assign n9264 = ~n9261 & ~n9263 ;
  assign n9265 = ~\ctl_rf_c2_rf_chsad_reg[3]/NET0131  & ~n8718 ;
  assign n9266 = n8718 & ~n9044 ;
  assign n9267 = ~n9043 & n9266 ;
  assign n9268 = ~n9265 & ~n9267 ;
  assign n9269 = ~\ctl_rf_c2_rf_chsad_reg[4]/NET0131  & ~n8718 ;
  assign n9270 = ~n8714 & n8718 ;
  assign n9271 = ~n8713 & n9270 ;
  assign n9272 = ~n9269 & ~n9271 ;
  assign n9273 = ~\ctl_rf_c2_rf_chsad_reg[5]/NET0131  & ~n8718 ;
  assign n9274 = ~n8587 & n8718 ;
  assign n9275 = ~n8586 & n9274 ;
  assign n9276 = ~n9273 & ~n9275 ;
  assign n9277 = ~\ctl_rf_c2_rf_chsad_reg[6]/NET0131  & ~n8718 ;
  assign n9278 = ~n8596 & n8718 ;
  assign n9279 = ~n8595 & n9278 ;
  assign n9280 = ~n9277 & ~n9279 ;
  assign n9281 = ~\ctl_rf_c2_rf_chsad_reg[9]/NET0131  & ~n9232 ;
  assign n9282 = ~n8808 & n9232 ;
  assign n9283 = ~n8807 & n9282 ;
  assign n9284 = ~n9281 & ~n9283 ;
  assign n9285 = ~\ctl_rf_c2_rf_chtsz_reg[4]/NET0131  & ~n8723 ;
  assign n9286 = ~n8714 & n8723 ;
  assign n9287 = ~n8713 & n9286 ;
  assign n9288 = ~n9285 & ~n9287 ;
  assign n9289 = n2235 & n2266 ;
  assign n9290 = ~\ctl_rf_c3_rf_chdad_reg[0]/NET0131  & ~n9289 ;
  assign n9291 = ~n3771 & n9289 ;
  assign n9292 = ~n3770 & n9291 ;
  assign n9293 = ~n9290 & ~n9292 ;
  assign n9294 = ~\ctl_rf_c3_rf_chdad_reg[1]/NET0131  & ~n9289 ;
  assign n9295 = ~n8992 & n9289 ;
  assign n9296 = ~n8991 & n9295 ;
  assign n9297 = ~n9294 & ~n9296 ;
  assign n9298 = ~\ctl_rf_c3_rf_chdad_reg[2]/NET0131  & ~n9289 ;
  assign n9299 = ~n9001 & n9289 ;
  assign n9300 = ~n9000 & n9299 ;
  assign n9301 = ~n9298 & ~n9300 ;
  assign n9302 = n2235 & n2274 ;
  assign n9303 = ~\ctl_rf_c5_rf_chdad_reg[0]/NET0131  & ~n9302 ;
  assign n9304 = ~n3771 & n9302 ;
  assign n9305 = ~n3770 & n9304 ;
  assign n9306 = ~n9303 & ~n9305 ;
  assign n9307 = ~\ctl_rf_c5_rf_chdad_reg[13]/NET0131  & ~n8881 ;
  assign n9308 = n8881 & ~n9018 ;
  assign n9309 = ~n9017 & n9308 ;
  assign n9310 = ~n9307 & ~n9309 ;
  assign n9311 = ~\ctl_rf_c5_rf_chdad_reg[2]/NET0131  & ~n9302 ;
  assign n9312 = ~n9001 & n9302 ;
  assign n9313 = ~n9000 & n9312 ;
  assign n9314 = ~n9311 & ~n9313 ;
  assign n9315 = ~\ctl_rf_c5_rf_chsad_reg[0]/NET0131  & ~n8641 ;
  assign n9316 = ~n3771 & n8641 ;
  assign n9317 = ~n3770 & n9316 ;
  assign n9318 = ~n9315 & ~n9317 ;
  assign n9319 = ~\ctl_rf_c5_rf_chsad_reg[14]/NET0131  & ~n8886 ;
  assign n9320 = n8886 & ~n9027 ;
  assign n9321 = ~n9026 & n9320 ;
  assign n9322 = ~n9319 & ~n9321 ;
  assign n9323 = ~\ctl_rf_c5_rf_chsad_reg[1]/NET0131  & ~n8641 ;
  assign n9324 = n8641 & ~n8992 ;
  assign n9325 = ~n8991 & n9324 ;
  assign n9326 = ~n9323 & ~n9325 ;
  assign n9327 = ~\ctl_rf_c5_rf_chsad_reg[2]/NET0131  & ~n8641 ;
  assign n9328 = n8641 & ~n9001 ;
  assign n9329 = ~n9000 & n9328 ;
  assign n9330 = ~n9327 & ~n9329 ;
  assign n9331 = ~\ctl_rf_c5_rf_chsad_reg[3]/NET0131  & ~n8641 ;
  assign n9332 = n8641 & ~n9044 ;
  assign n9333 = ~n9043 & n9332 ;
  assign n9334 = ~n9331 & ~n9333 ;
  assign n9335 = ~\ctl_rf_c5_rf_chsad_reg[4]/NET0131  & ~n8641 ;
  assign n9336 = n8641 & ~n8714 ;
  assign n9337 = ~n8713 & n9336 ;
  assign n9338 = ~n9335 & ~n9337 ;
  assign n9339 = n2235 & n2289 ;
  assign n9340 = ~\ctl_rf_c7_rf_chdad_reg[0]/NET0131  & ~n9339 ;
  assign n9341 = ~n3771 & n9339 ;
  assign n9342 = ~n3770 & n9341 ;
  assign n9343 = ~n9340 & ~n9342 ;
  assign n9344 = ~\ctl_rf_c7_rf_chdad_reg[13]/NET0131  & ~n8949 ;
  assign n9345 = n8949 & ~n9018 ;
  assign n9346 = ~n9017 & n9345 ;
  assign n9347 = ~n9344 & ~n9346 ;
  assign n9348 = ~\ctl_rf_c7_rf_chdad_reg[14]/NET0131  & ~n8949 ;
  assign n9349 = n8949 & ~n9027 ;
  assign n9350 = ~n9026 & n9349 ;
  assign n9351 = ~n9348 & ~n9350 ;
  assign n9352 = ~\ctl_rf_c7_rf_chdad_reg[1]/NET0131  & ~n9339 ;
  assign n9353 = ~n8992 & n9339 ;
  assign n9354 = ~n8991 & n9353 ;
  assign n9355 = ~n9352 & ~n9354 ;
  assign n9356 = ~\ctl_rf_c7_rf_chdad_reg[2]/NET0131  & ~n9339 ;
  assign n9357 = ~n9001 & n9339 ;
  assign n9358 = ~n9000 & n9357 ;
  assign n9359 = ~n9356 & ~n9358 ;
  assign n9360 = ~\ctl_rf_c7_rf_chsad_reg[0]/NET0131  & ~n8672 ;
  assign n9361 = ~n3771 & n8672 ;
  assign n9362 = ~n3770 & n9361 ;
  assign n9363 = ~n9360 & ~n9362 ;
  assign n9364 = ~\ctl_rf_c7_rf_chsad_reg[1]/NET0131  & ~n8672 ;
  assign n9365 = n8672 & ~n8992 ;
  assign n9366 = ~n8991 & n9365 ;
  assign n9367 = ~n9364 & ~n9366 ;
  assign n9368 = ~\ctl_rf_c7_rf_chsad_reg[2]/NET0131  & ~n8672 ;
  assign n9369 = n8672 & ~n9001 ;
  assign n9370 = ~n9000 & n9369 ;
  assign n9371 = ~n9368 & ~n9370 ;
  assign n9372 = ~\ctl_rf_c7_rf_chsad_reg[3]/NET0131  & ~n8672 ;
  assign n9373 = n8672 & ~n9044 ;
  assign n9374 = ~n9043 & n9373 ;
  assign n9375 = ~n9372 & ~n9374 ;
  assign n9376 = ~\ctl_rf_c7_rf_chsad_reg[4]/NET0131  & ~n8672 ;
  assign n9377 = n8672 & ~n8714 ;
  assign n9378 = ~n8713 & n9377 ;
  assign n9379 = ~n9376 & ~n9378 ;
  assign n9380 = ~\ctl_rf_c0_rf_chdad_reg[0]/NET0131  & ~n9134 ;
  assign n9381 = ~n3771 & n9134 ;
  assign n9382 = ~n3770 & n9381 ;
  assign n9383 = ~n9380 & ~n9382 ;
  assign n9384 = ~\ctl_rf_c0_rf_chdad_reg[11]/NET0131  & ~n9143 ;
  assign n9385 = ~n8791 & n9143 ;
  assign n9386 = ~n8790 & n9385 ;
  assign n9387 = ~n9384 & ~n9386 ;
  assign n9388 = ~\ctl_rf_c0_rf_chdad_reg[12]/NET0131  & ~n9143 ;
  assign n9389 = ~n8768 & n9143 ;
  assign n9390 = ~n8767 & n9389 ;
  assign n9391 = ~n9388 & ~n9390 ;
  assign n9392 = ~\ctl_rf_c0_rf_chdad_reg[14]/NET0131  & ~n9143 ;
  assign n9393 = ~n9027 & n9143 ;
  assign n9394 = ~n9026 & n9393 ;
  assign n9395 = ~n9392 & ~n9394 ;
  assign n9396 = ~\ctl_rf_c0_rf_chdad_reg[15]/NET0131  & ~n9143 ;
  assign n9397 = ~n3763 & n9143 ;
  assign n9398 = ~n3762 & n9397 ;
  assign n9399 = ~n9396 & ~n9398 ;
  assign n9400 = \m1_mux_hrp_df_reg[0]/NET0131  & n2830 ;
  assign n9401 = \m1_mux_hrp_df_reg[0]/NET0131  & n2764 ;
  assign n9402 = n2798 & n9401 ;
  assign n9403 = ~n9400 & ~n9402 ;
  assign n9404 = ~\ctl_rf_c4dmabs_reg[16]/NET0131  & \ctl_rf_c4dmabs_reg[22]/NET0131  ;
  assign n9405 = \ctl_rf_c4dmabs_reg[17]/NET0131  & ~n9404 ;
  assign n9406 = ~\ctl_rf_c4dmabs_reg[16]/NET0131  & \ctl_rf_c4dmabs_reg[20]/NET0131  ;
  assign n9407 = ~\ctl_rf_c4dmabs_reg[21]/NET0131  & ~\ctl_rf_c4dmabs_reg[22]/NET0131  ;
  assign n9408 = ~n9406 & n9407 ;
  assign n9409 = ~n9405 & ~n9408 ;
  assign n9410 = ~\ctl_rf_c4dmabs_reg[23]/NET0131  & ~n9409 ;
  assign n9411 = ~\ctl_rf_c4dmabs_reg[18]/NET0131  & ~\ctl_rf_c4dmabs_reg[19]/NET0131  ;
  assign n9412 = ~n9410 & n9411 ;
  assign n9413 = ~\ctl_rf_c4dmabs_reg[28]/NET0131  & ~\ctl_rf_c4dmabs_reg[29]/NET0131  ;
  assign n9414 = ~\ctl_rf_c4dmabs_reg[30]/NET0131  & ~\ctl_rf_c4dmabs_reg[31]/NET0131  ;
  assign n9415 = n9413 & n9414 ;
  assign n9416 = ~\ctl_rf_c4dmabs_reg[24]/NET0131  & ~\ctl_rf_c4dmabs_reg[25]/NET0131  ;
  assign n9417 = ~\ctl_rf_c4dmabs_reg[26]/NET0131  & ~\ctl_rf_c4dmabs_reg[27]/NET0131  ;
  assign n9418 = n9416 & n9417 ;
  assign n9419 = n9415 & n9418 ;
  assign n9420 = ~n9412 & n9419 ;
  assign n9421 = ~\ctl_rf_c6dmabs_reg[16]/NET0131  & \ctl_rf_c6dmabs_reg[22]/NET0131  ;
  assign n9422 = \ctl_rf_c6dmabs_reg[17]/NET0131  & ~n9421 ;
  assign n9423 = ~\ctl_rf_c6dmabs_reg[16]/NET0131  & \ctl_rf_c6dmabs_reg[20]/NET0131  ;
  assign n9424 = ~\ctl_rf_c6dmabs_reg[21]/NET0131  & ~\ctl_rf_c6dmabs_reg[22]/NET0131  ;
  assign n9425 = ~n9423 & n9424 ;
  assign n9426 = ~n9422 & ~n9425 ;
  assign n9427 = ~\ctl_rf_c6dmabs_reg[23]/NET0131  & ~n9426 ;
  assign n9428 = ~\ctl_rf_c6dmabs_reg[18]/NET0131  & ~\ctl_rf_c6dmabs_reg[19]/NET0131  ;
  assign n9429 = ~n9427 & n9428 ;
  assign n9430 = ~\ctl_rf_c6dmabs_reg[28]/NET0131  & ~\ctl_rf_c6dmabs_reg[29]/NET0131  ;
  assign n9431 = ~\ctl_rf_c6dmabs_reg[30]/NET0131  & ~\ctl_rf_c6dmabs_reg[31]/NET0131  ;
  assign n9432 = n9430 & n9431 ;
  assign n9433 = ~\ctl_rf_c6dmabs_reg[24]/NET0131  & ~\ctl_rf_c6dmabs_reg[25]/NET0131  ;
  assign n9434 = ~\ctl_rf_c6dmabs_reg[26]/NET0131  & ~\ctl_rf_c6dmabs_reg[27]/NET0131  ;
  assign n9435 = n9433 & n9434 ;
  assign n9436 = n9432 & n9435 ;
  assign n9437 = ~n9429 & n9436 ;
  assign n9438 = ~n9420 & ~n9437 ;
  assign n9439 = ~\ctl_rf_c3dmabs_reg[16]/NET0131  & \ctl_rf_c3dmabs_reg[22]/NET0131  ;
  assign n9440 = \ctl_rf_c3dmabs_reg[17]/NET0131  & ~n9439 ;
  assign n9441 = ~\ctl_rf_c3dmabs_reg[16]/NET0131  & \ctl_rf_c3dmabs_reg[20]/NET0131  ;
  assign n9442 = ~\ctl_rf_c3dmabs_reg[21]/NET0131  & ~\ctl_rf_c3dmabs_reg[22]/NET0131  ;
  assign n9443 = ~n9441 & n9442 ;
  assign n9444 = ~n9440 & ~n9443 ;
  assign n9445 = ~\ctl_rf_c3dmabs_reg[23]/NET0131  & ~n9444 ;
  assign n9446 = ~\ctl_rf_c3dmabs_reg[18]/NET0131  & ~\ctl_rf_c3dmabs_reg[19]/NET0131  ;
  assign n9447 = ~n9445 & n9446 ;
  assign n9448 = ~\ctl_rf_c3dmabs_reg[28]/NET0131  & ~\ctl_rf_c3dmabs_reg[29]/NET0131  ;
  assign n9449 = ~\ctl_rf_c3dmabs_reg[30]/NET0131  & ~\ctl_rf_c3dmabs_reg[31]/NET0131  ;
  assign n9450 = n9448 & n9449 ;
  assign n9451 = ~\ctl_rf_c3dmabs_reg[24]/NET0131  & ~\ctl_rf_c3dmabs_reg[25]/NET0131  ;
  assign n9452 = ~\ctl_rf_c3dmabs_reg[26]/NET0131  & ~\ctl_rf_c3dmabs_reg[27]/NET0131  ;
  assign n9453 = n9451 & n9452 ;
  assign n9454 = n9450 & n9453 ;
  assign n9455 = ~n9447 & n9454 ;
  assign n9456 = n9438 & ~n9455 ;
  assign n9457 = ~\ctl_rf_c5dmabs_reg[16]/NET0131  & \ctl_rf_c5dmabs_reg[22]/NET0131  ;
  assign n9458 = \ctl_rf_c5dmabs_reg[17]/NET0131  & ~n9457 ;
  assign n9459 = ~\ctl_rf_c5dmabs_reg[16]/NET0131  & \ctl_rf_c5dmabs_reg[20]/NET0131  ;
  assign n9460 = ~\ctl_rf_c5dmabs_reg[21]/NET0131  & ~\ctl_rf_c5dmabs_reg[22]/NET0131  ;
  assign n9461 = ~n9459 & n9460 ;
  assign n9462 = ~n9458 & ~n9461 ;
  assign n9463 = ~\ctl_rf_c5dmabs_reg[23]/NET0131  & ~n9462 ;
  assign n9464 = ~\ctl_rf_c5dmabs_reg[18]/NET0131  & ~\ctl_rf_c5dmabs_reg[19]/NET0131  ;
  assign n9465 = ~n9463 & n9464 ;
  assign n9466 = ~\ctl_rf_c5dmabs_reg[28]/NET0131  & ~\ctl_rf_c5dmabs_reg[29]/NET0131  ;
  assign n9467 = ~\ctl_rf_c5dmabs_reg[30]/NET0131  & ~\ctl_rf_c5dmabs_reg[31]/NET0131  ;
  assign n9468 = n9466 & n9467 ;
  assign n9469 = ~\ctl_rf_c5dmabs_reg[24]/NET0131  & ~\ctl_rf_c5dmabs_reg[25]/NET0131  ;
  assign n9470 = ~\ctl_rf_c5dmabs_reg[26]/NET0131  & ~\ctl_rf_c5dmabs_reg[27]/NET0131  ;
  assign n9471 = n9469 & n9470 ;
  assign n9472 = n9468 & n9471 ;
  assign n9473 = ~n9465 & n9472 ;
  assign n9474 = ~\ctl_rf_c7dmabs_reg[16]/NET0131  & \ctl_rf_c7dmabs_reg[22]/NET0131  ;
  assign n9475 = \ctl_rf_c7dmabs_reg[17]/NET0131  & ~n9474 ;
  assign n9476 = ~\ctl_rf_c7dmabs_reg[16]/NET0131  & \ctl_rf_c7dmabs_reg[20]/NET0131  ;
  assign n9477 = ~\ctl_rf_c7dmabs_reg[21]/NET0131  & ~\ctl_rf_c7dmabs_reg[22]/NET0131  ;
  assign n9478 = ~n9476 & n9477 ;
  assign n9479 = ~n9475 & ~n9478 ;
  assign n9480 = ~\ctl_rf_c7dmabs_reg[23]/NET0131  & ~n9479 ;
  assign n9481 = ~\ctl_rf_c7dmabs_reg[18]/NET0131  & ~\ctl_rf_c7dmabs_reg[19]/NET0131  ;
  assign n9482 = ~n9480 & n9481 ;
  assign n9483 = ~\ctl_rf_c7dmabs_reg[28]/NET0131  & ~\ctl_rf_c7dmabs_reg[29]/NET0131  ;
  assign n9484 = ~\ctl_rf_c7dmabs_reg[30]/NET0131  & ~\ctl_rf_c7dmabs_reg[31]/NET0131  ;
  assign n9485 = n9483 & n9484 ;
  assign n9486 = ~\ctl_rf_c7dmabs_reg[24]/NET0131  & ~\ctl_rf_c7dmabs_reg[25]/NET0131  ;
  assign n9487 = ~\ctl_rf_c7dmabs_reg[26]/NET0131  & ~\ctl_rf_c7dmabs_reg[27]/NET0131  ;
  assign n9488 = n9486 & n9487 ;
  assign n9489 = n9485 & n9488 ;
  assign n9490 = ~n9482 & n9489 ;
  assign n9491 = ~n9473 & ~n9490 ;
  assign n9492 = ~\ctl_rf_c2dmabs_reg[16]/NET0131  & \ctl_rf_c2dmabs_reg[22]/NET0131  ;
  assign n9493 = \ctl_rf_c2dmabs_reg[17]/NET0131  & ~n9492 ;
  assign n9494 = ~\ctl_rf_c2dmabs_reg[16]/NET0131  & \ctl_rf_c2dmabs_reg[20]/NET0131  ;
  assign n9495 = ~\ctl_rf_c2dmabs_reg[21]/NET0131  & ~\ctl_rf_c2dmabs_reg[22]/NET0131  ;
  assign n9496 = ~n9494 & n9495 ;
  assign n9497 = ~n9493 & ~n9496 ;
  assign n9498 = ~\ctl_rf_c2dmabs_reg[23]/NET0131  & ~n9497 ;
  assign n9499 = ~\ctl_rf_c2dmabs_reg[18]/NET0131  & ~\ctl_rf_c2dmabs_reg[19]/NET0131  ;
  assign n9500 = ~n9498 & n9499 ;
  assign n9501 = ~\ctl_rf_c2dmabs_reg[28]/NET0131  & ~\ctl_rf_c2dmabs_reg[29]/NET0131  ;
  assign n9502 = ~\ctl_rf_c2dmabs_reg[30]/NET0131  & ~\ctl_rf_c2dmabs_reg[31]/NET0131  ;
  assign n9503 = n9501 & n9502 ;
  assign n9504 = ~\ctl_rf_c2dmabs_reg[24]/NET0131  & ~\ctl_rf_c2dmabs_reg[25]/NET0131  ;
  assign n9505 = ~\ctl_rf_c2dmabs_reg[26]/NET0131  & ~\ctl_rf_c2dmabs_reg[27]/NET0131  ;
  assign n9506 = n9504 & n9505 ;
  assign n9507 = n9503 & n9506 ;
  assign n9508 = ~n9500 & n9507 ;
  assign n9509 = ~\ctl_rf_c1dmabs_reg[16]/NET0131  & \ctl_rf_c1dmabs_reg[22]/NET0131  ;
  assign n9510 = \ctl_rf_c1dmabs_reg[17]/NET0131  & ~n9509 ;
  assign n9511 = ~\ctl_rf_c1dmabs_reg[16]/NET0131  & \ctl_rf_c1dmabs_reg[20]/NET0131  ;
  assign n9512 = ~\ctl_rf_c1dmabs_reg[21]/NET0131  & ~\ctl_rf_c1dmabs_reg[22]/NET0131  ;
  assign n9513 = ~n9511 & n9512 ;
  assign n9514 = ~n9510 & ~n9513 ;
  assign n9515 = ~\ctl_rf_c1dmabs_reg[23]/NET0131  & ~n9514 ;
  assign n9516 = ~\ctl_rf_c1dmabs_reg[18]/NET0131  & ~\ctl_rf_c1dmabs_reg[19]/NET0131  ;
  assign n9517 = ~n9515 & n9516 ;
  assign n9518 = ~\ctl_rf_c1dmabs_reg[28]/NET0131  & ~\ctl_rf_c1dmabs_reg[29]/NET0131  ;
  assign n9519 = ~\ctl_rf_c1dmabs_reg[30]/NET0131  & ~\ctl_rf_c1dmabs_reg[31]/NET0131  ;
  assign n9520 = n9518 & n9519 ;
  assign n9521 = ~\ctl_rf_c1dmabs_reg[24]/NET0131  & ~\ctl_rf_c1dmabs_reg[25]/NET0131  ;
  assign n9522 = ~\ctl_rf_c1dmabs_reg[26]/NET0131  & ~\ctl_rf_c1dmabs_reg[27]/NET0131  ;
  assign n9523 = n9521 & n9522 ;
  assign n9524 = n9520 & n9523 ;
  assign n9525 = ~n9517 & n9524 ;
  assign n9526 = ~n9508 & ~n9525 ;
  assign n9527 = n9491 & n9526 ;
  assign n9528 = n9456 & n9527 ;
  assign n9529 = ~\ctl_rf_c0dmabs_reg[16]/NET0131  & \ctl_rf_c0dmabs_reg[22]/NET0131  ;
  assign n9530 = \ctl_rf_c0dmabs_reg[17]/NET0131  & ~n9529 ;
  assign n9531 = ~\ctl_rf_c0dmabs_reg[16]/NET0131  & \ctl_rf_c0dmabs_reg[20]/NET0131  ;
  assign n9532 = ~\ctl_rf_c0dmabs_reg[21]/NET0131  & ~\ctl_rf_c0dmabs_reg[22]/NET0131  ;
  assign n9533 = ~n9531 & n9532 ;
  assign n9534 = ~n9530 & ~n9533 ;
  assign n9535 = ~\ctl_rf_c0dmabs_reg[23]/NET0131  & ~n9534 ;
  assign n9536 = ~\ctl_rf_c0dmabs_reg[18]/NET0131  & ~\ctl_rf_c0dmabs_reg[19]/NET0131  ;
  assign n9537 = ~n9535 & n9536 ;
  assign n9538 = ~\ctl_rf_c0dmabs_reg[28]/NET0131  & ~\ctl_rf_c0dmabs_reg[29]/NET0131  ;
  assign n9539 = ~\ctl_rf_c0dmabs_reg[30]/NET0131  & ~\ctl_rf_c0dmabs_reg[31]/NET0131  ;
  assign n9540 = n9538 & n9539 ;
  assign n9541 = ~\ctl_rf_c0dmabs_reg[24]/NET0131  & ~\ctl_rf_c0dmabs_reg[25]/NET0131  ;
  assign n9542 = ~\ctl_rf_c0dmabs_reg[26]/NET0131  & ~\ctl_rf_c0dmabs_reg[27]/NET0131  ;
  assign n9543 = n9541 & n9542 ;
  assign n9544 = n9540 & n9543 ;
  assign n9545 = ~n9537 & n9544 ;
  assign n9546 = ~\ctl_rf_c0brbs_reg[16]/NET0131  & \ctl_rf_c0brbs_reg[22]/NET0131  ;
  assign n9547 = \ctl_rf_c0brbs_reg[17]/NET0131  & ~n9546 ;
  assign n9548 = ~\ctl_rf_c0brbs_reg[16]/NET0131  & \ctl_rf_c0brbs_reg[20]/NET0131  ;
  assign n9549 = ~\ctl_rf_c0brbs_reg[21]/NET0131  & ~\ctl_rf_c0brbs_reg[22]/NET0131  ;
  assign n9550 = ~n9548 & n9549 ;
  assign n9551 = ~n9547 & ~n9550 ;
  assign n9552 = ~\ctl_rf_c0brbs_reg[23]/NET0131  & ~n9551 ;
  assign n9553 = ~\ctl_rf_c0brbs_reg[18]/NET0131  & ~\ctl_rf_c0brbs_reg[19]/NET0131  ;
  assign n9554 = ~n9552 & n9553 ;
  assign n9555 = ~\ctl_rf_c0brbs_reg[28]/NET0131  & ~\ctl_rf_c0brbs_reg[29]/NET0131  ;
  assign n9556 = ~\ctl_rf_c0brbs_reg[30]/NET0131  & ~\ctl_rf_c0brbs_reg[31]/NET0131  ;
  assign n9557 = n9555 & n9556 ;
  assign n9558 = ~\ctl_rf_c0brbs_reg[24]/NET0131  & ~\ctl_rf_c0brbs_reg[25]/NET0131  ;
  assign n9559 = ~\ctl_rf_c0brbs_reg[26]/NET0131  & ~\ctl_rf_c0brbs_reg[27]/NET0131  ;
  assign n9560 = n9558 & n9559 ;
  assign n9561 = n9557 & n9560 ;
  assign n9562 = ~n9554 & n9561 ;
  assign n9563 = ~n9545 & ~n9562 ;
  assign n9564 = ~\ctl_rf_c1brbs_reg[16]/NET0131  & \ctl_rf_c1brbs_reg[22]/NET0131  ;
  assign n9565 = \ctl_rf_c1brbs_reg[17]/NET0131  & ~n9564 ;
  assign n9566 = ~\ctl_rf_c1brbs_reg[16]/NET0131  & \ctl_rf_c1brbs_reg[20]/NET0131  ;
  assign n9567 = ~\ctl_rf_c1brbs_reg[21]/NET0131  & ~\ctl_rf_c1brbs_reg[22]/NET0131  ;
  assign n9568 = ~n9566 & n9567 ;
  assign n9569 = ~n9565 & ~n9568 ;
  assign n9570 = ~\ctl_rf_c1brbs_reg[23]/NET0131  & ~n9569 ;
  assign n9571 = ~\ctl_rf_c1brbs_reg[18]/NET0131  & ~\ctl_rf_c1brbs_reg[19]/NET0131  ;
  assign n9572 = ~n9570 & n9571 ;
  assign n9573 = ~\ctl_rf_c1brbs_reg[28]/NET0131  & ~\ctl_rf_c1brbs_reg[29]/NET0131  ;
  assign n9574 = ~\ctl_rf_c1brbs_reg[30]/NET0131  & ~\ctl_rf_c1brbs_reg[31]/NET0131  ;
  assign n9575 = n9573 & n9574 ;
  assign n9576 = ~\ctl_rf_c1brbs_reg[24]/NET0131  & ~\ctl_rf_c1brbs_reg[25]/NET0131  ;
  assign n9577 = ~\ctl_rf_c1brbs_reg[26]/NET0131  & ~\ctl_rf_c1brbs_reg[27]/NET0131  ;
  assign n9578 = n9576 & n9577 ;
  assign n9579 = n9575 & n9578 ;
  assign n9580 = ~n9572 & n9579 ;
  assign n9581 = ~\ctl_rf_c2brbs_reg[16]/NET0131  & \ctl_rf_c2brbs_reg[22]/NET0131  ;
  assign n9582 = \ctl_rf_c2brbs_reg[17]/NET0131  & ~n9581 ;
  assign n9583 = ~\ctl_rf_c2brbs_reg[16]/NET0131  & \ctl_rf_c2brbs_reg[20]/NET0131  ;
  assign n9584 = ~\ctl_rf_c2brbs_reg[21]/NET0131  & ~\ctl_rf_c2brbs_reg[22]/NET0131  ;
  assign n9585 = ~n9583 & n9584 ;
  assign n9586 = ~n9582 & ~n9585 ;
  assign n9587 = ~\ctl_rf_c2brbs_reg[23]/NET0131  & ~n9586 ;
  assign n9588 = ~\ctl_rf_c2brbs_reg[18]/NET0131  & ~\ctl_rf_c2brbs_reg[19]/NET0131  ;
  assign n9589 = ~n9587 & n9588 ;
  assign n9590 = ~\ctl_rf_c2brbs_reg[28]/NET0131  & ~\ctl_rf_c2brbs_reg[29]/NET0131  ;
  assign n9591 = ~\ctl_rf_c2brbs_reg[30]/NET0131  & ~\ctl_rf_c2brbs_reg[31]/NET0131  ;
  assign n9592 = n9590 & n9591 ;
  assign n9593 = ~\ctl_rf_c2brbs_reg[24]/NET0131  & ~\ctl_rf_c2brbs_reg[25]/NET0131  ;
  assign n9594 = ~\ctl_rf_c2brbs_reg[26]/NET0131  & ~\ctl_rf_c2brbs_reg[27]/NET0131  ;
  assign n9595 = n9593 & n9594 ;
  assign n9596 = n9592 & n9595 ;
  assign n9597 = ~n9589 & n9596 ;
  assign n9598 = ~n9580 & ~n9597 ;
  assign n9599 = n9563 & n9598 ;
  assign n9600 = n9528 & n9599 ;
  assign n9601 = ~n2799 & ~n2830 ;
  assign n9602 = ~\ctl_rf_c6brbs_reg[16]/NET0131  & \ctl_rf_c6brbs_reg[22]/NET0131  ;
  assign n9603 = \ctl_rf_c6brbs_reg[17]/NET0131  & ~n9602 ;
  assign n9604 = ~\ctl_rf_c6brbs_reg[16]/NET0131  & \ctl_rf_c6brbs_reg[20]/NET0131  ;
  assign n9605 = ~\ctl_rf_c6brbs_reg[21]/NET0131  & ~\ctl_rf_c6brbs_reg[22]/NET0131  ;
  assign n9606 = ~n9604 & n9605 ;
  assign n9607 = ~n9603 & ~n9606 ;
  assign n9608 = ~\ctl_rf_c6brbs_reg[23]/NET0131  & ~n9607 ;
  assign n9609 = ~\ctl_rf_c6brbs_reg[18]/NET0131  & ~\ctl_rf_c6brbs_reg[19]/NET0131  ;
  assign n9610 = ~n9608 & n9609 ;
  assign n9611 = ~\ctl_rf_c6brbs_reg[28]/NET0131  & ~\ctl_rf_c6brbs_reg[29]/NET0131  ;
  assign n9612 = ~\ctl_rf_c6brbs_reg[30]/NET0131  & ~\ctl_rf_c6brbs_reg[31]/NET0131  ;
  assign n9613 = n9611 & n9612 ;
  assign n9614 = ~\ctl_rf_c6brbs_reg[24]/NET0131  & ~\ctl_rf_c6brbs_reg[25]/NET0131  ;
  assign n9615 = ~\ctl_rf_c6brbs_reg[26]/NET0131  & ~\ctl_rf_c6brbs_reg[27]/NET0131  ;
  assign n9616 = n9614 & n9615 ;
  assign n9617 = n9613 & n9616 ;
  assign n9618 = ~n9610 & n9617 ;
  assign n9619 = ~\ctl_rf_c7brbs_reg[16]/NET0131  & \ctl_rf_c7brbs_reg[22]/NET0131  ;
  assign n9620 = \ctl_rf_c7brbs_reg[17]/NET0131  & ~n9619 ;
  assign n9621 = ~\ctl_rf_c7brbs_reg[16]/NET0131  & \ctl_rf_c7brbs_reg[20]/NET0131  ;
  assign n9622 = ~\ctl_rf_c7brbs_reg[21]/NET0131  & ~\ctl_rf_c7brbs_reg[22]/NET0131  ;
  assign n9623 = ~n9621 & n9622 ;
  assign n9624 = ~n9620 & ~n9623 ;
  assign n9625 = ~\ctl_rf_c7brbs_reg[23]/NET0131  & ~n9624 ;
  assign n9626 = ~\ctl_rf_c7brbs_reg[18]/NET0131  & ~\ctl_rf_c7brbs_reg[19]/NET0131  ;
  assign n9627 = ~n9625 & n9626 ;
  assign n9628 = ~\ctl_rf_c7brbs_reg[28]/NET0131  & ~\ctl_rf_c7brbs_reg[29]/NET0131  ;
  assign n9629 = ~\ctl_rf_c7brbs_reg[30]/NET0131  & ~\ctl_rf_c7brbs_reg[31]/NET0131  ;
  assign n9630 = n9628 & n9629 ;
  assign n9631 = ~\ctl_rf_c7brbs_reg[24]/NET0131  & ~\ctl_rf_c7brbs_reg[25]/NET0131  ;
  assign n9632 = ~\ctl_rf_c7brbs_reg[26]/NET0131  & ~\ctl_rf_c7brbs_reg[27]/NET0131  ;
  assign n9633 = n9631 & n9632 ;
  assign n9634 = n9630 & n9633 ;
  assign n9635 = ~n9627 & n9634 ;
  assign n9636 = ~n9618 & ~n9635 ;
  assign n9637 = ~\ctl_rf_c5brbs_reg[16]/NET0131  & \ctl_rf_c5brbs_reg[22]/NET0131  ;
  assign n9638 = \ctl_rf_c5brbs_reg[17]/NET0131  & ~n9637 ;
  assign n9639 = ~\ctl_rf_c5brbs_reg[16]/NET0131  & \ctl_rf_c5brbs_reg[20]/NET0131  ;
  assign n9640 = ~\ctl_rf_c5brbs_reg[21]/NET0131  & ~\ctl_rf_c5brbs_reg[22]/NET0131  ;
  assign n9641 = ~n9639 & n9640 ;
  assign n9642 = ~n9638 & ~n9641 ;
  assign n9643 = ~\ctl_rf_c5brbs_reg[23]/NET0131  & ~n9642 ;
  assign n9644 = ~\ctl_rf_c5brbs_reg[18]/NET0131  & ~\ctl_rf_c5brbs_reg[19]/NET0131  ;
  assign n9645 = ~n9643 & n9644 ;
  assign n9646 = ~\ctl_rf_c5brbs_reg[28]/NET0131  & ~\ctl_rf_c5brbs_reg[29]/NET0131  ;
  assign n9647 = ~\ctl_rf_c5brbs_reg[30]/NET0131  & ~\ctl_rf_c5brbs_reg[31]/NET0131  ;
  assign n9648 = n9646 & n9647 ;
  assign n9649 = ~\ctl_rf_c5brbs_reg[24]/NET0131  & ~\ctl_rf_c5brbs_reg[25]/NET0131  ;
  assign n9650 = ~\ctl_rf_c5brbs_reg[26]/NET0131  & ~\ctl_rf_c5brbs_reg[27]/NET0131  ;
  assign n9651 = n9649 & n9650 ;
  assign n9652 = n9648 & n9651 ;
  assign n9653 = ~n9645 & n9652 ;
  assign n9654 = n9636 & ~n9653 ;
  assign n9655 = ~\ctl_rf_c3brbs_reg[16]/NET0131  & \ctl_rf_c3brbs_reg[22]/NET0131  ;
  assign n9656 = \ctl_rf_c3brbs_reg[17]/NET0131  & ~n9655 ;
  assign n9657 = ~\ctl_rf_c3brbs_reg[16]/NET0131  & \ctl_rf_c3brbs_reg[20]/NET0131  ;
  assign n9658 = ~\ctl_rf_c3brbs_reg[21]/NET0131  & ~\ctl_rf_c3brbs_reg[22]/NET0131  ;
  assign n9659 = ~n9657 & n9658 ;
  assign n9660 = ~n9656 & ~n9659 ;
  assign n9661 = ~\ctl_rf_c3brbs_reg[23]/NET0131  & ~n9660 ;
  assign n9662 = ~\ctl_rf_c3brbs_reg[18]/NET0131  & ~\ctl_rf_c3brbs_reg[19]/NET0131  ;
  assign n9663 = ~n9661 & n9662 ;
  assign n9664 = ~\ctl_rf_c3brbs_reg[28]/NET0131  & ~\ctl_rf_c3brbs_reg[29]/NET0131  ;
  assign n9665 = ~\ctl_rf_c3brbs_reg[30]/NET0131  & ~\ctl_rf_c3brbs_reg[31]/NET0131  ;
  assign n9666 = n9664 & n9665 ;
  assign n9667 = ~\ctl_rf_c3brbs_reg[24]/NET0131  & ~\ctl_rf_c3brbs_reg[25]/NET0131  ;
  assign n9668 = ~\ctl_rf_c3brbs_reg[26]/NET0131  & ~\ctl_rf_c3brbs_reg[27]/NET0131  ;
  assign n9669 = n9667 & n9668 ;
  assign n9670 = n9666 & n9669 ;
  assign n9671 = ~n9663 & n9670 ;
  assign n9672 = ~\ctl_rf_c4brbs_reg[16]/NET0131  & \ctl_rf_c4brbs_reg[22]/NET0131  ;
  assign n9673 = \ctl_rf_c4brbs_reg[17]/NET0131  & ~n9672 ;
  assign n9674 = ~\ctl_rf_c4brbs_reg[16]/NET0131  & \ctl_rf_c4brbs_reg[20]/NET0131  ;
  assign n9675 = ~\ctl_rf_c4brbs_reg[21]/NET0131  & ~\ctl_rf_c4brbs_reg[22]/NET0131  ;
  assign n9676 = ~n9674 & n9675 ;
  assign n9677 = ~n9673 & ~n9676 ;
  assign n9678 = ~\ctl_rf_c4brbs_reg[23]/NET0131  & ~n9677 ;
  assign n9679 = ~\ctl_rf_c4brbs_reg[18]/NET0131  & ~\ctl_rf_c4brbs_reg[19]/NET0131  ;
  assign n9680 = ~n9678 & n9679 ;
  assign n9681 = ~\ctl_rf_c4brbs_reg[28]/NET0131  & ~\ctl_rf_c4brbs_reg[29]/NET0131  ;
  assign n9682 = ~\ctl_rf_c4brbs_reg[30]/NET0131  & ~\ctl_rf_c4brbs_reg[31]/NET0131  ;
  assign n9683 = n9681 & n9682 ;
  assign n9684 = ~\ctl_rf_c4brbs_reg[24]/NET0131  & ~\ctl_rf_c4brbs_reg[25]/NET0131  ;
  assign n9685 = ~\ctl_rf_c4brbs_reg[26]/NET0131  & ~\ctl_rf_c4brbs_reg[27]/NET0131  ;
  assign n9686 = n9684 & n9685 ;
  assign n9687 = n9683 & n9686 ;
  assign n9688 = ~n9680 & n9687 ;
  assign n9689 = ~n9671 & ~n9688 ;
  assign n9690 = n9654 & n9689 ;
  assign n9691 = n9601 & n9690 ;
  assign n9692 = n9600 & n9691 ;
  assign n9693 = ~n2846 & n9692 ;
  assign n9694 = n9403 & ~n9693 ;
  assign n9695 = n9528 & n9563 ;
  assign n9696 = n9671 & ~n9688 ;
  assign n9697 = n9654 & n9696 ;
  assign n9698 = n9598 & n9697 ;
  assign n9699 = n9636 & n9653 ;
  assign n9700 = ~n9618 & n9635 ;
  assign n9701 = ~n9653 & n9700 ;
  assign n9702 = ~n9699 & ~n9701 ;
  assign n9703 = n9598 & n9689 ;
  assign n9704 = ~n9702 & n9703 ;
  assign n9705 = ~n9698 & ~n9704 ;
  assign n9706 = n9580 & ~n9597 ;
  assign n9707 = n9689 & n9706 ;
  assign n9708 = n9654 & n9707 ;
  assign n9709 = n9705 & ~n9708 ;
  assign n9710 = n9695 & ~n9709 ;
  assign n9711 = n9438 & n9455 ;
  assign n9712 = n9491 & n9711 ;
  assign n9713 = n9473 & n9490 ;
  assign n9714 = ~n9491 & ~n9713 ;
  assign n9715 = n9456 & n9714 ;
  assign n9716 = ~n9525 & ~n9715 ;
  assign n9717 = ~n9712 & n9716 ;
  assign n9718 = ~n9528 & ~n9545 ;
  assign n9719 = n9491 & ~n9508 ;
  assign n9720 = n9456 & n9719 ;
  assign n9721 = ~n9526 & ~n9720 ;
  assign n9722 = n9718 & ~n9721 ;
  assign n9723 = ~n9717 & n9722 ;
  assign n9724 = ~n9710 & ~n9723 ;
  assign n9725 = n2230 & n2232 ;
  assign n9726 = \ctl_rf_be_d1_reg[1]/P0001  & n9725 ;
  assign n9727 = n8578 & n9726 ;
  assign n9728 = ~\ctl_rf_c1_rf_chllp_reg[10]/NET0131  & ~n9727 ;
  assign n9729 = ~n8759 & n9727 ;
  assign n9730 = ~n8758 & n9729 ;
  assign n9731 = ~n9728 & ~n9730 ;
  assign n9732 = ~\ctl_rf_c1_rf_chllp_reg[11]/NET0131  & ~n9727 ;
  assign n9733 = ~n8791 & n9727 ;
  assign n9734 = ~n8790 & n9733 ;
  assign n9735 = ~n9732 & ~n9734 ;
  assign n9736 = ~\ctl_rf_c1_rf_chllp_reg[12]/NET0131  & ~n9727 ;
  assign n9737 = ~n8768 & n9727 ;
  assign n9738 = ~n8767 & n9737 ;
  assign n9739 = ~n9736 & ~n9738 ;
  assign n9740 = ~\ctl_rf_c1_rf_chllp_reg[13]/NET0131  & ~n9727 ;
  assign n9741 = ~n9018 & n9727 ;
  assign n9742 = ~n9017 & n9741 ;
  assign n9743 = ~n9740 & ~n9742 ;
  assign n9744 = ~\ctl_rf_c1_rf_chllp_reg[14]/NET0131  & ~n9727 ;
  assign n9745 = ~n9027 & n9727 ;
  assign n9746 = ~n9026 & n9745 ;
  assign n9747 = ~n9744 & ~n9746 ;
  assign n9748 = ~\ctl_rf_c1_rf_chllp_reg[15]/NET0131  & ~n9727 ;
  assign n9749 = ~n3763 & n9727 ;
  assign n9750 = ~n3762 & n9749 ;
  assign n9751 = ~n9748 & ~n9750 ;
  assign n9752 = \ctl_rf_be_d1_reg[2]/P0001  & n9725 ;
  assign n9753 = n8578 & n9752 ;
  assign n9754 = ~\ctl_rf_c1_rf_chllp_reg[16]/NET0131  & ~n9753 ;
  assign n9755 = ~n2680 & n9753 ;
  assign n9756 = ~n2679 & n9755 ;
  assign n9757 = ~n9754 & ~n9756 ;
  assign n9758 = ~\ctl_rf_c1_rf_chllp_reg[17]/NET0131  & ~n9753 ;
  assign n9759 = ~n2260 & n9753 ;
  assign n9760 = ~n2259 & n9759 ;
  assign n9761 = ~n9758 & ~n9760 ;
  assign n9762 = ~\ctl_rf_c1_rf_chllp_reg[18]/NET0131  & ~n9753 ;
  assign n9763 = ~n2400 & n9753 ;
  assign n9764 = ~n2399 & n9763 ;
  assign n9765 = ~n9762 & ~n9764 ;
  assign n9766 = ~\ctl_rf_c1_rf_chllp_reg[19]/NET0131  & ~n9753 ;
  assign n9767 = ~n2409 & n9753 ;
  assign n9768 = ~n2408 & n9767 ;
  assign n9769 = ~n9766 & ~n9768 ;
  assign n9770 = ~\ctl_rf_c1_rf_chllp_reg[21]/NET0131  & ~n9753 ;
  assign n9771 = ~n2366 & n9753 ;
  assign n9772 = ~n2365 & n9771 ;
  assign n9773 = ~n9770 & ~n9772 ;
  assign n9774 = ~\ctl_rf_c1_rf_chllp_reg[22]/NET0131  & ~n9753 ;
  assign n9775 = ~n2500 & n9753 ;
  assign n9776 = ~n2499 & n9775 ;
  assign n9777 = ~n9774 & ~n9776 ;
  assign n9778 = ~\ctl_rf_c1_rf_chllp_reg[23]/NET0131  & ~n9753 ;
  assign n9779 = ~n2529 & n9753 ;
  assign n9780 = ~n2528 & n9779 ;
  assign n9781 = ~n9778 & ~n9780 ;
  assign n9782 = \ctl_rf_be_d1_reg[3]/P0001  & n9725 ;
  assign n9783 = n8578 & n9782 ;
  assign n9784 = ~\ctl_rf_c1_rf_chllp_reg[25]/NET0131  & ~n9783 ;
  assign n9785 = \hwdata[25]_pad  & ~n2242 ;
  assign n9786 = \hwdata[1]_pad  & n2242 ;
  assign n9787 = ~n9785 & ~n9786 ;
  assign n9788 = ~n2240 & ~n9787 ;
  assign n9789 = \hwdata[9]_pad  & n2240 ;
  assign n9790 = n9783 & ~n9789 ;
  assign n9791 = ~n9788 & n9790 ;
  assign n9792 = ~n9784 & ~n9791 ;
  assign n9793 = ~\ctl_rf_c1_rf_chllp_reg[26]/NET0131  & ~n9783 ;
  assign n9794 = \hwdata[26]_pad  & ~n2242 ;
  assign n9795 = \hwdata[2]_pad  & n2242 ;
  assign n9796 = ~n9794 & ~n9795 ;
  assign n9797 = ~n2240 & ~n9796 ;
  assign n9798 = \hwdata[10]_pad  & n2240 ;
  assign n9799 = n9783 & ~n9798 ;
  assign n9800 = ~n9797 & n9799 ;
  assign n9801 = ~n9793 & ~n9800 ;
  assign n9802 = ~\ctl_rf_c1_rf_chllp_reg[27]/NET0131  & ~n9783 ;
  assign n9803 = \hwdata[27]_pad  & ~n2242 ;
  assign n9804 = \hwdata[3]_pad  & n2242 ;
  assign n9805 = ~n9803 & ~n9804 ;
  assign n9806 = ~n2240 & ~n9805 ;
  assign n9807 = \hwdata[11]_pad  & n2240 ;
  assign n9808 = n9783 & ~n9807 ;
  assign n9809 = ~n9806 & n9808 ;
  assign n9810 = ~n9802 & ~n9809 ;
  assign n9811 = ~\ctl_rf_c1_rf_chllp_reg[28]/NET0131  & ~n9783 ;
  assign n9812 = \hwdata[28]_pad  & ~n2242 ;
  assign n9813 = \hwdata[4]_pad  & n2242 ;
  assign n9814 = ~n9812 & ~n9813 ;
  assign n9815 = ~n2240 & ~n9814 ;
  assign n9816 = \hwdata[12]_pad  & n2240 ;
  assign n9817 = n9783 & ~n9816 ;
  assign n9818 = ~n9815 & n9817 ;
  assign n9819 = ~n9811 & ~n9818 ;
  assign n9820 = \ctl_rf_be_d1_reg[0]/P0001  & n9725 ;
  assign n9821 = n8578 & n9820 ;
  assign n9822 = ~\ctl_rf_c1_rf_chllp_reg[4]/NET0131  & ~n9821 ;
  assign n9823 = ~n8714 & n9821 ;
  assign n9824 = ~n8713 & n9823 ;
  assign n9825 = ~n9822 & ~n9824 ;
  assign n9826 = ~\ctl_rf_c1_rf_chllp_reg[5]/NET0131  & ~n9821 ;
  assign n9827 = ~n8587 & n9821 ;
  assign n9828 = ~n8586 & n9827 ;
  assign n9829 = ~n9826 & ~n9828 ;
  assign n9830 = ~\ctl_rf_c1_rf_chllp_reg[6]/NET0131  & ~n9821 ;
  assign n9831 = ~n8596 & n9821 ;
  assign n9832 = ~n8595 & n9831 ;
  assign n9833 = ~n9830 & ~n9832 ;
  assign n9834 = ~\ctl_rf_c1_rf_chllp_reg[7]/NET0131  & ~n9821 ;
  assign n9835 = ~n2247 & n9821 ;
  assign n9836 = ~n2246 & n9835 ;
  assign n9837 = ~n9834 & ~n9836 ;
  assign n9838 = ~\ctl_rf_c1_rf_chllp_reg[8]/NET0131  & ~n9727 ;
  assign n9839 = ~n8781 & n9727 ;
  assign n9840 = ~n8780 & n9839 ;
  assign n9841 = ~n9838 & ~n9840 ;
  assign n9842 = ~\ctl_rf_c1_rf_chllp_reg[9]/NET0131  & ~n9727 ;
  assign n9843 = ~n8808 & n9727 ;
  assign n9844 = ~n8807 & n9843 ;
  assign n9845 = ~n9842 & ~n9844 ;
  assign n9846 = n8609 & n9726 ;
  assign n9847 = ~\ctl_rf_c3_rf_chllp_reg[10]/NET0131  & ~n9846 ;
  assign n9848 = ~n8759 & n9846 ;
  assign n9849 = ~n8758 & n9848 ;
  assign n9850 = ~n9847 & ~n9849 ;
  assign n9851 = ~\ctl_rf_c3_rf_chllp_reg[11]/NET0131  & ~n9846 ;
  assign n9852 = ~n8791 & n9846 ;
  assign n9853 = ~n8790 & n9852 ;
  assign n9854 = ~n9851 & ~n9853 ;
  assign n9855 = ~\ctl_rf_c3_rf_chllp_reg[12]/NET0131  & ~n9846 ;
  assign n9856 = ~n8768 & n9846 ;
  assign n9857 = ~n8767 & n9856 ;
  assign n9858 = ~n9855 & ~n9857 ;
  assign n9859 = ~\ctl_rf_c3_rf_chllp_reg[14]/NET0131  & ~n9846 ;
  assign n9860 = ~n9027 & n9846 ;
  assign n9861 = ~n9026 & n9860 ;
  assign n9862 = ~n9859 & ~n9861 ;
  assign n9863 = ~\ctl_rf_c3_rf_chllp_reg[13]/NET0131  & ~n9846 ;
  assign n9864 = ~n9018 & n9846 ;
  assign n9865 = ~n9017 & n9864 ;
  assign n9866 = ~n9863 & ~n9865 ;
  assign n9867 = ~\ctl_rf_c3_rf_chllp_reg[15]/NET0131  & ~n9846 ;
  assign n9868 = ~n3763 & n9846 ;
  assign n9869 = ~n3762 & n9868 ;
  assign n9870 = ~n9867 & ~n9869 ;
  assign n9871 = n8609 & n9752 ;
  assign n9872 = ~\ctl_rf_c3_rf_chllp_reg[16]/NET0131  & ~n9871 ;
  assign n9873 = ~n2680 & n9871 ;
  assign n9874 = ~n2679 & n9873 ;
  assign n9875 = ~n9872 & ~n9874 ;
  assign n9876 = ~\ctl_rf_c3_rf_chllp_reg[17]/NET0131  & ~n9871 ;
  assign n9877 = ~n2260 & n9871 ;
  assign n9878 = ~n2259 & n9877 ;
  assign n9879 = ~n9876 & ~n9878 ;
  assign n9880 = ~\ctl_rf_c3_rf_chllp_reg[18]/NET0131  & ~n9871 ;
  assign n9881 = ~n2400 & n9871 ;
  assign n9882 = ~n2399 & n9881 ;
  assign n9883 = ~n9880 & ~n9882 ;
  assign n9884 = ~\ctl_rf_c3_rf_chllp_reg[19]/NET0131  & ~n9871 ;
  assign n9885 = ~n2409 & n9871 ;
  assign n9886 = ~n2408 & n9885 ;
  assign n9887 = ~n9884 & ~n9886 ;
  assign n9888 = ~\ctl_rf_c3_rf_chllp_reg[22]/NET0131  & ~n9871 ;
  assign n9889 = ~n2500 & n9871 ;
  assign n9890 = ~n2499 & n9889 ;
  assign n9891 = ~n9888 & ~n9890 ;
  assign n9892 = ~\ctl_rf_c3_rf_chllp_reg[23]/NET0131  & ~n9871 ;
  assign n9893 = ~n2529 & n9871 ;
  assign n9894 = ~n2528 & n9893 ;
  assign n9895 = ~n9892 & ~n9894 ;
  assign n9896 = n8609 & n9782 ;
  assign n9897 = ~\ctl_rf_c3_rf_chllp_reg[25]/NET0131  & ~n9896 ;
  assign n9898 = ~n9789 & n9896 ;
  assign n9899 = ~n9788 & n9898 ;
  assign n9900 = ~n9897 & ~n9899 ;
  assign n9901 = ~\ctl_rf_c3_rf_chllp_reg[26]/NET0131  & ~n9896 ;
  assign n9902 = ~n9798 & n9896 ;
  assign n9903 = ~n9797 & n9902 ;
  assign n9904 = ~n9901 & ~n9903 ;
  assign n9905 = ~\ctl_rf_c3_rf_chllp_reg[27]/NET0131  & ~n9896 ;
  assign n9906 = ~n9807 & n9896 ;
  assign n9907 = ~n9806 & n9906 ;
  assign n9908 = ~n9905 & ~n9907 ;
  assign n9909 = ~\ctl_rf_c3_rf_chllp_reg[28]/NET0131  & ~n9896 ;
  assign n9910 = ~n9816 & n9896 ;
  assign n9911 = ~n9815 & n9910 ;
  assign n9912 = ~n9909 & ~n9911 ;
  assign n9913 = n8609 & n9820 ;
  assign n9914 = ~\ctl_rf_c3_rf_chllp_reg[4]/NET0131  & ~n9913 ;
  assign n9915 = ~n8714 & n9913 ;
  assign n9916 = ~n8713 & n9915 ;
  assign n9917 = ~n9914 & ~n9916 ;
  assign n9918 = ~\ctl_rf_c3_rf_chllp_reg[5]/NET0131  & ~n9913 ;
  assign n9919 = ~n8587 & n9913 ;
  assign n9920 = ~n8586 & n9919 ;
  assign n9921 = ~n9918 & ~n9920 ;
  assign n9922 = ~\ctl_rf_c3_rf_chllp_reg[6]/NET0131  & ~n9913 ;
  assign n9923 = ~n8596 & n9913 ;
  assign n9924 = ~n8595 & n9923 ;
  assign n9925 = ~n9922 & ~n9924 ;
  assign n9926 = ~\ctl_rf_c3_rf_chllp_reg[7]/NET0131  & ~n9913 ;
  assign n9927 = ~n2247 & n9913 ;
  assign n9928 = ~n2246 & n9927 ;
  assign n9929 = ~n9926 & ~n9928 ;
  assign n9930 = ~\ctl_rf_c3_rf_chllp_reg[8]/NET0131  & ~n9846 ;
  assign n9931 = ~n8781 & n9846 ;
  assign n9932 = ~n8780 & n9931 ;
  assign n9933 = ~n9930 & ~n9932 ;
  assign n9934 = ~\ctl_rf_c3_rf_chllp_reg[9]/NET0131  & ~n9846 ;
  assign n9935 = ~n8808 & n9846 ;
  assign n9936 = ~n8807 & n9935 ;
  assign n9937 = ~n9934 & ~n9936 ;
  assign n9938 = ~\ahb_slv_slv_ad_d1o_reg[2]/NET0131  & \ahb_slv_slv_ad_d1o_reg[8]/NET0131  ;
  assign n9939 = n2275 & n9938 ;
  assign n9940 = \ctl_rf_be_d1_reg[1]/P0001  & n9939 ;
  assign n9941 = n8629 & n9940 ;
  assign n9942 = ~\ctl_rf_c4_rf_chllp_reg[10]/NET0131  & ~n9941 ;
  assign n9943 = ~n8759 & n9941 ;
  assign n9944 = ~n8758 & n9943 ;
  assign n9945 = ~n9942 & ~n9944 ;
  assign n9946 = ~\ctl_rf_c4_rf_chllp_reg[11]/NET0131  & ~n9941 ;
  assign n9947 = ~n8791 & n9941 ;
  assign n9948 = ~n8790 & n9947 ;
  assign n9949 = ~n9946 & ~n9948 ;
  assign n9950 = ~\ctl_rf_c4_rf_chllp_reg[12]/NET0131  & ~n9941 ;
  assign n9951 = ~n8768 & n9941 ;
  assign n9952 = ~n8767 & n9951 ;
  assign n9953 = ~n9950 & ~n9952 ;
  assign n9954 = ~\ctl_rf_c4_rf_chllp_reg[13]/NET0131  & ~n9941 ;
  assign n9955 = ~n9018 & n9941 ;
  assign n9956 = ~n9017 & n9955 ;
  assign n9957 = ~n9954 & ~n9956 ;
  assign n9958 = ~\ctl_rf_c4_rf_chllp_reg[14]/NET0131  & ~n9941 ;
  assign n9959 = ~n9027 & n9941 ;
  assign n9960 = ~n9026 & n9959 ;
  assign n9961 = ~n9958 & ~n9960 ;
  assign n9962 = ~\ctl_rf_c4_rf_chllp_reg[15]/NET0131  & ~n9941 ;
  assign n9963 = ~n3763 & n9941 ;
  assign n9964 = ~n3762 & n9963 ;
  assign n9965 = ~n9962 & ~n9964 ;
  assign n9966 = \ctl_rf_be_d1_reg[2]/P0001  & n9939 ;
  assign n9967 = n8629 & n9966 ;
  assign n9968 = ~\ctl_rf_c4_rf_chllp_reg[16]/NET0131  & ~n9967 ;
  assign n9969 = ~n2680 & n9967 ;
  assign n9970 = ~n2679 & n9969 ;
  assign n9971 = ~n9968 & ~n9970 ;
  assign n9972 = ~\ctl_rf_c4_rf_chllp_reg[17]/NET0131  & ~n9967 ;
  assign n9973 = ~n2260 & n9967 ;
  assign n9974 = ~n2259 & n9973 ;
  assign n9975 = ~n9972 & ~n9974 ;
  assign n9976 = ~\ctl_rf_c4_rf_chllp_reg[18]/NET0131  & ~n9967 ;
  assign n9977 = ~n2400 & n9967 ;
  assign n9978 = ~n2399 & n9977 ;
  assign n9979 = ~n9976 & ~n9978 ;
  assign n9980 = ~\ctl_rf_c4_rf_chllp_reg[19]/NET0131  & ~n9967 ;
  assign n9981 = ~n2409 & n9967 ;
  assign n9982 = ~n2408 & n9981 ;
  assign n9983 = ~n9980 & ~n9982 ;
  assign n9984 = ~\ctl_rf_c4_rf_chllp_reg[21]/NET0131  & ~n9967 ;
  assign n9985 = ~n2366 & n9967 ;
  assign n9986 = ~n2365 & n9985 ;
  assign n9987 = ~n9984 & ~n9986 ;
  assign n9988 = ~\ctl_rf_c4_rf_chllp_reg[22]/NET0131  & ~n9967 ;
  assign n9989 = ~n2500 & n9967 ;
  assign n9990 = ~n2499 & n9989 ;
  assign n9991 = ~n9988 & ~n9990 ;
  assign n9992 = ~\ctl_rf_c4_rf_chllp_reg[23]/NET0131  & ~n9967 ;
  assign n9993 = ~n2529 & n9967 ;
  assign n9994 = ~n2528 & n9993 ;
  assign n9995 = ~n9992 & ~n9994 ;
  assign n9996 = \ctl_rf_be_d1_reg[3]/P0001  & n9939 ;
  assign n9997 = n8629 & n9996 ;
  assign n9998 = ~\ctl_rf_c4_rf_chllp_reg[25]/NET0131  & ~n9997 ;
  assign n9999 = ~n9789 & n9997 ;
  assign n10000 = ~n9788 & n9999 ;
  assign n10001 = ~n9998 & ~n10000 ;
  assign n10002 = ~\ctl_rf_c4_rf_chllp_reg[26]/NET0131  & ~n9997 ;
  assign n10003 = ~n9798 & n9997 ;
  assign n10004 = ~n9797 & n10003 ;
  assign n10005 = ~n10002 & ~n10004 ;
  assign n10006 = ~\ctl_rf_c4_rf_chllp_reg[27]/NET0131  & ~n9997 ;
  assign n10007 = ~n9807 & n9997 ;
  assign n10008 = ~n9806 & n10007 ;
  assign n10009 = ~n10006 & ~n10008 ;
  assign n10010 = ~\ctl_rf_c4_rf_chllp_reg[28]/NET0131  & ~n9997 ;
  assign n10011 = ~n9816 & n9997 ;
  assign n10012 = ~n9815 & n10011 ;
  assign n10013 = ~n10010 & ~n10012 ;
  assign n10014 = \ctl_rf_be_d1_reg[0]/P0001  & n9939 ;
  assign n10015 = n8629 & n10014 ;
  assign n10016 = ~\ctl_rf_c4_rf_chllp_reg[4]/NET0131  & ~n10015 ;
  assign n10017 = ~n8714 & n10015 ;
  assign n10018 = ~n8713 & n10017 ;
  assign n10019 = ~n10016 & ~n10018 ;
  assign n10020 = ~\ctl_rf_c4_rf_chllp_reg[5]/NET0131  & ~n10015 ;
  assign n10021 = ~n8587 & n10015 ;
  assign n10022 = ~n8586 & n10021 ;
  assign n10023 = ~n10020 & ~n10022 ;
  assign n10024 = ~\ctl_rf_c4_rf_chllp_reg[6]/NET0131  & ~n10015 ;
  assign n10025 = ~n8596 & n10015 ;
  assign n10026 = ~n8595 & n10025 ;
  assign n10027 = ~n10024 & ~n10026 ;
  assign n10028 = ~\ctl_rf_c4_rf_chllp_reg[7]/NET0131  & ~n10015 ;
  assign n10029 = ~n2247 & n10015 ;
  assign n10030 = ~n2246 & n10029 ;
  assign n10031 = ~n10028 & ~n10030 ;
  assign n10032 = ~\ctl_rf_c4_rf_chllp_reg[8]/NET0131  & ~n9941 ;
  assign n10033 = ~n8781 & n9941 ;
  assign n10034 = ~n8780 & n10033 ;
  assign n10035 = ~n10032 & ~n10034 ;
  assign n10036 = ~\ctl_rf_c4_rf_chllp_reg[9]/NET0131  & ~n9941 ;
  assign n10037 = ~n8808 & n9941 ;
  assign n10038 = ~n8807 & n10037 ;
  assign n10039 = ~n10036 & ~n10038 ;
  assign n10040 = n8629 & n9726 ;
  assign n10041 = ~\ctl_rf_c5_rf_chllp_reg[10]/NET0131  & ~n10040 ;
  assign n10042 = ~n8759 & n10040 ;
  assign n10043 = ~n8758 & n10042 ;
  assign n10044 = ~n10041 & ~n10043 ;
  assign n10045 = ~\ctl_rf_c5_rf_chllp_reg[11]/NET0131  & ~n10040 ;
  assign n10046 = ~n8791 & n10040 ;
  assign n10047 = ~n8790 & n10046 ;
  assign n10048 = ~n10045 & ~n10047 ;
  assign n10049 = ~\ctl_rf_c5_rf_chllp_reg[12]/NET0131  & ~n10040 ;
  assign n10050 = ~n8768 & n10040 ;
  assign n10051 = ~n8767 & n10050 ;
  assign n10052 = ~n10049 & ~n10051 ;
  assign n10053 = ~\ctl_rf_c5_rf_chllp_reg[13]/NET0131  & ~n10040 ;
  assign n10054 = ~n9018 & n10040 ;
  assign n10055 = ~n9017 & n10054 ;
  assign n10056 = ~n10053 & ~n10055 ;
  assign n10057 = ~\ctl_rf_c5_rf_chllp_reg[14]/NET0131  & ~n10040 ;
  assign n10058 = ~n9027 & n10040 ;
  assign n10059 = ~n9026 & n10058 ;
  assign n10060 = ~n10057 & ~n10059 ;
  assign n10061 = ~\ctl_rf_c5_rf_chllp_reg[15]/NET0131  & ~n10040 ;
  assign n10062 = ~n3763 & n10040 ;
  assign n10063 = ~n3762 & n10062 ;
  assign n10064 = ~n10061 & ~n10063 ;
  assign n10065 = n8629 & n9752 ;
  assign n10066 = ~\ctl_rf_c5_rf_chllp_reg[16]/NET0131  & ~n10065 ;
  assign n10067 = ~n2680 & n10065 ;
  assign n10068 = ~n2679 & n10067 ;
  assign n10069 = ~n10066 & ~n10068 ;
  assign n10070 = ~\ctl_rf_c5_rf_chllp_reg[17]/NET0131  & ~n10065 ;
  assign n10071 = ~n2260 & n10065 ;
  assign n10072 = ~n2259 & n10071 ;
  assign n10073 = ~n10070 & ~n10072 ;
  assign n10074 = ~\ctl_rf_c5_rf_chllp_reg[18]/NET0131  & ~n10065 ;
  assign n10075 = ~n2400 & n10065 ;
  assign n10076 = ~n2399 & n10075 ;
  assign n10077 = ~n10074 & ~n10076 ;
  assign n10078 = ~\ctl_rf_c5_rf_chllp_reg[19]/NET0131  & ~n10065 ;
  assign n10079 = ~n2409 & n10065 ;
  assign n10080 = ~n2408 & n10079 ;
  assign n10081 = ~n10078 & ~n10080 ;
  assign n10082 = ~\ctl_rf_c5_rf_chllp_reg[21]/NET0131  & ~n10065 ;
  assign n10083 = ~n2366 & n10065 ;
  assign n10084 = ~n2365 & n10083 ;
  assign n10085 = ~n10082 & ~n10084 ;
  assign n10086 = ~\ctl_rf_c5_rf_chllp_reg[22]/NET0131  & ~n10065 ;
  assign n10087 = ~n2500 & n10065 ;
  assign n10088 = ~n2499 & n10087 ;
  assign n10089 = ~n10086 & ~n10088 ;
  assign n10090 = ~\ctl_rf_c5_rf_chllp_reg[23]/NET0131  & ~n10065 ;
  assign n10091 = ~n2529 & n10065 ;
  assign n10092 = ~n2528 & n10091 ;
  assign n10093 = ~n10090 & ~n10092 ;
  assign n10094 = n8629 & n9782 ;
  assign n10095 = ~\ctl_rf_c5_rf_chllp_reg[25]/NET0131  & ~n10094 ;
  assign n10096 = ~n9789 & n10094 ;
  assign n10097 = ~n9788 & n10096 ;
  assign n10098 = ~n10095 & ~n10097 ;
  assign n10099 = ~\ctl_rf_c5_rf_chllp_reg[26]/NET0131  & ~n10094 ;
  assign n10100 = ~n9798 & n10094 ;
  assign n10101 = ~n9797 & n10100 ;
  assign n10102 = ~n10099 & ~n10101 ;
  assign n10103 = ~\ctl_rf_c5_rf_chllp_reg[27]/NET0131  & ~n10094 ;
  assign n10104 = ~n9807 & n10094 ;
  assign n10105 = ~n9806 & n10104 ;
  assign n10106 = ~n10103 & ~n10105 ;
  assign n10107 = ~\ctl_rf_c5_rf_chllp_reg[28]/NET0131  & ~n10094 ;
  assign n10108 = ~n9816 & n10094 ;
  assign n10109 = ~n9815 & n10108 ;
  assign n10110 = ~n10107 & ~n10109 ;
  assign n10111 = n8629 & n9820 ;
  assign n10112 = ~\ctl_rf_c5_rf_chllp_reg[4]/NET0131  & ~n10111 ;
  assign n10113 = ~n8714 & n10111 ;
  assign n10114 = ~n8713 & n10113 ;
  assign n10115 = ~n10112 & ~n10114 ;
  assign n10116 = ~\ctl_rf_c5_rf_chllp_reg[5]/NET0131  & ~n10111 ;
  assign n10117 = ~n8587 & n10111 ;
  assign n10118 = ~n8586 & n10117 ;
  assign n10119 = ~n10116 & ~n10118 ;
  assign n10120 = ~\ctl_rf_c5_rf_chllp_reg[6]/NET0131  & ~n10111 ;
  assign n10121 = ~n8596 & n10111 ;
  assign n10122 = ~n8595 & n10121 ;
  assign n10123 = ~n10120 & ~n10122 ;
  assign n10124 = \hrdata_reg[17]_pad  & ~n4569 ;
  assign n10125 = n4745 & n5771 ;
  assign n10126 = n5744 & n10125 ;
  assign n10127 = ~n4746 & ~n10126 ;
  assign n10128 = ~n4573 & ~n10127 ;
  assign n10129 = ~n5370 & ~n5425 ;
  assign n10130 = ~n4573 & ~n4745 ;
  assign n10131 = ~n10129 & n10130 ;
  assign n10132 = ~n10128 & ~n10131 ;
  assign n10133 = n4573 & ~n5670 ;
  assign n10134 = ~n5651 & n10133 ;
  assign n10135 = n4569 & ~n10134 ;
  assign n10136 = n10132 & n10135 ;
  assign n10137 = ~n10124 & ~n10136 ;
  assign n10138 = ~\ctl_rf_c5_rf_chllp_reg[7]/NET0131  & ~n10111 ;
  assign n10139 = ~n2247 & n10111 ;
  assign n10140 = ~n2246 & n10139 ;
  assign n10141 = ~n10138 & ~n10140 ;
  assign n10142 = ~\ctl_rf_c5_rf_chllp_reg[8]/NET0131  & ~n10040 ;
  assign n10143 = ~n8781 & n10040 ;
  assign n10144 = ~n8780 & n10143 ;
  assign n10145 = ~n10142 & ~n10144 ;
  assign n10146 = ~\ctl_rf_c5_rf_chllp_reg[9]/NET0131  & ~n10040 ;
  assign n10147 = ~n8808 & n10040 ;
  assign n10148 = ~n8807 & n10147 ;
  assign n10149 = ~n10146 & ~n10148 ;
  assign n10150 = \hrdata_reg[18]_pad  & ~n4569 ;
  assign n10151 = n4745 & n5881 ;
  assign n10152 = n5854 & n10151 ;
  assign n10153 = ~n4746 & ~n10152 ;
  assign n10154 = ~n4573 & ~n10153 ;
  assign n10155 = ~n7154 & ~n7209 ;
  assign n10156 = n10130 & ~n10155 ;
  assign n10157 = ~n10154 & ~n10156 ;
  assign n10158 = n4573 & ~n6125 ;
  assign n10159 = ~n6108 & n10158 ;
  assign n10160 = n4569 & ~n10159 ;
  assign n10161 = n10157 & n10160 ;
  assign n10162 = ~n10150 & ~n10161 ;
  assign n10163 = n2230 & n8577 ;
  assign n10164 = \ctl_rf_be_d1_reg[1]/P0001  & n10163 ;
  assign n10165 = n8656 & n10164 ;
  assign n10166 = ~\ctl_rf_c6_rf_chllp_reg[10]/NET0131  & ~n10165 ;
  assign n10167 = ~n8759 & n10165 ;
  assign n10168 = ~n8758 & n10167 ;
  assign n10169 = ~n10166 & ~n10168 ;
  assign n10170 = ~\ctl_rf_c6_rf_chllp_reg[11]/NET0131  & ~n10165 ;
  assign n10171 = ~n8791 & n10165 ;
  assign n10172 = ~n8790 & n10171 ;
  assign n10173 = ~n10170 & ~n10172 ;
  assign n10174 = ~\ctl_rf_c6_rf_chllp_reg[12]/NET0131  & ~n10165 ;
  assign n10175 = ~n8768 & n10165 ;
  assign n10176 = ~n8767 & n10175 ;
  assign n10177 = ~n10174 & ~n10176 ;
  assign n10178 = ~\ctl_rf_c6_rf_chllp_reg[13]/NET0131  & ~n10165 ;
  assign n10179 = ~n9018 & n10165 ;
  assign n10180 = ~n9017 & n10179 ;
  assign n10181 = ~n10178 & ~n10180 ;
  assign n10182 = ~\ctl_rf_c6_rf_chllp_reg[14]/NET0131  & ~n10165 ;
  assign n10183 = ~n9027 & n10165 ;
  assign n10184 = ~n9026 & n10183 ;
  assign n10185 = ~n10182 & ~n10184 ;
  assign n10186 = ~\ctl_rf_c6_rf_chllp_reg[15]/NET0131  & ~n10165 ;
  assign n10187 = ~n3763 & n10165 ;
  assign n10188 = ~n3762 & n10187 ;
  assign n10189 = ~n10186 & ~n10188 ;
  assign n10190 = \ctl_rf_be_d1_reg[2]/P0001  & n10163 ;
  assign n10191 = n8656 & n10190 ;
  assign n10192 = ~\ctl_rf_c6_rf_chllp_reg[16]/NET0131  & ~n10191 ;
  assign n10193 = ~n2680 & n10191 ;
  assign n10194 = ~n2679 & n10193 ;
  assign n10195 = ~n10192 & ~n10194 ;
  assign n10196 = ~\ctl_rf_c6_rf_chllp_reg[17]/NET0131  & ~n10191 ;
  assign n10197 = ~n2260 & n10191 ;
  assign n10198 = ~n2259 & n10197 ;
  assign n10199 = ~n10196 & ~n10198 ;
  assign n10200 = ~\ctl_rf_c6_rf_chllp_reg[19]/NET0131  & ~n10191 ;
  assign n10201 = ~n2409 & n10191 ;
  assign n10202 = ~n2408 & n10201 ;
  assign n10203 = ~n10200 & ~n10202 ;
  assign n10204 = ~\ctl_rf_c6_rf_chllp_reg[21]/NET0131  & ~n10191 ;
  assign n10205 = ~n2366 & n10191 ;
  assign n10206 = ~n2365 & n10205 ;
  assign n10207 = ~n10204 & ~n10206 ;
  assign n10208 = ~\ctl_rf_c6_rf_chllp_reg[23]/NET0131  & ~n10191 ;
  assign n10209 = ~n2529 & n10191 ;
  assign n10210 = ~n2528 & n10209 ;
  assign n10211 = ~n10208 & ~n10210 ;
  assign n10212 = \ctl_rf_be_d1_reg[3]/P0001  & n10163 ;
  assign n10213 = n8656 & n10212 ;
  assign n10214 = ~\ctl_rf_c6_rf_chllp_reg[25]/NET0131  & ~n10213 ;
  assign n10215 = ~n9789 & n10213 ;
  assign n10216 = ~n9788 & n10215 ;
  assign n10217 = ~n10214 & ~n10216 ;
  assign n10218 = ~\ctl_rf_c6_rf_chllp_reg[26]/NET0131  & ~n10213 ;
  assign n10219 = ~n9798 & n10213 ;
  assign n10220 = ~n9797 & n10219 ;
  assign n10221 = ~n10218 & ~n10220 ;
  assign n10222 = ~\ctl_rf_c6_rf_chllp_reg[27]/NET0131  & ~n10213 ;
  assign n10223 = ~n9807 & n10213 ;
  assign n10224 = ~n9806 & n10223 ;
  assign n10225 = ~n10222 & ~n10224 ;
  assign n10226 = ~\ctl_rf_c6_rf_chllp_reg[28]/NET0131  & ~n10213 ;
  assign n10227 = ~n9816 & n10213 ;
  assign n10228 = ~n9815 & n10227 ;
  assign n10229 = ~n10226 & ~n10228 ;
  assign n10230 = \ctl_rf_be_d1_reg[0]/P0001  & n10163 ;
  assign n10231 = n8656 & n10230 ;
  assign n10232 = ~\ctl_rf_c6_rf_chllp_reg[4]/NET0131  & ~n10231 ;
  assign n10233 = ~n8714 & n10231 ;
  assign n10234 = ~n8713 & n10233 ;
  assign n10235 = ~n10232 & ~n10234 ;
  assign n10236 = ~\ctl_rf_c6_rf_chllp_reg[5]/NET0131  & ~n10231 ;
  assign n10237 = ~n8587 & n10231 ;
  assign n10238 = ~n8586 & n10237 ;
  assign n10239 = ~n10236 & ~n10238 ;
  assign n10240 = ~\ctl_rf_c6_rf_chllp_reg[6]/NET0131  & ~n10231 ;
  assign n10241 = ~n8596 & n10231 ;
  assign n10242 = ~n8595 & n10241 ;
  assign n10243 = ~n10240 & ~n10242 ;
  assign n10244 = ~\ctl_rf_c6_rf_chllp_reg[7]/NET0131  & ~n10231 ;
  assign n10245 = ~n2247 & n10231 ;
  assign n10246 = ~n2246 & n10245 ;
  assign n10247 = ~n10244 & ~n10246 ;
  assign n10248 = ~\ctl_rf_c6_rf_chllp_reg[8]/NET0131  & ~n10165 ;
  assign n10249 = ~n8781 & n10165 ;
  assign n10250 = ~n8780 & n10249 ;
  assign n10251 = ~n10248 & ~n10250 ;
  assign n10252 = ~\ctl_rf_c6_rf_chllp_reg[9]/NET0131  & ~n10165 ;
  assign n10253 = ~n8808 & n10165 ;
  assign n10254 = ~n8807 & n10253 ;
  assign n10255 = ~n10252 & ~n10254 ;
  assign n10256 = \hrdata_reg[19]_pad  & ~n4569 ;
  assign n10257 = n4745 & n6226 ;
  assign n10258 = n6199 & n10257 ;
  assign n10259 = ~n4746 & ~n10258 ;
  assign n10260 = ~n4573 & ~n10259 ;
  assign n10261 = ~n7935 & ~n7990 ;
  assign n10262 = n10130 & ~n10261 ;
  assign n10263 = ~n10260 & ~n10262 ;
  assign n10264 = n4573 & ~n6451 ;
  assign n10265 = ~n6437 & n10264 ;
  assign n10266 = n4569 & ~n10265 ;
  assign n10267 = n10263 & n10266 ;
  assign n10268 = ~n10256 & ~n10267 ;
  assign n10269 = \hrdata_reg[20]_pad  & ~n4569 ;
  assign n10270 = ~n4745 & ~n8134 ;
  assign n10271 = ~n8079 & n10270 ;
  assign n10272 = n6513 & ~n6529 ;
  assign n10273 = \haddr[8]_pad  & n4745 ;
  assign n10274 = ~n10272 & n10273 ;
  assign n10275 = ~n4573 & ~n10274 ;
  assign n10276 = ~n10271 & n10275 ;
  assign n10277 = n4573 & ~n6754 ;
  assign n10278 = ~n6740 & n10277 ;
  assign n10279 = n4569 & ~n10278 ;
  assign n10280 = ~n10276 & n10279 ;
  assign n10281 = ~n10269 & ~n10280 ;
  assign n10282 = \hrdata_reg[21]_pad  & ~n4569 ;
  assign n10283 = ~n4745 & ~n8278 ;
  assign n10284 = ~n8223 & n10283 ;
  assign n10285 = n6816 & ~n6832 ;
  assign n10286 = n10273 & ~n10285 ;
  assign n10287 = ~n4573 & ~n10286 ;
  assign n10288 = ~n10284 & n10287 ;
  assign n10289 = n4573 & ~n7057 ;
  assign n10290 = ~n7043 & n10289 ;
  assign n10291 = n4569 & ~n10290 ;
  assign n10292 = ~n10288 & n10291 ;
  assign n10293 = ~n10282 & ~n10292 ;
  assign n10294 = n8677 & n10164 ;
  assign n10295 = ~\ctl_rf_c7_rf_chllp_reg[10]/NET0131  & ~n10294 ;
  assign n10296 = ~n8759 & n10294 ;
  assign n10297 = ~n8758 & n10296 ;
  assign n10298 = ~n10295 & ~n10297 ;
  assign n10299 = ~\ctl_rf_c7_rf_chllp_reg[11]/NET0131  & ~n10294 ;
  assign n10300 = ~n8791 & n10294 ;
  assign n10301 = ~n8790 & n10300 ;
  assign n10302 = ~n10299 & ~n10301 ;
  assign n10303 = ~\ctl_rf_c7_rf_chllp_reg[12]/NET0131  & ~n10294 ;
  assign n10304 = ~n8768 & n10294 ;
  assign n10305 = ~n8767 & n10304 ;
  assign n10306 = ~n10303 & ~n10305 ;
  assign n10307 = ~\ctl_rf_c7_rf_chllp_reg[13]/NET0131  & ~n10294 ;
  assign n10308 = ~n9018 & n10294 ;
  assign n10309 = ~n9017 & n10308 ;
  assign n10310 = ~n10307 & ~n10309 ;
  assign n10311 = ~\ctl_rf_c7_rf_chllp_reg[14]/NET0131  & ~n10294 ;
  assign n10312 = ~n9027 & n10294 ;
  assign n10313 = ~n9026 & n10312 ;
  assign n10314 = ~n10311 & ~n10313 ;
  assign n10315 = ~\ctl_rf_c7_rf_chllp_reg[15]/NET0131  & ~n10294 ;
  assign n10316 = ~n3763 & n10294 ;
  assign n10317 = ~n3762 & n10316 ;
  assign n10318 = ~n10315 & ~n10317 ;
  assign n10319 = n8677 & n10190 ;
  assign n10320 = ~\ctl_rf_c7_rf_chllp_reg[16]/NET0131  & ~n10319 ;
  assign n10321 = ~n2680 & n10319 ;
  assign n10322 = ~n2679 & n10321 ;
  assign n10323 = ~n10320 & ~n10322 ;
  assign n10324 = ~\ctl_rf_c7_rf_chllp_reg[17]/NET0131  & ~n10319 ;
  assign n10325 = ~n2260 & n10319 ;
  assign n10326 = ~n2259 & n10325 ;
  assign n10327 = ~n10324 & ~n10326 ;
  assign n10328 = ~\ctl_rf_c7_rf_chllp_reg[18]/NET0131  & ~n10319 ;
  assign n10329 = ~n2400 & n10319 ;
  assign n10330 = ~n2399 & n10329 ;
  assign n10331 = ~n10328 & ~n10330 ;
  assign n10332 = ~\ctl_rf_c7_rf_chllp_reg[19]/NET0131  & ~n10319 ;
  assign n10333 = ~n2409 & n10319 ;
  assign n10334 = ~n2408 & n10333 ;
  assign n10335 = ~n10332 & ~n10334 ;
  assign n10336 = ~\ctl_rf_c7_rf_chllp_reg[21]/NET0131  & ~n10319 ;
  assign n10337 = ~n2366 & n10319 ;
  assign n10338 = ~n2365 & n10337 ;
  assign n10339 = ~n10336 & ~n10338 ;
  assign n10340 = ~\ctl_rf_c7_rf_chllp_reg[22]/NET0131  & ~n10319 ;
  assign n10341 = ~n2500 & n10319 ;
  assign n10342 = ~n2499 & n10341 ;
  assign n10343 = ~n10340 & ~n10342 ;
  assign n10344 = ~\ctl_rf_c7_rf_chllp_reg[23]/NET0131  & ~n10319 ;
  assign n10345 = ~n2529 & n10319 ;
  assign n10346 = ~n2528 & n10345 ;
  assign n10347 = ~n10344 & ~n10346 ;
  assign n10348 = n8677 & n10212 ;
  assign n10349 = ~\ctl_rf_c7_rf_chllp_reg[25]/NET0131  & ~n10348 ;
  assign n10350 = ~n9789 & n10348 ;
  assign n10351 = ~n9788 & n10350 ;
  assign n10352 = ~n10349 & ~n10351 ;
  assign n10353 = ~\ctl_rf_c7_rf_chllp_reg[26]/NET0131  & ~n10348 ;
  assign n10354 = ~n9798 & n10348 ;
  assign n10355 = ~n9797 & n10354 ;
  assign n10356 = ~n10353 & ~n10355 ;
  assign n10357 = ~\ctl_rf_c7_rf_chllp_reg[27]/NET0131  & ~n10348 ;
  assign n10358 = ~n9807 & n10348 ;
  assign n10359 = ~n9806 & n10358 ;
  assign n10360 = ~n10357 & ~n10359 ;
  assign n10361 = ~\ctl_rf_c7_rf_chllp_reg[28]/NET0131  & ~n10348 ;
  assign n10362 = ~n9816 & n10348 ;
  assign n10363 = ~n9815 & n10362 ;
  assign n10364 = ~n10361 & ~n10363 ;
  assign n10365 = n8677 & n10230 ;
  assign n10366 = ~\ctl_rf_c7_rf_chllp_reg[4]/NET0131  & ~n10365 ;
  assign n10367 = ~n8714 & n10365 ;
  assign n10368 = ~n8713 & n10367 ;
  assign n10369 = ~n10366 & ~n10368 ;
  assign n10370 = ~\ctl_rf_c7_rf_chllp_reg[5]/NET0131  & ~n10365 ;
  assign n10371 = ~n8587 & n10365 ;
  assign n10372 = ~n8586 & n10371 ;
  assign n10373 = ~n10370 & ~n10372 ;
  assign n10374 = ~\ctl_rf_c7_rf_chllp_reg[6]/NET0131  & ~n10365 ;
  assign n10375 = ~n8596 & n10365 ;
  assign n10376 = ~n8595 & n10375 ;
  assign n10377 = ~n10374 & ~n10376 ;
  assign n10378 = ~\ctl_rf_c7_rf_chllp_reg[7]/NET0131  & ~n10365 ;
  assign n10379 = ~n2247 & n10365 ;
  assign n10380 = ~n2246 & n10379 ;
  assign n10381 = ~n10378 & ~n10380 ;
  assign n10382 = ~\ctl_rf_c7_rf_chllp_reg[8]/NET0131  & ~n10294 ;
  assign n10383 = ~n8781 & n10294 ;
  assign n10384 = ~n8780 & n10383 ;
  assign n10385 = ~n10382 & ~n10384 ;
  assign n10386 = ~\ctl_rf_c7_rf_chllp_reg[9]/NET0131  & ~n10294 ;
  assign n10387 = ~n8808 & n10294 ;
  assign n10388 = ~n8807 & n10387 ;
  assign n10389 = ~n10386 & ~n10388 ;
  assign n10390 = \hrdata_reg[22]_pad  & ~n4569 ;
  assign n10391 = ~n4745 & ~n8422 ;
  assign n10392 = ~n8367 & n10391 ;
  assign n10393 = n7279 & ~n7295 ;
  assign n10394 = n10273 & ~n10393 ;
  assign n10395 = ~n4573 & ~n10394 ;
  assign n10396 = ~n10392 & n10395 ;
  assign n10397 = n4573 & ~n7520 ;
  assign n10398 = ~n7506 & n10397 ;
  assign n10399 = n4569 & ~n10398 ;
  assign n10400 = ~n10396 & n10399 ;
  assign n10401 = ~n10390 & ~n10400 ;
  assign n10402 = \hrdata_reg[23]_pad  & ~n4569 ;
  assign n10403 = ~n4745 & ~n8565 ;
  assign n10404 = ~n8510 & n10403 ;
  assign n10405 = n7582 & ~n7598 ;
  assign n10406 = n10273 & ~n10405 ;
  assign n10407 = ~n4573 & ~n10406 ;
  assign n10408 = ~n10404 & n10407 ;
  assign n10409 = n4573 & ~n7839 ;
  assign n10410 = ~n7825 & n10409 ;
  assign n10411 = n4569 & ~n10410 ;
  assign n10412 = ~n10408 & n10411 ;
  assign n10413 = ~n10402 & ~n10412 ;
  assign n10414 = ~n2830 & ~n9692 ;
  assign n10415 = n8578 & n9940 ;
  assign n10416 = ~\ctl_rf_c0_rf_chllp_reg[10]/NET0131  & ~n10415 ;
  assign n10417 = ~n8759 & n10415 ;
  assign n10418 = ~n8758 & n10417 ;
  assign n10419 = ~n10416 & ~n10418 ;
  assign n10420 = ~\ctl_rf_c0_rf_chllp_reg[11]/NET0131  & ~n10415 ;
  assign n10421 = ~n8791 & n10415 ;
  assign n10422 = ~n8790 & n10421 ;
  assign n10423 = ~n10420 & ~n10422 ;
  assign n10424 = ~\ctl_rf_c0_rf_chllp_reg[12]/NET0131  & ~n10415 ;
  assign n10425 = ~n8768 & n10415 ;
  assign n10426 = ~n8767 & n10425 ;
  assign n10427 = ~n10424 & ~n10426 ;
  assign n10428 = ~\ctl_rf_c0_rf_chllp_reg[15]/NET0131  & ~n10415 ;
  assign n10429 = ~n3763 & n10415 ;
  assign n10430 = ~n3762 & n10429 ;
  assign n10431 = ~n10428 & ~n10430 ;
  assign n10432 = n8578 & n9996 ;
  assign n10433 = ~\ctl_rf_c0_rf_chllp_reg[28]/NET0131  & ~n10432 ;
  assign n10434 = ~n9816 & n10432 ;
  assign n10435 = ~n9815 & n10434 ;
  assign n10436 = ~n10433 & ~n10435 ;
  assign n10437 = n8578 & n10014 ;
  assign n10438 = ~\ctl_rf_c0_rf_chllp_reg[5]/NET0131  & ~n10437 ;
  assign n10439 = ~n8587 & n10437 ;
  assign n10440 = ~n8586 & n10439 ;
  assign n10441 = ~n10438 & ~n10440 ;
  assign n10442 = ~\ctl_rf_c0_rf_chllp_reg[6]/NET0131  & ~n10437 ;
  assign n10443 = ~n8596 & n10437 ;
  assign n10444 = ~n8595 & n10443 ;
  assign n10445 = ~n10442 & ~n10444 ;
  assign n10446 = ~\ctl_rf_c0_rf_chllp_reg[7]/NET0131  & ~n10437 ;
  assign n10447 = ~n2247 & n10437 ;
  assign n10448 = ~n2246 & n10447 ;
  assign n10449 = ~n10446 & ~n10448 ;
  assign n10450 = ~\ctl_rf_c0_rf_chllp_reg[8]/NET0131  & ~n10415 ;
  assign n10451 = ~n8781 & n10415 ;
  assign n10452 = ~n8780 & n10451 ;
  assign n10453 = ~n10450 & ~n10452 ;
  assign n10454 = ~\ctl_rf_c0_rf_chllp_reg[9]/NET0131  & ~n10415 ;
  assign n10455 = ~n8808 & n10415 ;
  assign n10456 = ~n8807 & n10455 ;
  assign n10457 = ~n10454 & ~n10456 ;
  assign n10458 = n8609 & n9940 ;
  assign n10459 = ~\ctl_rf_c2_rf_chllp_reg[10]/NET0131  & ~n10458 ;
  assign n10460 = ~n8759 & n10458 ;
  assign n10461 = ~n8758 & n10460 ;
  assign n10462 = ~n10459 & ~n10461 ;
  assign n10463 = ~\ctl_rf_c2_rf_chllp_reg[11]/NET0131  & ~n10458 ;
  assign n10464 = ~n8791 & n10458 ;
  assign n10465 = ~n8790 & n10464 ;
  assign n10466 = ~n10463 & ~n10465 ;
  assign n10467 = ~\ctl_rf_c2_rf_chllp_reg[12]/NET0131  & ~n10458 ;
  assign n10468 = ~n8768 & n10458 ;
  assign n10469 = ~n8767 & n10468 ;
  assign n10470 = ~n10467 & ~n10469 ;
  assign n10471 = ~\ctl_rf_c2_rf_chllp_reg[15]/NET0131  & ~n10458 ;
  assign n10472 = ~n3763 & n10458 ;
  assign n10473 = ~n3762 & n10472 ;
  assign n10474 = ~n10471 & ~n10473 ;
  assign n10475 = n8609 & n9966 ;
  assign n10476 = ~\ctl_rf_c2_rf_chllp_reg[21]/NET0131  & ~n10475 ;
  assign n10477 = ~n2366 & n10475 ;
  assign n10478 = ~n2365 & n10477 ;
  assign n10479 = ~n10476 & ~n10478 ;
  assign n10480 = ~\ctl_rf_c2_rf_chllp_reg[22]/NET0131  & ~n10475 ;
  assign n10481 = ~n2500 & n10475 ;
  assign n10482 = ~n2499 & n10481 ;
  assign n10483 = ~n10480 & ~n10482 ;
  assign n10484 = n8609 & n9996 ;
  assign n10485 = ~\ctl_rf_c2_rf_chllp_reg[28]/NET0131  & ~n10484 ;
  assign n10486 = ~n9816 & n10484 ;
  assign n10487 = ~n9815 & n10486 ;
  assign n10488 = ~n10485 & ~n10487 ;
  assign n10489 = n8609 & n10014 ;
  assign n10490 = ~\ctl_rf_c2_rf_chllp_reg[5]/NET0131  & ~n10489 ;
  assign n10491 = ~n8587 & n10489 ;
  assign n10492 = ~n8586 & n10491 ;
  assign n10493 = ~n10490 & ~n10492 ;
  assign n10494 = ~\ctl_rf_c2_rf_chllp_reg[6]/NET0131  & ~n10489 ;
  assign n10495 = ~n8596 & n10489 ;
  assign n10496 = ~n8595 & n10495 ;
  assign n10497 = ~n10494 & ~n10496 ;
  assign n10498 = ~\ctl_rf_c2_rf_chllp_reg[7]/NET0131  & ~n10489 ;
  assign n10499 = ~n2247 & n10489 ;
  assign n10500 = ~n2246 & n10499 ;
  assign n10501 = ~n10498 & ~n10500 ;
  assign n10502 = ~\ctl_rf_c2_rf_chllp_reg[8]/NET0131  & ~n10458 ;
  assign n10503 = ~n8781 & n10458 ;
  assign n10504 = ~n8780 & n10503 ;
  assign n10505 = ~n10502 & ~n10504 ;
  assign n10506 = ~\ctl_rf_c2_rf_chllp_reg[9]/NET0131  & ~n10458 ;
  assign n10507 = ~n8808 & n10458 ;
  assign n10508 = ~n8807 & n10507 ;
  assign n10509 = ~n10506 & ~n10508 ;
  assign n10510 = ~n9636 & ~n9653 ;
  assign n10511 = n9618 & n9635 ;
  assign n10512 = n9689 & ~n10511 ;
  assign n10513 = n10510 & n10512 ;
  assign n10514 = ~n9597 & ~n9697 ;
  assign n10515 = ~n10513 & n10514 ;
  assign n10516 = ~n9580 & n9689 ;
  assign n10517 = n9654 & n10516 ;
  assign n10518 = ~n9598 & ~n10517 ;
  assign n10519 = n9695 & ~n10518 ;
  assign n10520 = ~n10515 & n10519 ;
  assign n10521 = ~n9420 & ~n9473 ;
  assign n10522 = n9437 & n9490 ;
  assign n10523 = n10521 & ~n10522 ;
  assign n10524 = ~n9437 & ~n9490 ;
  assign n10525 = ~n9455 & ~n10524 ;
  assign n10526 = n10523 & n10525 ;
  assign n10527 = ~n9508 & ~n9712 ;
  assign n10528 = ~n10526 & n10527 ;
  assign n10529 = n9491 & ~n9525 ;
  assign n10530 = n9456 & n10529 ;
  assign n10531 = ~n9526 & ~n10530 ;
  assign n10532 = n9718 & ~n10531 ;
  assign n10533 = ~n10528 & n10532 ;
  assign n10534 = ~n10520 & ~n10533 ;
  assign n10535 = ~\ctl_rf_c0_rf_chllp_reg[13]/NET0131  & ~n10415 ;
  assign n10536 = ~n9018 & n10415 ;
  assign n10537 = ~n9017 & n10536 ;
  assign n10538 = ~n10535 & ~n10537 ;
  assign n10539 = ~\ctl_rf_c0_rf_chllp_reg[14]/NET0131  & ~n10415 ;
  assign n10540 = ~n9027 & n10415 ;
  assign n10541 = ~n9026 & n10540 ;
  assign n10542 = ~n10539 & ~n10541 ;
  assign n10543 = n8578 & n9966 ;
  assign n10544 = ~\ctl_rf_c0_rf_chllp_reg[16]/NET0131  & ~n10543 ;
  assign n10545 = ~n2680 & n10543 ;
  assign n10546 = ~n2679 & n10545 ;
  assign n10547 = ~n10544 & ~n10546 ;
  assign n10548 = ~\ctl_rf_c0_rf_chllp_reg[19]/NET0131  & ~n10543 ;
  assign n10549 = ~n2409 & n10543 ;
  assign n10550 = ~n2408 & n10549 ;
  assign n10551 = ~n10548 & ~n10550 ;
  assign n10552 = ~\ctl_rf_c0_rf_chllp_reg[25]/NET0131  & ~n10432 ;
  assign n10553 = ~n9789 & n10432 ;
  assign n10554 = ~n9788 & n10553 ;
  assign n10555 = ~n10552 & ~n10554 ;
  assign n10556 = ~\ctl_rf_c0_rf_chllp_reg[26]/NET0131  & ~n10432 ;
  assign n10557 = ~n9798 & n10432 ;
  assign n10558 = ~n9797 & n10557 ;
  assign n10559 = ~n10556 & ~n10558 ;
  assign n10560 = ~\ctl_rf_c0_rf_chllp_reg[27]/NET0131  & ~n10432 ;
  assign n10561 = ~n9807 & n10432 ;
  assign n10562 = ~n9806 & n10561 ;
  assign n10563 = ~n10560 & ~n10562 ;
  assign n10564 = ~\ctl_rf_c0_rf_chllp_reg[4]/NET0131  & ~n10437 ;
  assign n10565 = ~n8714 & n10437 ;
  assign n10566 = ~n8713 & n10565 ;
  assign n10567 = ~n10564 & ~n10566 ;
  assign n10568 = ~\ctl_rf_c1_rf_chllp_reg[20]/NET0131  & ~n9753 ;
  assign n10569 = ~n2566 & n9753 ;
  assign n10570 = ~n2565 & n10569 ;
  assign n10571 = ~n10568 & ~n10570 ;
  assign n10572 = ~\ctl_rf_c1_rf_chllp_reg[24]/NET0131  & ~n9783 ;
  assign n10573 = ~n2575 & n9783 ;
  assign n10574 = ~n2574 & n10573 ;
  assign n10575 = ~n10572 & ~n10574 ;
  assign n10576 = ~\ctl_rf_c1_rf_chllp_reg[29]/NET0131  & ~n9783 ;
  assign n10577 = \hwdata[29]_pad  & ~n2242 ;
  assign n10578 = \hwdata[5]_pad  & n2242 ;
  assign n10579 = ~n10577 & ~n10578 ;
  assign n10580 = ~n2240 & ~n10579 ;
  assign n10581 = \hwdata[13]_pad  & n2240 ;
  assign n10582 = n9783 & ~n10581 ;
  assign n10583 = ~n10580 & n10582 ;
  assign n10584 = ~n10576 & ~n10583 ;
  assign n10585 = ~\ctl_rf_c1_rf_chllp_reg[2]/NET0131  & ~n9821 ;
  assign n10586 = ~n9001 & n9821 ;
  assign n10587 = ~n9000 & n10586 ;
  assign n10588 = ~n10585 & ~n10587 ;
  assign n10589 = ~\ctl_rf_c1_rf_chllp_reg[30]/NET0131  & ~n9783 ;
  assign n10590 = \hwdata[30]_pad  & ~n2242 ;
  assign n10591 = \hwdata[6]_pad  & n2242 ;
  assign n10592 = ~n10590 & ~n10591 ;
  assign n10593 = ~n2240 & ~n10592 ;
  assign n10594 = \hwdata[14]_pad  & n2240 ;
  assign n10595 = n9783 & ~n10594 ;
  assign n10596 = ~n10593 & n10595 ;
  assign n10597 = ~n10589 & ~n10596 ;
  assign n10598 = ~\ctl_rf_c1_rf_chllp_reg[31]/NET0131  & ~n9783 ;
  assign n10599 = ~n2307 & n9783 ;
  assign n10600 = ~n2306 & n10599 ;
  assign n10601 = ~n10598 & ~n10600 ;
  assign n10602 = ~\ctl_rf_c1_rf_chllp_reg[3]/NET0131  & ~n9821 ;
  assign n10603 = ~n9044 & n9821 ;
  assign n10604 = ~n9043 & n10603 ;
  assign n10605 = ~n10602 & ~n10604 ;
  assign n10606 = ~\ctl_rf_c2_rf_chllp_reg[13]/NET0131  & ~n10458 ;
  assign n10607 = ~n9018 & n10458 ;
  assign n10608 = ~n9017 & n10607 ;
  assign n10609 = ~n10606 & ~n10608 ;
  assign n10610 = ~\ctl_rf_c2_rf_chllp_reg[14]/NET0131  & ~n10458 ;
  assign n10611 = ~n9027 & n10458 ;
  assign n10612 = ~n9026 & n10611 ;
  assign n10613 = ~n10610 & ~n10612 ;
  assign n10614 = ~\ctl_rf_c2_rf_chllp_reg[16]/NET0131  & ~n10475 ;
  assign n10615 = ~n2680 & n10475 ;
  assign n10616 = ~n2679 & n10615 ;
  assign n10617 = ~n10614 & ~n10616 ;
  assign n10618 = ~\ctl_rf_c2_rf_chllp_reg[17]/NET0131  & ~n10475 ;
  assign n10619 = ~n2260 & n10475 ;
  assign n10620 = ~n2259 & n10619 ;
  assign n10621 = ~n10618 & ~n10620 ;
  assign n10622 = ~\ctl_rf_c2_rf_chllp_reg[18]/NET0131  & ~n10475 ;
  assign n10623 = ~n2400 & n10475 ;
  assign n10624 = ~n2399 & n10623 ;
  assign n10625 = ~n10622 & ~n10624 ;
  assign n10626 = ~\ctl_rf_c2_rf_chllp_reg[19]/NET0131  & ~n10475 ;
  assign n10627 = ~n2409 & n10475 ;
  assign n10628 = ~n2408 & n10627 ;
  assign n10629 = ~n10626 & ~n10628 ;
  assign n10630 = ~\ctl_rf_c2_rf_chllp_reg[25]/NET0131  & ~n10484 ;
  assign n10631 = ~n9789 & n10484 ;
  assign n10632 = ~n9788 & n10631 ;
  assign n10633 = ~n10630 & ~n10632 ;
  assign n10634 = ~\ctl_rf_c2_rf_chllp_reg[26]/NET0131  & ~n10484 ;
  assign n10635 = ~n9798 & n10484 ;
  assign n10636 = ~n9797 & n10635 ;
  assign n10637 = ~n10634 & ~n10636 ;
  assign n10638 = ~\ctl_rf_c2_rf_chllp_reg[27]/NET0131  & ~n10484 ;
  assign n10639 = ~n9807 & n10484 ;
  assign n10640 = ~n9806 & n10639 ;
  assign n10641 = ~n10638 & ~n10640 ;
  assign n10642 = ~\ctl_rf_c2_rf_chllp_reg[4]/NET0131  & ~n10489 ;
  assign n10643 = ~n8714 & n10489 ;
  assign n10644 = ~n8713 & n10643 ;
  assign n10645 = ~n10642 & ~n10644 ;
  assign n10646 = ~\ctl_rf_c3_rf_chllp_reg[20]/NET0131  & ~n9871 ;
  assign n10647 = ~n2566 & n9871 ;
  assign n10648 = ~n2565 & n10647 ;
  assign n10649 = ~n10646 & ~n10648 ;
  assign n10650 = ~\ctl_rf_c3_rf_chllp_reg[24]/NET0131  & ~n9896 ;
  assign n10651 = ~n2575 & n9896 ;
  assign n10652 = ~n2574 & n10651 ;
  assign n10653 = ~n10650 & ~n10652 ;
  assign n10654 = ~\ctl_rf_c3_rf_chllp_reg[29]/NET0131  & ~n9896 ;
  assign n10655 = n9896 & ~n10581 ;
  assign n10656 = ~n10580 & n10655 ;
  assign n10657 = ~n10654 & ~n10656 ;
  assign n10658 = ~\ctl_rf_c3_rf_chllp_reg[2]/NET0131  & ~n9913 ;
  assign n10659 = ~n9001 & n9913 ;
  assign n10660 = ~n9000 & n10659 ;
  assign n10661 = ~n10658 & ~n10660 ;
  assign n10662 = ~\ctl_rf_c3_rf_chllp_reg[30]/NET0131  & ~n9896 ;
  assign n10663 = n9896 & ~n10594 ;
  assign n10664 = ~n10593 & n10663 ;
  assign n10665 = ~n10662 & ~n10664 ;
  assign n10666 = ~\ctl_rf_c3_rf_chllp_reg[31]/NET0131  & ~n9896 ;
  assign n10667 = ~n2307 & n9896 ;
  assign n10668 = ~n2306 & n10667 ;
  assign n10669 = ~n10666 & ~n10668 ;
  assign n10670 = ~\ctl_rf_c3_rf_chllp_reg[3]/NET0131  & ~n9913 ;
  assign n10671 = ~n9044 & n9913 ;
  assign n10672 = ~n9043 & n10671 ;
  assign n10673 = ~n10670 & ~n10672 ;
  assign n10674 = ~\ctl_rf_c4_rf_chllp_reg[20]/NET0131  & ~n9967 ;
  assign n10675 = ~n2566 & n9967 ;
  assign n10676 = ~n2565 & n10675 ;
  assign n10677 = ~n10674 & ~n10676 ;
  assign n10678 = ~\ctl_rf_c4_rf_chllp_reg[24]/NET0131  & ~n9997 ;
  assign n10679 = ~n2575 & n9997 ;
  assign n10680 = ~n2574 & n10679 ;
  assign n10681 = ~n10678 & ~n10680 ;
  assign n10682 = ~\ctl_rf_c4_rf_chllp_reg[29]/NET0131  & ~n9997 ;
  assign n10683 = n9997 & ~n10581 ;
  assign n10684 = ~n10580 & n10683 ;
  assign n10685 = ~n10682 & ~n10684 ;
  assign n10686 = ~\ctl_rf_c4_rf_chllp_reg[2]/NET0131  & ~n10015 ;
  assign n10687 = ~n9001 & n10015 ;
  assign n10688 = ~n9000 & n10687 ;
  assign n10689 = ~n10686 & ~n10688 ;
  assign n10690 = ~\ctl_rf_c4_rf_chllp_reg[30]/NET0131  & ~n9997 ;
  assign n10691 = n9997 & ~n10594 ;
  assign n10692 = ~n10593 & n10691 ;
  assign n10693 = ~n10690 & ~n10692 ;
  assign n10694 = ~\ctl_rf_c4_rf_chllp_reg[31]/NET0131  & ~n9997 ;
  assign n10695 = ~n2307 & n9997 ;
  assign n10696 = ~n2306 & n10695 ;
  assign n10697 = ~n10694 & ~n10696 ;
  assign n10698 = ~\ctl_rf_c4_rf_chllp_reg[3]/NET0131  & ~n10015 ;
  assign n10699 = ~n9044 & n10015 ;
  assign n10700 = ~n9043 & n10699 ;
  assign n10701 = ~n10698 & ~n10700 ;
  assign n10702 = ~\ctl_rf_c5_rf_chllp_reg[20]/NET0131  & ~n10065 ;
  assign n10703 = ~n2566 & n10065 ;
  assign n10704 = ~n2565 & n10703 ;
  assign n10705 = ~n10702 & ~n10704 ;
  assign n10706 = ~\ctl_rf_c5_rf_chllp_reg[24]/NET0131  & ~n10094 ;
  assign n10707 = ~n2575 & n10094 ;
  assign n10708 = ~n2574 & n10707 ;
  assign n10709 = ~n10706 & ~n10708 ;
  assign n10710 = ~\ctl_rf_c5_rf_chllp_reg[29]/NET0131  & ~n10094 ;
  assign n10711 = n10094 & ~n10581 ;
  assign n10712 = ~n10580 & n10711 ;
  assign n10713 = ~n10710 & ~n10712 ;
  assign n10714 = ~\ctl_rf_c5_rf_chllp_reg[2]/NET0131  & ~n10111 ;
  assign n10715 = ~n9001 & n10111 ;
  assign n10716 = ~n9000 & n10715 ;
  assign n10717 = ~n10714 & ~n10716 ;
  assign n10718 = ~\ctl_rf_c5_rf_chllp_reg[30]/NET0131  & ~n10094 ;
  assign n10719 = n10094 & ~n10594 ;
  assign n10720 = ~n10593 & n10719 ;
  assign n10721 = ~n10718 & ~n10720 ;
  assign n10722 = ~\ctl_rf_c5_rf_chllp_reg[31]/NET0131  & ~n10094 ;
  assign n10723 = ~n2307 & n10094 ;
  assign n10724 = ~n2306 & n10723 ;
  assign n10725 = ~n10722 & ~n10724 ;
  assign n10726 = ~\ctl_rf_c5_rf_chllp_reg[3]/NET0131  & ~n10111 ;
  assign n10727 = ~n9044 & n10111 ;
  assign n10728 = ~n9043 & n10727 ;
  assign n10729 = ~n10726 & ~n10728 ;
  assign n10730 = ~\ctl_rf_c6_rf_chllp_reg[20]/NET0131  & ~n10191 ;
  assign n10731 = ~n2566 & n10191 ;
  assign n10732 = ~n2565 & n10731 ;
  assign n10733 = ~n10730 & ~n10732 ;
  assign n10734 = ~\ctl_rf_c6_rf_chllp_reg[24]/NET0131  & ~n10213 ;
  assign n10735 = ~n2575 & n10213 ;
  assign n10736 = ~n2574 & n10735 ;
  assign n10737 = ~n10734 & ~n10736 ;
  assign n10738 = ~\ctl_rf_c6_rf_chllp_reg[29]/NET0131  & ~n10213 ;
  assign n10739 = n10213 & ~n10581 ;
  assign n10740 = ~n10580 & n10739 ;
  assign n10741 = ~n10738 & ~n10740 ;
  assign n10742 = ~\ctl_rf_c6_rf_chllp_reg[2]/NET0131  & ~n10231 ;
  assign n10743 = ~n9001 & n10231 ;
  assign n10744 = ~n9000 & n10743 ;
  assign n10745 = ~n10742 & ~n10744 ;
  assign n10746 = ~\ctl_rf_c6_rf_chllp_reg[30]/NET0131  & ~n10213 ;
  assign n10747 = n10213 & ~n10594 ;
  assign n10748 = ~n10593 & n10747 ;
  assign n10749 = ~n10746 & ~n10748 ;
  assign n10750 = ~\ctl_rf_c6_rf_chllp_reg[31]/NET0131  & ~n10213 ;
  assign n10751 = ~n2307 & n10213 ;
  assign n10752 = ~n2306 & n10751 ;
  assign n10753 = ~n10750 & ~n10752 ;
  assign n10754 = ~\ctl_rf_c6_rf_chllp_reg[3]/NET0131  & ~n10231 ;
  assign n10755 = ~n9044 & n10231 ;
  assign n10756 = ~n9043 & n10755 ;
  assign n10757 = ~n10754 & ~n10756 ;
  assign n10758 = ~\ctl_rf_c7_rf_chllp_reg[20]/NET0131  & ~n10319 ;
  assign n10759 = ~n2566 & n10319 ;
  assign n10760 = ~n2565 & n10759 ;
  assign n10761 = ~n10758 & ~n10760 ;
  assign n10762 = ~\ctl_rf_c7_rf_chllp_reg[24]/NET0131  & ~n10348 ;
  assign n10763 = ~n2575 & n10348 ;
  assign n10764 = ~n2574 & n10763 ;
  assign n10765 = ~n10762 & ~n10764 ;
  assign n10766 = ~\ctl_rf_c7_rf_chllp_reg[29]/NET0131  & ~n10348 ;
  assign n10767 = n10348 & ~n10581 ;
  assign n10768 = ~n10580 & n10767 ;
  assign n10769 = ~n10766 & ~n10768 ;
  assign n10770 = ~\ctl_rf_c7_rf_chllp_reg[2]/NET0131  & ~n10365 ;
  assign n10771 = ~n9001 & n10365 ;
  assign n10772 = ~n9000 & n10771 ;
  assign n10773 = ~n10770 & ~n10772 ;
  assign n10774 = ~\ctl_rf_c7_rf_chllp_reg[30]/NET0131  & ~n10348 ;
  assign n10775 = n10348 & ~n10594 ;
  assign n10776 = ~n10593 & n10775 ;
  assign n10777 = ~n10774 & ~n10776 ;
  assign n10778 = ~\ctl_rf_c7_rf_chllp_reg[31]/NET0131  & ~n10348 ;
  assign n10779 = ~n2307 & n10348 ;
  assign n10780 = ~n2306 & n10779 ;
  assign n10781 = ~n10778 & ~n10780 ;
  assign n10782 = ~\ctl_rf_c7_rf_chllp_reg[3]/NET0131  & ~n10365 ;
  assign n10783 = ~n9044 & n10365 ;
  assign n10784 = ~n9043 & n10783 ;
  assign n10785 = ~n10782 & ~n10784 ;
  assign n10786 = ~\ctl_rf_c0_rf_chllp_reg[23]/NET0131  & ~n10543 ;
  assign n10787 = ~n2529 & n10543 ;
  assign n10788 = ~n2528 & n10787 ;
  assign n10789 = ~n10786 & ~n10788 ;
  assign n10790 = ~\ctl_rf_c2_rf_chllp_reg[23]/NET0131  & ~n10475 ;
  assign n10791 = ~n2529 & n10475 ;
  assign n10792 = ~n2528 & n10791 ;
  assign n10793 = ~n10790 & ~n10792 ;
  assign n10794 = \de_de_st_reg[1]/NET0131  & \de_st_rd_msk_reg/NET0131  ;
  assign n10795 = \ch_sel_arb_chcsr_reg_reg[17]/NET0131  & n10794 ;
  assign n10796 = \ch_sel_arb_chcsr_reg_reg[15]/NET0131  & \ch_sel_arb_chcsr_reg_reg[16]/NET0131  ;
  assign n10797 = n10795 & n10796 ;
  assign n10798 = \de_bst_cnt_reg[8]/NET0131  & ~n10794 ;
  assign n10799 = ~n10797 & ~n10798 ;
  assign n10800 = ~\ctl_rf_c0_rf_chllp_reg[20]/NET0131  & ~n10543 ;
  assign n10801 = ~n2566 & n10543 ;
  assign n10802 = ~n2565 & n10801 ;
  assign n10803 = ~n10800 & ~n10802 ;
  assign n10804 = ~\ctl_rf_c0_rf_chllp_reg[24]/NET0131  & ~n10432 ;
  assign n10805 = ~n2575 & n10432 ;
  assign n10806 = ~n2574 & n10805 ;
  assign n10807 = ~n10804 & ~n10806 ;
  assign n10808 = ~\ctl_rf_c0_rf_chllp_reg[29]/NET0131  & ~n10432 ;
  assign n10809 = n10432 & ~n10581 ;
  assign n10810 = ~n10580 & n10809 ;
  assign n10811 = ~n10808 & ~n10810 ;
  assign n10812 = ~\ctl_rf_c0_rf_chllp_reg[2]/NET0131  & ~n10437 ;
  assign n10813 = ~n9001 & n10437 ;
  assign n10814 = ~n9000 & n10813 ;
  assign n10815 = ~n10812 & ~n10814 ;
  assign n10816 = ~\ctl_rf_c0_rf_chllp_reg[30]/NET0131  & ~n10432 ;
  assign n10817 = n10432 & ~n10594 ;
  assign n10818 = ~n10593 & n10817 ;
  assign n10819 = ~n10816 & ~n10818 ;
  assign n10820 = ~\ctl_rf_c0_rf_chllp_reg[31]/NET0131  & ~n10432 ;
  assign n10821 = ~n2307 & n10432 ;
  assign n10822 = ~n2306 & n10821 ;
  assign n10823 = ~n10820 & ~n10822 ;
  assign n10824 = ~\ctl_rf_c0_rf_chllp_reg[3]/NET0131  & ~n10437 ;
  assign n10825 = ~n9044 & n10437 ;
  assign n10826 = ~n9043 & n10825 ;
  assign n10827 = ~n10824 & ~n10826 ;
  assign n10828 = ~\ctl_rf_c2_rf_chllp_reg[20]/NET0131  & ~n10475 ;
  assign n10829 = ~n2566 & n10475 ;
  assign n10830 = ~n2565 & n10829 ;
  assign n10831 = ~n10828 & ~n10830 ;
  assign n10832 = ~\ctl_rf_c2_rf_chllp_reg[29]/NET0131  & ~n10484 ;
  assign n10833 = n10484 & ~n10581 ;
  assign n10834 = ~n10580 & n10833 ;
  assign n10835 = ~n10832 & ~n10834 ;
  assign n10836 = ~\ctl_rf_c2_rf_chllp_reg[2]/NET0131  & ~n10489 ;
  assign n10837 = ~n9001 & n10489 ;
  assign n10838 = ~n9000 & n10837 ;
  assign n10839 = ~n10836 & ~n10838 ;
  assign n10840 = ~\ctl_rf_c2_rf_chllp_reg[30]/NET0131  & ~n10484 ;
  assign n10841 = n10484 & ~n10594 ;
  assign n10842 = ~n10593 & n10841 ;
  assign n10843 = ~n10840 & ~n10842 ;
  assign n10844 = ~\ctl_rf_c2_rf_chllp_reg[31]/NET0131  & ~n10484 ;
  assign n10845 = ~n2307 & n10484 ;
  assign n10846 = ~n2306 & n10845 ;
  assign n10847 = ~n10844 & ~n10846 ;
  assign n10848 = ~\ctl_rf_c2_rf_chllp_reg[3]/NET0131  & ~n10489 ;
  assign n10849 = ~n9044 & n10489 ;
  assign n10850 = ~n9043 & n10849 ;
  assign n10851 = ~n10848 & ~n10850 ;
  assign n10852 = \h1size[1]_pad  & ~n3493 ;
  assign n10853 = n3491 & n10852 ;
  assign n10854 = \ch_sel_arb_chcsr_reg_reg[12]/NET0131  & \ch_sel_arb_chcsr_reg_reg[2]/NET0131  ;
  assign n10855 = ~n2815 & n10854 ;
  assign n10856 = n3487 & n10855 ;
  assign n10857 = \ch_sel_arb_chcsr_reg_reg[9]/NET0131  & ~\de_m1_is_llp_reg/NET0131  ;
  assign n10858 = n3486 & n10857 ;
  assign n10859 = ~n2816 & n10858 ;
  assign n10860 = ~n3490 & ~n10859 ;
  assign n10861 = ~n10856 & n10860 ;
  assign n10862 = ~n10853 & n10861 ;
  assign n10863 = ~\de_m1_arb_st_reg[1]/NET0131  & ~n10862 ;
  assign n10864 = \ahb_slv_slv_sz_d1o_reg[1]/NET0131  & \de_m1_arb_st_reg[1]/NET0131  ;
  assign n10865 = ~n10863 & ~n10864 ;
  assign n10866 = ~\de_m1_arb_st_reg[1]/NET0131  & ~n2801 ;
  assign n10867 = n10510 & ~n10511 ;
  assign n10868 = ~n9688 & ~n9699 ;
  assign n10869 = ~n10867 & n10868 ;
  assign n10870 = ~n9653 & ~n9671 ;
  assign n10871 = n9636 & n10870 ;
  assign n10872 = ~n9689 & ~n10871 ;
  assign n10873 = ~n10869 & ~n10872 ;
  assign n10874 = n9600 & n10873 ;
  assign n10875 = n10523 & ~n10524 ;
  assign n10876 = n9420 & n9473 ;
  assign n10877 = ~n10521 & n10524 ;
  assign n10878 = ~n10876 & n10877 ;
  assign n10879 = ~n10875 & ~n10878 ;
  assign n10880 = ~n9455 & n9526 ;
  assign n10881 = ~n9545 & n10880 ;
  assign n10882 = ~n9528 & n10881 ;
  assign n10883 = ~n10879 & n10882 ;
  assign n10884 = ~n10874 & ~n10883 ;
  assign n10885 = \de_de_st_reg[5]/NET0131  & ~\de_m1_arb_st_reg[1]/NET0131  ;
  assign n10886 = ~n2801 & n10885 ;
  assign n10887 = \de_m1_arb_st_reg[0]/NET0131  & ~n10886 ;
  assign n10888 = ~n2801 & n2914 ;
  assign n10889 = n4540 & n10888 ;
  assign n10890 = ~n10887 & ~n10889 ;
  assign n10891 = \hrdata_reg[10]_pad  & ~n4569 ;
  assign n10892 = ~n4745 & n5881 ;
  assign n10893 = n5854 & n10892 ;
  assign n10894 = ~n5145 & ~n10893 ;
  assign n10895 = ~n4573 & ~n10894 ;
  assign n10896 = ~n4573 & n4745 ;
  assign n10897 = ~n10155 & n10896 ;
  assign n10898 = ~n10895 & ~n10897 ;
  assign n10899 = n4573 & n5936 ;
  assign n10900 = n4573 & ~n5993 ;
  assign n10901 = n5977 & n10900 ;
  assign n10902 = ~n10899 & ~n10901 ;
  assign n10903 = n4569 & n10902 ;
  assign n10904 = n10898 & n10903 ;
  assign n10905 = ~n10891 & ~n10904 ;
  assign n10906 = \hrdata_reg[11]_pad  & ~n4569 ;
  assign n10907 = ~n4745 & n6226 ;
  assign n10908 = n6199 & n10907 ;
  assign n10909 = ~n5145 & ~n10908 ;
  assign n10910 = ~n4573 & ~n10909 ;
  assign n10911 = ~n10261 & n10896 ;
  assign n10912 = ~n10910 & ~n10911 ;
  assign n10913 = n4573 & n6281 ;
  assign n10914 = n4573 & ~n6338 ;
  assign n10915 = n6322 & n10914 ;
  assign n10916 = ~n10913 & ~n10915 ;
  assign n10917 = n4569 & n10916 ;
  assign n10918 = n10912 & n10917 ;
  assign n10919 = ~n10906 & ~n10918 ;
  assign n10920 = \hrdata_reg[12]_pad  & ~n4569 ;
  assign n10921 = n4573 & n6584 ;
  assign n10922 = n4573 & ~n6641 ;
  assign n10923 = n6625 & n10922 ;
  assign n10924 = ~n10921 & ~n10923 ;
  assign n10925 = n4569 & n10924 ;
  assign n10926 = ~n10920 & ~n10925 ;
  assign n10927 = n4745 & ~n8134 ;
  assign n10928 = ~n8079 & n10927 ;
  assign n10929 = ~n4573 & ~n10928 ;
  assign n10930 = \haddr[8]_pad  & ~n4745 ;
  assign n10931 = ~n10272 & n10930 ;
  assign n10932 = ~n10920 & ~n10931 ;
  assign n10933 = n10929 & n10932 ;
  assign n10934 = ~n10926 & ~n10933 ;
  assign n10935 = \hrdata_reg[13]_pad  & ~n4569 ;
  assign n10936 = n4573 & n6887 ;
  assign n10937 = n4573 & ~n6944 ;
  assign n10938 = n6928 & n10937 ;
  assign n10939 = ~n10936 & ~n10938 ;
  assign n10940 = n4569 & n10939 ;
  assign n10941 = ~n10935 & ~n10940 ;
  assign n10942 = n4745 & ~n8278 ;
  assign n10943 = ~n8223 & n10942 ;
  assign n10944 = ~n4573 & ~n10943 ;
  assign n10945 = ~n10285 & n10930 ;
  assign n10946 = ~n10935 & ~n10945 ;
  assign n10947 = n10944 & n10946 ;
  assign n10948 = ~n10941 & ~n10947 ;
  assign n10949 = \hrdata_reg[14]_pad  & ~n4569 ;
  assign n10950 = n4573 & n7350 ;
  assign n10951 = n4573 & ~n7407 ;
  assign n10952 = n7391 & n10951 ;
  assign n10953 = ~n10950 & ~n10952 ;
  assign n10954 = n4569 & n10953 ;
  assign n10955 = ~n10949 & ~n10954 ;
  assign n10956 = n4745 & ~n8422 ;
  assign n10957 = ~n8367 & n10956 ;
  assign n10958 = ~n4573 & ~n10957 ;
  assign n10959 = ~n10393 & n10930 ;
  assign n10960 = ~n10949 & ~n10959 ;
  assign n10961 = n10958 & n10960 ;
  assign n10962 = ~n10955 & ~n10961 ;
  assign n10963 = \hrdata_reg[15]_pad  & ~n4569 ;
  assign n10964 = n4569 & ~n7727 ;
  assign n10965 = ~n7677 & n10964 ;
  assign n10966 = ~n7065 & ~n10965 ;
  assign n10967 = ~n10963 & n10966 ;
  assign n10968 = n4745 & ~n8565 ;
  assign n10969 = ~n8510 & n10968 ;
  assign n10970 = ~n4573 & ~n10969 ;
  assign n10971 = ~n10405 & n10930 ;
  assign n10972 = ~n10963 & ~n10971 ;
  assign n10973 = n10970 & n10972 ;
  assign n10974 = ~n10967 & ~n10973 ;
  assign n10975 = \hrdata_reg[9]_pad  & ~n4569 ;
  assign n10976 = ~n4745 & n5771 ;
  assign n10977 = n5744 & n10976 ;
  assign n10978 = ~n5145 & ~n10977 ;
  assign n10979 = ~n4573 & ~n10978 ;
  assign n10980 = ~n10129 & n10896 ;
  assign n10981 = ~n10979 & ~n10980 ;
  assign n10982 = n4573 & n5479 ;
  assign n10983 = n4573 & ~n5536 ;
  assign n10984 = n5520 & n10983 ;
  assign n10985 = ~n10982 & ~n10984 ;
  assign n10986 = n4569 & n10985 ;
  assign n10987 = n10981 & n10986 ;
  assign n10988 = ~n10975 & ~n10987 ;
  assign n10989 = \ahb_slv_slv_sz_d1o_reg[0]/NET0131  & \de_m1_arb_st_reg[1]/NET0131  ;
  assign n10990 = \de_m1_arb_st_reg[1]/NET0131  & ~n10989 ;
  assign n10991 = \h1size[0]_pad  & ~n3493 ;
  assign n10992 = n3491 & n10991 ;
  assign n10993 = \ch_sel_arb_chcsr_reg_reg[8]/NET0131  & ~\de_m1_is_llp_reg/NET0131  ;
  assign n10994 = n3486 & n10993 ;
  assign n10995 = ~n2816 & n10994 ;
  assign n10996 = \ch_sel_arb_chcsr_reg_reg[11]/NET0131  & \ch_sel_arb_chcsr_reg_reg[2]/NET0131  ;
  assign n10997 = ~n2815 & n10996 ;
  assign n10998 = n3487 & n10997 ;
  assign n10999 = ~n10995 & ~n10998 ;
  assign n11000 = ~n10989 & n10999 ;
  assign n11001 = ~n10992 & n11000 ;
  assign n11002 = ~n10990 & ~n11001 ;
  assign n11003 = \ahb_mst0_m0_m1_diff_tx_reg/NET0131  & ~\ch_sel_arb_chcsr_reg_reg[1]/NET0131  ;
  assign n11004 = ~\de_m0_is_llp_reg/NET0131  & ~n11003 ;
  assign n11005 = n2937 & n11004 ;
  assign n11006 = \de_m0_is_llp_reg/NET0131  & ~n11003 ;
  assign n11007 = ~n2937 & n11006 ;
  assign n11008 = ~n11005 & ~n11007 ;
  assign n11009 = ~\de_m0_is_llp_reg/NET0131  & n11003 ;
  assign n11010 = ~n2937 & n11009 ;
  assign n11011 = \ahb_mst0_hsizeo_reg[1]/NET0131  & ~n11010 ;
  assign n11012 = n11008 & n11011 ;
  assign n11013 = \ch_sel_arb_chcsr_reg_reg[9]/NET0131  & ~\de_m0_is_llp_reg/NET0131  ;
  assign n11014 = n11003 & n11013 ;
  assign n11015 = ~n2937 & n11014 ;
  assign n11016 = \ch_sel_arb_chcsr_reg_reg[12]/NET0131  & ~\ch_sel_arb_chcsr_reg_reg[2]/NET0131  ;
  assign n11017 = ~n2815 & n11016 ;
  assign n11018 = n11004 & n11017 ;
  assign n11019 = ~n11007 & ~n11018 ;
  assign n11020 = ~n11015 & n11019 ;
  assign n11021 = ~n11012 & n11020 ;
  assign n11022 = \ahb_slv_br_st_reg[2]/NET0131  & n2830 ;
  assign n11023 = \ahb_slv_br_st_reg[2]/NET0131  & n2764 ;
  assign n11024 = n2798 & n11023 ;
  assign n11025 = ~n11022 & ~n11024 ;
  assign n11026 = hreadyin_pad & hsel_br_pad ;
  assign n11027 = ~\htrans[0]_pad  & \htrans[1]_pad  ;
  assign n11028 = n11026 & n11027 ;
  assign n11029 = ~\ahb_slv_br_st_reg[2]/NET0131  & ~hreadyout_br_pad ;
  assign n11030 = ~\hresp_br[0]_pad  & \hresp_br[1]_pad  ;
  assign n11031 = \hresp_br[0]_pad  & ~\hresp_br[1]_pad  ;
  assign n11032 = ~n11030 & ~n11031 ;
  assign n11033 = n11029 & n11032 ;
  assign n11034 = hreadyout_br_pad & hsel_br_pad ;
  assign n11035 = \htrans[0]_pad  & \htrans[1]_pad  ;
  assign n11036 = n11034 & n11035 ;
  assign n11037 = ~\ahb_slv_br_st_reg[1]/NET0131  & ~n11036 ;
  assign n11038 = ~n11033 & n11037 ;
  assign n11039 = ~n11028 & n11038 ;
  assign n11040 = n11025 & n11039 ;
  assign n11041 = ~\ch_sel_arb_chcsr_reg_reg[17]/NET0131  & n10794 ;
  assign n11042 = ~\ch_sel_arb_chcsr_reg_reg[15]/NET0131  & ~\ch_sel_arb_chcsr_reg_reg[16]/NET0131  ;
  assign n11043 = n11041 & n11042 ;
  assign n11044 = \de_bst_cnt_reg[0]/NET0131  & ~n10794 ;
  assign n11045 = ~n11043 & ~n11044 ;
  assign n11046 = \de_bst_cnt_reg[2]/NET0131  & ~n10794 ;
  assign n11047 = \ch_sel_arb_chcsr_reg_reg[15]/NET0131  & ~\ch_sel_arb_chcsr_reg_reg[16]/NET0131  ;
  assign n11048 = n11041 & n11047 ;
  assign n11049 = ~n11046 & ~n11048 ;
  assign n11050 = \de_bst_cnt_reg[3]/NET0131  & ~n10794 ;
  assign n11051 = ~\ch_sel_arb_chcsr_reg_reg[15]/NET0131  & \ch_sel_arb_chcsr_reg_reg[16]/NET0131  ;
  assign n11052 = n11041 & n11051 ;
  assign n11053 = ~n11050 & ~n11052 ;
  assign n11054 = \de_bst_cnt_reg[4]/NET0131  & ~n10794 ;
  assign n11055 = n10796 & n11041 ;
  assign n11056 = ~n11054 & ~n11055 ;
  assign n11057 = \de_bst_cnt_reg[5]/NET0131  & ~n10794 ;
  assign n11058 = n10795 & n11042 ;
  assign n11059 = ~n11057 & ~n11058 ;
  assign n11060 = n10795 & n11051 ;
  assign n11061 = \de_bst_cnt_reg[7]/NET0131  & ~n10794 ;
  assign n11062 = ~n11060 & ~n11061 ;
  assign n11063 = n10795 & n11047 ;
  assign n11064 = \de_bst_cnt_reg[6]/NET0131  & ~n10794 ;
  assign n11065 = ~n11063 & ~n11064 ;
  assign n11066 = \ahb_mst0_hsizeo_reg[0]/NET0131  & ~n11010 ;
  assign n11067 = n11008 & n11066 ;
  assign n11068 = \ch_sel_arb_chcsr_reg_reg[8]/NET0131  & ~\de_m0_is_llp_reg/NET0131  ;
  assign n11069 = n11003 & n11068 ;
  assign n11070 = ~n2937 & n11069 ;
  assign n11071 = \ch_sel_arb_chcsr_reg_reg[11]/NET0131  & ~\ch_sel_arb_chcsr_reg_reg[2]/NET0131  ;
  assign n11072 = ~n2815 & n11071 ;
  assign n11073 = n11004 & n11072 ;
  assign n11074 = ~n11070 & ~n11073 ;
  assign n11075 = ~n11067 & n11074 ;
  assign n11076 = \ahb_mst0_hsizeo_reg[2]/NET0131  & ~n11010 ;
  assign n11077 = n11008 & n11076 ;
  assign n11078 = \ch_sel_arb_chcsr_reg_reg[13]/NET0131  & ~\ch_sel_arb_chcsr_reg_reg[2]/NET0131  ;
  assign n11079 = ~n2815 & n11078 ;
  assign n11080 = n11004 & n11079 ;
  assign n11081 = \ch_sel_arb_chcsr_reg_reg[10]/NET0131  & ~\de_m0_is_llp_reg/NET0131  ;
  assign n11082 = n11003 & n11081 ;
  assign n11083 = ~n2937 & n11082 ;
  assign n11084 = ~n11080 & ~n11083 ;
  assign n11085 = ~n11077 & n11084 ;
  assign n11086 = \ch_sel_arb_chcsr_reg_reg[2]/NET0131  & \de_de_st_reg[1]/NET0131  ;
  assign n11087 = ~\de_m1_arb_st_reg[1]/NET0131  & ~n2826 ;
  assign n11088 = ~n11086 & n11087 ;
  assign n11089 = ~n2830 & ~n11088 ;
  assign n11090 = ~n2799 & n11089 ;
  assign n11091 = \h1write_pad  & ~n11090 ;
  assign n11092 = \ahb_slv_slv_wr_d1o_reg/NET0131  & \de_m1_arb_st_reg[1]/NET0131  ;
  assign n11093 = ~\ch_sel_arb_chcsr_reg_reg[2]/NET0131  & ~\de_m1_arb_st_reg[1]/NET0131  ;
  assign n11094 = n3486 & n11093 ;
  assign n11095 = ~n11092 & ~n11094 ;
  assign n11096 = ~n2830 & ~n11095 ;
  assign n11097 = ~n2799 & n11096 ;
  assign n11098 = ~n11091 & ~n11097 ;
  assign n11099 = \ch_sel_arb_chcsr_reg_reg[19]/NET0131  & ~\de_m1_arb_st_reg[1]/NET0131  ;
  assign n11100 = \ahb_slv_slv_pt_d1o_reg[2]/NET0131  & \de_m1_arb_st_reg[1]/NET0131  ;
  assign n11101 = ~n11099 & ~n11100 ;
  assign n11102 = \ch_sel_arb_chcsr_reg_reg[20]/NET0131  & ~\de_m1_arb_st_reg[1]/NET0131  ;
  assign n11103 = \ahb_slv_slv_pt_d1o_reg[3]/NET0131  & \de_m1_arb_st_reg[1]/NET0131  ;
  assign n11104 = ~n11102 & ~n11103 ;
  assign n11105 = \ch_sel_arb_chcsr_reg_reg[18]/NET0131  & ~\de_m1_arb_st_reg[1]/NET0131  ;
  assign n11106 = \ahb_slv_slv_pt_d1o_reg[1]/NET0131  & \de_m1_arb_st_reg[1]/NET0131  ;
  assign n11107 = ~n11105 & ~n11106 ;
  assign n11108 = ~n3762 & ~n3763 ;
  assign n11109 = \ctl_rf_be_d1_reg[2]/P0001  & n4065 ;
  assign n11110 = n2231 & n11109 ;
  assign n11111 = ~n11108 & n11110 ;
  assign n11112 = n5173 & ~n11110 ;
  assign n11113 = n3776 & n11112 ;
  assign n11114 = ~n11111 & ~n11113 ;
  assign n11115 = \ctl_rf_be_d1_reg[2]/P0001  & n3756 ;
  assign n11116 = n2311 & n11115 ;
  assign n11117 = ~n11108 & n11116 ;
  assign n11118 = n5173 & ~n11116 ;
  assign n11119 = n3792 & n11118 ;
  assign n11120 = ~n11117 & ~n11119 ;
  assign n11121 = n2311 & n11109 ;
  assign n11122 = ~n11108 & n11121 ;
  assign n11123 = n5173 & ~n11121 ;
  assign n11124 = n3794 & n11123 ;
  assign n11125 = ~n11122 & ~n11124 ;
  assign n11126 = n2231 & n11115 ;
  assign n11127 = ~n11108 & n11126 ;
  assign n11128 = n5173 & ~n11126 ;
  assign n11129 = n3783 & n11128 ;
  assign n11130 = ~n11127 & ~n11129 ;
  assign n11131 = n2317 & n11115 ;
  assign n11132 = ~n11108 & n11131 ;
  assign n11133 = n5173 & ~n11131 ;
  assign n11134 = n3778 & n11133 ;
  assign n11135 = ~n11132 & ~n11134 ;
  assign n11136 = n2317 & n11109 ;
  assign n11137 = ~n11108 & n11136 ;
  assign n11138 = n5173 & ~n11136 ;
  assign n11139 = n3787 & n11138 ;
  assign n11140 = ~n11137 & ~n11139 ;
  assign n11141 = n2324 & n11115 ;
  assign n11142 = ~n11108 & n11141 ;
  assign n11143 = n5173 & ~n11141 ;
  assign n11144 = n3789 & n11143 ;
  assign n11145 = ~n11142 & ~n11144 ;
  assign n11146 = n2324 & n11109 ;
  assign n11147 = ~n11108 & n11146 ;
  assign n11148 = n5173 & ~n11146 ;
  assign n11149 = n3781 & n11148 ;
  assign n11150 = ~n11147 & ~n11149 ;
  assign n11151 = ~\ahb_slv_br_st_reg[2]/NET0131  & \ahb_slv_slv_br_req_reg/NET0131  ;
  assign n11152 = ~n11028 & ~n11151 ;
  assign n11153 = ~n2913 & ~n11028 ;
  assign n11154 = n2881 & n11153 ;
  assign n11155 = ~n11152 & ~n11154 ;
  assign n11156 = ~\de_de_st_reg[5]/NET0131  & \de_m1_is_llp_reg/NET0131  ;
  assign n11157 = ~\de_de_st_reg[6]/NET0131  & ~n11156 ;
  assign n11158 = \ctl_rf_c2_rf_chllp_reg[0]/P0002  & n2983 ;
  assign n11159 = n3024 & n11158 ;
  assign n11160 = \ctl_rf_c0_rf_chllp_reg[0]/P0002  & n2983 ;
  assign n11161 = n3050 & n11160 ;
  assign n11162 = \ctl_rf_c5_rf_chllp_reg[0]/P0002  & ~n2983 ;
  assign n11163 = n2999 & n11162 ;
  assign n11164 = ~n11161 & ~n11163 ;
  assign n11165 = ~n11159 & n11164 ;
  assign n11166 = \ctl_rf_c6_rf_chllp_reg[0]/P0002  & n2983 ;
  assign n11167 = n3011 & n11166 ;
  assign n11168 = \de_de_st_reg[6]/NET0131  & ~n11167 ;
  assign n11169 = \ctl_rf_c4_rf_chllp_reg[0]/P0002  & n2983 ;
  assign n11170 = n2999 & n11169 ;
  assign n11171 = \ctl_rf_c3_rf_chllp_reg[0]/P0002  & ~n2983 ;
  assign n11172 = n3024 & n11171 ;
  assign n11173 = ~n11170 & ~n11172 ;
  assign n11174 = \ctl_rf_c1_rf_chllp_reg[0]/P0002  & ~n2983 ;
  assign n11175 = n3050 & n11174 ;
  assign n11176 = \ctl_rf_c7_rf_chllp_reg[0]/P0002  & ~n2983 ;
  assign n11177 = n3011 & n11176 ;
  assign n11178 = ~n11175 & ~n11177 ;
  assign n11179 = n11173 & n11178 ;
  assign n11180 = n11168 & n11179 ;
  assign n11181 = n11165 & n11180 ;
  assign n11182 = ~n11157 & ~n11181 ;
  assign n11183 = ~\ahb_slv_br_st_reg[0]/NET0131  & ~\ahb_slv_br_st_reg[1]/NET0131  ;
  assign n11184 = \ahb_slv_br_st_reg[2]/NET0131  & n11183 ;
  assign n11185 = ~\ahb_slv_br_st_reg[0]/NET0131  & \ahb_slv_br_st_reg[1]/NET0131  ;
  assign n11186 = ~\ahb_slv_br_st_reg[2]/NET0131  & n11185 ;
  assign n11187 = \ahb_slv_br_st_reg[0]/NET0131  & ~\ahb_slv_br_st_reg[2]/NET0131  ;
  assign n11188 = ~\ahb_slv_br_st_reg[1]/NET0131  & n11187 ;
  assign n11189 = n11028 & n11188 ;
  assign n11190 = ~n11186 & ~n11189 ;
  assign n11191 = ~n11184 & n11190 ;
  assign n11192 = ~n2913 & n11190 ;
  assign n11193 = n2881 & n11192 ;
  assign n11194 = ~n11191 & ~n11193 ;
  assign n11195 = \de_m0_is_llp_reg/NET0131  & n4472 ;
  assign n11196 = ~n11181 & ~n11195 ;
  assign n11197 = \ahb_slv_br_st_reg[0]/NET0131  & ~\ahb_slv_br_st_reg[1]/NET0131  ;
  assign n11198 = ~\ahb_slv_br_st_reg[2]/NET0131  & n11197 ;
  assign n11199 = n11028 & n11198 ;
  assign n11200 = ~n11186 & ~n11199 ;
  assign n11201 = ~\ahb_mst1_mx_cmd_st_reg[0]/NET0131  & n2802 ;
  assign n11202 = \ahb_mst1_mx_cmd_st_reg[1]/NET0131  & ~n2830 ;
  assign n11203 = n11201 & n11202 ;
  assign n11204 = ~n2799 & n11203 ;
  assign n11205 = ~n11199 & n11204 ;
  assign n11206 = ~n11200 & ~n11205 ;
  assign n11207 = n2881 & ~n2913 ;
  assign n11208 = n11184 & ~n11207 ;
  assign n11209 = n11186 & n11204 ;
  assign n11210 = ~n11208 & ~n11209 ;
  assign n11211 = \ctl_rf_c0_rf_chllp_on_reg/NET0131  & \de_de_st_reg[5]/NET0131  ;
  assign n11212 = n2983 & n11211 ;
  assign n11213 = n3050 & n11212 ;
  assign n11214 = ~\ctl_rf_c0_rf_chabt_reg/NET0131  & ~n2814 ;
  assign n11215 = \ctl_rf_c0_rf_chllp_cnt_reg[0]/NET0131  & \ctl_rf_c0_rf_chllp_cnt_reg[1]/NET0131  ;
  assign n11216 = ~n11214 & n11215 ;
  assign n11217 = n11213 & n11216 ;
  assign n11218 = \ctl_rf_c0_rf_chllp_cnt_reg[2]/NET0131  & n11217 ;
  assign n11219 = \ctl_rf_be_d1_reg[0]/P0001  & ~\ctl_rf_c0_rf_ch_en_reg/NET0131  ;
  assign n11220 = ~n3772 & n11219 ;
  assign n11221 = ~n4173 & n11220 ;
  assign n11222 = ~\ctl_rf_c0_rf_chllp_cnt_reg[2]/NET0131  & ~n11217 ;
  assign n11223 = ~n11221 & ~n11222 ;
  assign n11224 = ~n11218 & n11223 ;
  assign n11225 = ~\ctl_rf_c0_rf_chllp_cnt_reg[3]/NET0131  & ~n11218 ;
  assign n11226 = \ctl_rf_c0_rf_chllp_cnt_reg[2]/NET0131  & \ctl_rf_c0_rf_chllp_cnt_reg[3]/NET0131  ;
  assign n11227 = n11217 & n11226 ;
  assign n11228 = ~n11221 & ~n11227 ;
  assign n11229 = ~n11225 & n11228 ;
  assign n11230 = \ctl_rf_c1_rf_chllp_on_reg/NET0131  & \de_de_st_reg[5]/NET0131  ;
  assign n11231 = ~n2983 & n11230 ;
  assign n11232 = n3050 & n11231 ;
  assign n11233 = ~\ctl_rf_c1_rf_chabt_reg/NET0131  & ~n2814 ;
  assign n11234 = \ctl_rf_c1_rf_chllp_cnt_reg[0]/NET0131  & \ctl_rf_c1_rf_chllp_cnt_reg[1]/NET0131  ;
  assign n11235 = ~n11233 & n11234 ;
  assign n11236 = n11232 & n11235 ;
  assign n11237 = \ctl_rf_c1_rf_chllp_cnt_reg[2]/NET0131  & n11236 ;
  assign n11238 = \ctl_rf_be_d1_reg[0]/P0001  & ~\ctl_rf_c1_rf_ch_en_reg/NET0131  ;
  assign n11239 = ~n3772 & n11238 ;
  assign n11240 = ~n4122 & n11239 ;
  assign n11241 = ~\ctl_rf_c1_rf_chllp_cnt_reg[2]/NET0131  & ~n11236 ;
  assign n11242 = ~n11240 & ~n11241 ;
  assign n11243 = ~n11237 & n11242 ;
  assign n11244 = ~\ctl_rf_c1_rf_chllp_cnt_reg[3]/NET0131  & ~n11237 ;
  assign n11245 = \ctl_rf_c1_rf_chllp_cnt_reg[2]/NET0131  & \ctl_rf_c1_rf_chllp_cnt_reg[3]/NET0131  ;
  assign n11246 = n11236 & n11245 ;
  assign n11247 = ~n11240 & ~n11246 ;
  assign n11248 = ~n11244 & n11247 ;
  assign n11249 = \ctl_rf_c2_rf_chllp_on_reg/NET0131  & \de_de_st_reg[5]/NET0131  ;
  assign n11250 = n2983 & n11249 ;
  assign n11251 = n3024 & n11250 ;
  assign n11252 = ~\ctl_rf_c2_rf_chabt_reg/NET0131  & ~n2814 ;
  assign n11253 = \ctl_rf_c2_rf_chllp_cnt_reg[0]/NET0131  & \ctl_rf_c2_rf_chllp_cnt_reg[1]/NET0131  ;
  assign n11254 = ~n11252 & n11253 ;
  assign n11255 = n11251 & n11254 ;
  assign n11256 = \ctl_rf_c2_rf_chllp_cnt_reg[2]/NET0131  & n11255 ;
  assign n11257 = \ctl_rf_be_d1_reg[0]/P0001  & ~\ctl_rf_c2_rf_ch_en_reg/NET0131  ;
  assign n11258 = ~n3772 & n11257 ;
  assign n11259 = ~n4139 & n11258 ;
  assign n11260 = ~\ctl_rf_c2_rf_chllp_cnt_reg[2]/NET0131  & ~n11255 ;
  assign n11261 = ~n11259 & ~n11260 ;
  assign n11262 = ~n11256 & n11261 ;
  assign n11263 = ~\ctl_rf_c2_rf_chllp_cnt_reg[3]/NET0131  & ~n11256 ;
  assign n11264 = \ctl_rf_c2_rf_chllp_cnt_reg[2]/NET0131  & \ctl_rf_c2_rf_chllp_cnt_reg[3]/NET0131  ;
  assign n11265 = n11255 & n11264 ;
  assign n11266 = ~n11259 & ~n11265 ;
  assign n11267 = ~n11263 & n11266 ;
  assign n11268 = \ctl_rf_c3_rf_chllp_on_reg/NET0131  & \de_de_st_reg[5]/NET0131  ;
  assign n11269 = ~n2983 & n11268 ;
  assign n11270 = n3024 & n11269 ;
  assign n11271 = ~\ctl_rf_c3_rf_chabt_reg/NET0131  & ~n2814 ;
  assign n11272 = \ctl_rf_c3_rf_chllp_cnt_reg[0]/NET0131  & \ctl_rf_c3_rf_chllp_cnt_reg[1]/NET0131  ;
  assign n11273 = ~n11271 & n11272 ;
  assign n11274 = n11270 & n11273 ;
  assign n11275 = \ctl_rf_c3_rf_chllp_cnt_reg[2]/NET0131  & n11274 ;
  assign n11276 = \ctl_rf_be_d1_reg[0]/P0001  & ~\ctl_rf_c3_rf_ch_en_reg/NET0131  ;
  assign n11277 = ~n3772 & n11276 ;
  assign n11278 = ~n4156 & n11277 ;
  assign n11279 = ~\ctl_rf_c3_rf_chllp_cnt_reg[2]/NET0131  & ~n11274 ;
  assign n11280 = ~n11278 & ~n11279 ;
  assign n11281 = ~n11275 & n11280 ;
  assign n11282 = ~\ctl_rf_c3_rf_chllp_cnt_reg[3]/NET0131  & ~n11275 ;
  assign n11283 = \ctl_rf_c3_rf_chllp_cnt_reg[2]/NET0131  & \ctl_rf_c3_rf_chllp_cnt_reg[3]/NET0131  ;
  assign n11284 = n11274 & n11283 ;
  assign n11285 = ~n11278 & ~n11284 ;
  assign n11286 = ~n11282 & n11285 ;
  assign n11287 = \ctl_rf_c4_rf_chllp_on_reg/NET0131  & \de_de_st_reg[5]/NET0131  ;
  assign n11288 = n2983 & n11287 ;
  assign n11289 = n2999 & n11288 ;
  assign n11290 = ~\ctl_rf_c4_rf_chabt_reg/NET0131  & ~n2814 ;
  assign n11291 = \ctl_rf_c4_rf_chllp_cnt_reg[0]/NET0131  & \ctl_rf_c4_rf_chllp_cnt_reg[1]/NET0131  ;
  assign n11292 = ~n11290 & n11291 ;
  assign n11293 = n11289 & n11292 ;
  assign n11294 = \ctl_rf_c4_rf_chllp_cnt_reg[2]/NET0131  & n11293 ;
  assign n11295 = \ctl_rf_be_d1_reg[0]/P0001  & ~\ctl_rf_c4_rf_ch_en_reg/NET0131  ;
  assign n11296 = ~n3772 & n11295 ;
  assign n11297 = ~n3766 & n11296 ;
  assign n11298 = ~\ctl_rf_c4_rf_chllp_cnt_reg[2]/NET0131  & ~n11293 ;
  assign n11299 = ~n11297 & ~n11298 ;
  assign n11300 = ~n11294 & n11299 ;
  assign n11301 = ~\ctl_rf_c4_rf_chllp_cnt_reg[3]/NET0131  & ~n11294 ;
  assign n11302 = \ctl_rf_c4_rf_chllp_cnt_reg[2]/NET0131  & \ctl_rf_c4_rf_chllp_cnt_reg[3]/NET0131  ;
  assign n11303 = n11293 & n11302 ;
  assign n11304 = ~n11297 & ~n11303 ;
  assign n11305 = ~n11301 & n11304 ;
  assign n11306 = \ctl_rf_c5_rf_chllp_on_reg/NET0131  & \de_de_st_reg[5]/NET0131  ;
  assign n11307 = ~n2983 & n11306 ;
  assign n11308 = n2999 & n11307 ;
  assign n11309 = ~\ctl_rf_c5_rf_chabt_reg/NET0131  & ~n2814 ;
  assign n11310 = \ctl_rf_c5_rf_chllp_cnt_reg[0]/NET0131  & \ctl_rf_c5_rf_chllp_cnt_reg[1]/NET0131  ;
  assign n11311 = ~n11309 & n11310 ;
  assign n11312 = n11308 & n11311 ;
  assign n11313 = \ctl_rf_c5_rf_chllp_cnt_reg[2]/NET0131  & n11312 ;
  assign n11314 = \ctl_rf_be_d1_reg[0]/P0001  & ~\ctl_rf_c5_rf_ch_en_reg/NET0131  ;
  assign n11315 = ~n3772 & n11314 ;
  assign n11316 = ~n4070 & n11315 ;
  assign n11317 = ~\ctl_rf_c5_rf_chllp_cnt_reg[2]/NET0131  & ~n11312 ;
  assign n11318 = ~n11316 & ~n11317 ;
  assign n11319 = ~n11313 & n11318 ;
  assign n11320 = ~\ctl_rf_c5_rf_chllp_cnt_reg[3]/NET0131  & ~n11313 ;
  assign n11321 = \ctl_rf_c5_rf_chllp_cnt_reg[2]/NET0131  & \ctl_rf_c5_rf_chllp_cnt_reg[3]/NET0131  ;
  assign n11322 = n11312 & n11321 ;
  assign n11323 = ~n11316 & ~n11322 ;
  assign n11324 = ~n11320 & n11323 ;
  assign n11325 = \ctl_rf_c6_rf_chllp_on_reg/NET0131  & \de_de_st_reg[5]/NET0131  ;
  assign n11326 = n2983 & n11325 ;
  assign n11327 = n3011 & n11326 ;
  assign n11328 = ~\ctl_rf_c6_rf_chabt_reg/NET0131  & ~n2814 ;
  assign n11329 = \ctl_rf_c6_rf_chllp_cnt_reg[0]/NET0131  & \ctl_rf_c6_rf_chllp_cnt_reg[1]/NET0131  ;
  assign n11330 = ~n11328 & n11329 ;
  assign n11331 = n11327 & n11330 ;
  assign n11332 = \ctl_rf_c6_rf_chllp_cnt_reg[2]/NET0131  & n11331 ;
  assign n11333 = \ctl_rf_be_d1_reg[0]/P0001  & ~\ctl_rf_c6_rf_ch_en_reg/NET0131  ;
  assign n11334 = ~n3772 & n11333 ;
  assign n11335 = ~n4088 & n11334 ;
  assign n11336 = ~\ctl_rf_c6_rf_chllp_cnt_reg[2]/NET0131  & ~n11331 ;
  assign n11337 = ~n11335 & ~n11336 ;
  assign n11338 = ~n11332 & n11337 ;
  assign n11339 = ~\ctl_rf_c6_rf_chllp_cnt_reg[3]/NET0131  & ~n11332 ;
  assign n11340 = \ctl_rf_c6_rf_chllp_cnt_reg[2]/NET0131  & \ctl_rf_c6_rf_chllp_cnt_reg[3]/NET0131  ;
  assign n11341 = n11331 & n11340 ;
  assign n11342 = ~n11335 & ~n11341 ;
  assign n11343 = ~n11339 & n11342 ;
  assign n11344 = \ctl_rf_c7_rf_chllp_on_reg/NET0131  & \de_de_st_reg[5]/NET0131  ;
  assign n11345 = ~n2983 & n11344 ;
  assign n11346 = n3011 & n11345 ;
  assign n11347 = ~\ctl_rf_c7_rf_chabt_reg/NET0131  & ~n2814 ;
  assign n11348 = \ctl_rf_c7_rf_chllp_cnt_reg[0]/NET0131  & \ctl_rf_c7_rf_chllp_cnt_reg[1]/NET0131  ;
  assign n11349 = ~n11347 & n11348 ;
  assign n11350 = n11346 & n11349 ;
  assign n11351 = \ctl_rf_c7_rf_chllp_cnt_reg[2]/NET0131  & n11350 ;
  assign n11352 = \ctl_rf_be_d1_reg[0]/P0001  & ~\ctl_rf_c7_rf_ch_en_reg/NET0131  ;
  assign n11353 = ~n3772 & n11352 ;
  assign n11354 = ~n4105 & n11353 ;
  assign n11355 = ~\ctl_rf_c7_rf_chllp_cnt_reg[2]/NET0131  & ~n11350 ;
  assign n11356 = ~n11354 & ~n11355 ;
  assign n11357 = ~n11351 & n11356 ;
  assign n11358 = ~\ctl_rf_c7_rf_chllp_cnt_reg[3]/NET0131  & ~n11351 ;
  assign n11359 = \ctl_rf_c7_rf_chllp_cnt_reg[2]/NET0131  & \ctl_rf_c7_rf_chllp_cnt_reg[3]/NET0131  ;
  assign n11360 = n11350 & n11359 ;
  assign n11361 = ~n11354 & ~n11360 ;
  assign n11362 = ~n11358 & n11361 ;
  assign n11363 = \ahb_slv_br_st_reg[2]/NET0131  & ~n2848 ;
  assign n11364 = ~n2880 & n11363 ;
  assign n11365 = \hresp_br[0]_pad  & n11029 ;
  assign n11366 = ~n11364 & ~n11365 ;
  assign n11367 = ~n11036 & ~n11366 ;
  assign n11368 = \ctl_rf_c0_rf_chllp_cnt_reg[0]/NET0131  & ~n11214 ;
  assign n11369 = n11213 & n11368 ;
  assign n11370 = n11213 & ~n11214 ;
  assign n11371 = ~\ctl_rf_c0_rf_chllp_cnt_reg[0]/NET0131  & ~n11370 ;
  assign n11372 = ~n11369 & ~n11371 ;
  assign n11373 = ~n11221 & n11372 ;
  assign n11374 = \ctl_rf_c1_rf_chllp_cnt_reg[0]/NET0131  & ~n11233 ;
  assign n11375 = n11232 & n11374 ;
  assign n11376 = n11232 & ~n11233 ;
  assign n11377 = ~\ctl_rf_c1_rf_chllp_cnt_reg[0]/NET0131  & ~n11376 ;
  assign n11378 = ~n11375 & ~n11377 ;
  assign n11379 = ~n11240 & n11378 ;
  assign n11380 = \ctl_rf_c5_rf_chllp_cnt_reg[0]/NET0131  & ~n11309 ;
  assign n11381 = n11308 & n11380 ;
  assign n11382 = n11308 & ~n11309 ;
  assign n11383 = ~\ctl_rf_c5_rf_chllp_cnt_reg[0]/NET0131  & ~n11382 ;
  assign n11384 = ~n11381 & ~n11383 ;
  assign n11385 = ~n11316 & n11384 ;
  assign n11386 = \ctl_rf_c2_rf_chllp_cnt_reg[0]/NET0131  & ~n11252 ;
  assign n11387 = n11251 & n11386 ;
  assign n11388 = n11251 & ~n11252 ;
  assign n11389 = ~\ctl_rf_c2_rf_chllp_cnt_reg[0]/NET0131  & ~n11388 ;
  assign n11390 = ~n11387 & ~n11389 ;
  assign n11391 = ~n11259 & n11390 ;
  assign n11392 = \ctl_rf_c3_rf_chllp_cnt_reg[0]/NET0131  & ~n11271 ;
  assign n11393 = n11270 & n11392 ;
  assign n11394 = n11270 & ~n11271 ;
  assign n11395 = ~\ctl_rf_c3_rf_chllp_cnt_reg[0]/NET0131  & ~n11394 ;
  assign n11396 = ~n11393 & ~n11395 ;
  assign n11397 = ~n11278 & n11396 ;
  assign n11398 = \ctl_rf_c4_rf_chllp_cnt_reg[0]/NET0131  & ~n11290 ;
  assign n11399 = n11289 & n11398 ;
  assign n11400 = n11289 & ~n11290 ;
  assign n11401 = ~\ctl_rf_c4_rf_chllp_cnt_reg[0]/NET0131  & ~n11400 ;
  assign n11402 = ~n11399 & ~n11401 ;
  assign n11403 = ~n11297 & n11402 ;
  assign n11404 = \ctl_rf_c6_rf_chllp_cnt_reg[0]/NET0131  & ~n11328 ;
  assign n11405 = n11327 & n11404 ;
  assign n11406 = n11327 & ~n11328 ;
  assign n11407 = ~\ctl_rf_c6_rf_chllp_cnt_reg[0]/NET0131  & ~n11406 ;
  assign n11408 = ~n11405 & ~n11407 ;
  assign n11409 = ~n11335 & n11408 ;
  assign n11410 = \ctl_rf_c7_rf_chllp_cnt_reg[0]/NET0131  & ~n11347 ;
  assign n11411 = n11346 & n11410 ;
  assign n11412 = n11346 & ~n11347 ;
  assign n11413 = ~\ctl_rf_c7_rf_chllp_cnt_reg[0]/NET0131  & ~n11412 ;
  assign n11414 = ~n11411 & ~n11413 ;
  assign n11415 = ~n11354 & n11414 ;
  assign n11416 = ~\ctl_rf_c0_rf_chllp_cnt_reg[1]/NET0131  & ~n11369 ;
  assign n11417 = ~n11217 & ~n11416 ;
  assign n11418 = ~n11221 & n11417 ;
  assign n11419 = ~\ctl_rf_c1_rf_chllp_cnt_reg[1]/NET0131  & ~n11375 ;
  assign n11420 = ~n11236 & ~n11419 ;
  assign n11421 = ~n11240 & n11420 ;
  assign n11422 = ~\ctl_rf_c2_rf_chllp_cnt_reg[1]/NET0131  & ~n11387 ;
  assign n11423 = ~n11255 & ~n11422 ;
  assign n11424 = ~n11259 & n11423 ;
  assign n11425 = ~\ctl_rf_c3_rf_chllp_cnt_reg[1]/NET0131  & ~n11393 ;
  assign n11426 = ~n11274 & ~n11425 ;
  assign n11427 = ~n11278 & n11426 ;
  assign n11428 = ~\ctl_rf_c4_rf_chllp_cnt_reg[1]/NET0131  & ~n11399 ;
  assign n11429 = ~n11293 & ~n11428 ;
  assign n11430 = ~n11297 & n11429 ;
  assign n11431 = ~\ctl_rf_c5_rf_chllp_cnt_reg[1]/NET0131  & ~n11381 ;
  assign n11432 = ~n11312 & ~n11431 ;
  assign n11433 = ~n11316 & n11432 ;
  assign n11434 = ~\ctl_rf_c6_rf_chllp_cnt_reg[1]/NET0131  & ~n11405 ;
  assign n11435 = ~n11331 & ~n11434 ;
  assign n11436 = ~n11335 & n11435 ;
  assign n11437 = ~\ctl_rf_c7_rf_chllp_cnt_reg[1]/NET0131  & ~n11411 ;
  assign n11438 = ~n11350 & ~n11437 ;
  assign n11439 = ~n11354 & n11438 ;
  assign n11440 = \ahb_slv_br_st_reg[2]/NET0131  & ~\m1_mux_hrmxnof_reg/NET0131  ;
  assign n11441 = ~n2912 & n11440 ;
  assign n11442 = \hresp_br[1]_pad  & n11029 ;
  assign n11443 = ~n11036 & ~n11442 ;
  assign n11444 = ~n11441 & n11443 ;
  assign n11445 = n9528 & ~n9545 ;
  assign n11446 = ~\ahb_slv_slv_ad_d1o_reg[8]/NET0131  & \ahb_slv_slv_wr_d1o_reg/NET0131  ;
  assign n11447 = n2228 & n11446 ;
  assign n11448 = ~\ahb_slv_slv_ad_d1o_reg[2]/NET0131  & n2275 ;
  assign n11449 = \ctl_rf_be_d1_reg[2]/P0001  & n8577 ;
  assign n11450 = n11448 & n11449 ;
  assign n11451 = n11447 & n11450 ;
  assign n11452 = \ctl_rf_abt_reg[0]/NET0131  & ~n11451 ;
  assign n11453 = \ctl_rf_abt_reg[0]/NET0131  & ~n2680 ;
  assign n11454 = ~n2679 & n11453 ;
  assign n11455 = ~n11452 & ~n11454 ;
  assign n11456 = ~n5176 & n11455 ;
  assign n11457 = \ctl_rf_abt_reg[2]/NET0131  & ~n11451 ;
  assign n11458 = \ctl_rf_abt_reg[2]/NET0131  & ~n2400 ;
  assign n11459 = ~n2399 & n11458 ;
  assign n11460 = ~n11457 & ~n11459 ;
  assign n11461 = ~n5197 & n11460 ;
  assign n11462 = \ctl_rf_abt_reg[1]/NET0131  & ~n11451 ;
  assign n11463 = \ctl_rf_abt_reg[1]/NET0131  & ~n2260 ;
  assign n11464 = ~n2259 & n11463 ;
  assign n11465 = ~n11462 & ~n11464 ;
  assign n11466 = ~n5187 & n11465 ;
  assign n11467 = \ctl_rf_abt_reg[3]/NET0131  & ~n11451 ;
  assign n11468 = \ctl_rf_abt_reg[3]/NET0131  & ~n2409 ;
  assign n11469 = ~n2408 & n11468 ;
  assign n11470 = ~n11467 & ~n11469 ;
  assign n11471 = ~n5207 & n11470 ;
  assign n11472 = \ctl_rf_abt_reg[4]/NET0131  & ~n11451 ;
  assign n11473 = \ctl_rf_abt_reg[4]/NET0131  & ~n2566 ;
  assign n11474 = ~n2565 & n11473 ;
  assign n11475 = ~n11472 & ~n11474 ;
  assign n11476 = ~n5217 & n11475 ;
  assign n11477 = \ctl_rf_abt_reg[5]/NET0131  & ~n11451 ;
  assign n11478 = \ctl_rf_abt_reg[5]/NET0131  & ~n2366 ;
  assign n11479 = ~n2365 & n11478 ;
  assign n11480 = ~n11477 & ~n11479 ;
  assign n11481 = ~n5227 & n11480 ;
  assign n11482 = \ctl_rf_abt_reg[6]/NET0131  & ~n11451 ;
  assign n11483 = \ctl_rf_abt_reg[6]/NET0131  & ~n2500 ;
  assign n11484 = ~n2499 & n11483 ;
  assign n11485 = ~n11482 & ~n11484 ;
  assign n11486 = ~n5237 & n11485 ;
  assign n11487 = \ctl_rf_abt_reg[7]/NET0131  & ~n11451 ;
  assign n11488 = \ctl_rf_abt_reg[7]/NET0131  & ~n2529 ;
  assign n11489 = ~n2528 & n11488 ;
  assign n11490 = ~n11487 & ~n11489 ;
  assign n11491 = ~n5247 & n11490 ;
  assign n11492 = \h1prot[0]_pad  & n2830 ;
  assign n11493 = \h1prot[0]_pad  & n2764 ;
  assign n11494 = n2798 & n11493 ;
  assign n11495 = ~n11492 & ~n11494 ;
  assign n11496 = \ahb_slv_slv_pt_d1o_reg[0]/NET0131  & \de_m1_arb_st_reg[1]/NET0131  ;
  assign n11497 = ~n2830 & n11496 ;
  assign n11498 = ~n2799 & n11497 ;
  assign n11499 = n11495 & ~n11498 ;
  assign n11500 = ~n2830 & ~n2846 ;
  assign n11501 = ~n2799 & n11500 ;
  assign n11502 = ~n2799 & n4518 ;
  assign n11503 = \ahb_mst1_mx_dtp_reg/NET0131  & n2830 ;
  assign n11504 = \ahb_mst1_mx_dtp_reg/NET0131  & n2764 ;
  assign n11505 = n2798 & n11504 ;
  assign n11506 = ~n11503 & ~n11505 ;
  assign n11507 = ~n11502 & n11506 ;
  assign n11508 = ~\ahb_slv_slv_ad_d1o_reg[2]/NET0131  & \ctl_rf_be_d1_reg[0]/P0001  ;
  assign n11509 = n2276 & n11508 ;
  assign n11510 = n11447 & n11509 ;
  assign n11511 = \ctl_rf_tc_reg[7]/NET0131  & ~n11510 ;
  assign n11512 = \ctl_rf_tc_reg[7]/NET0131  & ~n2247 ;
  assign n11513 = ~n2246 & n11512 ;
  assign n11514 = ~n11511 & ~n11513 ;
  assign n11515 = \de_de_st_reg[5]/NET0131  & n2814 ;
  assign n11516 = ~\ctl_rf_c7_rf_int_tc_msk_reg/NET0131  & ~n2983 ;
  assign n11517 = n3011 & n11516 ;
  assign n11518 = n11515 & n11517 ;
  assign n11519 = n11514 & ~n11518 ;
  assign n11520 = \ctl_rf_tc_reg[3]/NET0131  & ~n11510 ;
  assign n11521 = \ctl_rf_tc_reg[3]/NET0131  & ~n9044 ;
  assign n11522 = ~n9043 & n11521 ;
  assign n11523 = ~n11520 & ~n11522 ;
  assign n11524 = ~\ctl_rf_c3_rf_int_tc_msk_reg/NET0131  & ~n2983 ;
  assign n11525 = n3024 & n11524 ;
  assign n11526 = n11515 & n11525 ;
  assign n11527 = n11523 & ~n11526 ;
  assign n11528 = \ctl_rf_tc_reg[0]/NET0131  & ~n11510 ;
  assign n11529 = \ctl_rf_tc_reg[0]/NET0131  & ~n3771 ;
  assign n11530 = ~n3770 & n11529 ;
  assign n11531 = ~n11528 & ~n11530 ;
  assign n11532 = ~\ctl_rf_c0_rf_int_tc_msk_reg/NET0131  & n2983 ;
  assign n11533 = n3050 & n11532 ;
  assign n11534 = n11515 & n11533 ;
  assign n11535 = n11531 & ~n11534 ;
  assign n11536 = \ctl_rf_tc_reg[1]/NET0131  & ~n11510 ;
  assign n11537 = \ctl_rf_tc_reg[1]/NET0131  & ~n8992 ;
  assign n11538 = ~n8991 & n11537 ;
  assign n11539 = ~n11536 & ~n11538 ;
  assign n11540 = ~\ctl_rf_c1_rf_int_tc_msk_reg/NET0131  & ~n2983 ;
  assign n11541 = n3050 & n11540 ;
  assign n11542 = n11515 & n11541 ;
  assign n11543 = n11539 & ~n11542 ;
  assign n11544 = \ctl_rf_tc_reg[4]/NET0131  & ~n11510 ;
  assign n11545 = \ctl_rf_tc_reg[4]/NET0131  & ~n8714 ;
  assign n11546 = ~n8713 & n11545 ;
  assign n11547 = ~n11544 & ~n11546 ;
  assign n11548 = ~\ctl_rf_c4_rf_int_tc_msk_reg/NET0131  & n2983 ;
  assign n11549 = n2999 & n11548 ;
  assign n11550 = n11515 & n11549 ;
  assign n11551 = n11547 & ~n11550 ;
  assign n11552 = \ctl_rf_tc_reg[2]/NET0131  & ~n11510 ;
  assign n11553 = \ctl_rf_tc_reg[2]/NET0131  & ~n9001 ;
  assign n11554 = ~n9000 & n11553 ;
  assign n11555 = ~n11552 & ~n11554 ;
  assign n11556 = ~\ctl_rf_c2_rf_int_tc_msk_reg/NET0131  & n2983 ;
  assign n11557 = n3024 & n11556 ;
  assign n11558 = n11515 & n11557 ;
  assign n11559 = n11555 & ~n11558 ;
  assign n11560 = \ctl_rf_tc_reg[6]/NET0131  & ~n11510 ;
  assign n11561 = \ctl_rf_tc_reg[6]/NET0131  & ~n8596 ;
  assign n11562 = ~n8595 & n11561 ;
  assign n11563 = ~n11560 & ~n11562 ;
  assign n11564 = ~\ctl_rf_c6_rf_int_tc_msk_reg/NET0131  & n2983 ;
  assign n11565 = n3011 & n11564 ;
  assign n11566 = n11515 & n11565 ;
  assign n11567 = n11563 & ~n11566 ;
  assign n11568 = \ctl_rf_tc_reg[5]/NET0131  & ~n11510 ;
  assign n11569 = \ctl_rf_tc_reg[5]/NET0131  & ~n8587 ;
  assign n11570 = ~n8586 & n11569 ;
  assign n11571 = ~n11568 & ~n11570 ;
  assign n11572 = ~\ctl_rf_c5_rf_int_tc_msk_reg/NET0131  & ~n2983 ;
  assign n11573 = n2999 & n11572 ;
  assign n11574 = n11515 & n11573 ;
  assign n11575 = n11571 & ~n11574 ;
  assign n11576 = \ctl_rf_c2_rf_dwidth_reg[2]/NET0131  & n2983 ;
  assign n11577 = n3024 & n11576 ;
  assign n11578 = \ctl_rf_c1_rf_dwidth_reg[2]/NET0131  & ~n2983 ;
  assign n11579 = n3050 & n11578 ;
  assign n11580 = ~n11577 & ~n11579 ;
  assign n11581 = \ctl_rf_c7_rf_dwidth_reg[2]/NET0131  & ~n2983 ;
  assign n11582 = n3011 & n11581 ;
  assign n11583 = \ctl_rf_c0_rf_dwidth_reg[2]/NET0131  & n2983 ;
  assign n11584 = n3050 & n11583 ;
  assign n11585 = ~n11582 & ~n11584 ;
  assign n11586 = n11580 & n11585 ;
  assign n11587 = \ctl_rf_c3_rf_dwidth_reg[2]/NET0131  & ~n2983 ;
  assign n11588 = n3024 & n11587 ;
  assign n11589 = \ctl_rf_c6_rf_dwidth_reg[2]/NET0131  & n2983 ;
  assign n11590 = n3011 & n11589 ;
  assign n11591 = ~n11588 & ~n11590 ;
  assign n11592 = \ctl_rf_c5_rf_dwidth_reg[2]/NET0131  & ~n2983 ;
  assign n11593 = n2999 & n11592 ;
  assign n11594 = \ctl_rf_c4_rf_dwidth_reg[2]/NET0131  & n2983 ;
  assign n11595 = n2999 & n11594 ;
  assign n11596 = ~n11593 & ~n11595 ;
  assign n11597 = n11591 & n11596 ;
  assign n11598 = n11586 & n11597 ;
  assign n11599 = \ctl_rf_c2_rf_dst_sel_reg/NET0131  & n2983 ;
  assign n11600 = n3024 & n11599 ;
  assign n11601 = \ctl_rf_c1_rf_dst_sel_reg/NET0131  & ~n2983 ;
  assign n11602 = n3050 & n11601 ;
  assign n11603 = ~n11600 & ~n11602 ;
  assign n11604 = \ctl_rf_c7_rf_dst_sel_reg/NET0131  & ~n2983 ;
  assign n11605 = n3011 & n11604 ;
  assign n11606 = \ctl_rf_c0_rf_dst_sel_reg/NET0131  & n2983 ;
  assign n11607 = n3050 & n11606 ;
  assign n11608 = ~n11605 & ~n11607 ;
  assign n11609 = n11603 & n11608 ;
  assign n11610 = \ctl_rf_c3_rf_dst_sel_reg/NET0131  & ~n2983 ;
  assign n11611 = n3024 & n11610 ;
  assign n11612 = \ctl_rf_c6_rf_dst_sel_reg/NET0131  & n2983 ;
  assign n11613 = n3011 & n11612 ;
  assign n11614 = ~n11611 & ~n11613 ;
  assign n11615 = \ctl_rf_c5_rf_dst_sel_reg/NET0131  & ~n2983 ;
  assign n11616 = n2999 & n11615 ;
  assign n11617 = \ctl_rf_c4_rf_dst_sel_reg/NET0131  & n2983 ;
  assign n11618 = n2999 & n11617 ;
  assign n11619 = ~n11616 & ~n11618 ;
  assign n11620 = n11614 & n11619 ;
  assign n11621 = n11609 & n11620 ;
  assign n11622 = \ctl_rf_c2_rf_swidth_reg[0]/NET0131  & n2983 ;
  assign n11623 = n3024 & n11622 ;
  assign n11624 = \ctl_rf_c1_rf_swidth_reg[0]/NET0131  & ~n2983 ;
  assign n11625 = n3050 & n11624 ;
  assign n11626 = ~n11623 & ~n11625 ;
  assign n11627 = \ctl_rf_c7_rf_swidth_reg[0]/NET0131  & ~n2983 ;
  assign n11628 = n3011 & n11627 ;
  assign n11629 = \ctl_rf_c0_rf_swidth_reg[0]/NET0131  & n2983 ;
  assign n11630 = n3050 & n11629 ;
  assign n11631 = ~n11628 & ~n11630 ;
  assign n11632 = n11626 & n11631 ;
  assign n11633 = \ctl_rf_c3_rf_swidth_reg[0]/NET0131  & ~n2983 ;
  assign n11634 = n3024 & n11633 ;
  assign n11635 = \ctl_rf_c6_rf_swidth_reg[0]/NET0131  & n2983 ;
  assign n11636 = n3011 & n11635 ;
  assign n11637 = ~n11634 & ~n11636 ;
  assign n11638 = \ctl_rf_c5_rf_swidth_reg[0]/NET0131  & ~n2983 ;
  assign n11639 = n2999 & n11638 ;
  assign n11640 = \ctl_rf_c4_rf_swidth_reg[0]/NET0131  & n2983 ;
  assign n11641 = n2999 & n11640 ;
  assign n11642 = ~n11639 & ~n11641 ;
  assign n11643 = n11637 & n11642 ;
  assign n11644 = n11632 & n11643 ;
  assign n11645 = \ctl_rf_c2_rf_dwidth_reg[1]/NET0131  & n2983 ;
  assign n11646 = n3024 & n11645 ;
  assign n11647 = \ctl_rf_c1_rf_dwidth_reg[1]/NET0131  & ~n2983 ;
  assign n11648 = n3050 & n11647 ;
  assign n11649 = ~n11646 & ~n11648 ;
  assign n11650 = \ctl_rf_c7_rf_dwidth_reg[1]/NET0131  & ~n2983 ;
  assign n11651 = n3011 & n11650 ;
  assign n11652 = \ctl_rf_c0_rf_dwidth_reg[1]/NET0131  & n2983 ;
  assign n11653 = n3050 & n11652 ;
  assign n11654 = ~n11651 & ~n11653 ;
  assign n11655 = n11649 & n11654 ;
  assign n11656 = \ctl_rf_c3_rf_dwidth_reg[1]/NET0131  & ~n2983 ;
  assign n11657 = n3024 & n11656 ;
  assign n11658 = \ctl_rf_c6_rf_dwidth_reg[1]/NET0131  & n2983 ;
  assign n11659 = n3011 & n11658 ;
  assign n11660 = ~n11657 & ~n11659 ;
  assign n11661 = \ctl_rf_c5_rf_dwidth_reg[1]/NET0131  & ~n2983 ;
  assign n11662 = n2999 & n11661 ;
  assign n11663 = \ctl_rf_c4_rf_dwidth_reg[1]/NET0131  & n2983 ;
  assign n11664 = n2999 & n11663 ;
  assign n11665 = ~n11662 & ~n11664 ;
  assign n11666 = n11660 & n11665 ;
  assign n11667 = n11655 & n11666 ;
  assign n11668 = \ctl_rf_c2_rf_prot1_reg/NET0131  & n2983 ;
  assign n11669 = n3024 & n11668 ;
  assign n11670 = \ctl_rf_c1_rf_prot1_reg/NET0131  & ~n2983 ;
  assign n11671 = n3050 & n11670 ;
  assign n11672 = ~n11669 & ~n11671 ;
  assign n11673 = \ctl_rf_c7_rf_prot1_reg/NET0131  & ~n2983 ;
  assign n11674 = n3011 & n11673 ;
  assign n11675 = \ctl_rf_c0_rf_prot1_reg/NET0131  & n2983 ;
  assign n11676 = n3050 & n11675 ;
  assign n11677 = ~n11674 & ~n11676 ;
  assign n11678 = n11672 & n11677 ;
  assign n11679 = \ctl_rf_c3_rf_prot1_reg/NET0131  & ~n2983 ;
  assign n11680 = n3024 & n11679 ;
  assign n11681 = \ctl_rf_c6_rf_prot1_reg/NET0131  & n2983 ;
  assign n11682 = n3011 & n11681 ;
  assign n11683 = ~n11680 & ~n11682 ;
  assign n11684 = \ctl_rf_c5_rf_prot1_reg/NET0131  & ~n2983 ;
  assign n11685 = n2999 & n11684 ;
  assign n11686 = \ctl_rf_c4_rf_prot1_reg/NET0131  & n2983 ;
  assign n11687 = n2999 & n11686 ;
  assign n11688 = ~n11685 & ~n11687 ;
  assign n11689 = n11683 & n11688 ;
  assign n11690 = n11678 & n11689 ;
  assign n11691 = \ctl_rf_c2_rf_sad_ctl1_reg/NET0131  & n2983 ;
  assign n11692 = n3024 & n11691 ;
  assign n11693 = \ctl_rf_c1_rf_sad_ctl1_reg/NET0131  & ~n2983 ;
  assign n11694 = n3050 & n11693 ;
  assign n11695 = ~n11692 & ~n11694 ;
  assign n11696 = \ctl_rf_c7_rf_sad_ctl1_reg/NET0131  & ~n2983 ;
  assign n11697 = n3011 & n11696 ;
  assign n11698 = \ctl_rf_c0_rf_sad_ctl1_reg/NET0131  & n2983 ;
  assign n11699 = n3050 & n11698 ;
  assign n11700 = ~n11697 & ~n11699 ;
  assign n11701 = n11695 & n11700 ;
  assign n11702 = \ctl_rf_c3_rf_sad_ctl1_reg/NET0131  & ~n2983 ;
  assign n11703 = n3024 & n11702 ;
  assign n11704 = \ctl_rf_c6_rf_sad_ctl1_reg/NET0131  & n2983 ;
  assign n11705 = n3011 & n11704 ;
  assign n11706 = ~n11703 & ~n11705 ;
  assign n11707 = \ctl_rf_c5_rf_sad_ctl1_reg/NET0131  & ~n2983 ;
  assign n11708 = n2999 & n11707 ;
  assign n11709 = \ctl_rf_c4_rf_sad_ctl1_reg/NET0131  & n2983 ;
  assign n11710 = n2999 & n11709 ;
  assign n11711 = ~n11708 & ~n11710 ;
  assign n11712 = n11706 & n11711 ;
  assign n11713 = n11701 & n11712 ;
  assign n11714 = \ctl_rf_c2_rf_swidth_reg[1]/NET0131  & n2983 ;
  assign n11715 = n3024 & n11714 ;
  assign n11716 = \ctl_rf_c1_rf_swidth_reg[1]/NET0131  & ~n2983 ;
  assign n11717 = n3050 & n11716 ;
  assign n11718 = ~n11715 & ~n11717 ;
  assign n11719 = \ctl_rf_c7_rf_swidth_reg[1]/NET0131  & ~n2983 ;
  assign n11720 = n3011 & n11719 ;
  assign n11721 = \ctl_rf_c0_rf_swidth_reg[1]/NET0131  & n2983 ;
  assign n11722 = n3050 & n11721 ;
  assign n11723 = ~n11720 & ~n11722 ;
  assign n11724 = n11718 & n11723 ;
  assign n11725 = \ctl_rf_c3_rf_swidth_reg[1]/NET0131  & ~n2983 ;
  assign n11726 = n3024 & n11725 ;
  assign n11727 = \ctl_rf_c6_rf_swidth_reg[1]/NET0131  & n2983 ;
  assign n11728 = n3011 & n11727 ;
  assign n11729 = ~n11726 & ~n11728 ;
  assign n11730 = \ctl_rf_c5_rf_swidth_reg[1]/NET0131  & ~n2983 ;
  assign n11731 = n2999 & n11730 ;
  assign n11732 = \ctl_rf_c4_rf_swidth_reg[1]/NET0131  & n2983 ;
  assign n11733 = n2999 & n11732 ;
  assign n11734 = ~n11731 & ~n11733 ;
  assign n11735 = n11729 & n11734 ;
  assign n11736 = n11724 & n11735 ;
  assign n11737 = \ctl_rf_c2_rf_swidth_reg[2]/NET0131  & n2983 ;
  assign n11738 = n3024 & n11737 ;
  assign n11739 = \ctl_rf_c1_rf_swidth_reg[2]/NET0131  & ~n2983 ;
  assign n11740 = n3050 & n11739 ;
  assign n11741 = ~n11738 & ~n11740 ;
  assign n11742 = \ctl_rf_c7_rf_swidth_reg[2]/NET0131  & ~n2983 ;
  assign n11743 = n3011 & n11742 ;
  assign n11744 = \ctl_rf_c0_rf_swidth_reg[2]/NET0131  & n2983 ;
  assign n11745 = n3050 & n11744 ;
  assign n11746 = ~n11743 & ~n11745 ;
  assign n11747 = n11741 & n11746 ;
  assign n11748 = \ctl_rf_c3_rf_swidth_reg[2]/NET0131  & ~n2983 ;
  assign n11749 = n3024 & n11748 ;
  assign n11750 = \ctl_rf_c6_rf_swidth_reg[2]/NET0131  & n2983 ;
  assign n11751 = n3011 & n11750 ;
  assign n11752 = ~n11749 & ~n11751 ;
  assign n11753 = \ctl_rf_c5_rf_swidth_reg[2]/NET0131  & ~n2983 ;
  assign n11754 = n2999 & n11753 ;
  assign n11755 = \ctl_rf_c4_rf_swidth_reg[2]/NET0131  & n2983 ;
  assign n11756 = n2999 & n11755 ;
  assign n11757 = ~n11754 & ~n11756 ;
  assign n11758 = n11752 & n11757 ;
  assign n11759 = n11747 & n11758 ;
  assign n11760 = \ctl_rf_c2_rf_src_sz_reg[0]/NET0131  & n2983 ;
  assign n11761 = n3024 & n11760 ;
  assign n11762 = \ctl_rf_c1_rf_src_sz_reg[0]/NET0131  & ~n2983 ;
  assign n11763 = n3050 & n11762 ;
  assign n11764 = ~n11761 & ~n11763 ;
  assign n11765 = \ctl_rf_c7_rf_src_sz_reg[0]/NET0131  & ~n2983 ;
  assign n11766 = n3011 & n11765 ;
  assign n11767 = \ctl_rf_c0_rf_src_sz_reg[0]/NET0131  & n2983 ;
  assign n11768 = n3050 & n11767 ;
  assign n11769 = ~n11766 & ~n11768 ;
  assign n11770 = n11764 & n11769 ;
  assign n11771 = \ctl_rf_c3_rf_src_sz_reg[0]/NET0131  & ~n2983 ;
  assign n11772 = n3024 & n11771 ;
  assign n11773 = \ctl_rf_c6_rf_src_sz_reg[0]/NET0131  & n2983 ;
  assign n11774 = n3011 & n11773 ;
  assign n11775 = ~n11772 & ~n11774 ;
  assign n11776 = \ctl_rf_c5_rf_src_sz_reg[0]/NET0131  & ~n2983 ;
  assign n11777 = n2999 & n11776 ;
  assign n11778 = \ctl_rf_c4_rf_src_sz_reg[0]/NET0131  & n2983 ;
  assign n11779 = n2999 & n11778 ;
  assign n11780 = ~n11777 & ~n11779 ;
  assign n11781 = n11775 & n11780 ;
  assign n11782 = n11770 & n11781 ;
  assign n11783 = \ctl_rf_c2_rf_src_sel_reg/NET0131  & n2983 ;
  assign n11784 = n3024 & n11783 ;
  assign n11785 = \ctl_rf_c1_rf_src_sel_reg/NET0131  & ~n2983 ;
  assign n11786 = n3050 & n11785 ;
  assign n11787 = ~n11784 & ~n11786 ;
  assign n11788 = \ctl_rf_c7_rf_src_sel_reg/NET0131  & ~n2983 ;
  assign n11789 = n3011 & n11788 ;
  assign n11790 = \ctl_rf_c0_rf_src_sel_reg/NET0131  & n2983 ;
  assign n11791 = n3050 & n11790 ;
  assign n11792 = ~n11789 & ~n11791 ;
  assign n11793 = n11787 & n11792 ;
  assign n11794 = \ctl_rf_c3_rf_src_sel_reg/NET0131  & ~n2983 ;
  assign n11795 = n3024 & n11794 ;
  assign n11796 = \ctl_rf_c6_rf_src_sel_reg/NET0131  & n2983 ;
  assign n11797 = n3011 & n11796 ;
  assign n11798 = ~n11795 & ~n11797 ;
  assign n11799 = \ctl_rf_c5_rf_src_sel_reg/NET0131  & ~n2983 ;
  assign n11800 = n2999 & n11799 ;
  assign n11801 = \ctl_rf_c4_rf_src_sel_reg/NET0131  & n2983 ;
  assign n11802 = n2999 & n11801 ;
  assign n11803 = ~n11800 & ~n11802 ;
  assign n11804 = n11798 & n11803 ;
  assign n11805 = n11793 & n11804 ;
  assign n11806 = \ctl_rf_c2_rf_dad_ctl0_reg/NET0131  & n2983 ;
  assign n11807 = n3024 & n11806 ;
  assign n11808 = \ctl_rf_c1_rf_dad_ctl0_reg/NET0131  & ~n2983 ;
  assign n11809 = n3050 & n11808 ;
  assign n11810 = ~n11807 & ~n11809 ;
  assign n11811 = \ctl_rf_c7_rf_dad_ctl0_reg/NET0131  & ~n2983 ;
  assign n11812 = n3011 & n11811 ;
  assign n11813 = \ctl_rf_c0_rf_dad_ctl0_reg/NET0131  & n2983 ;
  assign n11814 = n3050 & n11813 ;
  assign n11815 = ~n11812 & ~n11814 ;
  assign n11816 = n11810 & n11815 ;
  assign n11817 = \ctl_rf_c3_rf_dad_ctl0_reg/NET0131  & ~n2983 ;
  assign n11818 = n3024 & n11817 ;
  assign n11819 = \ctl_rf_c6_rf_dad_ctl0_reg/NET0131  & n2983 ;
  assign n11820 = n3011 & n11819 ;
  assign n11821 = ~n11818 & ~n11820 ;
  assign n11822 = \ctl_rf_c5_rf_dad_ctl0_reg/NET0131  & ~n2983 ;
  assign n11823 = n2999 & n11822 ;
  assign n11824 = \ctl_rf_c4_rf_dad_ctl0_reg/NET0131  & n2983 ;
  assign n11825 = n2999 & n11824 ;
  assign n11826 = ~n11823 & ~n11825 ;
  assign n11827 = n11821 & n11826 ;
  assign n11828 = n11816 & n11827 ;
  assign n11829 = \ctl_rf_c2_rf_dad_ctl1_reg/NET0131  & n2983 ;
  assign n11830 = n3024 & n11829 ;
  assign n11831 = \ctl_rf_c1_rf_dad_ctl1_reg/NET0131  & ~n2983 ;
  assign n11832 = n3050 & n11831 ;
  assign n11833 = ~n11830 & ~n11832 ;
  assign n11834 = \ctl_rf_c7_rf_dad_ctl1_reg/NET0131  & ~n2983 ;
  assign n11835 = n3011 & n11834 ;
  assign n11836 = \ctl_rf_c0_rf_dad_ctl1_reg/NET0131  & n2983 ;
  assign n11837 = n3050 & n11836 ;
  assign n11838 = ~n11835 & ~n11837 ;
  assign n11839 = n11833 & n11838 ;
  assign n11840 = \ctl_rf_c3_rf_dad_ctl1_reg/NET0131  & ~n2983 ;
  assign n11841 = n3024 & n11840 ;
  assign n11842 = \ctl_rf_c6_rf_dad_ctl1_reg/NET0131  & n2983 ;
  assign n11843 = n3011 & n11842 ;
  assign n11844 = ~n11841 & ~n11843 ;
  assign n11845 = \ctl_rf_c5_rf_dad_ctl1_reg/NET0131  & ~n2983 ;
  assign n11846 = n2999 & n11845 ;
  assign n11847 = \ctl_rf_c4_rf_dad_ctl1_reg/NET0131  & n2983 ;
  assign n11848 = n2999 & n11847 ;
  assign n11849 = ~n11846 & ~n11848 ;
  assign n11850 = n11844 & n11849 ;
  assign n11851 = n11839 & n11850 ;
  assign n11852 = \ctl_rf_c2_rf_sad_ctl0_reg/NET0131  & n2983 ;
  assign n11853 = n3024 & n11852 ;
  assign n11854 = \ctl_rf_c1_rf_sad_ctl0_reg/NET0131  & ~n2983 ;
  assign n11855 = n3050 & n11854 ;
  assign n11856 = ~n11853 & ~n11855 ;
  assign n11857 = \ctl_rf_c7_rf_sad_ctl0_reg/NET0131  & ~n2983 ;
  assign n11858 = n3011 & n11857 ;
  assign n11859 = \ctl_rf_c0_rf_sad_ctl0_reg/NET0131  & n2983 ;
  assign n11860 = n3050 & n11859 ;
  assign n11861 = ~n11858 & ~n11860 ;
  assign n11862 = n11856 & n11861 ;
  assign n11863 = \ctl_rf_c3_rf_sad_ctl0_reg/NET0131  & ~n2983 ;
  assign n11864 = n3024 & n11863 ;
  assign n11865 = \ctl_rf_c6_rf_sad_ctl0_reg/NET0131  & n2983 ;
  assign n11866 = n3011 & n11865 ;
  assign n11867 = ~n11864 & ~n11866 ;
  assign n11868 = \ctl_rf_c5_rf_sad_ctl0_reg/NET0131  & ~n2983 ;
  assign n11869 = n2999 & n11868 ;
  assign n11870 = \ctl_rf_c4_rf_sad_ctl0_reg/NET0131  & n2983 ;
  assign n11871 = n2999 & n11870 ;
  assign n11872 = ~n11869 & ~n11871 ;
  assign n11873 = n11867 & n11872 ;
  assign n11874 = n11862 & n11873 ;
  assign n11875 = \ctl_rf_c2_rf_dwidth_reg[0]/NET0131  & n2983 ;
  assign n11876 = n3024 & n11875 ;
  assign n11877 = \ctl_rf_c1_rf_dwidth_reg[0]/NET0131  & ~n2983 ;
  assign n11878 = n3050 & n11877 ;
  assign n11879 = ~n11876 & ~n11878 ;
  assign n11880 = \ctl_rf_c7_rf_dwidth_reg[0]/NET0131  & ~n2983 ;
  assign n11881 = n3011 & n11880 ;
  assign n11882 = \ctl_rf_c0_rf_dwidth_reg[0]/NET0131  & n2983 ;
  assign n11883 = n3050 & n11882 ;
  assign n11884 = ~n11881 & ~n11883 ;
  assign n11885 = n11879 & n11884 ;
  assign n11886 = \ctl_rf_c3_rf_dwidth_reg[0]/NET0131  & ~n2983 ;
  assign n11887 = n3024 & n11886 ;
  assign n11888 = \ctl_rf_c6_rf_dwidth_reg[0]/NET0131  & n2983 ;
  assign n11889 = n3011 & n11888 ;
  assign n11890 = ~n11887 & ~n11889 ;
  assign n11891 = \ctl_rf_c5_rf_dwidth_reg[0]/NET0131  & ~n2983 ;
  assign n11892 = n2999 & n11891 ;
  assign n11893 = \ctl_rf_c4_rf_dwidth_reg[0]/NET0131  & n2983 ;
  assign n11894 = n2999 & n11893 ;
  assign n11895 = ~n11892 & ~n11894 ;
  assign n11896 = n11890 & n11895 ;
  assign n11897 = n11885 & n11896 ;
  assign n11898 = \ctl_rf_c2_rf_prot2_reg/NET0131  & n2983 ;
  assign n11899 = n3024 & n11898 ;
  assign n11900 = \ctl_rf_c1_rf_prot2_reg/NET0131  & ~n2983 ;
  assign n11901 = n3050 & n11900 ;
  assign n11902 = ~n11899 & ~n11901 ;
  assign n11903 = \ctl_rf_c7_rf_prot2_reg/NET0131  & ~n2983 ;
  assign n11904 = n3011 & n11903 ;
  assign n11905 = \ctl_rf_c0_rf_prot2_reg/NET0131  & n2983 ;
  assign n11906 = n3050 & n11905 ;
  assign n11907 = ~n11904 & ~n11906 ;
  assign n11908 = n11902 & n11907 ;
  assign n11909 = \ctl_rf_c3_rf_prot2_reg/NET0131  & ~n2983 ;
  assign n11910 = n3024 & n11909 ;
  assign n11911 = \ctl_rf_c6_rf_prot2_reg/NET0131  & n2983 ;
  assign n11912 = n3011 & n11911 ;
  assign n11913 = ~n11910 & ~n11912 ;
  assign n11914 = \ctl_rf_c5_rf_prot2_reg/NET0131  & ~n2983 ;
  assign n11915 = n2999 & n11914 ;
  assign n11916 = \ctl_rf_c4_rf_prot2_reg/NET0131  & n2983 ;
  assign n11917 = n2999 & n11916 ;
  assign n11918 = ~n11915 & ~n11917 ;
  assign n11919 = n11913 & n11918 ;
  assign n11920 = n11908 & n11919 ;
  assign n11921 = \ctl_rf_c2_rf_src_sz_reg[1]/NET0131  & n2983 ;
  assign n11922 = n3024 & n11921 ;
  assign n11923 = \ctl_rf_c1_rf_src_sz_reg[1]/NET0131  & ~n2983 ;
  assign n11924 = n3050 & n11923 ;
  assign n11925 = ~n11922 & ~n11924 ;
  assign n11926 = \ctl_rf_c7_rf_src_sz_reg[1]/NET0131  & ~n2983 ;
  assign n11927 = n3011 & n11926 ;
  assign n11928 = \ctl_rf_c0_rf_src_sz_reg[1]/NET0131  & n2983 ;
  assign n11929 = n3050 & n11928 ;
  assign n11930 = ~n11927 & ~n11929 ;
  assign n11931 = n11925 & n11930 ;
  assign n11932 = \ctl_rf_c3_rf_src_sz_reg[1]/NET0131  & ~n2983 ;
  assign n11933 = n3024 & n11932 ;
  assign n11934 = \ctl_rf_c6_rf_src_sz_reg[1]/NET0131  & n2983 ;
  assign n11935 = n3011 & n11934 ;
  assign n11936 = ~n11933 & ~n11935 ;
  assign n11937 = \ctl_rf_c5_rf_src_sz_reg[1]/NET0131  & ~n2983 ;
  assign n11938 = n2999 & n11937 ;
  assign n11939 = \ctl_rf_c4_rf_src_sz_reg[1]/NET0131  & n2983 ;
  assign n11940 = n2999 & n11939 ;
  assign n11941 = ~n11938 & ~n11940 ;
  assign n11942 = n11936 & n11941 ;
  assign n11943 = n11931 & n11942 ;
  assign n11944 = \ctl_rf_c2_rf_prot3_reg/NET0131  & n2983 ;
  assign n11945 = n3024 & n11944 ;
  assign n11946 = \ctl_rf_c1_rf_prot3_reg/NET0131  & ~n2983 ;
  assign n11947 = n3050 & n11946 ;
  assign n11948 = ~n11945 & ~n11947 ;
  assign n11949 = \ctl_rf_c7_rf_prot3_reg/NET0131  & ~n2983 ;
  assign n11950 = n3011 & n11949 ;
  assign n11951 = \ctl_rf_c0_rf_prot3_reg/NET0131  & n2983 ;
  assign n11952 = n3050 & n11951 ;
  assign n11953 = ~n11950 & ~n11952 ;
  assign n11954 = n11948 & n11953 ;
  assign n11955 = \ctl_rf_c3_rf_prot3_reg/NET0131  & ~n2983 ;
  assign n11956 = n3024 & n11955 ;
  assign n11957 = \ctl_rf_c6_rf_prot3_reg/NET0131  & n2983 ;
  assign n11958 = n3011 & n11957 ;
  assign n11959 = ~n11956 & ~n11958 ;
  assign n11960 = \ctl_rf_c5_rf_prot3_reg/NET0131  & ~n2983 ;
  assign n11961 = n2999 & n11960 ;
  assign n11962 = \ctl_rf_c4_rf_prot3_reg/NET0131  & n2983 ;
  assign n11963 = n2999 & n11962 ;
  assign n11964 = ~n11961 & ~n11963 ;
  assign n11965 = n11959 & n11964 ;
  assign n11966 = n11954 & n11965 ;
  assign n11967 = \ctl_rf_c2_rf_src_sz_reg[2]/NET0131  & n2983 ;
  assign n11968 = n3024 & n11967 ;
  assign n11969 = \ctl_rf_c1_rf_src_sz_reg[2]/NET0131  & ~n2983 ;
  assign n11970 = n3050 & n11969 ;
  assign n11971 = ~n11968 & ~n11970 ;
  assign n11972 = \ctl_rf_c7_rf_src_sz_reg[2]/NET0131  & ~n2983 ;
  assign n11973 = n3011 & n11972 ;
  assign n11974 = \ctl_rf_c0_rf_src_sz_reg[2]/NET0131  & n2983 ;
  assign n11975 = n3050 & n11974 ;
  assign n11976 = ~n11973 & ~n11975 ;
  assign n11977 = n11971 & n11976 ;
  assign n11978 = \ctl_rf_c3_rf_src_sz_reg[2]/NET0131  & ~n2983 ;
  assign n11979 = n3024 & n11978 ;
  assign n11980 = \ctl_rf_c6_rf_src_sz_reg[2]/NET0131  & n2983 ;
  assign n11981 = n3011 & n11980 ;
  assign n11982 = ~n11979 & ~n11981 ;
  assign n11983 = \ctl_rf_c5_rf_src_sz_reg[2]/NET0131  & ~n2983 ;
  assign n11984 = n2999 & n11983 ;
  assign n11985 = \ctl_rf_c4_rf_src_sz_reg[2]/NET0131  & n2983 ;
  assign n11986 = n2999 & n11985 ;
  assign n11987 = ~n11984 & ~n11986 ;
  assign n11988 = n11982 & n11987 ;
  assign n11989 = n11977 & n11988 ;
  assign n11990 = \h1rdt1_br[13]_pad  & n2767 ;
  assign n11991 = \h1rdt0_dma[13]_pad  & n2793 ;
  assign n11992 = ~n11990 & ~n11991 ;
  assign n11993 = \h1rdt2_dma[13]_pad  & n2786 ;
  assign n11994 = \h1rdt4_br[13]_pad  & n2777 ;
  assign n11995 = ~n11993 & ~n11994 ;
  assign n11996 = n11992 & n11995 ;
  assign n11997 = \h1rdt5_dma[13]_pad  & n2770 ;
  assign n11998 = \h1rdt7_br[13]_pad  & n2751 ;
  assign n11999 = ~n11997 & ~n11998 ;
  assign n12000 = \h1rdt1_dma[13]_pad  & n2760 ;
  assign n12001 = \h1rdt6_br[13]_pad  & n2753 ;
  assign n12002 = ~n12000 & ~n12001 ;
  assign n12003 = n11999 & n12002 ;
  assign n12004 = n11996 & n12003 ;
  assign n12005 = \h1rdt5_br[13]_pad  & n2782 ;
  assign n12006 = \h1rdt4_dma[13]_pad  & n2788 ;
  assign n12007 = ~n12005 & ~n12006 ;
  assign n12008 = \h1rdt6_dma[13]_pad  & n2791 ;
  assign n12009 = \h1rdt3_dma[13]_pad  & n2757 ;
  assign n12010 = ~n12008 & ~n12009 ;
  assign n12011 = n12007 & n12010 ;
  assign n12012 = \h1rdt3_br[13]_pad  & n2765 ;
  assign n12013 = \h1rdt0_br[13]_pad  & n2780 ;
  assign n12014 = ~n12012 & ~n12013 ;
  assign n12015 = \h1rdt2_br[13]_pad  & n2746 ;
  assign n12016 = \h1rdt7_dma[13]_pad  & n2774 ;
  assign n12017 = ~n12015 & ~n12016 ;
  assign n12018 = n12014 & n12017 ;
  assign n12019 = n12011 & n12018 ;
  assign n12020 = n12004 & n12019 ;
  assign n12021 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & n2238 ;
  assign n12022 = \ctl_rf_m0end_reg/NET0131  & ~\ctl_rf_m1end_reg/NET0131  ;
  assign n12023 = ~\ctl_rf_m0end_reg/NET0131  & \ctl_rf_m1end_reg/NET0131  ;
  assign n12024 = ~n12022 & ~n12023 ;
  assign n12025 = n12021 & ~n12024 ;
  assign n12026 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & n2241 ;
  assign n12027 = ~n12024 & n12026 ;
  assign n12028 = ~n12025 & ~n12027 ;
  assign n12029 = ~n12020 & n12028 ;
  assign n12030 = \h1rdt6_dma[21]_pad  & n2791 ;
  assign n12031 = \h1rdt1_br[21]_pad  & n2767 ;
  assign n12032 = ~n12030 & ~n12031 ;
  assign n12033 = \h1rdt5_dma[21]_pad  & n2770 ;
  assign n12034 = \h1rdt5_br[21]_pad  & n2782 ;
  assign n12035 = ~n12033 & ~n12034 ;
  assign n12036 = n12032 & n12035 ;
  assign n12037 = \h1rdt0_br[21]_pad  & n2780 ;
  assign n12038 = \h1rdt3_br[21]_pad  & n2765 ;
  assign n12039 = ~n12037 & ~n12038 ;
  assign n12040 = \h1rdt3_dma[21]_pad  & n2757 ;
  assign n12041 = \h1rdt2_br[21]_pad  & n2746 ;
  assign n12042 = ~n12040 & ~n12041 ;
  assign n12043 = n12039 & n12042 ;
  assign n12044 = n12036 & n12043 ;
  assign n12045 = \h1rdt2_dma[21]_pad  & n2786 ;
  assign n12046 = \h1rdt1_dma[21]_pad  & n2760 ;
  assign n12047 = ~n12045 & ~n12046 ;
  assign n12048 = \h1rdt4_br[21]_pad  & n2777 ;
  assign n12049 = \h1rdt6_br[21]_pad  & n2753 ;
  assign n12050 = ~n12048 & ~n12049 ;
  assign n12051 = n12047 & n12050 ;
  assign n12052 = \h1rdt7_br[21]_pad  & n2751 ;
  assign n12053 = \h1rdt4_dma[21]_pad  & n2788 ;
  assign n12054 = ~n12052 & ~n12053 ;
  assign n12055 = \h1rdt0_dma[21]_pad  & n2793 ;
  assign n12056 = \h1rdt7_dma[21]_pad  & n2774 ;
  assign n12057 = ~n12055 & ~n12056 ;
  assign n12058 = n12054 & n12057 ;
  assign n12059 = n12051 & n12058 ;
  assign n12060 = n12044 & n12059 ;
  assign n12061 = ~n12025 & n12027 ;
  assign n12062 = ~n12060 & n12061 ;
  assign n12063 = ~n12029 & ~n12062 ;
  assign n12064 = \h1rdt2_br[29]_pad  & n2746 ;
  assign n12065 = \h1rdt1_br[29]_pad  & n2767 ;
  assign n12066 = ~n12064 & ~n12065 ;
  assign n12067 = \h1rdt6_br[29]_pad  & n2753 ;
  assign n12068 = \h1rdt4_dma[29]_pad  & n2788 ;
  assign n12069 = ~n12067 & ~n12068 ;
  assign n12070 = n12066 & n12069 ;
  assign n12071 = \h1rdt1_dma[29]_pad  & n2760 ;
  assign n12072 = \h1rdt7_br[29]_pad  & n2751 ;
  assign n12073 = ~n12071 & ~n12072 ;
  assign n12074 = \h1rdt4_br[29]_pad  & n2777 ;
  assign n12075 = \h1rdt0_dma[29]_pad  & n2793 ;
  assign n12076 = ~n12074 & ~n12075 ;
  assign n12077 = n12073 & n12076 ;
  assign n12078 = n12070 & n12077 ;
  assign n12079 = \h1rdt7_dma[29]_pad  & n2774 ;
  assign n12080 = \h1rdt3_dma[29]_pad  & n2757 ;
  assign n12081 = ~n12079 & ~n12080 ;
  assign n12082 = \h1rdt5_dma[29]_pad  & n2770 ;
  assign n12083 = \h1rdt2_dma[29]_pad  & n2786 ;
  assign n12084 = ~n12082 & ~n12083 ;
  assign n12085 = n12081 & n12084 ;
  assign n12086 = \h1rdt3_br[29]_pad  & n2765 ;
  assign n12087 = \h1rdt6_dma[29]_pad  & n2791 ;
  assign n12088 = ~n12086 & ~n12087 ;
  assign n12089 = \h1rdt5_br[29]_pad  & n2782 ;
  assign n12090 = \h1rdt0_br[29]_pad  & n2780 ;
  assign n12091 = ~n12089 & ~n12090 ;
  assign n12092 = n12088 & n12091 ;
  assign n12093 = n12085 & n12092 ;
  assign n12094 = n12078 & n12093 ;
  assign n12095 = n12025 & ~n12094 ;
  assign n12096 = n12063 & ~n12095 ;
  assign n12097 = \h1rdt0_br[14]_pad  & n2780 ;
  assign n12098 = \h1rdt2_br[14]_pad  & n2746 ;
  assign n12099 = ~n12097 & ~n12098 ;
  assign n12100 = \h1rdt6_br[14]_pad  & n2753 ;
  assign n12101 = \h1rdt4_dma[14]_pad  & n2788 ;
  assign n12102 = ~n12100 & ~n12101 ;
  assign n12103 = n12099 & n12102 ;
  assign n12104 = \h1rdt1_br[14]_pad  & n2767 ;
  assign n12105 = \h1rdt7_br[14]_pad  & n2751 ;
  assign n12106 = ~n12104 & ~n12105 ;
  assign n12107 = \h1rdt0_dma[14]_pad  & n2793 ;
  assign n12108 = \h1rdt7_dma[14]_pad  & n2774 ;
  assign n12109 = ~n12107 & ~n12108 ;
  assign n12110 = n12106 & n12109 ;
  assign n12111 = n12103 & n12110 ;
  assign n12112 = \h1rdt4_br[14]_pad  & n2777 ;
  assign n12113 = \h1rdt5_br[14]_pad  & n2782 ;
  assign n12114 = ~n12112 & ~n12113 ;
  assign n12115 = \h1rdt2_dma[14]_pad  & n2786 ;
  assign n12116 = \h1rdt1_dma[14]_pad  & n2760 ;
  assign n12117 = ~n12115 & ~n12116 ;
  assign n12118 = n12114 & n12117 ;
  assign n12119 = \h1rdt3_br[14]_pad  & n2765 ;
  assign n12120 = \h1rdt3_dma[14]_pad  & n2757 ;
  assign n12121 = ~n12119 & ~n12120 ;
  assign n12122 = \h1rdt5_dma[14]_pad  & n2770 ;
  assign n12123 = \h1rdt6_dma[14]_pad  & n2791 ;
  assign n12124 = ~n12122 & ~n12123 ;
  assign n12125 = n12121 & n12124 ;
  assign n12126 = n12118 & n12125 ;
  assign n12127 = n12111 & n12126 ;
  assign n12128 = n12028 & ~n12127 ;
  assign n12129 = \h1rdt1_dma[22]_pad  & n2760 ;
  assign n12130 = \h1rdt5_br[22]_pad  & n2782 ;
  assign n12131 = ~n12129 & ~n12130 ;
  assign n12132 = \h1rdt7_dma[22]_pad  & n2774 ;
  assign n12133 = \h1rdt4_dma[22]_pad  & n2788 ;
  assign n12134 = ~n12132 & ~n12133 ;
  assign n12135 = n12131 & n12134 ;
  assign n12136 = \h1rdt3_dma[22]_pad  & n2757 ;
  assign n12137 = \h1rdt3_br[22]_pad  & n2765 ;
  assign n12138 = ~n12136 & ~n12137 ;
  assign n12139 = \h1rdt6_dma[22]_pad  & n2791 ;
  assign n12140 = \h1rdt0_dma[22]_pad  & n2793 ;
  assign n12141 = ~n12139 & ~n12140 ;
  assign n12142 = n12138 & n12141 ;
  assign n12143 = n12135 & n12142 ;
  assign n12144 = \h1rdt0_br[22]_pad  & n2780 ;
  assign n12145 = \h1rdt6_br[22]_pad  & n2753 ;
  assign n12146 = ~n12144 & ~n12145 ;
  assign n12147 = \h1rdt4_br[22]_pad  & n2777 ;
  assign n12148 = \h1rdt5_dma[22]_pad  & n2770 ;
  assign n12149 = ~n12147 & ~n12148 ;
  assign n12150 = n12146 & n12149 ;
  assign n12151 = \h1rdt7_br[22]_pad  & n2751 ;
  assign n12152 = \h1rdt2_br[22]_pad  & n2746 ;
  assign n12153 = ~n12151 & ~n12152 ;
  assign n12154 = \h1rdt1_br[22]_pad  & n2767 ;
  assign n12155 = \h1rdt2_dma[22]_pad  & n2786 ;
  assign n12156 = ~n12154 & ~n12155 ;
  assign n12157 = n12153 & n12156 ;
  assign n12158 = n12150 & n12157 ;
  assign n12159 = n12143 & n12158 ;
  assign n12160 = n12061 & ~n12159 ;
  assign n12161 = ~n12128 & ~n12160 ;
  assign n12162 = \h1rdt5_dma[30]_pad  & n2770 ;
  assign n12163 = \h1rdt0_br[30]_pad  & n2780 ;
  assign n12164 = ~n12162 & ~n12163 ;
  assign n12165 = \h1rdt0_dma[30]_pad  & n2793 ;
  assign n12166 = \h1rdt6_br[30]_pad  & n2753 ;
  assign n12167 = ~n12165 & ~n12166 ;
  assign n12168 = n12164 & n12167 ;
  assign n12169 = \h1rdt5_br[30]_pad  & n2782 ;
  assign n12170 = \h1rdt7_br[30]_pad  & n2751 ;
  assign n12171 = ~n12169 & ~n12170 ;
  assign n12172 = \h1rdt4_dma[30]_pad  & n2788 ;
  assign n12173 = \h1rdt4_br[30]_pad  & n2777 ;
  assign n12174 = ~n12172 & ~n12173 ;
  assign n12175 = n12171 & n12174 ;
  assign n12176 = n12168 & n12175 ;
  assign n12177 = \h1rdt7_dma[30]_pad  & n2774 ;
  assign n12178 = \h1rdt6_dma[30]_pad  & n2791 ;
  assign n12179 = ~n12177 & ~n12178 ;
  assign n12180 = \h1rdt2_br[30]_pad  & n2746 ;
  assign n12181 = \h1rdt1_br[30]_pad  & n2767 ;
  assign n12182 = ~n12180 & ~n12181 ;
  assign n12183 = n12179 & n12182 ;
  assign n12184 = \h1rdt3_br[30]_pad  & n2765 ;
  assign n12185 = \h1rdt2_dma[30]_pad  & n2786 ;
  assign n12186 = ~n12184 & ~n12185 ;
  assign n12187 = \h1rdt1_dma[30]_pad  & n2760 ;
  assign n12188 = \h1rdt3_dma[30]_pad  & n2757 ;
  assign n12189 = ~n12187 & ~n12188 ;
  assign n12190 = n12186 & n12189 ;
  assign n12191 = n12183 & n12190 ;
  assign n12192 = n12176 & n12191 ;
  assign n12193 = n12025 & ~n12192 ;
  assign n12194 = n12161 & ~n12193 ;
  assign n12195 = \h1rdt6_br[15]_pad  & n2753 ;
  assign n12196 = \h1rdt4_br[15]_pad  & n2777 ;
  assign n12197 = ~n12195 & ~n12196 ;
  assign n12198 = \h1rdt2_br[15]_pad  & n2746 ;
  assign n12199 = \h1rdt1_dma[15]_pad  & n2760 ;
  assign n12200 = ~n12198 & ~n12199 ;
  assign n12201 = n12197 & n12200 ;
  assign n12202 = \h1rdt0_dma[15]_pad  & n2793 ;
  assign n12203 = \h1rdt7_br[15]_pad  & n2751 ;
  assign n12204 = ~n12202 & ~n12203 ;
  assign n12205 = \h1rdt1_br[15]_pad  & n2767 ;
  assign n12206 = \h1rdt2_dma[15]_pad  & n2786 ;
  assign n12207 = ~n12205 & ~n12206 ;
  assign n12208 = n12204 & n12207 ;
  assign n12209 = n12201 & n12208 ;
  assign n12210 = \h1rdt5_br[15]_pad  & n2782 ;
  assign n12211 = \h1rdt6_dma[15]_pad  & n2791 ;
  assign n12212 = ~n12210 & ~n12211 ;
  assign n12213 = \h1rdt7_dma[15]_pad  & n2774 ;
  assign n12214 = \h1rdt4_dma[15]_pad  & n2788 ;
  assign n12215 = ~n12213 & ~n12214 ;
  assign n12216 = n12212 & n12215 ;
  assign n12217 = \h1rdt3_br[15]_pad  & n2765 ;
  assign n12218 = \h1rdt5_dma[15]_pad  & n2770 ;
  assign n12219 = ~n12217 & ~n12218 ;
  assign n12220 = \h1rdt3_dma[15]_pad  & n2757 ;
  assign n12221 = \h1rdt0_br[15]_pad  & n2780 ;
  assign n12222 = ~n12220 & ~n12221 ;
  assign n12223 = n12219 & n12222 ;
  assign n12224 = n12216 & n12223 ;
  assign n12225 = n12209 & n12224 ;
  assign n12226 = n12028 & ~n12225 ;
  assign n12227 = \h1rdt5_dma[23]_pad  & n2770 ;
  assign n12228 = \h1rdt3_dma[23]_pad  & n2757 ;
  assign n12229 = ~n12227 & ~n12228 ;
  assign n12230 = \h1rdt5_br[23]_pad  & n2782 ;
  assign n12231 = \h1rdt0_dma[23]_pad  & n2793 ;
  assign n12232 = ~n12230 & ~n12231 ;
  assign n12233 = n12229 & n12232 ;
  assign n12234 = \h1rdt4_br[23]_pad  & n2777 ;
  assign n12235 = \h1rdt3_br[23]_pad  & n2765 ;
  assign n12236 = ~n12234 & ~n12235 ;
  assign n12237 = \h1rdt1_dma[23]_pad  & n2760 ;
  assign n12238 = \h1rdt4_dma[23]_pad  & n2788 ;
  assign n12239 = ~n12237 & ~n12238 ;
  assign n12240 = n12236 & n12239 ;
  assign n12241 = n12233 & n12240 ;
  assign n12242 = \h1rdt0_br[23]_pad  & n2780 ;
  assign n12243 = \h1rdt6_dma[23]_pad  & n2791 ;
  assign n12244 = ~n12242 & ~n12243 ;
  assign n12245 = \h1rdt7_dma[23]_pad  & n2774 ;
  assign n12246 = \h1rdt2_dma[23]_pad  & n2786 ;
  assign n12247 = ~n12245 & ~n12246 ;
  assign n12248 = n12244 & n12247 ;
  assign n12249 = \h1rdt7_br[23]_pad  & n2751 ;
  assign n12250 = \h1rdt1_br[23]_pad  & n2767 ;
  assign n12251 = ~n12249 & ~n12250 ;
  assign n12252 = \h1rdt2_br[23]_pad  & n2746 ;
  assign n12253 = \h1rdt6_br[23]_pad  & n2753 ;
  assign n12254 = ~n12252 & ~n12253 ;
  assign n12255 = n12251 & n12254 ;
  assign n12256 = n12248 & n12255 ;
  assign n12257 = n12241 & n12256 ;
  assign n12258 = n12061 & ~n12257 ;
  assign n12259 = ~n12226 & ~n12258 ;
  assign n12260 = \h1rdt5_dma[31]_pad  & n2770 ;
  assign n12261 = \h1rdt0_br[31]_pad  & n2780 ;
  assign n12262 = ~n12260 & ~n12261 ;
  assign n12263 = \h1rdt1_br[31]_pad  & n2767 ;
  assign n12264 = \h1rdt6_br[31]_pad  & n2753 ;
  assign n12265 = ~n12263 & ~n12264 ;
  assign n12266 = n12262 & n12265 ;
  assign n12267 = \h1rdt7_dma[31]_pad  & n2774 ;
  assign n12268 = \h1rdt7_br[31]_pad  & n2751 ;
  assign n12269 = ~n12267 & ~n12268 ;
  assign n12270 = \h1rdt2_br[31]_pad  & n2746 ;
  assign n12271 = \h1rdt4_br[31]_pad  & n2777 ;
  assign n12272 = ~n12270 & ~n12271 ;
  assign n12273 = n12269 & n12272 ;
  assign n12274 = n12266 & n12273 ;
  assign n12275 = \h1rdt4_dma[31]_pad  & n2788 ;
  assign n12276 = \h1rdt0_dma[31]_pad  & n2793 ;
  assign n12277 = ~n12275 & ~n12276 ;
  assign n12278 = \h1rdt5_br[31]_pad  & n2782 ;
  assign n12279 = \h1rdt6_dma[31]_pad  & n2791 ;
  assign n12280 = ~n12278 & ~n12279 ;
  assign n12281 = n12277 & n12280 ;
  assign n12282 = \h1rdt3_br[31]_pad  & n2765 ;
  assign n12283 = \h1rdt2_dma[31]_pad  & n2786 ;
  assign n12284 = ~n12282 & ~n12283 ;
  assign n12285 = \h1rdt1_dma[31]_pad  & n2760 ;
  assign n12286 = \h1rdt3_dma[31]_pad  & n2757 ;
  assign n12287 = ~n12285 & ~n12286 ;
  assign n12288 = n12284 & n12287 ;
  assign n12289 = n12281 & n12288 ;
  assign n12290 = n12274 & n12289 ;
  assign n12291 = n12025 & ~n12290 ;
  assign n12292 = n12259 & ~n12291 ;
  assign n12293 = \h1rdt6_dma[16]_pad  & n2791 ;
  assign n12294 = \h1rdt2_br[16]_pad  & n2746 ;
  assign n12295 = ~n12293 & ~n12294 ;
  assign n12296 = \h1rdt0_dma[16]_pad  & n2793 ;
  assign n12297 = \h1rdt5_br[16]_pad  & n2782 ;
  assign n12298 = ~n12296 & ~n12297 ;
  assign n12299 = n12295 & n12298 ;
  assign n12300 = \h1rdt6_br[16]_pad  & n2753 ;
  assign n12301 = \h1rdt3_br[16]_pad  & n2765 ;
  assign n12302 = ~n12300 & ~n12301 ;
  assign n12303 = \h1rdt4_dma[16]_pad  & n2788 ;
  assign n12304 = \h1rdt1_br[16]_pad  & n2767 ;
  assign n12305 = ~n12303 & ~n12304 ;
  assign n12306 = n12302 & n12305 ;
  assign n12307 = n12299 & n12306 ;
  assign n12308 = \h1rdt3_dma[16]_pad  & n2757 ;
  assign n12309 = \h1rdt5_dma[16]_pad  & n2770 ;
  assign n12310 = ~n12308 & ~n12309 ;
  assign n12311 = \h1rdt2_dma[16]_pad  & n2786 ;
  assign n12312 = \h1rdt1_dma[16]_pad  & n2760 ;
  assign n12313 = ~n12311 & ~n12312 ;
  assign n12314 = n12310 & n12313 ;
  assign n12315 = \h1rdt7_br[16]_pad  & n2751 ;
  assign n12316 = \h1rdt4_br[16]_pad  & n2777 ;
  assign n12317 = ~n12315 & ~n12316 ;
  assign n12318 = \h1rdt0_br[16]_pad  & n2780 ;
  assign n12319 = \h1rdt7_dma[16]_pad  & n2774 ;
  assign n12320 = ~n12318 & ~n12319 ;
  assign n12321 = n12317 & n12320 ;
  assign n12322 = n12314 & n12321 ;
  assign n12323 = n12307 & n12322 ;
  assign n12324 = n12028 & ~n12323 ;
  assign n12325 = \h1rdt1_br[8]_pad  & n2767 ;
  assign n12326 = \h1rdt5_br[8]_pad  & n2782 ;
  assign n12327 = ~n12325 & ~n12326 ;
  assign n12328 = \h1rdt0_dma[8]_pad  & n2793 ;
  assign n12329 = \h1rdt6_dma[8]_pad  & n2791 ;
  assign n12330 = ~n12328 & ~n12329 ;
  assign n12331 = n12327 & n12330 ;
  assign n12332 = \h1rdt0_br[8]_pad  & n2780 ;
  assign n12333 = \h1rdt3_br[8]_pad  & n2765 ;
  assign n12334 = ~n12332 & ~n12333 ;
  assign n12335 = \h1rdt4_dma[8]_pad  & n2788 ;
  assign n12336 = \h1rdt7_dma[8]_pad  & n2774 ;
  assign n12337 = ~n12335 & ~n12336 ;
  assign n12338 = n12334 & n12337 ;
  assign n12339 = n12331 & n12338 ;
  assign n12340 = \h1rdt2_dma[8]_pad  & n2786 ;
  assign n12341 = \h1rdt1_dma[8]_pad  & n2760 ;
  assign n12342 = ~n12340 & ~n12341 ;
  assign n12343 = \h1rdt3_dma[8]_pad  & n2757 ;
  assign n12344 = \h1rdt5_dma[8]_pad  & n2770 ;
  assign n12345 = ~n12343 & ~n12344 ;
  assign n12346 = n12342 & n12345 ;
  assign n12347 = \h1rdt7_br[8]_pad  & n2751 ;
  assign n12348 = \h1rdt6_br[8]_pad  & n2753 ;
  assign n12349 = ~n12347 & ~n12348 ;
  assign n12350 = \h1rdt4_br[8]_pad  & n2777 ;
  assign n12351 = \h1rdt2_br[8]_pad  & n2746 ;
  assign n12352 = ~n12350 & ~n12351 ;
  assign n12353 = n12349 & n12352 ;
  assign n12354 = n12346 & n12353 ;
  assign n12355 = n12339 & n12354 ;
  assign n12356 = n12061 & ~n12355 ;
  assign n12357 = ~n12324 & ~n12356 ;
  assign n12358 = \h1rdt5_dma[0]_pad  & n2770 ;
  assign n12359 = \h1rdt0_br[0]_pad  & n2780 ;
  assign n12360 = ~n12358 & ~n12359 ;
  assign n12361 = \h1rdt0_dma[0]_pad  & n2793 ;
  assign n12362 = \h1rdt4_br[0]_pad  & n2777 ;
  assign n12363 = ~n12361 & ~n12362 ;
  assign n12364 = n12360 & n12363 ;
  assign n12365 = \h1rdt2_br[0]_pad  & n2746 ;
  assign n12366 = \h1rdt7_br[0]_pad  & n2751 ;
  assign n12367 = ~n12365 & ~n12366 ;
  assign n12368 = \h1rdt4_dma[0]_pad  & n2788 ;
  assign n12369 = \h1rdt6_br[0]_pad  & n2753 ;
  assign n12370 = ~n12368 & ~n12369 ;
  assign n12371 = n12367 & n12370 ;
  assign n12372 = n12364 & n12371 ;
  assign n12373 = \h1rdt6_dma[0]_pad  & n2791 ;
  assign n12374 = \h1rdt7_dma[0]_pad  & n2774 ;
  assign n12375 = ~n12373 & ~n12374 ;
  assign n12376 = \h1rdt5_br[0]_pad  & n2782 ;
  assign n12377 = \h1rdt1_br[0]_pad  & n2767 ;
  assign n12378 = ~n12376 & ~n12377 ;
  assign n12379 = n12375 & n12378 ;
  assign n12380 = \h1rdt3_br[0]_pad  & n2765 ;
  assign n12381 = \h1rdt2_dma[0]_pad  & n2786 ;
  assign n12382 = ~n12380 & ~n12381 ;
  assign n12383 = \h1rdt1_dma[0]_pad  & n2760 ;
  assign n12384 = \h1rdt3_dma[0]_pad  & n2757 ;
  assign n12385 = ~n12383 & ~n12384 ;
  assign n12386 = n12382 & n12385 ;
  assign n12387 = n12379 & n12386 ;
  assign n12388 = n12372 & n12387 ;
  assign n12389 = n12025 & ~n12388 ;
  assign n12390 = n12357 & ~n12389 ;
  assign n12391 = \h1rdt2_br[17]_pad  & n2746 ;
  assign n12392 = \h1rdt6_dma[17]_pad  & n2791 ;
  assign n12393 = ~n12391 & ~n12392 ;
  assign n12394 = \h1rdt5_dma[17]_pad  & n2770 ;
  assign n12395 = \h1rdt5_br[17]_pad  & n2782 ;
  assign n12396 = ~n12394 & ~n12395 ;
  assign n12397 = n12393 & n12396 ;
  assign n12398 = \h1rdt2_dma[17]_pad  & n2786 ;
  assign n12399 = \h1rdt3_br[17]_pad  & n2765 ;
  assign n12400 = ~n12398 & ~n12399 ;
  assign n12401 = \h1rdt3_dma[17]_pad  & n2757 ;
  assign n12402 = \h1rdt7_dma[17]_pad  & n2774 ;
  assign n12403 = ~n12401 & ~n12402 ;
  assign n12404 = n12400 & n12403 ;
  assign n12405 = n12397 & n12404 ;
  assign n12406 = \h1rdt6_br[17]_pad  & n2753 ;
  assign n12407 = \h1rdt4_br[17]_pad  & n2777 ;
  assign n12408 = ~n12406 & ~n12407 ;
  assign n12409 = \h1rdt0_br[17]_pad  & n2780 ;
  assign n12410 = \h1rdt1_dma[17]_pad  & n2760 ;
  assign n12411 = ~n12409 & ~n12410 ;
  assign n12412 = n12408 & n12411 ;
  assign n12413 = \h1rdt7_br[17]_pad  & n2751 ;
  assign n12414 = \h1rdt4_dma[17]_pad  & n2788 ;
  assign n12415 = ~n12413 & ~n12414 ;
  assign n12416 = \h1rdt0_dma[17]_pad  & n2793 ;
  assign n12417 = \h1rdt1_br[17]_pad  & n2767 ;
  assign n12418 = ~n12416 & ~n12417 ;
  assign n12419 = n12415 & n12418 ;
  assign n12420 = n12412 & n12419 ;
  assign n12421 = n12405 & n12420 ;
  assign n12422 = n12028 & ~n12421 ;
  assign n12423 = \h1rdt2_dma[9]_pad  & n2786 ;
  assign n12424 = \h1rdt1_dma[9]_pad  & n2760 ;
  assign n12425 = ~n12423 & ~n12424 ;
  assign n12426 = \h1rdt4_dma[9]_pad  & n2788 ;
  assign n12427 = \h1rdt3_dma[9]_pad  & n2757 ;
  assign n12428 = ~n12426 & ~n12427 ;
  assign n12429 = n12425 & n12428 ;
  assign n12430 = \h1rdt5_br[9]_pad  & n2782 ;
  assign n12431 = \h1rdt7_br[9]_pad  & n2751 ;
  assign n12432 = ~n12430 & ~n12431 ;
  assign n12433 = \h1rdt0_dma[9]_pad  & n2793 ;
  assign n12434 = \h1rdt5_dma[9]_pad  & n2770 ;
  assign n12435 = ~n12433 & ~n12434 ;
  assign n12436 = n12432 & n12435 ;
  assign n12437 = n12429 & n12436 ;
  assign n12438 = \h1rdt6_dma[9]_pad  & n2791 ;
  assign n12439 = \h1rdt7_dma[9]_pad  & n2774 ;
  assign n12440 = ~n12438 & ~n12439 ;
  assign n12441 = \h1rdt2_br[9]_pad  & n2746 ;
  assign n12442 = \h1rdt1_br[9]_pad  & n2767 ;
  assign n12443 = ~n12441 & ~n12442 ;
  assign n12444 = n12440 & n12443 ;
  assign n12445 = \h1rdt3_br[9]_pad  & n2765 ;
  assign n12446 = \h1rdt0_br[9]_pad  & n2780 ;
  assign n12447 = ~n12445 & ~n12446 ;
  assign n12448 = \h1rdt6_br[9]_pad  & n2753 ;
  assign n12449 = \h1rdt4_br[9]_pad  & n2777 ;
  assign n12450 = ~n12448 & ~n12449 ;
  assign n12451 = n12447 & n12450 ;
  assign n12452 = n12444 & n12451 ;
  assign n12453 = n12437 & n12452 ;
  assign n12454 = n12061 & ~n12453 ;
  assign n12455 = ~n12422 & ~n12454 ;
  assign n12456 = \h1rdt2_dma[1]_pad  & n2786 ;
  assign n12457 = \h1rdt1_dma[1]_pad  & n2760 ;
  assign n12458 = ~n12456 & ~n12457 ;
  assign n12459 = \h1rdt6_dma[1]_pad  & n2791 ;
  assign n12460 = \h1rdt3_dma[1]_pad  & n2757 ;
  assign n12461 = ~n12459 & ~n12460 ;
  assign n12462 = n12458 & n12461 ;
  assign n12463 = \h1rdt0_dma[1]_pad  & n2793 ;
  assign n12464 = \h1rdt7_br[1]_pad  & n2751 ;
  assign n12465 = ~n12463 & ~n12464 ;
  assign n12466 = \h1rdt7_dma[1]_pad  & n2774 ;
  assign n12467 = \h1rdt5_dma[1]_pad  & n2770 ;
  assign n12468 = ~n12466 & ~n12467 ;
  assign n12469 = n12465 & n12468 ;
  assign n12470 = n12462 & n12469 ;
  assign n12471 = \h1rdt2_br[1]_pad  & n2746 ;
  assign n12472 = \h1rdt1_br[1]_pad  & n2767 ;
  assign n12473 = ~n12471 & ~n12472 ;
  assign n12474 = \h1rdt5_br[1]_pad  & n2782 ;
  assign n12475 = \h1rdt4_dma[1]_pad  & n2788 ;
  assign n12476 = ~n12474 & ~n12475 ;
  assign n12477 = n12473 & n12476 ;
  assign n12478 = \h1rdt3_br[1]_pad  & n2765 ;
  assign n12479 = \h1rdt0_br[1]_pad  & n2780 ;
  assign n12480 = ~n12478 & ~n12479 ;
  assign n12481 = \h1rdt4_br[1]_pad  & n2777 ;
  assign n12482 = \h1rdt6_br[1]_pad  & n2753 ;
  assign n12483 = ~n12481 & ~n12482 ;
  assign n12484 = n12480 & n12483 ;
  assign n12485 = n12477 & n12484 ;
  assign n12486 = n12470 & n12485 ;
  assign n12487 = n12025 & ~n12486 ;
  assign n12488 = n12455 & ~n12487 ;
  assign n12489 = \h1rdt1_br[18]_pad  & n2767 ;
  assign n12490 = \h1rdt7_dma[18]_pad  & n2774 ;
  assign n12491 = ~n12489 & ~n12490 ;
  assign n12492 = \h1rdt0_dma[18]_pad  & n2793 ;
  assign n12493 = \h1rdt5_br[18]_pad  & n2782 ;
  assign n12494 = ~n12492 & ~n12493 ;
  assign n12495 = n12491 & n12494 ;
  assign n12496 = \h1rdt6_br[18]_pad  & n2753 ;
  assign n12497 = \h1rdt3_br[18]_pad  & n2765 ;
  assign n12498 = ~n12496 & ~n12497 ;
  assign n12499 = \h1rdt4_dma[18]_pad  & n2788 ;
  assign n12500 = \h1rdt6_dma[18]_pad  & n2791 ;
  assign n12501 = ~n12499 & ~n12500 ;
  assign n12502 = n12498 & n12501 ;
  assign n12503 = n12495 & n12502 ;
  assign n12504 = \h1rdt3_dma[18]_pad  & n2757 ;
  assign n12505 = \h1rdt5_dma[18]_pad  & n2770 ;
  assign n12506 = ~n12504 & ~n12505 ;
  assign n12507 = \h1rdt2_dma[18]_pad  & n2786 ;
  assign n12508 = \h1rdt1_dma[18]_pad  & n2760 ;
  assign n12509 = ~n12507 & ~n12508 ;
  assign n12510 = n12506 & n12509 ;
  assign n12511 = \h1rdt7_br[18]_pad  & n2751 ;
  assign n12512 = \h1rdt4_br[18]_pad  & n2777 ;
  assign n12513 = ~n12511 & ~n12512 ;
  assign n12514 = \h1rdt0_br[18]_pad  & n2780 ;
  assign n12515 = \h1rdt2_br[18]_pad  & n2746 ;
  assign n12516 = ~n12514 & ~n12515 ;
  assign n12517 = n12513 & n12516 ;
  assign n12518 = n12510 & n12517 ;
  assign n12519 = n12503 & n12518 ;
  assign n12520 = n12028 & ~n12519 ;
  assign n12521 = \h1rdt2_dma[10]_pad  & n2786 ;
  assign n12522 = \h1rdt0_dma[10]_pad  & n2793 ;
  assign n12523 = ~n12521 & ~n12522 ;
  assign n12524 = \h1rdt3_dma[10]_pad  & n2757 ;
  assign n12525 = \h1rdt1_dma[10]_pad  & n2760 ;
  assign n12526 = ~n12524 & ~n12525 ;
  assign n12527 = n12523 & n12526 ;
  assign n12528 = \h1rdt6_br[10]_pad  & n2753 ;
  assign n12529 = \h1rdt3_br[10]_pad  & n2765 ;
  assign n12530 = ~n12528 & ~n12529 ;
  assign n12531 = \h1rdt5_dma[10]_pad  & n2770 ;
  assign n12532 = \h1rdt4_br[10]_pad  & n2777 ;
  assign n12533 = ~n12531 & ~n12532 ;
  assign n12534 = n12530 & n12533 ;
  assign n12535 = n12527 & n12534 ;
  assign n12536 = \h1rdt7_dma[10]_pad  & n2774 ;
  assign n12537 = \h1rdt6_dma[10]_pad  & n2791 ;
  assign n12538 = ~n12536 & ~n12537 ;
  assign n12539 = \h1rdt0_br[10]_pad  & n2780 ;
  assign n12540 = \h1rdt5_br[10]_pad  & n2782 ;
  assign n12541 = ~n12539 & ~n12540 ;
  assign n12542 = n12538 & n12541 ;
  assign n12543 = \h1rdt7_br[10]_pad  & n2751 ;
  assign n12544 = \h1rdt2_br[10]_pad  & n2746 ;
  assign n12545 = ~n12543 & ~n12544 ;
  assign n12546 = \h1rdt4_dma[10]_pad  & n2788 ;
  assign n12547 = \h1rdt1_br[10]_pad  & n2767 ;
  assign n12548 = ~n12546 & ~n12547 ;
  assign n12549 = n12545 & n12548 ;
  assign n12550 = n12542 & n12549 ;
  assign n12551 = n12535 & n12550 ;
  assign n12552 = n12061 & ~n12551 ;
  assign n12553 = ~n12520 & ~n12552 ;
  assign n12554 = \h1rdt5_dma[2]_pad  & n2770 ;
  assign n12555 = \h1rdt3_dma[2]_pad  & n2757 ;
  assign n12556 = ~n12554 & ~n12555 ;
  assign n12557 = \h1rdt6_br[2]_pad  & n2753 ;
  assign n12558 = \h1rdt2_dma[2]_pad  & n2786 ;
  assign n12559 = ~n12557 & ~n12558 ;
  assign n12560 = n12556 & n12559 ;
  assign n12561 = \h1rdt2_br[2]_pad  & n2746 ;
  assign n12562 = \h1rdt7_br[2]_pad  & n2751 ;
  assign n12563 = ~n12561 & ~n12562 ;
  assign n12564 = \h1rdt4_br[2]_pad  & n2777 ;
  assign n12565 = \h1rdt6_dma[2]_pad  & n2791 ;
  assign n12566 = ~n12564 & ~n12565 ;
  assign n12567 = n12563 & n12566 ;
  assign n12568 = n12560 & n12567 ;
  assign n12569 = \h1rdt0_dma[2]_pad  & n2793 ;
  assign n12570 = \h1rdt1_dma[2]_pad  & n2760 ;
  assign n12571 = ~n12569 & ~n12570 ;
  assign n12572 = \h1rdt4_dma[2]_pad  & n2788 ;
  assign n12573 = \h1rdt7_dma[2]_pad  & n2774 ;
  assign n12574 = ~n12572 & ~n12573 ;
  assign n12575 = n12571 & n12574 ;
  assign n12576 = \h1rdt3_br[2]_pad  & n2765 ;
  assign n12577 = \h1rdt5_br[2]_pad  & n2782 ;
  assign n12578 = ~n12576 & ~n12577 ;
  assign n12579 = \h1rdt0_br[2]_pad  & n2780 ;
  assign n12580 = \h1rdt1_br[2]_pad  & n2767 ;
  assign n12581 = ~n12579 & ~n12580 ;
  assign n12582 = n12578 & n12581 ;
  assign n12583 = n12575 & n12582 ;
  assign n12584 = n12568 & n12583 ;
  assign n12585 = n12025 & ~n12584 ;
  assign n12586 = n12553 & ~n12585 ;
  assign n12587 = \h1rdt2_br[19]_pad  & n2746 ;
  assign n12588 = \h1rdt7_dma[19]_pad  & n2774 ;
  assign n12589 = ~n12587 & ~n12588 ;
  assign n12590 = \h1rdt3_dma[19]_pad  & n2757 ;
  assign n12591 = \h1rdt5_br[19]_pad  & n2782 ;
  assign n12592 = ~n12590 & ~n12591 ;
  assign n12593 = n12589 & n12592 ;
  assign n12594 = \h1rdt6_br[19]_pad  & n2753 ;
  assign n12595 = \h1rdt7_br[19]_pad  & n2751 ;
  assign n12596 = ~n12594 & ~n12595 ;
  assign n12597 = \h1rdt6_dma[19]_pad  & n2791 ;
  assign n12598 = \h1rdt0_br[19]_pad  & n2780 ;
  assign n12599 = ~n12597 & ~n12598 ;
  assign n12600 = n12596 & n12599 ;
  assign n12601 = n12593 & n12600 ;
  assign n12602 = \h1rdt5_dma[19]_pad  & n2770 ;
  assign n12603 = \h1rdt0_dma[19]_pad  & n2793 ;
  assign n12604 = ~n12602 & ~n12603 ;
  assign n12605 = \h1rdt2_dma[19]_pad  & n2786 ;
  assign n12606 = \h1rdt1_dma[19]_pad  & n2760 ;
  assign n12607 = ~n12605 & ~n12606 ;
  assign n12608 = n12604 & n12607 ;
  assign n12609 = \h1rdt3_br[19]_pad  & n2765 ;
  assign n12610 = \h1rdt4_br[19]_pad  & n2777 ;
  assign n12611 = ~n12609 & ~n12610 ;
  assign n12612 = \h1rdt4_dma[19]_pad  & n2788 ;
  assign n12613 = \h1rdt1_br[19]_pad  & n2767 ;
  assign n12614 = ~n12612 & ~n12613 ;
  assign n12615 = n12611 & n12614 ;
  assign n12616 = n12608 & n12615 ;
  assign n12617 = n12601 & n12616 ;
  assign n12618 = n12028 & ~n12617 ;
  assign n12619 = \h1rdt3_dma[11]_pad  & n2757 ;
  assign n12620 = \h1rdt0_br[11]_pad  & n2780 ;
  assign n12621 = ~n12619 & ~n12620 ;
  assign n12622 = \h1rdt6_dma[11]_pad  & n2791 ;
  assign n12623 = \h1rdt6_br[11]_pad  & n2753 ;
  assign n12624 = ~n12622 & ~n12623 ;
  assign n12625 = n12621 & n12624 ;
  assign n12626 = \h1rdt0_dma[11]_pad  & n2793 ;
  assign n12627 = \h1rdt7_br[11]_pad  & n2751 ;
  assign n12628 = ~n12626 & ~n12627 ;
  assign n12629 = \h1rdt7_dma[11]_pad  & n2774 ;
  assign n12630 = \h1rdt4_br[11]_pad  & n2777 ;
  assign n12631 = ~n12629 & ~n12630 ;
  assign n12632 = n12628 & n12631 ;
  assign n12633 = n12625 & n12632 ;
  assign n12634 = \h1rdt2_br[11]_pad  & n2746 ;
  assign n12635 = \h1rdt1_br[11]_pad  & n2767 ;
  assign n12636 = ~n12634 & ~n12635 ;
  assign n12637 = \h1rdt5_br[11]_pad  & n2782 ;
  assign n12638 = \h1rdt4_dma[11]_pad  & n2788 ;
  assign n12639 = ~n12637 & ~n12638 ;
  assign n12640 = n12636 & n12639 ;
  assign n12641 = \h1rdt3_br[11]_pad  & n2765 ;
  assign n12642 = \h1rdt2_dma[11]_pad  & n2786 ;
  assign n12643 = ~n12641 & ~n12642 ;
  assign n12644 = \h1rdt1_dma[11]_pad  & n2760 ;
  assign n12645 = \h1rdt5_dma[11]_pad  & n2770 ;
  assign n12646 = ~n12644 & ~n12645 ;
  assign n12647 = n12643 & n12646 ;
  assign n12648 = n12640 & n12647 ;
  assign n12649 = n12633 & n12648 ;
  assign n12650 = n12061 & ~n12649 ;
  assign n12651 = ~n12618 & ~n12650 ;
  assign n12652 = \h1rdt5_dma[3]_pad  & n2770 ;
  assign n12653 = \h1rdt3_dma[3]_pad  & n2757 ;
  assign n12654 = ~n12652 & ~n12653 ;
  assign n12655 = \h1rdt6_dma[3]_pad  & n2791 ;
  assign n12656 = \h1rdt5_br[3]_pad  & n2782 ;
  assign n12657 = ~n12655 & ~n12656 ;
  assign n12658 = n12654 & n12657 ;
  assign n12659 = \h1rdt6_br[3]_pad  & n2753 ;
  assign n12660 = \h1rdt3_br[3]_pad  & n2765 ;
  assign n12661 = ~n12659 & ~n12660 ;
  assign n12662 = \h1rdt7_dma[3]_pad  & n2774 ;
  assign n12663 = \h1rdt4_dma[3]_pad  & n2788 ;
  assign n12664 = ~n12662 & ~n12663 ;
  assign n12665 = n12661 & n12664 ;
  assign n12666 = n12658 & n12665 ;
  assign n12667 = \h1rdt2_br[3]_pad  & n2746 ;
  assign n12668 = \h1rdt1_br[3]_pad  & n2767 ;
  assign n12669 = ~n12667 & ~n12668 ;
  assign n12670 = \h1rdt0_dma[3]_pad  & n2793 ;
  assign n12671 = \h1rdt4_br[3]_pad  & n2777 ;
  assign n12672 = ~n12670 & ~n12671 ;
  assign n12673 = n12669 & n12672 ;
  assign n12674 = \h1rdt7_br[3]_pad  & n2751 ;
  assign n12675 = \h1rdt0_br[3]_pad  & n2780 ;
  assign n12676 = ~n12674 & ~n12675 ;
  assign n12677 = \h1rdt2_dma[3]_pad  & n2786 ;
  assign n12678 = \h1rdt1_dma[3]_pad  & n2760 ;
  assign n12679 = ~n12677 & ~n12678 ;
  assign n12680 = n12676 & n12679 ;
  assign n12681 = n12673 & n12680 ;
  assign n12682 = n12666 & n12681 ;
  assign n12683 = n12025 & ~n12682 ;
  assign n12684 = n12651 & ~n12683 ;
  assign n12685 = \h1rdt0_br[25]_pad  & n2780 ;
  assign n12686 = \h1rdt4_br[25]_pad  & n2777 ;
  assign n12687 = ~n12685 & ~n12686 ;
  assign n12688 = \h1rdt2_dma[25]_pad  & n2786 ;
  assign n12689 = \h1rdt4_dma[25]_pad  & n2788 ;
  assign n12690 = ~n12688 & ~n12689 ;
  assign n12691 = n12687 & n12690 ;
  assign n12692 = \h1rdt5_br[25]_pad  & n2782 ;
  assign n12693 = \h1rdt7_br[25]_pad  & n2751 ;
  assign n12694 = ~n12692 & ~n12693 ;
  assign n12695 = \h1rdt1_dma[25]_pad  & n2760 ;
  assign n12696 = \h1rdt6_br[25]_pad  & n2753 ;
  assign n12697 = ~n12695 & ~n12696 ;
  assign n12698 = n12694 & n12697 ;
  assign n12699 = n12691 & n12698 ;
  assign n12700 = \h1rdt7_dma[25]_pad  & n2774 ;
  assign n12701 = \h1rdt2_br[25]_pad  & n2746 ;
  assign n12702 = ~n12700 & ~n12701 ;
  assign n12703 = \h1rdt6_dma[25]_pad  & n2791 ;
  assign n12704 = \h1rdt1_br[25]_pad  & n2767 ;
  assign n12705 = ~n12703 & ~n12704 ;
  assign n12706 = n12702 & n12705 ;
  assign n12707 = \h1rdt3_br[25]_pad  & n2765 ;
  assign n12708 = \h1rdt0_dma[25]_pad  & n2793 ;
  assign n12709 = ~n12707 & ~n12708 ;
  assign n12710 = \h1rdt5_dma[25]_pad  & n2770 ;
  assign n12711 = \h1rdt3_dma[25]_pad  & n2757 ;
  assign n12712 = ~n12710 & ~n12711 ;
  assign n12713 = n12709 & n12712 ;
  assign n12714 = n12706 & n12713 ;
  assign n12715 = n12699 & n12714 ;
  assign n12716 = n12061 & ~n12715 ;
  assign n12717 = n12028 & ~n12486 ;
  assign n12718 = ~n12716 & ~n12717 ;
  assign n12719 = n12025 & ~n12421 ;
  assign n12720 = n12718 & ~n12719 ;
  assign n12721 = \h1rdt5_dma[20]_pad  & n2770 ;
  assign n12722 = \h1rdt3_dma[20]_pad  & n2757 ;
  assign n12723 = ~n12721 & ~n12722 ;
  assign n12724 = \h1rdt4_br[20]_pad  & n2777 ;
  assign n12725 = \h1rdt4_dma[20]_pad  & n2788 ;
  assign n12726 = ~n12724 & ~n12725 ;
  assign n12727 = n12723 & n12726 ;
  assign n12728 = \h1rdt1_dma[20]_pad  & n2760 ;
  assign n12729 = \h1rdt3_br[20]_pad  & n2765 ;
  assign n12730 = ~n12728 & ~n12729 ;
  assign n12731 = \h1rdt6_br[20]_pad  & n2753 ;
  assign n12732 = \h1rdt5_br[20]_pad  & n2782 ;
  assign n12733 = ~n12731 & ~n12732 ;
  assign n12734 = n12730 & n12733 ;
  assign n12735 = n12727 & n12734 ;
  assign n12736 = \h1rdt0_br[20]_pad  & n2780 ;
  assign n12737 = \h1rdt2_br[20]_pad  & n2746 ;
  assign n12738 = ~n12736 & ~n12737 ;
  assign n12739 = \h1rdt1_br[20]_pad  & n2767 ;
  assign n12740 = \h1rdt2_dma[20]_pad  & n2786 ;
  assign n12741 = ~n12739 & ~n12740 ;
  assign n12742 = n12738 & n12741 ;
  assign n12743 = \h1rdt7_br[20]_pad  & n2751 ;
  assign n12744 = \h1rdt0_dma[20]_pad  & n2793 ;
  assign n12745 = ~n12743 & ~n12744 ;
  assign n12746 = \h1rdt6_dma[20]_pad  & n2791 ;
  assign n12747 = \h1rdt7_dma[20]_pad  & n2774 ;
  assign n12748 = ~n12746 & ~n12747 ;
  assign n12749 = n12745 & n12748 ;
  assign n12750 = n12742 & n12749 ;
  assign n12751 = n12735 & n12750 ;
  assign n12752 = n12028 & ~n12751 ;
  assign n12753 = \h1rdt0_dma[12]_pad  & n2793 ;
  assign n12754 = \h1rdt4_br[12]_pad  & n2777 ;
  assign n12755 = ~n12753 & ~n12754 ;
  assign n12756 = \h1rdt2_dma[12]_pad  & n2786 ;
  assign n12757 = \h1rdt4_dma[12]_pad  & n2788 ;
  assign n12758 = ~n12756 & ~n12757 ;
  assign n12759 = n12755 & n12758 ;
  assign n12760 = \h1rdt3_dma[12]_pad  & n2757 ;
  assign n12761 = \h1rdt3_br[12]_pad  & n2765 ;
  assign n12762 = ~n12760 & ~n12761 ;
  assign n12763 = \h1rdt6_dma[12]_pad  & n2791 ;
  assign n12764 = \h1rdt6_br[12]_pad  & n2753 ;
  assign n12765 = ~n12763 & ~n12764 ;
  assign n12766 = n12762 & n12765 ;
  assign n12767 = n12759 & n12766 ;
  assign n12768 = \h1rdt1_dma[12]_pad  & n2760 ;
  assign n12769 = \h1rdt2_br[12]_pad  & n2746 ;
  assign n12770 = ~n12768 & ~n12769 ;
  assign n12771 = \h1rdt1_br[12]_pad  & n2767 ;
  assign n12772 = \h1rdt5_dma[12]_pad  & n2770 ;
  assign n12773 = ~n12771 & ~n12772 ;
  assign n12774 = n12770 & n12773 ;
  assign n12775 = \h1rdt7_br[12]_pad  & n2751 ;
  assign n12776 = \h1rdt0_br[12]_pad  & n2780 ;
  assign n12777 = ~n12775 & ~n12776 ;
  assign n12778 = \h1rdt5_br[12]_pad  & n2782 ;
  assign n12779 = \h1rdt7_dma[12]_pad  & n2774 ;
  assign n12780 = ~n12778 & ~n12779 ;
  assign n12781 = n12777 & n12780 ;
  assign n12782 = n12774 & n12781 ;
  assign n12783 = n12767 & n12782 ;
  assign n12784 = n12061 & ~n12783 ;
  assign n12785 = ~n12752 & ~n12784 ;
  assign n12786 = \h1rdt6_dma[4]_pad  & n2791 ;
  assign n12787 = \h1rdt5_br[4]_pad  & n2782 ;
  assign n12788 = ~n12786 & ~n12787 ;
  assign n12789 = \h1rdt5_dma[4]_pad  & n2770 ;
  assign n12790 = \h1rdt1_br[4]_pad  & n2767 ;
  assign n12791 = ~n12789 & ~n12790 ;
  assign n12792 = n12788 & n12791 ;
  assign n12793 = \h1rdt0_br[4]_pad  & n2780 ;
  assign n12794 = \h1rdt3_br[4]_pad  & n2765 ;
  assign n12795 = ~n12793 & ~n12794 ;
  assign n12796 = \h1rdt3_dma[4]_pad  & n2757 ;
  assign n12797 = \h1rdt2_br[4]_pad  & n2746 ;
  assign n12798 = ~n12796 & ~n12797 ;
  assign n12799 = n12795 & n12798 ;
  assign n12800 = n12792 & n12799 ;
  assign n12801 = \h1rdt2_dma[4]_pad  & n2786 ;
  assign n12802 = \h1rdt1_dma[4]_pad  & n2760 ;
  assign n12803 = ~n12801 & ~n12802 ;
  assign n12804 = \h1rdt6_br[4]_pad  & n2753 ;
  assign n12805 = \h1rdt4_br[4]_pad  & n2777 ;
  assign n12806 = ~n12804 & ~n12805 ;
  assign n12807 = n12803 & n12806 ;
  assign n12808 = \h1rdt7_br[4]_pad  & n2751 ;
  assign n12809 = \h1rdt4_dma[4]_pad  & n2788 ;
  assign n12810 = ~n12808 & ~n12809 ;
  assign n12811 = \h1rdt0_dma[4]_pad  & n2793 ;
  assign n12812 = \h1rdt7_dma[4]_pad  & n2774 ;
  assign n12813 = ~n12811 & ~n12812 ;
  assign n12814 = n12810 & n12813 ;
  assign n12815 = n12807 & n12814 ;
  assign n12816 = n12800 & n12815 ;
  assign n12817 = n12025 & ~n12816 ;
  assign n12818 = n12785 & ~n12817 ;
  assign n12819 = ~n12020 & n12061 ;
  assign n12820 = n12028 & ~n12060 ;
  assign n12821 = ~n12819 & ~n12820 ;
  assign n12822 = \h1rdt6_dma[5]_pad  & n2791 ;
  assign n12823 = \h1rdt2_br[5]_pad  & n2746 ;
  assign n12824 = ~n12822 & ~n12823 ;
  assign n12825 = \h1rdt5_dma[5]_pad  & n2770 ;
  assign n12826 = \h1rdt5_br[5]_pad  & n2782 ;
  assign n12827 = ~n12825 & ~n12826 ;
  assign n12828 = n12824 & n12827 ;
  assign n12829 = \h1rdt0_br[5]_pad  & n2780 ;
  assign n12830 = \h1rdt3_br[5]_pad  & n2765 ;
  assign n12831 = ~n12829 & ~n12830 ;
  assign n12832 = \h1rdt3_dma[5]_pad  & n2757 ;
  assign n12833 = \h1rdt1_br[5]_pad  & n2767 ;
  assign n12834 = ~n12832 & ~n12833 ;
  assign n12835 = n12831 & n12834 ;
  assign n12836 = n12828 & n12835 ;
  assign n12837 = \h1rdt2_dma[5]_pad  & n2786 ;
  assign n12838 = \h1rdt1_dma[5]_pad  & n2760 ;
  assign n12839 = ~n12837 & ~n12838 ;
  assign n12840 = \h1rdt4_br[5]_pad  & n2777 ;
  assign n12841 = \h1rdt6_br[5]_pad  & n2753 ;
  assign n12842 = ~n12840 & ~n12841 ;
  assign n12843 = n12839 & n12842 ;
  assign n12844 = \h1rdt7_br[5]_pad  & n2751 ;
  assign n12845 = \h1rdt4_dma[5]_pad  & n2788 ;
  assign n12846 = ~n12844 & ~n12845 ;
  assign n12847 = \h1rdt0_dma[5]_pad  & n2793 ;
  assign n12848 = \h1rdt7_dma[5]_pad  & n2774 ;
  assign n12849 = ~n12847 & ~n12848 ;
  assign n12850 = n12846 & n12849 ;
  assign n12851 = n12843 & n12850 ;
  assign n12852 = n12836 & n12851 ;
  assign n12853 = n12025 & ~n12852 ;
  assign n12854 = n12821 & ~n12853 ;
  assign n12855 = n12061 & ~n12127 ;
  assign n12856 = n12028 & ~n12159 ;
  assign n12857 = ~n12855 & ~n12856 ;
  assign n12858 = \h1rdt6_dma[6]_pad  & n2791 ;
  assign n12859 = \h1rdt6_br[6]_pad  & n2753 ;
  assign n12860 = ~n12858 & ~n12859 ;
  assign n12861 = \h1rdt0_br[6]_pad  & n2780 ;
  assign n12862 = \h1rdt1_br[6]_pad  & n2767 ;
  assign n12863 = ~n12861 & ~n12862 ;
  assign n12864 = n12860 & n12863 ;
  assign n12865 = \h1rdt5_br[6]_pad  & n2782 ;
  assign n12866 = \h1rdt7_br[6]_pad  & n2751 ;
  assign n12867 = ~n12865 & ~n12866 ;
  assign n12868 = \h1rdt0_dma[6]_pad  & n2793 ;
  assign n12869 = \h1rdt2_br[6]_pad  & n2746 ;
  assign n12870 = ~n12868 & ~n12869 ;
  assign n12871 = n12867 & n12870 ;
  assign n12872 = n12864 & n12871 ;
  assign n12873 = \h1rdt4_br[6]_pad  & n2777 ;
  assign n12874 = \h1rdt4_dma[6]_pad  & n2788 ;
  assign n12875 = ~n12873 & ~n12874 ;
  assign n12876 = \h1rdt1_dma[6]_pad  & n2760 ;
  assign n12877 = \h1rdt2_dma[6]_pad  & n2786 ;
  assign n12878 = ~n12876 & ~n12877 ;
  assign n12879 = n12875 & n12878 ;
  assign n12880 = \h1rdt3_br[6]_pad  & n2765 ;
  assign n12881 = \h1rdt5_dma[6]_pad  & n2770 ;
  assign n12882 = ~n12880 & ~n12881 ;
  assign n12883 = \h1rdt3_dma[6]_pad  & n2757 ;
  assign n12884 = \h1rdt7_dma[6]_pad  & n2774 ;
  assign n12885 = ~n12883 & ~n12884 ;
  assign n12886 = n12882 & n12885 ;
  assign n12887 = n12879 & n12886 ;
  assign n12888 = n12872 & n12887 ;
  assign n12889 = n12025 & ~n12888 ;
  assign n12890 = n12857 & ~n12889 ;
  assign n12891 = n12061 & ~n12225 ;
  assign n12892 = n12028 & ~n12257 ;
  assign n12893 = ~n12891 & ~n12892 ;
  assign n12894 = \h1rdt1_dma[7]_pad  & n2760 ;
  assign n12895 = \h1rdt3_dma[7]_pad  & n2757 ;
  assign n12896 = ~n12894 & ~n12895 ;
  assign n12897 = \h1rdt0_dma[7]_pad  & n2793 ;
  assign n12898 = \h1rdt0_br[7]_pad  & n2780 ;
  assign n12899 = ~n12897 & ~n12898 ;
  assign n12900 = n12896 & n12899 ;
  assign n12901 = \h1rdt2_br[7]_pad  & n2746 ;
  assign n12902 = \h1rdt7_br[7]_pad  & n2751 ;
  assign n12903 = ~n12901 & ~n12902 ;
  assign n12904 = \h1rdt4_dma[7]_pad  & n2788 ;
  assign n12905 = \h1rdt5_dma[7]_pad  & n2770 ;
  assign n12906 = ~n12904 & ~n12905 ;
  assign n12907 = n12903 & n12906 ;
  assign n12908 = n12900 & n12907 ;
  assign n12909 = \h1rdt5_br[7]_pad  & n2782 ;
  assign n12910 = \h1rdt6_br[7]_pad  & n2753 ;
  assign n12911 = ~n12909 & ~n12910 ;
  assign n12912 = \h1rdt4_br[7]_pad  & n2777 ;
  assign n12913 = \h1rdt1_br[7]_pad  & n2767 ;
  assign n12914 = ~n12912 & ~n12913 ;
  assign n12915 = n12911 & n12914 ;
  assign n12916 = \h1rdt3_br[7]_pad  & n2765 ;
  assign n12917 = \h1rdt6_dma[7]_pad  & n2791 ;
  assign n12918 = ~n12916 & ~n12917 ;
  assign n12919 = \h1rdt7_dma[7]_pad  & n2774 ;
  assign n12920 = \h1rdt2_dma[7]_pad  & n2786 ;
  assign n12921 = ~n12919 & ~n12920 ;
  assign n12922 = n12918 & n12921 ;
  assign n12923 = n12915 & n12922 ;
  assign n12924 = n12908 & n12923 ;
  assign n12925 = n12025 & ~n12924 ;
  assign n12926 = n12893 & ~n12925 ;
  assign n12927 = \h1rdt4_br[24]_pad  & n2777 ;
  assign n12928 = \h1rdt0_br[24]_pad  & n2780 ;
  assign n12929 = ~n12927 & ~n12928 ;
  assign n12930 = \h1rdt5_br[24]_pad  & n2782 ;
  assign n12931 = \h1rdt2_br[24]_pad  & n2746 ;
  assign n12932 = ~n12930 & ~n12931 ;
  assign n12933 = n12929 & n12932 ;
  assign n12934 = \h1rdt6_dma[24]_pad  & n2791 ;
  assign n12935 = \h1rdt7_br[24]_pad  & n2751 ;
  assign n12936 = ~n12934 & ~n12935 ;
  assign n12937 = \h1rdt0_dma[24]_pad  & n2793 ;
  assign n12938 = \h1rdt1_br[24]_pad  & n2767 ;
  assign n12939 = ~n12937 & ~n12938 ;
  assign n12940 = n12936 & n12939 ;
  assign n12941 = n12933 & n12940 ;
  assign n12942 = \h1rdt7_dma[24]_pad  & n2774 ;
  assign n12943 = \h1rdt4_dma[24]_pad  & n2788 ;
  assign n12944 = ~n12942 & ~n12943 ;
  assign n12945 = \h1rdt5_dma[24]_pad  & n2770 ;
  assign n12946 = \h1rdt3_dma[24]_pad  & n2757 ;
  assign n12947 = ~n12945 & ~n12946 ;
  assign n12948 = n12944 & n12947 ;
  assign n12949 = \h1rdt3_br[24]_pad  & n2765 ;
  assign n12950 = \h1rdt2_dma[24]_pad  & n2786 ;
  assign n12951 = ~n12949 & ~n12950 ;
  assign n12952 = \h1rdt1_dma[24]_pad  & n2760 ;
  assign n12953 = \h1rdt6_br[24]_pad  & n2753 ;
  assign n12954 = ~n12952 & ~n12953 ;
  assign n12955 = n12951 & n12954 ;
  assign n12956 = n12948 & n12955 ;
  assign n12957 = n12941 & n12956 ;
  assign n12958 = n12028 & ~n12957 ;
  assign n12959 = n12061 & ~n12388 ;
  assign n12960 = ~n12958 & ~n12959 ;
  assign n12961 = n12025 & ~n12355 ;
  assign n12962 = n12960 & ~n12961 ;
  assign n12963 = n12028 & ~n12715 ;
  assign n12964 = n12061 & ~n12486 ;
  assign n12965 = ~n12963 & ~n12964 ;
  assign n12966 = n12025 & ~n12453 ;
  assign n12967 = n12965 & ~n12966 ;
  assign n12968 = \h1rdt0_br[26]_pad  & n2780 ;
  assign n12969 = \h1rdt4_dma[26]_pad  & n2788 ;
  assign n12970 = ~n12968 & ~n12969 ;
  assign n12971 = \h1rdt2_dma[26]_pad  & n2786 ;
  assign n12972 = \h1rdt6_br[26]_pad  & n2753 ;
  assign n12973 = ~n12971 & ~n12972 ;
  assign n12974 = n12970 & n12973 ;
  assign n12975 = \h1rdt1_br[26]_pad  & n2767 ;
  assign n12976 = \h1rdt3_br[26]_pad  & n2765 ;
  assign n12977 = ~n12975 & ~n12976 ;
  assign n12978 = \h1rdt0_dma[26]_pad  & n2793 ;
  assign n12979 = \h1rdt5_br[26]_pad  & n2782 ;
  assign n12980 = ~n12978 & ~n12979 ;
  assign n12981 = n12977 & n12980 ;
  assign n12982 = n12974 & n12981 ;
  assign n12983 = \h1rdt1_dma[26]_pad  & n2760 ;
  assign n12984 = \h1rdt5_dma[26]_pad  & n2770 ;
  assign n12985 = ~n12983 & ~n12984 ;
  assign n12986 = \h1rdt3_dma[26]_pad  & n2757 ;
  assign n12987 = \h1rdt2_br[26]_pad  & n2746 ;
  assign n12988 = ~n12986 & ~n12987 ;
  assign n12989 = n12985 & n12988 ;
  assign n12990 = \h1rdt7_br[26]_pad  & n2751 ;
  assign n12991 = \h1rdt7_dma[26]_pad  & n2774 ;
  assign n12992 = ~n12990 & ~n12991 ;
  assign n12993 = \h1rdt6_dma[26]_pad  & n2791 ;
  assign n12994 = \h1rdt4_br[26]_pad  & n2777 ;
  assign n12995 = ~n12993 & ~n12994 ;
  assign n12996 = n12992 & n12995 ;
  assign n12997 = n12989 & n12996 ;
  assign n12998 = n12982 & n12997 ;
  assign n12999 = n12028 & ~n12998 ;
  assign n13000 = n12061 & ~n12584 ;
  assign n13001 = ~n12999 & ~n13000 ;
  assign n13002 = n12025 & ~n12551 ;
  assign n13003 = n13001 & ~n13002 ;
  assign n13004 = \h1rdt6_dma[27]_pad  & n2791 ;
  assign n13005 = \h1rdt2_br[27]_pad  & n2746 ;
  assign n13006 = ~n13004 & ~n13005 ;
  assign n13007 = \h1rdt3_dma[27]_pad  & n2757 ;
  assign n13008 = \h1rdt1_dma[27]_pad  & n2760 ;
  assign n13009 = ~n13007 & ~n13008 ;
  assign n13010 = n13006 & n13009 ;
  assign n13011 = \h1rdt0_br[27]_pad  & n2780 ;
  assign n13012 = \h1rdt7_br[27]_pad  & n2751 ;
  assign n13013 = ~n13011 & ~n13012 ;
  assign n13014 = \h1rdt5_dma[27]_pad  & n2770 ;
  assign n13015 = \h1rdt2_dma[27]_pad  & n2786 ;
  assign n13016 = ~n13014 & ~n13015 ;
  assign n13017 = n13013 & n13016 ;
  assign n13018 = n13010 & n13017 ;
  assign n13019 = \h1rdt6_br[27]_pad  & n2753 ;
  assign n13020 = \h1rdt4_br[27]_pad  & n2777 ;
  assign n13021 = ~n13019 & ~n13020 ;
  assign n13022 = \h1rdt5_br[27]_pad  & n2782 ;
  assign n13023 = \h1rdt0_dma[27]_pad  & n2793 ;
  assign n13024 = ~n13022 & ~n13023 ;
  assign n13025 = n13021 & n13024 ;
  assign n13026 = \h1rdt3_br[27]_pad  & n2765 ;
  assign n13027 = \h1rdt1_br[27]_pad  & n2767 ;
  assign n13028 = ~n13026 & ~n13027 ;
  assign n13029 = \h1rdt7_dma[27]_pad  & n2774 ;
  assign n13030 = \h1rdt4_dma[27]_pad  & n2788 ;
  assign n13031 = ~n13029 & ~n13030 ;
  assign n13032 = n13028 & n13031 ;
  assign n13033 = n13025 & n13032 ;
  assign n13034 = n13018 & n13033 ;
  assign n13035 = n12028 & ~n13034 ;
  assign n13036 = n12061 & ~n12682 ;
  assign n13037 = ~n13035 & ~n13036 ;
  assign n13038 = n12025 & ~n12649 ;
  assign n13039 = n13037 & ~n13038 ;
  assign n13040 = \h1rdt6_dma[28]_pad  & n2791 ;
  assign n13041 = \h1rdt2_br[28]_pad  & n2746 ;
  assign n13042 = ~n13040 & ~n13041 ;
  assign n13043 = \h1rdt3_dma[28]_pad  & n2757 ;
  assign n13044 = \h1rdt5_br[28]_pad  & n2782 ;
  assign n13045 = ~n13043 & ~n13044 ;
  assign n13046 = n13042 & n13045 ;
  assign n13047 = \h1rdt0_br[28]_pad  & n2780 ;
  assign n13048 = \h1rdt3_br[28]_pad  & n2765 ;
  assign n13049 = ~n13047 & ~n13048 ;
  assign n13050 = \h1rdt5_dma[28]_pad  & n2770 ;
  assign n13051 = \h1rdt1_br[28]_pad  & n2767 ;
  assign n13052 = ~n13050 & ~n13051 ;
  assign n13053 = n13049 & n13052 ;
  assign n13054 = n13046 & n13053 ;
  assign n13055 = \h1rdt2_dma[28]_pad  & n2786 ;
  assign n13056 = \h1rdt1_dma[28]_pad  & n2760 ;
  assign n13057 = ~n13055 & ~n13056 ;
  assign n13058 = \h1rdt4_br[28]_pad  & n2777 ;
  assign n13059 = \h1rdt6_br[28]_pad  & n2753 ;
  assign n13060 = ~n13058 & ~n13059 ;
  assign n13061 = n13057 & n13060 ;
  assign n13062 = \h1rdt7_br[28]_pad  & n2751 ;
  assign n13063 = \h1rdt4_dma[28]_pad  & n2788 ;
  assign n13064 = ~n13062 & ~n13063 ;
  assign n13065 = \h1rdt0_dma[28]_pad  & n2793 ;
  assign n13066 = \h1rdt7_dma[28]_pad  & n2774 ;
  assign n13067 = ~n13065 & ~n13066 ;
  assign n13068 = n13064 & n13067 ;
  assign n13069 = n13061 & n13068 ;
  assign n13070 = n13054 & n13069 ;
  assign n13071 = n12028 & ~n13070 ;
  assign n13072 = n12061 & ~n12816 ;
  assign n13073 = ~n13071 & ~n13072 ;
  assign n13074 = n12025 & ~n12783 ;
  assign n13075 = n13073 & ~n13074 ;
  assign n13076 = n12061 & ~n12852 ;
  assign n13077 = n12028 & ~n12094 ;
  assign n13078 = ~n13076 & ~n13077 ;
  assign n13079 = ~n12020 & n12025 ;
  assign n13080 = n13078 & ~n13079 ;
  assign n13081 = n12061 & ~n12998 ;
  assign n13082 = n12028 & ~n12584 ;
  assign n13083 = ~n13081 & ~n13082 ;
  assign n13084 = n12025 & ~n12519 ;
  assign n13085 = n13083 & ~n13084 ;
  assign n13086 = n12061 & ~n12888 ;
  assign n13087 = n12028 & ~n12192 ;
  assign n13088 = ~n13086 & ~n13087 ;
  assign n13089 = n12025 & ~n12127 ;
  assign n13090 = n13088 & ~n13089 ;
  assign n13091 = n12061 & ~n12924 ;
  assign n13092 = n12028 & ~n12290 ;
  assign n13093 = ~n13091 & ~n13092 ;
  assign n13094 = n12025 & ~n12225 ;
  assign n13095 = n13093 & ~n13094 ;
  assign n13096 = n12061 & ~n13034 ;
  assign n13097 = n12028 & ~n12682 ;
  assign n13098 = ~n13096 & ~n13097 ;
  assign n13099 = n12025 & ~n12617 ;
  assign n13100 = n13098 & ~n13099 ;
  assign n13101 = n12061 & ~n13070 ;
  assign n13102 = n12028 & ~n12816 ;
  assign n13103 = ~n13101 & ~n13102 ;
  assign n13104 = n12025 & ~n12751 ;
  assign n13105 = n13103 & ~n13104 ;
  assign n13106 = n12028 & ~n12852 ;
  assign n13107 = n12061 & ~n12094 ;
  assign n13108 = ~n13106 & ~n13107 ;
  assign n13109 = n12025 & ~n12060 ;
  assign n13110 = n13108 & ~n13109 ;
  assign n13111 = n12028 & ~n12888 ;
  assign n13112 = n12061 & ~n12192 ;
  assign n13113 = ~n13111 & ~n13112 ;
  assign n13114 = n12025 & ~n12159 ;
  assign n13115 = n13113 & ~n13114 ;
  assign n13116 = n12028 & ~n12924 ;
  assign n13117 = n12061 & ~n12290 ;
  assign n13118 = ~n13116 & ~n13117 ;
  assign n13119 = n12025 & ~n12257 ;
  assign n13120 = n13118 & ~n13119 ;
  assign n13121 = n12061 & ~n12323 ;
  assign n13122 = n12028 & ~n12355 ;
  assign n13123 = ~n13121 & ~n13122 ;
  assign n13124 = n12025 & ~n12957 ;
  assign n13125 = n13123 & ~n13124 ;
  assign n13126 = n12061 & ~n12421 ;
  assign n13127 = n12028 & ~n12453 ;
  assign n13128 = ~n13126 & ~n13127 ;
  assign n13129 = n12025 & ~n12715 ;
  assign n13130 = n13128 & ~n13129 ;
  assign n13131 = n12061 & ~n12957 ;
  assign n13132 = n12028 & ~n12388 ;
  assign n13133 = ~n13131 & ~n13132 ;
  assign n13134 = n12025 & ~n12323 ;
  assign n13135 = n13133 & ~n13134 ;
  assign n13136 = n12061 & ~n12519 ;
  assign n13137 = n12028 & ~n12551 ;
  assign n13138 = ~n13136 & ~n13137 ;
  assign n13139 = n12025 & ~n12998 ;
  assign n13140 = n13138 & ~n13139 ;
  assign n13141 = n12061 & ~n12617 ;
  assign n13142 = n12028 & ~n12649 ;
  assign n13143 = ~n13141 & ~n13142 ;
  assign n13144 = n12025 & ~n13034 ;
  assign n13145 = n13143 & ~n13144 ;
  assign n13146 = n12061 & ~n12751 ;
  assign n13147 = n12028 & ~n12783 ;
  assign n13148 = ~n13146 & ~n13147 ;
  assign n13149 = n12025 & ~n13070 ;
  assign n13150 = n13148 & ~n13149 ;
  assign n13151 = \dma_ack[4]_pad  & n3003 ;
  assign n13152 = ~\ctl_rf_c4_rf_chabt_reg/NET0131  & \ctl_rf_c4_rf_mode_reg/NET0131  ;
  assign n13153 = \de_de_st_reg[5]/NET0131  & ~\dma_ack[4]_pad  ;
  assign n13154 = n13152 & n13153 ;
  assign n13155 = n2983 & n13154 ;
  assign n13156 = n2999 & n13155 ;
  assign n13157 = ~n13151 & ~n13156 ;
  assign n13158 = \dma_ack[1]_pad  & n3077 ;
  assign n13159 = ~\ctl_rf_c1_rf_chabt_reg/NET0131  & \ctl_rf_c1_rf_mode_reg/NET0131  ;
  assign n13160 = \de_de_st_reg[5]/NET0131  & ~\dma_ack[1]_pad  ;
  assign n13161 = n13159 & n13160 ;
  assign n13162 = ~n2983 & n13161 ;
  assign n13163 = n3050 & n13162 ;
  assign n13164 = ~n13158 & ~n13163 ;
  assign n13165 = \de_de_st_reg[1]/NET0131  & n4506 ;
  assign n13166 = ~\ahb_mst0_m0_m1_diff_tx_reg/NET0131  & ~n13165 ;
  assign n13167 = ~\ahb_mst0_m0_m1_diff_tx_reg/NET0131  & ~n2823 ;
  assign n13168 = ~n2814 & n13167 ;
  assign n13169 = ~n13166 & ~n13168 ;
  assign n13170 = ~\de_de_st_reg[5]/NET0131  & n13169 ;
  assign n13171 = \dma_ack[7]_pad  & n3088 ;
  assign n13172 = ~\ctl_rf_c7_rf_chabt_reg/NET0131  & \ctl_rf_c7_rf_mode_reg/NET0131  ;
  assign n13173 = \de_de_st_reg[5]/NET0131  & ~\dma_ack[7]_pad  ;
  assign n13174 = n13172 & n13173 ;
  assign n13175 = ~n2983 & n13174 ;
  assign n13176 = n3011 & n13175 ;
  assign n13177 = ~n13171 & ~n13176 ;
  assign n13178 = \dma_ack[2]_pad  & n3065 ;
  assign n13179 = ~\ctl_rf_c2_rf_chabt_reg/NET0131  & \ctl_rf_c2_rf_mode_reg/NET0131  ;
  assign n13180 = \de_de_st_reg[5]/NET0131  & ~\dma_ack[2]_pad  ;
  assign n13181 = n13179 & n13180 ;
  assign n13182 = n2983 & n13181 ;
  assign n13183 = n3024 & n13182 ;
  assign n13184 = ~n13178 & ~n13183 ;
  assign n13185 = \dma_ack[3]_pad  & n3029 ;
  assign n13186 = ~\ctl_rf_c3_rf_chabt_reg/NET0131  & \ctl_rf_c3_rf_mode_reg/NET0131  ;
  assign n13187 = \de_de_st_reg[5]/NET0131  & ~\dma_ack[3]_pad  ;
  assign n13188 = n13186 & n13187 ;
  assign n13189 = ~n2983 & n13188 ;
  assign n13190 = n3024 & n13189 ;
  assign n13191 = ~n13185 & ~n13190 ;
  assign n13192 = \dma_ack[5]_pad  & n3040 ;
  assign n13193 = ~\ctl_rf_c5_rf_chabt_reg/NET0131  & \ctl_rf_c5_rf_mode_reg/NET0131  ;
  assign n13194 = \de_de_st_reg[5]/NET0131  & ~\dma_ack[5]_pad  ;
  assign n13195 = n13193 & n13194 ;
  assign n13196 = ~n2983 & n13195 ;
  assign n13197 = n2999 & n13196 ;
  assign n13198 = ~n13192 & ~n13197 ;
  assign n13199 = \dma_ack[6]_pad  & n3015 ;
  assign n13200 = ~\ctl_rf_c6_rf_chabt_reg/NET0131  & \ctl_rf_c6_rf_mode_reg/NET0131  ;
  assign n13201 = \de_de_st_reg[5]/NET0131  & ~\dma_ack[6]_pad  ;
  assign n13202 = n13200 & n13201 ;
  assign n13203 = n2983 & n13202 ;
  assign n13204 = n3011 & n13203 ;
  assign n13205 = ~n13199 & ~n13204 ;
  assign n13206 = \dma_ack[0]_pad  & n3054 ;
  assign n13207 = ~\ctl_rf_c0_rf_chabt_reg/NET0131  & \ctl_rf_c0_rf_mode_reg/NET0131  ;
  assign n13208 = \de_de_st_reg[5]/NET0131  & ~\dma_ack[0]_pad  ;
  assign n13209 = n13207 & n13208 ;
  assign n13210 = n2983 & n13209 ;
  assign n13211 = n3050 & n13210 ;
  assign n13212 = ~n13206 & ~n13211 ;
  assign n13213 = \dma_tc[2]_pad  & n3065 ;
  assign n13214 = n2983 & n13179 ;
  assign n13215 = n3024 & n13214 ;
  assign n13216 = \de_de_st_reg[5]/NET0131  & ~\dma_tc[2]_pad  ;
  assign n13217 = n2814 & n13216 ;
  assign n13218 = n13215 & n13217 ;
  assign n13219 = ~n13213 & ~n13218 ;
  assign n13220 = \dma_tc[7]_pad  & n3088 ;
  assign n13221 = ~n2983 & n13172 ;
  assign n13222 = n3011 & n13221 ;
  assign n13223 = \de_de_st_reg[5]/NET0131  & ~\dma_tc[7]_pad  ;
  assign n13224 = n2814 & n13223 ;
  assign n13225 = n13222 & n13224 ;
  assign n13226 = ~n13220 & ~n13225 ;
  assign n13227 = \dma_tc[3]_pad  & n3029 ;
  assign n13228 = ~n2983 & n13186 ;
  assign n13229 = n3024 & n13228 ;
  assign n13230 = \de_de_st_reg[5]/NET0131  & ~\dma_tc[3]_pad  ;
  assign n13231 = n2814 & n13230 ;
  assign n13232 = n13229 & n13231 ;
  assign n13233 = ~n13227 & ~n13232 ;
  assign n13234 = \dma_tc[5]_pad  & n3040 ;
  assign n13235 = ~n2983 & n13193 ;
  assign n13236 = n2999 & n13235 ;
  assign n13237 = \de_de_st_reg[5]/NET0131  & ~\dma_tc[5]_pad  ;
  assign n13238 = n2814 & n13237 ;
  assign n13239 = n13236 & n13238 ;
  assign n13240 = ~n13234 & ~n13239 ;
  assign n13241 = \dma_tc[0]_pad  & n3054 ;
  assign n13242 = n2983 & n13207 ;
  assign n13243 = n3050 & n13242 ;
  assign n13244 = \de_de_st_reg[5]/NET0131  & ~\dma_tc[0]_pad  ;
  assign n13245 = n2814 & n13244 ;
  assign n13246 = n13243 & n13245 ;
  assign n13247 = ~n13241 & ~n13246 ;
  assign n13248 = \dma_tc[1]_pad  & n3077 ;
  assign n13249 = ~n2983 & n13159 ;
  assign n13250 = n3050 & n13249 ;
  assign n13251 = \de_de_st_reg[5]/NET0131  & ~\dma_tc[1]_pad  ;
  assign n13252 = n2814 & n13251 ;
  assign n13253 = n13250 & n13252 ;
  assign n13254 = ~n13248 & ~n13253 ;
  assign n13255 = \dma_tc[4]_pad  & n3003 ;
  assign n13256 = n2983 & n13152 ;
  assign n13257 = n2999 & n13256 ;
  assign n13258 = \de_de_st_reg[5]/NET0131  & ~\dma_tc[4]_pad  ;
  assign n13259 = n2814 & n13258 ;
  assign n13260 = n13257 & n13259 ;
  assign n13261 = ~n13255 & ~n13260 ;
  assign n13262 = \dma_tc[6]_pad  & n3015 ;
  assign n13263 = n2983 & n13200 ;
  assign n13264 = n3011 & n13263 ;
  assign n13265 = \de_de_st_reg[5]/NET0131  & ~\dma_tc[6]_pad  ;
  assign n13266 = n2814 & n13265 ;
  assign n13267 = n13264 & n13266 ;
  assign n13268 = ~n13262 & ~n13267 ;
  assign n13269 = \ctl_rf_be_d1_reg[0]/P0001  & n3756 ;
  assign n13270 = n2274 & n13269 ;
  assign n13271 = \ctl_rf_be_d1_reg[0]/P0001  & n4065 ;
  assign n13272 = n2274 & n13271 ;
  assign n13273 = n2289 & n13271 ;
  assign n13274 = n2289 & n13269 ;
  assign n13275 = ~n3763 & n11126 ;
  assign n13276 = ~n3762 & n13275 ;
  assign n13277 = \ctl_rf_be_d1_reg[1]/P0001  & ~n4105 ;
  assign n13278 = n2252 & n13269 ;
  assign n13279 = n2252 & n13271 ;
  assign n13280 = \ctl_rf_be_d1_reg[3]/P0001  & ~n4070 ;
  assign n13281 = ~n3763 & n11116 ;
  assign n13282 = ~n3762 & n13281 ;
  assign n13283 = \ctl_rf_be_d1_reg[1]/P0001  & ~n4070 ;
  assign n13284 = ~n3763 & n11121 ;
  assign n13285 = ~n3762 & n13284 ;
  assign n13286 = ~n3763 & n11110 ;
  assign n13287 = ~n3762 & n13286 ;
  assign n13288 = ~n3763 & n11136 ;
  assign n13289 = ~n3762 & n13288 ;
  assign n13290 = n2266 & n13271 ;
  assign n13291 = n2266 & n13269 ;
  assign n13292 = ~n3763 & n11146 ;
  assign n13293 = ~n3762 & n13292 ;
  assign n13294 = \ctl_rf_be_d1_reg[3]/P0001  & ~n4105 ;
  assign n13295 = ~n3763 & n11131 ;
  assign n13296 = ~n3762 & n13295 ;
  assign n13297 = ~n3763 & n11141 ;
  assign n13298 = ~n3762 & n13297 ;
  assign n13299 = \ctl_rf_be_d1_reg[1]/P0001  & ~n3766 ;
  assign n13300 = \ctl_rf_be_d1_reg[3]/P0001  & ~n3766 ;
  assign n13301 = \ctl_rf_be_d1_reg[1]/P0001  & ~n4088 ;
  assign n13302 = \ctl_rf_be_d1_reg[3]/P0001  & ~n4088 ;
  assign n13303 = \ctl_rf_be_d1_reg[3]/P0001  & ~n4139 ;
  assign n13304 = \ctl_rf_be_d1_reg[3]/P0001  & ~n4173 ;
  assign n13305 = \ctl_rf_be_d1_reg[1]/P0001  & ~n4122 ;
  assign n13306 = \ctl_rf_be_d1_reg[1]/P0001  & ~n4139 ;
  assign n13307 = \ctl_rf_be_d1_reg[1]/P0001  & ~n4156 ;
  assign n13308 = \ctl_rf_be_d1_reg[3]/P0001  & ~n4156 ;
  assign n13309 = ~\ctl_rf_c6_rf_int_tc1_msk_reg/NET0131  & \ctl_rf_tc_reg[6]/NET0131  ;
  assign n13310 = ~n4722 & ~n13309 ;
  assign n13311 = ~n6440 & ~n7828 ;
  assign n13312 = n13310 & n13311 ;
  assign n13313 = ~n5661 & ~n6116 ;
  assign n13314 = ~n6743 & ~n7046 ;
  assign n13315 = n13313 & n13314 ;
  assign n13316 = n13312 & n13315 ;
  assign n13317 = ~n6746 & ~n7049 ;
  assign n13318 = ~n7512 & ~n7831 ;
  assign n13319 = n13317 & n13318 ;
  assign n13320 = ~n4732 & ~n5662 ;
  assign n13321 = ~n6117 & ~n6443 ;
  assign n13322 = n13320 & n13321 ;
  assign n13323 = n13319 & n13322 ;
  assign n13324 = n13316 & n13323 ;
  assign n13325 = \ctl_rf_be_d1_reg[3]/P0001  & ~n4122 ;
  assign n13326 = \ctl_rf_be_d1_reg[1]/P0001  & ~n4173 ;
  assign n13327 = \ahb_slv_slv_ad_d1o_reg[2]/NET0131  & n11447 ;
  assign n13328 = n13271 & n13327 ;
  assign n13329 = n2234 & n11508 ;
  assign n13330 = n11447 & n13329 ;
  assign n13331 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[20]_pad  ;
  assign n13332 = n2238 & n13331 ;
  assign n13333 = ~n12024 & n13332 ;
  assign n13334 = n12025 & ~n13333 ;
  assign n13335 = \hwdata[4]_pad  & ~n12027 ;
  assign n13336 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[28]_pad  ;
  assign n13337 = n2241 & n13336 ;
  assign n13338 = ~n12024 & n13337 ;
  assign n13339 = ~n13333 & ~n13338 ;
  assign n13340 = ~n13335 & n13339 ;
  assign n13341 = ~n13334 & ~n13340 ;
  assign n13342 = ~\de_m0_arb_st_reg/NET0131  & n13341 ;
  assign n13343 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[16]_pad  ;
  assign n13344 = n2238 & n13343 ;
  assign n13345 = ~n12024 & n13344 ;
  assign n13346 = n12025 & ~n13345 ;
  assign n13347 = \hwdata[0]_pad  & ~n12027 ;
  assign n13348 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[24]_pad  ;
  assign n13349 = n2241 & n13348 ;
  assign n13350 = ~n12024 & n13349 ;
  assign n13351 = ~n13345 & ~n13350 ;
  assign n13352 = ~n13347 & n13351 ;
  assign n13353 = ~n13346 & ~n13352 ;
  assign n13354 = ~\de_m0_arb_st_reg/NET0131  & n13353 ;
  assign n13355 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[3]_pad  ;
  assign n13356 = n2238 & n13355 ;
  assign n13357 = ~n12024 & n13356 ;
  assign n13358 = n12025 & ~n13357 ;
  assign n13359 = \hwdata[19]_pad  & ~n12027 ;
  assign n13360 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[11]_pad  ;
  assign n13361 = n2241 & n13360 ;
  assign n13362 = ~n12024 & n13361 ;
  assign n13363 = ~n13357 & ~n13362 ;
  assign n13364 = ~n13359 & n13363 ;
  assign n13365 = ~n13358 & ~n13364 ;
  assign n13366 = ~\de_m0_arb_st_reg/NET0131  & n13365 ;
  assign n13367 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[7]_pad  ;
  assign n13368 = n2238 & n13367 ;
  assign n13369 = ~n12024 & n13368 ;
  assign n13370 = n12025 & ~n13369 ;
  assign n13371 = \hwdata[23]_pad  & ~n12027 ;
  assign n13372 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[15]_pad  ;
  assign n13373 = n2241 & n13372 ;
  assign n13374 = ~n12024 & n13373 ;
  assign n13375 = ~n13369 & ~n13374 ;
  assign n13376 = ~n13371 & n13375 ;
  assign n13377 = ~n13370 & ~n13376 ;
  assign n13378 = ~\de_m0_arb_st_reg/NET0131  & n13377 ;
  assign n13379 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[26]_pad  ;
  assign n13380 = n2238 & n13379 ;
  assign n13381 = ~n12024 & n13380 ;
  assign n13382 = n12025 & ~n13381 ;
  assign n13383 = \hwdata[10]_pad  & ~n12027 ;
  assign n13384 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[18]_pad  ;
  assign n13385 = n2241 & n13384 ;
  assign n13386 = ~n12024 & n13385 ;
  assign n13387 = ~n13381 & ~n13386 ;
  assign n13388 = ~n13383 & n13387 ;
  assign n13389 = ~n13382 & ~n13388 ;
  assign n13390 = ~\de_m0_arb_st_reg/NET0131  & n13389 ;
  assign n13391 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[27]_pad  ;
  assign n13392 = n2238 & n13391 ;
  assign n13393 = ~n12024 & n13392 ;
  assign n13394 = n12025 & ~n13393 ;
  assign n13395 = \hwdata[11]_pad  & ~n12027 ;
  assign n13396 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[19]_pad  ;
  assign n13397 = n2241 & n13396 ;
  assign n13398 = ~n12024 & n13397 ;
  assign n13399 = ~n13393 & ~n13398 ;
  assign n13400 = ~n13395 & n13399 ;
  assign n13401 = ~n13394 & ~n13400 ;
  assign n13402 = ~\de_m0_arb_st_reg/NET0131  & n13401 ;
  assign n13403 = n2238 & n13336 ;
  assign n13404 = ~n12024 & n13403 ;
  assign n13405 = n12025 & ~n13404 ;
  assign n13406 = \hwdata[12]_pad  & ~n12027 ;
  assign n13407 = n2241 & n13331 ;
  assign n13408 = ~n12024 & n13407 ;
  assign n13409 = ~n13404 & ~n13408 ;
  assign n13410 = ~n13406 & n13409 ;
  assign n13411 = ~n13405 & ~n13410 ;
  assign n13412 = ~\de_m0_arb_st_reg/NET0131  & n13411 ;
  assign n13413 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[29]_pad  ;
  assign n13414 = n2238 & n13413 ;
  assign n13415 = ~n12024 & n13414 ;
  assign n13416 = n12025 & ~n13415 ;
  assign n13417 = \hwdata[13]_pad  & ~n12027 ;
  assign n13418 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[21]_pad  ;
  assign n13419 = n2241 & n13418 ;
  assign n13420 = ~n12024 & n13419 ;
  assign n13421 = ~n13415 & ~n13420 ;
  assign n13422 = ~n13417 & n13421 ;
  assign n13423 = ~n13416 & ~n13422 ;
  assign n13424 = ~\de_m0_arb_st_reg/NET0131  & n13423 ;
  assign n13425 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[30]_pad  ;
  assign n13426 = n2238 & n13425 ;
  assign n13427 = ~n12024 & n13426 ;
  assign n13428 = n12025 & ~n13427 ;
  assign n13429 = \hwdata[14]_pad  & ~n12027 ;
  assign n13430 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[22]_pad  ;
  assign n13431 = n2241 & n13430 ;
  assign n13432 = ~n12024 & n13431 ;
  assign n13433 = ~n13427 & ~n13432 ;
  assign n13434 = ~n13429 & n13433 ;
  assign n13435 = ~n13428 & ~n13434 ;
  assign n13436 = ~\de_m0_arb_st_reg/NET0131  & n13435 ;
  assign n13437 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[10]_pad  ;
  assign n13438 = n2238 & n13437 ;
  assign n13439 = ~n12024 & n13438 ;
  assign n13440 = n12025 & ~n13439 ;
  assign n13441 = \hwdata[26]_pad  & ~n12027 ;
  assign n13442 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[2]_pad  ;
  assign n13443 = n2241 & n13442 ;
  assign n13444 = ~n12024 & n13443 ;
  assign n13445 = ~n13439 & ~n13444 ;
  assign n13446 = ~n13441 & n13445 ;
  assign n13447 = ~n13440 & ~n13446 ;
  assign n13448 = ~\de_m0_arb_st_reg/NET0131  & n13447 ;
  assign n13449 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[31]_pad  ;
  assign n13450 = n2238 & n13449 ;
  assign n13451 = ~n12024 & n13450 ;
  assign n13452 = n12025 & ~n13451 ;
  assign n13453 = \hwdata[15]_pad  & ~n12027 ;
  assign n13454 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[23]_pad  ;
  assign n13455 = n2241 & n13454 ;
  assign n13456 = ~n12024 & n13455 ;
  assign n13457 = ~n13451 & ~n13456 ;
  assign n13458 = ~n13453 & n13457 ;
  assign n13459 = ~n13452 & ~n13458 ;
  assign n13460 = ~\de_m0_arb_st_reg/NET0131  & n13459 ;
  assign n13461 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[0]_pad  ;
  assign n13462 = n2238 & n13461 ;
  assign n13463 = ~n12024 & n13462 ;
  assign n13464 = n12025 & ~n13463 ;
  assign n13465 = \hwdata[16]_pad  & ~n12027 ;
  assign n13466 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[8]_pad  ;
  assign n13467 = n2241 & n13466 ;
  assign n13468 = ~n12024 & n13467 ;
  assign n13469 = ~n13463 & ~n13468 ;
  assign n13470 = ~n13465 & n13469 ;
  assign n13471 = ~n13464 & ~n13470 ;
  assign n13472 = ~\de_m0_arb_st_reg/NET0131  & n13471 ;
  assign n13473 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[1]_pad  ;
  assign n13474 = n2238 & n13473 ;
  assign n13475 = ~n12024 & n13474 ;
  assign n13476 = n12025 & ~n13475 ;
  assign n13477 = \hwdata[17]_pad  & ~n12027 ;
  assign n13478 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[9]_pad  ;
  assign n13479 = n2241 & n13478 ;
  assign n13480 = ~n12024 & n13479 ;
  assign n13481 = ~n13475 & ~n13480 ;
  assign n13482 = ~n13477 & n13481 ;
  assign n13483 = ~n13476 & ~n13482 ;
  assign n13484 = ~\de_m0_arb_st_reg/NET0131  & n13483 ;
  assign n13485 = n2238 & n13442 ;
  assign n13486 = ~n12024 & n13485 ;
  assign n13487 = n12025 & ~n13486 ;
  assign n13488 = \hwdata[18]_pad  & ~n12027 ;
  assign n13489 = n2241 & n13437 ;
  assign n13490 = ~n12024 & n13489 ;
  assign n13491 = ~n13486 & ~n13490 ;
  assign n13492 = ~n13488 & n13491 ;
  assign n13493 = ~n13487 & ~n13492 ;
  assign n13494 = ~\de_m0_arb_st_reg/NET0131  & n13493 ;
  assign n13495 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[17]_pad  ;
  assign n13496 = n2238 & n13495 ;
  assign n13497 = ~n12024 & n13496 ;
  assign n13498 = n12025 & ~n13497 ;
  assign n13499 = \hwdata[1]_pad  & ~n12027 ;
  assign n13500 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[25]_pad  ;
  assign n13501 = n2241 & n13500 ;
  assign n13502 = ~n12024 & n13501 ;
  assign n13503 = ~n13497 & ~n13502 ;
  assign n13504 = ~n13499 & n13503 ;
  assign n13505 = ~n13498 & ~n13504 ;
  assign n13506 = ~\de_m0_arb_st_reg/NET0131  & n13505 ;
  assign n13507 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[4]_pad  ;
  assign n13508 = n2238 & n13507 ;
  assign n13509 = ~n12024 & n13508 ;
  assign n13510 = n12025 & ~n13509 ;
  assign n13511 = \hwdata[20]_pad  & ~n12027 ;
  assign n13512 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[12]_pad  ;
  assign n13513 = n2241 & n13512 ;
  assign n13514 = ~n12024 & n13513 ;
  assign n13515 = ~n13509 & ~n13514 ;
  assign n13516 = ~n13511 & n13515 ;
  assign n13517 = ~n13510 & ~n13516 ;
  assign n13518 = ~\de_m0_arb_st_reg/NET0131  & n13517 ;
  assign n13519 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[5]_pad  ;
  assign n13520 = n2238 & n13519 ;
  assign n13521 = ~n12024 & n13520 ;
  assign n13522 = n12025 & ~n13521 ;
  assign n13523 = \hwdata[21]_pad  & ~n12027 ;
  assign n13524 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[13]_pad  ;
  assign n13525 = n2241 & n13524 ;
  assign n13526 = ~n12024 & n13525 ;
  assign n13527 = ~n13521 & ~n13526 ;
  assign n13528 = ~n13523 & n13527 ;
  assign n13529 = ~n13522 & ~n13528 ;
  assign n13530 = ~\de_m0_arb_st_reg/NET0131  & n13529 ;
  assign n13531 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[6]_pad  ;
  assign n13532 = n2238 & n13531 ;
  assign n13533 = ~n12024 & n13532 ;
  assign n13534 = n12025 & ~n13533 ;
  assign n13535 = \hwdata[22]_pad  & ~n12027 ;
  assign n13536 = ~\ahb_slv_slv_sz_d1o_reg[2]/NET0131  & \hwdata[14]_pad  ;
  assign n13537 = n2241 & n13536 ;
  assign n13538 = ~n12024 & n13537 ;
  assign n13539 = ~n13533 & ~n13538 ;
  assign n13540 = ~n13535 & n13539 ;
  assign n13541 = ~n13534 & ~n13540 ;
  assign n13542 = ~\de_m0_arb_st_reg/NET0131  & n13541 ;
  assign n13543 = n2238 & n13466 ;
  assign n13544 = ~n12024 & n13543 ;
  assign n13545 = n12025 & ~n13544 ;
  assign n13546 = \hwdata[24]_pad  & ~n12027 ;
  assign n13547 = n2241 & n13461 ;
  assign n13548 = ~n12024 & n13547 ;
  assign n13549 = ~n13544 & ~n13548 ;
  assign n13550 = ~n13546 & n13549 ;
  assign n13551 = ~n13545 & ~n13550 ;
  assign n13552 = ~\de_m0_arb_st_reg/NET0131  & n13551 ;
  assign n13553 = n2238 & n13360 ;
  assign n13554 = ~n12024 & n13553 ;
  assign n13555 = n12025 & ~n13554 ;
  assign n13556 = \hwdata[27]_pad  & ~n12027 ;
  assign n13557 = n2241 & n13355 ;
  assign n13558 = ~n12024 & n13557 ;
  assign n13559 = ~n13554 & ~n13558 ;
  assign n13560 = ~n13556 & n13559 ;
  assign n13561 = ~n13555 & ~n13560 ;
  assign n13562 = ~\de_m0_arb_st_reg/NET0131  & n13561 ;
  assign n13563 = n2238 & n13512 ;
  assign n13564 = ~n12024 & n13563 ;
  assign n13565 = n12025 & ~n13564 ;
  assign n13566 = \hwdata[28]_pad  & ~n12027 ;
  assign n13567 = n2241 & n13507 ;
  assign n13568 = ~n12024 & n13567 ;
  assign n13569 = ~n13564 & ~n13568 ;
  assign n13570 = ~n13566 & n13569 ;
  assign n13571 = ~n13565 & ~n13570 ;
  assign n13572 = ~\de_m0_arb_st_reg/NET0131  & n13571 ;
  assign n13573 = n2238 & n13384 ;
  assign n13574 = ~n12024 & n13573 ;
  assign n13575 = n12025 & ~n13574 ;
  assign n13576 = \hwdata[2]_pad  & ~n12027 ;
  assign n13577 = n2241 & n13379 ;
  assign n13578 = ~n12024 & n13577 ;
  assign n13579 = ~n13574 & ~n13578 ;
  assign n13580 = ~n13576 & n13579 ;
  assign n13581 = ~n13575 & ~n13580 ;
  assign n13582 = ~\de_m0_arb_st_reg/NET0131  & n13581 ;
  assign n13583 = n2238 & n13536 ;
  assign n13584 = ~n12024 & n13583 ;
  assign n13585 = n12025 & ~n13584 ;
  assign n13586 = \hwdata[30]_pad  & ~n12027 ;
  assign n13587 = n2241 & n13531 ;
  assign n13588 = ~n12024 & n13587 ;
  assign n13589 = ~n13584 & ~n13588 ;
  assign n13590 = ~n13586 & n13589 ;
  assign n13591 = ~n13585 & ~n13590 ;
  assign n13592 = ~\de_m0_arb_st_reg/NET0131  & n13591 ;
  assign n13593 = n2238 & n13372 ;
  assign n13594 = ~n12024 & n13593 ;
  assign n13595 = n12025 & ~n13594 ;
  assign n13596 = \hwdata[31]_pad  & ~n12027 ;
  assign n13597 = n2241 & n13367 ;
  assign n13598 = ~n12024 & n13597 ;
  assign n13599 = ~n13594 & ~n13598 ;
  assign n13600 = ~n13596 & n13599 ;
  assign n13601 = ~n13595 & ~n13600 ;
  assign n13602 = ~\de_m0_arb_st_reg/NET0131  & n13601 ;
  assign n13603 = n2238 & n13418 ;
  assign n13604 = ~n12024 & n13603 ;
  assign n13605 = n12025 & ~n13604 ;
  assign n13606 = \hwdata[5]_pad  & ~n12027 ;
  assign n13607 = n2241 & n13413 ;
  assign n13608 = ~n12024 & n13607 ;
  assign n13609 = ~n13604 & ~n13608 ;
  assign n13610 = ~n13606 & n13609 ;
  assign n13611 = ~n13605 & ~n13610 ;
  assign n13612 = ~\de_m0_arb_st_reg/NET0131  & n13611 ;
  assign n13613 = n2238 & n13430 ;
  assign n13614 = ~n12024 & n13613 ;
  assign n13615 = n12025 & ~n13614 ;
  assign n13616 = \hwdata[6]_pad  & ~n12027 ;
  assign n13617 = n2241 & n13425 ;
  assign n13618 = ~n12024 & n13617 ;
  assign n13619 = ~n13614 & ~n13618 ;
  assign n13620 = ~n13616 & n13619 ;
  assign n13621 = ~n13615 & ~n13620 ;
  assign n13622 = ~\de_m0_arb_st_reg/NET0131  & n13621 ;
  assign n13623 = n2238 & n13454 ;
  assign n13624 = ~n12024 & n13623 ;
  assign n13625 = n12025 & ~n13624 ;
  assign n13626 = \hwdata[7]_pad  & ~n12027 ;
  assign n13627 = n2241 & n13449 ;
  assign n13628 = ~n12024 & n13627 ;
  assign n13629 = ~n13624 & ~n13628 ;
  assign n13630 = ~n13626 & n13629 ;
  assign n13631 = ~n13625 & ~n13630 ;
  assign n13632 = ~\de_m0_arb_st_reg/NET0131  & n13631 ;
  assign n13633 = n2238 & n13348 ;
  assign n13634 = ~n12024 & n13633 ;
  assign n13635 = n12025 & ~n13634 ;
  assign n13636 = \hwdata[8]_pad  & ~n12027 ;
  assign n13637 = n2241 & n13343 ;
  assign n13638 = ~n12024 & n13637 ;
  assign n13639 = ~n13634 & ~n13638 ;
  assign n13640 = ~n13636 & n13639 ;
  assign n13641 = ~n13635 & ~n13640 ;
  assign n13642 = ~\de_m0_arb_st_reg/NET0131  & n13641 ;
  assign n13643 = n2238 & n13500 ;
  assign n13644 = ~n12024 & n13643 ;
  assign n13645 = n12025 & ~n13644 ;
  assign n13646 = \hwdata[9]_pad  & ~n12027 ;
  assign n13647 = n2241 & n13495 ;
  assign n13648 = ~n12024 & n13647 ;
  assign n13649 = ~n13644 & ~n13648 ;
  assign n13650 = ~n13646 & n13649 ;
  assign n13651 = ~n13645 & ~n13650 ;
  assign n13652 = ~\de_m0_arb_st_reg/NET0131  & n13651 ;
  assign n13653 = n2238 & n13478 ;
  assign n13654 = ~n12024 & n13653 ;
  assign n13655 = n12025 & ~n13654 ;
  assign n13656 = \hwdata[25]_pad  & ~n12027 ;
  assign n13657 = n2241 & n13473 ;
  assign n13658 = ~n12024 & n13657 ;
  assign n13659 = ~n13654 & ~n13658 ;
  assign n13660 = ~n13656 & n13659 ;
  assign n13661 = ~n13655 & ~n13660 ;
  assign n13662 = ~\de_m0_arb_st_reg/NET0131  & n13661 ;
  assign n13663 = n2238 & n13524 ;
  assign n13664 = ~n12024 & n13663 ;
  assign n13665 = n12025 & ~n13664 ;
  assign n13666 = \hwdata[29]_pad  & ~n12027 ;
  assign n13667 = n2241 & n13519 ;
  assign n13668 = ~n12024 & n13667 ;
  assign n13669 = ~n13664 & ~n13668 ;
  assign n13670 = ~n13666 & n13669 ;
  assign n13671 = ~n13665 & ~n13670 ;
  assign n13672 = ~\de_m0_arb_st_reg/NET0131  & n13671 ;
  assign n13673 = n2238 & n13396 ;
  assign n13674 = ~n12024 & n13673 ;
  assign n13675 = n12025 & ~n13674 ;
  assign n13676 = \hwdata[3]_pad  & ~n12027 ;
  assign n13677 = n2241 & n13391 ;
  assign n13678 = ~n12024 & n13677 ;
  assign n13679 = ~n13674 & ~n13678 ;
  assign n13680 = ~n13676 & n13679 ;
  assign n13681 = ~n13675 & ~n13680 ;
  assign n13682 = ~\de_m0_arb_st_reg/NET0131  & n13681 ;
  assign n13683 = ~\ahb_slv_slv_ad_d1o_reg[8]/NET0131  & n2275 ;
  assign n13684 = ~\ahb_slv_slv_ad_d1o_reg[2]/NET0131  & \ahb_slv_slv_wr_d1o_reg/NET0131  ;
  assign n13685 = n2272 & n13684 ;
  assign n13686 = n13683 & n13685 ;
  assign n13687 = \ctl_rf_be_d1_reg[2]/P0001  & n3755 ;
  assign n13688 = n13686 & n13687 ;
  assign n13689 = \ahb_slv_slv_ad_d1o_reg[4]/NET0131  & \ahb_slv_slv_wr_d1o_reg/NET0131  ;
  assign n13690 = n2272 & n13689 ;
  assign n13691 = n13683 & n13690 ;
  assign n13692 = \ahb_slv_slv_ad_d1o_reg[2]/NET0131  & ~\ahb_slv_slv_ad_d1o_reg[3]/NET0131  ;
  assign n13693 = \ctl_rf_be_d1_reg[2]/P0001  & n13692 ;
  assign n13694 = n13691 & n13693 ;
  assign n13695 = ~\ahb_slv_slv_ad_d1o_reg[4]/NET0131  & \ahb_slv_slv_wr_d1o_reg/NET0131  ;
  assign n13696 = n2272 & n13695 ;
  assign n13697 = n13683 & n13696 ;
  assign n13698 = \ahb_slv_slv_ad_d1o_reg[2]/NET0131  & \ahb_slv_slv_ad_d1o_reg[3]/NET0131  ;
  assign n13699 = \ctl_rf_be_d1_reg[2]/P0001  & n13698 ;
  assign n13700 = n13697 & n13699 ;
  assign n13701 = \ctl_rf_be_d1_reg[3]/P0001  & n13698 ;
  assign n13702 = n13697 & n13701 ;
  assign n13703 = ~\ahb_slv_slv_ad_d1o_reg[2]/NET0131  & ~\ahb_slv_slv_ad_d1o_reg[7]/NET0131  ;
  assign n13704 = n2264 & n13703 ;
  assign n13705 = n13683 & n13704 ;
  assign n13706 = n11449 & n13705 ;
  assign n13707 = \ctl_rf_be_d1_reg[3]/P0001  & n8577 ;
  assign n13708 = n13705 & n13707 ;
  assign n13709 = \ctl_rf_be_d1_reg[3]/P0001  & n3755 ;
  assign n13710 = n13686 & n13709 ;
  assign n13711 = \ctl_rf_be_d1_reg[3]/P0001  & n13692 ;
  assign n13712 = n13691 & n13711 ;
  assign n13713 = ~n2922 & n13353 ;
  assign n13714 = ~n2922 & n13671 ;
  assign n13715 = ~n2922 & n13581 ;
  assign n13716 = ~n2922 & n13601 ;
  assign n13717 = ~n2922 & n13483 ;
  assign n13718 = ~n2922 & n13661 ;
  assign n13719 = ~n2922 & n13681 ;
  assign n13720 = ~n2922 & n13459 ;
  assign n13721 = ~n2922 & n13591 ;
  assign n13722 = ~n2922 & n13571 ;
  assign n13723 = ~n2922 & n13611 ;
  assign n13724 = ~n2922 & n13423 ;
  assign n13725 = ~n2922 & n13631 ;
  assign n13726 = ~n2922 & n13621 ;
  assign n13727 = ~n2922 & n13641 ;
  assign n13728 = ~n2922 & n13389 ;
  assign n13729 = ~n2922 & n13471 ;
  assign n13730 = ~n2922 & n13561 ;
  assign n13731 = ~n2922 & n13365 ;
  assign n13732 = ~n2922 & n13411 ;
  assign n13733 = ~n2922 & n13493 ;
  assign n13734 = ~n2922 & n13377 ;
  assign n13735 = ~n2922 & n13529 ;
  assign n13736 = ~n2922 & n13447 ;
  assign n13737 = ~n2922 & n13401 ;
  assign n13738 = ~n2922 & n13435 ;
  assign n13739 = ~n2922 & n13505 ;
  assign n13740 = ~n2922 & n13517 ;
  assign n13741 = ~n2922 & n13541 ;
  assign n13742 = ~n2922 & n13551 ;
  assign n13743 = ~n2922 & n13341 ;
  assign n13744 = ~n2922 & n13651 ;
  assign n13745 = n2252 & n2318 ;
  assign n13746 = n11449 & n13686 ;
  assign n13747 = \ctl_rf_be_d1_reg[1]/P0001  & n8630 ;
  assign n13748 = n8578 & n13747 ;
  assign n13749 = n13687 & n13705 ;
  assign n13750 = n13705 & n13709 ;
  assign n13751 = n2252 & n2300 ;
  assign n13752 = n13697 & n13711 ;
  assign n13753 = \ahb_slv_slv_ad_d1o_reg[2]/NET0131  & ~\ahb_slv_slv_ad_d1o_reg[7]/NET0131  ;
  assign n13754 = n2264 & n13753 ;
  assign n13755 = n13683 & n13754 ;
  assign n13756 = n13707 & n13755 ;
  assign n13757 = n2266 & n2318 ;
  assign n13758 = \ahb_slv_slv_ad_d1o_reg[3]/NET0131  & \ahb_slv_slv_ad_d1o_reg[4]/NET0131  ;
  assign n13759 = \ctl_rf_be_d1_reg[3]/P0001  & n13758 ;
  assign n13760 = n13705 & n13759 ;
  assign n13761 = n13755 & n13759 ;
  assign n13762 = n8609 & n13747 ;
  assign n13763 = \ctl_rf_be_d1_reg[2]/P0001  & n2233 ;
  assign n13764 = n13686 & n13763 ;
  assign n13765 = \ctl_rf_be_d1_reg[3]/P0001  & n2233 ;
  assign n13766 = n13686 & n13765 ;
  assign n13767 = n13705 & n13763 ;
  assign n13768 = n2266 & n2300 ;
  assign n13769 = n13755 & n13763 ;
  assign n13770 = n13755 & n13765 ;
  assign n13771 = n8629 & n13747 ;
  assign n13772 = n2274 & n2300 ;
  assign n13773 = n13705 & n13765 ;
  assign n13774 = \ctl_rf_be_d1_reg[1]/P0001  & n8579 ;
  assign n13775 = n8629 & n13774 ;
  assign n13776 = n13693 & n13697 ;
  assign n13777 = n11449 & n13755 ;
  assign n13778 = \ctl_rf_be_d1_reg[1]/P0001  & n8657 ;
  assign n13779 = n8656 & n13778 ;
  assign n13780 = \ctl_rf_be_d1_reg[2]/P0001  & n13758 ;
  assign n13781 = n13686 & n13780 ;
  assign n13782 = n13686 & n13759 ;
  assign n13783 = n13705 & n13780 ;
  assign n13784 = n2289 & n2300 ;
  assign n13785 = n8677 & n13778 ;
  assign n13786 = n13686 & n13707 ;
  assign n13787 = n13687 & n13755 ;
  assign n13788 = n13755 & n13780 ;
  assign n13789 = n13691 & n13701 ;
  assign n13790 = n13691 & n13699 ;
  assign n13791 = n13709 & n13755 ;
  assign n13792 = ~\ctl_rf_c0_rf_chllp_on_reg/NET0131  & n4018 ;
  assign n13793 = \ctl_rf_c0_rf_ch_en_reg/NET0131  & ~n13792 ;
  assign n13794 = ~\ctl_rf_c1_rf_chllp_on_reg/NET0131  & n3891 ;
  assign n13795 = \ctl_rf_c1_rf_ch_en_reg/NET0131  & ~n13794 ;
  assign n13796 = n8578 & n13774 ;
  assign n13797 = ~\ctl_rf_c2_rf_chllp_on_reg/NET0131  & n3828 ;
  assign n13798 = \ctl_rf_c2_rf_ch_en_reg/NET0131  & ~n13797 ;
  assign n13799 = ~\ctl_rf_c3_rf_chllp_on_reg/NET0131  & n3922 ;
  assign n13800 = \ctl_rf_c3_rf_ch_en_reg/NET0131  & ~n13799 ;
  assign n13801 = n8609 & n13774 ;
  assign n13802 = n2274 & n2318 ;
  assign n13803 = ~\ctl_rf_c4_rf_chllp_on_reg/NET0131  & n3859 ;
  assign n13804 = \ctl_rf_c4_rf_ch_en_reg/NET0131  & ~n13803 ;
  assign n13805 = ~\ctl_rf_c5_rf_chllp_on_reg/NET0131  & n3986 ;
  assign n13806 = \ctl_rf_c5_rf_ch_en_reg/NET0131  & ~n13805 ;
  assign n13807 = n2289 & n2318 ;
  assign n13808 = ~\ctl_rf_c6_rf_chllp_on_reg/NET0131  & n4049 ;
  assign n13809 = \ctl_rf_c6_rf_ch_en_reg/NET0131  & ~n13808 ;
  assign n13810 = ~\ctl_rf_c7_rf_chllp_on_reg/NET0131  & n3955 ;
  assign n13811 = \ctl_rf_c7_rf_ch_en_reg/NET0131  & ~n13810 ;
  assign n13812 = ~n2940 & ~n4539 ;
  assign n13813 = \h0readyin_pad  & ~n13812 ;
  assign n13814 = \h0write_pad  & ~n13813 ;
  assign n13815 = \ch_sel_arb_chcsr_reg_reg[2]/NET0131  & \h0readyin_pad  ;
  assign n13816 = n11003 & n13815 ;
  assign n13817 = ~n13814 & ~n13816 ;
  assign n13818 = ~n8991 & ~n8992 ;
  assign n13819 = ~n2574 & ~n2575 ;
  assign n13820 = ~n9788 & ~n9789 ;
  assign n13821 = ~n9797 & ~n9798 ;
  assign n13822 = ~n9806 & ~n9807 ;
  assign n13823 = ~n9815 & ~n9816 ;
  assign n13824 = ~n10580 & ~n10581 ;
  assign n13825 = ~n9000 & ~n9001 ;
  assign n13826 = ~n10593 & ~n10594 ;
  assign n13827 = ~n2306 & ~n2307 ;
  assign n13828 = ~n9043 & ~n9044 ;
  assign n13829 = ~n8713 & ~n8714 ;
  assign n13830 = ~n8586 & ~n8587 ;
  assign n13831 = ~n8595 & ~n8596 ;
  assign n13832 = ~n2246 & ~n2247 ;
  assign n13833 = ~n8780 & ~n8781 ;
  assign n13834 = ~n8807 & ~n8808 ;
  assign n13835 = ~n2679 & ~n2680 ;
  assign n13836 = ~n8767 & ~n8768 ;
  assign n13837 = ~n2259 & ~n2260 ;
  assign n13838 = ~n2399 & ~n2400 ;
  assign n13839 = ~n2408 & ~n2409 ;
  assign n13840 = ~n2565 & ~n2566 ;
  assign n13841 = ~n2365 & ~n2366 ;
  assign n13842 = ~n2499 & ~n2500 ;
  assign n13843 = ~n2528 & ~n2529 ;
  assign n13844 = ~n9026 & ~n9027 ;
  assign n13845 = ~n8758 & ~n8759 ;
  assign n13846 = ~n8790 & ~n8791 ;
  assign n13847 = ~n9017 & ~n9018 ;
  assign n13848 = ~\ahb_slv_slv_ad_d1o_reg[4]/NET0131  & ~\haddr[4]_pad  ;
  assign n13849 = \ahb_slv_slv_ad_d1o_reg[4]/NET0131  & \haddr[4]_pad  ;
  assign n13850 = ~n13848 & ~n13849 ;
  assign n13851 = ~\ahb_slv_slv_ad_d1o_reg[8]/NET0131  & ~\haddr[8]_pad  ;
  assign n13852 = \ahb_slv_slv_ad_d1o_reg[8]/NET0131  & \haddr[8]_pad  ;
  assign n13853 = ~n13851 & ~n13852 ;
  assign n13854 = hreadyin_pad & n4569 ;
  assign n13855 = ~n13853 & n13854 ;
  assign n13856 = ~n13850 & n13855 ;
  assign n13857 = \ahb_slv_slv_ad_d1o_reg[7]/NET0131  & ~\haddr[7]_pad  ;
  assign n13858 = ~\ahb_slv_slv_ad_d1o_reg[3]/NET0131  & \haddr[3]_pad  ;
  assign n13859 = ~\ahb_slv_slv_ad_d1o_reg[5]/NET0131  & \haddr[5]_pad  ;
  assign n13860 = ~n13858 & ~n13859 ;
  assign n13861 = ~n13857 & n13860 ;
  assign n13862 = ~\ahb_slv_slv_ad_d1o_reg[7]/NET0131  & \haddr[7]_pad  ;
  assign n13863 = \ahb_slv_slv_ad_d1o_reg[5]/NET0131  & ~\haddr[5]_pad  ;
  assign n13864 = ~n13862 & ~n13863 ;
  assign n13865 = \ahb_slv_slv_ad_d1o_reg[6]/NET0131  & ~\haddr[6]_pad  ;
  assign n13866 = \ahb_slv_slv_ad_d1o_reg[2]/NET0131  & ~\haddr[2]_pad  ;
  assign n13867 = ~n13865 & ~n13866 ;
  assign n13868 = n13864 & n13867 ;
  assign n13869 = ~\ahb_slv_slv_ad_d1o_reg[2]/NET0131  & \haddr[2]_pad  ;
  assign n13870 = hwrite_pad & ~n13869 ;
  assign n13871 = ~\ahb_slv_slv_ad_d1o_reg[6]/NET0131  & \haddr[6]_pad  ;
  assign n13872 = \ahb_slv_slv_ad_d1o_reg[3]/NET0131  & ~\haddr[3]_pad  ;
  assign n13873 = ~n13871 & ~n13872 ;
  assign n13874 = n13870 & n13873 ;
  assign n13875 = n13868 & n13874 ;
  assign n13876 = n13861 & n13875 ;
  assign n13877 = n13856 & n13876 ;
  assign n13878 = ~\de_de_st_reg[5]/NET0131  & \de_m0_arb_st_reg/NET0131  ;
  assign n13879 = ~\ch_sel_arb_chcsr_reg_reg[1]/NET0131  & n11086 ;
  assign n13880 = ~n13878 & ~n13879 ;
  assign n13881 = ~\hsize[0]_pad  & \hsize[1]_pad  ;
  assign n13882 = ~\hsize[2]_pad  & n13881 ;
  assign n13883 = ~\haddr[1]_pad  & \hsize[0]_pad  ;
  assign n13884 = n4571 & n13883 ;
  assign n13885 = ~n13882 & ~n13884 ;
  assign n13886 = ~\hsize[0]_pad  & n4571 ;
  assign n13887 = ~\haddr[0]_pad  & ~\haddr[1]_pad  ;
  assign n13888 = n13886 & n13887 ;
  assign n13889 = n13885 & ~n13888 ;
  assign n13890 = \haddr[0]_pad  & ~\haddr[1]_pad  ;
  assign n13891 = n13886 & n13890 ;
  assign n13892 = n13885 & ~n13891 ;
  assign n13893 = \haddr[1]_pad  & ~\hsize[0]_pad  ;
  assign n13894 = n4571 & n13893 ;
  assign n13895 = ~\haddr[0]_pad  & n13894 ;
  assign n13896 = \haddr[1]_pad  & \hsize[0]_pad  ;
  assign n13897 = n4571 & n13896 ;
  assign n13898 = ~n13882 & ~n13897 ;
  assign n13899 = ~n13895 & n13898 ;
  assign n13900 = \haddr[0]_pad  & n13894 ;
  assign n13901 = n13898 & ~n13900 ;
  assign n13902 = hreadyin_pad & \htrans[1]_pad  ;
  assign n13903 = ~hsel_br_pad & ~hsel_reg_pad ;
  assign n13904 = n13902 & ~n13903 ;
  assign n13905 = \ch_sel_dma_reqd1_reg[5]/NET0131  & \ctl_rf_sync_reg[5]/NET0131  ;
  assign n13906 = \ch_sel_dma_reqd1_reg[7]/NET0131  & \ctl_rf_sync_reg[7]/NET0131  ;
  assign n13907 = \ch_sel_dma_reqd1_reg[1]/NET0131  & \ctl_rf_sync_reg[1]/NET0131  ;
  assign n13908 = \ch_sel_dma_reqd1_reg[0]/NET0131  & \ctl_rf_sync_reg[0]/NET0131  ;
  assign n13909 = \ch_sel_dma_reqd1_reg[4]/NET0131  & \ctl_rf_sync_reg[4]/NET0131  ;
  assign n13910 = \ch_sel_dma_reqd1_reg[3]/NET0131  & \ctl_rf_sync_reg[3]/NET0131  ;
  assign n13911 = \ch_sel_dma_reqd1_reg[6]/NET0131  & \ctl_rf_sync_reg[6]/NET0131  ;
  assign n13912 = \ch_sel_dma_reqd1_reg[2]/NET0131  & \ctl_rf_sync_reg[2]/NET0131  ;
  assign n13913 = \ahb_mst0_mx_dtp_reg/NET0131  & ~\h0readyin_pad  ;
  assign n13914 = ~n4521 & ~n13913 ;
  assign n13915 = ~\de_de_st_reg[5]/NET0131  & ~\de_st_rd_msk_reg/NET0131  ;
  assign n13916 = ~n10794 & ~n13915 ;
  assign n13917 = ~\ctl_rf_c7_rf_chdad_reg[18]/NET0131  & ~n2295 ;
  assign n13918 = n2295 & ~n2400 ;
  assign n13919 = ~n2399 & n13918 ;
  assign n13920 = ~n13917 & ~n13919 ;
  assign n13921 = ~\ctl_rf_c7_rf_chdad_reg[19]/NET0131  & ~n2295 ;
  assign n13922 = n2295 & ~n2409 ;
  assign n13923 = ~n2408 & n13922 ;
  assign n13924 = ~n13921 & ~n13923 ;
  assign n13925 = ~\ctl_rf_c2_rf_chllp_reg[24]/NET0131  & ~n10484 ;
  assign n13926 = ~n2575 & n10484 ;
  assign n13927 = ~n2574 & n13926 ;
  assign n13928 = ~n13925 & ~n13927 ;
  assign n13929 = ~\ctl_rf_c1_rf_chsad_reg[18]/NET0131  & ~n2360 ;
  assign n13930 = n2360 & ~n2400 ;
  assign n13931 = ~n2399 & n13930 ;
  assign n13932 = ~n13929 & ~n13931 ;
  assign n13933 = ~\ctl_rf_c5_rf_chdad_reg[1]/NET0131  & ~n9302 ;
  assign n13934 = ~n8992 & n9302 ;
  assign n13935 = ~n8991 & n13934 ;
  assign n13936 = ~n13933 & ~n13935 ;
  assign n13937 = ~\ctl_rf_c5_rf_chtsz_reg[7]/NET0131  & ~n8646 ;
  assign n13938 = ~n2247 & n8646 ;
  assign n13939 = ~n2246 & n13938 ;
  assign n13940 = ~n13937 & ~n13939 ;
  assign n13941 = ~\ctl_rf_c5_rf_chtsz_reg[5]/NET0131  & ~n8646 ;
  assign n13942 = ~n8587 & n8646 ;
  assign n13943 = ~n8586 & n13942 ;
  assign n13944 = ~n13941 & ~n13943 ;
  assign n13945 = ~\ctl_rf_c5_rf_chtsz_reg[4]/NET0131  & ~n8646 ;
  assign n13946 = n8646 & ~n8714 ;
  assign n13947 = ~n8713 & n13946 ;
  assign n13948 = ~n13945 & ~n13947 ;
  assign n13949 = ~\ctl_rf_c6_rf_chsad_reg[17]/NET0131  & ~n2385 ;
  assign n13950 = ~n2260 & n2385 ;
  assign n13951 = ~n2259 & n13950 ;
  assign n13952 = ~n13949 & ~n13951 ;
  assign n13953 = ~\ctl_rf_c7_rf_chsad_reg[17]/NET0131  & ~n2390 ;
  assign n13954 = ~n2260 & n2390 ;
  assign n13955 = ~n2259 & n13954 ;
  assign n13956 = ~n13953 & ~n13955 ;
  assign n13957 = ~\ctl_rf_c3_rf_chsad_reg[17]/NET0131  & ~n2370 ;
  assign n13958 = ~n2260 & n2370 ;
  assign n13959 = ~n2259 & n13958 ;
  assign n13960 = ~n13957 & ~n13959 ;
  assign n13961 = ~\ctl_rf_c4_rf_chsad_reg[17]/NET0131  & ~n2375 ;
  assign n13962 = ~n2260 & n2375 ;
  assign n13963 = ~n2259 & n13962 ;
  assign n13964 = ~n13961 & ~n13963 ;
  assign n13965 = ~\ctl_rf_c5_rf_chsad_reg[17]/NET0131  & ~n2380 ;
  assign n13966 = ~n2260 & n2380 ;
  assign n13967 = ~n2259 & n13966 ;
  assign n13968 = ~n13965 & ~n13967 ;
  assign n13969 = ~\ctl_rf_c1_rf_chsad_reg[17]/NET0131  & ~n2360 ;
  assign n13970 = ~n2260 & n2360 ;
  assign n13971 = ~n2259 & n13970 ;
  assign n13972 = ~n13969 & ~n13971 ;
  assign n13973 = ~\ctl_rf_c0_rf_chsad_reg[17]/NET0131  & ~n2485 ;
  assign n13974 = ~n2260 & n2485 ;
  assign n13975 = ~n2259 & n13974 ;
  assign n13976 = ~n13973 & ~n13975 ;
  assign n13977 = ~\ctl_rf_c2_rf_chsad_reg[17]/NET0131  & ~n2490 ;
  assign n13978 = ~n2260 & n2490 ;
  assign n13979 = ~n2259 & n13978 ;
  assign n13980 = ~n13977 & ~n13979 ;
  assign n13981 = ~\ctl_rf_c4_rf_chtsz_reg[7]/NET0131  & ~n8632 ;
  assign n13982 = ~n2247 & n8632 ;
  assign n13983 = ~n2246 & n13982 ;
  assign n13984 = ~n13981 & ~n13983 ;
  assign n13985 = ~\ctl_rf_c2_rf_chsad_reg[15]/NET0131  & ~n9232 ;
  assign n13986 = ~n3763 & n9232 ;
  assign n13987 = ~n3762 & n13986 ;
  assign n13988 = ~n13985 & ~n13987 ;
  assign n13989 = ~\ctl_rf_c6_rf_chllp_reg[18]/NET0131  & ~n10191 ;
  assign n13990 = ~n2400 & n10191 ;
  assign n13991 = ~n2399 & n13990 ;
  assign n13992 = ~n13989 & ~n13991 ;
  assign n13993 = ~\ctl_rf_c0_rf_chllp_reg[18]/NET0131  & ~n10543 ;
  assign n13994 = ~n2400 & n10543 ;
  assign n13995 = ~n2399 & n13994 ;
  assign n13996 = ~n13993 & ~n13995 ;
  assign n13997 = ~\ctl_rf_c6_rf_chllp_reg[22]/NET0131  & ~n10191 ;
  assign n13998 = ~n2500 & n10191 ;
  assign n13999 = ~n2499 & n13998 ;
  assign n14000 = ~n13997 & ~n13999 ;
  assign n14001 = ~\ctl_rf_c0_rf_chllp_reg[22]/NET0131  & ~n10543 ;
  assign n14002 = ~n2500 & n10543 ;
  assign n14003 = ~n2499 & n14002 ;
  assign n14004 = ~n14001 & ~n14003 ;
  assign n14005 = ~\ctl_rf_c0_rf_chllp_reg[21]/NET0131  & ~n10543 ;
  assign n14006 = ~n2366 & n10543 ;
  assign n14007 = ~n2365 & n14006 ;
  assign n14008 = ~n14005 & ~n14007 ;
  assign n14009 = ~\ctl_rf_c0_rf_chllp_reg[17]/NET0131  & ~n10543 ;
  assign n14010 = ~n2260 & n10543 ;
  assign n14011 = ~n2259 & n14010 ;
  assign n14012 = ~n14009 & ~n14011 ;
  assign n14013 = ~\ctl_rf_c1_rf_chsad_reg[19]/NET0131  & ~n2360 ;
  assign n14014 = n2360 & ~n2409 ;
  assign n14015 = ~n2408 & n14014 ;
  assign n14016 = ~n14013 & ~n14015 ;
  assign n14017 = ~\ctl_rf_c1_rf_chsad_reg[3]/NET0131  & ~n2236 ;
  assign n14018 = n2236 & ~n9044 ;
  assign n14019 = ~n9043 & n14018 ;
  assign n14020 = ~n14017 & ~n14019 ;
  assign n14021 = ~\ctl_rf_c3_rf_chllp_reg[21]/NET0131  & ~n9871 ;
  assign n14022 = ~n2366 & n9871 ;
  assign n14023 = ~n2365 & n14022 ;
  assign n14024 = ~n14021 & ~n14023 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g16/_0_  = n2250 ;
  assign \g58487/_0_  = n2263 ;
  assign \g58489/_0_  = n2271 ;
  assign \g58491/_0_  = n2282 ;
  assign \g58493/_0_  = n2287 ;
  assign \g58495/_0_  = n2294 ;
  assign \g58497/_0_  = n2299 ;
  assign \g58499/_0_  = n2310 ;
  assign \g58500/_0_  = n2316 ;
  assign \g58501/_0_  = n2323 ;
  assign \g58502/_0_  = n2329 ;
  assign \g58504/_0_  = n2334 ;
  assign \g58505/_0_  = n2339 ;
  assign \g58507/_0_  = n2344 ;
  assign \g58508/_0_  = n2349 ;
  assign \g58509/_0_  = n2354 ;
  assign \g58510/_0_  = n2359 ;
  assign \g58556/_0_  = n2369 ;
  assign \g58557/_0_  = n2374 ;
  assign \g58558/_0_  = n2379 ;
  assign \g58559/_0_  = n2384 ;
  assign \g58560/_0_  = n2389 ;
  assign \g58561/_0_  = n2394 ;
  assign \g58562/_0_  = n2403 ;
  assign \g58563/_0_  = n2412 ;
  assign \g58566/_0_  = n2416 ;
  assign \g58567/_0_  = n2420 ;
  assign \g58568/_0_  = n2424 ;
  assign \g58569/_0_  = n2428 ;
  assign \g58570/_0_  = n2432 ;
  assign \g58571/_0_  = n2436 ;
  assign \g58572/_0_  = n2440 ;
  assign \g58573/_0_  = n2444 ;
  assign \g58574/_0_  = n2448 ;
  assign \g58575/_0_  = n2452 ;
  assign \g58576/_0_  = n2456 ;
  assign \g58577/_0_  = n2460 ;
  assign \g58578/_0_  = n2464 ;
  assign \g58579/_0_  = n2468 ;
  assign \g58580/_0_  = n2472 ;
  assign \g58581/_0_  = n2476 ;
  assign \g58584/_0_  = n2480 ;
  assign \g58585/_0_  = n2484 ;
  assign \g58586/_0_  = n2489 ;
  assign \g58587/_0_  = n2494 ;
  assign \g58588/_0_  = n2503 ;
  assign \g58589/_0_  = n2507 ;
  assign \g58590/_0_  = n2511 ;
  assign \g58591/_0_  = n2515 ;
  assign \g58592/_0_  = n2519 ;
  assign \g58593/_0_  = n2523 ;
  assign \g58594/_0_  = n2532 ;
  assign \g58595/_0_  = n2536 ;
  assign \g58596/_0_  = n2540 ;
  assign \g58597/_0_  = n2544 ;
  assign \g58598/_0_  = n2548 ;
  assign \g58599/_0_  = n2552 ;
  assign \g58600/_0_  = n2556 ;
  assign \g58601/_0_  = n2560 ;
  assign \g58602/_0_  = n2569 ;
  assign \g58603/_0_  = n2578 ;
  assign \g58604/_0_  = n2582 ;
  assign \g58605/_0_  = n2586 ;
  assign \g58606/_0_  = n2590 ;
  assign \g58607/_0_  = n2594 ;
  assign \g58608/_0_  = n2598 ;
  assign \g58609/_0_  = n2602 ;
  assign \g58610/_0_  = n2606 ;
  assign \g58611/_0_  = n2610 ;
  assign \g58612/_0_  = n2614 ;
  assign \g58613/_0_  = n2618 ;
  assign \g58614/_0_  = n2622 ;
  assign \g58615/_0_  = n2626 ;
  assign \g58616/_0_  = n2630 ;
  assign \g58617/_0_  = n2634 ;
  assign \g58618/_0_  = n2638 ;
  assign \g58619/_0_  = n2642 ;
  assign \g58620/_0_  = n2646 ;
  assign \g58621/_0_  = n2650 ;
  assign \g58622/_0_  = n2654 ;
  assign \g58623/_0_  = n2658 ;
  assign \g58624/_0_  = n2662 ;
  assign \g58625/_0_  = n2666 ;
  assign \g58626/_0_  = n2670 ;
  assign \g58627/_0_  = n2674 ;
  assign \g58723/_0_  = n2683 ;
  assign \g58734/_0_  = n2687 ;
  assign \g58737/_0_  = n2691 ;
  assign \g58741/_0_  = n2695 ;
  assign \g58749/_0_  = n2699 ;
  assign \g58754/_0_  = n2703 ;
  assign \g58762/_0_  = n2707 ;
  assign \g58763/_0_  = n2711 ;
  assign \g58764/_0_  = n2715 ;
  assign \g58765/_0_  = n2719 ;
  assign \g58766/_0_  = n2723 ;
  assign \g58767/_0_  = n2727 ;
  assign \g58768/_0_  = n2731 ;
  assign \g58769/_0_  = n2735 ;
  assign \g58770/_0_  = n2739 ;
  assign \g58771/_0_  = n2743 ;
  assign \g59788/_0_  = n2845 ;
  assign \g59832/_0_  = ~n2931 ;
  assign \g59873/_0_  = n2952 ;
  assign \g59874/_0_  = ~n2968 ;
  assign \g59893/_0_  = ~n3207 ;
  assign \g59894/_0_  = ~n3302 ;
  assign \g59895/_0_  = ~n3389 ;
  assign \g59896/_0_  = ~n3484 ;
  assign \g59923/_0_  = n3508 ;
  assign \g60031/_0_  = ~n3549 ;
  assign \g60032/_0_  = ~n3589 ;
  assign \g60033/_0_  = ~n3641 ;
  assign \g60036/_0_  = ~n3661 ;
  assign \g60037/_0_  = ~n3679 ;
  assign \g60038/_0_  = ~n3697 ;
  assign \g60165/_0_  = ~n3734 ;
  assign \g60186/_2__syn_2  = n3735 ;
  assign \g60187/_0_  = ~n3752 ;
  assign \g60188/_0_  = ~n3754 ;
  assign \g60258/_0_  = ~n4064 ;
  assign \g60259/_0_  = ~n4083 ;
  assign \g60260/_0_  = ~n4100 ;
  assign \g60261/_0_  = ~n4117 ;
  assign \g60263/_0_  = ~n4134 ;
  assign \g60264/_0_  = ~n4151 ;
  assign \g60265/_0_  = ~n4168 ;
  assign \g60266/_0_  = ~n4185 ;
  assign \g60267/_0_  = n4503 ;
  assign \g60303/_3_  = ~n4532 ;
  assign \g60360/_0_  = n4537 ;
  assign \g60361/_0_  = ~n4546 ;
  assign \g60401/_00_  = ~n4553 ;
  assign \g60428/_0_  = ~n4563 ;
  assign \g60429/_0_  = n4568 ;
  assign \g60448/_0_  = ~n5015 ;
  assign \g60449/_0_  = ~n5153 ;
  assign \g60974/_0_  = ~n5167 ;
  assign \g61072/_0_  = ~n5179 ;
  assign \g61073/_0_  = ~n5190 ;
  assign \g61074/_0_  = ~n5200 ;
  assign \g61075/_0_  = ~n5210 ;
  assign \g61076/_0_  = ~n5220 ;
  assign \g61077/_0_  = ~n5230 ;
  assign \g61078/_0_  = ~n5240 ;
  assign \g61079/_0_  = ~n5250 ;
  assign \g61486/_0_  = ~n5255 ;
  assign \g61502/_3_  = n5262 ;
  assign \g61879/_0_  = ~n5268 ;
  assign \g62077/_0_  = n5280 ;
  assign \g62078/_0_  = n5676 ;
  assign \g62079/_0_  = n5786 ;
  assign \g62080/_0_  = n6131 ;
  assign \g62081/_0_  = n6457 ;
  assign \g62082/_0_  = n6760 ;
  assign \g62083/_0_  = n7063 ;
  assign \g62084/_0_  = n7223 ;
  assign \g62085/_0_  = n7526 ;
  assign \g62086/_0_  = n7845 ;
  assign \g62087/_0_  = n8004 ;
  assign \g62088/_0_  = n8148 ;
  assign \g62089/_0_  = n8292 ;
  assign \g62090/_0_  = n8436 ;
  assign \g62091/_0_  = n8576 ;
  assign \g62629/_0_  = n8590 ;
  assign \g62630/_0_  = n8599 ;
  assign \g62631/_0_  = n8603 ;
  assign \g62632/_0_  = n8608 ;
  assign \g62633/_0_  = n8614 ;
  assign \g62634/_0_  = n8618 ;
  assign \g62635/_0_  = n8622 ;
  assign \g62637/_0_  = n8628 ;
  assign \g62638/_0_  = n8636 ;
  assign \g62639/_0_  = n8640 ;
  assign \g62641/_0_  = n8645 ;
  assign \g62643/_0_  = n8650 ;
  assign \g62645/_0_  = n8655 ;
  assign \g62646/_0_  = n8663 ;
  assign \g62647/_0_  = n8667 ;
  assign \g62648/_0_  = n8671 ;
  assign \g62649/_0_  = n8676 ;
  assign \g62650/_0_  = n8682 ;
  assign \g62651/_0_  = n8686 ;
  assign \g62652/_0_  = n8690 ;
  assign \g62655/_0_  = n8695 ;
  assign \g62656/_0_  = n8700 ;
  assign \g62657/_0_  = n8704 ;
  assign \g62658/_0_  = n8708 ;
  assign \g62659/_0_  = n8717 ;
  assign \g62660/_0_  = n8722 ;
  assign \g62661/_0_  = n8727 ;
  assign \g62662/_0_  = n8731 ;
  assign \g62663/_0_  = n8735 ;
  assign \g62664/_0_  = n8739 ;
  assign \g62665/_0_  = n8743 ;
  assign \g62667/_0_  = n8747 ;
  assign \g62668/_0_  = n8751 ;
  assign \g62669/_0_  = n8762 ;
  assign \g62670/_0_  = n8771 ;
  assign \g62671/_0_  = n8775 ;
  assign \g62672/_0_  = n8784 ;
  assign \g62673/_0_  = n8794 ;
  assign \g62674/_0_  = n8798 ;
  assign \g62675/_0_  = n8802 ;
  assign \g62676/_0_  = n8811 ;
  assign \g62677/_0_  = n8816 ;
  assign \g62678/_0_  = n8820 ;
  assign \g62679/_0_  = n8824 ;
  assign \g62680/_0_  = n8828 ;
  assign \g62681/_0_  = n8832 ;
  assign \g62682/_0_  = n8836 ;
  assign \g62683/_0_  = n8840 ;
  assign \g62684/_0_  = n8845 ;
  assign \g62685/_0_  = n8851 ;
  assign \g62686/_0_  = n8856 ;
  assign \g62687/_0_  = n8860 ;
  assign \g62688/_0_  = n8864 ;
  assign \g62689/_0_  = n8868 ;
  assign \g62690/_0_  = n8872 ;
  assign \g62691/_0_  = n8876 ;
  assign \g62692/_0_  = n8880 ;
  assign \g62693/_0_  = n8885 ;
  assign \g62694/_0_  = n8890 ;
  assign \g62695/_0_  = n8894 ;
  assign \g62696/_0_  = n8898 ;
  assign \g62697/_0_  = n8902 ;
  assign \g62698/_0_  = n8906 ;
  assign \g62699/_0_  = n8910 ;
  assign \g62700/_0_  = n8914 ;
  assign \g62701/_0_  = n8919 ;
  assign \g62702/_0_  = n8923 ;
  assign \g62703/_0_  = n8928 ;
  assign \g62704/_0_  = n8932 ;
  assign \g62705/_0_  = n8936 ;
  assign \g62706/_0_  = n8940 ;
  assign \g62707/_0_  = n8944 ;
  assign \g62708/_0_  = n8948 ;
  assign \g62709/_0_  = n8953 ;
  assign \g62710/_0_  = n8957 ;
  assign \g62711/_0_  = n8961 ;
  assign \g62712/_0_  = n8966 ;
  assign \g62713/_0_  = n8970 ;
  assign \g62714/_0_  = n8974 ;
  assign \g62715/_0_  = n8978 ;
  assign \g62716/_0_  = n8982 ;
  assign \g62721/_0_  = n8986 ;
  assign \g62722/_0_  = n8995 ;
  assign \g62723/_0_  = n9004 ;
  assign \g62725/_0_  = n9008 ;
  assign \g62726/_0_  = n9012 ;
  assign \g62727/_0_  = n9021 ;
  assign \g62728/_0_  = n9030 ;
  assign \g62729/_0_  = n9034 ;
  assign \g62730/_0_  = n9038 ;
  assign \g62731/_0_  = n9047 ;
  assign \g62732/_0_  = n9051 ;
  assign \g62733/_0_  = n9056 ;
  assign \g62734/_0_  = n9060 ;
  assign \g62735/_0_  = n9064 ;
  assign \g62736/_0_  = n9068 ;
  assign \g62737/_0_  = n9072 ;
  assign \g62738/_0_  = n9076 ;
  assign \g62739/_0_  = n9080 ;
  assign \g62740/_0_  = n9084 ;
  assign \g62741/_0_  = n9088 ;
  assign \g62742/_0_  = n9092 ;
  assign \g62743/_0_  = n9097 ;
  assign \g62744/_0_  = n9101 ;
  assign \g62745/_0_  = n9105 ;
  assign \g62746/_0_  = n9109 ;
  assign \g62747/_0_  = n9113 ;
  assign \g62748/_0_  = n9117 ;
  assign \g62749/_0_  = n9121 ;
  assign \g62750/_0_  = n9125 ;
  assign \g62751/_0_  = n9129 ;
  assign \g62752/_0_  = n9133 ;
  assign \g62753/_0_  = n9138 ;
  assign \g62754/_0_  = n9142 ;
  assign \g62755/_0_  = n9147 ;
  assign \g62756/_0_  = n9151 ;
  assign \g62757/_0_  = n9156 ;
  assign \g62758/_0_  = n9160 ;
  assign \g62759/_0_  = n9164 ;
  assign \g62760/_0_  = n9168 ;
  assign \g62761/_0_  = n9172 ;
  assign \g62762/_0_  = n9176 ;
  assign \g62763/_0_  = n9180 ;
  assign \g62764/_0_  = n9184 ;
  assign \g62765/_0_  = n9188 ;
  assign \g62766/_0_  = n9192 ;
  assign \g62767/_0_  = n9197 ;
  assign \g62768/_0_  = n9201 ;
  assign \g62769/_0_  = n9205 ;
  assign \g62770/_0_  = n9209 ;
  assign \g62771/_0_  = n9213 ;
  assign \g62772/_0_  = n9218 ;
  assign \g62773/_0_  = n9222 ;
  assign \g62774/_0_  = n9226 ;
  assign \g62775/_0_  = n9231 ;
  assign \g62776/_0_  = n9236 ;
  assign \g62777/_0_  = n9240 ;
  assign \g62778/_0_  = n9244 ;
  assign \g62779/_0_  = n9248 ;
  assign \g62780/_0_  = n9252 ;
  assign \g62781/_0_  = n9256 ;
  assign \g62783/_0_  = n9260 ;
  assign \g62784/_0_  = n9264 ;
  assign \g62785/_0_  = n9268 ;
  assign \g62786/_0_  = n9272 ;
  assign \g62787/_0_  = n9276 ;
  assign \g62788/_0_  = n9280 ;
  assign \g62789/_0_  = n9284 ;
  assign \g62790/_0_  = n9288 ;
  assign \g62791/_0_  = n9293 ;
  assign \g62792/_0_  = n9297 ;
  assign \g62793/_0_  = n9301 ;
  assign \g62794/_0_  = n9306 ;
  assign \g62795/_0_  = n9310 ;
  assign \g62797/_0_  = n9314 ;
  assign \g62798/_0_  = n9318 ;
  assign \g62799/_0_  = n9322 ;
  assign \g62800/_0_  = n9326 ;
  assign \g62801/_0_  = n9330 ;
  assign \g62802/_0_  = n9334 ;
  assign \g62803/_0_  = n9338 ;
  assign \g62804/_0_  = n9343 ;
  assign \g62805/_0_  = n9347 ;
  assign \g62806/_0_  = n9351 ;
  assign \g62807/_0_  = n9355 ;
  assign \g62808/_0_  = n9359 ;
  assign \g62809/_0_  = n9363 ;
  assign \g62810/_0_  = n9367 ;
  assign \g62811/_0_  = n9371 ;
  assign \g62812/_0_  = n9375 ;
  assign \g62813/_0_  = n9379 ;
  assign \g62814/_0_  = n9383 ;
  assign \g62815/_0_  = n9387 ;
  assign \g62816/_0_  = n9391 ;
  assign \g62817/_0_  = n9395 ;
  assign \g62818/_0_  = n9399 ;
  assign \g63108/_0_  = ~n9694 ;
  assign \g63117/_0_  = ~n9724 ;
  assign \g63125/_0_  = n9731 ;
  assign \g63126/_0_  = n9735 ;
  assign \g63127/_0_  = n9739 ;
  assign \g63128/_0_  = n9743 ;
  assign \g63129/_0_  = n9747 ;
  assign \g63130/_0_  = n9751 ;
  assign \g63131/_0_  = n9757 ;
  assign \g63132/_0_  = n9761 ;
  assign \g63133/_0_  = n9765 ;
  assign \g63134/_0_  = n9769 ;
  assign \g63135/_0_  = n9773 ;
  assign \g63136/_0_  = n9777 ;
  assign \g63137/_0_  = n9781 ;
  assign \g63138/_0_  = n9792 ;
  assign \g63139/_0_  = n9801 ;
  assign \g63140/_0_  = n9810 ;
  assign \g63141/_0_  = n9819 ;
  assign \g63142/_0_  = n9825 ;
  assign \g63143/_0_  = n9829 ;
  assign \g63144/_0_  = n9833 ;
  assign \g63145/_0_  = n9837 ;
  assign \g63146/_0_  = n9841 ;
  assign \g63147/_0_  = n9845 ;
  assign \g63148/_0_  = n9850 ;
  assign \g63149/_0_  = n9854 ;
  assign \g63150/_0_  = n9858 ;
  assign \g63151/_0_  = n9862 ;
  assign \g63152/_0_  = n9866 ;
  assign \g63153/_0_  = n9870 ;
  assign \g63154/_0_  = n9875 ;
  assign \g63155/_0_  = n9879 ;
  assign \g63156/_0_  = n9883 ;
  assign \g63157/_0_  = n9887 ;
  assign \g63159/_0_  = n9891 ;
  assign \g63160/_0_  = n9895 ;
  assign \g63161/_0_  = n9900 ;
  assign \g63162/_0_  = n9904 ;
  assign \g63163/_0_  = n9908 ;
  assign \g63164/_0_  = n9912 ;
  assign \g63165/_0_  = n9917 ;
  assign \g63166/_0_  = n9921 ;
  assign \g63167/_0_  = n9925 ;
  assign \g63168/_0_  = n9929 ;
  assign \g63169/_0_  = n9933 ;
  assign \g63170/_0_  = n9937 ;
  assign \g63171/_0_  = n9945 ;
  assign \g63172/_0_  = n9949 ;
  assign \g63173/_0_  = n9953 ;
  assign \g63174/_0_  = n9957 ;
  assign \g63175/_0_  = n9961 ;
  assign \g63176/_0_  = n9965 ;
  assign \g63177/_0_  = n9971 ;
  assign \g63178/_0_  = n9975 ;
  assign \g63179/_0_  = n9979 ;
  assign \g63180/_0_  = n9983 ;
  assign \g63181/_0_  = n9987 ;
  assign \g63182/_0_  = n9991 ;
  assign \g63183/_0_  = n9995 ;
  assign \g63184/_0_  = n10001 ;
  assign \g63185/_0_  = n10005 ;
  assign \g63186/_0_  = n10009 ;
  assign \g63187/_0_  = n10013 ;
  assign \g63188/_0_  = n10019 ;
  assign \g63189/_0_  = n10023 ;
  assign \g63190/_0_  = n10027 ;
  assign \g63191/_0_  = n10031 ;
  assign \g63192/_0_  = n10035 ;
  assign \g63193/_0_  = n10039 ;
  assign \g63194/_0_  = n10044 ;
  assign \g63195/_0_  = n10048 ;
  assign \g63196/_0_  = n10052 ;
  assign \g63197/_0_  = n10056 ;
  assign \g63198/_0_  = n10060 ;
  assign \g63199/_0_  = n10064 ;
  assign \g63200/_0_  = n10069 ;
  assign \g63201/_0_  = n10073 ;
  assign \g63202/_0_  = n10077 ;
  assign \g63203/_0_  = n10081 ;
  assign \g63204/_0_  = n10085 ;
  assign \g63205/_0_  = n10089 ;
  assign \g63206/_0_  = n10093 ;
  assign \g63207/_0_  = n10098 ;
  assign \g63208/_0_  = n10102 ;
  assign \g63209/_0_  = n10106 ;
  assign \g63210/_0_  = n10110 ;
  assign \g63211/_0_  = n10115 ;
  assign \g63212/_0_  = n10119 ;
  assign \g63213/_0_  = n10123 ;
  assign \g63214/_0_  = ~n10137 ;
  assign \g63215/_0_  = n10141 ;
  assign \g63216/_0_  = n10145 ;
  assign \g63217/_0_  = n10149 ;
  assign \g63218/_0_  = ~n10162 ;
  assign \g63219/_0_  = n10169 ;
  assign \g63220/_0_  = n10173 ;
  assign \g63221/_0_  = n10177 ;
  assign \g63222/_0_  = n10181 ;
  assign \g63223/_0_  = n10185 ;
  assign \g63224/_0_  = n10189 ;
  assign \g63225/_0_  = n10195 ;
  assign \g63226/_0_  = n10199 ;
  assign \g63228/_0_  = n10203 ;
  assign \g63229/_0_  = n10207 ;
  assign \g63231/_0_  = n10211 ;
  assign \g63232/_0_  = n10217 ;
  assign \g63233/_0_  = n10221 ;
  assign \g63234/_0_  = n10225 ;
  assign \g63235/_0_  = n10229 ;
  assign \g63236/_0_  = n10235 ;
  assign \g63237/_0_  = n10239 ;
  assign \g63238/_0_  = n10243 ;
  assign \g63239/_0_  = n10247 ;
  assign \g63240/_0_  = n10251 ;
  assign \g63241/_0_  = n10255 ;
  assign \g63242/_0_  = ~n10268 ;
  assign \g63244/_0_  = ~n10281 ;
  assign \g63246/_0_  = ~n10293 ;
  assign \g63247/_0_  = n10298 ;
  assign \g63248/_0_  = n10302 ;
  assign \g63249/_0_  = n10306 ;
  assign \g63250/_0_  = n10310 ;
  assign \g63251/_0_  = n10314 ;
  assign \g63252/_0_  = n10318 ;
  assign \g63253/_0_  = n10323 ;
  assign \g63254/_0_  = n10327 ;
  assign \g63255/_0_  = n10331 ;
  assign \g63256/_0_  = n10335 ;
  assign \g63257/_0_  = n10339 ;
  assign \g63258/_0_  = n10343 ;
  assign \g63259/_0_  = n10347 ;
  assign \g63260/_0_  = n10352 ;
  assign \g63261/_0_  = n10356 ;
  assign \g63262/_0_  = n10360 ;
  assign \g63263/_0_  = n10364 ;
  assign \g63264/_0_  = n10369 ;
  assign \g63265/_0_  = n10373 ;
  assign \g63266/_0_  = n10377 ;
  assign \g63267/_0_  = n10381 ;
  assign \g63268/_0_  = n10385 ;
  assign \g63269/_0_  = n10389 ;
  assign \g63270/_0_  = ~n10401 ;
  assign \g63272/_0_  = ~n10413 ;
  assign \g63291/_0_  = ~n10414 ;
  assign \g63292/_0_  = n10419 ;
  assign \g63293/_0_  = n10423 ;
  assign \g63294/_0_  = n10427 ;
  assign \g63295/_0_  = n10431 ;
  assign \g63298/_0_  = n10436 ;
  assign \g63299/_0_  = n10441 ;
  assign \g63300/_0_  = n10445 ;
  assign \g63301/_0_  = n10449 ;
  assign \g63302/_0_  = n10453 ;
  assign \g63303/_0_  = n10457 ;
  assign \g63304/_0_  = n10462 ;
  assign \g63305/_0_  = n10466 ;
  assign \g63306/_0_  = n10470 ;
  assign \g63307/_0_  = n10474 ;
  assign \g63308/_0_  = n10479 ;
  assign \g63309/_0_  = n10483 ;
  assign \g63310/_0_  = n10488 ;
  assign \g63311/_0_  = n10493 ;
  assign \g63312/_0_  = n10497 ;
  assign \g63313/_0_  = n10501 ;
  assign \g63314/_0_  = n10505 ;
  assign \g63315/_0_  = n10509 ;
  assign \g63316/_0_  = ~n10534 ;
  assign \g63317/_0_  = n10538 ;
  assign \g63318/_0_  = n10542 ;
  assign \g63320/_0_  = n10547 ;
  assign \g63322/_0_  = n10551 ;
  assign \g63323/_0_  = n10555 ;
  assign \g63324/_0_  = n10559 ;
  assign \g63325/_0_  = n10563 ;
  assign \g63326/_0_  = n10567 ;
  assign \g63327/_0_  = n10571 ;
  assign \g63328/_0_  = n10575 ;
  assign \g63329/_0_  = n10584 ;
  assign \g63330/_0_  = n10588 ;
  assign \g63331/_0_  = n10597 ;
  assign \g63332/_0_  = n10601 ;
  assign \g63333/_0_  = n10605 ;
  assign \g63334/_0_  = n10609 ;
  assign \g63335/_0_  = n10613 ;
  assign \g63336/_0_  = n10617 ;
  assign \g63337/_0_  = n10621 ;
  assign \g63338/_0_  = n10625 ;
  assign \g63339/_0_  = n10629 ;
  assign \g63340/_0_  = n10633 ;
  assign \g63341/_0_  = n10637 ;
  assign \g63342/_0_  = n10641 ;
  assign \g63343/_0_  = n10645 ;
  assign \g63344/_0_  = n10649 ;
  assign \g63345/_0_  = n10653 ;
  assign \g63346/_0_  = n10657 ;
  assign \g63347/_0_  = n10661 ;
  assign \g63348/_0_  = n10665 ;
  assign \g63349/_0_  = n10669 ;
  assign \g63350/_0_  = n10673 ;
  assign \g63351/_0_  = n10677 ;
  assign \g63352/_0_  = n10681 ;
  assign \g63353/_0_  = n10685 ;
  assign \g63354/_0_  = n10689 ;
  assign \g63355/_0_  = n10693 ;
  assign \g63356/_0_  = n10697 ;
  assign \g63357/_0_  = n10701 ;
  assign \g63358/_0_  = n10705 ;
  assign \g63359/_0_  = n10709 ;
  assign \g63360/_0_  = n10713 ;
  assign \g63361/_0_  = n10717 ;
  assign \g63362/_0_  = n10721 ;
  assign \g63363/_0_  = n10725 ;
  assign \g63364/_0_  = n10729 ;
  assign \g63365/_0_  = n10733 ;
  assign \g63366/_0_  = n10737 ;
  assign \g63367/_0_  = n10741 ;
  assign \g63368/_0_  = n10745 ;
  assign \g63369/_0_  = n10749 ;
  assign \g63370/_0_  = n10753 ;
  assign \g63371/_0_  = n10757 ;
  assign \g63372/_0_  = n10761 ;
  assign \g63373/_0_  = n10765 ;
  assign \g63374/_0_  = n10769 ;
  assign \g63375/_0_  = n10773 ;
  assign \g63376/_0_  = n10777 ;
  assign \g63377/_0_  = n10781 ;
  assign \g63378/_0_  = n10785 ;
  assign \g63379/_0_  = n10789 ;
  assign \g63380/_0_  = n10793 ;
  assign \g63383/_3_  = ~n10799 ;
  assign \g63386/_0_  = n10803 ;
  assign \g63387/_0_  = n10807 ;
  assign \g63388/_0_  = n10811 ;
  assign \g63389/_0_  = n10815 ;
  assign \g63390/_0_  = n10819 ;
  assign \g63391/_0_  = n10823 ;
  assign \g63392/_0_  = n10827 ;
  assign \g63419/_0_  = n10831 ;
  assign \g63421/_0_  = n10835 ;
  assign \g63422/_0_  = n10839 ;
  assign \g63423/_0_  = n10843 ;
  assign \g63424/_0_  = n10847 ;
  assign \g63425/_0_  = n10851 ;
  assign \g63536/_3_  = ~n10865 ;
  assign \g63625/_0_  = ~n10866 ;
  assign \g63628/_0_  = ~n9693 ;
  assign \g63871/_0_  = ~n10884 ;
  assign \g63874/_0_  = ~n3095 ;
  assign \g63889/_0_  = ~n10890 ;
  assign \g63933/_0_  = ~n10905 ;
  assign \g63945/_0_  = ~n10919 ;
  assign \g63959/_0_  = n10934 ;
  assign \g63962/_0_  = n10948 ;
  assign \g63974/_0_  = n10962 ;
  assign \g63977/_0_  = n10974 ;
  assign \g64035/_0_  = ~n10988 ;
  assign \g64435/_3_  = n11002 ;
  assign \g64939/_0_  = ~n11021 ;
  assign \g65149/_0_  = n11040 ;
  assign \g65632/_3_  = ~n11045 ;
  assign \g65633/_0_  = ~n11049 ;
  assign \g65634/_0_  = ~n11053 ;
  assign \g65635/_0_  = ~n11056 ;
  assign \g65636/_0_  = ~n11059 ;
  assign \g65638/_3_  = ~n11062 ;
  assign \g65640/_3_  = ~n11065 ;
  assign \g65999/_0_  = ~n11075 ;
  assign \g66912/_0_  = ~n11085 ;
  assign \g66914/_0_  = ~n11098 ;
  assign \g67555/_3_  = ~n11101 ;
  assign \g67564/_3_  = ~n11104 ;
  assign \g67567/_3_  = ~n11107 ;
  assign \g67735/_0_  = ~n11114 ;
  assign \g67736/_0_  = ~n11120 ;
  assign \g67737/_0_  = ~n11125 ;
  assign \g67738/_0_  = ~n11130 ;
  assign \g67758/_0_  = ~n11135 ;
  assign \g67760/_0_  = ~n11140 ;
  assign \g67761/_0_  = ~n11145 ;
  assign \g67763/_0_  = ~n11150 ;
  assign \g67766/_0_  = n11155 ;
  assign \g67810/_0_  = n11182 ;
  assign \g67816/_0_  = ~n11194 ;
  assign \g67902/_0_  = ~n11196 ;
  assign \g67927/_0_  = n11206 ;
  assign \g67936/_0_  = ~n11210 ;
  assign \g68067/_0_  = n11224 ;
  assign \g68068/_0_  = n11229 ;
  assign \g68069/_0_  = n11243 ;
  assign \g68070/_0_  = n11248 ;
  assign \g68071/_0_  = n11262 ;
  assign \g68072/_0_  = n11267 ;
  assign \g68073/_0_  = n11281 ;
  assign \g68074/_0_  = n11286 ;
  assign \g68075/_0_  = n11300 ;
  assign \g68076/_0_  = n11305 ;
  assign \g68077/_0_  = n11319 ;
  assign \g68078/_0_  = n11324 ;
  assign \g68079/_0_  = n11338 ;
  assign \g68080/_0_  = n11343 ;
  assign \g68081/_0_  = n11357 ;
  assign \g68082/_0_  = n11362 ;
  assign \g68083/_0_  = n11367 ;
  assign \g68084/_0_  = n11373 ;
  assign \g68085/_0_  = n11379 ;
  assign \g68086/_0_  = n11385 ;
  assign \g68087/_0_  = n11391 ;
  assign \g68088/_0_  = n11397 ;
  assign \g68089/_0_  = n11403 ;
  assign \g68090/_0_  = n11409 ;
  assign \g68091/_0_  = n11415 ;
  assign \g68096/_0_  = n11418 ;
  assign \g68160/_0_  = n11421 ;
  assign \g68218/_0_  = n11424 ;
  assign \g68219/_0_  = n11427 ;
  assign \g68220/_0_  = n11430 ;
  assign \g68221/_0_  = n11433 ;
  assign \g68222/_0_  = n11436 ;
  assign \g68226/_0_  = n11439 ;
  assign \g68247/_0_  = ~n11444 ;
  assign \g68252/_0_  = n11445 ;
  assign \g68632/_0_  = ~n11456 ;
  assign \g68633/_0_  = ~n11461 ;
  assign \g68635/_0_  = ~n11466 ;
  assign \g68640/_0_  = ~n11471 ;
  assign \g68642/_0_  = ~n11476 ;
  assign \g68643/_0_  = ~n11481 ;
  assign \g68644/_0_  = ~n11486 ;
  assign \g68645/_0_  = ~n11491 ;
  assign \g68649/_0_  = ~n11499 ;
  assign \g68668/_2_  = n11501 ;
  assign \g68670/_0_  = ~n11507 ;
  assign \g68681/_3_  = ~n11519 ;
  assign \g68689/_0_  = ~n11527 ;
  assign \g68690/_0_  = ~n11535 ;
  assign \g68691/_0_  = ~n11543 ;
  assign \g68692/_0_  = ~n11551 ;
  assign \g68693/_0_  = ~n11559 ;
  assign \g68694/_0_  = ~n11567 ;
  assign \g68695/_0_  = ~n11575 ;
  assign \g68737/_0_  = ~n11598 ;
  assign \g68742/_0_  = ~n11621 ;
  assign \g68745/_0_  = ~n11644 ;
  assign \g68750/_0_  = ~n11667 ;
  assign \g68759/_0_  = ~n11690 ;
  assign \g68761/_0_  = ~n11713 ;
  assign \g68774/_0_  = ~n4278 ;
  assign \g68775/_0_  = ~n4446 ;
  assign \g68776/_0_  = ~n4399 ;
  assign \g68777/_0_  = ~n4231 ;
  assign \g68778/_0_  = ~n4303 ;
  assign \g68780/_0_  = ~n4469 ;
  assign \g68781/_0_  = ~n4422 ;
  assign \g68782/_0_  = ~n4498 ;
  assign \g68783/_0_  = ~n4373 ;
  assign \g68784/_0_  = ~n4350 ;
  assign \g68785/_0_  = ~n4255 ;
  assign \g68786/_0_  = ~n4208 ;
  assign \g68787/_0_  = ~n11736 ;
  assign \g68790/_0_  = ~n11759 ;
  assign \g68791/_0_  = ~n11782 ;
  assign \g68793/_0_  = ~n11805 ;
  assign \g68794/_0_  = ~n11828 ;
  assign \g68795/_0_  = ~n11851 ;
  assign \g68796/_0_  = ~n11874 ;
  assign \g68797/_0_  = ~n11897 ;
  assign \g68804/_0_  = ~n11920 ;
  assign \g68805/_0_  = ~n11943 ;
  assign \g68807/_0_  = ~n11966 ;
  assign \g68809/_0_  = ~n11989 ;
  assign \g68864/_3_  = ~n12096 ;
  assign \g68865/_3_  = ~n12194 ;
  assign \g68866/_3_  = ~n12292 ;
  assign \g68867/_3_  = ~n12390 ;
  assign \g68868/_3_  = ~n12488 ;
  assign \g68869/_3_  = ~n12586 ;
  assign \g68870/_3_  = ~n12684 ;
  assign \g68871/_3_  = ~n12720 ;
  assign \g68872/_3_  = ~n12818 ;
  assign \g68873/_3_  = ~n12854 ;
  assign \g68874/_3_  = ~n12890 ;
  assign \g68875/_3_  = ~n12926 ;
  assign \g68876/_3_  = ~n12962 ;
  assign \g68877/_3_  = ~n12967 ;
  assign \g68878/_3_  = ~n13003 ;
  assign \g68879/_3_  = ~n13039 ;
  assign \g68880/_3_  = ~n13075 ;
  assign \g68881/_3_  = ~n13080 ;
  assign \g68882/_3_  = ~n13085 ;
  assign \g68883/_3_  = ~n13090 ;
  assign \g68884/_3_  = ~n13095 ;
  assign \g68885/_3_  = ~n13100 ;
  assign \g68886/_3_  = ~n13105 ;
  assign \g68887/_3_  = ~n13110 ;
  assign \g68888/_3_  = ~n13115 ;
  assign \g68889/_3_  = ~n13120 ;
  assign \g68890/_3_  = ~n13125 ;
  assign \g68891/_3_  = ~n13130 ;
  assign \g68892/_3_  = ~n13135 ;
  assign \g68893/_3_  = ~n13140 ;
  assign \g68894/_3_  = ~n13145 ;
  assign \g68895/_3_  = ~n13150 ;
  assign \g69037/_1__syn_2  = n11502 ;
  assign \g69077/_0_  = ~n13157 ;
  assign \g69081/_0_  = ~n13164 ;
  assign \g69084/_0_  = n13170 ;
  assign \g69085/_0_  = ~n13177 ;
  assign \g69086/_0_  = ~n13184 ;
  assign \g69088/_0_  = ~n13191 ;
  assign \g69094/_0_  = ~n13198 ;
  assign \g69095/_0_  = ~n13205 ;
  assign \g69097/_0_  = ~n13212 ;
  assign \g69114/_3_  = ~n13219 ;
  assign \g69116/_3_  = ~n13226 ;
  assign \g69118/_3_  = ~n13233 ;
  assign \g69120/_3_  = ~n13240 ;
  assign \g69122/_3_  = ~n13247 ;
  assign \g69124/_3_  = ~n13254 ;
  assign \g69126/_3_  = ~n13261 ;
  assign \g69128/_3_  = ~n13268 ;
  assign \g69581/_3_  = n9525 ;
  assign \g70303/_1__syn_2  = n13270 ;
  assign \g70304/_1__syn_2  = n13272 ;
  assign \g70305/_1__syn_2  = n13273 ;
  assign \g70306/_1__syn_2  = n13274 ;
  assign \g70353/_1__syn_2  = n13276 ;
  assign \g70359/_2_  = n13277 ;
  assign \g70364/_1__syn_2  = n13278 ;
  assign \g70375/_1__syn_2  = n13279 ;
  assign \g70380/_2_  = n13280 ;
  assign \g70383/_1__syn_2  = n13282 ;
  assign \g70394/_2_  = n13283 ;
  assign \g70395/_2_  = n4076 ;
  assign \g70396/_1__syn_2  = n13285 ;
  assign \g70398/_1__syn_2  = n13287 ;
  assign \g70407/_1_  = n13289 ;
  assign \g70416/_1__syn_2  = n13290 ;
  assign \g70418/_1__syn_2  = n13291 ;
  assign \g70419/_2_  = n4111 ;
  assign \g70424/_1_  = n13293 ;
  assign \g70465/_2_  = n13294 ;
  assign \g70511/_1_  = n13296 ;
  assign \g70512/_1_  = n13298 ;
  assign \g70513/_2_  = n13299 ;
  assign \g70514/_2_  = n4057 ;
  assign \g70516/_2_  = n13300 ;
  assign \g70518/_2_  = n13301 ;
  assign \g70519/_2_  = n4094 ;
  assign \g70520/_2_  = n13302 ;
  assign \g70530/_2_  = n13303 ;
  assign \g70534/_3_  = n9671 ;
  assign \g70536/_3_  = n9688 ;
  assign \g70540/_3_  = n9455 ;
  assign \g70541/_2_  = n13304 ;
  assign \g70545/_3_  = n9508 ;
  assign \g70546/_2_  = n13305 ;
  assign \g70547/_2_  = n4128 ;
  assign \g70550/_3_  = n9597 ;
  assign \g70551/_2_  = n13306 ;
  assign \g70552/_2_  = n4145 ;
  assign \g70558/_3_  = n9580 ;
  assign \g70559/_2_  = n4162 ;
  assign \g70560/_2_  = n13307 ;
  assign \g70562/_3_  = n9437 ;
  assign \g70564/_3_  = n9562 ;
  assign \g70567/_3_  = n9618 ;
  assign \g70568/_2_  = n13308 ;
  assign \g70571/_3_  = n9473 ;
  assign \g70577/_0_  = ~n13324 ;
  assign \g70578/_2_  = n13325 ;
  assign \g70585/_3_  = n9653 ;
  assign \g70586/_2_  = n13326 ;
  assign \g70587/_2_  = n4179 ;
  assign \g70588/_3_  = n13328 ;
  assign \g70602/_3_  = n13330 ;
  assign \g70841/_0_  = n13342 ;
  assign \g70842/_0_  = n13354 ;
  assign \g70843/_0_  = n13366 ;
  assign \g70844/_0_  = n13378 ;
  assign \g70845/_0_  = n13390 ;
  assign \g70846/_0_  = n13402 ;
  assign \g70847/_0_  = n13412 ;
  assign \g70848/_0_  = n13424 ;
  assign \g70849/_0_  = n13436 ;
  assign \g70850/_0_  = n13448 ;
  assign \g70851/_0_  = n13460 ;
  assign \g70852/_0_  = n13472 ;
  assign \g70853/_0_  = n13484 ;
  assign \g70854/_0_  = n13494 ;
  assign \g70855/_0_  = n13506 ;
  assign \g70856/_0_  = n13518 ;
  assign \g70857/_0_  = n13530 ;
  assign \g70858/_0_  = n13542 ;
  assign \g70859/_0_  = n13552 ;
  assign \g70860/_0_  = n13562 ;
  assign \g70861/_0_  = n13572 ;
  assign \g70862/_0_  = n13582 ;
  assign \g70863/_0_  = n13592 ;
  assign \g70864/_0_  = n13602 ;
  assign \g70865/_0_  = n13612 ;
  assign \g70866/_0_  = n13622 ;
  assign \g70867/_0_  = n13632 ;
  assign \g70868/_0_  = n13642 ;
  assign \g70869/_0_  = n13652 ;
  assign \g70870/_0_  = n13662 ;
  assign \g70871/_0_  = n13672 ;
  assign \g70872/_0_  = n13682 ;
  assign \g70944/_1__syn_2  = n13688 ;
  assign \g71042/_1__syn_2  = n13694 ;
  assign \g71064/_1__syn_2  = n13700 ;
  assign \g71065/_1__syn_2  = n13702 ;
  assign \g71076/_1__syn_2  = n13706 ;
  assign \g71077/_1__syn_2  = n13708 ;
  assign \g71202/_1__syn_2  = n13710 ;
  assign \g71204/_1__syn_2  = n13712 ;
  assign \g71236/_0_  = n13713 ;
  assign \g71237/_0_  = n13714 ;
  assign \g71241/_0_  = n13715 ;
  assign \g71242/_0_  = n13716 ;
  assign \g71245/_0_  = n13717 ;
  assign \g71246/_0_  = n13718 ;
  assign \g71306/_0_  = n13719 ;
  assign \g71308/_0_  = n13720 ;
  assign \g71309/_0_  = n13721 ;
  assign \g71310/_0_  = n13722 ;
  assign \g71355/_0_  = n13723 ;
  assign \g71416/_0_  = n13724 ;
  assign \g71417/_0_  = n13725 ;
  assign \g71420/_0_  = n13726 ;
  assign \g71432/_0_  = n13727 ;
  assign \g71434/_0_  = n13728 ;
  assign \g71435/_0_  = n13729 ;
  assign \g71436/_0_  = n13730 ;
  assign \g71446/_0_  = n13731 ;
  assign \g71449/_0_  = n13732 ;
  assign \g71451/_0_  = n13733 ;
  assign \g71452/_0_  = n13734 ;
  assign \g71485/_0_  = n13735 ;
  assign \g71494/_0_  = n13736 ;
  assign \g71499/_0_  = n13737 ;
  assign \g71500/_0_  = n13738 ;
  assign \g71501/_0_  = n13739 ;
  assign \g71502/_0_  = n13740 ;
  assign \g71503/_0_  = n13741 ;
  assign \g71504/_0_  = n13742 ;
  assign \g71505/_0_  = n13743 ;
  assign \g71506/_0_  = n13744 ;
  assign \g71815/_0_  = n13745 ;
  assign \g71823/_0_  = n10437 ;
  assign \g71832/_0_  = n9152 ;
  assign \g71833/_0__syn_2  = n13746 ;
  assign \g71837/_0_  = n8696 ;
  assign \g71838/_0_  = n13748 ;
  assign \g71846/_1__syn_2  = n13749 ;
  assign \g71847/_1__syn_2  = n13750 ;
  assign \g71849/_0_  = n9193 ;
  assign \g71854/_0_  = n8753 ;
  assign \g71858/_1__syn_2  = n2254 ;
  assign \g71859/_1__syn_2  = n13751 ;
  assign \g71863/_0_  = n8812 ;
  assign \g71867/_0_  = n9214 ;
  assign \g71869/_0_  = n9227 ;
  assign \g71872/_1_  = n2335 ;
  assign \g71873/_1__syn_2  = n13752 ;
  assign \g71874/_1__syn_2  = n13756 ;
  assign \g71875/_0_  = n13757 ;
  assign \g71877/_1__syn_2  = n13760 ;
  assign \g71881/_0_  = n10489 ;
  assign \g71906/_0_  = n2340 ;
  assign \g71907/_1__syn_2  = n13761 ;
  assign \g71910/_0_  = n8723 ;
  assign \g71911/_0_  = n13762 ;
  assign \g71912/_1__syn_2  = n13764 ;
  assign \g71913/_1__syn_2  = n13766 ;
  assign \g71914/_1__syn_2  = n13767 ;
  assign \g71918/_0_  = n9289 ;
  assign \g71921/_0_  = n2267 ;
  assign \g71922/_0_  = n13768 ;
  assign \g71929/_1__syn_2  = n13769 ;
  assign \g71931/_1__syn_2  = n13770 ;
  assign \g71938/_1__syn_2  = n13771 ;
  assign \g71942/_0_  = n8881 ;
  assign \g71946/_1__syn_2  = n8678 ;
  assign \g71947/_0_  = n13772 ;
  assign \g71951/_0_  = n10111 ;
  assign \g71958/_1__syn_2  = n13773 ;
  assign \g71965/_0_  = n8886 ;
  assign \g71970/_1__syn_2  = n13775 ;
  assign \g71972/_1__syn_2  = n13776 ;
  assign \g71973/_1__syn_2  = n13777 ;
  assign \g71986/_1__syn_2  = n8659 ;
  assign \g71987/_1__syn_2  = n13779 ;
  assign \g71990/_1__syn_2  = n13781 ;
  assign \g71991/_1__syn_2  = n13782 ;
  assign \g71992/_1__syn_2  = n13783 ;
  assign \g71994/_1__syn_2  = n9339 ;
  assign \g71997/_1__syn_2  = n8949 ;
  assign \g72001/_1__syn_2  = n13784 ;
  assign \g72013/_1__syn_2  = n8962 ;
  assign \g72021/_1__syn_2  = n13785 ;
  assign \g72030/_0_  = n2283 ;
  assign \g72031/_0__syn_2  = n13786 ;
  assign \g72036/_1__syn_2  = n13787 ;
  assign \g72038/_0_  = n2330 ;
  assign \g72042/_1__syn_2  = n13788 ;
  assign \g72047/_1__syn_2  = n2350 ;
  assign \g72048/_1__syn_2  = n13789 ;
  assign \g72049/_1__syn_2  = n13790 ;
  assign \g72056/_0_  = n2345 ;
  assign \g72064/_1__syn_2  = n10365 ;
  assign \g72073/_1__syn_2  = n13791 ;
  assign \g72075/_0_  = n9134 ;
  assign \g72078/_0_  = n9143 ;
  assign \g72081/_0_  = n2355 ;
  assign \g72091/_0_  = n13793 ;
  assign \g72096/_0_  = n13795 ;
  assign \g72100/_1__syn_2  = n9821 ;
  assign \g72113/_0_  = n8785 ;
  assign \g72118/_0_  = n2301 ;
  assign \g72121/_1__syn_2  = n8581 ;
  assign \g72122/_1__syn_2  = n13796 ;
  assign \g72125/_1__syn_2  = n8915 ;
  assign \g72128/_0_  = n13798 ;
  assign \g72140/_0_  = n13800 ;
  assign \g72144/_1__syn_2  = n9913 ;
  assign \g72154/_1__syn_2  = n9052 ;
  assign \g72159/_0_  = n2312 ;
  assign \g72164/_1__syn_2  = n8610 ;
  assign \g72165/_1__syn_2  = n13801 ;
  assign \g72167/_1__syn_2  = n8847 ;
  assign \g72170/_1__syn_2  = n2278 ;
  assign \g72172/_1__syn_2  = n13802 ;
  assign \g72173/_0_  = n13804 ;
  assign \g72177/_1__syn_2  = n10015 ;
  assign \g72189/_0_  = n8852 ;
  assign \g72194/_0_  = n2319 ;
  assign \g72196/_0_  = n8841 ;
  assign \g72198/_0_  = n13806 ;
  assign \g72206/_1__syn_2  = n9093 ;
  assign \g72209/_1__syn_2  = n2290 ;
  assign \g72210/_1__syn_2  = n13807 ;
  assign \g72211/_0_  = n13809 ;
  assign \g72215/_0_  = n10231 ;
  assign \g72227/_1__syn_2  = n8924 ;
  assign \g72229/_1__syn_2  = n2325 ;
  assign \g72230/_0_  = n13811 ;
  assign \g72239/_0_  = ~n13817 ;
  assign \g72250/_3_  = ~n13818 ;
  assign \g72251/_3_  = ~n13819 ;
  assign \g72252/_3_  = ~n13820 ;
  assign \g72253/_3_  = ~n13821 ;
  assign \g72254/_3_  = ~n13822 ;
  assign \g72255/_3_  = ~n13823 ;
  assign \g72256/_3_  = ~n13824 ;
  assign \g72257/_3_  = ~n13825 ;
  assign \g72259/_3_  = ~n13826 ;
  assign \g72260/_3_  = ~n13827 ;
  assign \g72261/_3_  = ~n13828 ;
  assign \g72262/_3_  = ~n13829 ;
  assign \g72263/_3_  = ~n13830 ;
  assign \g72264/_3_  = ~n13831 ;
  assign \g72265/_3_  = ~n13832 ;
  assign \g72266/_3_  = ~n13833 ;
  assign \g72267/_3_  = ~n13834 ;
  assign \g72273/_3_  = ~n13835 ;
  assign \g72275/_3_  = ~n13836 ;
  assign \g72282/_3_  = ~n13837 ;
  assign \g72285/_3_  = ~n13838 ;
  assign \g72293/_3_  = ~n13839 ;
  assign \g72304/_3_  = ~n13840 ;
  assign \g72305/_3_  = ~n13841 ;
  assign \g72306/_3_  = ~n13842 ;
  assign \g72307/_3_  = ~n13843 ;
  assign \g72309/_3_  = ~n11108 ;
  assign \g72310/_3_  = ~n13844 ;
  assign \g72324/_3_  = ~n3772 ;
  assign \g72325/_3_  = ~n13845 ;
  assign \g72326/_3_  = ~n13846 ;
  assign \g72327/_3_  = ~n13847 ;
  assign \g72711/_0_  = ~n13877 ;
  assign \g72763/_0_  = ~n13880 ;
  assign \g72966/_0_  = ~n13889 ;
  assign \g72967/_0_  = ~n13892 ;
  assign \g73018/_0_  = ~n2983 ;
  assign \g73058/_0_  = ~n2998 ;
  assign \g73062/_0_  = ~n2991 ;
  assign \g73067/_0_  = ~n13899 ;
  assign \g73068/_0_  = ~n13901 ;
  assign \g73207/_0_  = ~n13316 ;
  assign \g75007/_1__syn_2  = n13904 ;
  assign \g75568/_1_  = n13854 ;
  assign \g75792/_0_  = n13905 ;
  assign \g75836/_0_  = n13906 ;
  assign \g76027/_0_  = n13907 ;
  assign \g76034/_0_  = n13908 ;
  assign \g76108/_0_  = n13909 ;
  assign \g76130/_0_  = n13910 ;
  assign \g76266/_0_  = n13911 ;
  assign \g76315/_0_  = n13912 ;
  assign \g76569/_0_  = ~n13914 ;
  assign \g76714/_0_  = n13916 ;
  assign \g77122/_1__syn_2  = n4521 ;
  assign \g77709/_1_  = n10794 ;
  assign \g81909/_0_  = n13920 ;
  assign \g81922/_0_  = n13924 ;
  assign \g81926/_1__syn_2  = n2295 ;
  assign \g82197/_1_  = n2834 ;
  assign \g82272/_0_  = n13928 ;
  assign \g82291/_0_  = n13932 ;
  assign \g82716/_0_  = n13936 ;
  assign \g82718/_0_  = n9302 ;
  assign \g82738/_0_  = n13940 ;
  assign \g82769/_0_  = n13944 ;
  assign \g82775/_0_  = n13948 ;
  assign \g82779/_1__syn_2  = n8646 ;
  assign \g82804/_0_  = n13952 ;
  assign \g82810/_0_  = n13956 ;
  assign \g82817/_0_  = n13960 ;
  assign \g82823/_0_  = n13964 ;
  assign \g82835/_0_  = n13968 ;
  assign \g82841/_0_  = n13972 ;
  assign \g82847/_0_  = n13976 ;
  assign \g82853/_0_  = n13980 ;
  assign \g82859/_0_  = n13984 ;
  assign \g82862/_1__syn_2  = n8632 ;
  assign \g82956/_0_  = n13988 ;
  assign \g82959/_1_  = n9232 ;
  assign \g83020/_0_  = n13992 ;
  assign \g83025/_0_  = n13996 ;
  assign \g83078/_0_  = n14000 ;
  assign \g83083/_0_  = n14004 ;
  assign \g83121/_0_  = n14008 ;
  assign \g83135/_0_  = n14012 ;
  assign \g83205/_0_  = n14016 ;
  assign \g83240/_0_  = n14020 ;
  assign \g83509/_1__syn_2  = n9601 ;
  assign \g83769/_0_  = n14024 ;
  assign \h0lock_pad  = 1'b0 ;
  assign \h1sel_br[7]_pad  = n9635 ;
  assign \h1sel_dma[0]_pad  = n9545 ;
  assign \h1sel_dma[4]_pad  = n9420 ;
  assign \h1sel_dma[7]_pad  = n9490 ;
endmodule
