module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  output f_pad ;
  output g_pad ;
  output h_pad ;
  wire n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 ;
  assign n6 = b_pad & ~c_pad ;
  assign n7 = ~b_pad & c_pad ;
  assign n8 = ~n6 & ~n7 ;
  assign n9 = a_pad & n8 ;
  assign n10 = ~a_pad & ~n8 ;
  assign n11 = ~n9 & ~n10 ;
  assign n12 = d_pad & e_pad ;
  assign n13 = ~d_pad & ~e_pad ;
  assign n14 = ~n12 & ~n13 ;
  assign n15 = a_pad & b_pad ;
  assign n16 = ~a_pad & ~b_pad ;
  assign n17 = c_pad & ~n16 ;
  assign n18 = ~n15 & ~n17 ;
  assign n19 = n14 & ~n18 ;
  assign n20 = ~n14 & n18 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = ~n13 & ~n18 ;
  assign n23 = ~n12 & ~n22 ;
  assign f_pad = ~n11 ;
  assign g_pad = n21 ;
  assign h_pad = ~n23 ;
endmodule
