module top( \101(0)_pad  , \104(1)_pad  , \107(2)_pad  , \110(3)_pad  , \113(4)_pad  , \116(5)_pad  , \119(6)_pad  , \122(7)_pad  , \125(8)_pad  , \128(9)_pad  , \131(10)_pad  , \134(11)_pad  , \137(12)_pad  , \140(13)_pad  , \143(14)_pad  , \146(15)_pad  , \210(16)_pad  , \214(17)_pad  , \217(18)_pad  , \221(19)_pad  , \224(20)_pad  , \227(21)_pad  , \234(22)_pad  , \237(23)_pad  , \469(24)_pad  , \472(25)_pad  , \475(26)_pad  , \478(27)_pad  , \898(28)_pad  , \900(29)_pad  , \902(30)_pad  , \952(31)_pad  , \953(32)_pad  , \12(862)_pad  , \15(861)_pad  , \18(860)_pad  , \21(859)_pad  , \24(858)_pad  , \27(857)_pad  , \3(865)_pad  , \30(856)_pad  , \33(855)_pad  , \36(854)_pad  , \39(853)_pad  , \42(852)_pad  , \45(851)_pad  , \48(850)_pad  , \51(899)_pad  , \54(900)_pad  , \57(912)_pad  , \6(864)_pad  , \60(901)_pad  , \63(902)_pad  , \66(903)_pad  , \69(908)_pad  , \72(909)_pad  , \75(866)_pad  , \9(863)_pad  );
  input \101(0)_pad  ;
  input \104(1)_pad  ;
  input \107(2)_pad  ;
  input \110(3)_pad  ;
  input \113(4)_pad  ;
  input \116(5)_pad  ;
  input \119(6)_pad  ;
  input \122(7)_pad  ;
  input \125(8)_pad  ;
  input \128(9)_pad  ;
  input \131(10)_pad  ;
  input \134(11)_pad  ;
  input \137(12)_pad  ;
  input \140(13)_pad  ;
  input \143(14)_pad  ;
  input \146(15)_pad  ;
  input \210(16)_pad  ;
  input \214(17)_pad  ;
  input \217(18)_pad  ;
  input \221(19)_pad  ;
  input \224(20)_pad  ;
  input \227(21)_pad  ;
  input \234(22)_pad  ;
  input \237(23)_pad  ;
  input \469(24)_pad  ;
  input \472(25)_pad  ;
  input \475(26)_pad  ;
  input \478(27)_pad  ;
  input \898(28)_pad  ;
  input \900(29)_pad  ;
  input \902(30)_pad  ;
  input \952(31)_pad  ;
  input \953(32)_pad  ;
  output \12(862)_pad  ;
  output \15(861)_pad  ;
  output \18(860)_pad  ;
  output \21(859)_pad  ;
  output \24(858)_pad  ;
  output \27(857)_pad  ;
  output \3(865)_pad  ;
  output \30(856)_pad  ;
  output \33(855)_pad  ;
  output \36(854)_pad  ;
  output \39(853)_pad  ;
  output \42(852)_pad  ;
  output \45(851)_pad  ;
  output \48(850)_pad  ;
  output \51(899)_pad  ;
  output \54(900)_pad  ;
  output \57(912)_pad  ;
  output \6(864)_pad  ;
  output \60(901)_pad  ;
  output \63(902)_pad  ;
  output \66(903)_pad  ;
  output \69(908)_pad  ;
  output \72(909)_pad  ;
  output \75(866)_pad  ;
  output \9(863)_pad  ;
  wire n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 ;
  assign n34 = ~\143(14)_pad  & ~\146(15)_pad  ;
  assign n35 = \143(14)_pad  & \146(15)_pad  ;
  assign n36 = ~n34 & ~n35 ;
  assign n37 = ~\128(9)_pad  & n36 ;
  assign n38 = \128(9)_pad  & ~n36 ;
  assign n39 = ~n37 & ~n38 ;
  assign n40 = \131(10)_pad  & ~\134(11)_pad  ;
  assign n41 = ~\131(10)_pad  & \134(11)_pad  ;
  assign n42 = ~n40 & ~n41 ;
  assign n43 = \137(12)_pad  & ~n42 ;
  assign n44 = ~\137(12)_pad  & n42 ;
  assign n45 = ~n43 & ~n44 ;
  assign n46 = n39 & n45 ;
  assign n47 = ~n39 & ~n45 ;
  assign n48 = ~n46 & ~n47 ;
  assign n49 = \227(21)_pad  & ~\953(32)_pad  ;
  assign n50 = n48 & n49 ;
  assign n51 = ~n48 & ~n49 ;
  assign n52 = ~n50 & ~n51 ;
  assign n53 = ~\104(1)_pad  & ~\107(2)_pad  ;
  assign n54 = \104(1)_pad  & \107(2)_pad  ;
  assign n55 = ~n53 & ~n54 ;
  assign n56 = ~\110(3)_pad  & ~\140(13)_pad  ;
  assign n57 = \110(3)_pad  & \140(13)_pad  ;
  assign n58 = ~n56 & ~n57 ;
  assign n59 = \101(0)_pad  & ~n58 ;
  assign n60 = ~\101(0)_pad  & n58 ;
  assign n61 = ~n59 & ~n60 ;
  assign n62 = n55 & ~n61 ;
  assign n63 = ~n55 & n61 ;
  assign n64 = ~n62 & ~n63 ;
  assign n65 = ~\902(30)_pad  & ~n64 ;
  assign n66 = ~n52 & n65 ;
  assign n67 = ~\902(30)_pad  & n64 ;
  assign n68 = n52 & n67 ;
  assign n69 = ~n66 & ~n68 ;
  assign n70 = ~\469(24)_pad  & n69 ;
  assign n71 = \469(24)_pad  & ~\902(30)_pad  ;
  assign n72 = ~n64 & n71 ;
  assign n73 = ~n52 & n72 ;
  assign n74 = n64 & n71 ;
  assign n75 = n52 & n74 ;
  assign n76 = ~n73 & ~n75 ;
  assign n77 = \234(22)_pad  & ~\902(30)_pad  ;
  assign n78 = \221(19)_pad  & ~n77 ;
  assign n79 = n76 & ~n78 ;
  assign n80 = ~n70 & n79 ;
  assign n81 = ~\101(0)_pad  & ~\119(6)_pad  ;
  assign n82 = \101(0)_pad  & \119(6)_pad  ;
  assign n83 = ~n81 & ~n82 ;
  assign n84 = \113(4)_pad  & ~\116(5)_pad  ;
  assign n85 = ~\113(4)_pad  & \116(5)_pad  ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = n83 & n86 ;
  assign n88 = ~n83 & ~n86 ;
  assign n89 = ~n87 & ~n88 ;
  assign n90 = \110(3)_pad  & ~\122(7)_pad  ;
  assign n91 = ~\110(3)_pad  & \122(7)_pad  ;
  assign n92 = ~n90 & ~n91 ;
  assign n93 = n55 & ~n92 ;
  assign n94 = ~n55 & n92 ;
  assign n95 = ~n93 & ~n94 ;
  assign n96 = n89 & n95 ;
  assign n97 = ~n89 & ~n95 ;
  assign n98 = ~n96 & ~n97 ;
  assign n99 = \224(20)_pad  & ~\953(32)_pad  ;
  assign n100 = \125(8)_pad  & ~n99 ;
  assign n101 = ~\125(8)_pad  & n99 ;
  assign n102 = ~n100 & ~n101 ;
  assign n103 = n39 & ~n102 ;
  assign n104 = ~n39 & n102 ;
  assign n105 = ~n103 & ~n104 ;
  assign n106 = n98 & n105 ;
  assign n107 = ~n98 & ~n105 ;
  assign n108 = ~n106 & ~n107 ;
  assign n109 = ~\902(30)_pad  & n108 ;
  assign n110 = ~\237(23)_pad  & ~\902(30)_pad  ;
  assign n111 = \210(16)_pad  & ~n110 ;
  assign n112 = \214(17)_pad  & ~n110 ;
  assign n113 = n111 & ~n112 ;
  assign n114 = ~n109 & n113 ;
  assign n115 = ~n111 & ~n112 ;
  assign n116 = n109 & n115 ;
  assign n117 = ~n114 & ~n116 ;
  assign n118 = n80 & ~n117 ;
  assign n119 = ~\237(23)_pad  & ~\953(32)_pad  ;
  assign n120 = \210(16)_pad  & n119 ;
  assign n121 = ~\902(30)_pad  & ~n120 ;
  assign n122 = n89 & n121 ;
  assign n123 = ~n48 & n122 ;
  assign n124 = ~n89 & n121 ;
  assign n125 = n48 & n124 ;
  assign n126 = ~n123 & ~n125 ;
  assign n127 = ~\902(30)_pad  & n120 ;
  assign n128 = ~n89 & n127 ;
  assign n129 = ~n48 & n128 ;
  assign n130 = n89 & n127 ;
  assign n131 = n48 & n130 ;
  assign n132 = ~n129 & ~n131 ;
  assign n133 = n126 & n132 ;
  assign n134 = \472(25)_pad  & n133 ;
  assign n135 = ~\472(25)_pad  & ~n133 ;
  assign n136 = ~n134 & ~n135 ;
  assign n137 = ~\125(8)_pad  & ~\140(13)_pad  ;
  assign n138 = \125(8)_pad  & \140(13)_pad  ;
  assign n139 = ~n137 & ~n138 ;
  assign n140 = ~\146(15)_pad  & ~n139 ;
  assign n141 = \146(15)_pad  & n139 ;
  assign n142 = ~n140 & ~n141 ;
  assign n143 = ~\119(6)_pad  & ~\128(9)_pad  ;
  assign n144 = \119(6)_pad  & \128(9)_pad  ;
  assign n145 = ~n143 & ~n144 ;
  assign n146 = \110(3)_pad  & ~\137(12)_pad  ;
  assign n147 = ~\110(3)_pad  & \137(12)_pad  ;
  assign n148 = ~n146 & ~n147 ;
  assign n149 = \234(22)_pad  & ~\953(32)_pad  ;
  assign n150 = \221(19)_pad  & n149 ;
  assign n151 = n148 & n150 ;
  assign n152 = ~n145 & n151 ;
  assign n153 = ~n142 & n152 ;
  assign n154 = n148 & ~n150 ;
  assign n155 = n145 & n154 ;
  assign n156 = ~n142 & n155 ;
  assign n157 = ~n153 & ~n156 ;
  assign n158 = ~n145 & n154 ;
  assign n159 = n142 & n158 ;
  assign n160 = n145 & n151 ;
  assign n161 = n142 & n160 ;
  assign n162 = ~n159 & ~n161 ;
  assign n163 = n157 & n162 ;
  assign n164 = ~n148 & ~n150 ;
  assign n165 = ~n145 & n164 ;
  assign n166 = ~n142 & n165 ;
  assign n167 = ~n148 & n150 ;
  assign n168 = n145 & n167 ;
  assign n169 = ~n142 & n168 ;
  assign n170 = ~n166 & ~n169 ;
  assign n171 = ~n145 & n167 ;
  assign n172 = n142 & n171 ;
  assign n173 = n145 & n164 ;
  assign n174 = n142 & n173 ;
  assign n175 = ~n172 & ~n174 ;
  assign n176 = n170 & n175 ;
  assign n177 = n163 & n176 ;
  assign n178 = \217(18)_pad  & ~n77 ;
  assign n179 = ~\902(30)_pad  & ~n178 ;
  assign n180 = ~n177 & n179 ;
  assign n181 = ~\902(30)_pad  & ~n177 ;
  assign n182 = n178 & ~n181 ;
  assign n183 = ~n180 & ~n182 ;
  assign n184 = n136 & ~n183 ;
  assign n185 = \122(7)_pad  & ~\146(15)_pad  ;
  assign n186 = ~n139 & n185 ;
  assign n187 = \122(7)_pad  & \146(15)_pad  ;
  assign n188 = n139 & n187 ;
  assign n189 = ~n186 & ~n188 ;
  assign n190 = ~\122(7)_pad  & \146(15)_pad  ;
  assign n191 = ~n139 & n190 ;
  assign n192 = ~\122(7)_pad  & ~\146(15)_pad  ;
  assign n193 = n139 & n192 ;
  assign n194 = ~n191 & ~n193 ;
  assign n195 = n189 & n194 ;
  assign n196 = \214(17)_pad  & n119 ;
  assign n197 = ~\104(1)_pad  & ~\113(4)_pad  ;
  assign n198 = \104(1)_pad  & \113(4)_pad  ;
  assign n199 = ~n197 & ~n198 ;
  assign n200 = n196 & ~n199 ;
  assign n201 = ~n196 & n199 ;
  assign n202 = ~n200 & ~n201 ;
  assign n203 = \131(10)_pad  & ~\143(14)_pad  ;
  assign n204 = ~\131(10)_pad  & \143(14)_pad  ;
  assign n205 = ~n203 & ~n204 ;
  assign n206 = ~\902(30)_pad  & ~n205 ;
  assign n207 = ~n202 & n206 ;
  assign n208 = ~n195 & n207 ;
  assign n209 = ~\902(30)_pad  & n205 ;
  assign n210 = n202 & n209 ;
  assign n211 = ~n195 & n210 ;
  assign n212 = ~n208 & ~n211 ;
  assign n213 = ~n202 & n209 ;
  assign n214 = n195 & n213 ;
  assign n215 = n202 & n206 ;
  assign n216 = n195 & n215 ;
  assign n217 = ~n214 & ~n216 ;
  assign n218 = n212 & n217 ;
  assign n219 = ~\475(26)_pad  & ~n218 ;
  assign n220 = \475(26)_pad  & n218 ;
  assign n221 = ~n219 & ~n220 ;
  assign n222 = \217(18)_pad  & n149 ;
  assign n223 = ~\134(11)_pad  & ~\143(14)_pad  ;
  assign n224 = \134(11)_pad  & \143(14)_pad  ;
  assign n225 = ~n223 & ~n224 ;
  assign n226 = n222 & ~n225 ;
  assign n227 = ~n222 & n225 ;
  assign n228 = ~n226 & ~n227 ;
  assign n229 = ~\116(5)_pad  & ~\122(7)_pad  ;
  assign n230 = \116(5)_pad  & \122(7)_pad  ;
  assign n231 = ~n229 & ~n230 ;
  assign n232 = \107(2)_pad  & ~\128(9)_pad  ;
  assign n233 = ~\107(2)_pad  & \128(9)_pad  ;
  assign n234 = ~n232 & ~n233 ;
  assign n235 = n231 & ~n234 ;
  assign n236 = ~n231 & n234 ;
  assign n237 = ~n235 & ~n236 ;
  assign n238 = n228 & n237 ;
  assign n239 = ~n228 & ~n237 ;
  assign n240 = ~n238 & ~n239 ;
  assign n241 = \478(27)_pad  & ~\902(30)_pad  ;
  assign n242 = ~n240 & n241 ;
  assign n243 = ~\902(30)_pad  & ~n240 ;
  assign n244 = ~\478(27)_pad  & ~n243 ;
  assign n245 = ~n242 & ~n244 ;
  assign n246 = \234(22)_pad  & \237(23)_pad  ;
  assign n247 = \902(30)_pad  & \953(32)_pad  ;
  assign n248 = ~n246 & n247 ;
  assign n249 = ~\898(28)_pad  & n248 ;
  assign n250 = \952(31)_pad  & ~\953(32)_pad  ;
  assign n251 = ~n246 & n250 ;
  assign n252 = ~n249 & ~n251 ;
  assign n253 = ~n245 & ~n252 ;
  assign n254 = n221 & n253 ;
  assign n255 = n184 & n254 ;
  assign n256 = n118 & n255 ;
  assign n257 = \110(3)_pad  & ~n256 ;
  assign n258 = ~\110(3)_pad  & ~n117 ;
  assign n259 = n80 & n258 ;
  assign n260 = n255 & n259 ;
  assign n261 = ~n257 & ~n260 ;
  assign n262 = ~\469(24)_pad  & ~n78 ;
  assign n263 = n69 & n262 ;
  assign n264 = \469(24)_pad  & ~n78 ;
  assign n265 = ~n69 & n264 ;
  assign n266 = ~n263 & ~n265 ;
  assign n267 = ~n117 & ~n266 ;
  assign n268 = ~n221 & n253 ;
  assign n269 = ~n136 & n183 ;
  assign n270 = n268 & n269 ;
  assign n271 = n267 & n270 ;
  assign n272 = \113(4)_pad  & ~n271 ;
  assign n273 = ~\113(4)_pad  & n268 ;
  assign n274 = n269 & n273 ;
  assign n275 = n267 & n274 ;
  assign n276 = ~n272 & ~n275 ;
  assign n277 = n245 & ~n252 ;
  assign n278 = n221 & n277 ;
  assign n279 = n269 & n278 ;
  assign n280 = n267 & n279 ;
  assign n281 = \116(5)_pad  & ~n280 ;
  assign n282 = ~\116(5)_pad  & n278 ;
  assign n283 = n269 & n282 ;
  assign n284 = n267 & n283 ;
  assign n285 = ~n281 & ~n284 ;
  assign n286 = ~n136 & ~n183 ;
  assign n287 = n254 & n286 ;
  assign n288 = n267 & n287 ;
  assign n289 = \119(6)_pad  & ~n288 ;
  assign n290 = ~\119(6)_pad  & ~n117 ;
  assign n291 = ~n266 & n290 ;
  assign n292 = n287 & n291 ;
  assign n293 = ~n289 & ~n292 ;
  assign n294 = n136 & n183 ;
  assign n295 = ~n221 & n277 ;
  assign n296 = n294 & n295 ;
  assign n297 = n267 & n296 ;
  assign n298 = \122(7)_pad  & ~n297 ;
  assign n299 = ~\122(7)_pad  & ~n117 ;
  assign n300 = ~n266 & n299 ;
  assign n301 = n296 & n300 ;
  assign n302 = ~n298 & ~n301 ;
  assign n303 = ~\900(29)_pad  & n248 ;
  assign n304 = ~n251 & ~n303 ;
  assign n305 = ~n245 & ~n304 ;
  assign n306 = ~n221 & n305 ;
  assign n307 = n184 & n306 ;
  assign n308 = n267 & n307 ;
  assign n309 = \125(8)_pad  & ~n308 ;
  assign n310 = ~\125(8)_pad  & ~n117 ;
  assign n311 = ~n266 & n310 ;
  assign n312 = n307 & n311 ;
  assign n313 = ~n309 & ~n312 ;
  assign n314 = n254 & n269 ;
  assign n315 = n118 & n314 ;
  assign n316 = \101(0)_pad  & ~n315 ;
  assign n317 = ~\101(0)_pad  & n254 ;
  assign n318 = n269 & n317 ;
  assign n319 = n118 & n318 ;
  assign n320 = ~n316 & ~n319 ;
  assign n321 = n245 & ~n304 ;
  assign n322 = n221 & n321 ;
  assign n323 = n286 & n322 ;
  assign n324 = n118 & n323 ;
  assign n325 = \128(9)_pad  & ~n324 ;
  assign n326 = ~\128(9)_pad  & n322 ;
  assign n327 = n286 & n326 ;
  assign n328 = n118 & n327 ;
  assign n329 = ~n325 & ~n328 ;
  assign n330 = ~n109 & n111 ;
  assign n331 = ~\902(30)_pad  & ~n111 ;
  assign n332 = n108 & n331 ;
  assign n333 = ~n112 & ~n332 ;
  assign n334 = ~n330 & n333 ;
  assign n335 = n80 & n334 ;
  assign n336 = n269 & n306 ;
  assign n337 = n335 & n336 ;
  assign n338 = \131(10)_pad  & ~n337 ;
  assign n339 = ~\131(10)_pad  & n306 ;
  assign n340 = n269 & n339 ;
  assign n341 = n335 & n340 ;
  assign n342 = ~n338 & ~n341 ;
  assign n343 = n269 & n322 ;
  assign n344 = n335 & n343 ;
  assign n345 = \134(11)_pad  & ~n344 ;
  assign n346 = ~\134(11)_pad  & n322 ;
  assign n347 = n269 & n346 ;
  assign n348 = n335 & n347 ;
  assign n349 = ~n345 & ~n348 ;
  assign n350 = n221 & n305 ;
  assign n351 = n286 & n350 ;
  assign n352 = n335 & n351 ;
  assign n353 = \137(12)_pad  & ~n352 ;
  assign n354 = ~\137(12)_pad  & n334 ;
  assign n355 = n80 & n354 ;
  assign n356 = n351 & n355 ;
  assign n357 = ~n353 & ~n356 ;
  assign n358 = n307 & n335 ;
  assign n359 = \140(13)_pad  & ~n358 ;
  assign n360 = ~\140(13)_pad  & n306 ;
  assign n361 = n184 & n360 ;
  assign n362 = n335 & n361 ;
  assign n363 = ~n359 & ~n362 ;
  assign n364 = ~n221 & n321 ;
  assign n365 = n269 & n364 ;
  assign n366 = n118 & n365 ;
  assign n367 = \143(14)_pad  & ~n366 ;
  assign n368 = ~\143(14)_pad  & n364 ;
  assign n369 = n269 & n368 ;
  assign n370 = n118 & n369 ;
  assign n371 = ~n367 & ~n370 ;
  assign n372 = n286 & n306 ;
  assign n373 = n118 & n372 ;
  assign n374 = \146(15)_pad  & ~n373 ;
  assign n375 = ~\146(15)_pad  & n306 ;
  assign n376 = n286 & n375 ;
  assign n377 = n118 & n376 ;
  assign n378 = ~n374 & ~n377 ;
  assign n379 = ~n352 & ~n358 ;
  assign n380 = ~n366 & ~n373 ;
  assign n381 = n379 & n380 ;
  assign n382 = ~n308 & ~n324 ;
  assign n383 = ~n337 & ~n344 ;
  assign n384 = n382 & n383 ;
  assign n385 = n381 & n384 ;
  assign n386 = ~n297 & ~n315 ;
  assign n387 = n278 & n294 ;
  assign n388 = n118 & n387 ;
  assign n389 = n268 & n294 ;
  assign n390 = n118 & n389 ;
  assign n391 = ~n388 & ~n390 ;
  assign n392 = n386 & n391 ;
  assign n393 = ~n256 & ~n271 ;
  assign n394 = ~n280 & ~n288 ;
  assign n395 = n393 & n394 ;
  assign n396 = n392 & n395 ;
  assign n397 = n385 & n396 ;
  assign n398 = \210(16)_pad  & \902(30)_pad  ;
  assign n399 = ~n397 & n398 ;
  assign n400 = ~n108 & ~n399 ;
  assign n401 = ~\952(31)_pad  & \953(32)_pad  ;
  assign n402 = n108 & n398 ;
  assign n403 = ~n397 & n402 ;
  assign n404 = ~n401 & ~n403 ;
  assign n405 = ~n400 & n404 ;
  assign n406 = n52 & n64 ;
  assign n407 = ~n52 & ~n64 ;
  assign n408 = ~n406 & ~n407 ;
  assign n409 = \469(24)_pad  & \902(30)_pad  ;
  assign n410 = ~n397 & n409 ;
  assign n411 = n408 & ~n410 ;
  assign n412 = ~n408 & n409 ;
  assign n413 = ~n397 & n412 ;
  assign n414 = ~n401 & ~n413 ;
  assign n415 = ~n411 & n414 ;
  assign n416 = n89 & ~n120 ;
  assign n417 = ~n48 & n416 ;
  assign n418 = n89 & n120 ;
  assign n419 = n48 & n418 ;
  assign n420 = ~n417 & ~n419 ;
  assign n421 = ~n89 & n120 ;
  assign n422 = ~n48 & n421 ;
  assign n423 = ~n89 & ~n120 ;
  assign n424 = n48 & n423 ;
  assign n425 = ~n422 & ~n424 ;
  assign n426 = n420 & n425 ;
  assign n427 = \472(25)_pad  & \902(30)_pad  ;
  assign n428 = ~n397 & n427 ;
  assign n429 = n426 & ~n428 ;
  assign n430 = ~n426 & n427 ;
  assign n431 = ~n397 & n430 ;
  assign n432 = ~n401 & ~n431 ;
  assign n433 = ~n429 & n432 ;
  assign n434 = \104(1)_pad  & ~n390 ;
  assign n435 = ~\104(1)_pad  & n268 ;
  assign n436 = n294 & n435 ;
  assign n437 = n118 & n436 ;
  assign n438 = ~n434 & ~n437 ;
  assign n439 = n202 & n205 ;
  assign n440 = ~n195 & n439 ;
  assign n441 = n202 & ~n205 ;
  assign n442 = n195 & n441 ;
  assign n443 = ~n440 & ~n442 ;
  assign n444 = ~n202 & ~n205 ;
  assign n445 = ~n195 & n444 ;
  assign n446 = ~n202 & n205 ;
  assign n447 = n195 & n446 ;
  assign n448 = ~n445 & ~n447 ;
  assign n449 = n443 & n448 ;
  assign n450 = \475(26)_pad  & \902(30)_pad  ;
  assign n451 = ~n397 & n450 ;
  assign n452 = n449 & ~n451 ;
  assign n453 = ~n449 & n450 ;
  assign n454 = ~n397 & n453 ;
  assign n455 = ~n401 & ~n454 ;
  assign n456 = ~n452 & n455 ;
  assign n457 = \478(27)_pad  & \902(30)_pad  ;
  assign n458 = ~n397 & n457 ;
  assign n459 = n240 & ~n458 ;
  assign n460 = ~n240 & n457 ;
  assign n461 = ~n397 & n460 ;
  assign n462 = ~n401 & ~n461 ;
  assign n463 = ~n459 & n462 ;
  assign n464 = \217(18)_pad  & \902(30)_pad  ;
  assign n465 = ~n397 & n464 ;
  assign n466 = n177 & ~n465 ;
  assign n467 = ~n177 & n464 ;
  assign n468 = ~n397 & n467 ;
  assign n469 = ~n401 & ~n468 ;
  assign n470 = ~n466 & n469 ;
  assign n471 = ~\953(32)_pad  & ~n396 ;
  assign n472 = ~\224(20)_pad  & \953(32)_pad  ;
  assign n473 = n98 & ~n472 ;
  assign n474 = ~n471 & n473 ;
  assign n475 = ~\898(28)_pad  & \953(32)_pad  ;
  assign n476 = ~n98 & n472 ;
  assign n477 = ~\953(32)_pad  & ~n98 ;
  assign n478 = ~n396 & n477 ;
  assign n479 = ~n476 & ~n478 ;
  assign n480 = ~n475 & n479 ;
  assign n481 = ~n474 & n480 ;
  assign n482 = ~\953(32)_pad  & ~n385 ;
  assign n483 = ~\227(21)_pad  & \953(32)_pad  ;
  assign n484 = n48 & n139 ;
  assign n485 = ~n48 & ~n139 ;
  assign n486 = ~n484 & ~n485 ;
  assign n487 = ~n483 & n486 ;
  assign n488 = ~n482 & n487 ;
  assign n489 = ~\900(29)_pad  & \953(32)_pad  ;
  assign n490 = n486 & ~n489 ;
  assign n491 = ~n483 & ~n489 ;
  assign n492 = ~n482 & n491 ;
  assign n493 = ~n490 & ~n492 ;
  assign n494 = ~n488 & ~n493 ;
  assign n495 = n221 & ~n245 ;
  assign n496 = n334 & n495 ;
  assign n497 = ~n266 & n496 ;
  assign n498 = n294 & n497 ;
  assign n499 = ~\953(32)_pad  & ~n498 ;
  assign n500 = ~\952(31)_pad  & n499 ;
  assign n501 = n267 & n495 ;
  assign n502 = n266 & n334 ;
  assign n503 = n76 & n78 ;
  assign n504 = ~n70 & n503 ;
  assign n505 = n495 & ~n504 ;
  assign n506 = n502 & n505 ;
  assign n507 = ~n501 & ~n506 ;
  assign n508 = n221 & n245 ;
  assign n509 = ~n112 & n245 ;
  assign n510 = ~\475(26)_pad  & ~n112 ;
  assign n511 = n218 & n510 ;
  assign n512 = \475(26)_pad  & ~n112 ;
  assign n513 = ~n218 & n512 ;
  assign n514 = ~n511 & ~n513 ;
  assign n515 = ~n509 & n514 ;
  assign n516 = ~n508 & ~n515 ;
  assign n517 = ~n330 & ~n332 ;
  assign n518 = n112 & n245 ;
  assign n519 = \475(26)_pad  & n112 ;
  assign n520 = n218 & n519 ;
  assign n521 = ~\475(26)_pad  & n112 ;
  assign n522 = ~n218 & n521 ;
  assign n523 = ~n520 & ~n522 ;
  assign n524 = ~n518 & n523 ;
  assign n525 = n517 & n524 ;
  assign n526 = ~n266 & n525 ;
  assign n527 = ~n516 & n526 ;
  assign n528 = n294 & ~n527 ;
  assign n529 = n507 & n528 ;
  assign n530 = ~n294 & ~n497 ;
  assign n531 = n251 & ~n286 ;
  assign n532 = ~n530 & n531 ;
  assign n533 = ~n529 & n532 ;
  assign n534 = n499 & ~n533 ;
  assign n535 = n397 & n534 ;
  assign n536 = ~n500 & ~n535 ;
  assign n537 = \107(2)_pad  & ~n388 ;
  assign n538 = ~\107(2)_pad  & n278 ;
  assign n539 = n294 & n538 ;
  assign n540 = n118 & n539 ;
  assign n541 = ~n537 & ~n540 ;
  assign \12(862)_pad  = ~n261 ;
  assign \15(861)_pad  = ~n276 ;
  assign \18(860)_pad  = ~n285 ;
  assign \21(859)_pad  = ~n293 ;
  assign \24(858)_pad  = ~n302 ;
  assign \27(857)_pad  = ~n313 ;
  assign \3(865)_pad  = ~n320 ;
  assign \30(856)_pad  = ~n329 ;
  assign \33(855)_pad  = ~n342 ;
  assign \36(854)_pad  = ~n349 ;
  assign \39(853)_pad  = ~n357 ;
  assign \42(852)_pad  = ~n363 ;
  assign \45(851)_pad  = ~n371 ;
  assign \48(850)_pad  = ~n378 ;
  assign \51(899)_pad  = n405 ;
  assign \54(900)_pad  = n415 ;
  assign \57(912)_pad  = n433 ;
  assign \6(864)_pad  = ~n438 ;
  assign \60(901)_pad  = n456 ;
  assign \63(902)_pad  = n463 ;
  assign \66(903)_pad  = n470 ;
  assign \69(908)_pad  = ~n481 ;
  assign \72(909)_pad  = ~n494 ;
  assign \75(866)_pad  = n536 ;
  assign \9(863)_pad  = ~n541 ;
endmodule
