module top (\102GAT(31)_pad , \105GAT(32)_pad , \108GAT(33)_pad , \112GAT(34)_pad , \115GAT(35)_pad , \11GAT(3)_pad , \14GAT(4)_pad , \17GAT(5)_pad , \1GAT(0)_pad , \21GAT(6)_pad , \24GAT(7)_pad , \27GAT(8)_pad , \30GAT(9)_pad , \34GAT(10)_pad , \37GAT(11)_pad , \40GAT(12)_pad , \43GAT(13)_pad , \47GAT(14)_pad , \4GAT(1)_pad , \50GAT(15)_pad , \53GAT(16)_pad , \56GAT(17)_pad , \60GAT(18)_pad , \63GAT(19)_pad , \66GAT(20)_pad , \69GAT(21)_pad , \73GAT(22)_pad , \76GAT(23)_pad , \79GAT(24)_pad , \82GAT(25)_pad , \86GAT(26)_pad , \89GAT(27)_pad , \8GAT(2)_pad , \92GAT(28)_pad , \95GAT(29)_pad , \99GAT(30)_pad , \203GAT(82) , \309GAT(131) , \360GAT(162) , \421GAT(188)_pad , \430GAT(193)_pad , \431GAT(194)_pad , \432GAT(195)_pad );
	input \102GAT(31)_pad  ;
	input \105GAT(32)_pad  ;
	input \108GAT(33)_pad  ;
	input \112GAT(34)_pad  ;
	input \115GAT(35)_pad  ;
	input \11GAT(3)_pad  ;
	input \14GAT(4)_pad  ;
	input \17GAT(5)_pad  ;
	input \1GAT(0)_pad  ;
	input \21GAT(6)_pad  ;
	input \24GAT(7)_pad  ;
	input \27GAT(8)_pad  ;
	input \30GAT(9)_pad  ;
	input \34GAT(10)_pad  ;
	input \37GAT(11)_pad  ;
	input \40GAT(12)_pad  ;
	input \43GAT(13)_pad  ;
	input \47GAT(14)_pad  ;
	input \4GAT(1)_pad  ;
	input \50GAT(15)_pad  ;
	input \53GAT(16)_pad  ;
	input \56GAT(17)_pad  ;
	input \60GAT(18)_pad  ;
	input \63GAT(19)_pad  ;
	input \66GAT(20)_pad  ;
	input \69GAT(21)_pad  ;
	input \73GAT(22)_pad  ;
	input \76GAT(23)_pad  ;
	input \79GAT(24)_pad  ;
	input \82GAT(25)_pad  ;
	input \86GAT(26)_pad  ;
	input \89GAT(27)_pad  ;
	input \8GAT(2)_pad  ;
	input \92GAT(28)_pad  ;
	input \95GAT(29)_pad  ;
	input \99GAT(30)_pad  ;
	output \203GAT(82)  ;
	output \309GAT(131)  ;
	output \360GAT(162)  ;
	output \421GAT(188)_pad  ;
	output \430GAT(193)_pad  ;
	output \431GAT(194)_pad  ;
	output \432GAT(195)_pad  ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\89GAT(27)_pad ,
		\95GAT(29)_pad ,
		_w38_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1 (
		\11GAT(3)_pad ,
		\17GAT(5)_pad ,
		\1GAT(0)_pad ,
		\4GAT(1)_pad ,
		_w39_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		_w38_,
		_w39_,
		_w40_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3 (
		\24GAT(7)_pad ,
		\30GAT(9)_pad ,
		\50GAT(15)_pad ,
		\56GAT(17)_pad ,
		_w41_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4 (
		\102GAT(31)_pad ,
		\108GAT(33)_pad ,
		\63GAT(19)_pad ,
		\69GAT(21)_pad ,
		_w42_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name5 (
		\37GAT(11)_pad ,
		\43GAT(13)_pad ,
		\76GAT(23)_pad ,
		\82GAT(25)_pad ,
		_w43_
	);
	LUT3 #(
		.INIT('h80)
	) name6 (
		_w41_,
		_w42_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h7)
	) name7 (
		_w40_,
		_w44_,
		_w45_
	);
	LUT3 #(
		.INIT('h2a)
	) name8 (
		\76GAT(23)_pad ,
		_w40_,
		_w44_,
		_w46_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\82GAT(25)_pad ,
		\86GAT(26)_pad ,
		_w47_
	);
	LUT4 #(
		.INIT('h9500)
	) name10 (
		\76GAT(23)_pad ,
		_w40_,
		_w44_,
		_w47_,
		_w48_
	);
	LUT4 #(
		.INIT('hc444)
	) name11 (
		\37GAT(11)_pad ,
		\43GAT(13)_pad ,
		_w40_,
		_w44_,
		_w49_
	);
	LUT4 #(
		.INIT('hc444)
	) name12 (
		\63GAT(19)_pad ,
		\69GAT(21)_pad ,
		_w40_,
		_w44_,
		_w50_
	);
	LUT4 #(
		.INIT('h8caf)
	) name13 (
		\47GAT(14)_pad ,
		\73GAT(22)_pad ,
		_w49_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		_w48_,
		_w51_,
		_w52_
	);
	LUT4 #(
		.INIT('hc444)
	) name15 (
		\1GAT(0)_pad ,
		\4GAT(1)_pad ,
		_w40_,
		_w44_,
		_w53_
	);
	LUT4 #(
		.INIT('hc444)
	) name16 (
		\50GAT(15)_pad ,
		\56GAT(17)_pad ,
		_w40_,
		_w44_,
		_w54_
	);
	LUT4 #(
		.INIT('h8acf)
	) name17 (
		\60GAT(18)_pad ,
		\8GAT(2)_pad ,
		_w53_,
		_w54_,
		_w55_
	);
	LUT4 #(
		.INIT('hc444)
	) name18 (
		\89GAT(27)_pad ,
		\95GAT(29)_pad ,
		_w39_,
		_w44_,
		_w56_
	);
	LUT4 #(
		.INIT('hc444)
	) name19 (
		\24GAT(7)_pad ,
		\30GAT(9)_pad ,
		_w40_,
		_w44_,
		_w57_
	);
	LUT4 #(
		.INIT('h8acf)
	) name20 (
		\34GAT(10)_pad ,
		\99GAT(30)_pad ,
		_w56_,
		_w57_,
		_w58_
	);
	LUT4 #(
		.INIT('hc444)
	) name21 (
		\11GAT(3)_pad ,
		\17GAT(5)_pad ,
		_w40_,
		_w44_,
		_w59_
	);
	LUT4 #(
		.INIT('hc444)
	) name22 (
		\102GAT(31)_pad ,
		\108GAT(33)_pad ,
		_w40_,
		_w44_,
		_w60_
	);
	LUT4 #(
		.INIT('h8acf)
	) name23 (
		\112GAT(34)_pad ,
		\21GAT(6)_pad ,
		_w59_,
		_w60_,
		_w61_
	);
	LUT3 #(
		.INIT('h80)
	) name24 (
		_w55_,
		_w58_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h7)
	) name25 (
		_w52_,
		_w62_,
		_w63_
	);
	LUT4 #(
		.INIT('ha222)
	) name26 (
		\82GAT(25)_pad ,
		\86GAT(26)_pad ,
		_w52_,
		_w62_,
		_w64_
	);
	LUT4 #(
		.INIT('h2111)
	) name27 (
		\76GAT(23)_pad ,
		\92GAT(28)_pad ,
		_w40_,
		_w44_,
		_w65_
	);
	LUT4 #(
		.INIT('h7f00)
	) name28 (
		_w48_,
		_w52_,
		_w62_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w64_,
		_w66_,
		_w67_
	);
	LUT4 #(
		.INIT('hc444)
	) name30 (
		\99GAT(30)_pad ,
		_w56_,
		_w52_,
		_w62_,
		_w68_
	);
	LUT4 #(
		.INIT('hc444)
	) name31 (
		\60GAT(18)_pad ,
		_w54_,
		_w52_,
		_w62_,
		_w69_
	);
	LUT4 #(
		.INIT('h8caf)
	) name32 (
		\105GAT(32)_pad ,
		\66GAT(20)_pad ,
		_w68_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		_w67_,
		_w70_,
		_w71_
	);
	LUT4 #(
		.INIT('hc444)
	) name34 (
		\34GAT(10)_pad ,
		_w57_,
		_w52_,
		_w62_,
		_w72_
	);
	LUT4 #(
		.INIT('hc444)
	) name35 (
		\21GAT(6)_pad ,
		_w59_,
		_w52_,
		_w62_,
		_w73_
	);
	LUT4 #(
		.INIT('h8acf)
	) name36 (
		\27GAT(8)_pad ,
		\40GAT(12)_pad ,
		_w72_,
		_w73_,
		_w74_
	);
	LUT4 #(
		.INIT('hc444)
	) name37 (
		\73GAT(22)_pad ,
		_w50_,
		_w52_,
		_w62_,
		_w75_
	);
	LUT4 #(
		.INIT('hc444)
	) name38 (
		\112GAT(34)_pad ,
		_w60_,
		_w52_,
		_w62_,
		_w76_
	);
	LUT4 #(
		.INIT('h8acf)
	) name39 (
		\115GAT(35)_pad ,
		\79GAT(24)_pad ,
		_w75_,
		_w76_,
		_w77_
	);
	LUT4 #(
		.INIT('hc444)
	) name40 (
		\47GAT(14)_pad ,
		_w49_,
		_w52_,
		_w62_,
		_w78_
	);
	LUT4 #(
		.INIT('hc444)
	) name41 (
		\8GAT(2)_pad ,
		_w53_,
		_w52_,
		_w62_,
		_w79_
	);
	LUT4 #(
		.INIT('h8acf)
	) name42 (
		\14GAT(4)_pad ,
		\53GAT(16)_pad ,
		_w78_,
		_w79_,
		_w80_
	);
	LUT3 #(
		.INIT('h80)
	) name43 (
		_w74_,
		_w77_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h7)
	) name44 (
		_w71_,
		_w81_,
		_w82_
	);
	LUT4 #(
		.INIT('hc444)
	) name45 (
		\66GAT(20)_pad ,
		_w69_,
		_w71_,
		_w81_,
		_w83_
	);
	LUT4 #(
		.INIT('hc444)
	) name46 (
		\53GAT(16)_pad ,
		_w78_,
		_w71_,
		_w81_,
		_w84_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w83_,
		_w84_,
		_w85_
	);
	LUT4 #(
		.INIT('hc444)
	) name48 (
		\40GAT(12)_pad ,
		_w72_,
		_w71_,
		_w81_,
		_w86_
	);
	LUT4 #(
		.INIT('hc444)
	) name49 (
		\27GAT(8)_pad ,
		_w73_,
		_w71_,
		_w81_,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		_w86_,
		_w87_,
		_w88_
	);
	LUT4 #(
		.INIT('h0001)
	) name51 (
		_w83_,
		_w84_,
		_w86_,
		_w87_,
		_w89_
	);
	LUT4 #(
		.INIT('hfffe)
	) name52 (
		_w83_,
		_w84_,
		_w86_,
		_w87_,
		_w90_
	);
	LUT4 #(
		.INIT('hc444)
	) name53 (
		\105GAT(32)_pad ,
		_w68_,
		_w71_,
		_w81_,
		_w91_
	);
	LUT4 #(
		.INIT('hc444)
	) name54 (
		\115GAT(35)_pad ,
		_w76_,
		_w71_,
		_w81_,
		_w92_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		_w46_,
		_w64_,
		_w93_
	);
	LUT4 #(
		.INIT('hd500)
	) name56 (
		\92GAT(28)_pad ,
		_w71_,
		_w81_,
		_w93_,
		_w94_
	);
	LUT4 #(
		.INIT('hc444)
	) name57 (
		\79GAT(24)_pad ,
		_w75_,
		_w71_,
		_w81_,
		_w95_
	);
	LUT4 #(
		.INIT('h0001)
	) name58 (
		_w91_,
		_w92_,
		_w94_,
		_w95_,
		_w96_
	);
	LUT4 #(
		.INIT('hc444)
	) name59 (
		\14GAT(4)_pad ,
		_w79_,
		_w71_,
		_w81_,
		_w97_
	);
	LUT3 #(
		.INIT('h07)
	) name60 (
		_w89_,
		_w96_,
		_w97_,
		_w98_
	);
	LUT3 #(
		.INIT('h23)
	) name61 (
		_w86_,
		_w94_,
		_w95_,
		_w99_
	);
	LUT3 #(
		.INIT('h3b)
	) name62 (
		_w85_,
		_w88_,
		_w99_,
		_w100_
	);
	LUT4 #(
		.INIT('h2232)
	) name63 (
		_w84_,
		_w86_,
		_w91_,
		_w94_,
		_w101_
	);
	LUT4 #(
		.INIT('h0100)
	) name64 (
		_w83_,
		_w84_,
		_w86_,
		_w95_,
		_w102_
	);
	LUT3 #(
		.INIT('hfe)
	) name65 (
		_w87_,
		_w101_,
		_w102_,
		_w103_
	);
	assign \203GAT(82)  = _w45_ ;
	assign \309GAT(131)  = _w63_ ;
	assign \360GAT(162)  = _w82_ ;
	assign \421GAT(188)_pad  = _w98_ ;
	assign \430GAT(193)_pad  = _w90_ ;
	assign \431GAT(194)_pad  = _w100_ ;
	assign \432GAT(195)_pad  = _w103_ ;
endmodule;