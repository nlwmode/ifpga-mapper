module top (\dcnt_reg[0]/P0001 , \dcnt_reg[1]/P0001 , \dcnt_reg[2]/P0001 , \dcnt_reg[3]/P0001 , \key[0]_pad , \key[100]_pad , \key[101]_pad , \key[102]_pad , \key[103]_pad , \key[104]_pad , \key[105]_pad , \key[106]_pad , \key[107]_pad , \key[108]_pad , \key[109]_pad , \key[10]_pad , \key[110]_pad , \key[111]_pad , \key[112]_pad , \key[113]_pad , \key[114]_pad , \key[115]_pad , \key[116]_pad , \key[117]_pad , \key[118]_pad , \key[119]_pad , \key[11]_pad , \key[120]_pad , \key[121]_pad , \key[122]_pad , \key[123]_pad , \key[124]_pad , \key[125]_pad , \key[126]_pad , \key[127]_pad , \key[12]_pad , \key[13]_pad , \key[14]_pad , \key[15]_pad , \key[16]_pad , \key[17]_pad , \key[18]_pad , \key[19]_pad , \key[1]_pad , \key[20]_pad , \key[21]_pad , \key[22]_pad , \key[23]_pad , \key[24]_pad , \key[25]_pad , \key[26]_pad , \key[27]_pad , \key[28]_pad , \key[29]_pad , \key[2]_pad , \key[30]_pad , \key[31]_pad , \key[32]_pad , \key[33]_pad , \key[34]_pad , \key[35]_pad , \key[36]_pad , \key[37]_pad , \key[38]_pad , \key[39]_pad , \key[3]_pad , \key[40]_pad , \key[41]_pad , \key[42]_pad , \key[43]_pad , \key[44]_pad , \key[45]_pad , \key[46]_pad , \key[47]_pad , \key[48]_pad , \key[49]_pad , \key[4]_pad , \key[50]_pad , \key[51]_pad , \key[52]_pad , \key[53]_pad , \key[54]_pad , \key[55]_pad , \key[56]_pad , \key[57]_pad , \key[58]_pad , \key[59]_pad , \key[5]_pad , \key[60]_pad , \key[61]_pad , \key[62]_pad , \key[63]_pad , \key[64]_pad , \key[65]_pad , \key[66]_pad , \key[67]_pad , \key[68]_pad , \key[69]_pad , \key[6]_pad , \key[70]_pad , \key[71]_pad , \key[72]_pad , \key[73]_pad , \key[74]_pad , \key[75]_pad , \key[76]_pad , \key[77]_pad , \key[78]_pad , \key[79]_pad , \key[7]_pad , \key[80]_pad , \key[81]_pad , \key[82]_pad , \key[83]_pad , \key[84]_pad , \key[85]_pad , \key[86]_pad , \key[87]_pad , \key[88]_pad , \key[89]_pad , \key[8]_pad , \key[90]_pad , \key[91]_pad , \key[92]_pad , \key[93]_pad , \key[94]_pad , \key[95]_pad , \key[96]_pad , \key[97]_pad , \key[98]_pad , \key[99]_pad , \key[9]_pad , ld_pad, \ld_r_reg/P0001 , rst_pad, \sa00_reg[0]/P0001 , \sa00_reg[1]/P0001 , \sa00_reg[2]/P0001 , \sa00_reg[3]/P0001 , \sa00_reg[4]/P0001 , \sa00_reg[5]/P0001 , \sa00_reg[6]/NET0131 , \sa00_reg[7]/NET0131 , \sa01_reg[0]/P0001 , \sa01_reg[1]/P0001 , \sa01_reg[2]/P0001 , \sa01_reg[3]/P0001 , \sa01_reg[4]/P0001 , \sa01_reg[5]/P0001 , \sa01_reg[6]/NET0131 , \sa01_reg[7]/NET0131 , \sa02_reg[0]/P0001 , \sa02_reg[1]/P0001 , \sa02_reg[2]/P0001 , \sa02_reg[3]/P0001 , \sa02_reg[4]/P0001 , \sa02_reg[5]/P0001 , \sa02_reg[6]/NET0131 , \sa02_reg[7]/NET0131 , \sa03_reg[0]/P0001 , \sa03_reg[1]/P0001 , \sa03_reg[2]/P0001 , \sa03_reg[3]/P0001 , \sa03_reg[4]/P0001 , \sa03_reg[5]/P0001 , \sa03_reg[6]/NET0131 , \sa03_reg[7]/NET0131 , \sa10_reg[0]/P0001 , \sa10_reg[1]/P0001 , \sa10_reg[2]/P0001 , \sa10_reg[3]/P0001 , \sa10_reg[4]/P0001 , \sa10_reg[5]/P0001 , \sa10_reg[6]/NET0131 , \sa10_reg[7]/NET0131 , \sa11_reg[0]/P0001 , \sa11_reg[1]/P0001 , \sa11_reg[2]/P0001 , \sa11_reg[3]/P0001 , \sa11_reg[4]/P0001 , \sa11_reg[5]/P0001 , \sa11_reg[6]/NET0131 , \sa11_reg[7]/NET0131 , \sa12_reg[0]/P0001 , \sa12_reg[1]/P0001 , \sa12_reg[2]/P0001 , \sa12_reg[3]/P0001 , \sa12_reg[4]/P0001 , \sa12_reg[5]/P0001 , \sa12_reg[6]/NET0131 , \sa12_reg[7]/NET0131 , \sa13_reg[0]/P0001 , \sa13_reg[1]/P0001 , \sa13_reg[2]/P0001 , \sa13_reg[3]/P0001 , \sa13_reg[4]/P0001 , \sa13_reg[5]/P0001 , \sa13_reg[6]/NET0131 , \sa13_reg[7]/NET0131 , \sa20_reg[0]/P0001 , \sa20_reg[1]/P0001 , \sa20_reg[2]/P0001 , \sa20_reg[3]/P0001 , \sa20_reg[4]/P0001 , \sa20_reg[5]/P0001 , \sa20_reg[6]/NET0131 , \sa20_reg[7]/NET0131 , \sa21_reg[0]/P0001 , \sa21_reg[1]/P0001 , \sa21_reg[2]/P0001 , \sa21_reg[3]/P0001 , \sa21_reg[4]/P0001 , \sa21_reg[5]/P0001 , \sa21_reg[6]/NET0131 , \sa21_reg[7]/P0001 , \sa22_reg[0]/P0001 , \sa22_reg[1]/P0001 , \sa22_reg[2]/P0001 , \sa22_reg[3]/P0001 , \sa22_reg[4]/P0001 , \sa22_reg[5]/P0001 , \sa22_reg[6]/NET0131 , \sa22_reg[7]/NET0131 , \sa23_reg[0]/P0001 , \sa23_reg[1]/P0001 , \sa23_reg[2]/P0001 , \sa23_reg[3]/P0001 , \sa23_reg[4]/P0001 , \sa23_reg[5]/P0001 , \sa23_reg[6]/NET0131 , \sa23_reg[7]/NET0131 , \sa30_reg[0]/P0002 , \sa30_reg[1]/P0001 , \sa30_reg[2]/P0001 , \sa30_reg[3]/P0001 , \sa30_reg[4]/P0001 , \sa30_reg[5]/P0001 , \sa30_reg[6]/NET0131 , \sa30_reg[7]/P0001 , \sa31_reg[0]/P0002 , \sa31_reg[1]/P0001 , \sa31_reg[2]/P0001 , \sa31_reg[3]/P0001 , \sa31_reg[4]/P0001 , \sa31_reg[5]/P0001 , \sa31_reg[6]/NET0131 , \sa31_reg[7]/P0001 , \sa32_reg[0]/P0002 , \sa32_reg[1]/P0001 , \sa32_reg[2]/P0001 , \sa32_reg[3]/P0001 , \sa32_reg[4]/P0001 , \sa32_reg[5]/P0001 , \sa32_reg[6]/NET0131 , \sa32_reg[7]/P0001 , \sa33_reg[0]/P0001 , \sa33_reg[1]/P0001 , \sa33_reg[2]/P0001 , \sa33_reg[3]/P0001 , \sa33_reg[4]/P0001 , \sa33_reg[5]/P0001 , \sa33_reg[6]/P0001 , \sa33_reg[7]/NET0131 , \text_in_r_reg[0]/P0001 , \text_in_r_reg[100]/P0001 , \text_in_r_reg[101]/P0001 , \text_in_r_reg[102]/P0001 , \text_in_r_reg[103]/P0001 , \text_in_r_reg[104]/P0001 , \text_in_r_reg[105]/P0001 , \text_in_r_reg[106]/P0001 , \text_in_r_reg[107]/P0001 , \text_in_r_reg[108]/P0001 , \text_in_r_reg[109]/P0001 , \text_in_r_reg[10]/P0001 , \text_in_r_reg[110]/P0001 , \text_in_r_reg[111]/P0001 , \text_in_r_reg[112]/P0001 , \text_in_r_reg[113]/P0001 , \text_in_r_reg[114]/P0001 , \text_in_r_reg[115]/P0001 , \text_in_r_reg[116]/P0001 , \text_in_r_reg[117]/P0001 , \text_in_r_reg[118]/P0001 , \text_in_r_reg[119]/P0001 , \text_in_r_reg[11]/P0001 , \text_in_r_reg[120]/P0001 , \text_in_r_reg[121]/P0001 , \text_in_r_reg[122]/P0001 , \text_in_r_reg[123]/P0001 , \text_in_r_reg[124]/P0001 , \text_in_r_reg[125]/P0001 , \text_in_r_reg[126]/P0001 , \text_in_r_reg[127]/P0001 , \text_in_r_reg[12]/P0001 , \text_in_r_reg[13]/P0001 , \text_in_r_reg[14]/P0001 , \text_in_r_reg[15]/P0001 , \text_in_r_reg[16]/P0001 , \text_in_r_reg[17]/P0001 , \text_in_r_reg[18]/P0001 , \text_in_r_reg[19]/P0001 , \text_in_r_reg[1]/P0001 , \text_in_r_reg[20]/P0001 , \text_in_r_reg[21]/P0001 , \text_in_r_reg[22]/P0001 , \text_in_r_reg[23]/P0001 , \text_in_r_reg[24]/P0001 , \text_in_r_reg[25]/P0001 , \text_in_r_reg[26]/P0001 , \text_in_r_reg[27]/P0001 , \text_in_r_reg[28]/P0001 , \text_in_r_reg[29]/P0001 , \text_in_r_reg[2]/P0001 , \text_in_r_reg[30]/P0001 , \text_in_r_reg[31]/P0001 , \text_in_r_reg[32]/P0001 , \text_in_r_reg[33]/P0001 , \text_in_r_reg[34]/P0001 , \text_in_r_reg[35]/P0001 , \text_in_r_reg[36]/P0001 , \text_in_r_reg[37]/P0001 , \text_in_r_reg[38]/P0001 , \text_in_r_reg[39]/P0001 , \text_in_r_reg[3]/P0001 , \text_in_r_reg[40]/P0001 , \text_in_r_reg[41]/P0001 , \text_in_r_reg[42]/P0001 , \text_in_r_reg[43]/P0001 , \text_in_r_reg[44]/P0001 , \text_in_r_reg[45]/P0001 , \text_in_r_reg[46]/P0001 , \text_in_r_reg[47]/P0001 , \text_in_r_reg[48]/P0001 , \text_in_r_reg[49]/P0001 , \text_in_r_reg[4]/P0001 , \text_in_r_reg[50]/P0001 , \text_in_r_reg[51]/P0001 , \text_in_r_reg[52]/P0001 , \text_in_r_reg[53]/P0001 , \text_in_r_reg[54]/P0001 , \text_in_r_reg[55]/P0001 , \text_in_r_reg[56]/P0001 , \text_in_r_reg[57]/P0001 , \text_in_r_reg[58]/P0001 , \text_in_r_reg[59]/P0001 , \text_in_r_reg[5]/P0001 , \text_in_r_reg[60]/P0001 , \text_in_r_reg[61]/P0001 , \text_in_r_reg[62]/P0001 , \text_in_r_reg[63]/P0001 , \text_in_r_reg[64]/P0001 , \text_in_r_reg[65]/P0001 , \text_in_r_reg[66]/P0001 , \text_in_r_reg[67]/P0001 , \text_in_r_reg[68]/P0001 , \text_in_r_reg[69]/P0001 , \text_in_r_reg[6]/P0001 , \text_in_r_reg[70]/P0001 , \text_in_r_reg[71]/P0001 , \text_in_r_reg[72]/P0001 , \text_in_r_reg[73]/P0001 , \text_in_r_reg[74]/P0001 , \text_in_r_reg[75]/P0001 , \text_in_r_reg[76]/P0001 , \text_in_r_reg[77]/P0001 , \text_in_r_reg[78]/P0001 , \text_in_r_reg[79]/P0001 , \text_in_r_reg[7]/P0001 , \text_in_r_reg[80]/P0001 , \text_in_r_reg[81]/P0001 , \text_in_r_reg[82]/P0001 , \text_in_r_reg[83]/P0001 , \text_in_r_reg[84]/P0001 , \text_in_r_reg[85]/P0001 , \text_in_r_reg[86]/P0001 , \text_in_r_reg[87]/P0001 , \text_in_r_reg[88]/P0001 , \text_in_r_reg[89]/P0001 , \text_in_r_reg[8]/P0001 , \text_in_r_reg[90]/P0001 , \text_in_r_reg[91]/P0001 , \text_in_r_reg[92]/P0001 , \text_in_r_reg[93]/P0001 , \text_in_r_reg[94]/P0001 , \text_in_r_reg[95]/P0001 , \text_in_r_reg[96]/P0001 , \text_in_r_reg[97]/P0001 , \text_in_r_reg[98]/P0001 , \text_in_r_reg[99]/P0001 , \text_in_r_reg[9]/P0001 , \u0_r0_out_reg[24]/P0001 , \u0_r0_out_reg[25]/P0001 , \u0_r0_out_reg[26]/P0001 , \u0_r0_out_reg[27]/P0001 , \u0_r0_out_reg[28]/P0001 , \u0_r0_out_reg[29]/P0001 , \u0_r0_out_reg[30]/P0001 , \u0_r0_out_reg[31]/P0001 , \u0_r0_rcnt_reg[0]/P0001 , \u0_r0_rcnt_reg[1]/P0001 , \u0_r0_rcnt_reg[2]/P0001 , \u0_r0_rcnt_reg[3]/P0001 , \u0_w_reg[0][0]/P0001 , \u0_w_reg[0][10]/P0001 , \u0_w_reg[0][11]/P0001 , \u0_w_reg[0][12]/P0001 , \u0_w_reg[0][13]/P0001 , \u0_w_reg[0][14]/P0001 , \u0_w_reg[0][15]/P0001 , \u0_w_reg[0][16]/P0001 , \u0_w_reg[0][17]/P0001 , \u0_w_reg[0][18]/P0001 , \u0_w_reg[0][19]/P0001 , \u0_w_reg[0][1]/P0001 , \u0_w_reg[0][20]/P0001 , \u0_w_reg[0][21]/P0001 , \u0_w_reg[0][22]/P0001 , \u0_w_reg[0][23]/P0001 , \u0_w_reg[0][24]/P0001 , \u0_w_reg[0][25]/P0001 , \u0_w_reg[0][26]/P0001 , \u0_w_reg[0][27]/P0001 , \u0_w_reg[0][28]/P0001 , \u0_w_reg[0][29]/P0001 , \u0_w_reg[0][2]/P0001 , \u0_w_reg[0][30]/P0001 , \u0_w_reg[0][31]/P0001 , \u0_w_reg[0][3]/P0001 , \u0_w_reg[0][4]/P0001 , \u0_w_reg[0][5]/P0001 , \u0_w_reg[0][6]/P0001 , \u0_w_reg[0][7]/P0001 , \u0_w_reg[0][8]/P0001 , \u0_w_reg[0][9]/P0001 , \u0_w_reg[1][0]/P0001 , \u0_w_reg[1][10]/P0001 , \u0_w_reg[1][11]/P0001 , \u0_w_reg[1][12]/P0001 , \u0_w_reg[1][13]/P0001 , \u0_w_reg[1][14]/P0001 , \u0_w_reg[1][15]/P0001 , \u0_w_reg[1][16]/P0001 , \u0_w_reg[1][17]/P0001 , \u0_w_reg[1][18]/P0001 , \u0_w_reg[1][19]/P0001 , \u0_w_reg[1][1]/P0001 , \u0_w_reg[1][20]/P0001 , \u0_w_reg[1][21]/P0001 , \u0_w_reg[1][22]/P0001 , \u0_w_reg[1][23]/P0001 , \u0_w_reg[1][24]/P0002 , \u0_w_reg[1][25]/P0001 , \u0_w_reg[1][26]/P0001 , \u0_w_reg[1][27]/P0001 , \u0_w_reg[1][28]/P0001 , \u0_w_reg[1][29]/P0002 , \u0_w_reg[1][2]/P0001 , \u0_w_reg[1][30]/P0001 , \u0_w_reg[1][31]/P0001 , \u0_w_reg[1][3]/P0001 , \u0_w_reg[1][4]/P0001 , \u0_w_reg[1][5]/P0001 , \u0_w_reg[1][6]/P0001 , \u0_w_reg[1][7]/P0001 , \u0_w_reg[1][8]/P0001 , \u0_w_reg[1][9]/P0001 , \u0_w_reg[2][0]/P0001 , \u0_w_reg[2][10]/P0001 , \u0_w_reg[2][11]/P0001 , \u0_w_reg[2][12]/P0001 , \u0_w_reg[2][13]/P0001 , \u0_w_reg[2][14]/P0001 , \u0_w_reg[2][15]/P0001 , \u0_w_reg[2][16]/P0001 , \u0_w_reg[2][17]/P0001 , \u0_w_reg[2][18]/P0001 , \u0_w_reg[2][19]/P0001 , \u0_w_reg[2][1]/P0001 , \u0_w_reg[2][20]/P0001 , \u0_w_reg[2][21]/P0001 , \u0_w_reg[2][22]/P0001 , \u0_w_reg[2][23]/P0001 , \u0_w_reg[2][24]/P0001 , \u0_w_reg[2][25]/P0001 , \u0_w_reg[2][26]/P0001 , \u0_w_reg[2][27]/P0001 , \u0_w_reg[2][28]/P0001 , \u0_w_reg[2][29]/P0001 , \u0_w_reg[2][2]/P0001 , \u0_w_reg[2][30]/P0001 , \u0_w_reg[2][31]/P0001 , \u0_w_reg[2][3]/P0001 , \u0_w_reg[2][4]/P0001 , \u0_w_reg[2][5]/P0001 , \u0_w_reg[2][6]/P0001 , \u0_w_reg[2][7]/P0001 , \u0_w_reg[2][8]/P0001 , \u0_w_reg[2][9]/P0001 , \u0_w_reg[3][0]/P0001 , \u0_w_reg[3][10]/P0001 , \u0_w_reg[3][11]/P0001 , \u0_w_reg[3][12]/P0001 , \u0_w_reg[3][13]/P0001 , \u0_w_reg[3][14]/P0001 , \u0_w_reg[3][15]/P0001 , \u0_w_reg[3][16]/P0001 , \u0_w_reg[3][17]/P0001 , \u0_w_reg[3][18]/P0001 , \u0_w_reg[3][19]/P0001 , \u0_w_reg[3][1]/P0001 , \u0_w_reg[3][20]/P0001 , \u0_w_reg[3][21]/P0001 , \u0_w_reg[3][22]/P0001 , \u0_w_reg[3][23]/P0001 , \u0_w_reg[3][24]/P0001 , \u0_w_reg[3][25]/P0001 , \u0_w_reg[3][26]/P0001 , \u0_w_reg[3][27]/P0001 , \u0_w_reg[3][28]/P0001 , \u0_w_reg[3][29]/P0001 , \u0_w_reg[3][2]/P0001 , \u0_w_reg[3][30]/P0001 , \u0_w_reg[3][31]/P0001 , \u0_w_reg[3][3]/P0001 , \u0_w_reg[3][4]/P0001 , \u0_w_reg[3][5]/P0001 , \u0_w_reg[3][6]/P0001 , \u0_w_reg[3][7]/P0001 , \u0_w_reg[3][8]/P0001 , \u0_w_reg[3][9]/P0001 , \_al_n0 , \_al_n1 , \g21/_0_ , \g56610/_0_ , \g56611/_0_ , \g56612/_0_ , \g56613/_0_ , \g56614/_0_ , \g56615/_0_ , \g56616/_0_ , \g56617/_0_ , \g56630/_0_ , \g56631/_0_ , \g56632/_0_ , \g56633/_0_ , \g56634/_0_ , \g56635/_0_ , \g56645/_0_ , \g56646/_0_ , \g56647/_0_ , \g56648/_0_ , \g56649/_0_ , \g56650/_0_ , \g56651/_0_ , \g56652/_0_ , \g56666/_0_ , \g56667/_0_ , \g56668/_0_ , \g56669/_0_ , \g56670/_0_ , \g56671/_0_ , \g56672/_0_ , \g56674/_0_ , \g56675/_0_ , \g56704/_0_ , \g56739/_0_ , \g56743/_0_ , \g56763/_0_ , \g56776/_0_ , \g56812/_0_ , \g56818/_0_ , \g56861/_0_ , \g56874/_0_ , \g56919/_0_ , \g56920/_0_ , \g56921/_0_ , \g56923/_0_ , \g56924/_0_ , \g56925/_0_ , \g56926/_0_ , \g56956/_0_ , \g56957/_0_ , \g56958/_0_ , \g56959/_0_ , \g56960/_0_ , \g56961/_0_ , \g56972/_0_ , \g56973/_0_ , \g56974/_0_ , \g56976/_0_ , \g56977/_0_ , \g56978/_0_ , \g56979/_0_ , \g56980/_0_ , \g57008/_0_ , \g57010/_0_ , \g57011/_0_ , \g57012/_0_ , \g57013/_0_ , \g57014/_0_ , \g57015/_0_ , \g57016/_0_ , \g57017/_0_ , \g57086/_0_ , \g57091/_0_ , \g57114/_0_ , \g57129/_0_ , \g57163/_0_ , \g57171/_0_ , \g57204/_0_ , \g57218/_0_ , \g57262/_0_ , \g57263/_0_ , \g57264/_0_ , \g57265/_0_ , \g57266/_0_ , \g57267/_0_ , \g57268/_0_ , \g57269/_0_ , \g57300/_0_ , \g57301/_0_ , \g57302/_0_ , \g57303/_0_ , \g57304/_0_ , \g57316/_0_ , \g57317/_0_ , \g57319/_0_ , \g57320/_0_ , \g57321/_0_ , \g57322/_0_ , \g57323/_0_ , \g57324/_0_ , \g57350/_0_ , \g57353/_0_ , \g57354/_0_ , \g57355/_0_ , \g57356/_0_ , \g57357/_0_ , \g57358/_0_ , \g57359/_0_ , \g57360/_0_ , \g57427/_0_ , \g57432/_0_ , \g57456/_0_ , \g57471/_0_ , \g57506/_0_ , \g57512/_0_ , \g57540/_0_ , \g57547/_0_ , \g57654/_0_ , \g57655/_0_ , \g57656/_0_ , \g57657/_0_ , \g57658/_0_ , \g57676/_0_ , \g57677/_0_ , \g57678/_0_ , \g57679/_0_ , \g57680/_0_ , \g57681/_0_ , \g57682/_0_ , \g57683/_0_ , \g57684/_0_ , \g57685/_0_ , \g57686/_0_ , \g57687/_0_ , \g57688/_0_ , \g57689/_0_ , \g57690/_0_ , \g57691/_0_ , \g57700/_0_ , \g57701/_0_ , \g57702/_0_ , \g57703/_0_ , \g57704/_0_ , \g57705/_0_ , \g57706/_0_ , \g57707/_0_ , \g57708/_0_ , \g57709/_3_ , \g57710/_3_ , \g57711/_0_ , \g57712/_3_ , \g57715/_3_ , \g57716/_3_ , \g57767/_0_ , \g57768/_3_ , \g57769/_3_ , \g57770/_3_ , \g57771/_3_ , \g57777/_3_ , \g57779/_3_ , \g57804/_3_ , \g57805/_3_ , \g57806/_3_ , \g57807/_3_ , \g57808/_3_ , \g57809/_3_ , \g57810/_3_ , \g57811/_3_ , \g57812/_3_ , \g57813/_3_ , \g57814/_3_ , \g57815/_3_ , \g57816/_0_ , \g57817/_3_ , \g57818/_3_ , \g57819/_3_ , \g57822/_3_ , \g57823/_3_ , \g57824/_3_ , \g57830/_3_ , \g57835/_3_ , \g57836/_3_ , \g57837/_3_ , \g57841/_3_ , \g57842/_3_ , \g57843/_3_ , \g57854/_3_ , \g57855/_3_ , \g57856/_3_ , \g57857/_3_ , \g57858/_3_ , \g57859/_3_ , \g57860/_3_ , \g57861/_3_ , \g57871/_3_ , \g57872/_3_ , \g57874/_3_ , \g57968/_3_ , \g57969/_3_ , \g57970/_3_ , \g57971/_3_ , \g57980/_3_ , \g57983/_3_ , \g57984/_3_ , \g57985/_3_ , \g58012/_3_ , \g58013/_3_ , \g58015/_3_ , \g58057/_3_ , \g58058/_3_ , \g58059/_3_ , \g58189/_3_ , \g58190/_3_ , \g58191/_3_ , \g58192/_3_ , \g58193/_3_ , \g58194/_3_ , \g58195/_3_ , \g58196/_3_ , \g58197/_3_ , \g58224/_3_ , \g58226/_3_ , \g58229/_3_ , \g58255/_3_ , \g58256/_3_ , \g58257/_3_ , \g58258/_3_ , \g58259/_3_ , \g58260/_3_ , \g58261/_3_ , \g58262/_3_ , \g58263/_3_ , \g58264/_3_ , \g58265/_3_ , \g58266/_3_ , \g58267/_3_ , \g58268/_3_ , \g58269/_3_ , \g58270/_0_ , \g58271/_3_ , \g58272/_3_ , \g58273/_3_ , \g58274/_3_ , \g58275/_3_ , \g58276/_3_ , \g58277/_3_ , \g58278/_3_ , \g58279/_3_ , \g58285/_3_ , \g58286/_3_ , \g58288/_3_ , \g58289/_3_ , \g58290/_3_ , \g58292/_3_ , \g58294/_3_ , \g58295/_3_ , \g58297/_3_ , \g58330/_0_ , \g58331/_0_ , \g58332/_0_ , \g58333/_0_ , \g58444/_3_ , \g58445/_3_ , \g58446/_3_ , \g58462/_0_ , \g58506/_0_ , \g58507/_0_ , \g58508/_0_ , \g58509/_0_ , \g58531/_0_ , \g58532/_0_ , \g58533/_0_ , \g58550/_0_ , \g58551/_0_ , \g58552/_0_ , \g58553/_0_ , \g58554/_0_ , \g58555/_0_ , \g58556/_0_ , \g58557/_0_ , \g58558/_0_ , \g58559/_0_ , \g58560/_0_ , \g58600/_3_ , \g58601/_3_ , \g58602/_3_ , \g58603/_3_ , \g58604/_3_ , \g58605/_3_ , \g58606/_3_ , \g58607/_3_ , \g58608/_3_ , \g58611/_0_ , \g58612/_0_ , \g58613/_0_ , \g58614/_0_ , \g58617/_0_ , \g58618/_0_ , \g58619/_0_ , \g58634/_0_ , \g58635/_0_ , \g58636/_0_ , \g58637/_0_ , \g58638/_0_ , \g58639/_0_ , \g58640/_0_ , \g58641/_0_ , \g58829/_3_ , \g58830/_3_ , \g58831/_3_ , \g58832/_3_ , \g58833/_3_ , \g58834/_3_ , \g58835/_0_ , \g58844/_0_ , \g58902/_0_ , \g58903/_0_ , \g58904/_0_ , \g58905/_0_ , \g58910/_0_ , \g58913/_0_ , \g58934/_0_ , \g58935/_0_ , \g58936/_0_ , \g58937/_0_ , \g58938/_0_ , \g58970/_0_ , \g58972/_0_ , \g58994/_0_ , \g58995/_0_ , \g58996/_0_ , \g58997/_0_ , \g58998/_0_ , \g58999/_0_ , \g59000/_0_ , \g59002/_0_ , \g59003/_0_ , \g59004/_0_ , \g59254/_0_ , \g59257/_0_ , \g59258/_0_ , \g59259/_0_ , \g59276/_0_ , \g59277/_0_ , \g59278/_0_ , \g59279/_0_ , \g59280/_0_ , \g59291/_0_ , \g59292/_0_ , \g59293/_0_ , \g59294/_0_ , \g59295/_0_ , \g59308/_0_ , \g59309/_0_ , \g59310/_0_ , \g59311/_0_ , \g59330/_0_ , \g59331/_0_ , \g59332/_0_ , \g59333/_0_ , \g59334/_0_ , \g59335/_0_ , \g59336/_0_ , \g59337/_0_ , \g59338/_0_ , \g59339/_0_ , \g59596/_0_ , \g59597/_0_ , \g59598/_0_ , \g59599/_0_ , \g59625/_0_ , \g59626/_0_ , \g59627/_0_ , \g59628/_0_ , \g59837/_0_ , \g59838/_0_ , \g59839/_0_ , \g59840/_0_ , \g60090/_0_ , \g60320/_0_ , \g60321/_0_ , \g60409/_0_ , \g60539/_0_ , \g60860/_0_ , \g60977/_0_ , \g61012/_0_ , \g61185/_0_ , \g61524/_2_ , \g61776/_0_ , \g61895/_0_ , \g61897/_0_ , \g62220/_0_ , \g65958/_0_ , \g72347/_3_ , \g77848/_0_ , \g85056/_0_ , \sa30_reg[0]/_05_ , \sa31_reg[0]/_05_ , \sa32_reg[0]/_05_ , \u0_w_reg[1][24]/_05_ , \u0_w_reg[1][29]/_05_ );
	input \dcnt_reg[0]/P0001  ;
	input \dcnt_reg[1]/P0001  ;
	input \dcnt_reg[2]/P0001  ;
	input \dcnt_reg[3]/P0001  ;
	input \key[0]_pad  ;
	input \key[100]_pad  ;
	input \key[101]_pad  ;
	input \key[102]_pad  ;
	input \key[103]_pad  ;
	input \key[104]_pad  ;
	input \key[105]_pad  ;
	input \key[106]_pad  ;
	input \key[107]_pad  ;
	input \key[108]_pad  ;
	input \key[109]_pad  ;
	input \key[10]_pad  ;
	input \key[110]_pad  ;
	input \key[111]_pad  ;
	input \key[112]_pad  ;
	input \key[113]_pad  ;
	input \key[114]_pad  ;
	input \key[115]_pad  ;
	input \key[116]_pad  ;
	input \key[117]_pad  ;
	input \key[118]_pad  ;
	input \key[119]_pad  ;
	input \key[11]_pad  ;
	input \key[120]_pad  ;
	input \key[121]_pad  ;
	input \key[122]_pad  ;
	input \key[123]_pad  ;
	input \key[124]_pad  ;
	input \key[125]_pad  ;
	input \key[126]_pad  ;
	input \key[127]_pad  ;
	input \key[12]_pad  ;
	input \key[13]_pad  ;
	input \key[14]_pad  ;
	input \key[15]_pad  ;
	input \key[16]_pad  ;
	input \key[17]_pad  ;
	input \key[18]_pad  ;
	input \key[19]_pad  ;
	input \key[1]_pad  ;
	input \key[20]_pad  ;
	input \key[21]_pad  ;
	input \key[22]_pad  ;
	input \key[23]_pad  ;
	input \key[24]_pad  ;
	input \key[25]_pad  ;
	input \key[26]_pad  ;
	input \key[27]_pad  ;
	input \key[28]_pad  ;
	input \key[29]_pad  ;
	input \key[2]_pad  ;
	input \key[30]_pad  ;
	input \key[31]_pad  ;
	input \key[32]_pad  ;
	input \key[33]_pad  ;
	input \key[34]_pad  ;
	input \key[35]_pad  ;
	input \key[36]_pad  ;
	input \key[37]_pad  ;
	input \key[38]_pad  ;
	input \key[39]_pad  ;
	input \key[3]_pad  ;
	input \key[40]_pad  ;
	input \key[41]_pad  ;
	input \key[42]_pad  ;
	input \key[43]_pad  ;
	input \key[44]_pad  ;
	input \key[45]_pad  ;
	input \key[46]_pad  ;
	input \key[47]_pad  ;
	input \key[48]_pad  ;
	input \key[49]_pad  ;
	input \key[4]_pad  ;
	input \key[50]_pad  ;
	input \key[51]_pad  ;
	input \key[52]_pad  ;
	input \key[53]_pad  ;
	input \key[54]_pad  ;
	input \key[55]_pad  ;
	input \key[56]_pad  ;
	input \key[57]_pad  ;
	input \key[58]_pad  ;
	input \key[59]_pad  ;
	input \key[5]_pad  ;
	input \key[60]_pad  ;
	input \key[61]_pad  ;
	input \key[62]_pad  ;
	input \key[63]_pad  ;
	input \key[64]_pad  ;
	input \key[65]_pad  ;
	input \key[66]_pad  ;
	input \key[67]_pad  ;
	input \key[68]_pad  ;
	input \key[69]_pad  ;
	input \key[6]_pad  ;
	input \key[70]_pad  ;
	input \key[71]_pad  ;
	input \key[72]_pad  ;
	input \key[73]_pad  ;
	input \key[74]_pad  ;
	input \key[75]_pad  ;
	input \key[76]_pad  ;
	input \key[77]_pad  ;
	input \key[78]_pad  ;
	input \key[79]_pad  ;
	input \key[7]_pad  ;
	input \key[80]_pad  ;
	input \key[81]_pad  ;
	input \key[82]_pad  ;
	input \key[83]_pad  ;
	input \key[84]_pad  ;
	input \key[85]_pad  ;
	input \key[86]_pad  ;
	input \key[87]_pad  ;
	input \key[88]_pad  ;
	input \key[89]_pad  ;
	input \key[8]_pad  ;
	input \key[90]_pad  ;
	input \key[91]_pad  ;
	input \key[92]_pad  ;
	input \key[93]_pad  ;
	input \key[94]_pad  ;
	input \key[95]_pad  ;
	input \key[96]_pad  ;
	input \key[97]_pad  ;
	input \key[98]_pad  ;
	input \key[99]_pad  ;
	input \key[9]_pad  ;
	input ld_pad ;
	input \ld_r_reg/P0001  ;
	input rst_pad ;
	input \sa00_reg[0]/P0001  ;
	input \sa00_reg[1]/P0001  ;
	input \sa00_reg[2]/P0001  ;
	input \sa00_reg[3]/P0001  ;
	input \sa00_reg[4]/P0001  ;
	input \sa00_reg[5]/P0001  ;
	input \sa00_reg[6]/NET0131  ;
	input \sa00_reg[7]/NET0131  ;
	input \sa01_reg[0]/P0001  ;
	input \sa01_reg[1]/P0001  ;
	input \sa01_reg[2]/P0001  ;
	input \sa01_reg[3]/P0001  ;
	input \sa01_reg[4]/P0001  ;
	input \sa01_reg[5]/P0001  ;
	input \sa01_reg[6]/NET0131  ;
	input \sa01_reg[7]/NET0131  ;
	input \sa02_reg[0]/P0001  ;
	input \sa02_reg[1]/P0001  ;
	input \sa02_reg[2]/P0001  ;
	input \sa02_reg[3]/P0001  ;
	input \sa02_reg[4]/P0001  ;
	input \sa02_reg[5]/P0001  ;
	input \sa02_reg[6]/NET0131  ;
	input \sa02_reg[7]/NET0131  ;
	input \sa03_reg[0]/P0001  ;
	input \sa03_reg[1]/P0001  ;
	input \sa03_reg[2]/P0001  ;
	input \sa03_reg[3]/P0001  ;
	input \sa03_reg[4]/P0001  ;
	input \sa03_reg[5]/P0001  ;
	input \sa03_reg[6]/NET0131  ;
	input \sa03_reg[7]/NET0131  ;
	input \sa10_reg[0]/P0001  ;
	input \sa10_reg[1]/P0001  ;
	input \sa10_reg[2]/P0001  ;
	input \sa10_reg[3]/P0001  ;
	input \sa10_reg[4]/P0001  ;
	input \sa10_reg[5]/P0001  ;
	input \sa10_reg[6]/NET0131  ;
	input \sa10_reg[7]/NET0131  ;
	input \sa11_reg[0]/P0001  ;
	input \sa11_reg[1]/P0001  ;
	input \sa11_reg[2]/P0001  ;
	input \sa11_reg[3]/P0001  ;
	input \sa11_reg[4]/P0001  ;
	input \sa11_reg[5]/P0001  ;
	input \sa11_reg[6]/NET0131  ;
	input \sa11_reg[7]/NET0131  ;
	input \sa12_reg[0]/P0001  ;
	input \sa12_reg[1]/P0001  ;
	input \sa12_reg[2]/P0001  ;
	input \sa12_reg[3]/P0001  ;
	input \sa12_reg[4]/P0001  ;
	input \sa12_reg[5]/P0001  ;
	input \sa12_reg[6]/NET0131  ;
	input \sa12_reg[7]/NET0131  ;
	input \sa13_reg[0]/P0001  ;
	input \sa13_reg[1]/P0001  ;
	input \sa13_reg[2]/P0001  ;
	input \sa13_reg[3]/P0001  ;
	input \sa13_reg[4]/P0001  ;
	input \sa13_reg[5]/P0001  ;
	input \sa13_reg[6]/NET0131  ;
	input \sa13_reg[7]/NET0131  ;
	input \sa20_reg[0]/P0001  ;
	input \sa20_reg[1]/P0001  ;
	input \sa20_reg[2]/P0001  ;
	input \sa20_reg[3]/P0001  ;
	input \sa20_reg[4]/P0001  ;
	input \sa20_reg[5]/P0001  ;
	input \sa20_reg[6]/NET0131  ;
	input \sa20_reg[7]/NET0131  ;
	input \sa21_reg[0]/P0001  ;
	input \sa21_reg[1]/P0001  ;
	input \sa21_reg[2]/P0001  ;
	input \sa21_reg[3]/P0001  ;
	input \sa21_reg[4]/P0001  ;
	input \sa21_reg[5]/P0001  ;
	input \sa21_reg[6]/NET0131  ;
	input \sa21_reg[7]/P0001  ;
	input \sa22_reg[0]/P0001  ;
	input \sa22_reg[1]/P0001  ;
	input \sa22_reg[2]/P0001  ;
	input \sa22_reg[3]/P0001  ;
	input \sa22_reg[4]/P0001  ;
	input \sa22_reg[5]/P0001  ;
	input \sa22_reg[6]/NET0131  ;
	input \sa22_reg[7]/NET0131  ;
	input \sa23_reg[0]/P0001  ;
	input \sa23_reg[1]/P0001  ;
	input \sa23_reg[2]/P0001  ;
	input \sa23_reg[3]/P0001  ;
	input \sa23_reg[4]/P0001  ;
	input \sa23_reg[5]/P0001  ;
	input \sa23_reg[6]/NET0131  ;
	input \sa23_reg[7]/NET0131  ;
	input \sa30_reg[0]/P0002  ;
	input \sa30_reg[1]/P0001  ;
	input \sa30_reg[2]/P0001  ;
	input \sa30_reg[3]/P0001  ;
	input \sa30_reg[4]/P0001  ;
	input \sa30_reg[5]/P0001  ;
	input \sa30_reg[6]/NET0131  ;
	input \sa30_reg[7]/P0001  ;
	input \sa31_reg[0]/P0002  ;
	input \sa31_reg[1]/P0001  ;
	input \sa31_reg[2]/P0001  ;
	input \sa31_reg[3]/P0001  ;
	input \sa31_reg[4]/P0001  ;
	input \sa31_reg[5]/P0001  ;
	input \sa31_reg[6]/NET0131  ;
	input \sa31_reg[7]/P0001  ;
	input \sa32_reg[0]/P0002  ;
	input \sa32_reg[1]/P0001  ;
	input \sa32_reg[2]/P0001  ;
	input \sa32_reg[3]/P0001  ;
	input \sa32_reg[4]/P0001  ;
	input \sa32_reg[5]/P0001  ;
	input \sa32_reg[6]/NET0131  ;
	input \sa32_reg[7]/P0001  ;
	input \sa33_reg[0]/P0001  ;
	input \sa33_reg[1]/P0001  ;
	input \sa33_reg[2]/P0001  ;
	input \sa33_reg[3]/P0001  ;
	input \sa33_reg[4]/P0001  ;
	input \sa33_reg[5]/P0001  ;
	input \sa33_reg[6]/P0001  ;
	input \sa33_reg[7]/NET0131  ;
	input \text_in_r_reg[0]/P0001  ;
	input \text_in_r_reg[100]/P0001  ;
	input \text_in_r_reg[101]/P0001  ;
	input \text_in_r_reg[102]/P0001  ;
	input \text_in_r_reg[103]/P0001  ;
	input \text_in_r_reg[104]/P0001  ;
	input \text_in_r_reg[105]/P0001  ;
	input \text_in_r_reg[106]/P0001  ;
	input \text_in_r_reg[107]/P0001  ;
	input \text_in_r_reg[108]/P0001  ;
	input \text_in_r_reg[109]/P0001  ;
	input \text_in_r_reg[10]/P0001  ;
	input \text_in_r_reg[110]/P0001  ;
	input \text_in_r_reg[111]/P0001  ;
	input \text_in_r_reg[112]/P0001  ;
	input \text_in_r_reg[113]/P0001  ;
	input \text_in_r_reg[114]/P0001  ;
	input \text_in_r_reg[115]/P0001  ;
	input \text_in_r_reg[116]/P0001  ;
	input \text_in_r_reg[117]/P0001  ;
	input \text_in_r_reg[118]/P0001  ;
	input \text_in_r_reg[119]/P0001  ;
	input \text_in_r_reg[11]/P0001  ;
	input \text_in_r_reg[120]/P0001  ;
	input \text_in_r_reg[121]/P0001  ;
	input \text_in_r_reg[122]/P0001  ;
	input \text_in_r_reg[123]/P0001  ;
	input \text_in_r_reg[124]/P0001  ;
	input \text_in_r_reg[125]/P0001  ;
	input \text_in_r_reg[126]/P0001  ;
	input \text_in_r_reg[127]/P0001  ;
	input \text_in_r_reg[12]/P0001  ;
	input \text_in_r_reg[13]/P0001  ;
	input \text_in_r_reg[14]/P0001  ;
	input \text_in_r_reg[15]/P0001  ;
	input \text_in_r_reg[16]/P0001  ;
	input \text_in_r_reg[17]/P0001  ;
	input \text_in_r_reg[18]/P0001  ;
	input \text_in_r_reg[19]/P0001  ;
	input \text_in_r_reg[1]/P0001  ;
	input \text_in_r_reg[20]/P0001  ;
	input \text_in_r_reg[21]/P0001  ;
	input \text_in_r_reg[22]/P0001  ;
	input \text_in_r_reg[23]/P0001  ;
	input \text_in_r_reg[24]/P0001  ;
	input \text_in_r_reg[25]/P0001  ;
	input \text_in_r_reg[26]/P0001  ;
	input \text_in_r_reg[27]/P0001  ;
	input \text_in_r_reg[28]/P0001  ;
	input \text_in_r_reg[29]/P0001  ;
	input \text_in_r_reg[2]/P0001  ;
	input \text_in_r_reg[30]/P0001  ;
	input \text_in_r_reg[31]/P0001  ;
	input \text_in_r_reg[32]/P0001  ;
	input \text_in_r_reg[33]/P0001  ;
	input \text_in_r_reg[34]/P0001  ;
	input \text_in_r_reg[35]/P0001  ;
	input \text_in_r_reg[36]/P0001  ;
	input \text_in_r_reg[37]/P0001  ;
	input \text_in_r_reg[38]/P0001  ;
	input \text_in_r_reg[39]/P0001  ;
	input \text_in_r_reg[3]/P0001  ;
	input \text_in_r_reg[40]/P0001  ;
	input \text_in_r_reg[41]/P0001  ;
	input \text_in_r_reg[42]/P0001  ;
	input \text_in_r_reg[43]/P0001  ;
	input \text_in_r_reg[44]/P0001  ;
	input \text_in_r_reg[45]/P0001  ;
	input \text_in_r_reg[46]/P0001  ;
	input \text_in_r_reg[47]/P0001  ;
	input \text_in_r_reg[48]/P0001  ;
	input \text_in_r_reg[49]/P0001  ;
	input \text_in_r_reg[4]/P0001  ;
	input \text_in_r_reg[50]/P0001  ;
	input \text_in_r_reg[51]/P0001  ;
	input \text_in_r_reg[52]/P0001  ;
	input \text_in_r_reg[53]/P0001  ;
	input \text_in_r_reg[54]/P0001  ;
	input \text_in_r_reg[55]/P0001  ;
	input \text_in_r_reg[56]/P0001  ;
	input \text_in_r_reg[57]/P0001  ;
	input \text_in_r_reg[58]/P0001  ;
	input \text_in_r_reg[59]/P0001  ;
	input \text_in_r_reg[5]/P0001  ;
	input \text_in_r_reg[60]/P0001  ;
	input \text_in_r_reg[61]/P0001  ;
	input \text_in_r_reg[62]/P0001  ;
	input \text_in_r_reg[63]/P0001  ;
	input \text_in_r_reg[64]/P0001  ;
	input \text_in_r_reg[65]/P0001  ;
	input \text_in_r_reg[66]/P0001  ;
	input \text_in_r_reg[67]/P0001  ;
	input \text_in_r_reg[68]/P0001  ;
	input \text_in_r_reg[69]/P0001  ;
	input \text_in_r_reg[6]/P0001  ;
	input \text_in_r_reg[70]/P0001  ;
	input \text_in_r_reg[71]/P0001  ;
	input \text_in_r_reg[72]/P0001  ;
	input \text_in_r_reg[73]/P0001  ;
	input \text_in_r_reg[74]/P0001  ;
	input \text_in_r_reg[75]/P0001  ;
	input \text_in_r_reg[76]/P0001  ;
	input \text_in_r_reg[77]/P0001  ;
	input \text_in_r_reg[78]/P0001  ;
	input \text_in_r_reg[79]/P0001  ;
	input \text_in_r_reg[7]/P0001  ;
	input \text_in_r_reg[80]/P0001  ;
	input \text_in_r_reg[81]/P0001  ;
	input \text_in_r_reg[82]/P0001  ;
	input \text_in_r_reg[83]/P0001  ;
	input \text_in_r_reg[84]/P0001  ;
	input \text_in_r_reg[85]/P0001  ;
	input \text_in_r_reg[86]/P0001  ;
	input \text_in_r_reg[87]/P0001  ;
	input \text_in_r_reg[88]/P0001  ;
	input \text_in_r_reg[89]/P0001  ;
	input \text_in_r_reg[8]/P0001  ;
	input \text_in_r_reg[90]/P0001  ;
	input \text_in_r_reg[91]/P0001  ;
	input \text_in_r_reg[92]/P0001  ;
	input \text_in_r_reg[93]/P0001  ;
	input \text_in_r_reg[94]/P0001  ;
	input \text_in_r_reg[95]/P0001  ;
	input \text_in_r_reg[96]/P0001  ;
	input \text_in_r_reg[97]/P0001  ;
	input \text_in_r_reg[98]/P0001  ;
	input \text_in_r_reg[99]/P0001  ;
	input \text_in_r_reg[9]/P0001  ;
	input \u0_r0_out_reg[24]/P0001  ;
	input \u0_r0_out_reg[25]/P0001  ;
	input \u0_r0_out_reg[26]/P0001  ;
	input \u0_r0_out_reg[27]/P0001  ;
	input \u0_r0_out_reg[28]/P0001  ;
	input \u0_r0_out_reg[29]/P0001  ;
	input \u0_r0_out_reg[30]/P0001  ;
	input \u0_r0_out_reg[31]/P0001  ;
	input \u0_r0_rcnt_reg[0]/P0001  ;
	input \u0_r0_rcnt_reg[1]/P0001  ;
	input \u0_r0_rcnt_reg[2]/P0001  ;
	input \u0_r0_rcnt_reg[3]/P0001  ;
	input \u0_w_reg[0][0]/P0001  ;
	input \u0_w_reg[0][10]/P0001  ;
	input \u0_w_reg[0][11]/P0001  ;
	input \u0_w_reg[0][12]/P0001  ;
	input \u0_w_reg[0][13]/P0001  ;
	input \u0_w_reg[0][14]/P0001  ;
	input \u0_w_reg[0][15]/P0001  ;
	input \u0_w_reg[0][16]/P0001  ;
	input \u0_w_reg[0][17]/P0001  ;
	input \u0_w_reg[0][18]/P0001  ;
	input \u0_w_reg[0][19]/P0001  ;
	input \u0_w_reg[0][1]/P0001  ;
	input \u0_w_reg[0][20]/P0001  ;
	input \u0_w_reg[0][21]/P0001  ;
	input \u0_w_reg[0][22]/P0001  ;
	input \u0_w_reg[0][23]/P0001  ;
	input \u0_w_reg[0][24]/P0001  ;
	input \u0_w_reg[0][25]/P0001  ;
	input \u0_w_reg[0][26]/P0001  ;
	input \u0_w_reg[0][27]/P0001  ;
	input \u0_w_reg[0][28]/P0001  ;
	input \u0_w_reg[0][29]/P0001  ;
	input \u0_w_reg[0][2]/P0001  ;
	input \u0_w_reg[0][30]/P0001  ;
	input \u0_w_reg[0][31]/P0001  ;
	input \u0_w_reg[0][3]/P0001  ;
	input \u0_w_reg[0][4]/P0001  ;
	input \u0_w_reg[0][5]/P0001  ;
	input \u0_w_reg[0][6]/P0001  ;
	input \u0_w_reg[0][7]/P0001  ;
	input \u0_w_reg[0][8]/P0001  ;
	input \u0_w_reg[0][9]/P0001  ;
	input \u0_w_reg[1][0]/P0001  ;
	input \u0_w_reg[1][10]/P0001  ;
	input \u0_w_reg[1][11]/P0001  ;
	input \u0_w_reg[1][12]/P0001  ;
	input \u0_w_reg[1][13]/P0001  ;
	input \u0_w_reg[1][14]/P0001  ;
	input \u0_w_reg[1][15]/P0001  ;
	input \u0_w_reg[1][16]/P0001  ;
	input \u0_w_reg[1][17]/P0001  ;
	input \u0_w_reg[1][18]/P0001  ;
	input \u0_w_reg[1][19]/P0001  ;
	input \u0_w_reg[1][1]/P0001  ;
	input \u0_w_reg[1][20]/P0001  ;
	input \u0_w_reg[1][21]/P0001  ;
	input \u0_w_reg[1][22]/P0001  ;
	input \u0_w_reg[1][23]/P0001  ;
	input \u0_w_reg[1][24]/P0002  ;
	input \u0_w_reg[1][25]/P0001  ;
	input \u0_w_reg[1][26]/P0001  ;
	input \u0_w_reg[1][27]/P0001  ;
	input \u0_w_reg[1][28]/P0001  ;
	input \u0_w_reg[1][29]/P0002  ;
	input \u0_w_reg[1][2]/P0001  ;
	input \u0_w_reg[1][30]/P0001  ;
	input \u0_w_reg[1][31]/P0001  ;
	input \u0_w_reg[1][3]/P0001  ;
	input \u0_w_reg[1][4]/P0001  ;
	input \u0_w_reg[1][5]/P0001  ;
	input \u0_w_reg[1][6]/P0001  ;
	input \u0_w_reg[1][7]/P0001  ;
	input \u0_w_reg[1][8]/P0001  ;
	input \u0_w_reg[1][9]/P0001  ;
	input \u0_w_reg[2][0]/P0001  ;
	input \u0_w_reg[2][10]/P0001  ;
	input \u0_w_reg[2][11]/P0001  ;
	input \u0_w_reg[2][12]/P0001  ;
	input \u0_w_reg[2][13]/P0001  ;
	input \u0_w_reg[2][14]/P0001  ;
	input \u0_w_reg[2][15]/P0001  ;
	input \u0_w_reg[2][16]/P0001  ;
	input \u0_w_reg[2][17]/P0001  ;
	input \u0_w_reg[2][18]/P0001  ;
	input \u0_w_reg[2][19]/P0001  ;
	input \u0_w_reg[2][1]/P0001  ;
	input \u0_w_reg[2][20]/P0001  ;
	input \u0_w_reg[2][21]/P0001  ;
	input \u0_w_reg[2][22]/P0001  ;
	input \u0_w_reg[2][23]/P0001  ;
	input \u0_w_reg[2][24]/P0001  ;
	input \u0_w_reg[2][25]/P0001  ;
	input \u0_w_reg[2][26]/P0001  ;
	input \u0_w_reg[2][27]/P0001  ;
	input \u0_w_reg[2][28]/P0001  ;
	input \u0_w_reg[2][29]/P0001  ;
	input \u0_w_reg[2][2]/P0001  ;
	input \u0_w_reg[2][30]/P0001  ;
	input \u0_w_reg[2][31]/P0001  ;
	input \u0_w_reg[2][3]/P0001  ;
	input \u0_w_reg[2][4]/P0001  ;
	input \u0_w_reg[2][5]/P0001  ;
	input \u0_w_reg[2][6]/P0001  ;
	input \u0_w_reg[2][7]/P0001  ;
	input \u0_w_reg[2][8]/P0001  ;
	input \u0_w_reg[2][9]/P0001  ;
	input \u0_w_reg[3][0]/P0001  ;
	input \u0_w_reg[3][10]/P0001  ;
	input \u0_w_reg[3][11]/P0001  ;
	input \u0_w_reg[3][12]/P0001  ;
	input \u0_w_reg[3][13]/P0001  ;
	input \u0_w_reg[3][14]/P0001  ;
	input \u0_w_reg[3][15]/P0001  ;
	input \u0_w_reg[3][16]/P0001  ;
	input \u0_w_reg[3][17]/P0001  ;
	input \u0_w_reg[3][18]/P0001  ;
	input \u0_w_reg[3][19]/P0001  ;
	input \u0_w_reg[3][1]/P0001  ;
	input \u0_w_reg[3][20]/P0001  ;
	input \u0_w_reg[3][21]/P0001  ;
	input \u0_w_reg[3][22]/P0001  ;
	input \u0_w_reg[3][23]/P0001  ;
	input \u0_w_reg[3][24]/P0001  ;
	input \u0_w_reg[3][25]/P0001  ;
	input \u0_w_reg[3][26]/P0001  ;
	input \u0_w_reg[3][27]/P0001  ;
	input \u0_w_reg[3][28]/P0001  ;
	input \u0_w_reg[3][29]/P0001  ;
	input \u0_w_reg[3][2]/P0001  ;
	input \u0_w_reg[3][30]/P0001  ;
	input \u0_w_reg[3][31]/P0001  ;
	input \u0_w_reg[3][3]/P0001  ;
	input \u0_w_reg[3][4]/P0001  ;
	input \u0_w_reg[3][5]/P0001  ;
	input \u0_w_reg[3][6]/P0001  ;
	input \u0_w_reg[3][7]/P0001  ;
	input \u0_w_reg[3][8]/P0001  ;
	input \u0_w_reg[3][9]/P0001  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g21/_0_  ;
	output \g56610/_0_  ;
	output \g56611/_0_  ;
	output \g56612/_0_  ;
	output \g56613/_0_  ;
	output \g56614/_0_  ;
	output \g56615/_0_  ;
	output \g56616/_0_  ;
	output \g56617/_0_  ;
	output \g56630/_0_  ;
	output \g56631/_0_  ;
	output \g56632/_0_  ;
	output \g56633/_0_  ;
	output \g56634/_0_  ;
	output \g56635/_0_  ;
	output \g56645/_0_  ;
	output \g56646/_0_  ;
	output \g56647/_0_  ;
	output \g56648/_0_  ;
	output \g56649/_0_  ;
	output \g56650/_0_  ;
	output \g56651/_0_  ;
	output \g56652/_0_  ;
	output \g56666/_0_  ;
	output \g56667/_0_  ;
	output \g56668/_0_  ;
	output \g56669/_0_  ;
	output \g56670/_0_  ;
	output \g56671/_0_  ;
	output \g56672/_0_  ;
	output \g56674/_0_  ;
	output \g56675/_0_  ;
	output \g56704/_0_  ;
	output \g56739/_0_  ;
	output \g56743/_0_  ;
	output \g56763/_0_  ;
	output \g56776/_0_  ;
	output \g56812/_0_  ;
	output \g56818/_0_  ;
	output \g56861/_0_  ;
	output \g56874/_0_  ;
	output \g56919/_0_  ;
	output \g56920/_0_  ;
	output \g56921/_0_  ;
	output \g56923/_0_  ;
	output \g56924/_0_  ;
	output \g56925/_0_  ;
	output \g56926/_0_  ;
	output \g56956/_0_  ;
	output \g56957/_0_  ;
	output \g56958/_0_  ;
	output \g56959/_0_  ;
	output \g56960/_0_  ;
	output \g56961/_0_  ;
	output \g56972/_0_  ;
	output \g56973/_0_  ;
	output \g56974/_0_  ;
	output \g56976/_0_  ;
	output \g56977/_0_  ;
	output \g56978/_0_  ;
	output \g56979/_0_  ;
	output \g56980/_0_  ;
	output \g57008/_0_  ;
	output \g57010/_0_  ;
	output \g57011/_0_  ;
	output \g57012/_0_  ;
	output \g57013/_0_  ;
	output \g57014/_0_  ;
	output \g57015/_0_  ;
	output \g57016/_0_  ;
	output \g57017/_0_  ;
	output \g57086/_0_  ;
	output \g57091/_0_  ;
	output \g57114/_0_  ;
	output \g57129/_0_  ;
	output \g57163/_0_  ;
	output \g57171/_0_  ;
	output \g57204/_0_  ;
	output \g57218/_0_  ;
	output \g57262/_0_  ;
	output \g57263/_0_  ;
	output \g57264/_0_  ;
	output \g57265/_0_  ;
	output \g57266/_0_  ;
	output \g57267/_0_  ;
	output \g57268/_0_  ;
	output \g57269/_0_  ;
	output \g57300/_0_  ;
	output \g57301/_0_  ;
	output \g57302/_0_  ;
	output \g57303/_0_  ;
	output \g57304/_0_  ;
	output \g57316/_0_  ;
	output \g57317/_0_  ;
	output \g57319/_0_  ;
	output \g57320/_0_  ;
	output \g57321/_0_  ;
	output \g57322/_0_  ;
	output \g57323/_0_  ;
	output \g57324/_0_  ;
	output \g57350/_0_  ;
	output \g57353/_0_  ;
	output \g57354/_0_  ;
	output \g57355/_0_  ;
	output \g57356/_0_  ;
	output \g57357/_0_  ;
	output \g57358/_0_  ;
	output \g57359/_0_  ;
	output \g57360/_0_  ;
	output \g57427/_0_  ;
	output \g57432/_0_  ;
	output \g57456/_0_  ;
	output \g57471/_0_  ;
	output \g57506/_0_  ;
	output \g57512/_0_  ;
	output \g57540/_0_  ;
	output \g57547/_0_  ;
	output \g57654/_0_  ;
	output \g57655/_0_  ;
	output \g57656/_0_  ;
	output \g57657/_0_  ;
	output \g57658/_0_  ;
	output \g57676/_0_  ;
	output \g57677/_0_  ;
	output \g57678/_0_  ;
	output \g57679/_0_  ;
	output \g57680/_0_  ;
	output \g57681/_0_  ;
	output \g57682/_0_  ;
	output \g57683/_0_  ;
	output \g57684/_0_  ;
	output \g57685/_0_  ;
	output \g57686/_0_  ;
	output \g57687/_0_  ;
	output \g57688/_0_  ;
	output \g57689/_0_  ;
	output \g57690/_0_  ;
	output \g57691/_0_  ;
	output \g57700/_0_  ;
	output \g57701/_0_  ;
	output \g57702/_0_  ;
	output \g57703/_0_  ;
	output \g57704/_0_  ;
	output \g57705/_0_  ;
	output \g57706/_0_  ;
	output \g57707/_0_  ;
	output \g57708/_0_  ;
	output \g57709/_3_  ;
	output \g57710/_3_  ;
	output \g57711/_0_  ;
	output \g57712/_3_  ;
	output \g57715/_3_  ;
	output \g57716/_3_  ;
	output \g57767/_0_  ;
	output \g57768/_3_  ;
	output \g57769/_3_  ;
	output \g57770/_3_  ;
	output \g57771/_3_  ;
	output \g57777/_3_  ;
	output \g57779/_3_  ;
	output \g57804/_3_  ;
	output \g57805/_3_  ;
	output \g57806/_3_  ;
	output \g57807/_3_  ;
	output \g57808/_3_  ;
	output \g57809/_3_  ;
	output \g57810/_3_  ;
	output \g57811/_3_  ;
	output \g57812/_3_  ;
	output \g57813/_3_  ;
	output \g57814/_3_  ;
	output \g57815/_3_  ;
	output \g57816/_0_  ;
	output \g57817/_3_  ;
	output \g57818/_3_  ;
	output \g57819/_3_  ;
	output \g57822/_3_  ;
	output \g57823/_3_  ;
	output \g57824/_3_  ;
	output \g57830/_3_  ;
	output \g57835/_3_  ;
	output \g57836/_3_  ;
	output \g57837/_3_  ;
	output \g57841/_3_  ;
	output \g57842/_3_  ;
	output \g57843/_3_  ;
	output \g57854/_3_  ;
	output \g57855/_3_  ;
	output \g57856/_3_  ;
	output \g57857/_3_  ;
	output \g57858/_3_  ;
	output \g57859/_3_  ;
	output \g57860/_3_  ;
	output \g57861/_3_  ;
	output \g57871/_3_  ;
	output \g57872/_3_  ;
	output \g57874/_3_  ;
	output \g57968/_3_  ;
	output \g57969/_3_  ;
	output \g57970/_3_  ;
	output \g57971/_3_  ;
	output \g57980/_3_  ;
	output \g57983/_3_  ;
	output \g57984/_3_  ;
	output \g57985/_3_  ;
	output \g58012/_3_  ;
	output \g58013/_3_  ;
	output \g58015/_3_  ;
	output \g58057/_3_  ;
	output \g58058/_3_  ;
	output \g58059/_3_  ;
	output \g58189/_3_  ;
	output \g58190/_3_  ;
	output \g58191/_3_  ;
	output \g58192/_3_  ;
	output \g58193/_3_  ;
	output \g58194/_3_  ;
	output \g58195/_3_  ;
	output \g58196/_3_  ;
	output \g58197/_3_  ;
	output \g58224/_3_  ;
	output \g58226/_3_  ;
	output \g58229/_3_  ;
	output \g58255/_3_  ;
	output \g58256/_3_  ;
	output \g58257/_3_  ;
	output \g58258/_3_  ;
	output \g58259/_3_  ;
	output \g58260/_3_  ;
	output \g58261/_3_  ;
	output \g58262/_3_  ;
	output \g58263/_3_  ;
	output \g58264/_3_  ;
	output \g58265/_3_  ;
	output \g58266/_3_  ;
	output \g58267/_3_  ;
	output \g58268/_3_  ;
	output \g58269/_3_  ;
	output \g58270/_0_  ;
	output \g58271/_3_  ;
	output \g58272/_3_  ;
	output \g58273/_3_  ;
	output \g58274/_3_  ;
	output \g58275/_3_  ;
	output \g58276/_3_  ;
	output \g58277/_3_  ;
	output \g58278/_3_  ;
	output \g58279/_3_  ;
	output \g58285/_3_  ;
	output \g58286/_3_  ;
	output \g58288/_3_  ;
	output \g58289/_3_  ;
	output \g58290/_3_  ;
	output \g58292/_3_  ;
	output \g58294/_3_  ;
	output \g58295/_3_  ;
	output \g58297/_3_  ;
	output \g58330/_0_  ;
	output \g58331/_0_  ;
	output \g58332/_0_  ;
	output \g58333/_0_  ;
	output \g58444/_3_  ;
	output \g58445/_3_  ;
	output \g58446/_3_  ;
	output \g58462/_0_  ;
	output \g58506/_0_  ;
	output \g58507/_0_  ;
	output \g58508/_0_  ;
	output \g58509/_0_  ;
	output \g58531/_0_  ;
	output \g58532/_0_  ;
	output \g58533/_0_  ;
	output \g58550/_0_  ;
	output \g58551/_0_  ;
	output \g58552/_0_  ;
	output \g58553/_0_  ;
	output \g58554/_0_  ;
	output \g58555/_0_  ;
	output \g58556/_0_  ;
	output \g58557/_0_  ;
	output \g58558/_0_  ;
	output \g58559/_0_  ;
	output \g58560/_0_  ;
	output \g58600/_3_  ;
	output \g58601/_3_  ;
	output \g58602/_3_  ;
	output \g58603/_3_  ;
	output \g58604/_3_  ;
	output \g58605/_3_  ;
	output \g58606/_3_  ;
	output \g58607/_3_  ;
	output \g58608/_3_  ;
	output \g58611/_0_  ;
	output \g58612/_0_  ;
	output \g58613/_0_  ;
	output \g58614/_0_  ;
	output \g58617/_0_  ;
	output \g58618/_0_  ;
	output \g58619/_0_  ;
	output \g58634/_0_  ;
	output \g58635/_0_  ;
	output \g58636/_0_  ;
	output \g58637/_0_  ;
	output \g58638/_0_  ;
	output \g58639/_0_  ;
	output \g58640/_0_  ;
	output \g58641/_0_  ;
	output \g58829/_3_  ;
	output \g58830/_3_  ;
	output \g58831/_3_  ;
	output \g58832/_3_  ;
	output \g58833/_3_  ;
	output \g58834/_3_  ;
	output \g58835/_0_  ;
	output \g58844/_0_  ;
	output \g58902/_0_  ;
	output \g58903/_0_  ;
	output \g58904/_0_  ;
	output \g58905/_0_  ;
	output \g58910/_0_  ;
	output \g58913/_0_  ;
	output \g58934/_0_  ;
	output \g58935/_0_  ;
	output \g58936/_0_  ;
	output \g58937/_0_  ;
	output \g58938/_0_  ;
	output \g58970/_0_  ;
	output \g58972/_0_  ;
	output \g58994/_0_  ;
	output \g58995/_0_  ;
	output \g58996/_0_  ;
	output \g58997/_0_  ;
	output \g58998/_0_  ;
	output \g58999/_0_  ;
	output \g59000/_0_  ;
	output \g59002/_0_  ;
	output \g59003/_0_  ;
	output \g59004/_0_  ;
	output \g59254/_0_  ;
	output \g59257/_0_  ;
	output \g59258/_0_  ;
	output \g59259/_0_  ;
	output \g59276/_0_  ;
	output \g59277/_0_  ;
	output \g59278/_0_  ;
	output \g59279/_0_  ;
	output \g59280/_0_  ;
	output \g59291/_0_  ;
	output \g59292/_0_  ;
	output \g59293/_0_  ;
	output \g59294/_0_  ;
	output \g59295/_0_  ;
	output \g59308/_0_  ;
	output \g59309/_0_  ;
	output \g59310/_0_  ;
	output \g59311/_0_  ;
	output \g59330/_0_  ;
	output \g59331/_0_  ;
	output \g59332/_0_  ;
	output \g59333/_0_  ;
	output \g59334/_0_  ;
	output \g59335/_0_  ;
	output \g59336/_0_  ;
	output \g59337/_0_  ;
	output \g59338/_0_  ;
	output \g59339/_0_  ;
	output \g59596/_0_  ;
	output \g59597/_0_  ;
	output \g59598/_0_  ;
	output \g59599/_0_  ;
	output \g59625/_0_  ;
	output \g59626/_0_  ;
	output \g59627/_0_  ;
	output \g59628/_0_  ;
	output \g59837/_0_  ;
	output \g59838/_0_  ;
	output \g59839/_0_  ;
	output \g59840/_0_  ;
	output \g60090/_0_  ;
	output \g60320/_0_  ;
	output \g60321/_0_  ;
	output \g60409/_0_  ;
	output \g60539/_0_  ;
	output \g60860/_0_  ;
	output \g60977/_0_  ;
	output \g61012/_0_  ;
	output \g61185/_0_  ;
	output \g61524/_2_  ;
	output \g61776/_0_  ;
	output \g61895/_0_  ;
	output \g61897/_0_  ;
	output \g62220/_0_  ;
	output \g65958/_0_  ;
	output \g72347/_3_  ;
	output \g77848/_0_  ;
	output \g85056/_0_  ;
	output \sa30_reg[0]/_05_  ;
	output \sa31_reg[0]/_05_  ;
	output \sa32_reg[0]/_05_  ;
	output \u0_w_reg[1][24]/_05_  ;
	output \u0_w_reg[1][29]/_05_  ;
	wire _w10982_ ;
	wire _w10981_ ;
	wire _w10980_ ;
	wire _w10979_ ;
	wire _w10978_ ;
	wire _w10977_ ;
	wire _w10976_ ;
	wire _w10975_ ;
	wire _w10974_ ;
	wire _w10973_ ;
	wire _w10972_ ;
	wire _w10971_ ;
	wire _w10970_ ;
	wire _w10969_ ;
	wire _w10968_ ;
	wire _w10967_ ;
	wire _w10966_ ;
	wire _w10965_ ;
	wire _w10964_ ;
	wire _w10963_ ;
	wire _w10962_ ;
	wire _w10961_ ;
	wire _w10960_ ;
	wire _w10959_ ;
	wire _w10958_ ;
	wire _w10957_ ;
	wire _w10956_ ;
	wire _w10955_ ;
	wire _w10954_ ;
	wire _w10953_ ;
	wire _w10952_ ;
	wire _w10951_ ;
	wire _w10950_ ;
	wire _w10949_ ;
	wire _w10948_ ;
	wire _w10947_ ;
	wire _w10946_ ;
	wire _w10945_ ;
	wire _w10944_ ;
	wire _w10943_ ;
	wire _w10942_ ;
	wire _w10941_ ;
	wire _w10940_ ;
	wire _w10939_ ;
	wire _w10938_ ;
	wire _w10937_ ;
	wire _w10936_ ;
	wire _w10935_ ;
	wire _w10934_ ;
	wire _w10933_ ;
	wire _w10932_ ;
	wire _w10931_ ;
	wire _w10930_ ;
	wire _w10929_ ;
	wire _w10928_ ;
	wire _w10927_ ;
	wire _w10926_ ;
	wire _w10925_ ;
	wire _w10924_ ;
	wire _w10923_ ;
	wire _w10922_ ;
	wire _w10921_ ;
	wire _w10920_ ;
	wire _w10919_ ;
	wire _w10918_ ;
	wire _w10917_ ;
	wire _w10916_ ;
	wire _w10915_ ;
	wire _w10914_ ;
	wire _w10913_ ;
	wire _w10912_ ;
	wire _w10911_ ;
	wire _w10910_ ;
	wire _w10909_ ;
	wire _w10908_ ;
	wire _w10907_ ;
	wire _w10906_ ;
	wire _w10905_ ;
	wire _w10904_ ;
	wire _w10903_ ;
	wire _w10902_ ;
	wire _w10901_ ;
	wire _w10900_ ;
	wire _w10899_ ;
	wire _w10898_ ;
	wire _w10897_ ;
	wire _w10896_ ;
	wire _w10895_ ;
	wire _w10894_ ;
	wire _w10893_ ;
	wire _w10892_ ;
	wire _w10891_ ;
	wire _w10890_ ;
	wire _w10889_ ;
	wire _w10888_ ;
	wire _w10887_ ;
	wire _w10886_ ;
	wire _w10885_ ;
	wire _w10884_ ;
	wire _w10883_ ;
	wire _w10882_ ;
	wire _w10881_ ;
	wire _w10880_ ;
	wire _w10879_ ;
	wire _w10878_ ;
	wire _w10877_ ;
	wire _w10876_ ;
	wire _w10875_ ;
	wire _w10874_ ;
	wire _w10873_ ;
	wire _w10872_ ;
	wire _w10871_ ;
	wire _w10870_ ;
	wire _w10869_ ;
	wire _w10868_ ;
	wire _w10867_ ;
	wire _w10866_ ;
	wire _w10865_ ;
	wire _w10864_ ;
	wire _w10863_ ;
	wire _w10862_ ;
	wire _w10861_ ;
	wire _w10860_ ;
	wire _w10859_ ;
	wire _w10858_ ;
	wire _w10857_ ;
	wire _w10856_ ;
	wire _w10855_ ;
	wire _w10854_ ;
	wire _w10853_ ;
	wire _w10852_ ;
	wire _w10851_ ;
	wire _w10850_ ;
	wire _w10849_ ;
	wire _w10848_ ;
	wire _w10847_ ;
	wire _w10846_ ;
	wire _w10845_ ;
	wire _w10844_ ;
	wire _w10843_ ;
	wire _w10842_ ;
	wire _w10841_ ;
	wire _w10840_ ;
	wire _w10839_ ;
	wire _w10838_ ;
	wire _w10837_ ;
	wire _w10836_ ;
	wire _w10835_ ;
	wire _w10834_ ;
	wire _w10833_ ;
	wire _w10832_ ;
	wire _w10831_ ;
	wire _w10830_ ;
	wire _w10829_ ;
	wire _w10828_ ;
	wire _w10827_ ;
	wire _w10826_ ;
	wire _w10825_ ;
	wire _w10824_ ;
	wire _w10823_ ;
	wire _w10822_ ;
	wire _w10821_ ;
	wire _w10820_ ;
	wire _w10819_ ;
	wire _w10818_ ;
	wire _w10817_ ;
	wire _w10816_ ;
	wire _w10815_ ;
	wire _w10814_ ;
	wire _w10813_ ;
	wire _w10812_ ;
	wire _w10811_ ;
	wire _w10810_ ;
	wire _w10809_ ;
	wire _w10808_ ;
	wire _w10807_ ;
	wire _w10806_ ;
	wire _w5619_ ;
	wire _w5618_ ;
	wire _w5617_ ;
	wire _w5616_ ;
	wire _w5615_ ;
	wire _w5614_ ;
	wire _w5613_ ;
	wire _w5612_ ;
	wire _w5611_ ;
	wire _w5610_ ;
	wire _w5609_ ;
	wire _w5608_ ;
	wire _w5607_ ;
	wire _w5606_ ;
	wire _w5605_ ;
	wire _w5604_ ;
	wire _w5603_ ;
	wire _w5602_ ;
	wire _w5601_ ;
	wire _w5600_ ;
	wire _w5599_ ;
	wire _w5598_ ;
	wire _w5597_ ;
	wire _w5596_ ;
	wire _w5595_ ;
	wire _w5594_ ;
	wire _w5593_ ;
	wire _w5592_ ;
	wire _w5591_ ;
	wire _w5590_ ;
	wire _w5589_ ;
	wire _w5588_ ;
	wire _w5587_ ;
	wire _w5586_ ;
	wire _w5585_ ;
	wire _w5584_ ;
	wire _w5583_ ;
	wire _w5582_ ;
	wire _w5581_ ;
	wire _w5580_ ;
	wire _w5579_ ;
	wire _w5578_ ;
	wire _w5577_ ;
	wire _w5576_ ;
	wire _w5575_ ;
	wire _w5574_ ;
	wire _w5573_ ;
	wire _w5572_ ;
	wire _w5571_ ;
	wire _w5570_ ;
	wire _w5569_ ;
	wire _w5568_ ;
	wire _w5567_ ;
	wire _w5566_ ;
	wire _w5565_ ;
	wire _w5564_ ;
	wire _w5563_ ;
	wire _w5562_ ;
	wire _w5561_ ;
	wire _w5560_ ;
	wire _w5559_ ;
	wire _w5558_ ;
	wire _w5557_ ;
	wire _w5556_ ;
	wire _w5555_ ;
	wire _w5554_ ;
	wire _w5553_ ;
	wire _w5552_ ;
	wire _w5551_ ;
	wire _w5550_ ;
	wire _w5549_ ;
	wire _w5548_ ;
	wire _w5547_ ;
	wire _w5546_ ;
	wire _w5545_ ;
	wire _w5544_ ;
	wire _w5543_ ;
	wire _w5542_ ;
	wire _w5541_ ;
	wire _w5540_ ;
	wire _w5539_ ;
	wire _w5538_ ;
	wire _w5537_ ;
	wire _w5536_ ;
	wire _w5535_ ;
	wire _w5534_ ;
	wire _w5533_ ;
	wire _w5532_ ;
	wire _w5531_ ;
	wire _w5530_ ;
	wire _w5529_ ;
	wire _w5528_ ;
	wire _w5527_ ;
	wire _w5526_ ;
	wire _w5525_ ;
	wire _w5524_ ;
	wire _w5523_ ;
	wire _w5522_ ;
	wire _w5521_ ;
	wire _w5520_ ;
	wire _w5519_ ;
	wire _w5518_ ;
	wire _w5517_ ;
	wire _w5516_ ;
	wire _w5515_ ;
	wire _w5514_ ;
	wire _w5513_ ;
	wire _w5512_ ;
	wire _w5511_ ;
	wire _w5510_ ;
	wire _w5509_ ;
	wire _w5508_ ;
	wire _w5507_ ;
	wire _w5506_ ;
	wire _w5505_ ;
	wire _w5504_ ;
	wire _w5503_ ;
	wire _w5502_ ;
	wire _w5501_ ;
	wire _w5500_ ;
	wire _w5499_ ;
	wire _w5498_ ;
	wire _w5497_ ;
	wire _w5496_ ;
	wire _w5495_ ;
	wire _w5494_ ;
	wire _w5493_ ;
	wire _w5492_ ;
	wire _w5491_ ;
	wire _w5490_ ;
	wire _w5489_ ;
	wire _w5488_ ;
	wire _w5487_ ;
	wire _w5486_ ;
	wire _w5485_ ;
	wire _w5484_ ;
	wire _w5483_ ;
	wire _w5482_ ;
	wire _w5481_ ;
	wire _w5480_ ;
	wire _w5479_ ;
	wire _w5478_ ;
	wire _w5477_ ;
	wire _w5476_ ;
	wire _w5475_ ;
	wire _w5474_ ;
	wire _w5473_ ;
	wire _w5472_ ;
	wire _w5471_ ;
	wire _w5470_ ;
	wire _w5469_ ;
	wire _w5468_ ;
	wire _w5467_ ;
	wire _w5466_ ;
	wire _w5465_ ;
	wire _w5464_ ;
	wire _w5463_ ;
	wire _w5462_ ;
	wire _w5461_ ;
	wire _w5460_ ;
	wire _w5459_ ;
	wire _w5458_ ;
	wire _w5457_ ;
	wire _w5456_ ;
	wire _w5455_ ;
	wire _w5454_ ;
	wire _w5453_ ;
	wire _w5452_ ;
	wire _w5451_ ;
	wire _w5450_ ;
	wire _w5449_ ;
	wire _w5448_ ;
	wire _w5447_ ;
	wire _w5446_ ;
	wire _w5445_ ;
	wire _w5444_ ;
	wire _w5443_ ;
	wire _w5442_ ;
	wire _w5441_ ;
	wire _w5440_ ;
	wire _w5439_ ;
	wire _w5438_ ;
	wire _w5437_ ;
	wire _w5436_ ;
	wire _w5435_ ;
	wire _w5434_ ;
	wire _w5433_ ;
	wire _w5432_ ;
	wire _w5431_ ;
	wire _w5430_ ;
	wire _w5429_ ;
	wire _w5428_ ;
	wire _w5427_ ;
	wire _w5426_ ;
	wire _w5425_ ;
	wire _w5424_ ;
	wire _w5423_ ;
	wire _w5422_ ;
	wire _w5421_ ;
	wire _w5420_ ;
	wire _w5419_ ;
	wire _w5418_ ;
	wire _w5417_ ;
	wire _w5416_ ;
	wire _w5415_ ;
	wire _w5414_ ;
	wire _w5413_ ;
	wire _w5412_ ;
	wire _w5411_ ;
	wire _w5410_ ;
	wire _w5409_ ;
	wire _w5408_ ;
	wire _w5407_ ;
	wire _w5406_ ;
	wire _w5405_ ;
	wire _w5404_ ;
	wire _w5403_ ;
	wire _w5402_ ;
	wire _w5401_ ;
	wire _w5400_ ;
	wire _w5399_ ;
	wire _w5398_ ;
	wire _w5397_ ;
	wire _w5396_ ;
	wire _w5395_ ;
	wire _w5394_ ;
	wire _w5393_ ;
	wire _w5392_ ;
	wire _w5391_ ;
	wire _w5390_ ;
	wire _w5389_ ;
	wire _w5388_ ;
	wire _w5387_ ;
	wire _w5386_ ;
	wire _w5385_ ;
	wire _w5384_ ;
	wire _w5383_ ;
	wire _w5382_ ;
	wire _w5381_ ;
	wire _w5380_ ;
	wire _w5379_ ;
	wire _w5378_ ;
	wire _w5377_ ;
	wire _w5376_ ;
	wire _w5375_ ;
	wire _w5374_ ;
	wire _w5373_ ;
	wire _w5372_ ;
	wire _w5371_ ;
	wire _w5370_ ;
	wire _w5369_ ;
	wire _w5368_ ;
	wire _w5367_ ;
	wire _w5366_ ;
	wire _w5365_ ;
	wire _w5364_ ;
	wire _w5363_ ;
	wire _w5362_ ;
	wire _w5361_ ;
	wire _w5360_ ;
	wire _w5359_ ;
	wire _w5358_ ;
	wire _w5357_ ;
	wire _w5356_ ;
	wire _w5355_ ;
	wire _w5354_ ;
	wire _w5353_ ;
	wire _w5352_ ;
	wire _w5351_ ;
	wire _w5350_ ;
	wire _w5349_ ;
	wire _w5348_ ;
	wire _w5347_ ;
	wire _w5346_ ;
	wire _w5345_ ;
	wire _w5344_ ;
	wire _w5343_ ;
	wire _w5342_ ;
	wire _w5341_ ;
	wire _w5340_ ;
	wire _w5339_ ;
	wire _w5338_ ;
	wire _w5337_ ;
	wire _w5336_ ;
	wire _w5335_ ;
	wire _w5334_ ;
	wire _w5333_ ;
	wire _w5332_ ;
	wire _w5331_ ;
	wire _w5330_ ;
	wire _w5329_ ;
	wire _w5328_ ;
	wire _w5327_ ;
	wire _w5326_ ;
	wire _w5325_ ;
	wire _w5324_ ;
	wire _w5323_ ;
	wire _w5322_ ;
	wire _w5321_ ;
	wire _w5320_ ;
	wire _w5319_ ;
	wire _w5318_ ;
	wire _w5317_ ;
	wire _w5316_ ;
	wire _w5315_ ;
	wire _w5314_ ;
	wire _w5313_ ;
	wire _w5312_ ;
	wire _w5311_ ;
	wire _w5310_ ;
	wire _w5309_ ;
	wire _w5308_ ;
	wire _w5307_ ;
	wire _w5306_ ;
	wire _w5305_ ;
	wire _w5304_ ;
	wire _w5303_ ;
	wire _w5302_ ;
	wire _w5301_ ;
	wire _w5300_ ;
	wire _w5299_ ;
	wire _w5298_ ;
	wire _w5297_ ;
	wire _w5296_ ;
	wire _w5295_ ;
	wire _w5294_ ;
	wire _w5293_ ;
	wire _w5292_ ;
	wire _w5291_ ;
	wire _w5290_ ;
	wire _w5289_ ;
	wire _w5288_ ;
	wire _w5287_ ;
	wire _w5286_ ;
	wire _w5285_ ;
	wire _w5284_ ;
	wire _w5283_ ;
	wire _w5282_ ;
	wire _w5281_ ;
	wire _w5280_ ;
	wire _w5279_ ;
	wire _w5278_ ;
	wire _w5277_ ;
	wire _w5276_ ;
	wire _w5275_ ;
	wire _w5274_ ;
	wire _w5273_ ;
	wire _w5272_ ;
	wire _w5271_ ;
	wire _w5270_ ;
	wire _w5269_ ;
	wire _w5268_ ;
	wire _w5267_ ;
	wire _w5266_ ;
	wire _w5265_ ;
	wire _w5264_ ;
	wire _w5263_ ;
	wire _w5262_ ;
	wire _w5261_ ;
	wire _w5260_ ;
	wire _w5259_ ;
	wire _w5258_ ;
	wire _w5257_ ;
	wire _w5256_ ;
	wire _w5255_ ;
	wire _w5254_ ;
	wire _w5253_ ;
	wire _w5252_ ;
	wire _w5251_ ;
	wire _w5250_ ;
	wire _w5249_ ;
	wire _w5248_ ;
	wire _w5247_ ;
	wire _w5246_ ;
	wire _w5245_ ;
	wire _w5244_ ;
	wire _w5243_ ;
	wire _w5242_ ;
	wire _w5241_ ;
	wire _w5240_ ;
	wire _w5239_ ;
	wire _w5238_ ;
	wire _w5237_ ;
	wire _w5236_ ;
	wire _w5235_ ;
	wire _w5234_ ;
	wire _w5233_ ;
	wire _w5232_ ;
	wire _w5231_ ;
	wire _w5230_ ;
	wire _w5229_ ;
	wire _w5228_ ;
	wire _w5227_ ;
	wire _w5226_ ;
	wire _w5225_ ;
	wire _w5224_ ;
	wire _w5223_ ;
	wire _w5222_ ;
	wire _w5221_ ;
	wire _w5220_ ;
	wire _w5219_ ;
	wire _w5218_ ;
	wire _w5217_ ;
	wire _w5216_ ;
	wire _w5215_ ;
	wire _w5214_ ;
	wire _w5213_ ;
	wire _w5212_ ;
	wire _w5211_ ;
	wire _w5210_ ;
	wire _w5209_ ;
	wire _w5208_ ;
	wire _w5207_ ;
	wire _w5206_ ;
	wire _w5205_ ;
	wire _w5204_ ;
	wire _w5203_ ;
	wire _w5202_ ;
	wire _w5201_ ;
	wire _w5200_ ;
	wire _w5199_ ;
	wire _w5198_ ;
	wire _w5197_ ;
	wire _w5196_ ;
	wire _w5195_ ;
	wire _w5194_ ;
	wire _w5193_ ;
	wire _w5192_ ;
	wire _w5191_ ;
	wire _w5190_ ;
	wire _w5189_ ;
	wire _w5188_ ;
	wire _w5187_ ;
	wire _w5186_ ;
	wire _w5185_ ;
	wire _w5184_ ;
	wire _w5183_ ;
	wire _w5182_ ;
	wire _w5181_ ;
	wire _w5180_ ;
	wire _w5179_ ;
	wire _w5178_ ;
	wire _w5177_ ;
	wire _w5176_ ;
	wire _w5175_ ;
	wire _w5174_ ;
	wire _w5173_ ;
	wire _w5172_ ;
	wire _w5171_ ;
	wire _w5170_ ;
	wire _w5169_ ;
	wire _w5168_ ;
	wire _w5167_ ;
	wire _w5166_ ;
	wire _w5165_ ;
	wire _w5164_ ;
	wire _w5163_ ;
	wire _w5162_ ;
	wire _w5161_ ;
	wire _w5160_ ;
	wire _w5159_ ;
	wire _w5158_ ;
	wire _w5157_ ;
	wire _w5156_ ;
	wire _w5155_ ;
	wire _w5154_ ;
	wire _w5153_ ;
	wire _w5152_ ;
	wire _w5151_ ;
	wire _w5150_ ;
	wire _w5149_ ;
	wire _w5148_ ;
	wire _w5147_ ;
	wire _w5146_ ;
	wire _w5145_ ;
	wire _w5144_ ;
	wire _w5143_ ;
	wire _w5142_ ;
	wire _w5141_ ;
	wire _w5140_ ;
	wire _w5139_ ;
	wire _w5138_ ;
	wire _w5137_ ;
	wire _w5136_ ;
	wire _w5135_ ;
	wire _w5134_ ;
	wire _w5133_ ;
	wire _w5132_ ;
	wire _w5131_ ;
	wire _w5130_ ;
	wire _w5129_ ;
	wire _w5128_ ;
	wire _w5127_ ;
	wire _w5126_ ;
	wire _w5125_ ;
	wire _w5124_ ;
	wire _w5123_ ;
	wire _w5122_ ;
	wire _w5121_ ;
	wire _w5120_ ;
	wire _w5119_ ;
	wire _w5118_ ;
	wire _w5117_ ;
	wire _w5116_ ;
	wire _w5115_ ;
	wire _w5114_ ;
	wire _w5113_ ;
	wire _w5112_ ;
	wire _w5111_ ;
	wire _w5110_ ;
	wire _w5109_ ;
	wire _w5108_ ;
	wire _w5107_ ;
	wire _w5106_ ;
	wire _w5105_ ;
	wire _w5104_ ;
	wire _w5103_ ;
	wire _w5102_ ;
	wire _w5101_ ;
	wire _w5100_ ;
	wire _w5099_ ;
	wire _w5098_ ;
	wire _w5097_ ;
	wire _w5096_ ;
	wire _w5095_ ;
	wire _w5094_ ;
	wire _w5093_ ;
	wire _w5092_ ;
	wire _w5091_ ;
	wire _w5090_ ;
	wire _w5089_ ;
	wire _w5088_ ;
	wire _w5087_ ;
	wire _w5086_ ;
	wire _w5085_ ;
	wire _w5084_ ;
	wire _w5083_ ;
	wire _w5082_ ;
	wire _w5081_ ;
	wire _w5080_ ;
	wire _w5079_ ;
	wire _w5078_ ;
	wire _w5077_ ;
	wire _w5076_ ;
	wire _w5075_ ;
	wire _w5074_ ;
	wire _w5073_ ;
	wire _w5072_ ;
	wire _w5071_ ;
	wire _w5070_ ;
	wire _w5069_ ;
	wire _w5068_ ;
	wire _w5067_ ;
	wire _w5066_ ;
	wire _w5065_ ;
	wire _w5064_ ;
	wire _w5063_ ;
	wire _w5062_ ;
	wire _w5061_ ;
	wire _w5060_ ;
	wire _w5059_ ;
	wire _w5058_ ;
	wire _w5057_ ;
	wire _w5056_ ;
	wire _w5055_ ;
	wire _w5054_ ;
	wire _w5053_ ;
	wire _w5052_ ;
	wire _w5051_ ;
	wire _w5050_ ;
	wire _w5049_ ;
	wire _w5048_ ;
	wire _w5047_ ;
	wire _w5046_ ;
	wire _w5045_ ;
	wire _w5044_ ;
	wire _w5043_ ;
	wire _w5042_ ;
	wire _w5041_ ;
	wire _w5040_ ;
	wire _w5039_ ;
	wire _w5038_ ;
	wire _w5037_ ;
	wire _w5036_ ;
	wire _w5035_ ;
	wire _w5034_ ;
	wire _w5033_ ;
	wire _w5032_ ;
	wire _w5031_ ;
	wire _w5030_ ;
	wire _w5029_ ;
	wire _w5028_ ;
	wire _w5027_ ;
	wire _w5026_ ;
	wire _w5025_ ;
	wire _w5024_ ;
	wire _w5023_ ;
	wire _w5022_ ;
	wire _w5021_ ;
	wire _w5020_ ;
	wire _w5019_ ;
	wire _w5018_ ;
	wire _w5017_ ;
	wire _w5016_ ;
	wire _w5015_ ;
	wire _w5014_ ;
	wire _w5013_ ;
	wire _w5012_ ;
	wire _w5011_ ;
	wire _w5010_ ;
	wire _w5009_ ;
	wire _w5008_ ;
	wire _w5007_ ;
	wire _w5006_ ;
	wire _w5005_ ;
	wire _w5004_ ;
	wire _w5003_ ;
	wire _w5002_ ;
	wire _w5001_ ;
	wire _w5000_ ;
	wire _w4999_ ;
	wire _w4998_ ;
	wire _w4997_ ;
	wire _w4996_ ;
	wire _w4995_ ;
	wire _w4994_ ;
	wire _w4993_ ;
	wire _w4992_ ;
	wire _w4991_ ;
	wire _w4990_ ;
	wire _w4989_ ;
	wire _w4988_ ;
	wire _w4987_ ;
	wire _w4986_ ;
	wire _w4985_ ;
	wire _w4984_ ;
	wire _w4983_ ;
	wire _w4982_ ;
	wire _w4981_ ;
	wire _w4980_ ;
	wire _w4979_ ;
	wire _w4978_ ;
	wire _w4977_ ;
	wire _w4976_ ;
	wire _w4975_ ;
	wire _w4974_ ;
	wire _w4973_ ;
	wire _w4972_ ;
	wire _w4971_ ;
	wire _w4970_ ;
	wire _w4969_ ;
	wire _w4968_ ;
	wire _w4967_ ;
	wire _w4966_ ;
	wire _w4965_ ;
	wire _w4964_ ;
	wire _w4963_ ;
	wire _w4962_ ;
	wire _w4961_ ;
	wire _w4960_ ;
	wire _w4959_ ;
	wire _w4958_ ;
	wire _w4957_ ;
	wire _w4956_ ;
	wire _w4955_ ;
	wire _w4954_ ;
	wire _w4953_ ;
	wire _w4952_ ;
	wire _w4951_ ;
	wire _w4950_ ;
	wire _w4949_ ;
	wire _w4948_ ;
	wire _w4947_ ;
	wire _w4946_ ;
	wire _w4945_ ;
	wire _w4944_ ;
	wire _w4943_ ;
	wire _w4942_ ;
	wire _w4941_ ;
	wire _w4940_ ;
	wire _w4939_ ;
	wire _w4938_ ;
	wire _w4937_ ;
	wire _w4936_ ;
	wire _w4935_ ;
	wire _w4934_ ;
	wire _w4933_ ;
	wire _w4932_ ;
	wire _w4931_ ;
	wire _w4930_ ;
	wire _w4929_ ;
	wire _w4928_ ;
	wire _w4927_ ;
	wire _w4926_ ;
	wire _w4925_ ;
	wire _w4924_ ;
	wire _w4923_ ;
	wire _w4922_ ;
	wire _w4921_ ;
	wire _w4920_ ;
	wire _w4919_ ;
	wire _w4918_ ;
	wire _w4917_ ;
	wire _w4916_ ;
	wire _w4915_ ;
	wire _w4914_ ;
	wire _w4913_ ;
	wire _w4912_ ;
	wire _w4911_ ;
	wire _w4910_ ;
	wire _w4909_ ;
	wire _w4908_ ;
	wire _w4907_ ;
	wire _w4906_ ;
	wire _w4905_ ;
	wire _w4904_ ;
	wire _w4903_ ;
	wire _w4902_ ;
	wire _w4901_ ;
	wire _w4900_ ;
	wire _w4899_ ;
	wire _w4898_ ;
	wire _w4897_ ;
	wire _w4896_ ;
	wire _w4895_ ;
	wire _w4894_ ;
	wire _w4893_ ;
	wire _w4892_ ;
	wire _w4891_ ;
	wire _w4890_ ;
	wire _w4889_ ;
	wire _w4888_ ;
	wire _w4887_ ;
	wire _w4886_ ;
	wire _w4885_ ;
	wire _w4884_ ;
	wire _w4883_ ;
	wire _w4882_ ;
	wire _w4881_ ;
	wire _w4880_ ;
	wire _w4879_ ;
	wire _w4878_ ;
	wire _w4877_ ;
	wire _w4876_ ;
	wire _w4875_ ;
	wire _w4874_ ;
	wire _w4873_ ;
	wire _w4872_ ;
	wire _w4871_ ;
	wire _w4870_ ;
	wire _w4869_ ;
	wire _w4868_ ;
	wire _w4867_ ;
	wire _w4866_ ;
	wire _w4865_ ;
	wire _w4864_ ;
	wire _w4863_ ;
	wire _w4862_ ;
	wire _w4861_ ;
	wire _w4860_ ;
	wire _w4859_ ;
	wire _w4858_ ;
	wire _w4857_ ;
	wire _w4856_ ;
	wire _w4855_ ;
	wire _w4854_ ;
	wire _w4853_ ;
	wire _w4852_ ;
	wire _w4851_ ;
	wire _w4850_ ;
	wire _w4849_ ;
	wire _w4848_ ;
	wire _w4847_ ;
	wire _w4846_ ;
	wire _w4845_ ;
	wire _w4844_ ;
	wire _w4843_ ;
	wire _w4842_ ;
	wire _w4841_ ;
	wire _w4840_ ;
	wire _w4839_ ;
	wire _w4838_ ;
	wire _w4837_ ;
	wire _w4836_ ;
	wire _w4835_ ;
	wire _w4834_ ;
	wire _w4833_ ;
	wire _w4832_ ;
	wire _w4831_ ;
	wire _w4830_ ;
	wire _w4829_ ;
	wire _w4828_ ;
	wire _w4827_ ;
	wire _w4826_ ;
	wire _w4825_ ;
	wire _w4824_ ;
	wire _w4823_ ;
	wire _w4822_ ;
	wire _w4821_ ;
	wire _w4820_ ;
	wire _w4819_ ;
	wire _w4818_ ;
	wire _w4817_ ;
	wire _w4816_ ;
	wire _w4815_ ;
	wire _w4814_ ;
	wire _w4813_ ;
	wire _w4812_ ;
	wire _w4811_ ;
	wire _w4810_ ;
	wire _w4809_ ;
	wire _w4808_ ;
	wire _w4807_ ;
	wire _w4806_ ;
	wire _w4805_ ;
	wire _w4804_ ;
	wire _w4803_ ;
	wire _w4802_ ;
	wire _w4801_ ;
	wire _w4800_ ;
	wire _w4799_ ;
	wire _w4798_ ;
	wire _w4797_ ;
	wire _w4796_ ;
	wire _w4795_ ;
	wire _w4794_ ;
	wire _w4793_ ;
	wire _w4792_ ;
	wire _w4791_ ;
	wire _w4790_ ;
	wire _w4789_ ;
	wire _w4788_ ;
	wire _w4787_ ;
	wire _w4786_ ;
	wire _w4785_ ;
	wire _w4784_ ;
	wire _w4783_ ;
	wire _w4782_ ;
	wire _w4781_ ;
	wire _w4780_ ;
	wire _w4779_ ;
	wire _w4778_ ;
	wire _w4777_ ;
	wire _w4776_ ;
	wire _w4775_ ;
	wire _w4774_ ;
	wire _w4773_ ;
	wire _w4772_ ;
	wire _w4771_ ;
	wire _w4770_ ;
	wire _w4769_ ;
	wire _w4768_ ;
	wire _w4767_ ;
	wire _w4766_ ;
	wire _w4765_ ;
	wire _w4764_ ;
	wire _w4763_ ;
	wire _w4762_ ;
	wire _w4761_ ;
	wire _w4760_ ;
	wire _w4759_ ;
	wire _w4758_ ;
	wire _w4757_ ;
	wire _w4756_ ;
	wire _w4755_ ;
	wire _w4754_ ;
	wire _w4753_ ;
	wire _w4752_ ;
	wire _w4751_ ;
	wire _w4750_ ;
	wire _w4749_ ;
	wire _w4748_ ;
	wire _w4747_ ;
	wire _w4746_ ;
	wire _w4745_ ;
	wire _w4744_ ;
	wire _w4743_ ;
	wire _w4742_ ;
	wire _w4741_ ;
	wire _w4740_ ;
	wire _w4739_ ;
	wire _w4738_ ;
	wire _w4737_ ;
	wire _w4736_ ;
	wire _w4735_ ;
	wire _w4734_ ;
	wire _w4733_ ;
	wire _w4732_ ;
	wire _w4731_ ;
	wire _w4730_ ;
	wire _w4729_ ;
	wire _w4728_ ;
	wire _w4727_ ;
	wire _w4726_ ;
	wire _w4725_ ;
	wire _w4724_ ;
	wire _w4723_ ;
	wire _w4722_ ;
	wire _w4721_ ;
	wire _w4720_ ;
	wire _w4719_ ;
	wire _w4718_ ;
	wire _w4717_ ;
	wire _w4716_ ;
	wire _w4715_ ;
	wire _w4714_ ;
	wire _w4713_ ;
	wire _w4712_ ;
	wire _w4711_ ;
	wire _w4710_ ;
	wire _w4709_ ;
	wire _w4708_ ;
	wire _w4707_ ;
	wire _w4706_ ;
	wire _w4705_ ;
	wire _w4704_ ;
	wire _w4703_ ;
	wire _w4702_ ;
	wire _w4701_ ;
	wire _w4700_ ;
	wire _w4699_ ;
	wire _w4698_ ;
	wire _w4697_ ;
	wire _w4696_ ;
	wire _w4695_ ;
	wire _w4694_ ;
	wire _w4693_ ;
	wire _w4692_ ;
	wire _w4691_ ;
	wire _w4690_ ;
	wire _w4689_ ;
	wire _w4688_ ;
	wire _w4687_ ;
	wire _w4686_ ;
	wire _w4685_ ;
	wire _w4684_ ;
	wire _w4683_ ;
	wire _w4682_ ;
	wire _w4681_ ;
	wire _w4680_ ;
	wire _w4679_ ;
	wire _w4678_ ;
	wire _w4677_ ;
	wire _w4676_ ;
	wire _w4675_ ;
	wire _w4674_ ;
	wire _w4673_ ;
	wire _w4672_ ;
	wire _w4671_ ;
	wire _w4670_ ;
	wire _w4669_ ;
	wire _w4668_ ;
	wire _w4667_ ;
	wire _w4666_ ;
	wire _w4665_ ;
	wire _w4664_ ;
	wire _w4663_ ;
	wire _w4662_ ;
	wire _w4661_ ;
	wire _w4660_ ;
	wire _w4659_ ;
	wire _w4658_ ;
	wire _w4657_ ;
	wire _w4656_ ;
	wire _w4655_ ;
	wire _w4654_ ;
	wire _w4653_ ;
	wire _w4652_ ;
	wire _w4651_ ;
	wire _w4650_ ;
	wire _w4649_ ;
	wire _w4648_ ;
	wire _w4647_ ;
	wire _w4646_ ;
	wire _w4645_ ;
	wire _w4644_ ;
	wire _w4643_ ;
	wire _w4642_ ;
	wire _w4641_ ;
	wire _w4640_ ;
	wire _w4639_ ;
	wire _w4638_ ;
	wire _w4637_ ;
	wire _w4636_ ;
	wire _w4635_ ;
	wire _w4634_ ;
	wire _w4633_ ;
	wire _w4632_ ;
	wire _w4631_ ;
	wire _w4630_ ;
	wire _w4629_ ;
	wire _w4628_ ;
	wire _w4627_ ;
	wire _w4626_ ;
	wire _w4625_ ;
	wire _w4624_ ;
	wire _w4623_ ;
	wire _w4622_ ;
	wire _w4621_ ;
	wire _w4620_ ;
	wire _w4619_ ;
	wire _w4618_ ;
	wire _w4617_ ;
	wire _w4616_ ;
	wire _w4615_ ;
	wire _w4614_ ;
	wire _w4613_ ;
	wire _w4612_ ;
	wire _w4611_ ;
	wire _w4610_ ;
	wire _w4609_ ;
	wire _w4608_ ;
	wire _w4607_ ;
	wire _w4606_ ;
	wire _w4605_ ;
	wire _w4604_ ;
	wire _w4603_ ;
	wire _w4602_ ;
	wire _w4601_ ;
	wire _w4600_ ;
	wire _w4599_ ;
	wire _w4598_ ;
	wire _w4597_ ;
	wire _w4596_ ;
	wire _w4595_ ;
	wire _w4594_ ;
	wire _w4593_ ;
	wire _w4592_ ;
	wire _w4591_ ;
	wire _w4590_ ;
	wire _w4589_ ;
	wire _w4588_ ;
	wire _w4587_ ;
	wire _w4586_ ;
	wire _w4585_ ;
	wire _w4584_ ;
	wire _w4583_ ;
	wire _w4582_ ;
	wire _w4581_ ;
	wire _w4580_ ;
	wire _w4579_ ;
	wire _w4578_ ;
	wire _w4577_ ;
	wire _w4576_ ;
	wire _w4575_ ;
	wire _w4574_ ;
	wire _w4573_ ;
	wire _w4572_ ;
	wire _w4571_ ;
	wire _w4570_ ;
	wire _w4569_ ;
	wire _w4568_ ;
	wire _w4567_ ;
	wire _w4566_ ;
	wire _w4565_ ;
	wire _w4564_ ;
	wire _w4563_ ;
	wire _w4562_ ;
	wire _w4561_ ;
	wire _w4560_ ;
	wire _w4559_ ;
	wire _w4558_ ;
	wire _w4557_ ;
	wire _w4556_ ;
	wire _w4555_ ;
	wire _w4554_ ;
	wire _w4553_ ;
	wire _w4552_ ;
	wire _w4551_ ;
	wire _w4550_ ;
	wire _w4549_ ;
	wire _w4548_ ;
	wire _w4547_ ;
	wire _w4546_ ;
	wire _w4545_ ;
	wire _w4544_ ;
	wire _w4543_ ;
	wire _w4542_ ;
	wire _w4541_ ;
	wire _w4540_ ;
	wire _w4539_ ;
	wire _w4538_ ;
	wire _w4537_ ;
	wire _w4536_ ;
	wire _w4535_ ;
	wire _w4534_ ;
	wire _w4533_ ;
	wire _w4532_ ;
	wire _w4531_ ;
	wire _w4530_ ;
	wire _w4529_ ;
	wire _w4528_ ;
	wire _w4527_ ;
	wire _w4526_ ;
	wire _w4525_ ;
	wire _w4524_ ;
	wire _w4523_ ;
	wire _w4522_ ;
	wire _w4521_ ;
	wire _w4520_ ;
	wire _w4519_ ;
	wire _w4518_ ;
	wire _w4517_ ;
	wire _w4516_ ;
	wire _w4515_ ;
	wire _w4514_ ;
	wire _w4513_ ;
	wire _w4512_ ;
	wire _w4511_ ;
	wire _w4510_ ;
	wire _w4509_ ;
	wire _w4508_ ;
	wire _w4507_ ;
	wire _w4506_ ;
	wire _w4505_ ;
	wire _w4504_ ;
	wire _w4503_ ;
	wire _w4502_ ;
	wire _w4501_ ;
	wire _w4500_ ;
	wire _w4499_ ;
	wire _w4498_ ;
	wire _w4497_ ;
	wire _w4496_ ;
	wire _w4495_ ;
	wire _w4494_ ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w5620_ ;
	wire _w5621_ ;
	wire _w5622_ ;
	wire _w5623_ ;
	wire _w5624_ ;
	wire _w5625_ ;
	wire _w5626_ ;
	wire _w5627_ ;
	wire _w5628_ ;
	wire _w5629_ ;
	wire _w5630_ ;
	wire _w5631_ ;
	wire _w5632_ ;
	wire _w5633_ ;
	wire _w5634_ ;
	wire _w5635_ ;
	wire _w5636_ ;
	wire _w5637_ ;
	wire _w5638_ ;
	wire _w5639_ ;
	wire _w5640_ ;
	wire _w5641_ ;
	wire _w5642_ ;
	wire _w5643_ ;
	wire _w5644_ ;
	wire _w5645_ ;
	wire _w5646_ ;
	wire _w5647_ ;
	wire _w5648_ ;
	wire _w5649_ ;
	wire _w5650_ ;
	wire _w5651_ ;
	wire _w5652_ ;
	wire _w5653_ ;
	wire _w5654_ ;
	wire _w5655_ ;
	wire _w5656_ ;
	wire _w5657_ ;
	wire _w5658_ ;
	wire _w5659_ ;
	wire _w5660_ ;
	wire _w5661_ ;
	wire _w5662_ ;
	wire _w5663_ ;
	wire _w5664_ ;
	wire _w5665_ ;
	wire _w5666_ ;
	wire _w5667_ ;
	wire _w5668_ ;
	wire _w5669_ ;
	wire _w5670_ ;
	wire _w5671_ ;
	wire _w5672_ ;
	wire _w5673_ ;
	wire _w5674_ ;
	wire _w5675_ ;
	wire _w5676_ ;
	wire _w5677_ ;
	wire _w5678_ ;
	wire _w5679_ ;
	wire _w5680_ ;
	wire _w5681_ ;
	wire _w5682_ ;
	wire _w5683_ ;
	wire _w5684_ ;
	wire _w5685_ ;
	wire _w5686_ ;
	wire _w5687_ ;
	wire _w5688_ ;
	wire _w5689_ ;
	wire _w5690_ ;
	wire _w5691_ ;
	wire _w5692_ ;
	wire _w5693_ ;
	wire _w5694_ ;
	wire _w5695_ ;
	wire _w5696_ ;
	wire _w5697_ ;
	wire _w5698_ ;
	wire _w5699_ ;
	wire _w5700_ ;
	wire _w5701_ ;
	wire _w5702_ ;
	wire _w5703_ ;
	wire _w5704_ ;
	wire _w5705_ ;
	wire _w5706_ ;
	wire _w5707_ ;
	wire _w5708_ ;
	wire _w5709_ ;
	wire _w5710_ ;
	wire _w5711_ ;
	wire _w5712_ ;
	wire _w5713_ ;
	wire _w5714_ ;
	wire _w5715_ ;
	wire _w5716_ ;
	wire _w5717_ ;
	wire _w5718_ ;
	wire _w5719_ ;
	wire _w5720_ ;
	wire _w5721_ ;
	wire _w5722_ ;
	wire _w5723_ ;
	wire _w5724_ ;
	wire _w5725_ ;
	wire _w5726_ ;
	wire _w5727_ ;
	wire _w5728_ ;
	wire _w5729_ ;
	wire _w5730_ ;
	wire _w5731_ ;
	wire _w5732_ ;
	wire _w5733_ ;
	wire _w5734_ ;
	wire _w5735_ ;
	wire _w5736_ ;
	wire _w5737_ ;
	wire _w5738_ ;
	wire _w5739_ ;
	wire _w5740_ ;
	wire _w5741_ ;
	wire _w5742_ ;
	wire _w5743_ ;
	wire _w5744_ ;
	wire _w5745_ ;
	wire _w5746_ ;
	wire _w5747_ ;
	wire _w5748_ ;
	wire _w5749_ ;
	wire _w5750_ ;
	wire _w5751_ ;
	wire _w5752_ ;
	wire _w5753_ ;
	wire _w5754_ ;
	wire _w5755_ ;
	wire _w5756_ ;
	wire _w5757_ ;
	wire _w5758_ ;
	wire _w5759_ ;
	wire _w5760_ ;
	wire _w5761_ ;
	wire _w5762_ ;
	wire _w5763_ ;
	wire _w5764_ ;
	wire _w5765_ ;
	wire _w5766_ ;
	wire _w5767_ ;
	wire _w5768_ ;
	wire _w5769_ ;
	wire _w5770_ ;
	wire _w5771_ ;
	wire _w5772_ ;
	wire _w5773_ ;
	wire _w5774_ ;
	wire _w5775_ ;
	wire _w5776_ ;
	wire _w5777_ ;
	wire _w5778_ ;
	wire _w5779_ ;
	wire _w5780_ ;
	wire _w5781_ ;
	wire _w5782_ ;
	wire _w5783_ ;
	wire _w5784_ ;
	wire _w5785_ ;
	wire _w5786_ ;
	wire _w5787_ ;
	wire _w5788_ ;
	wire _w5789_ ;
	wire _w5790_ ;
	wire _w5791_ ;
	wire _w5792_ ;
	wire _w5793_ ;
	wire _w5794_ ;
	wire _w5795_ ;
	wire _w5796_ ;
	wire _w5797_ ;
	wire _w5798_ ;
	wire _w5799_ ;
	wire _w5800_ ;
	wire _w5801_ ;
	wire _w5802_ ;
	wire _w5803_ ;
	wire _w5804_ ;
	wire _w5805_ ;
	wire _w5806_ ;
	wire _w5807_ ;
	wire _w5808_ ;
	wire _w5809_ ;
	wire _w5810_ ;
	wire _w5811_ ;
	wire _w5812_ ;
	wire _w5813_ ;
	wire _w5814_ ;
	wire _w5815_ ;
	wire _w5816_ ;
	wire _w5817_ ;
	wire _w5818_ ;
	wire _w5819_ ;
	wire _w5820_ ;
	wire _w5821_ ;
	wire _w5822_ ;
	wire _w5823_ ;
	wire _w5824_ ;
	wire _w5825_ ;
	wire _w5826_ ;
	wire _w5827_ ;
	wire _w5828_ ;
	wire _w5829_ ;
	wire _w5830_ ;
	wire _w5831_ ;
	wire _w5832_ ;
	wire _w5833_ ;
	wire _w5834_ ;
	wire _w5835_ ;
	wire _w5836_ ;
	wire _w5837_ ;
	wire _w5838_ ;
	wire _w5839_ ;
	wire _w5840_ ;
	wire _w5841_ ;
	wire _w5842_ ;
	wire _w5843_ ;
	wire _w5844_ ;
	wire _w5845_ ;
	wire _w5846_ ;
	wire _w5847_ ;
	wire _w5848_ ;
	wire _w5849_ ;
	wire _w5850_ ;
	wire _w5851_ ;
	wire _w5852_ ;
	wire _w5853_ ;
	wire _w5854_ ;
	wire _w5855_ ;
	wire _w5856_ ;
	wire _w5857_ ;
	wire _w5858_ ;
	wire _w5859_ ;
	wire _w5860_ ;
	wire _w5861_ ;
	wire _w5862_ ;
	wire _w5863_ ;
	wire _w5864_ ;
	wire _w5865_ ;
	wire _w5866_ ;
	wire _w5867_ ;
	wire _w5868_ ;
	wire _w5869_ ;
	wire _w5870_ ;
	wire _w5871_ ;
	wire _w5872_ ;
	wire _w5873_ ;
	wire _w5874_ ;
	wire _w5875_ ;
	wire _w5876_ ;
	wire _w5877_ ;
	wire _w5878_ ;
	wire _w5879_ ;
	wire _w5880_ ;
	wire _w5881_ ;
	wire _w5882_ ;
	wire _w5883_ ;
	wire _w5884_ ;
	wire _w5885_ ;
	wire _w5886_ ;
	wire _w5887_ ;
	wire _w5888_ ;
	wire _w5889_ ;
	wire _w5890_ ;
	wire _w5891_ ;
	wire _w5892_ ;
	wire _w5893_ ;
	wire _w5894_ ;
	wire _w5895_ ;
	wire _w5896_ ;
	wire _w5897_ ;
	wire _w5898_ ;
	wire _w5899_ ;
	wire _w5900_ ;
	wire _w5901_ ;
	wire _w5902_ ;
	wire _w5903_ ;
	wire _w5904_ ;
	wire _w5905_ ;
	wire _w5906_ ;
	wire _w5907_ ;
	wire _w5908_ ;
	wire _w5909_ ;
	wire _w5910_ ;
	wire _w5911_ ;
	wire _w5912_ ;
	wire _w5913_ ;
	wire _w5914_ ;
	wire _w5915_ ;
	wire _w5916_ ;
	wire _w5917_ ;
	wire _w5918_ ;
	wire _w5919_ ;
	wire _w5920_ ;
	wire _w5921_ ;
	wire _w5922_ ;
	wire _w5923_ ;
	wire _w5924_ ;
	wire _w5925_ ;
	wire _w5926_ ;
	wire _w5927_ ;
	wire _w5928_ ;
	wire _w5929_ ;
	wire _w5930_ ;
	wire _w5931_ ;
	wire _w5932_ ;
	wire _w5933_ ;
	wire _w5934_ ;
	wire _w5935_ ;
	wire _w5936_ ;
	wire _w5937_ ;
	wire _w5938_ ;
	wire _w5939_ ;
	wire _w5940_ ;
	wire _w5941_ ;
	wire _w5942_ ;
	wire _w5943_ ;
	wire _w5944_ ;
	wire _w5945_ ;
	wire _w5946_ ;
	wire _w5947_ ;
	wire _w5948_ ;
	wire _w5949_ ;
	wire _w5950_ ;
	wire _w5951_ ;
	wire _w5952_ ;
	wire _w5953_ ;
	wire _w5954_ ;
	wire _w5955_ ;
	wire _w5956_ ;
	wire _w5957_ ;
	wire _w5958_ ;
	wire _w5959_ ;
	wire _w5960_ ;
	wire _w5961_ ;
	wire _w5962_ ;
	wire _w5963_ ;
	wire _w5964_ ;
	wire _w5965_ ;
	wire _w5966_ ;
	wire _w5967_ ;
	wire _w5968_ ;
	wire _w5969_ ;
	wire _w5970_ ;
	wire _w5971_ ;
	wire _w5972_ ;
	wire _w5973_ ;
	wire _w5974_ ;
	wire _w5975_ ;
	wire _w5976_ ;
	wire _w5977_ ;
	wire _w5978_ ;
	wire _w5979_ ;
	wire _w5980_ ;
	wire _w5981_ ;
	wire _w5982_ ;
	wire _w5983_ ;
	wire _w5984_ ;
	wire _w5985_ ;
	wire _w5986_ ;
	wire _w5987_ ;
	wire _w5988_ ;
	wire _w5989_ ;
	wire _w5990_ ;
	wire _w5991_ ;
	wire _w5992_ ;
	wire _w5993_ ;
	wire _w5994_ ;
	wire _w5995_ ;
	wire _w5996_ ;
	wire _w5997_ ;
	wire _w5998_ ;
	wire _w5999_ ;
	wire _w6000_ ;
	wire _w6001_ ;
	wire _w6002_ ;
	wire _w6003_ ;
	wire _w6004_ ;
	wire _w6005_ ;
	wire _w6006_ ;
	wire _w6007_ ;
	wire _w6008_ ;
	wire _w6009_ ;
	wire _w6010_ ;
	wire _w6011_ ;
	wire _w6012_ ;
	wire _w6013_ ;
	wire _w6014_ ;
	wire _w6015_ ;
	wire _w6016_ ;
	wire _w6017_ ;
	wire _w6018_ ;
	wire _w6019_ ;
	wire _w6020_ ;
	wire _w6021_ ;
	wire _w6022_ ;
	wire _w6023_ ;
	wire _w6024_ ;
	wire _w6025_ ;
	wire _w6026_ ;
	wire _w6027_ ;
	wire _w6028_ ;
	wire _w6029_ ;
	wire _w6030_ ;
	wire _w6031_ ;
	wire _w6032_ ;
	wire _w6033_ ;
	wire _w6034_ ;
	wire _w6035_ ;
	wire _w6036_ ;
	wire _w6037_ ;
	wire _w6038_ ;
	wire _w6039_ ;
	wire _w6040_ ;
	wire _w6041_ ;
	wire _w6042_ ;
	wire _w6043_ ;
	wire _w6044_ ;
	wire _w6045_ ;
	wire _w6046_ ;
	wire _w6047_ ;
	wire _w6048_ ;
	wire _w6049_ ;
	wire _w6050_ ;
	wire _w6051_ ;
	wire _w6052_ ;
	wire _w6053_ ;
	wire _w6054_ ;
	wire _w6055_ ;
	wire _w6056_ ;
	wire _w6057_ ;
	wire _w6058_ ;
	wire _w6059_ ;
	wire _w6060_ ;
	wire _w6061_ ;
	wire _w6062_ ;
	wire _w6063_ ;
	wire _w6064_ ;
	wire _w6065_ ;
	wire _w6066_ ;
	wire _w6067_ ;
	wire _w6068_ ;
	wire _w6069_ ;
	wire _w6070_ ;
	wire _w6071_ ;
	wire _w6072_ ;
	wire _w6073_ ;
	wire _w6074_ ;
	wire _w6075_ ;
	wire _w6076_ ;
	wire _w6077_ ;
	wire _w6078_ ;
	wire _w6079_ ;
	wire _w6080_ ;
	wire _w6081_ ;
	wire _w6082_ ;
	wire _w6083_ ;
	wire _w6084_ ;
	wire _w6085_ ;
	wire _w6086_ ;
	wire _w6087_ ;
	wire _w6088_ ;
	wire _w6089_ ;
	wire _w6090_ ;
	wire _w6091_ ;
	wire _w6092_ ;
	wire _w6093_ ;
	wire _w6094_ ;
	wire _w6095_ ;
	wire _w6096_ ;
	wire _w6097_ ;
	wire _w6098_ ;
	wire _w6099_ ;
	wire _w6100_ ;
	wire _w6101_ ;
	wire _w6102_ ;
	wire _w6103_ ;
	wire _w6104_ ;
	wire _w6105_ ;
	wire _w6106_ ;
	wire _w6107_ ;
	wire _w6108_ ;
	wire _w6109_ ;
	wire _w6110_ ;
	wire _w6111_ ;
	wire _w6112_ ;
	wire _w6113_ ;
	wire _w6114_ ;
	wire _w6115_ ;
	wire _w6116_ ;
	wire _w6117_ ;
	wire _w6118_ ;
	wire _w6119_ ;
	wire _w6120_ ;
	wire _w6121_ ;
	wire _w6122_ ;
	wire _w6123_ ;
	wire _w6124_ ;
	wire _w6125_ ;
	wire _w6126_ ;
	wire _w6127_ ;
	wire _w6128_ ;
	wire _w6129_ ;
	wire _w6130_ ;
	wire _w6131_ ;
	wire _w6132_ ;
	wire _w6133_ ;
	wire _w6134_ ;
	wire _w6135_ ;
	wire _w6136_ ;
	wire _w6137_ ;
	wire _w6138_ ;
	wire _w6139_ ;
	wire _w6140_ ;
	wire _w6141_ ;
	wire _w6142_ ;
	wire _w6143_ ;
	wire _w6144_ ;
	wire _w6145_ ;
	wire _w6146_ ;
	wire _w6147_ ;
	wire _w6148_ ;
	wire _w6149_ ;
	wire _w6150_ ;
	wire _w6151_ ;
	wire _w6152_ ;
	wire _w6153_ ;
	wire _w6154_ ;
	wire _w6155_ ;
	wire _w6156_ ;
	wire _w6157_ ;
	wire _w6158_ ;
	wire _w6159_ ;
	wire _w6160_ ;
	wire _w6161_ ;
	wire _w6162_ ;
	wire _w6163_ ;
	wire _w6164_ ;
	wire _w6165_ ;
	wire _w6166_ ;
	wire _w6167_ ;
	wire _w6168_ ;
	wire _w6169_ ;
	wire _w6170_ ;
	wire _w6171_ ;
	wire _w6172_ ;
	wire _w6173_ ;
	wire _w6174_ ;
	wire _w6175_ ;
	wire _w6176_ ;
	wire _w6177_ ;
	wire _w6178_ ;
	wire _w6179_ ;
	wire _w6180_ ;
	wire _w6181_ ;
	wire _w6182_ ;
	wire _w6183_ ;
	wire _w6184_ ;
	wire _w6185_ ;
	wire _w6186_ ;
	wire _w6187_ ;
	wire _w6188_ ;
	wire _w6189_ ;
	wire _w6190_ ;
	wire _w6191_ ;
	wire _w6192_ ;
	wire _w6193_ ;
	wire _w6194_ ;
	wire _w6195_ ;
	wire _w6196_ ;
	wire _w6197_ ;
	wire _w6198_ ;
	wire _w6199_ ;
	wire _w6200_ ;
	wire _w6201_ ;
	wire _w6202_ ;
	wire _w6203_ ;
	wire _w6204_ ;
	wire _w6205_ ;
	wire _w6206_ ;
	wire _w6207_ ;
	wire _w6208_ ;
	wire _w6209_ ;
	wire _w6210_ ;
	wire _w6211_ ;
	wire _w6212_ ;
	wire _w6213_ ;
	wire _w6214_ ;
	wire _w6215_ ;
	wire _w6216_ ;
	wire _w6217_ ;
	wire _w6218_ ;
	wire _w6219_ ;
	wire _w6220_ ;
	wire _w6221_ ;
	wire _w6222_ ;
	wire _w6223_ ;
	wire _w6224_ ;
	wire _w6225_ ;
	wire _w6226_ ;
	wire _w6227_ ;
	wire _w6228_ ;
	wire _w6229_ ;
	wire _w6230_ ;
	wire _w6231_ ;
	wire _w6232_ ;
	wire _w6233_ ;
	wire _w6234_ ;
	wire _w6235_ ;
	wire _w6236_ ;
	wire _w6237_ ;
	wire _w6238_ ;
	wire _w6239_ ;
	wire _w6240_ ;
	wire _w6241_ ;
	wire _w6242_ ;
	wire _w6243_ ;
	wire _w6244_ ;
	wire _w6245_ ;
	wire _w6246_ ;
	wire _w6247_ ;
	wire _w6248_ ;
	wire _w6249_ ;
	wire _w6250_ ;
	wire _w6251_ ;
	wire _w6252_ ;
	wire _w6253_ ;
	wire _w6254_ ;
	wire _w6255_ ;
	wire _w6256_ ;
	wire _w6257_ ;
	wire _w6258_ ;
	wire _w6259_ ;
	wire _w6260_ ;
	wire _w6261_ ;
	wire _w6262_ ;
	wire _w6263_ ;
	wire _w6264_ ;
	wire _w6265_ ;
	wire _w6266_ ;
	wire _w6267_ ;
	wire _w6268_ ;
	wire _w6269_ ;
	wire _w6270_ ;
	wire _w6271_ ;
	wire _w6272_ ;
	wire _w6273_ ;
	wire _w6274_ ;
	wire _w6275_ ;
	wire _w6276_ ;
	wire _w6277_ ;
	wire _w6278_ ;
	wire _w6279_ ;
	wire _w6280_ ;
	wire _w6281_ ;
	wire _w6282_ ;
	wire _w6283_ ;
	wire _w6284_ ;
	wire _w6285_ ;
	wire _w6286_ ;
	wire _w6287_ ;
	wire _w6288_ ;
	wire _w6289_ ;
	wire _w6290_ ;
	wire _w6291_ ;
	wire _w6292_ ;
	wire _w6293_ ;
	wire _w6294_ ;
	wire _w6295_ ;
	wire _w6296_ ;
	wire _w6297_ ;
	wire _w6298_ ;
	wire _w6299_ ;
	wire _w6300_ ;
	wire _w6301_ ;
	wire _w6302_ ;
	wire _w6303_ ;
	wire _w6304_ ;
	wire _w6305_ ;
	wire _w6306_ ;
	wire _w6307_ ;
	wire _w6308_ ;
	wire _w6309_ ;
	wire _w6310_ ;
	wire _w6311_ ;
	wire _w6312_ ;
	wire _w6313_ ;
	wire _w6314_ ;
	wire _w6315_ ;
	wire _w6316_ ;
	wire _w6317_ ;
	wire _w6318_ ;
	wire _w6319_ ;
	wire _w6320_ ;
	wire _w6321_ ;
	wire _w6322_ ;
	wire _w6323_ ;
	wire _w6324_ ;
	wire _w6325_ ;
	wire _w6326_ ;
	wire _w6327_ ;
	wire _w6328_ ;
	wire _w6329_ ;
	wire _w6330_ ;
	wire _w6331_ ;
	wire _w6332_ ;
	wire _w6333_ ;
	wire _w6334_ ;
	wire _w6335_ ;
	wire _w6336_ ;
	wire _w6337_ ;
	wire _w6338_ ;
	wire _w6339_ ;
	wire _w6340_ ;
	wire _w6341_ ;
	wire _w6342_ ;
	wire _w6343_ ;
	wire _w6344_ ;
	wire _w6345_ ;
	wire _w6346_ ;
	wire _w6347_ ;
	wire _w6348_ ;
	wire _w6349_ ;
	wire _w6350_ ;
	wire _w6351_ ;
	wire _w6352_ ;
	wire _w6353_ ;
	wire _w6354_ ;
	wire _w6355_ ;
	wire _w6356_ ;
	wire _w6357_ ;
	wire _w6358_ ;
	wire _w6359_ ;
	wire _w6360_ ;
	wire _w6361_ ;
	wire _w6362_ ;
	wire _w6363_ ;
	wire _w6364_ ;
	wire _w6365_ ;
	wire _w6366_ ;
	wire _w6367_ ;
	wire _w6368_ ;
	wire _w6369_ ;
	wire _w6370_ ;
	wire _w6371_ ;
	wire _w6372_ ;
	wire _w6373_ ;
	wire _w6374_ ;
	wire _w6375_ ;
	wire _w6376_ ;
	wire _w6377_ ;
	wire _w6378_ ;
	wire _w6379_ ;
	wire _w6380_ ;
	wire _w6381_ ;
	wire _w6382_ ;
	wire _w6383_ ;
	wire _w6384_ ;
	wire _w6385_ ;
	wire _w6386_ ;
	wire _w6387_ ;
	wire _w6388_ ;
	wire _w6389_ ;
	wire _w6390_ ;
	wire _w6391_ ;
	wire _w6392_ ;
	wire _w6393_ ;
	wire _w6394_ ;
	wire _w6395_ ;
	wire _w6396_ ;
	wire _w6397_ ;
	wire _w6398_ ;
	wire _w6399_ ;
	wire _w6400_ ;
	wire _w6401_ ;
	wire _w6402_ ;
	wire _w6403_ ;
	wire _w6404_ ;
	wire _w6405_ ;
	wire _w6406_ ;
	wire _w6407_ ;
	wire _w6408_ ;
	wire _w6409_ ;
	wire _w6410_ ;
	wire _w6411_ ;
	wire _w6412_ ;
	wire _w6413_ ;
	wire _w6414_ ;
	wire _w6415_ ;
	wire _w6416_ ;
	wire _w6417_ ;
	wire _w6418_ ;
	wire _w6419_ ;
	wire _w6420_ ;
	wire _w6421_ ;
	wire _w6422_ ;
	wire _w6423_ ;
	wire _w6424_ ;
	wire _w6425_ ;
	wire _w6426_ ;
	wire _w6427_ ;
	wire _w6428_ ;
	wire _w6429_ ;
	wire _w6430_ ;
	wire _w6431_ ;
	wire _w6432_ ;
	wire _w6433_ ;
	wire _w6434_ ;
	wire _w6435_ ;
	wire _w6436_ ;
	wire _w6437_ ;
	wire _w6438_ ;
	wire _w6439_ ;
	wire _w6440_ ;
	wire _w6441_ ;
	wire _w6442_ ;
	wire _w6443_ ;
	wire _w6444_ ;
	wire _w6445_ ;
	wire _w6446_ ;
	wire _w6447_ ;
	wire _w6448_ ;
	wire _w6449_ ;
	wire _w6450_ ;
	wire _w6451_ ;
	wire _w6452_ ;
	wire _w6453_ ;
	wire _w6454_ ;
	wire _w6455_ ;
	wire _w6456_ ;
	wire _w6457_ ;
	wire _w6458_ ;
	wire _w6459_ ;
	wire _w6460_ ;
	wire _w6461_ ;
	wire _w6462_ ;
	wire _w6463_ ;
	wire _w6464_ ;
	wire _w6465_ ;
	wire _w6466_ ;
	wire _w6467_ ;
	wire _w6468_ ;
	wire _w6469_ ;
	wire _w6470_ ;
	wire _w6471_ ;
	wire _w6472_ ;
	wire _w6473_ ;
	wire _w6474_ ;
	wire _w6475_ ;
	wire _w6476_ ;
	wire _w6477_ ;
	wire _w6478_ ;
	wire _w6479_ ;
	wire _w6480_ ;
	wire _w6481_ ;
	wire _w6482_ ;
	wire _w6483_ ;
	wire _w6484_ ;
	wire _w6485_ ;
	wire _w6486_ ;
	wire _w6487_ ;
	wire _w6488_ ;
	wire _w6489_ ;
	wire _w6490_ ;
	wire _w6491_ ;
	wire _w6492_ ;
	wire _w6493_ ;
	wire _w6494_ ;
	wire _w6495_ ;
	wire _w6496_ ;
	wire _w6497_ ;
	wire _w6498_ ;
	wire _w6499_ ;
	wire _w6500_ ;
	wire _w6501_ ;
	wire _w6502_ ;
	wire _w6503_ ;
	wire _w6504_ ;
	wire _w6505_ ;
	wire _w6506_ ;
	wire _w6507_ ;
	wire _w6508_ ;
	wire _w6509_ ;
	wire _w6510_ ;
	wire _w6511_ ;
	wire _w6512_ ;
	wire _w6513_ ;
	wire _w6514_ ;
	wire _w6515_ ;
	wire _w6516_ ;
	wire _w6517_ ;
	wire _w6518_ ;
	wire _w6519_ ;
	wire _w6520_ ;
	wire _w6521_ ;
	wire _w6522_ ;
	wire _w6523_ ;
	wire _w6524_ ;
	wire _w6525_ ;
	wire _w6526_ ;
	wire _w6527_ ;
	wire _w6528_ ;
	wire _w6529_ ;
	wire _w6530_ ;
	wire _w6531_ ;
	wire _w6532_ ;
	wire _w6533_ ;
	wire _w6534_ ;
	wire _w6535_ ;
	wire _w6536_ ;
	wire _w6537_ ;
	wire _w6538_ ;
	wire _w6539_ ;
	wire _w6540_ ;
	wire _w6541_ ;
	wire _w6542_ ;
	wire _w6543_ ;
	wire _w6544_ ;
	wire _w6545_ ;
	wire _w6546_ ;
	wire _w6547_ ;
	wire _w6548_ ;
	wire _w6549_ ;
	wire _w6550_ ;
	wire _w6551_ ;
	wire _w6552_ ;
	wire _w6553_ ;
	wire _w6554_ ;
	wire _w6555_ ;
	wire _w6556_ ;
	wire _w6557_ ;
	wire _w6558_ ;
	wire _w6559_ ;
	wire _w6560_ ;
	wire _w6561_ ;
	wire _w6562_ ;
	wire _w6563_ ;
	wire _w6564_ ;
	wire _w6565_ ;
	wire _w6566_ ;
	wire _w6567_ ;
	wire _w6568_ ;
	wire _w6569_ ;
	wire _w6570_ ;
	wire _w6571_ ;
	wire _w6572_ ;
	wire _w6573_ ;
	wire _w6574_ ;
	wire _w6575_ ;
	wire _w6576_ ;
	wire _w6577_ ;
	wire _w6578_ ;
	wire _w6579_ ;
	wire _w6580_ ;
	wire _w6581_ ;
	wire _w6582_ ;
	wire _w6583_ ;
	wire _w6584_ ;
	wire _w6585_ ;
	wire _w6586_ ;
	wire _w6587_ ;
	wire _w6588_ ;
	wire _w6589_ ;
	wire _w6590_ ;
	wire _w6591_ ;
	wire _w6592_ ;
	wire _w6593_ ;
	wire _w6594_ ;
	wire _w6595_ ;
	wire _w6596_ ;
	wire _w6597_ ;
	wire _w6598_ ;
	wire _w6599_ ;
	wire _w6600_ ;
	wire _w6601_ ;
	wire _w6602_ ;
	wire _w6603_ ;
	wire _w6604_ ;
	wire _w6605_ ;
	wire _w6606_ ;
	wire _w6607_ ;
	wire _w6608_ ;
	wire _w6609_ ;
	wire _w6610_ ;
	wire _w6611_ ;
	wire _w6612_ ;
	wire _w6613_ ;
	wire _w6614_ ;
	wire _w6615_ ;
	wire _w6616_ ;
	wire _w6617_ ;
	wire _w6618_ ;
	wire _w6619_ ;
	wire _w6620_ ;
	wire _w6621_ ;
	wire _w6622_ ;
	wire _w6623_ ;
	wire _w6624_ ;
	wire _w6625_ ;
	wire _w6626_ ;
	wire _w6627_ ;
	wire _w6628_ ;
	wire _w6629_ ;
	wire _w6630_ ;
	wire _w6631_ ;
	wire _w6632_ ;
	wire _w6633_ ;
	wire _w6634_ ;
	wire _w6635_ ;
	wire _w6636_ ;
	wire _w6637_ ;
	wire _w6638_ ;
	wire _w6639_ ;
	wire _w6640_ ;
	wire _w6641_ ;
	wire _w6642_ ;
	wire _w6643_ ;
	wire _w6644_ ;
	wire _w6645_ ;
	wire _w6646_ ;
	wire _w6647_ ;
	wire _w6648_ ;
	wire _w6649_ ;
	wire _w6650_ ;
	wire _w6651_ ;
	wire _w6652_ ;
	wire _w6653_ ;
	wire _w6654_ ;
	wire _w6655_ ;
	wire _w6656_ ;
	wire _w6657_ ;
	wire _w6658_ ;
	wire _w6659_ ;
	wire _w6660_ ;
	wire _w6661_ ;
	wire _w6662_ ;
	wire _w6663_ ;
	wire _w6664_ ;
	wire _w6665_ ;
	wire _w6666_ ;
	wire _w6667_ ;
	wire _w6668_ ;
	wire _w6669_ ;
	wire _w6670_ ;
	wire _w6671_ ;
	wire _w6672_ ;
	wire _w6673_ ;
	wire _w6674_ ;
	wire _w6675_ ;
	wire _w6676_ ;
	wire _w6677_ ;
	wire _w6678_ ;
	wire _w6679_ ;
	wire _w6680_ ;
	wire _w6681_ ;
	wire _w6682_ ;
	wire _w6683_ ;
	wire _w6684_ ;
	wire _w6685_ ;
	wire _w6686_ ;
	wire _w6687_ ;
	wire _w6688_ ;
	wire _w6689_ ;
	wire _w6690_ ;
	wire _w6691_ ;
	wire _w6692_ ;
	wire _w6693_ ;
	wire _w6694_ ;
	wire _w6695_ ;
	wire _w6696_ ;
	wire _w6697_ ;
	wire _w6698_ ;
	wire _w6699_ ;
	wire _w6700_ ;
	wire _w6701_ ;
	wire _w6702_ ;
	wire _w6703_ ;
	wire _w6704_ ;
	wire _w6705_ ;
	wire _w6706_ ;
	wire _w6707_ ;
	wire _w6708_ ;
	wire _w6709_ ;
	wire _w6710_ ;
	wire _w6711_ ;
	wire _w6712_ ;
	wire _w6713_ ;
	wire _w6714_ ;
	wire _w6715_ ;
	wire _w6716_ ;
	wire _w6717_ ;
	wire _w6718_ ;
	wire _w6719_ ;
	wire _w6720_ ;
	wire _w6721_ ;
	wire _w6722_ ;
	wire _w6723_ ;
	wire _w6724_ ;
	wire _w6725_ ;
	wire _w6726_ ;
	wire _w6727_ ;
	wire _w6728_ ;
	wire _w6729_ ;
	wire _w6730_ ;
	wire _w6731_ ;
	wire _w6732_ ;
	wire _w6733_ ;
	wire _w6734_ ;
	wire _w6735_ ;
	wire _w6736_ ;
	wire _w6737_ ;
	wire _w6738_ ;
	wire _w6739_ ;
	wire _w6740_ ;
	wire _w6741_ ;
	wire _w6742_ ;
	wire _w6743_ ;
	wire _w6744_ ;
	wire _w6745_ ;
	wire _w6746_ ;
	wire _w6747_ ;
	wire _w6748_ ;
	wire _w6749_ ;
	wire _w6750_ ;
	wire _w6751_ ;
	wire _w6752_ ;
	wire _w6753_ ;
	wire _w6754_ ;
	wire _w6755_ ;
	wire _w6756_ ;
	wire _w6757_ ;
	wire _w6758_ ;
	wire _w6759_ ;
	wire _w6760_ ;
	wire _w6761_ ;
	wire _w6762_ ;
	wire _w6763_ ;
	wire _w6764_ ;
	wire _w6765_ ;
	wire _w6766_ ;
	wire _w6767_ ;
	wire _w6768_ ;
	wire _w6769_ ;
	wire _w6770_ ;
	wire _w6771_ ;
	wire _w6772_ ;
	wire _w6773_ ;
	wire _w6774_ ;
	wire _w6775_ ;
	wire _w6776_ ;
	wire _w6777_ ;
	wire _w6778_ ;
	wire _w6779_ ;
	wire _w6780_ ;
	wire _w6781_ ;
	wire _w6782_ ;
	wire _w6783_ ;
	wire _w6784_ ;
	wire _w6785_ ;
	wire _w6786_ ;
	wire _w6787_ ;
	wire _w6788_ ;
	wire _w6789_ ;
	wire _w6790_ ;
	wire _w6791_ ;
	wire _w6792_ ;
	wire _w6793_ ;
	wire _w6794_ ;
	wire _w6795_ ;
	wire _w6796_ ;
	wire _w6797_ ;
	wire _w6798_ ;
	wire _w6799_ ;
	wire _w6800_ ;
	wire _w6801_ ;
	wire _w6802_ ;
	wire _w6803_ ;
	wire _w6804_ ;
	wire _w6805_ ;
	wire _w6806_ ;
	wire _w6807_ ;
	wire _w6808_ ;
	wire _w6809_ ;
	wire _w6810_ ;
	wire _w6811_ ;
	wire _w6812_ ;
	wire _w6813_ ;
	wire _w6814_ ;
	wire _w6815_ ;
	wire _w6816_ ;
	wire _w6817_ ;
	wire _w6818_ ;
	wire _w6819_ ;
	wire _w6820_ ;
	wire _w6821_ ;
	wire _w6822_ ;
	wire _w6823_ ;
	wire _w6824_ ;
	wire _w6825_ ;
	wire _w6826_ ;
	wire _w6827_ ;
	wire _w6828_ ;
	wire _w6829_ ;
	wire _w6830_ ;
	wire _w6831_ ;
	wire _w6832_ ;
	wire _w6833_ ;
	wire _w6834_ ;
	wire _w6835_ ;
	wire _w6836_ ;
	wire _w6837_ ;
	wire _w6838_ ;
	wire _w6839_ ;
	wire _w6840_ ;
	wire _w6841_ ;
	wire _w6842_ ;
	wire _w6843_ ;
	wire _w6844_ ;
	wire _w6845_ ;
	wire _w6846_ ;
	wire _w6847_ ;
	wire _w6848_ ;
	wire _w6849_ ;
	wire _w6850_ ;
	wire _w6851_ ;
	wire _w6852_ ;
	wire _w6853_ ;
	wire _w6854_ ;
	wire _w6855_ ;
	wire _w6856_ ;
	wire _w6857_ ;
	wire _w6858_ ;
	wire _w6859_ ;
	wire _w6860_ ;
	wire _w6861_ ;
	wire _w6862_ ;
	wire _w6863_ ;
	wire _w6864_ ;
	wire _w6865_ ;
	wire _w6866_ ;
	wire _w6867_ ;
	wire _w6868_ ;
	wire _w6869_ ;
	wire _w6870_ ;
	wire _w6871_ ;
	wire _w6872_ ;
	wire _w6873_ ;
	wire _w6874_ ;
	wire _w6875_ ;
	wire _w6876_ ;
	wire _w6877_ ;
	wire _w6878_ ;
	wire _w6879_ ;
	wire _w6880_ ;
	wire _w6881_ ;
	wire _w6882_ ;
	wire _w6883_ ;
	wire _w6884_ ;
	wire _w6885_ ;
	wire _w6886_ ;
	wire _w6887_ ;
	wire _w6888_ ;
	wire _w6889_ ;
	wire _w6890_ ;
	wire _w6891_ ;
	wire _w6892_ ;
	wire _w6893_ ;
	wire _w6894_ ;
	wire _w6895_ ;
	wire _w6896_ ;
	wire _w6897_ ;
	wire _w6898_ ;
	wire _w6899_ ;
	wire _w6900_ ;
	wire _w6901_ ;
	wire _w6902_ ;
	wire _w6903_ ;
	wire _w6904_ ;
	wire _w6905_ ;
	wire _w6906_ ;
	wire _w6907_ ;
	wire _w6908_ ;
	wire _w6909_ ;
	wire _w6910_ ;
	wire _w6911_ ;
	wire _w6912_ ;
	wire _w6913_ ;
	wire _w6914_ ;
	wire _w6915_ ;
	wire _w6916_ ;
	wire _w6917_ ;
	wire _w6918_ ;
	wire _w6919_ ;
	wire _w6920_ ;
	wire _w6921_ ;
	wire _w6922_ ;
	wire _w6923_ ;
	wire _w6924_ ;
	wire _w6925_ ;
	wire _w6926_ ;
	wire _w6927_ ;
	wire _w6928_ ;
	wire _w6929_ ;
	wire _w6930_ ;
	wire _w6931_ ;
	wire _w6932_ ;
	wire _w6933_ ;
	wire _w6934_ ;
	wire _w6935_ ;
	wire _w6936_ ;
	wire _w6937_ ;
	wire _w6938_ ;
	wire _w6939_ ;
	wire _w6940_ ;
	wire _w6941_ ;
	wire _w6942_ ;
	wire _w6943_ ;
	wire _w6944_ ;
	wire _w6945_ ;
	wire _w6946_ ;
	wire _w6947_ ;
	wire _w6948_ ;
	wire _w6949_ ;
	wire _w6950_ ;
	wire _w6951_ ;
	wire _w6952_ ;
	wire _w6953_ ;
	wire _w6954_ ;
	wire _w6955_ ;
	wire _w6956_ ;
	wire _w6957_ ;
	wire _w6958_ ;
	wire _w6959_ ;
	wire _w6960_ ;
	wire _w6961_ ;
	wire _w6962_ ;
	wire _w6963_ ;
	wire _w6964_ ;
	wire _w6965_ ;
	wire _w6966_ ;
	wire _w6967_ ;
	wire _w6968_ ;
	wire _w6969_ ;
	wire _w6970_ ;
	wire _w6971_ ;
	wire _w6972_ ;
	wire _w6973_ ;
	wire _w6974_ ;
	wire _w6975_ ;
	wire _w6976_ ;
	wire _w6977_ ;
	wire _w6978_ ;
	wire _w6979_ ;
	wire _w6980_ ;
	wire _w6981_ ;
	wire _w6982_ ;
	wire _w6983_ ;
	wire _w6984_ ;
	wire _w6985_ ;
	wire _w6986_ ;
	wire _w6987_ ;
	wire _w6988_ ;
	wire _w6989_ ;
	wire _w6990_ ;
	wire _w6991_ ;
	wire _w6992_ ;
	wire _w6993_ ;
	wire _w6994_ ;
	wire _w6995_ ;
	wire _w6996_ ;
	wire _w6997_ ;
	wire _w6998_ ;
	wire _w6999_ ;
	wire _w7000_ ;
	wire _w7001_ ;
	wire _w7002_ ;
	wire _w7003_ ;
	wire _w7004_ ;
	wire _w7005_ ;
	wire _w7006_ ;
	wire _w7007_ ;
	wire _w7008_ ;
	wire _w7009_ ;
	wire _w7010_ ;
	wire _w7011_ ;
	wire _w7012_ ;
	wire _w7013_ ;
	wire _w7014_ ;
	wire _w7015_ ;
	wire _w7016_ ;
	wire _w7017_ ;
	wire _w7018_ ;
	wire _w7019_ ;
	wire _w7020_ ;
	wire _w7021_ ;
	wire _w7022_ ;
	wire _w7023_ ;
	wire _w7024_ ;
	wire _w7025_ ;
	wire _w7026_ ;
	wire _w7027_ ;
	wire _w7028_ ;
	wire _w7029_ ;
	wire _w7030_ ;
	wire _w7031_ ;
	wire _w7032_ ;
	wire _w7033_ ;
	wire _w7034_ ;
	wire _w7035_ ;
	wire _w7036_ ;
	wire _w7037_ ;
	wire _w7038_ ;
	wire _w7039_ ;
	wire _w7040_ ;
	wire _w7041_ ;
	wire _w7042_ ;
	wire _w7043_ ;
	wire _w7044_ ;
	wire _w7045_ ;
	wire _w7046_ ;
	wire _w7047_ ;
	wire _w7048_ ;
	wire _w7049_ ;
	wire _w7050_ ;
	wire _w7051_ ;
	wire _w7052_ ;
	wire _w7053_ ;
	wire _w7054_ ;
	wire _w7055_ ;
	wire _w7056_ ;
	wire _w7057_ ;
	wire _w7058_ ;
	wire _w7059_ ;
	wire _w7060_ ;
	wire _w7061_ ;
	wire _w7062_ ;
	wire _w7063_ ;
	wire _w7064_ ;
	wire _w7065_ ;
	wire _w7066_ ;
	wire _w7067_ ;
	wire _w7068_ ;
	wire _w7069_ ;
	wire _w7070_ ;
	wire _w7071_ ;
	wire _w7072_ ;
	wire _w7073_ ;
	wire _w7074_ ;
	wire _w7075_ ;
	wire _w7076_ ;
	wire _w7077_ ;
	wire _w7078_ ;
	wire _w7079_ ;
	wire _w7080_ ;
	wire _w7081_ ;
	wire _w7082_ ;
	wire _w7083_ ;
	wire _w7084_ ;
	wire _w7085_ ;
	wire _w7086_ ;
	wire _w7087_ ;
	wire _w7088_ ;
	wire _w7089_ ;
	wire _w7090_ ;
	wire _w7091_ ;
	wire _w7092_ ;
	wire _w7093_ ;
	wire _w7094_ ;
	wire _w7095_ ;
	wire _w7096_ ;
	wire _w7097_ ;
	wire _w7098_ ;
	wire _w7099_ ;
	wire _w7100_ ;
	wire _w7101_ ;
	wire _w7102_ ;
	wire _w7103_ ;
	wire _w7104_ ;
	wire _w7105_ ;
	wire _w7106_ ;
	wire _w7107_ ;
	wire _w7108_ ;
	wire _w7109_ ;
	wire _w7110_ ;
	wire _w7111_ ;
	wire _w7112_ ;
	wire _w7113_ ;
	wire _w7114_ ;
	wire _w7115_ ;
	wire _w7116_ ;
	wire _w7117_ ;
	wire _w7118_ ;
	wire _w7119_ ;
	wire _w7120_ ;
	wire _w7121_ ;
	wire _w7122_ ;
	wire _w7123_ ;
	wire _w7124_ ;
	wire _w7125_ ;
	wire _w7126_ ;
	wire _w7127_ ;
	wire _w7128_ ;
	wire _w7129_ ;
	wire _w7130_ ;
	wire _w7131_ ;
	wire _w7132_ ;
	wire _w7133_ ;
	wire _w7134_ ;
	wire _w7135_ ;
	wire _w7136_ ;
	wire _w7137_ ;
	wire _w7138_ ;
	wire _w7139_ ;
	wire _w7140_ ;
	wire _w7141_ ;
	wire _w7142_ ;
	wire _w7143_ ;
	wire _w7144_ ;
	wire _w7145_ ;
	wire _w7146_ ;
	wire _w7147_ ;
	wire _w7148_ ;
	wire _w7149_ ;
	wire _w7150_ ;
	wire _w7151_ ;
	wire _w7152_ ;
	wire _w7153_ ;
	wire _w7154_ ;
	wire _w7155_ ;
	wire _w7156_ ;
	wire _w7157_ ;
	wire _w7158_ ;
	wire _w7159_ ;
	wire _w7160_ ;
	wire _w7161_ ;
	wire _w7162_ ;
	wire _w7163_ ;
	wire _w7164_ ;
	wire _w7165_ ;
	wire _w7166_ ;
	wire _w7167_ ;
	wire _w7168_ ;
	wire _w7169_ ;
	wire _w7170_ ;
	wire _w7171_ ;
	wire _w7172_ ;
	wire _w7173_ ;
	wire _w7174_ ;
	wire _w7175_ ;
	wire _w7176_ ;
	wire _w7177_ ;
	wire _w7178_ ;
	wire _w7179_ ;
	wire _w7180_ ;
	wire _w7181_ ;
	wire _w7182_ ;
	wire _w7183_ ;
	wire _w7184_ ;
	wire _w7185_ ;
	wire _w7186_ ;
	wire _w7187_ ;
	wire _w7188_ ;
	wire _w7189_ ;
	wire _w7190_ ;
	wire _w7191_ ;
	wire _w7192_ ;
	wire _w7193_ ;
	wire _w7194_ ;
	wire _w7195_ ;
	wire _w7196_ ;
	wire _w7197_ ;
	wire _w7198_ ;
	wire _w7199_ ;
	wire _w7200_ ;
	wire _w7201_ ;
	wire _w7202_ ;
	wire _w7203_ ;
	wire _w7204_ ;
	wire _w7205_ ;
	wire _w7206_ ;
	wire _w7207_ ;
	wire _w7208_ ;
	wire _w7209_ ;
	wire _w7210_ ;
	wire _w7211_ ;
	wire _w7212_ ;
	wire _w7213_ ;
	wire _w7214_ ;
	wire _w7215_ ;
	wire _w7216_ ;
	wire _w7217_ ;
	wire _w7218_ ;
	wire _w7219_ ;
	wire _w7220_ ;
	wire _w7221_ ;
	wire _w7222_ ;
	wire _w7223_ ;
	wire _w7224_ ;
	wire _w7225_ ;
	wire _w7226_ ;
	wire _w7227_ ;
	wire _w7228_ ;
	wire _w7229_ ;
	wire _w7230_ ;
	wire _w7231_ ;
	wire _w7232_ ;
	wire _w7233_ ;
	wire _w7234_ ;
	wire _w7235_ ;
	wire _w7236_ ;
	wire _w7237_ ;
	wire _w7238_ ;
	wire _w7239_ ;
	wire _w7240_ ;
	wire _w7241_ ;
	wire _w7242_ ;
	wire _w7243_ ;
	wire _w7244_ ;
	wire _w7245_ ;
	wire _w7246_ ;
	wire _w7247_ ;
	wire _w7248_ ;
	wire _w7249_ ;
	wire _w7250_ ;
	wire _w7251_ ;
	wire _w7252_ ;
	wire _w7253_ ;
	wire _w7254_ ;
	wire _w7255_ ;
	wire _w7256_ ;
	wire _w7257_ ;
	wire _w7258_ ;
	wire _w7259_ ;
	wire _w7260_ ;
	wire _w7261_ ;
	wire _w7262_ ;
	wire _w7263_ ;
	wire _w7264_ ;
	wire _w7265_ ;
	wire _w7266_ ;
	wire _w7267_ ;
	wire _w7268_ ;
	wire _w7269_ ;
	wire _w7270_ ;
	wire _w7271_ ;
	wire _w7272_ ;
	wire _w7273_ ;
	wire _w7274_ ;
	wire _w7275_ ;
	wire _w7276_ ;
	wire _w7277_ ;
	wire _w7278_ ;
	wire _w7279_ ;
	wire _w7280_ ;
	wire _w7281_ ;
	wire _w7282_ ;
	wire _w7283_ ;
	wire _w7284_ ;
	wire _w7285_ ;
	wire _w7286_ ;
	wire _w7287_ ;
	wire _w7288_ ;
	wire _w7289_ ;
	wire _w7290_ ;
	wire _w7291_ ;
	wire _w7292_ ;
	wire _w7293_ ;
	wire _w7294_ ;
	wire _w7295_ ;
	wire _w7296_ ;
	wire _w7297_ ;
	wire _w7298_ ;
	wire _w7299_ ;
	wire _w7300_ ;
	wire _w7301_ ;
	wire _w7302_ ;
	wire _w7303_ ;
	wire _w7304_ ;
	wire _w7305_ ;
	wire _w7306_ ;
	wire _w7307_ ;
	wire _w7308_ ;
	wire _w7309_ ;
	wire _w7310_ ;
	wire _w7311_ ;
	wire _w7312_ ;
	wire _w7313_ ;
	wire _w7314_ ;
	wire _w7315_ ;
	wire _w7316_ ;
	wire _w7317_ ;
	wire _w7318_ ;
	wire _w7319_ ;
	wire _w7320_ ;
	wire _w7321_ ;
	wire _w7322_ ;
	wire _w7323_ ;
	wire _w7324_ ;
	wire _w7325_ ;
	wire _w7326_ ;
	wire _w7327_ ;
	wire _w7328_ ;
	wire _w7329_ ;
	wire _w7330_ ;
	wire _w7331_ ;
	wire _w7332_ ;
	wire _w7333_ ;
	wire _w7334_ ;
	wire _w7335_ ;
	wire _w7336_ ;
	wire _w7337_ ;
	wire _w7338_ ;
	wire _w7339_ ;
	wire _w7340_ ;
	wire _w7341_ ;
	wire _w7342_ ;
	wire _w7343_ ;
	wire _w7344_ ;
	wire _w7345_ ;
	wire _w7346_ ;
	wire _w7347_ ;
	wire _w7348_ ;
	wire _w7349_ ;
	wire _w7350_ ;
	wire _w7351_ ;
	wire _w7352_ ;
	wire _w7353_ ;
	wire _w7354_ ;
	wire _w7355_ ;
	wire _w7356_ ;
	wire _w7357_ ;
	wire _w7358_ ;
	wire _w7359_ ;
	wire _w7360_ ;
	wire _w7361_ ;
	wire _w7362_ ;
	wire _w7363_ ;
	wire _w7364_ ;
	wire _w7365_ ;
	wire _w7366_ ;
	wire _w7367_ ;
	wire _w7368_ ;
	wire _w7369_ ;
	wire _w7370_ ;
	wire _w7371_ ;
	wire _w7372_ ;
	wire _w7373_ ;
	wire _w7374_ ;
	wire _w7375_ ;
	wire _w7376_ ;
	wire _w7377_ ;
	wire _w7378_ ;
	wire _w7379_ ;
	wire _w7380_ ;
	wire _w7381_ ;
	wire _w7382_ ;
	wire _w7383_ ;
	wire _w7384_ ;
	wire _w7385_ ;
	wire _w7386_ ;
	wire _w7387_ ;
	wire _w7388_ ;
	wire _w7389_ ;
	wire _w7390_ ;
	wire _w7391_ ;
	wire _w7392_ ;
	wire _w7393_ ;
	wire _w7394_ ;
	wire _w7395_ ;
	wire _w7396_ ;
	wire _w7397_ ;
	wire _w7398_ ;
	wire _w7399_ ;
	wire _w7400_ ;
	wire _w7401_ ;
	wire _w7402_ ;
	wire _w7403_ ;
	wire _w7404_ ;
	wire _w7405_ ;
	wire _w7406_ ;
	wire _w7407_ ;
	wire _w7408_ ;
	wire _w7409_ ;
	wire _w7410_ ;
	wire _w7411_ ;
	wire _w7412_ ;
	wire _w7413_ ;
	wire _w7414_ ;
	wire _w7415_ ;
	wire _w7416_ ;
	wire _w7417_ ;
	wire _w7418_ ;
	wire _w7419_ ;
	wire _w7420_ ;
	wire _w7421_ ;
	wire _w7422_ ;
	wire _w7423_ ;
	wire _w7424_ ;
	wire _w7425_ ;
	wire _w7426_ ;
	wire _w7427_ ;
	wire _w7428_ ;
	wire _w7429_ ;
	wire _w7430_ ;
	wire _w7431_ ;
	wire _w7432_ ;
	wire _w7433_ ;
	wire _w7434_ ;
	wire _w7435_ ;
	wire _w7436_ ;
	wire _w7437_ ;
	wire _w7438_ ;
	wire _w7439_ ;
	wire _w7440_ ;
	wire _w7441_ ;
	wire _w7442_ ;
	wire _w7443_ ;
	wire _w7444_ ;
	wire _w7445_ ;
	wire _w7446_ ;
	wire _w7447_ ;
	wire _w7448_ ;
	wire _w7449_ ;
	wire _w7450_ ;
	wire _w7451_ ;
	wire _w7452_ ;
	wire _w7453_ ;
	wire _w7454_ ;
	wire _w7455_ ;
	wire _w7456_ ;
	wire _w7457_ ;
	wire _w7458_ ;
	wire _w7459_ ;
	wire _w7460_ ;
	wire _w7461_ ;
	wire _w7462_ ;
	wire _w7463_ ;
	wire _w7464_ ;
	wire _w7465_ ;
	wire _w7466_ ;
	wire _w7467_ ;
	wire _w7468_ ;
	wire _w7469_ ;
	wire _w7470_ ;
	wire _w7471_ ;
	wire _w7472_ ;
	wire _w7473_ ;
	wire _w7474_ ;
	wire _w7475_ ;
	wire _w7476_ ;
	wire _w7477_ ;
	wire _w7478_ ;
	wire _w7479_ ;
	wire _w7480_ ;
	wire _w7481_ ;
	wire _w7482_ ;
	wire _w7483_ ;
	wire _w7484_ ;
	wire _w7485_ ;
	wire _w7486_ ;
	wire _w7487_ ;
	wire _w7488_ ;
	wire _w7489_ ;
	wire _w7490_ ;
	wire _w7491_ ;
	wire _w7492_ ;
	wire _w7493_ ;
	wire _w7494_ ;
	wire _w7495_ ;
	wire _w7496_ ;
	wire _w7497_ ;
	wire _w7498_ ;
	wire _w7499_ ;
	wire _w7500_ ;
	wire _w7501_ ;
	wire _w7502_ ;
	wire _w7503_ ;
	wire _w7504_ ;
	wire _w7505_ ;
	wire _w7506_ ;
	wire _w7507_ ;
	wire _w7508_ ;
	wire _w7509_ ;
	wire _w7510_ ;
	wire _w7511_ ;
	wire _w7512_ ;
	wire _w7513_ ;
	wire _w7514_ ;
	wire _w7515_ ;
	wire _w7516_ ;
	wire _w7517_ ;
	wire _w7518_ ;
	wire _w7519_ ;
	wire _w7520_ ;
	wire _w7521_ ;
	wire _w7522_ ;
	wire _w7523_ ;
	wire _w7524_ ;
	wire _w7525_ ;
	wire _w7526_ ;
	wire _w7527_ ;
	wire _w7528_ ;
	wire _w7529_ ;
	wire _w7530_ ;
	wire _w7531_ ;
	wire _w7532_ ;
	wire _w7533_ ;
	wire _w7534_ ;
	wire _w7535_ ;
	wire _w7536_ ;
	wire _w7537_ ;
	wire _w7538_ ;
	wire _w7539_ ;
	wire _w7540_ ;
	wire _w7541_ ;
	wire _w7542_ ;
	wire _w7543_ ;
	wire _w7544_ ;
	wire _w7545_ ;
	wire _w7546_ ;
	wire _w7547_ ;
	wire _w7548_ ;
	wire _w7549_ ;
	wire _w7550_ ;
	wire _w7551_ ;
	wire _w7552_ ;
	wire _w7553_ ;
	wire _w7554_ ;
	wire _w7555_ ;
	wire _w7556_ ;
	wire _w7557_ ;
	wire _w7558_ ;
	wire _w7559_ ;
	wire _w7560_ ;
	wire _w7561_ ;
	wire _w7562_ ;
	wire _w7563_ ;
	wire _w7564_ ;
	wire _w7565_ ;
	wire _w7566_ ;
	wire _w7567_ ;
	wire _w7568_ ;
	wire _w7569_ ;
	wire _w7570_ ;
	wire _w7571_ ;
	wire _w7572_ ;
	wire _w7573_ ;
	wire _w7574_ ;
	wire _w7575_ ;
	wire _w7576_ ;
	wire _w7577_ ;
	wire _w7578_ ;
	wire _w7579_ ;
	wire _w7580_ ;
	wire _w7581_ ;
	wire _w7582_ ;
	wire _w7583_ ;
	wire _w7584_ ;
	wire _w7585_ ;
	wire _w7586_ ;
	wire _w7587_ ;
	wire _w7588_ ;
	wire _w7589_ ;
	wire _w7590_ ;
	wire _w7591_ ;
	wire _w7592_ ;
	wire _w7593_ ;
	wire _w7594_ ;
	wire _w7595_ ;
	wire _w7596_ ;
	wire _w7597_ ;
	wire _w7598_ ;
	wire _w7599_ ;
	wire _w7600_ ;
	wire _w7601_ ;
	wire _w7602_ ;
	wire _w7603_ ;
	wire _w7604_ ;
	wire _w7605_ ;
	wire _w7606_ ;
	wire _w7607_ ;
	wire _w7608_ ;
	wire _w7609_ ;
	wire _w7610_ ;
	wire _w7611_ ;
	wire _w7612_ ;
	wire _w7613_ ;
	wire _w7614_ ;
	wire _w7615_ ;
	wire _w7616_ ;
	wire _w7617_ ;
	wire _w7618_ ;
	wire _w7619_ ;
	wire _w7620_ ;
	wire _w7621_ ;
	wire _w7622_ ;
	wire _w7623_ ;
	wire _w7624_ ;
	wire _w7625_ ;
	wire _w7626_ ;
	wire _w7627_ ;
	wire _w7628_ ;
	wire _w7629_ ;
	wire _w7630_ ;
	wire _w7631_ ;
	wire _w7632_ ;
	wire _w7633_ ;
	wire _w7634_ ;
	wire _w7635_ ;
	wire _w7636_ ;
	wire _w7637_ ;
	wire _w7638_ ;
	wire _w7639_ ;
	wire _w7640_ ;
	wire _w7641_ ;
	wire _w7642_ ;
	wire _w7643_ ;
	wire _w7644_ ;
	wire _w7645_ ;
	wire _w7646_ ;
	wire _w7647_ ;
	wire _w7648_ ;
	wire _w7649_ ;
	wire _w7650_ ;
	wire _w7651_ ;
	wire _w7652_ ;
	wire _w7653_ ;
	wire _w7654_ ;
	wire _w7655_ ;
	wire _w7656_ ;
	wire _w7657_ ;
	wire _w7658_ ;
	wire _w7659_ ;
	wire _w7660_ ;
	wire _w7661_ ;
	wire _w7662_ ;
	wire _w7663_ ;
	wire _w7664_ ;
	wire _w7665_ ;
	wire _w7666_ ;
	wire _w7667_ ;
	wire _w7668_ ;
	wire _w7669_ ;
	wire _w7670_ ;
	wire _w7671_ ;
	wire _w7672_ ;
	wire _w7673_ ;
	wire _w7674_ ;
	wire _w7675_ ;
	wire _w7676_ ;
	wire _w7677_ ;
	wire _w7678_ ;
	wire _w7679_ ;
	wire _w7680_ ;
	wire _w7681_ ;
	wire _w7682_ ;
	wire _w7683_ ;
	wire _w7684_ ;
	wire _w7685_ ;
	wire _w7686_ ;
	wire _w7687_ ;
	wire _w7688_ ;
	wire _w7689_ ;
	wire _w7690_ ;
	wire _w7691_ ;
	wire _w7692_ ;
	wire _w7693_ ;
	wire _w7694_ ;
	wire _w7695_ ;
	wire _w7696_ ;
	wire _w7697_ ;
	wire _w7698_ ;
	wire _w7699_ ;
	wire _w7700_ ;
	wire _w7701_ ;
	wire _w7702_ ;
	wire _w7703_ ;
	wire _w7704_ ;
	wire _w7705_ ;
	wire _w7706_ ;
	wire _w7707_ ;
	wire _w7708_ ;
	wire _w7709_ ;
	wire _w7710_ ;
	wire _w7711_ ;
	wire _w7712_ ;
	wire _w7713_ ;
	wire _w7714_ ;
	wire _w7715_ ;
	wire _w7716_ ;
	wire _w7717_ ;
	wire _w7718_ ;
	wire _w7719_ ;
	wire _w7720_ ;
	wire _w7721_ ;
	wire _w7722_ ;
	wire _w7723_ ;
	wire _w7724_ ;
	wire _w7725_ ;
	wire _w7726_ ;
	wire _w7727_ ;
	wire _w7728_ ;
	wire _w7729_ ;
	wire _w7730_ ;
	wire _w7731_ ;
	wire _w7732_ ;
	wire _w7733_ ;
	wire _w7734_ ;
	wire _w7735_ ;
	wire _w7736_ ;
	wire _w7737_ ;
	wire _w7738_ ;
	wire _w7739_ ;
	wire _w7740_ ;
	wire _w7741_ ;
	wire _w7742_ ;
	wire _w7743_ ;
	wire _w7744_ ;
	wire _w7745_ ;
	wire _w7746_ ;
	wire _w7747_ ;
	wire _w7748_ ;
	wire _w7749_ ;
	wire _w7750_ ;
	wire _w7751_ ;
	wire _w7752_ ;
	wire _w7753_ ;
	wire _w7754_ ;
	wire _w7755_ ;
	wire _w7756_ ;
	wire _w7757_ ;
	wire _w7758_ ;
	wire _w7759_ ;
	wire _w7760_ ;
	wire _w7761_ ;
	wire _w7762_ ;
	wire _w7763_ ;
	wire _w7764_ ;
	wire _w7765_ ;
	wire _w7766_ ;
	wire _w7767_ ;
	wire _w7768_ ;
	wire _w7769_ ;
	wire _w7770_ ;
	wire _w7771_ ;
	wire _w7772_ ;
	wire _w7773_ ;
	wire _w7774_ ;
	wire _w7775_ ;
	wire _w7776_ ;
	wire _w7777_ ;
	wire _w7778_ ;
	wire _w7779_ ;
	wire _w7780_ ;
	wire _w7781_ ;
	wire _w7782_ ;
	wire _w7783_ ;
	wire _w7784_ ;
	wire _w7785_ ;
	wire _w7786_ ;
	wire _w7787_ ;
	wire _w7788_ ;
	wire _w7789_ ;
	wire _w7790_ ;
	wire _w7791_ ;
	wire _w7792_ ;
	wire _w7793_ ;
	wire _w7794_ ;
	wire _w7795_ ;
	wire _w7796_ ;
	wire _w7797_ ;
	wire _w7798_ ;
	wire _w7799_ ;
	wire _w7800_ ;
	wire _w7801_ ;
	wire _w7802_ ;
	wire _w7803_ ;
	wire _w7804_ ;
	wire _w7805_ ;
	wire _w7806_ ;
	wire _w7807_ ;
	wire _w7808_ ;
	wire _w7809_ ;
	wire _w7810_ ;
	wire _w7811_ ;
	wire _w7812_ ;
	wire _w7813_ ;
	wire _w7814_ ;
	wire _w7815_ ;
	wire _w7816_ ;
	wire _w7817_ ;
	wire _w7818_ ;
	wire _w7819_ ;
	wire _w7820_ ;
	wire _w7821_ ;
	wire _w7822_ ;
	wire _w7823_ ;
	wire _w7824_ ;
	wire _w7825_ ;
	wire _w7826_ ;
	wire _w7827_ ;
	wire _w7828_ ;
	wire _w7829_ ;
	wire _w7830_ ;
	wire _w7831_ ;
	wire _w7832_ ;
	wire _w7833_ ;
	wire _w7834_ ;
	wire _w7835_ ;
	wire _w7836_ ;
	wire _w7837_ ;
	wire _w7838_ ;
	wire _w7839_ ;
	wire _w7840_ ;
	wire _w7841_ ;
	wire _w7842_ ;
	wire _w7843_ ;
	wire _w7844_ ;
	wire _w7845_ ;
	wire _w7846_ ;
	wire _w7847_ ;
	wire _w7848_ ;
	wire _w7849_ ;
	wire _w7850_ ;
	wire _w7851_ ;
	wire _w7852_ ;
	wire _w7853_ ;
	wire _w7854_ ;
	wire _w7855_ ;
	wire _w7856_ ;
	wire _w7857_ ;
	wire _w7858_ ;
	wire _w7859_ ;
	wire _w7860_ ;
	wire _w7861_ ;
	wire _w7862_ ;
	wire _w7863_ ;
	wire _w7864_ ;
	wire _w7865_ ;
	wire _w7866_ ;
	wire _w7867_ ;
	wire _w7868_ ;
	wire _w7869_ ;
	wire _w7870_ ;
	wire _w7871_ ;
	wire _w7872_ ;
	wire _w7873_ ;
	wire _w7874_ ;
	wire _w7875_ ;
	wire _w7876_ ;
	wire _w7877_ ;
	wire _w7878_ ;
	wire _w7879_ ;
	wire _w7880_ ;
	wire _w7881_ ;
	wire _w7882_ ;
	wire _w7883_ ;
	wire _w7884_ ;
	wire _w7885_ ;
	wire _w7886_ ;
	wire _w7887_ ;
	wire _w7888_ ;
	wire _w7889_ ;
	wire _w7890_ ;
	wire _w7891_ ;
	wire _w7892_ ;
	wire _w7893_ ;
	wire _w7894_ ;
	wire _w7895_ ;
	wire _w7896_ ;
	wire _w7897_ ;
	wire _w7898_ ;
	wire _w7899_ ;
	wire _w7900_ ;
	wire _w7901_ ;
	wire _w7902_ ;
	wire _w7903_ ;
	wire _w7904_ ;
	wire _w7905_ ;
	wire _w7906_ ;
	wire _w7907_ ;
	wire _w7908_ ;
	wire _w7909_ ;
	wire _w7910_ ;
	wire _w7911_ ;
	wire _w7912_ ;
	wire _w7913_ ;
	wire _w7914_ ;
	wire _w7915_ ;
	wire _w7916_ ;
	wire _w7917_ ;
	wire _w7918_ ;
	wire _w7919_ ;
	wire _w7920_ ;
	wire _w7921_ ;
	wire _w7922_ ;
	wire _w7923_ ;
	wire _w7924_ ;
	wire _w7925_ ;
	wire _w7926_ ;
	wire _w7927_ ;
	wire _w7928_ ;
	wire _w7929_ ;
	wire _w7930_ ;
	wire _w7931_ ;
	wire _w7932_ ;
	wire _w7933_ ;
	wire _w7934_ ;
	wire _w7935_ ;
	wire _w7936_ ;
	wire _w7937_ ;
	wire _w7938_ ;
	wire _w7939_ ;
	wire _w7940_ ;
	wire _w7941_ ;
	wire _w7942_ ;
	wire _w7943_ ;
	wire _w7944_ ;
	wire _w7945_ ;
	wire _w7946_ ;
	wire _w7947_ ;
	wire _w7948_ ;
	wire _w7949_ ;
	wire _w7950_ ;
	wire _w7951_ ;
	wire _w7952_ ;
	wire _w7953_ ;
	wire _w7954_ ;
	wire _w7955_ ;
	wire _w7956_ ;
	wire _w7957_ ;
	wire _w7958_ ;
	wire _w7959_ ;
	wire _w7960_ ;
	wire _w7961_ ;
	wire _w7962_ ;
	wire _w7963_ ;
	wire _w7964_ ;
	wire _w7965_ ;
	wire _w7966_ ;
	wire _w7967_ ;
	wire _w7968_ ;
	wire _w7969_ ;
	wire _w7970_ ;
	wire _w7971_ ;
	wire _w7972_ ;
	wire _w7973_ ;
	wire _w7974_ ;
	wire _w7975_ ;
	wire _w7976_ ;
	wire _w7977_ ;
	wire _w7978_ ;
	wire _w7979_ ;
	wire _w7980_ ;
	wire _w7981_ ;
	wire _w7982_ ;
	wire _w7983_ ;
	wire _w7984_ ;
	wire _w7985_ ;
	wire _w7986_ ;
	wire _w7987_ ;
	wire _w7988_ ;
	wire _w7989_ ;
	wire _w7990_ ;
	wire _w7991_ ;
	wire _w7992_ ;
	wire _w7993_ ;
	wire _w7994_ ;
	wire _w7995_ ;
	wire _w7996_ ;
	wire _w7997_ ;
	wire _w7998_ ;
	wire _w7999_ ;
	wire _w8000_ ;
	wire _w8001_ ;
	wire _w8002_ ;
	wire _w8003_ ;
	wire _w8004_ ;
	wire _w8005_ ;
	wire _w8006_ ;
	wire _w8007_ ;
	wire _w8008_ ;
	wire _w8009_ ;
	wire _w8010_ ;
	wire _w8011_ ;
	wire _w8012_ ;
	wire _w8013_ ;
	wire _w8014_ ;
	wire _w8015_ ;
	wire _w8016_ ;
	wire _w8017_ ;
	wire _w8018_ ;
	wire _w8019_ ;
	wire _w8020_ ;
	wire _w8021_ ;
	wire _w8022_ ;
	wire _w8023_ ;
	wire _w8024_ ;
	wire _w8025_ ;
	wire _w8026_ ;
	wire _w8027_ ;
	wire _w8028_ ;
	wire _w8029_ ;
	wire _w8030_ ;
	wire _w8031_ ;
	wire _w8032_ ;
	wire _w8033_ ;
	wire _w8034_ ;
	wire _w8035_ ;
	wire _w8036_ ;
	wire _w8037_ ;
	wire _w8038_ ;
	wire _w8039_ ;
	wire _w8040_ ;
	wire _w8041_ ;
	wire _w8042_ ;
	wire _w8043_ ;
	wire _w8044_ ;
	wire _w8045_ ;
	wire _w8046_ ;
	wire _w8047_ ;
	wire _w8048_ ;
	wire _w8049_ ;
	wire _w8050_ ;
	wire _w8051_ ;
	wire _w8052_ ;
	wire _w8053_ ;
	wire _w8054_ ;
	wire _w8055_ ;
	wire _w8056_ ;
	wire _w8057_ ;
	wire _w8058_ ;
	wire _w8059_ ;
	wire _w8060_ ;
	wire _w8061_ ;
	wire _w8062_ ;
	wire _w8063_ ;
	wire _w8064_ ;
	wire _w8065_ ;
	wire _w8066_ ;
	wire _w8067_ ;
	wire _w8068_ ;
	wire _w8069_ ;
	wire _w8070_ ;
	wire _w8071_ ;
	wire _w8072_ ;
	wire _w8073_ ;
	wire _w8074_ ;
	wire _w8075_ ;
	wire _w8076_ ;
	wire _w8077_ ;
	wire _w8078_ ;
	wire _w8079_ ;
	wire _w8080_ ;
	wire _w8081_ ;
	wire _w8082_ ;
	wire _w8083_ ;
	wire _w8084_ ;
	wire _w8085_ ;
	wire _w8086_ ;
	wire _w8087_ ;
	wire _w8088_ ;
	wire _w8089_ ;
	wire _w8090_ ;
	wire _w8091_ ;
	wire _w8092_ ;
	wire _w8093_ ;
	wire _w8094_ ;
	wire _w8095_ ;
	wire _w8096_ ;
	wire _w8097_ ;
	wire _w8098_ ;
	wire _w8099_ ;
	wire _w8100_ ;
	wire _w8101_ ;
	wire _w8102_ ;
	wire _w8103_ ;
	wire _w8104_ ;
	wire _w8105_ ;
	wire _w8106_ ;
	wire _w8107_ ;
	wire _w8108_ ;
	wire _w8109_ ;
	wire _w8110_ ;
	wire _w8111_ ;
	wire _w8112_ ;
	wire _w8113_ ;
	wire _w8114_ ;
	wire _w8115_ ;
	wire _w8116_ ;
	wire _w8117_ ;
	wire _w8118_ ;
	wire _w8119_ ;
	wire _w8120_ ;
	wire _w8121_ ;
	wire _w8122_ ;
	wire _w8123_ ;
	wire _w8124_ ;
	wire _w8125_ ;
	wire _w8126_ ;
	wire _w8127_ ;
	wire _w8128_ ;
	wire _w8129_ ;
	wire _w8130_ ;
	wire _w8131_ ;
	wire _w8132_ ;
	wire _w8133_ ;
	wire _w8134_ ;
	wire _w8135_ ;
	wire _w8136_ ;
	wire _w8137_ ;
	wire _w8138_ ;
	wire _w8139_ ;
	wire _w8140_ ;
	wire _w8141_ ;
	wire _w8142_ ;
	wire _w8143_ ;
	wire _w8144_ ;
	wire _w8145_ ;
	wire _w8146_ ;
	wire _w8147_ ;
	wire _w8148_ ;
	wire _w8149_ ;
	wire _w8150_ ;
	wire _w8151_ ;
	wire _w8152_ ;
	wire _w8153_ ;
	wire _w8154_ ;
	wire _w8155_ ;
	wire _w8156_ ;
	wire _w8157_ ;
	wire _w8158_ ;
	wire _w8159_ ;
	wire _w8160_ ;
	wire _w8161_ ;
	wire _w8162_ ;
	wire _w8163_ ;
	wire _w8164_ ;
	wire _w8165_ ;
	wire _w8166_ ;
	wire _w8167_ ;
	wire _w8168_ ;
	wire _w8169_ ;
	wire _w8170_ ;
	wire _w8171_ ;
	wire _w8172_ ;
	wire _w8173_ ;
	wire _w8174_ ;
	wire _w8175_ ;
	wire _w8176_ ;
	wire _w8177_ ;
	wire _w8178_ ;
	wire _w8179_ ;
	wire _w8180_ ;
	wire _w8181_ ;
	wire _w8182_ ;
	wire _w8183_ ;
	wire _w8184_ ;
	wire _w8185_ ;
	wire _w8186_ ;
	wire _w8187_ ;
	wire _w8188_ ;
	wire _w8189_ ;
	wire _w8190_ ;
	wire _w8191_ ;
	wire _w8192_ ;
	wire _w8193_ ;
	wire _w8194_ ;
	wire _w8195_ ;
	wire _w8196_ ;
	wire _w8197_ ;
	wire _w8198_ ;
	wire _w8199_ ;
	wire _w8200_ ;
	wire _w8201_ ;
	wire _w8202_ ;
	wire _w8203_ ;
	wire _w8204_ ;
	wire _w8205_ ;
	wire _w8206_ ;
	wire _w8207_ ;
	wire _w8208_ ;
	wire _w8209_ ;
	wire _w8210_ ;
	wire _w8211_ ;
	wire _w8212_ ;
	wire _w8213_ ;
	wire _w8214_ ;
	wire _w8215_ ;
	wire _w8216_ ;
	wire _w8217_ ;
	wire _w8218_ ;
	wire _w8219_ ;
	wire _w8220_ ;
	wire _w8221_ ;
	wire _w8222_ ;
	wire _w8223_ ;
	wire _w8224_ ;
	wire _w8225_ ;
	wire _w8226_ ;
	wire _w8227_ ;
	wire _w8228_ ;
	wire _w8229_ ;
	wire _w8230_ ;
	wire _w8231_ ;
	wire _w8232_ ;
	wire _w8233_ ;
	wire _w8234_ ;
	wire _w8235_ ;
	wire _w8236_ ;
	wire _w8237_ ;
	wire _w8238_ ;
	wire _w8239_ ;
	wire _w8240_ ;
	wire _w8241_ ;
	wire _w8242_ ;
	wire _w8243_ ;
	wire _w8244_ ;
	wire _w8245_ ;
	wire _w8246_ ;
	wire _w8247_ ;
	wire _w8248_ ;
	wire _w8249_ ;
	wire _w8250_ ;
	wire _w8251_ ;
	wire _w8252_ ;
	wire _w8253_ ;
	wire _w8254_ ;
	wire _w8255_ ;
	wire _w8256_ ;
	wire _w8257_ ;
	wire _w8258_ ;
	wire _w8259_ ;
	wire _w8260_ ;
	wire _w8261_ ;
	wire _w8262_ ;
	wire _w8263_ ;
	wire _w8264_ ;
	wire _w8265_ ;
	wire _w8266_ ;
	wire _w8267_ ;
	wire _w8268_ ;
	wire _w8269_ ;
	wire _w8270_ ;
	wire _w8271_ ;
	wire _w8272_ ;
	wire _w8273_ ;
	wire _w8274_ ;
	wire _w8275_ ;
	wire _w8276_ ;
	wire _w8277_ ;
	wire _w8278_ ;
	wire _w8279_ ;
	wire _w8280_ ;
	wire _w8281_ ;
	wire _w8282_ ;
	wire _w8283_ ;
	wire _w8284_ ;
	wire _w8285_ ;
	wire _w8286_ ;
	wire _w8287_ ;
	wire _w8288_ ;
	wire _w8289_ ;
	wire _w8290_ ;
	wire _w8291_ ;
	wire _w8292_ ;
	wire _w8293_ ;
	wire _w8294_ ;
	wire _w8295_ ;
	wire _w8296_ ;
	wire _w8297_ ;
	wire _w8298_ ;
	wire _w8299_ ;
	wire _w8300_ ;
	wire _w8301_ ;
	wire _w8302_ ;
	wire _w8303_ ;
	wire _w8304_ ;
	wire _w8305_ ;
	wire _w8306_ ;
	wire _w8307_ ;
	wire _w8308_ ;
	wire _w8309_ ;
	wire _w8310_ ;
	wire _w8311_ ;
	wire _w8312_ ;
	wire _w8313_ ;
	wire _w8314_ ;
	wire _w8315_ ;
	wire _w8316_ ;
	wire _w8317_ ;
	wire _w8318_ ;
	wire _w8319_ ;
	wire _w8320_ ;
	wire _w8321_ ;
	wire _w8322_ ;
	wire _w8323_ ;
	wire _w8324_ ;
	wire _w8325_ ;
	wire _w8326_ ;
	wire _w8327_ ;
	wire _w8328_ ;
	wire _w8329_ ;
	wire _w8330_ ;
	wire _w8331_ ;
	wire _w8332_ ;
	wire _w8333_ ;
	wire _w8334_ ;
	wire _w8335_ ;
	wire _w8336_ ;
	wire _w8337_ ;
	wire _w8338_ ;
	wire _w8339_ ;
	wire _w8340_ ;
	wire _w8341_ ;
	wire _w8342_ ;
	wire _w8343_ ;
	wire _w8344_ ;
	wire _w8345_ ;
	wire _w8346_ ;
	wire _w8347_ ;
	wire _w8348_ ;
	wire _w8349_ ;
	wire _w8350_ ;
	wire _w8351_ ;
	wire _w8352_ ;
	wire _w8353_ ;
	wire _w8354_ ;
	wire _w8355_ ;
	wire _w8356_ ;
	wire _w8357_ ;
	wire _w8358_ ;
	wire _w8359_ ;
	wire _w8360_ ;
	wire _w8361_ ;
	wire _w8362_ ;
	wire _w8363_ ;
	wire _w8364_ ;
	wire _w8365_ ;
	wire _w8366_ ;
	wire _w8367_ ;
	wire _w8368_ ;
	wire _w8369_ ;
	wire _w8370_ ;
	wire _w8371_ ;
	wire _w8372_ ;
	wire _w8373_ ;
	wire _w8374_ ;
	wire _w8375_ ;
	wire _w8376_ ;
	wire _w8377_ ;
	wire _w8378_ ;
	wire _w8379_ ;
	wire _w8380_ ;
	wire _w8381_ ;
	wire _w8382_ ;
	wire _w8383_ ;
	wire _w8384_ ;
	wire _w8385_ ;
	wire _w8386_ ;
	wire _w8387_ ;
	wire _w8388_ ;
	wire _w8389_ ;
	wire _w8390_ ;
	wire _w8391_ ;
	wire _w8392_ ;
	wire _w8393_ ;
	wire _w8394_ ;
	wire _w8395_ ;
	wire _w8396_ ;
	wire _w8397_ ;
	wire _w8398_ ;
	wire _w8399_ ;
	wire _w8400_ ;
	wire _w8401_ ;
	wire _w8402_ ;
	wire _w8403_ ;
	wire _w8404_ ;
	wire _w8405_ ;
	wire _w8406_ ;
	wire _w8407_ ;
	wire _w8408_ ;
	wire _w8409_ ;
	wire _w8410_ ;
	wire _w8411_ ;
	wire _w8412_ ;
	wire _w8413_ ;
	wire _w8414_ ;
	wire _w8415_ ;
	wire _w8416_ ;
	wire _w8417_ ;
	wire _w8418_ ;
	wire _w8419_ ;
	wire _w8420_ ;
	wire _w8421_ ;
	wire _w8422_ ;
	wire _w8423_ ;
	wire _w8424_ ;
	wire _w8425_ ;
	wire _w8426_ ;
	wire _w8427_ ;
	wire _w8428_ ;
	wire _w8429_ ;
	wire _w8430_ ;
	wire _w8431_ ;
	wire _w8432_ ;
	wire _w8433_ ;
	wire _w8434_ ;
	wire _w8435_ ;
	wire _w8436_ ;
	wire _w8437_ ;
	wire _w8438_ ;
	wire _w8439_ ;
	wire _w8440_ ;
	wire _w8441_ ;
	wire _w8442_ ;
	wire _w8443_ ;
	wire _w8444_ ;
	wire _w8445_ ;
	wire _w8446_ ;
	wire _w8447_ ;
	wire _w8448_ ;
	wire _w8449_ ;
	wire _w8450_ ;
	wire _w8451_ ;
	wire _w8452_ ;
	wire _w8453_ ;
	wire _w8454_ ;
	wire _w8455_ ;
	wire _w8456_ ;
	wire _w8457_ ;
	wire _w8458_ ;
	wire _w8459_ ;
	wire _w8460_ ;
	wire _w8461_ ;
	wire _w8462_ ;
	wire _w8463_ ;
	wire _w8464_ ;
	wire _w8465_ ;
	wire _w8466_ ;
	wire _w8467_ ;
	wire _w8468_ ;
	wire _w8469_ ;
	wire _w8470_ ;
	wire _w8471_ ;
	wire _w8472_ ;
	wire _w8473_ ;
	wire _w8474_ ;
	wire _w8475_ ;
	wire _w8476_ ;
	wire _w8477_ ;
	wire _w8478_ ;
	wire _w8479_ ;
	wire _w8480_ ;
	wire _w8481_ ;
	wire _w8482_ ;
	wire _w8483_ ;
	wire _w8484_ ;
	wire _w8485_ ;
	wire _w8486_ ;
	wire _w8487_ ;
	wire _w8488_ ;
	wire _w8489_ ;
	wire _w8490_ ;
	wire _w8491_ ;
	wire _w8492_ ;
	wire _w8493_ ;
	wire _w8494_ ;
	wire _w8495_ ;
	wire _w8496_ ;
	wire _w8497_ ;
	wire _w8498_ ;
	wire _w8499_ ;
	wire _w8500_ ;
	wire _w8501_ ;
	wire _w8502_ ;
	wire _w8503_ ;
	wire _w8504_ ;
	wire _w8505_ ;
	wire _w8506_ ;
	wire _w8507_ ;
	wire _w8508_ ;
	wire _w8509_ ;
	wire _w8510_ ;
	wire _w8511_ ;
	wire _w8512_ ;
	wire _w8513_ ;
	wire _w8514_ ;
	wire _w8515_ ;
	wire _w8516_ ;
	wire _w8517_ ;
	wire _w8518_ ;
	wire _w8519_ ;
	wire _w8520_ ;
	wire _w8521_ ;
	wire _w8522_ ;
	wire _w8523_ ;
	wire _w8524_ ;
	wire _w8525_ ;
	wire _w8526_ ;
	wire _w8527_ ;
	wire _w8528_ ;
	wire _w8529_ ;
	wire _w8530_ ;
	wire _w8531_ ;
	wire _w8532_ ;
	wire _w8533_ ;
	wire _w8534_ ;
	wire _w8535_ ;
	wire _w8536_ ;
	wire _w8537_ ;
	wire _w8538_ ;
	wire _w8539_ ;
	wire _w8540_ ;
	wire _w8541_ ;
	wire _w8542_ ;
	wire _w8543_ ;
	wire _w8544_ ;
	wire _w8545_ ;
	wire _w8546_ ;
	wire _w8547_ ;
	wire _w8548_ ;
	wire _w8549_ ;
	wire _w8550_ ;
	wire _w8551_ ;
	wire _w8552_ ;
	wire _w8553_ ;
	wire _w8554_ ;
	wire _w8555_ ;
	wire _w8556_ ;
	wire _w8557_ ;
	wire _w8558_ ;
	wire _w8559_ ;
	wire _w8560_ ;
	wire _w8561_ ;
	wire _w8562_ ;
	wire _w8563_ ;
	wire _w8564_ ;
	wire _w8565_ ;
	wire _w8566_ ;
	wire _w8567_ ;
	wire _w8568_ ;
	wire _w8569_ ;
	wire _w8570_ ;
	wire _w8571_ ;
	wire _w8572_ ;
	wire _w8573_ ;
	wire _w8574_ ;
	wire _w8575_ ;
	wire _w8576_ ;
	wire _w8577_ ;
	wire _w8578_ ;
	wire _w8579_ ;
	wire _w8580_ ;
	wire _w8581_ ;
	wire _w8582_ ;
	wire _w8583_ ;
	wire _w8584_ ;
	wire _w8585_ ;
	wire _w8586_ ;
	wire _w8587_ ;
	wire _w8588_ ;
	wire _w8589_ ;
	wire _w8590_ ;
	wire _w8591_ ;
	wire _w8592_ ;
	wire _w8593_ ;
	wire _w8594_ ;
	wire _w8595_ ;
	wire _w8596_ ;
	wire _w8597_ ;
	wire _w8598_ ;
	wire _w8599_ ;
	wire _w8600_ ;
	wire _w8601_ ;
	wire _w8602_ ;
	wire _w8603_ ;
	wire _w8604_ ;
	wire _w8605_ ;
	wire _w8606_ ;
	wire _w8607_ ;
	wire _w8608_ ;
	wire _w8609_ ;
	wire _w8610_ ;
	wire _w8611_ ;
	wire _w8612_ ;
	wire _w8613_ ;
	wire _w8614_ ;
	wire _w8615_ ;
	wire _w8616_ ;
	wire _w8617_ ;
	wire _w8618_ ;
	wire _w8619_ ;
	wire _w8620_ ;
	wire _w8621_ ;
	wire _w8622_ ;
	wire _w8623_ ;
	wire _w8624_ ;
	wire _w8625_ ;
	wire _w8626_ ;
	wire _w8627_ ;
	wire _w8628_ ;
	wire _w8629_ ;
	wire _w8630_ ;
	wire _w8631_ ;
	wire _w8632_ ;
	wire _w8633_ ;
	wire _w8634_ ;
	wire _w8635_ ;
	wire _w8636_ ;
	wire _w8637_ ;
	wire _w8638_ ;
	wire _w8639_ ;
	wire _w8640_ ;
	wire _w8641_ ;
	wire _w8642_ ;
	wire _w8643_ ;
	wire _w8644_ ;
	wire _w8645_ ;
	wire _w8646_ ;
	wire _w8647_ ;
	wire _w8648_ ;
	wire _w8649_ ;
	wire _w8650_ ;
	wire _w8651_ ;
	wire _w8652_ ;
	wire _w8653_ ;
	wire _w8654_ ;
	wire _w8655_ ;
	wire _w8656_ ;
	wire _w8657_ ;
	wire _w8658_ ;
	wire _w8659_ ;
	wire _w8660_ ;
	wire _w8661_ ;
	wire _w8662_ ;
	wire _w8663_ ;
	wire _w8664_ ;
	wire _w8665_ ;
	wire _w8666_ ;
	wire _w8667_ ;
	wire _w8668_ ;
	wire _w8669_ ;
	wire _w8670_ ;
	wire _w8671_ ;
	wire _w8672_ ;
	wire _w8673_ ;
	wire _w8674_ ;
	wire _w8675_ ;
	wire _w8676_ ;
	wire _w8677_ ;
	wire _w8678_ ;
	wire _w8679_ ;
	wire _w8680_ ;
	wire _w8681_ ;
	wire _w8682_ ;
	wire _w8683_ ;
	wire _w8684_ ;
	wire _w8685_ ;
	wire _w8686_ ;
	wire _w8687_ ;
	wire _w8688_ ;
	wire _w8689_ ;
	wire _w8690_ ;
	wire _w8691_ ;
	wire _w8692_ ;
	wire _w8693_ ;
	wire _w8694_ ;
	wire _w8695_ ;
	wire _w8696_ ;
	wire _w8697_ ;
	wire _w8698_ ;
	wire _w8699_ ;
	wire _w8700_ ;
	wire _w8701_ ;
	wire _w8702_ ;
	wire _w8703_ ;
	wire _w8704_ ;
	wire _w8705_ ;
	wire _w8706_ ;
	wire _w8707_ ;
	wire _w8708_ ;
	wire _w8709_ ;
	wire _w8710_ ;
	wire _w8711_ ;
	wire _w8712_ ;
	wire _w8713_ ;
	wire _w8714_ ;
	wire _w8715_ ;
	wire _w8716_ ;
	wire _w8717_ ;
	wire _w8718_ ;
	wire _w8719_ ;
	wire _w8720_ ;
	wire _w8721_ ;
	wire _w8722_ ;
	wire _w8723_ ;
	wire _w8724_ ;
	wire _w8725_ ;
	wire _w8726_ ;
	wire _w8727_ ;
	wire _w8728_ ;
	wire _w8729_ ;
	wire _w8730_ ;
	wire _w8731_ ;
	wire _w8732_ ;
	wire _w8733_ ;
	wire _w8734_ ;
	wire _w8735_ ;
	wire _w8736_ ;
	wire _w8737_ ;
	wire _w8738_ ;
	wire _w8739_ ;
	wire _w8740_ ;
	wire _w8741_ ;
	wire _w8742_ ;
	wire _w8743_ ;
	wire _w8744_ ;
	wire _w8745_ ;
	wire _w8746_ ;
	wire _w8747_ ;
	wire _w8748_ ;
	wire _w8749_ ;
	wire _w8750_ ;
	wire _w8751_ ;
	wire _w8752_ ;
	wire _w8753_ ;
	wire _w8754_ ;
	wire _w8755_ ;
	wire _w8756_ ;
	wire _w8757_ ;
	wire _w8758_ ;
	wire _w8759_ ;
	wire _w8760_ ;
	wire _w8761_ ;
	wire _w8762_ ;
	wire _w8763_ ;
	wire _w8764_ ;
	wire _w8765_ ;
	wire _w8766_ ;
	wire _w8767_ ;
	wire _w8768_ ;
	wire _w8769_ ;
	wire _w8770_ ;
	wire _w8771_ ;
	wire _w8772_ ;
	wire _w8773_ ;
	wire _w8774_ ;
	wire _w8775_ ;
	wire _w8776_ ;
	wire _w8777_ ;
	wire _w8778_ ;
	wire _w8779_ ;
	wire _w8780_ ;
	wire _w8781_ ;
	wire _w8782_ ;
	wire _w8783_ ;
	wire _w8784_ ;
	wire _w8785_ ;
	wire _w8786_ ;
	wire _w8787_ ;
	wire _w8788_ ;
	wire _w8789_ ;
	wire _w8790_ ;
	wire _w8791_ ;
	wire _w8792_ ;
	wire _w8793_ ;
	wire _w8794_ ;
	wire _w8795_ ;
	wire _w8796_ ;
	wire _w8797_ ;
	wire _w8798_ ;
	wire _w8799_ ;
	wire _w8800_ ;
	wire _w8801_ ;
	wire _w8802_ ;
	wire _w8803_ ;
	wire _w8804_ ;
	wire _w8805_ ;
	wire _w8806_ ;
	wire _w8807_ ;
	wire _w8808_ ;
	wire _w8809_ ;
	wire _w8810_ ;
	wire _w8811_ ;
	wire _w8812_ ;
	wire _w8813_ ;
	wire _w8814_ ;
	wire _w8815_ ;
	wire _w8816_ ;
	wire _w8817_ ;
	wire _w8818_ ;
	wire _w8819_ ;
	wire _w8820_ ;
	wire _w8821_ ;
	wire _w8822_ ;
	wire _w8823_ ;
	wire _w8824_ ;
	wire _w8825_ ;
	wire _w8826_ ;
	wire _w8827_ ;
	wire _w8828_ ;
	wire _w8829_ ;
	wire _w8830_ ;
	wire _w8831_ ;
	wire _w8832_ ;
	wire _w8833_ ;
	wire _w8834_ ;
	wire _w8835_ ;
	wire _w8836_ ;
	wire _w8837_ ;
	wire _w8838_ ;
	wire _w8839_ ;
	wire _w8840_ ;
	wire _w8841_ ;
	wire _w8842_ ;
	wire _w8843_ ;
	wire _w8844_ ;
	wire _w8845_ ;
	wire _w8846_ ;
	wire _w8847_ ;
	wire _w8848_ ;
	wire _w8849_ ;
	wire _w8850_ ;
	wire _w8851_ ;
	wire _w8852_ ;
	wire _w8853_ ;
	wire _w8854_ ;
	wire _w8855_ ;
	wire _w8856_ ;
	wire _w8857_ ;
	wire _w8858_ ;
	wire _w8859_ ;
	wire _w8860_ ;
	wire _w8861_ ;
	wire _w8862_ ;
	wire _w8863_ ;
	wire _w8864_ ;
	wire _w8865_ ;
	wire _w8866_ ;
	wire _w8867_ ;
	wire _w8868_ ;
	wire _w8869_ ;
	wire _w8870_ ;
	wire _w8871_ ;
	wire _w8872_ ;
	wire _w8873_ ;
	wire _w8874_ ;
	wire _w8875_ ;
	wire _w8876_ ;
	wire _w8877_ ;
	wire _w8878_ ;
	wire _w8879_ ;
	wire _w8880_ ;
	wire _w8881_ ;
	wire _w8882_ ;
	wire _w8883_ ;
	wire _w8884_ ;
	wire _w8885_ ;
	wire _w8886_ ;
	wire _w8887_ ;
	wire _w8888_ ;
	wire _w8889_ ;
	wire _w8890_ ;
	wire _w8891_ ;
	wire _w8892_ ;
	wire _w8893_ ;
	wire _w8894_ ;
	wire _w8895_ ;
	wire _w8896_ ;
	wire _w8897_ ;
	wire _w8898_ ;
	wire _w8899_ ;
	wire _w8900_ ;
	wire _w8901_ ;
	wire _w8902_ ;
	wire _w8903_ ;
	wire _w8904_ ;
	wire _w8905_ ;
	wire _w8906_ ;
	wire _w8907_ ;
	wire _w8908_ ;
	wire _w8909_ ;
	wire _w8910_ ;
	wire _w8911_ ;
	wire _w8912_ ;
	wire _w8913_ ;
	wire _w8914_ ;
	wire _w8915_ ;
	wire _w8916_ ;
	wire _w8917_ ;
	wire _w8918_ ;
	wire _w8919_ ;
	wire _w8920_ ;
	wire _w8921_ ;
	wire _w8922_ ;
	wire _w8923_ ;
	wire _w8924_ ;
	wire _w8925_ ;
	wire _w8926_ ;
	wire _w8927_ ;
	wire _w8928_ ;
	wire _w8929_ ;
	wire _w8930_ ;
	wire _w8931_ ;
	wire _w8932_ ;
	wire _w8933_ ;
	wire _w8934_ ;
	wire _w8935_ ;
	wire _w8936_ ;
	wire _w8937_ ;
	wire _w8938_ ;
	wire _w8939_ ;
	wire _w8940_ ;
	wire _w8941_ ;
	wire _w8942_ ;
	wire _w8943_ ;
	wire _w8944_ ;
	wire _w8945_ ;
	wire _w8946_ ;
	wire _w8947_ ;
	wire _w8948_ ;
	wire _w8949_ ;
	wire _w8950_ ;
	wire _w8951_ ;
	wire _w8952_ ;
	wire _w8953_ ;
	wire _w8954_ ;
	wire _w8955_ ;
	wire _w8956_ ;
	wire _w8957_ ;
	wire _w8958_ ;
	wire _w8959_ ;
	wire _w8960_ ;
	wire _w8961_ ;
	wire _w8962_ ;
	wire _w8963_ ;
	wire _w8964_ ;
	wire _w8965_ ;
	wire _w8966_ ;
	wire _w8967_ ;
	wire _w8968_ ;
	wire _w8969_ ;
	wire _w8970_ ;
	wire _w8971_ ;
	wire _w8972_ ;
	wire _w8973_ ;
	wire _w8974_ ;
	wire _w8975_ ;
	wire _w8976_ ;
	wire _w8977_ ;
	wire _w8978_ ;
	wire _w8979_ ;
	wire _w8980_ ;
	wire _w8981_ ;
	wire _w8982_ ;
	wire _w8983_ ;
	wire _w8984_ ;
	wire _w8985_ ;
	wire _w8986_ ;
	wire _w8987_ ;
	wire _w8988_ ;
	wire _w8989_ ;
	wire _w8990_ ;
	wire _w8991_ ;
	wire _w8992_ ;
	wire _w8993_ ;
	wire _w8994_ ;
	wire _w8995_ ;
	wire _w8996_ ;
	wire _w8997_ ;
	wire _w8998_ ;
	wire _w8999_ ;
	wire _w9000_ ;
	wire _w9001_ ;
	wire _w9002_ ;
	wire _w9003_ ;
	wire _w9004_ ;
	wire _w9005_ ;
	wire _w9006_ ;
	wire _w9007_ ;
	wire _w9008_ ;
	wire _w9009_ ;
	wire _w9010_ ;
	wire _w9011_ ;
	wire _w9012_ ;
	wire _w9013_ ;
	wire _w9014_ ;
	wire _w9015_ ;
	wire _w9016_ ;
	wire _w9017_ ;
	wire _w9018_ ;
	wire _w9019_ ;
	wire _w9020_ ;
	wire _w9021_ ;
	wire _w9022_ ;
	wire _w9023_ ;
	wire _w9024_ ;
	wire _w9025_ ;
	wire _w9026_ ;
	wire _w9027_ ;
	wire _w9028_ ;
	wire _w9029_ ;
	wire _w9030_ ;
	wire _w9031_ ;
	wire _w9032_ ;
	wire _w9033_ ;
	wire _w9034_ ;
	wire _w9035_ ;
	wire _w9036_ ;
	wire _w9037_ ;
	wire _w9038_ ;
	wire _w9039_ ;
	wire _w9040_ ;
	wire _w9041_ ;
	wire _w9042_ ;
	wire _w9043_ ;
	wire _w9044_ ;
	wire _w9045_ ;
	wire _w9046_ ;
	wire _w9047_ ;
	wire _w9048_ ;
	wire _w9049_ ;
	wire _w9050_ ;
	wire _w9051_ ;
	wire _w9052_ ;
	wire _w9053_ ;
	wire _w9054_ ;
	wire _w9055_ ;
	wire _w9056_ ;
	wire _w9057_ ;
	wire _w9058_ ;
	wire _w9059_ ;
	wire _w9060_ ;
	wire _w9061_ ;
	wire _w9062_ ;
	wire _w9063_ ;
	wire _w9064_ ;
	wire _w9065_ ;
	wire _w9066_ ;
	wire _w9067_ ;
	wire _w9068_ ;
	wire _w9069_ ;
	wire _w9070_ ;
	wire _w9071_ ;
	wire _w9072_ ;
	wire _w9073_ ;
	wire _w9074_ ;
	wire _w9075_ ;
	wire _w9076_ ;
	wire _w9077_ ;
	wire _w9078_ ;
	wire _w9079_ ;
	wire _w9080_ ;
	wire _w9081_ ;
	wire _w9082_ ;
	wire _w9083_ ;
	wire _w9084_ ;
	wire _w9085_ ;
	wire _w9086_ ;
	wire _w9087_ ;
	wire _w9088_ ;
	wire _w9089_ ;
	wire _w9090_ ;
	wire _w9091_ ;
	wire _w9092_ ;
	wire _w9093_ ;
	wire _w9094_ ;
	wire _w9095_ ;
	wire _w9096_ ;
	wire _w9097_ ;
	wire _w9098_ ;
	wire _w9099_ ;
	wire _w9100_ ;
	wire _w9101_ ;
	wire _w9102_ ;
	wire _w9103_ ;
	wire _w9104_ ;
	wire _w9105_ ;
	wire _w9106_ ;
	wire _w9107_ ;
	wire _w9108_ ;
	wire _w9109_ ;
	wire _w9110_ ;
	wire _w9111_ ;
	wire _w9112_ ;
	wire _w9113_ ;
	wire _w9114_ ;
	wire _w9115_ ;
	wire _w9116_ ;
	wire _w9117_ ;
	wire _w9118_ ;
	wire _w9119_ ;
	wire _w9120_ ;
	wire _w9121_ ;
	wire _w9122_ ;
	wire _w9123_ ;
	wire _w9124_ ;
	wire _w9125_ ;
	wire _w9126_ ;
	wire _w9127_ ;
	wire _w9128_ ;
	wire _w9129_ ;
	wire _w9130_ ;
	wire _w9131_ ;
	wire _w9132_ ;
	wire _w9133_ ;
	wire _w9134_ ;
	wire _w9135_ ;
	wire _w9136_ ;
	wire _w9137_ ;
	wire _w9138_ ;
	wire _w9139_ ;
	wire _w9140_ ;
	wire _w9141_ ;
	wire _w9142_ ;
	wire _w9143_ ;
	wire _w9144_ ;
	wire _w9145_ ;
	wire _w9146_ ;
	wire _w9147_ ;
	wire _w9148_ ;
	wire _w9149_ ;
	wire _w9150_ ;
	wire _w9151_ ;
	wire _w9152_ ;
	wire _w9153_ ;
	wire _w9154_ ;
	wire _w9155_ ;
	wire _w9156_ ;
	wire _w9157_ ;
	wire _w9158_ ;
	wire _w9159_ ;
	wire _w9160_ ;
	wire _w9161_ ;
	wire _w9162_ ;
	wire _w9163_ ;
	wire _w9164_ ;
	wire _w9165_ ;
	wire _w9166_ ;
	wire _w9167_ ;
	wire _w9168_ ;
	wire _w9169_ ;
	wire _w9170_ ;
	wire _w9171_ ;
	wire _w9172_ ;
	wire _w9173_ ;
	wire _w9174_ ;
	wire _w9175_ ;
	wire _w9176_ ;
	wire _w9177_ ;
	wire _w9178_ ;
	wire _w9179_ ;
	wire _w9180_ ;
	wire _w9181_ ;
	wire _w9182_ ;
	wire _w9183_ ;
	wire _w9184_ ;
	wire _w9185_ ;
	wire _w9186_ ;
	wire _w9187_ ;
	wire _w9188_ ;
	wire _w9189_ ;
	wire _w9190_ ;
	wire _w9191_ ;
	wire _w9192_ ;
	wire _w9193_ ;
	wire _w9194_ ;
	wire _w9195_ ;
	wire _w9196_ ;
	wire _w9197_ ;
	wire _w9198_ ;
	wire _w9199_ ;
	wire _w9200_ ;
	wire _w9201_ ;
	wire _w9202_ ;
	wire _w9203_ ;
	wire _w9204_ ;
	wire _w9205_ ;
	wire _w9206_ ;
	wire _w9207_ ;
	wire _w9208_ ;
	wire _w9209_ ;
	wire _w9210_ ;
	wire _w9211_ ;
	wire _w9212_ ;
	wire _w9213_ ;
	wire _w9214_ ;
	wire _w9215_ ;
	wire _w9216_ ;
	wire _w9217_ ;
	wire _w9218_ ;
	wire _w9219_ ;
	wire _w9220_ ;
	wire _w9221_ ;
	wire _w9222_ ;
	wire _w9223_ ;
	wire _w9224_ ;
	wire _w9225_ ;
	wire _w9226_ ;
	wire _w9227_ ;
	wire _w9228_ ;
	wire _w9229_ ;
	wire _w9230_ ;
	wire _w9231_ ;
	wire _w9232_ ;
	wire _w9233_ ;
	wire _w9234_ ;
	wire _w9235_ ;
	wire _w9236_ ;
	wire _w9237_ ;
	wire _w9238_ ;
	wire _w9239_ ;
	wire _w9240_ ;
	wire _w9241_ ;
	wire _w9242_ ;
	wire _w9243_ ;
	wire _w9244_ ;
	wire _w9245_ ;
	wire _w9246_ ;
	wire _w9247_ ;
	wire _w9248_ ;
	wire _w9249_ ;
	wire _w9250_ ;
	wire _w9251_ ;
	wire _w9252_ ;
	wire _w9253_ ;
	wire _w9254_ ;
	wire _w9255_ ;
	wire _w9256_ ;
	wire _w9257_ ;
	wire _w9258_ ;
	wire _w9259_ ;
	wire _w9260_ ;
	wire _w9261_ ;
	wire _w9262_ ;
	wire _w9263_ ;
	wire _w9264_ ;
	wire _w9265_ ;
	wire _w9266_ ;
	wire _w9267_ ;
	wire _w9268_ ;
	wire _w9269_ ;
	wire _w9270_ ;
	wire _w9271_ ;
	wire _w9272_ ;
	wire _w9273_ ;
	wire _w9274_ ;
	wire _w9275_ ;
	wire _w9276_ ;
	wire _w9277_ ;
	wire _w9278_ ;
	wire _w9279_ ;
	wire _w9280_ ;
	wire _w9281_ ;
	wire _w9282_ ;
	wire _w9283_ ;
	wire _w9284_ ;
	wire _w9285_ ;
	wire _w9286_ ;
	wire _w9287_ ;
	wire _w9288_ ;
	wire _w9289_ ;
	wire _w9290_ ;
	wire _w9291_ ;
	wire _w9292_ ;
	wire _w9293_ ;
	wire _w9294_ ;
	wire _w9295_ ;
	wire _w9296_ ;
	wire _w9297_ ;
	wire _w9298_ ;
	wire _w9299_ ;
	wire _w9300_ ;
	wire _w9301_ ;
	wire _w9302_ ;
	wire _w9303_ ;
	wire _w9304_ ;
	wire _w9305_ ;
	wire _w9306_ ;
	wire _w9307_ ;
	wire _w9308_ ;
	wire _w9309_ ;
	wire _w9310_ ;
	wire _w9311_ ;
	wire _w9312_ ;
	wire _w9313_ ;
	wire _w9314_ ;
	wire _w9315_ ;
	wire _w9316_ ;
	wire _w9317_ ;
	wire _w9318_ ;
	wire _w9319_ ;
	wire _w9320_ ;
	wire _w9321_ ;
	wire _w9322_ ;
	wire _w9323_ ;
	wire _w9324_ ;
	wire _w9325_ ;
	wire _w9326_ ;
	wire _w9327_ ;
	wire _w9328_ ;
	wire _w9329_ ;
	wire _w9330_ ;
	wire _w9331_ ;
	wire _w9332_ ;
	wire _w9333_ ;
	wire _w9334_ ;
	wire _w9335_ ;
	wire _w9336_ ;
	wire _w9337_ ;
	wire _w9338_ ;
	wire _w9339_ ;
	wire _w9340_ ;
	wire _w9341_ ;
	wire _w9342_ ;
	wire _w9343_ ;
	wire _w9344_ ;
	wire _w9345_ ;
	wire _w9346_ ;
	wire _w9347_ ;
	wire _w9348_ ;
	wire _w9349_ ;
	wire _w9350_ ;
	wire _w9351_ ;
	wire _w9352_ ;
	wire _w9353_ ;
	wire _w9354_ ;
	wire _w9355_ ;
	wire _w9356_ ;
	wire _w9357_ ;
	wire _w9358_ ;
	wire _w9359_ ;
	wire _w9360_ ;
	wire _w9361_ ;
	wire _w9362_ ;
	wire _w9363_ ;
	wire _w9364_ ;
	wire _w9365_ ;
	wire _w9366_ ;
	wire _w9367_ ;
	wire _w9368_ ;
	wire _w9369_ ;
	wire _w9370_ ;
	wire _w9371_ ;
	wire _w9372_ ;
	wire _w9373_ ;
	wire _w9374_ ;
	wire _w9375_ ;
	wire _w9376_ ;
	wire _w9377_ ;
	wire _w9378_ ;
	wire _w9379_ ;
	wire _w9380_ ;
	wire _w9381_ ;
	wire _w9382_ ;
	wire _w9383_ ;
	wire _w9384_ ;
	wire _w9385_ ;
	wire _w9386_ ;
	wire _w9387_ ;
	wire _w9388_ ;
	wire _w9389_ ;
	wire _w9390_ ;
	wire _w9391_ ;
	wire _w9392_ ;
	wire _w9393_ ;
	wire _w9394_ ;
	wire _w9395_ ;
	wire _w9396_ ;
	wire _w9397_ ;
	wire _w9398_ ;
	wire _w9399_ ;
	wire _w9400_ ;
	wire _w9401_ ;
	wire _w9402_ ;
	wire _w9403_ ;
	wire _w9404_ ;
	wire _w9405_ ;
	wire _w9406_ ;
	wire _w9407_ ;
	wire _w9408_ ;
	wire _w9409_ ;
	wire _w9410_ ;
	wire _w9411_ ;
	wire _w9412_ ;
	wire _w9413_ ;
	wire _w9414_ ;
	wire _w9415_ ;
	wire _w9416_ ;
	wire _w9417_ ;
	wire _w9418_ ;
	wire _w9419_ ;
	wire _w9420_ ;
	wire _w9421_ ;
	wire _w9422_ ;
	wire _w9423_ ;
	wire _w9424_ ;
	wire _w9425_ ;
	wire _w9426_ ;
	wire _w9427_ ;
	wire _w9428_ ;
	wire _w9429_ ;
	wire _w9430_ ;
	wire _w9431_ ;
	wire _w9432_ ;
	wire _w9433_ ;
	wire _w9434_ ;
	wire _w9435_ ;
	wire _w9436_ ;
	wire _w9437_ ;
	wire _w9438_ ;
	wire _w9439_ ;
	wire _w9440_ ;
	wire _w9441_ ;
	wire _w9442_ ;
	wire _w9443_ ;
	wire _w9444_ ;
	wire _w9445_ ;
	wire _w9446_ ;
	wire _w9447_ ;
	wire _w9448_ ;
	wire _w9449_ ;
	wire _w9450_ ;
	wire _w9451_ ;
	wire _w9452_ ;
	wire _w9453_ ;
	wire _w9454_ ;
	wire _w9455_ ;
	wire _w9456_ ;
	wire _w9457_ ;
	wire _w9458_ ;
	wire _w9459_ ;
	wire _w9460_ ;
	wire _w9461_ ;
	wire _w9462_ ;
	wire _w9463_ ;
	wire _w9464_ ;
	wire _w9465_ ;
	wire _w9466_ ;
	wire _w9467_ ;
	wire _w9468_ ;
	wire _w9469_ ;
	wire _w9470_ ;
	wire _w9471_ ;
	wire _w9472_ ;
	wire _w9473_ ;
	wire _w9474_ ;
	wire _w9475_ ;
	wire _w9476_ ;
	wire _w9477_ ;
	wire _w9478_ ;
	wire _w9479_ ;
	wire _w9480_ ;
	wire _w9481_ ;
	wire _w9482_ ;
	wire _w9483_ ;
	wire _w9484_ ;
	wire _w9485_ ;
	wire _w9486_ ;
	wire _w9487_ ;
	wire _w9488_ ;
	wire _w9489_ ;
	wire _w9490_ ;
	wire _w9491_ ;
	wire _w9492_ ;
	wire _w9493_ ;
	wire _w9494_ ;
	wire _w9495_ ;
	wire _w9496_ ;
	wire _w9497_ ;
	wire _w9498_ ;
	wire _w9499_ ;
	wire _w9500_ ;
	wire _w9501_ ;
	wire _w9502_ ;
	wire _w9503_ ;
	wire _w9504_ ;
	wire _w9505_ ;
	wire _w9506_ ;
	wire _w9507_ ;
	wire _w9508_ ;
	wire _w9509_ ;
	wire _w9510_ ;
	wire _w9511_ ;
	wire _w9512_ ;
	wire _w9513_ ;
	wire _w9514_ ;
	wire _w9515_ ;
	wire _w9516_ ;
	wire _w9517_ ;
	wire _w9518_ ;
	wire _w9519_ ;
	wire _w9520_ ;
	wire _w9521_ ;
	wire _w9522_ ;
	wire _w9523_ ;
	wire _w9524_ ;
	wire _w9525_ ;
	wire _w9526_ ;
	wire _w9527_ ;
	wire _w9528_ ;
	wire _w9529_ ;
	wire _w9530_ ;
	wire _w9531_ ;
	wire _w9532_ ;
	wire _w9533_ ;
	wire _w9534_ ;
	wire _w9535_ ;
	wire _w9536_ ;
	wire _w9537_ ;
	wire _w9538_ ;
	wire _w9539_ ;
	wire _w9540_ ;
	wire _w9541_ ;
	wire _w9542_ ;
	wire _w9543_ ;
	wire _w9544_ ;
	wire _w9545_ ;
	wire _w9546_ ;
	wire _w9547_ ;
	wire _w9548_ ;
	wire _w9549_ ;
	wire _w9550_ ;
	wire _w9551_ ;
	wire _w9552_ ;
	wire _w9553_ ;
	wire _w9554_ ;
	wire _w9555_ ;
	wire _w9556_ ;
	wire _w9557_ ;
	wire _w9558_ ;
	wire _w9559_ ;
	wire _w9560_ ;
	wire _w9561_ ;
	wire _w9562_ ;
	wire _w9563_ ;
	wire _w9564_ ;
	wire _w9565_ ;
	wire _w9566_ ;
	wire _w9567_ ;
	wire _w9568_ ;
	wire _w9569_ ;
	wire _w9570_ ;
	wire _w9571_ ;
	wire _w9572_ ;
	wire _w9573_ ;
	wire _w9574_ ;
	wire _w9575_ ;
	wire _w9576_ ;
	wire _w9577_ ;
	wire _w9578_ ;
	wire _w9579_ ;
	wire _w9580_ ;
	wire _w9581_ ;
	wire _w9582_ ;
	wire _w9583_ ;
	wire _w9584_ ;
	wire _w9585_ ;
	wire _w9586_ ;
	wire _w9587_ ;
	wire _w9588_ ;
	wire _w9589_ ;
	wire _w9590_ ;
	wire _w9591_ ;
	wire _w9592_ ;
	wire _w9593_ ;
	wire _w9594_ ;
	wire _w9595_ ;
	wire _w9596_ ;
	wire _w9597_ ;
	wire _w9598_ ;
	wire _w9599_ ;
	wire _w9600_ ;
	wire _w9601_ ;
	wire _w9602_ ;
	wire _w9603_ ;
	wire _w9604_ ;
	wire _w9605_ ;
	wire _w9606_ ;
	wire _w9607_ ;
	wire _w9608_ ;
	wire _w9609_ ;
	wire _w9610_ ;
	wire _w9611_ ;
	wire _w9612_ ;
	wire _w9613_ ;
	wire _w9614_ ;
	wire _w9615_ ;
	wire _w9616_ ;
	wire _w9617_ ;
	wire _w9618_ ;
	wire _w9619_ ;
	wire _w9620_ ;
	wire _w9621_ ;
	wire _w9622_ ;
	wire _w9623_ ;
	wire _w9624_ ;
	wire _w9625_ ;
	wire _w9626_ ;
	wire _w9627_ ;
	wire _w9628_ ;
	wire _w9629_ ;
	wire _w9630_ ;
	wire _w9631_ ;
	wire _w9632_ ;
	wire _w9633_ ;
	wire _w9634_ ;
	wire _w9635_ ;
	wire _w9636_ ;
	wire _w9637_ ;
	wire _w9638_ ;
	wire _w9639_ ;
	wire _w9640_ ;
	wire _w9641_ ;
	wire _w9642_ ;
	wire _w9643_ ;
	wire _w9644_ ;
	wire _w9645_ ;
	wire _w9646_ ;
	wire _w9647_ ;
	wire _w9648_ ;
	wire _w9649_ ;
	wire _w9650_ ;
	wire _w9651_ ;
	wire _w9652_ ;
	wire _w9653_ ;
	wire _w9654_ ;
	wire _w9655_ ;
	wire _w9656_ ;
	wire _w9657_ ;
	wire _w9658_ ;
	wire _w9659_ ;
	wire _w9660_ ;
	wire _w9661_ ;
	wire _w9662_ ;
	wire _w9663_ ;
	wire _w9664_ ;
	wire _w9665_ ;
	wire _w9666_ ;
	wire _w9667_ ;
	wire _w9668_ ;
	wire _w9669_ ;
	wire _w9670_ ;
	wire _w9671_ ;
	wire _w9672_ ;
	wire _w9673_ ;
	wire _w9674_ ;
	wire _w9675_ ;
	wire _w9676_ ;
	wire _w9677_ ;
	wire _w9678_ ;
	wire _w9679_ ;
	wire _w9680_ ;
	wire _w9681_ ;
	wire _w9682_ ;
	wire _w9683_ ;
	wire _w9684_ ;
	wire _w9685_ ;
	wire _w9686_ ;
	wire _w9687_ ;
	wire _w9688_ ;
	wire _w9689_ ;
	wire _w9690_ ;
	wire _w9691_ ;
	wire _w9692_ ;
	wire _w9693_ ;
	wire _w9694_ ;
	wire _w9695_ ;
	wire _w9696_ ;
	wire _w9697_ ;
	wire _w9698_ ;
	wire _w9699_ ;
	wire _w9700_ ;
	wire _w9701_ ;
	wire _w9702_ ;
	wire _w9703_ ;
	wire _w9704_ ;
	wire _w9705_ ;
	wire _w9706_ ;
	wire _w9707_ ;
	wire _w9708_ ;
	wire _w9709_ ;
	wire _w9710_ ;
	wire _w9711_ ;
	wire _w9712_ ;
	wire _w9713_ ;
	wire _w9714_ ;
	wire _w9715_ ;
	wire _w9716_ ;
	wire _w9717_ ;
	wire _w9718_ ;
	wire _w9719_ ;
	wire _w9720_ ;
	wire _w9721_ ;
	wire _w9722_ ;
	wire _w9723_ ;
	wire _w9724_ ;
	wire _w9725_ ;
	wire _w9726_ ;
	wire _w9727_ ;
	wire _w9728_ ;
	wire _w9729_ ;
	wire _w9730_ ;
	wire _w9731_ ;
	wire _w9732_ ;
	wire _w9733_ ;
	wire _w9734_ ;
	wire _w9735_ ;
	wire _w9736_ ;
	wire _w9737_ ;
	wire _w9738_ ;
	wire _w9739_ ;
	wire _w9740_ ;
	wire _w9741_ ;
	wire _w9742_ ;
	wire _w9743_ ;
	wire _w9744_ ;
	wire _w9745_ ;
	wire _w9746_ ;
	wire _w9747_ ;
	wire _w9748_ ;
	wire _w9749_ ;
	wire _w9750_ ;
	wire _w9751_ ;
	wire _w9752_ ;
	wire _w9753_ ;
	wire _w9754_ ;
	wire _w9755_ ;
	wire _w9756_ ;
	wire _w9757_ ;
	wire _w9758_ ;
	wire _w9759_ ;
	wire _w9760_ ;
	wire _w9761_ ;
	wire _w9762_ ;
	wire _w9763_ ;
	wire _w9764_ ;
	wire _w9765_ ;
	wire _w9766_ ;
	wire _w9767_ ;
	wire _w9768_ ;
	wire _w9769_ ;
	wire _w9770_ ;
	wire _w9771_ ;
	wire _w9772_ ;
	wire _w9773_ ;
	wire _w9774_ ;
	wire _w9775_ ;
	wire _w9776_ ;
	wire _w9777_ ;
	wire _w9778_ ;
	wire _w9779_ ;
	wire _w9780_ ;
	wire _w9781_ ;
	wire _w9782_ ;
	wire _w9783_ ;
	wire _w9784_ ;
	wire _w9785_ ;
	wire _w9786_ ;
	wire _w9787_ ;
	wire _w9788_ ;
	wire _w9789_ ;
	wire _w9790_ ;
	wire _w9791_ ;
	wire _w9792_ ;
	wire _w9793_ ;
	wire _w9794_ ;
	wire _w9795_ ;
	wire _w9796_ ;
	wire _w9797_ ;
	wire _w9798_ ;
	wire _w9799_ ;
	wire _w9800_ ;
	wire _w9801_ ;
	wire _w9802_ ;
	wire _w9803_ ;
	wire _w9804_ ;
	wire _w9805_ ;
	wire _w9806_ ;
	wire _w9807_ ;
	wire _w9808_ ;
	wire _w9809_ ;
	wire _w9810_ ;
	wire _w9811_ ;
	wire _w9812_ ;
	wire _w9813_ ;
	wire _w9814_ ;
	wire _w9815_ ;
	wire _w9816_ ;
	wire _w9817_ ;
	wire _w9818_ ;
	wire _w9819_ ;
	wire _w9820_ ;
	wire _w9821_ ;
	wire _w9822_ ;
	wire _w9823_ ;
	wire _w9824_ ;
	wire _w9825_ ;
	wire _w9826_ ;
	wire _w9827_ ;
	wire _w9828_ ;
	wire _w9829_ ;
	wire _w9830_ ;
	wire _w9831_ ;
	wire _w9832_ ;
	wire _w9833_ ;
	wire _w9834_ ;
	wire _w9835_ ;
	wire _w9836_ ;
	wire _w9837_ ;
	wire _w9838_ ;
	wire _w9839_ ;
	wire _w9840_ ;
	wire _w9841_ ;
	wire _w9842_ ;
	wire _w9843_ ;
	wire _w9844_ ;
	wire _w9845_ ;
	wire _w9846_ ;
	wire _w9847_ ;
	wire _w9848_ ;
	wire _w9849_ ;
	wire _w9850_ ;
	wire _w9851_ ;
	wire _w9852_ ;
	wire _w9853_ ;
	wire _w9854_ ;
	wire _w9855_ ;
	wire _w9856_ ;
	wire _w9857_ ;
	wire _w9858_ ;
	wire _w9859_ ;
	wire _w9860_ ;
	wire _w9861_ ;
	wire _w9862_ ;
	wire _w9863_ ;
	wire _w9864_ ;
	wire _w9865_ ;
	wire _w9866_ ;
	wire _w9867_ ;
	wire _w9868_ ;
	wire _w9869_ ;
	wire _w9870_ ;
	wire _w9871_ ;
	wire _w9872_ ;
	wire _w9873_ ;
	wire _w9874_ ;
	wire _w9875_ ;
	wire _w9876_ ;
	wire _w9877_ ;
	wire _w9878_ ;
	wire _w9879_ ;
	wire _w9880_ ;
	wire _w9881_ ;
	wire _w9882_ ;
	wire _w9883_ ;
	wire _w9884_ ;
	wire _w9885_ ;
	wire _w9886_ ;
	wire _w9887_ ;
	wire _w9888_ ;
	wire _w9889_ ;
	wire _w9890_ ;
	wire _w9891_ ;
	wire _w9892_ ;
	wire _w9893_ ;
	wire _w9894_ ;
	wire _w9895_ ;
	wire _w9896_ ;
	wire _w9897_ ;
	wire _w9898_ ;
	wire _w9899_ ;
	wire _w9900_ ;
	wire _w9901_ ;
	wire _w9902_ ;
	wire _w9903_ ;
	wire _w9904_ ;
	wire _w9905_ ;
	wire _w9906_ ;
	wire _w9907_ ;
	wire _w9908_ ;
	wire _w9909_ ;
	wire _w9910_ ;
	wire _w9911_ ;
	wire _w9912_ ;
	wire _w9913_ ;
	wire _w9914_ ;
	wire _w9915_ ;
	wire _w9916_ ;
	wire _w9917_ ;
	wire _w9918_ ;
	wire _w9919_ ;
	wire _w9920_ ;
	wire _w9921_ ;
	wire _w9922_ ;
	wire _w9923_ ;
	wire _w9924_ ;
	wire _w9925_ ;
	wire _w9926_ ;
	wire _w9927_ ;
	wire _w9928_ ;
	wire _w9929_ ;
	wire _w9930_ ;
	wire _w9931_ ;
	wire _w9932_ ;
	wire _w9933_ ;
	wire _w9934_ ;
	wire _w9935_ ;
	wire _w9936_ ;
	wire _w9937_ ;
	wire _w9938_ ;
	wire _w9939_ ;
	wire _w9940_ ;
	wire _w9941_ ;
	wire _w9942_ ;
	wire _w9943_ ;
	wire _w9944_ ;
	wire _w9945_ ;
	wire _w9946_ ;
	wire _w9947_ ;
	wire _w9948_ ;
	wire _w9949_ ;
	wire _w9950_ ;
	wire _w9951_ ;
	wire _w9952_ ;
	wire _w9953_ ;
	wire _w9954_ ;
	wire _w9955_ ;
	wire _w9956_ ;
	wire _w9957_ ;
	wire _w9958_ ;
	wire _w9959_ ;
	wire _w9960_ ;
	wire _w9961_ ;
	wire _w9962_ ;
	wire _w9963_ ;
	wire _w9964_ ;
	wire _w9965_ ;
	wire _w9966_ ;
	wire _w9967_ ;
	wire _w9968_ ;
	wire _w9969_ ;
	wire _w9970_ ;
	wire _w9971_ ;
	wire _w9972_ ;
	wire _w9973_ ;
	wire _w9974_ ;
	wire _w9975_ ;
	wire _w9976_ ;
	wire _w9977_ ;
	wire _w9978_ ;
	wire _w9979_ ;
	wire _w9980_ ;
	wire _w9981_ ;
	wire _w9982_ ;
	wire _w9983_ ;
	wire _w9984_ ;
	wire _w9985_ ;
	wire _w9986_ ;
	wire _w9987_ ;
	wire _w9988_ ;
	wire _w9989_ ;
	wire _w9990_ ;
	wire _w9991_ ;
	wire _w9992_ ;
	wire _w9993_ ;
	wire _w9994_ ;
	wire _w9995_ ;
	wire _w9996_ ;
	wire _w9997_ ;
	wire _w9998_ ;
	wire _w9999_ ;
	wire _w10000_ ;
	wire _w10001_ ;
	wire _w10002_ ;
	wire _w10003_ ;
	wire _w10004_ ;
	wire _w10005_ ;
	wire _w10006_ ;
	wire _w10007_ ;
	wire _w10008_ ;
	wire _w10009_ ;
	wire _w10010_ ;
	wire _w10011_ ;
	wire _w10012_ ;
	wire _w10013_ ;
	wire _w10014_ ;
	wire _w10015_ ;
	wire _w10016_ ;
	wire _w10017_ ;
	wire _w10018_ ;
	wire _w10019_ ;
	wire _w10020_ ;
	wire _w10021_ ;
	wire _w10022_ ;
	wire _w10023_ ;
	wire _w10024_ ;
	wire _w10025_ ;
	wire _w10026_ ;
	wire _w10027_ ;
	wire _w10028_ ;
	wire _w10029_ ;
	wire _w10030_ ;
	wire _w10031_ ;
	wire _w10032_ ;
	wire _w10033_ ;
	wire _w10034_ ;
	wire _w10035_ ;
	wire _w10036_ ;
	wire _w10037_ ;
	wire _w10038_ ;
	wire _w10039_ ;
	wire _w10040_ ;
	wire _w10041_ ;
	wire _w10042_ ;
	wire _w10043_ ;
	wire _w10044_ ;
	wire _w10045_ ;
	wire _w10046_ ;
	wire _w10047_ ;
	wire _w10048_ ;
	wire _w10049_ ;
	wire _w10050_ ;
	wire _w10051_ ;
	wire _w10052_ ;
	wire _w10053_ ;
	wire _w10054_ ;
	wire _w10055_ ;
	wire _w10056_ ;
	wire _w10057_ ;
	wire _w10058_ ;
	wire _w10059_ ;
	wire _w10060_ ;
	wire _w10061_ ;
	wire _w10062_ ;
	wire _w10063_ ;
	wire _w10064_ ;
	wire _w10065_ ;
	wire _w10066_ ;
	wire _w10067_ ;
	wire _w10068_ ;
	wire _w10069_ ;
	wire _w10070_ ;
	wire _w10071_ ;
	wire _w10072_ ;
	wire _w10073_ ;
	wire _w10074_ ;
	wire _w10075_ ;
	wire _w10076_ ;
	wire _w10077_ ;
	wire _w10078_ ;
	wire _w10079_ ;
	wire _w10080_ ;
	wire _w10081_ ;
	wire _w10082_ ;
	wire _w10083_ ;
	wire _w10084_ ;
	wire _w10085_ ;
	wire _w10086_ ;
	wire _w10087_ ;
	wire _w10088_ ;
	wire _w10089_ ;
	wire _w10090_ ;
	wire _w10091_ ;
	wire _w10092_ ;
	wire _w10093_ ;
	wire _w10094_ ;
	wire _w10095_ ;
	wire _w10096_ ;
	wire _w10097_ ;
	wire _w10098_ ;
	wire _w10099_ ;
	wire _w10100_ ;
	wire _w10101_ ;
	wire _w10102_ ;
	wire _w10103_ ;
	wire _w10104_ ;
	wire _w10105_ ;
	wire _w10106_ ;
	wire _w10107_ ;
	wire _w10108_ ;
	wire _w10109_ ;
	wire _w10110_ ;
	wire _w10111_ ;
	wire _w10112_ ;
	wire _w10113_ ;
	wire _w10114_ ;
	wire _w10115_ ;
	wire _w10116_ ;
	wire _w10117_ ;
	wire _w10118_ ;
	wire _w10119_ ;
	wire _w10120_ ;
	wire _w10121_ ;
	wire _w10122_ ;
	wire _w10123_ ;
	wire _w10124_ ;
	wire _w10125_ ;
	wire _w10126_ ;
	wire _w10127_ ;
	wire _w10128_ ;
	wire _w10129_ ;
	wire _w10130_ ;
	wire _w10131_ ;
	wire _w10132_ ;
	wire _w10133_ ;
	wire _w10134_ ;
	wire _w10135_ ;
	wire _w10136_ ;
	wire _w10137_ ;
	wire _w10138_ ;
	wire _w10139_ ;
	wire _w10140_ ;
	wire _w10141_ ;
	wire _w10142_ ;
	wire _w10143_ ;
	wire _w10144_ ;
	wire _w10145_ ;
	wire _w10146_ ;
	wire _w10147_ ;
	wire _w10148_ ;
	wire _w10149_ ;
	wire _w10150_ ;
	wire _w10151_ ;
	wire _w10152_ ;
	wire _w10153_ ;
	wire _w10154_ ;
	wire _w10155_ ;
	wire _w10156_ ;
	wire _w10157_ ;
	wire _w10158_ ;
	wire _w10159_ ;
	wire _w10160_ ;
	wire _w10161_ ;
	wire _w10162_ ;
	wire _w10163_ ;
	wire _w10164_ ;
	wire _w10165_ ;
	wire _w10166_ ;
	wire _w10167_ ;
	wire _w10168_ ;
	wire _w10169_ ;
	wire _w10170_ ;
	wire _w10171_ ;
	wire _w10172_ ;
	wire _w10173_ ;
	wire _w10174_ ;
	wire _w10175_ ;
	wire _w10176_ ;
	wire _w10177_ ;
	wire _w10178_ ;
	wire _w10179_ ;
	wire _w10180_ ;
	wire _w10181_ ;
	wire _w10182_ ;
	wire _w10183_ ;
	wire _w10184_ ;
	wire _w10185_ ;
	wire _w10186_ ;
	wire _w10187_ ;
	wire _w10188_ ;
	wire _w10189_ ;
	wire _w10190_ ;
	wire _w10191_ ;
	wire _w10192_ ;
	wire _w10193_ ;
	wire _w10194_ ;
	wire _w10195_ ;
	wire _w10196_ ;
	wire _w10197_ ;
	wire _w10198_ ;
	wire _w10199_ ;
	wire _w10200_ ;
	wire _w10201_ ;
	wire _w10202_ ;
	wire _w10203_ ;
	wire _w10204_ ;
	wire _w10205_ ;
	wire _w10206_ ;
	wire _w10207_ ;
	wire _w10208_ ;
	wire _w10209_ ;
	wire _w10210_ ;
	wire _w10211_ ;
	wire _w10212_ ;
	wire _w10213_ ;
	wire _w10214_ ;
	wire _w10215_ ;
	wire _w10216_ ;
	wire _w10217_ ;
	wire _w10218_ ;
	wire _w10219_ ;
	wire _w10220_ ;
	wire _w10221_ ;
	wire _w10222_ ;
	wire _w10223_ ;
	wire _w10224_ ;
	wire _w10225_ ;
	wire _w10226_ ;
	wire _w10227_ ;
	wire _w10228_ ;
	wire _w10229_ ;
	wire _w10230_ ;
	wire _w10231_ ;
	wire _w10232_ ;
	wire _w10233_ ;
	wire _w10234_ ;
	wire _w10235_ ;
	wire _w10236_ ;
	wire _w10237_ ;
	wire _w10238_ ;
	wire _w10239_ ;
	wire _w10240_ ;
	wire _w10241_ ;
	wire _w10242_ ;
	wire _w10243_ ;
	wire _w10244_ ;
	wire _w10245_ ;
	wire _w10246_ ;
	wire _w10247_ ;
	wire _w10248_ ;
	wire _w10249_ ;
	wire _w10250_ ;
	wire _w10251_ ;
	wire _w10252_ ;
	wire _w10253_ ;
	wire _w10254_ ;
	wire _w10255_ ;
	wire _w10256_ ;
	wire _w10257_ ;
	wire _w10258_ ;
	wire _w10259_ ;
	wire _w10260_ ;
	wire _w10261_ ;
	wire _w10262_ ;
	wire _w10263_ ;
	wire _w10264_ ;
	wire _w10265_ ;
	wire _w10266_ ;
	wire _w10267_ ;
	wire _w10268_ ;
	wire _w10269_ ;
	wire _w10270_ ;
	wire _w10271_ ;
	wire _w10272_ ;
	wire _w10273_ ;
	wire _w10274_ ;
	wire _w10275_ ;
	wire _w10276_ ;
	wire _w10277_ ;
	wire _w10278_ ;
	wire _w10279_ ;
	wire _w10280_ ;
	wire _w10281_ ;
	wire _w10282_ ;
	wire _w10283_ ;
	wire _w10284_ ;
	wire _w10285_ ;
	wire _w10286_ ;
	wire _w10287_ ;
	wire _w10288_ ;
	wire _w10289_ ;
	wire _w10290_ ;
	wire _w10291_ ;
	wire _w10292_ ;
	wire _w10293_ ;
	wire _w10294_ ;
	wire _w10295_ ;
	wire _w10296_ ;
	wire _w10297_ ;
	wire _w10298_ ;
	wire _w10299_ ;
	wire _w10300_ ;
	wire _w10301_ ;
	wire _w10302_ ;
	wire _w10303_ ;
	wire _w10304_ ;
	wire _w10305_ ;
	wire _w10306_ ;
	wire _w10307_ ;
	wire _w10308_ ;
	wire _w10309_ ;
	wire _w10310_ ;
	wire _w10311_ ;
	wire _w10312_ ;
	wire _w10313_ ;
	wire _w10314_ ;
	wire _w10315_ ;
	wire _w10316_ ;
	wire _w10317_ ;
	wire _w10318_ ;
	wire _w10319_ ;
	wire _w10320_ ;
	wire _w10321_ ;
	wire _w10322_ ;
	wire _w10323_ ;
	wire _w10324_ ;
	wire _w10325_ ;
	wire _w10326_ ;
	wire _w10327_ ;
	wire _w10328_ ;
	wire _w10329_ ;
	wire _w10330_ ;
	wire _w10331_ ;
	wire _w10332_ ;
	wire _w10333_ ;
	wire _w10334_ ;
	wire _w10335_ ;
	wire _w10336_ ;
	wire _w10337_ ;
	wire _w10338_ ;
	wire _w10339_ ;
	wire _w10340_ ;
	wire _w10341_ ;
	wire _w10342_ ;
	wire _w10343_ ;
	wire _w10344_ ;
	wire _w10345_ ;
	wire _w10346_ ;
	wire _w10347_ ;
	wire _w10348_ ;
	wire _w10349_ ;
	wire _w10350_ ;
	wire _w10351_ ;
	wire _w10352_ ;
	wire _w10353_ ;
	wire _w10354_ ;
	wire _w10355_ ;
	wire _w10356_ ;
	wire _w10357_ ;
	wire _w10358_ ;
	wire _w10359_ ;
	wire _w10360_ ;
	wire _w10361_ ;
	wire _w10362_ ;
	wire _w10363_ ;
	wire _w10364_ ;
	wire _w10365_ ;
	wire _w10366_ ;
	wire _w10367_ ;
	wire _w10368_ ;
	wire _w10369_ ;
	wire _w10370_ ;
	wire _w10371_ ;
	wire _w10372_ ;
	wire _w10373_ ;
	wire _w10374_ ;
	wire _w10375_ ;
	wire _w10376_ ;
	wire _w10377_ ;
	wire _w10378_ ;
	wire _w10379_ ;
	wire _w10380_ ;
	wire _w10381_ ;
	wire _w10382_ ;
	wire _w10383_ ;
	wire _w10384_ ;
	wire _w10385_ ;
	wire _w10386_ ;
	wire _w10387_ ;
	wire _w10388_ ;
	wire _w10389_ ;
	wire _w10390_ ;
	wire _w10391_ ;
	wire _w10392_ ;
	wire _w10393_ ;
	wire _w10394_ ;
	wire _w10395_ ;
	wire _w10396_ ;
	wire _w10397_ ;
	wire _w10398_ ;
	wire _w10399_ ;
	wire _w10400_ ;
	wire _w10401_ ;
	wire _w10402_ ;
	wire _w10403_ ;
	wire _w10404_ ;
	wire _w10405_ ;
	wire _w10406_ ;
	wire _w10407_ ;
	wire _w10408_ ;
	wire _w10409_ ;
	wire _w10410_ ;
	wire _w10411_ ;
	wire _w10412_ ;
	wire _w10413_ ;
	wire _w10414_ ;
	wire _w10415_ ;
	wire _w10416_ ;
	wire _w10417_ ;
	wire _w10418_ ;
	wire _w10419_ ;
	wire _w10420_ ;
	wire _w10421_ ;
	wire _w10422_ ;
	wire _w10423_ ;
	wire _w10424_ ;
	wire _w10425_ ;
	wire _w10426_ ;
	wire _w10427_ ;
	wire _w10428_ ;
	wire _w10429_ ;
	wire _w10430_ ;
	wire _w10431_ ;
	wire _w10432_ ;
	wire _w10433_ ;
	wire _w10434_ ;
	wire _w10435_ ;
	wire _w10436_ ;
	wire _w10437_ ;
	wire _w10438_ ;
	wire _w10439_ ;
	wire _w10440_ ;
	wire _w10441_ ;
	wire _w10442_ ;
	wire _w10443_ ;
	wire _w10444_ ;
	wire _w10445_ ;
	wire _w10446_ ;
	wire _w10447_ ;
	wire _w10448_ ;
	wire _w10449_ ;
	wire _w10450_ ;
	wire _w10451_ ;
	wire _w10452_ ;
	wire _w10453_ ;
	wire _w10454_ ;
	wire _w10455_ ;
	wire _w10456_ ;
	wire _w10457_ ;
	wire _w10458_ ;
	wire _w10459_ ;
	wire _w10460_ ;
	wire _w10461_ ;
	wire _w10462_ ;
	wire _w10463_ ;
	wire _w10464_ ;
	wire _w10465_ ;
	wire _w10466_ ;
	wire _w10467_ ;
	wire _w10468_ ;
	wire _w10469_ ;
	wire _w10470_ ;
	wire _w10471_ ;
	wire _w10472_ ;
	wire _w10473_ ;
	wire _w10474_ ;
	wire _w10475_ ;
	wire _w10476_ ;
	wire _w10477_ ;
	wire _w10478_ ;
	wire _w10479_ ;
	wire _w10480_ ;
	wire _w10481_ ;
	wire _w10482_ ;
	wire _w10483_ ;
	wire _w10484_ ;
	wire _w10485_ ;
	wire _w10486_ ;
	wire _w10487_ ;
	wire _w10488_ ;
	wire _w10489_ ;
	wire _w10490_ ;
	wire _w10491_ ;
	wire _w10492_ ;
	wire _w10493_ ;
	wire _w10494_ ;
	wire _w10495_ ;
	wire _w10496_ ;
	wire _w10497_ ;
	wire _w10498_ ;
	wire _w10499_ ;
	wire _w10500_ ;
	wire _w10501_ ;
	wire _w10502_ ;
	wire _w10503_ ;
	wire _w10504_ ;
	wire _w10505_ ;
	wire _w10506_ ;
	wire _w10507_ ;
	wire _w10508_ ;
	wire _w10509_ ;
	wire _w10510_ ;
	wire _w10511_ ;
	wire _w10512_ ;
	wire _w10513_ ;
	wire _w10514_ ;
	wire _w10515_ ;
	wire _w10516_ ;
	wire _w10517_ ;
	wire _w10518_ ;
	wire _w10519_ ;
	wire _w10520_ ;
	wire _w10521_ ;
	wire _w10522_ ;
	wire _w10523_ ;
	wire _w10524_ ;
	wire _w10525_ ;
	wire _w10526_ ;
	wire _w10527_ ;
	wire _w10528_ ;
	wire _w10529_ ;
	wire _w10530_ ;
	wire _w10531_ ;
	wire _w10532_ ;
	wire _w10533_ ;
	wire _w10534_ ;
	wire _w10535_ ;
	wire _w10536_ ;
	wire _w10537_ ;
	wire _w10538_ ;
	wire _w10539_ ;
	wire _w10540_ ;
	wire _w10541_ ;
	wire _w10542_ ;
	wire _w10543_ ;
	wire _w10544_ ;
	wire _w10545_ ;
	wire _w10546_ ;
	wire _w10547_ ;
	wire _w10548_ ;
	wire _w10549_ ;
	wire _w10550_ ;
	wire _w10551_ ;
	wire _w10552_ ;
	wire _w10553_ ;
	wire _w10554_ ;
	wire _w10555_ ;
	wire _w10556_ ;
	wire _w10557_ ;
	wire _w10558_ ;
	wire _w10559_ ;
	wire _w10560_ ;
	wire _w10561_ ;
	wire _w10562_ ;
	wire _w10563_ ;
	wire _w10564_ ;
	wire _w10565_ ;
	wire _w10566_ ;
	wire _w10567_ ;
	wire _w10568_ ;
	wire _w10569_ ;
	wire _w10570_ ;
	wire _w10571_ ;
	wire _w10572_ ;
	wire _w10573_ ;
	wire _w10574_ ;
	wire _w10575_ ;
	wire _w10576_ ;
	wire _w10577_ ;
	wire _w10578_ ;
	wire _w10579_ ;
	wire _w10580_ ;
	wire _w10581_ ;
	wire _w10582_ ;
	wire _w10583_ ;
	wire _w10584_ ;
	wire _w10585_ ;
	wire _w10586_ ;
	wire _w10587_ ;
	wire _w10588_ ;
	wire _w10589_ ;
	wire _w10590_ ;
	wire _w10591_ ;
	wire _w10592_ ;
	wire _w10593_ ;
	wire _w10594_ ;
	wire _w10595_ ;
	wire _w10596_ ;
	wire _w10597_ ;
	wire _w10598_ ;
	wire _w10599_ ;
	wire _w10600_ ;
	wire _w10601_ ;
	wire _w10602_ ;
	wire _w10603_ ;
	wire _w10604_ ;
	wire _w10605_ ;
	wire _w10606_ ;
	wire _w10607_ ;
	wire _w10608_ ;
	wire _w10609_ ;
	wire _w10610_ ;
	wire _w10611_ ;
	wire _w10612_ ;
	wire _w10613_ ;
	wire _w10614_ ;
	wire _w10615_ ;
	wire _w10616_ ;
	wire _w10617_ ;
	wire _w10618_ ;
	wire _w10619_ ;
	wire _w10620_ ;
	wire _w10621_ ;
	wire _w10622_ ;
	wire _w10623_ ;
	wire _w10624_ ;
	wire _w10625_ ;
	wire _w10626_ ;
	wire _w10627_ ;
	wire _w10628_ ;
	wire _w10629_ ;
	wire _w10630_ ;
	wire _w10631_ ;
	wire _w10632_ ;
	wire _w10633_ ;
	wire _w10634_ ;
	wire _w10635_ ;
	wire _w10636_ ;
	wire _w10637_ ;
	wire _w10638_ ;
	wire _w10639_ ;
	wire _w10640_ ;
	wire _w10641_ ;
	wire _w10642_ ;
	wire _w10643_ ;
	wire _w10644_ ;
	wire _w10645_ ;
	wire _w10646_ ;
	wire _w10647_ ;
	wire _w10648_ ;
	wire _w10649_ ;
	wire _w10650_ ;
	wire _w10651_ ;
	wire _w10652_ ;
	wire _w10653_ ;
	wire _w10654_ ;
	wire _w10655_ ;
	wire _w10656_ ;
	wire _w10657_ ;
	wire _w10658_ ;
	wire _w10659_ ;
	wire _w10660_ ;
	wire _w10661_ ;
	wire _w10662_ ;
	wire _w10663_ ;
	wire _w10664_ ;
	wire _w10665_ ;
	wire _w10666_ ;
	wire _w10667_ ;
	wire _w10668_ ;
	wire _w10669_ ;
	wire _w10670_ ;
	wire _w10671_ ;
	wire _w10672_ ;
	wire _w10673_ ;
	wire _w10674_ ;
	wire _w10675_ ;
	wire _w10676_ ;
	wire _w10677_ ;
	wire _w10678_ ;
	wire _w10679_ ;
	wire _w10680_ ;
	wire _w10681_ ;
	wire _w10682_ ;
	wire _w10683_ ;
	wire _w10684_ ;
	wire _w10685_ ;
	wire _w10686_ ;
	wire _w10687_ ;
	wire _w10688_ ;
	wire _w10689_ ;
	wire _w10690_ ;
	wire _w10691_ ;
	wire _w10692_ ;
	wire _w10693_ ;
	wire _w10694_ ;
	wire _w10695_ ;
	wire _w10696_ ;
	wire _w10697_ ;
	wire _w10698_ ;
	wire _w10699_ ;
	wire _w10700_ ;
	wire _w10701_ ;
	wire _w10702_ ;
	wire _w10703_ ;
	wire _w10704_ ;
	wire _w10705_ ;
	wire _w10706_ ;
	wire _w10707_ ;
	wire _w10708_ ;
	wire _w10709_ ;
	wire _w10710_ ;
	wire _w10711_ ;
	wire _w10712_ ;
	wire _w10713_ ;
	wire _w10714_ ;
	wire _w10715_ ;
	wire _w10716_ ;
	wire _w10717_ ;
	wire _w10718_ ;
	wire _w10719_ ;
	wire _w10720_ ;
	wire _w10721_ ;
	wire _w10722_ ;
	wire _w10723_ ;
	wire _w10724_ ;
	wire _w10725_ ;
	wire _w10726_ ;
	wire _w10727_ ;
	wire _w10728_ ;
	wire _w10729_ ;
	wire _w10730_ ;
	wire _w10731_ ;
	wire _w10732_ ;
	wire _w10733_ ;
	wire _w10734_ ;
	wire _w10735_ ;
	wire _w10736_ ;
	wire _w10737_ ;
	wire _w10738_ ;
	wire _w10739_ ;
	wire _w10740_ ;
	wire _w10741_ ;
	wire _w10742_ ;
	wire _w10743_ ;
	wire _w10744_ ;
	wire _w10745_ ;
	wire _w10746_ ;
	wire _w10747_ ;
	wire _w10748_ ;
	wire _w10749_ ;
	wire _w10750_ ;
	wire _w10751_ ;
	wire _w10752_ ;
	wire _w10753_ ;
	wire _w10754_ ;
	wire _w10755_ ;
	wire _w10756_ ;
	wire _w10757_ ;
	wire _w10758_ ;
	wire _w10759_ ;
	wire _w10760_ ;
	wire _w10761_ ;
	wire _w10762_ ;
	wire _w10763_ ;
	wire _w10764_ ;
	wire _w10765_ ;
	wire _w10766_ ;
	wire _w10767_ ;
	wire _w10768_ ;
	wire _w10769_ ;
	wire _w10770_ ;
	wire _w10771_ ;
	wire _w10772_ ;
	wire _w10773_ ;
	wire _w10774_ ;
	wire _w10775_ ;
	wire _w10776_ ;
	wire _w10777_ ;
	wire _w10778_ ;
	wire _w10779_ ;
	wire _w10780_ ;
	wire _w10781_ ;
	wire _w10782_ ;
	wire _w10783_ ;
	wire _w10784_ ;
	wire _w10785_ ;
	wire _w10786_ ;
	wire _w10787_ ;
	wire _w10788_ ;
	wire _w10789_ ;
	wire _w10790_ ;
	wire _w10791_ ;
	wire _w10792_ ;
	wire _w10793_ ;
	wire _w10794_ ;
	wire _w10795_ ;
	wire _w10796_ ;
	wire _w10797_ ;
	wire _w10798_ ;
	wire _w10799_ ;
	wire _w10800_ ;
	wire _w10801_ ;
	wire _w10802_ ;
	wire _w10803_ ;
	wire _w10804_ ;
	wire _w10805_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w533_
	);
	LUT4 #(
		.INIT('h1000)
	) name1 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w534_
	);
	LUT2 #(
		.INIT('h2)
	) name2 (
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w535_
	);
	LUT3 #(
		.INIT('h08)
	) name3 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w536_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w537_
	);
	LUT3 #(
		.INIT('h20)
	) name5 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w538_
	);
	LUT4 #(
		.INIT('h0400)
	) name6 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w539_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name7 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w540_
	);
	LUT4 #(
		.INIT('h20aa)
	) name8 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w534_,
		_w540_,
		_w541_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w542_
	);
	LUT3 #(
		.INIT('h02)
	) name10 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w543_
	);
	LUT3 #(
		.INIT('h80)
	) name11 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w544_
	);
	LUT4 #(
		.INIT('h2000)
	) name12 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w545_
	);
	LUT3 #(
		.INIT('h07)
	) name13 (
		_w542_,
		_w543_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[5]/P0001 ,
		_w547_
	);
	LUT3 #(
		.INIT('h01)
	) name15 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		_w548_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		_w533_,
		_w548_,
		_w549_
	);
	LUT4 #(
		.INIT('haaa2)
	) name17 (
		\sa13_reg[1]/P0001 ,
		_w546_,
		_w549_,
		_w541_,
		_w550_
	);
	LUT4 #(
		.INIT('h0004)
	) name18 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		\sa13_reg[2]/P0001 ,
		_w551_,
		_w552_
	);
	LUT3 #(
		.INIT('h80)
	) name20 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w553_
	);
	LUT3 #(
		.INIT('h04)
	) name21 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w554_
	);
	LUT4 #(
		.INIT('heee4)
	) name22 (
		\sa13_reg[2]/P0001 ,
		_w551_,
		_w554_,
		_w553_,
		_w555_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w556_
	);
	LUT3 #(
		.INIT('h02)
	) name24 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w557_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w558_
	);
	LUT3 #(
		.INIT('h40)
	) name26 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w559_
	);
	LUT4 #(
		.INIT('h153f)
	) name27 (
		_w547_,
		_w557_,
		_w558_,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w561_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w562_
	);
	LUT4 #(
		.INIT('h0800)
	) name30 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w563_
	);
	LUT4 #(
		.INIT('h5551)
	) name31 (
		\sa13_reg[1]/P0001 ,
		_w560_,
		_w563_,
		_w555_,
		_w564_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w565_
	);
	LUT4 #(
		.INIT('h0040)
	) name33 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w566_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w567_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w568_
	);
	LUT4 #(
		.INIT('h0040)
	) name36 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w569_
	);
	LUT3 #(
		.INIT('h54)
	) name37 (
		\sa13_reg[2]/P0001 ,
		_w566_,
		_w569_,
		_w570_
	);
	LUT3 #(
		.INIT('h80)
	) name38 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w571_
	);
	LUT4 #(
		.INIT('h4000)
	) name39 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w572_
	);
	LUT3 #(
		.INIT('h08)
	) name40 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w573_
	);
	LUT4 #(
		.INIT('h0080)
	) name41 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w574_
	);
	LUT3 #(
		.INIT('h07)
	) name42 (
		\sa13_reg[4]/P0001 ,
		_w572_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w576_
	);
	LUT4 #(
		.INIT('h0001)
	) name44 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w577_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		_w578_
	);
	LUT4 #(
		.INIT('h0200)
	) name46 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w579_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w577_,
		_w579_,
		_w580_
	);
	LUT4 #(
		.INIT('h3111)
	) name48 (
		\sa13_reg[2]/P0001 ,
		_w570_,
		_w575_,
		_w580_,
		_w581_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name49 (
		\sa13_reg[0]/P0001 ,
		_w550_,
		_w564_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w583_
	);
	LUT3 #(
		.INIT('h01)
	) name51 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w584_
	);
	LUT3 #(
		.INIT('h80)
	) name52 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w585_
	);
	LUT3 #(
		.INIT('h7e)
	) name53 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w586_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		_w583_,
		_w586_,
		_w587_
	);
	LUT3 #(
		.INIT('h01)
	) name55 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w588_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w589_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w588_,
		_w589_,
		_w590_
	);
	LUT3 #(
		.INIT('h80)
	) name58 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		_w591_
	);
	LUT3 #(
		.INIT('h2a)
	) name59 (
		\sa13_reg[1]/P0001 ,
		_w535_,
		_w591_,
		_w592_
	);
	LUT3 #(
		.INIT('h10)
	) name60 (
		_w587_,
		_w590_,
		_w592_,
		_w593_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w594_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		_w543_,
		_w594_,
		_w595_
	);
	LUT4 #(
		.INIT('h4000)
	) name63 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w596_
	);
	LUT3 #(
		.INIT('h01)
	) name64 (
		\sa13_reg[1]/P0001 ,
		_w569_,
		_w596_,
		_w597_
	);
	LUT3 #(
		.INIT('h10)
	) name65 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w598_
	);
	LUT4 #(
		.INIT('hd8ff)
	) name66 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w599_
	);
	LUT4 #(
		.INIT('h0400)
	) name67 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w600_
	);
	LUT4 #(
		.INIT('h32fa)
	) name68 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w599_,
		_w600_,
		_w601_
	);
	LUT3 #(
		.INIT('h40)
	) name69 (
		_w595_,
		_w597_,
		_w601_,
		_w602_
	);
	LUT4 #(
		.INIT('h0004)
	) name70 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w603_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		\sa13_reg[2]/P0001 ,
		_w603_,
		_w604_
	);
	LUT4 #(
		.INIT('h2220)
	) name72 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w605_
	);
	LUT3 #(
		.INIT('h2a)
	) name73 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w606_
	);
	LUT3 #(
		.INIT('h04)
	) name74 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w607_
	);
	LUT4 #(
		.INIT('h51f3)
	) name75 (
		_w567_,
		_w605_,
		_w606_,
		_w607_,
		_w608_
	);
	LUT4 #(
		.INIT('h0001)
	) name76 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w609_
	);
	LUT4 #(
		.INIT('h002a)
	) name77 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w600_,
		_w609_,
		_w610_
	);
	LUT3 #(
		.INIT('h07)
	) name78 (
		_w604_,
		_w608_,
		_w610_,
		_w611_
	);
	LUT4 #(
		.INIT('h5501)
	) name79 (
		\sa13_reg[0]/P0001 ,
		_w593_,
		_w602_,
		_w611_,
		_w612_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w613_
	);
	LUT3 #(
		.INIT('h20)
	) name81 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		_w614_
	);
	LUT4 #(
		.INIT('h0002)
	) name82 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w615_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w616_
	);
	LUT4 #(
		.INIT('h0001)
	) name84 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w617_
	);
	LUT4 #(
		.INIT('h0103)
	) name85 (
		_w537_,
		_w615_,
		_w617_,
		_w614_,
		_w618_
	);
	LUT4 #(
		.INIT('h0020)
	) name86 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w619_
	);
	LUT4 #(
		.INIT('h0001)
	) name87 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w620_
	);
	LUT3 #(
		.INIT('h07)
	) name88 (
		\sa13_reg[4]/P0001 ,
		_w619_,
		_w620_,
		_w621_
	);
	LUT4 #(
		.INIT('h08cc)
	) name89 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[2]/P0001 ,
		_w618_,
		_w621_,
		_w622_
	);
	LUT4 #(
		.INIT('h0020)
	) name90 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w623_
	);
	LUT4 #(
		.INIT('h5504)
	) name91 (
		\sa13_reg[2]/P0001 ,
		_w538_,
		_w616_,
		_w623_,
		_w624_
	);
	LUT4 #(
		.INIT('h1000)
	) name92 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w625_
	);
	LUT4 #(
		.INIT('h0800)
	) name93 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w626_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w625_,
		_w626_,
		_w627_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w628_
	);
	LUT3 #(
		.INIT('h01)
	) name96 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w629_
	);
	LUT4 #(
		.INIT('h135f)
	) name97 (
		_w571_,
		_w594_,
		_w628_,
		_w629_,
		_w630_
	);
	LUT4 #(
		.INIT('h4555)
	) name98 (
		\sa13_reg[1]/P0001 ,
		_w624_,
		_w627_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h2)
	) name99 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[2]/P0001 ,
		_w632_
	);
	LUT3 #(
		.INIT('h80)
	) name100 (
		_w543_,
		_w613_,
		_w632_,
		_w633_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name101 (
		\sa13_reg[5]/P0001 ,
		_w558_,
		_w563_,
		_w617_,
		_w634_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		_w633_,
		_w634_,
		_w635_
	);
	LUT3 #(
		.INIT('h10)
	) name103 (
		_w622_,
		_w631_,
		_w635_,
		_w636_
	);
	LUT3 #(
		.INIT('h10)
	) name104 (
		_w582_,
		_w612_,
		_w636_,
		_w637_
	);
	LUT2 #(
		.INIT('h4)
	) name105 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w638_
	);
	LUT2 #(
		.INIT('h4)
	) name106 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w639_
	);
	LUT4 #(
		.INIT('h1000)
	) name107 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w640_
	);
	LUT3 #(
		.INIT('h08)
	) name108 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w641_
	);
	LUT2 #(
		.INIT('h4)
	) name109 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		_w642_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w643_
	);
	LUT4 #(
		.INIT('h0400)
	) name111 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w644_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name112 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w645_
	);
	LUT4 #(
		.INIT('h20aa)
	) name113 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w640_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w647_
	);
	LUT3 #(
		.INIT('h08)
	) name115 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w648_
	);
	LUT4 #(
		.INIT('h0080)
	) name116 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w649_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		\sa20_reg[7]/NET0131 ,
		_w649_,
		_w650_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w651_
	);
	LUT2 #(
		.INIT('h2)
	) name119 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w652_
	);
	LUT4 #(
		.INIT('h2000)
	) name120 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w653_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		_w654_
	);
	LUT2 #(
		.INIT('h4)
	) name122 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w655_
	);
	LUT3 #(
		.INIT('h23)
	) name123 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w656_
	);
	LUT3 #(
		.INIT('h15)
	) name124 (
		_w653_,
		_w654_,
		_w656_,
		_w657_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name125 (
		\sa20_reg[1]/P0001 ,
		_w646_,
		_w650_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w659_
	);
	LUT4 #(
		.INIT('h0008)
	) name127 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w660_
	);
	LUT4 #(
		.INIT('h1000)
	) name128 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w661_
	);
	LUT3 #(
		.INIT('h02)
	) name129 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w662_
	);
	LUT4 #(
		.INIT('h0004)
	) name130 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w663_
	);
	LUT4 #(
		.INIT('h5554)
	) name131 (
		\sa20_reg[2]/P0001 ,
		_w660_,
		_w661_,
		_w663_,
		_w664_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w665_
	);
	LUT4 #(
		.INIT('h0800)
	) name133 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w666_
	);
	LUT3 #(
		.INIT('h04)
	) name134 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w667_
	);
	LUT3 #(
		.INIT('h80)
	) name135 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w668_
	);
	LUT4 #(
		.INIT('h1113)
	) name136 (
		\sa20_reg[2]/P0001 ,
		_w666_,
		_w667_,
		_w668_,
		_w669_
	);
	LUT3 #(
		.INIT('h45)
	) name137 (
		\sa20_reg[1]/P0001 ,
		_w664_,
		_w669_,
		_w670_
	);
	LUT2 #(
		.INIT('h4)
	) name138 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w671_
	);
	LUT4 #(
		.INIT('h0040)
	) name139 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w672_
	);
	LUT4 #(
		.INIT('h0040)
	) name140 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w673_
	);
	LUT3 #(
		.INIT('h54)
	) name141 (
		\sa20_reg[2]/P0001 ,
		_w672_,
		_w673_,
		_w674_
	);
	LUT3 #(
		.INIT('h08)
	) name142 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w675_
	);
	LUT4 #(
		.INIT('h0080)
	) name143 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w676_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w677_
	);
	LUT4 #(
		.INIT('h4000)
	) name145 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w678_
	);
	LUT3 #(
		.INIT('h13)
	) name146 (
		\sa20_reg[7]/NET0131 ,
		_w676_,
		_w678_,
		_w679_
	);
	LUT4 #(
		.INIT('h0200)
	) name147 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w680_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w681_
	);
	LUT4 #(
		.INIT('h0001)
	) name149 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w682_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		_w680_,
		_w682_,
		_w683_
	);
	LUT4 #(
		.INIT('h3111)
	) name151 (
		\sa20_reg[2]/P0001 ,
		_w674_,
		_w679_,
		_w683_,
		_w684_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name152 (
		\sa20_reg[0]/P0001 ,
		_w670_,
		_w658_,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		_w686_
	);
	LUT4 #(
		.INIT('h4000)
	) name154 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w687_
	);
	LUT4 #(
		.INIT('h0200)
	) name155 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w688_
	);
	LUT4 #(
		.INIT('h0001)
	) name156 (
		\sa20_reg[1]/P0001 ,
		_w673_,
		_w687_,
		_w688_,
		_w689_
	);
	LUT3 #(
		.INIT('h10)
	) name157 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w690_
	);
	LUT4 #(
		.INIT('h0100)
	) name158 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w691_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		_w692_
	);
	LUT3 #(
		.INIT('h20)
	) name160 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w693_
	);
	LUT4 #(
		.INIT('h135f)
	) name161 (
		_w662_,
		_w639_,
		_w692_,
		_w693_,
		_w694_
	);
	LUT3 #(
		.INIT('h40)
	) name162 (
		_w691_,
		_w689_,
		_w694_,
		_w695_
	);
	LUT3 #(
		.INIT('h80)
	) name163 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w696_
	);
	LUT3 #(
		.INIT('h01)
	) name164 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w697_
	);
	LUT3 #(
		.INIT('h7e)
	) name165 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w698_
	);
	LUT4 #(
		.INIT('h0072)
	) name166 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		_w682_,
		_w698_,
		_w699_
	);
	LUT2 #(
		.INIT('h2)
	) name167 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w700_
	);
	LUT4 #(
		.INIT('h0080)
	) name168 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w701_
	);
	LUT3 #(
		.INIT('h2a)
	) name169 (
		\sa20_reg[1]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h4)
	) name170 (
		_w699_,
		_w702_,
		_w703_
	);
	LUT3 #(
		.INIT('h02)
	) name171 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w704_
	);
	LUT4 #(
		.INIT('h2220)
	) name172 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w705_
	);
	LUT3 #(
		.INIT('h54)
	) name173 (
		_w647_,
		_w704_,
		_w705_,
		_w706_
	);
	LUT3 #(
		.INIT('h04)
	) name174 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w707_
	);
	LUT4 #(
		.INIT('h2000)
	) name175 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w708_
	);
	LUT4 #(
		.INIT('h0015)
	) name176 (
		\sa20_reg[2]/P0001 ,
		_w677_,
		_w707_,
		_w708_,
		_w709_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w710_
	);
	LUT4 #(
		.INIT('h0001)
	) name178 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w711_
	);
	LUT4 #(
		.INIT('h002a)
	) name179 (
		\sa20_reg[2]/P0001 ,
		_w639_,
		_w693_,
		_w711_,
		_w712_
	);
	LUT3 #(
		.INIT('h0b)
	) name180 (
		_w706_,
		_w709_,
		_w712_,
		_w713_
	);
	LUT4 #(
		.INIT('h5501)
	) name181 (
		\sa20_reg[0]/P0001 ,
		_w695_,
		_w703_,
		_w713_,
		_w714_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w715_
	);
	LUT4 #(
		.INIT('h4000)
	) name183 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w716_
	);
	LUT2 #(
		.INIT('h2)
	) name184 (
		\sa20_reg[2]/P0001 ,
		_w716_,
		_w717_
	);
	LUT4 #(
		.INIT('h0002)
	) name185 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w718_
	);
	LUT3 #(
		.INIT('h02)
	) name186 (
		\sa20_reg[2]/P0001 ,
		_w716_,
		_w718_,
		_w719_
	);
	LUT4 #(
		.INIT('h0800)
	) name187 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w720_
	);
	LUT4 #(
		.INIT('h0020)
	) name188 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w721_
	);
	LUT4 #(
		.INIT('h0001)
	) name189 (
		\sa20_reg[2]/P0001 ,
		_w666_,
		_w721_,
		_w720_,
		_w722_
	);
	LUT4 #(
		.INIT('h1000)
	) name190 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w723_
	);
	LUT4 #(
		.INIT('h0800)
	) name191 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w724_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		_w723_,
		_w724_,
		_w725_
	);
	LUT4 #(
		.INIT('h0155)
	) name193 (
		\sa20_reg[1]/P0001 ,
		_w719_,
		_w722_,
		_w725_,
		_w726_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		\sa20_reg[1]/P0001 ,
		\sa20_reg[2]/P0001 ,
		_w727_
	);
	LUT3 #(
		.INIT('h20)
	) name195 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		_w728_
	);
	LUT3 #(
		.INIT('h02)
	) name196 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w729_
	);
	LUT4 #(
		.INIT('h0002)
	) name197 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w730_
	);
	LUT4 #(
		.INIT('h0001)
	) name198 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w731_
	);
	LUT4 #(
		.INIT('h0103)
	) name199 (
		_w643_,
		_w730_,
		_w731_,
		_w728_,
		_w732_
	);
	LUT2 #(
		.INIT('h2)
	) name200 (
		_w727_,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		_w666_,
		_w686_,
		_w734_
	);
	LUT2 #(
		.INIT('h2)
	) name202 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		_w735_
	);
	LUT3 #(
		.INIT('h01)
	) name203 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w736_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		\sa20_reg[7]/NET0131 ,
		_w711_,
		_w737_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name205 (
		\sa20_reg[7]/NET0131 ,
		_w711_,
		_w735_,
		_w736_,
		_w738_
	);
	LUT2 #(
		.INIT('h2)
	) name206 (
		\sa20_reg[1]/P0001 ,
		\sa20_reg[2]/P0001 ,
		_w739_
	);
	LUT3 #(
		.INIT('h02)
	) name207 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w740_
	);
	LUT3 #(
		.INIT('h80)
	) name208 (
		_w700_,
		_w739_,
		_w740_,
		_w741_
	);
	LUT3 #(
		.INIT('h80)
	) name209 (
		\sa20_reg[2]/P0001 ,
		_w647_,
		_w667_,
		_w742_
	);
	LUT4 #(
		.INIT('h0100)
	) name210 (
		_w741_,
		_w742_,
		_w734_,
		_w738_,
		_w743_
	);
	LUT3 #(
		.INIT('h10)
	) name211 (
		_w733_,
		_w726_,
		_w743_,
		_w744_
	);
	LUT3 #(
		.INIT('h10)
	) name212 (
		_w685_,
		_w714_,
		_w744_,
		_w745_
	);
	LUT2 #(
		.INIT('h9)
	) name213 (
		_w637_,
		_w745_,
		_w746_
	);
	LUT3 #(
		.INIT('h08)
	) name214 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w747_
	);
	LUT4 #(
		.INIT('h0040)
	) name215 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w748_
	);
	LUT2 #(
		.INIT('h4)
	) name216 (
		\sa13_reg[4]/P0001 ,
		_w748_,
		_w749_
	);
	LUT4 #(
		.INIT('h0002)
	) name217 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w750_
	);
	LUT4 #(
		.INIT('h1000)
	) name218 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w751_
	);
	LUT4 #(
		.INIT('h8000)
	) name219 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w752_
	);
	LUT4 #(
		.INIT('h0001)
	) name220 (
		_w539_,
		_w750_,
		_w751_,
		_w752_,
		_w753_
	);
	LUT4 #(
		.INIT('h0080)
	) name221 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w754_
	);
	LUT3 #(
		.INIT('ha8)
	) name222 (
		\sa13_reg[2]/P0001 ,
		_w544_,
		_w754_,
		_w755_
	);
	LUT4 #(
		.INIT('h0010)
	) name223 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w756_
	);
	LUT3 #(
		.INIT('h20)
	) name224 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w757_
	);
	LUT4 #(
		.INIT('h5554)
	) name225 (
		\sa13_reg[2]/P0001 ,
		_w566_,
		_w757_,
		_w756_,
		_w758_
	);
	LUT4 #(
		.INIT('h0100)
	) name226 (
		_w755_,
		_w749_,
		_w758_,
		_w753_,
		_w759_
	);
	LUT2 #(
		.INIT('h2)
	) name227 (
		\sa13_reg[1]/P0001 ,
		_w759_,
		_w760_
	);
	LUT3 #(
		.INIT('h08)
	) name228 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w761_
	);
	LUT4 #(
		.INIT('hc7f7)
	) name229 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w762_
	);
	LUT2 #(
		.INIT('h2)
	) name230 (
		_w576_,
		_w762_,
		_w763_
	);
	LUT4 #(
		.INIT('h0002)
	) name231 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w764_
	);
	LUT4 #(
		.INIT('h4000)
	) name232 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w765_
	);
	LUT3 #(
		.INIT('h54)
	) name233 (
		\sa13_reg[3]/P0001 ,
		_w764_,
		_w765_,
		_w766_
	);
	LUT3 #(
		.INIT('h54)
	) name234 (
		\sa13_reg[1]/P0001 ,
		_w763_,
		_w766_,
		_w767_
	);
	LUT4 #(
		.INIT('h0010)
	) name235 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w768_
	);
	LUT3 #(
		.INIT('h32)
	) name236 (
		_w584_,
		_w616_,
		_w768_,
		_w769_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w629_,
		_w752_,
		_w770_
	);
	LUT3 #(
		.INIT('h8a)
	) name238 (
		\sa13_reg[2]/P0001 ,
		_w769_,
		_w770_,
		_w771_
	);
	LUT3 #(
		.INIT('h23)
	) name239 (
		\sa13_reg[2]/P0001 ,
		_w577_,
		_w563_,
		_w772_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		_w560_,
		_w772_,
		_w773_
	);
	LUT3 #(
		.INIT('h10)
	) name241 (
		_w771_,
		_w767_,
		_w773_,
		_w774_
	);
	LUT3 #(
		.INIT('h45)
	) name242 (
		\sa13_reg[0]/P0001 ,
		_w760_,
		_w774_,
		_w775_
	);
	LUT4 #(
		.INIT('h0080)
	) name243 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w776_
	);
	LUT3 #(
		.INIT('h07)
	) name244 (
		\sa13_reg[4]/P0001 ,
		_w572_,
		_w776_,
		_w777_
	);
	LUT4 #(
		.INIT('hfd3f)
	) name245 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w778_
	);
	LUT3 #(
		.INIT('h10)
	) name246 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w779_
	);
	LUT4 #(
		.INIT('h0008)
	) name247 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w780_
	);
	LUT4 #(
		.INIT('h444e)
	) name248 (
		\sa13_reg[2]/P0001 ,
		_w778_,
		_w779_,
		_w780_,
		_w781_
	);
	LUT3 #(
		.INIT('h15)
	) name249 (
		\sa13_reg[1]/P0001 ,
		_w777_,
		_w781_,
		_w782_
	);
	LUT2 #(
		.INIT('h4)
	) name250 (
		\sa13_reg[3]/P0001 ,
		_w615_,
		_w783_
	);
	LUT3 #(
		.INIT('h04)
	) name251 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w784_
	);
	LUT2 #(
		.INIT('h8)
	) name252 (
		_w562_,
		_w784_,
		_w785_
	);
	LUT4 #(
		.INIT('h0200)
	) name253 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w786_
	);
	LUT3 #(
		.INIT('h07)
	) name254 (
		_w542_,
		_w543_,
		_w786_,
		_w787_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name255 (
		\sa13_reg[1]/P0001 ,
		_w783_,
		_w785_,
		_w787_,
		_w788_
	);
	LUT3 #(
		.INIT('h04)
	) name256 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w789_
	);
	LUT4 #(
		.INIT('h0020)
	) name257 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w790_
	);
	LUT4 #(
		.INIT('h5554)
	) name258 (
		\sa13_reg[2]/P0001 ,
		_w789_,
		_w776_,
		_w790_,
		_w791_
	);
	LUT4 #(
		.INIT('hfedc)
	) name259 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w792_
	);
	LUT3 #(
		.INIT('h8c)
	) name260 (
		_w614_,
		_w632_,
		_w792_,
		_w793_
	);
	LUT4 #(
		.INIT('h8000)
	) name261 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w794_
	);
	LUT4 #(
		.INIT('h0010)
	) name262 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w795_
	);
	LUT4 #(
		.INIT('h7fef)
	) name263 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w796_
	);
	LUT2 #(
		.INIT('h2)
	) name264 (
		_w583_,
		_w796_,
		_w797_
	);
	LUT4 #(
		.INIT('h2000)
	) name265 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w798_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name266 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w569_,
		_w798_,
		_w799_
	);
	LUT4 #(
		.INIT('h0100)
	) name267 (
		_w791_,
		_w797_,
		_w793_,
		_w799_,
		_w800_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name268 (
		\sa13_reg[0]/P0001 ,
		_w788_,
		_w782_,
		_w800_,
		_w801_
	);
	LUT3 #(
		.INIT('h14)
	) name269 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w802_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		_w565_,
		_w802_,
		_w803_
	);
	LUT3 #(
		.INIT('h08)
	) name271 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w804_
	);
	LUT4 #(
		.INIT('h0080)
	) name272 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w805_
	);
	LUT3 #(
		.INIT('h07)
	) name273 (
		\sa13_reg[4]/P0001 ,
		_w572_,
		_w805_,
		_w806_
	);
	LUT4 #(
		.INIT('h1311)
	) name274 (
		\sa13_reg[2]/P0001 ,
		_w617_,
		_w803_,
		_w806_,
		_w807_
	);
	LUT2 #(
		.INIT('h1)
	) name275 (
		\sa13_reg[1]/P0001 ,
		_w807_,
		_w808_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[2]/P0001 ,
		_w809_
	);
	LUT4 #(
		.INIT('h1000)
	) name277 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w810_
	);
	LUT4 #(
		.INIT('h0007)
	) name278 (
		_w535_,
		_w591_,
		_w798_,
		_w810_,
		_w811_
	);
	LUT2 #(
		.INIT('h2)
	) name279 (
		_w809_,
		_w811_,
		_w812_
	);
	LUT2 #(
		.INIT('h8)
	) name280 (
		_w583_,
		_w754_,
		_w813_
	);
	LUT3 #(
		.INIT('h02)
	) name281 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w814_
	);
	LUT4 #(
		.INIT('h23af)
	) name282 (
		\sa13_reg[2]/P0001 ,
		_w568_,
		_w563_,
		_w814_,
		_w815_
	);
	LUT3 #(
		.INIT('h8a)
	) name283 (
		\sa13_reg[1]/P0001 ,
		_w813_,
		_w815_,
		_w816_
	);
	LUT3 #(
		.INIT('h80)
	) name284 (
		\sa13_reg[4]/P0001 ,
		_w543_,
		_w594_,
		_w817_
	);
	LUT4 #(
		.INIT('h5540)
	) name285 (
		\sa13_reg[2]/P0001 ,
		_w543_,
		_w613_,
		_w751_,
		_w818_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		_w817_,
		_w818_,
		_w819_
	);
	LUT3 #(
		.INIT('h10)
	) name287 (
		_w816_,
		_w812_,
		_w819_,
		_w820_
	);
	LUT3 #(
		.INIT('h10)
	) name288 (
		_w801_,
		_w808_,
		_w820_,
		_w821_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w822_
	);
	LUT3 #(
		.INIT('h10)
	) name290 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w823_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w824_
	);
	LUT4 #(
		.INIT('h0008)
	) name292 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w825_
	);
	LUT3 #(
		.INIT('ha8)
	) name293 (
		\sa02_reg[2]/P0001 ,
		_w823_,
		_w825_,
		_w826_
	);
	LUT2 #(
		.INIT('h4)
	) name294 (
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w827_
	);
	LUT3 #(
		.INIT('h10)
	) name295 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w828_
	);
	LUT2 #(
		.INIT('h4)
	) name296 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		_w829_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		_w828_,
		_w829_,
		_w830_
	);
	LUT3 #(
		.INIT('h80)
	) name298 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w831_
	);
	LUT2 #(
		.INIT('h4)
	) name299 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w832_
	);
	LUT2 #(
		.INIT('h2)
	) name300 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		_w833_
	);
	LUT3 #(
		.INIT('h08)
	) name301 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w834_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name302 (
		_w831_,
		_w833_,
		_w832_,
		_w834_,
		_w835_
	);
	LUT4 #(
		.INIT('h5455)
	) name303 (
		\sa02_reg[1]/P0001 ,
		_w826_,
		_w830_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h2)
	) name304 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w837_
	);
	LUT3 #(
		.INIT('h20)
	) name305 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		_w838_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w839_
	);
	LUT3 #(
		.INIT('h01)
	) name307 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w840_
	);
	LUT2 #(
		.INIT('h2)
	) name308 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w841_
	);
	LUT4 #(
		.INIT('hfedc)
	) name309 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w842_
	);
	LUT3 #(
		.INIT('h8a)
	) name310 (
		\sa02_reg[1]/P0001 ,
		_w838_,
		_w842_,
		_w843_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w844_
	);
	LUT2 #(
		.INIT('h8)
	) name312 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w845_
	);
	LUT4 #(
		.INIT('h0020)
	) name313 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w846_
	);
	LUT2 #(
		.INIT('h2)
	) name314 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w847_
	);
	LUT4 #(
		.INIT('h0080)
	) name315 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w848_
	);
	LUT3 #(
		.INIT('h04)
	) name316 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w849_
	);
	LUT3 #(
		.INIT('h01)
	) name317 (
		_w846_,
		_w848_,
		_w849_,
		_w850_
	);
	LUT3 #(
		.INIT('h45)
	) name318 (
		\sa02_reg[2]/P0001 ,
		_w843_,
		_w850_,
		_w851_
	);
	LUT4 #(
		.INIT('h0080)
	) name319 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w852_
	);
	LUT4 #(
		.INIT('h0200)
	) name320 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w853_
	);
	LUT3 #(
		.INIT('h0b)
	) name321 (
		\sa02_reg[6]/NET0131 ,
		_w852_,
		_w853_,
		_w854_
	);
	LUT4 #(
		.INIT('h0004)
	) name322 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w855_
	);
	LUT2 #(
		.INIT('h8)
	) name323 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w856_
	);
	LUT2 #(
		.INIT('h2)
	) name324 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w857_
	);
	LUT3 #(
		.INIT('h04)
	) name325 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w858_
	);
	LUT4 #(
		.INIT('h47cf)
	) name326 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w855_,
		_w858_,
		_w859_
	);
	LUT3 #(
		.INIT('h2a)
	) name327 (
		\sa02_reg[1]/P0001 ,
		_w854_,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w861_
	);
	LUT4 #(
		.INIT('h0010)
	) name329 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w862_
	);
	LUT4 #(
		.INIT('haabf)
	) name330 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w831_,
		_w862_,
		_w863_
	);
	LUT4 #(
		.INIT('h2000)
	) name331 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w864_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name332 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		_w846_,
		_w864_,
		_w865_
	);
	LUT3 #(
		.INIT('hd0)
	) name333 (
		\sa02_reg[2]/P0001 ,
		_w863_,
		_w865_,
		_w866_
	);
	LUT4 #(
		.INIT('h0100)
	) name334 (
		_w860_,
		_w851_,
		_w836_,
		_w866_,
		_w867_
	);
	LUT4 #(
		.INIT('h0040)
	) name335 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w868_
	);
	LUT3 #(
		.INIT('h20)
	) name336 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w869_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w870_
	);
	LUT4 #(
		.INIT('hf5ef)
	) name338 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w871_
	);
	LUT3 #(
		.INIT('h10)
	) name339 (
		\sa02_reg[2]/P0001 ,
		_w868_,
		_w871_,
		_w872_
	);
	LUT4 #(
		.INIT('h0080)
	) name340 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w873_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w874_
	);
	LUT3 #(
		.INIT('h80)
	) name342 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w875_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name343 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w876_
	);
	LUT2 #(
		.INIT('h4)
	) name344 (
		_w873_,
		_w876_,
		_w877_
	);
	LUT3 #(
		.INIT('h80)
	) name345 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w878_
	);
	LUT4 #(
		.INIT('h77ef)
	) name346 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w879_
	);
	LUT3 #(
		.INIT('h20)
	) name347 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w880_
	);
	LUT4 #(
		.INIT('h0400)
	) name348 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w881_
	);
	LUT3 #(
		.INIT('h40)
	) name349 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w882_
	);
	LUT4 #(
		.INIT('h1000)
	) name350 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w883_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		_w884_
	);
	LUT4 #(
		.INIT('h0002)
	) name352 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w885_
	);
	LUT4 #(
		.INIT('heffd)
	) name353 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w886_
	);
	LUT4 #(
		.INIT('h0d00)
	) name354 (
		\sa02_reg[5]/P0001 ,
		_w879_,
		_w881_,
		_w886_,
		_w887_
	);
	LUT4 #(
		.INIT('h02aa)
	) name355 (
		\sa02_reg[1]/P0001 ,
		_w872_,
		_w877_,
		_w887_,
		_w888_
	);
	LUT3 #(
		.INIT('h01)
	) name356 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w889_
	);
	LUT4 #(
		.INIT('h0777)
	) name357 (
		_w870_,
		_w831_,
		_w833_,
		_w889_,
		_w890_
	);
	LUT2 #(
		.INIT('h8)
	) name358 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		_w891_
	);
	LUT4 #(
		.INIT('h153f)
	) name359 (
		\sa02_reg[7]/NET0131 ,
		_w840_,
		_w891_,
		_w855_,
		_w892_
	);
	LUT3 #(
		.INIT('h15)
	) name360 (
		\sa02_reg[1]/P0001 ,
		_w890_,
		_w892_,
		_w893_
	);
	LUT2 #(
		.INIT('h4)
	) name361 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w894_
	);
	LUT4 #(
		.INIT('h1000)
	) name362 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w895_
	);
	LUT4 #(
		.INIT('h0008)
	) name363 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w896_
	);
	LUT3 #(
		.INIT('h54)
	) name364 (
		\sa02_reg[2]/P0001 ,
		_w895_,
		_w896_,
		_w897_
	);
	LUT4 #(
		.INIT('h0400)
	) name365 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w898_
	);
	LUT3 #(
		.INIT('h20)
	) name366 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w898_,
		_w899_
	);
	LUT3 #(
		.INIT('h80)
	) name367 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w900_
	);
	LUT3 #(
		.INIT('h01)
	) name368 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w901_
	);
	LUT3 #(
		.INIT('h7e)
	) name369 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w902_
	);
	LUT2 #(
		.INIT('h2)
	) name370 (
		_w891_,
		_w902_,
		_w903_
	);
	LUT4 #(
		.INIT('h0800)
	) name371 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w904_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w905_
	);
	LUT3 #(
		.INIT('hf4)
	) name373 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w906_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name374 (
		\sa02_reg[2]/P0001 ,
		_w904_,
		_w844_,
		_w906_,
		_w907_
	);
	LUT4 #(
		.INIT('h0100)
	) name375 (
		_w903_,
		_w897_,
		_w899_,
		_w907_,
		_w908_
	);
	LUT3 #(
		.INIT('h10)
	) name376 (
		_w893_,
		_w888_,
		_w908_,
		_w909_
	);
	LUT3 #(
		.INIT('h10)
	) name377 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w910_
	);
	LUT4 #(
		.INIT('h0080)
	) name378 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w911_
	);
	LUT4 #(
		.INIT('hee7f)
	) name379 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w912_
	);
	LUT4 #(
		.INIT('h5054)
	) name380 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		_w864_,
		_w912_,
		_w913_
	);
	LUT4 #(
		.INIT('h0001)
	) name381 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w914_
	);
	LUT3 #(
		.INIT('h04)
	) name382 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w915_
	);
	LUT4 #(
		.INIT('h1445)
	) name383 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w916_
	);
	LUT2 #(
		.INIT('h8)
	) name384 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w917_
	);
	LUT3 #(
		.INIT('ha2)
	) name385 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w918_
	);
	LUT4 #(
		.INIT('h5551)
	) name386 (
		_w914_,
		_w917_,
		_w918_,
		_w916_,
		_w919_
	);
	LUT3 #(
		.INIT('h45)
	) name387 (
		\sa02_reg[1]/P0001 ,
		_w913_,
		_w919_,
		_w920_
	);
	LUT3 #(
		.INIT('h8a)
	) name388 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w852_,
		_w921_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		\sa02_reg[2]/P0001 ,
		_w883_,
		_w922_
	);
	LUT3 #(
		.INIT('h02)
	) name390 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w923_
	);
	LUT2 #(
		.INIT('h8)
	) name391 (
		_w847_,
		_w923_,
		_w924_
	);
	LUT4 #(
		.INIT('h0111)
	) name392 (
		\sa02_reg[2]/P0001 ,
		_w883_,
		_w847_,
		_w923_,
		_w925_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		_w921_,
		_w925_,
		_w926_
	);
	LUT4 #(
		.INIT('h0020)
	) name394 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w927_
	);
	LUT3 #(
		.INIT('h80)
	) name395 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		_w927_,
		_w928_
	);
	LUT4 #(
		.INIT('h0002)
	) name396 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w929_
	);
	LUT4 #(
		.INIT('h8caf)
	) name397 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		_w904_,
		_w929_,
		_w930_
	);
	LUT3 #(
		.INIT('h8a)
	) name398 (
		\sa02_reg[1]/P0001 ,
		_w928_,
		_w930_,
		_w931_
	);
	LUT3 #(
		.INIT('h01)
	) name399 (
		_w926_,
		_w931_,
		_w920_,
		_w932_
	);
	LUT4 #(
		.INIT('he400)
	) name400 (
		\sa02_reg[0]/P0001 ,
		_w909_,
		_w867_,
		_w932_,
		_w933_
	);
	LUT2 #(
		.INIT('h4)
	) name401 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w934_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w935_
	);
	LUT3 #(
		.INIT('h10)
	) name403 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w936_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w937_
	);
	LUT3 #(
		.INIT('h20)
	) name405 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w938_
	);
	LUT4 #(
		.INIT('h0400)
	) name406 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w939_
	);
	LUT2 #(
		.INIT('h2)
	) name407 (
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w940_
	);
	LUT3 #(
		.INIT('h08)
	) name408 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w941_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name409 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w942_
	);
	LUT4 #(
		.INIT('h80aa)
	) name410 (
		\sa31_reg[2]/P0001 ,
		_w934_,
		_w936_,
		_w942_,
		_w943_
	);
	LUT2 #(
		.INIT('h8)
	) name411 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w944_
	);
	LUT3 #(
		.INIT('h80)
	) name412 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w945_
	);
	LUT4 #(
		.INIT('h2000)
	) name413 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w946_
	);
	LUT2 #(
		.INIT('h2)
	) name414 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w947_
	);
	LUT3 #(
		.INIT('h08)
	) name415 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w948_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		_w949_
	);
	LUT3 #(
		.INIT('h23)
	) name417 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w950_
	);
	LUT4 #(
		.INIT('h0777)
	) name418 (
		_w947_,
		_w948_,
		_w949_,
		_w950_,
		_w951_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name419 (
		\sa31_reg[1]/P0001 ,
		_w943_,
		_w946_,
		_w951_,
		_w952_
	);
	LUT4 #(
		.INIT('h0008)
	) name420 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w953_
	);
	LUT2 #(
		.INIT('h4)
	) name421 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w954_
	);
	LUT4 #(
		.INIT('h1000)
	) name422 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w955_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		_w953_,
		_w955_,
		_w956_
	);
	LUT3 #(
		.INIT('h54)
	) name424 (
		\sa31_reg[2]/P0001 ,
		_w953_,
		_w955_,
		_w957_
	);
	LUT3 #(
		.INIT('h04)
	) name425 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w958_
	);
	LUT3 #(
		.INIT('h80)
	) name426 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w959_
	);
	LUT3 #(
		.INIT('ha8)
	) name427 (
		\sa31_reg[2]/P0001 ,
		_w958_,
		_w959_,
		_w960_
	);
	LUT2 #(
		.INIT('h2)
	) name428 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w961_
	);
	LUT4 #(
		.INIT('h0800)
	) name429 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w962_
	);
	LUT2 #(
		.INIT('h1)
	) name430 (
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w963_
	);
	LUT3 #(
		.INIT('h02)
	) name431 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w964_
	);
	LUT3 #(
		.INIT('h13)
	) name432 (
		_w949_,
		_w962_,
		_w964_,
		_w965_
	);
	LUT4 #(
		.INIT('h5455)
	) name433 (
		\sa31_reg[1]/P0001 ,
		_w960_,
		_w957_,
		_w965_,
		_w966_
	);
	LUT3 #(
		.INIT('h08)
	) name434 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w967_
	);
	LUT4 #(
		.INIT('h0040)
	) name435 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w968_
	);
	LUT2 #(
		.INIT('h4)
	) name436 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w969_
	);
	LUT4 #(
		.INIT('h0040)
	) name437 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w970_
	);
	LUT3 #(
		.INIT('h54)
	) name438 (
		\sa31_reg[2]/P0001 ,
		_w968_,
		_w970_,
		_w971_
	);
	LUT4 #(
		.INIT('h0080)
	) name439 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w972_
	);
	LUT3 #(
		.INIT('h80)
	) name440 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w973_
	);
	LUT3 #(
		.INIT('h13)
	) name441 (
		_w969_,
		_w972_,
		_w973_,
		_w974_
	);
	LUT3 #(
		.INIT('h01)
	) name442 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w975_
	);
	LUT4 #(
		.INIT('h0001)
	) name443 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w976_
	);
	LUT4 #(
		.INIT('h0200)
	) name444 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w977_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		_w976_,
		_w977_,
		_w978_
	);
	LUT4 #(
		.INIT('h3111)
	) name446 (
		\sa31_reg[2]/P0001 ,
		_w971_,
		_w974_,
		_w978_,
		_w979_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name447 (
		\sa31_reg[0]/P0002 ,
		_w952_,
		_w966_,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		_w981_
	);
	LUT4 #(
		.INIT('h4000)
	) name449 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w982_
	);
	LUT4 #(
		.INIT('h0105)
	) name450 (
		\sa31_reg[1]/P0001 ,
		_w964_,
		_w982_,
		_w981_,
		_w983_
	);
	LUT2 #(
		.INIT('h2)
	) name451 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w984_
	);
	LUT3 #(
		.INIT('h40)
	) name452 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w985_
	);
	LUT3 #(
		.INIT('h9d)
	) name453 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w986_
	);
	LUT3 #(
		.INIT('h10)
	) name454 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w987_
	);
	LUT4 #(
		.INIT('hfa3f)
	) name455 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w988_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name456 (
		\sa31_reg[4]/P0001 ,
		_w954_,
		_w986_,
		_w988_,
		_w989_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		_w983_,
		_w989_,
		_w990_
	);
	LUT2 #(
		.INIT('h4)
	) name458 (
		\sa31_reg[2]/P0001 ,
		_w976_,
		_w991_
	);
	LUT2 #(
		.INIT('h2)
	) name459 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		_w992_
	);
	LUT3 #(
		.INIT('h80)
	) name460 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w993_
	);
	LUT3 #(
		.INIT('h7e)
	) name461 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w994_
	);
	LUT2 #(
		.INIT('h2)
	) name462 (
		_w992_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h2)
	) name463 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w996_
	);
	LUT3 #(
		.INIT('h80)
	) name464 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w997_
	);
	LUT3 #(
		.INIT('h2a)
	) name465 (
		\sa31_reg[1]/P0001 ,
		_w996_,
		_w997_,
		_w998_
	);
	LUT3 #(
		.INIT('h10)
	) name466 (
		_w995_,
		_w991_,
		_w998_,
		_w999_
	);
	LUT2 #(
		.INIT('h8)
	) name467 (
		_w947_,
		_w985_,
		_w1000_
	);
	LUT2 #(
		.INIT('h1)
	) name468 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w1001_
	);
	LUT4 #(
		.INIT('h0004)
	) name469 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w1002_
	);
	LUT2 #(
		.INIT('h8)
	) name470 (
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w1003_
	);
	LUT3 #(
		.INIT('h2a)
	) name471 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w1004_
	);
	LUT4 #(
		.INIT('h2220)
	) name472 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w1005_
	);
	LUT3 #(
		.INIT('h45)
	) name473 (
		_w1002_,
		_w1004_,
		_w1005_,
		_w1006_
	);
	LUT3 #(
		.INIT('h20)
	) name474 (
		_w950_,
		_w1004_,
		_w992_,
		_w1007_
	);
	LUT4 #(
		.INIT('h00ba)
	) name475 (
		\sa31_reg[2]/P0001 ,
		_w1000_,
		_w1006_,
		_w1007_,
		_w1008_
	);
	LUT4 #(
		.INIT('h0155)
	) name476 (
		\sa31_reg[0]/P0002 ,
		_w990_,
		_w999_,
		_w1008_,
		_w1009_
	);
	LUT4 #(
		.INIT('h0800)
	) name477 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w1010_
	);
	LUT4 #(
		.INIT('h0020)
	) name478 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w1011_
	);
	LUT4 #(
		.INIT('hf7df)
	) name479 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w1012_
	);
	LUT3 #(
		.INIT('h45)
	) name480 (
		\sa31_reg[2]/P0001 ,
		_w1010_,
		_w1012_,
		_w1013_
	);
	LUT2 #(
		.INIT('h2)
	) name481 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w1014_
	);
	LUT3 #(
		.INIT('h08)
	) name482 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w1015_
	);
	LUT2 #(
		.INIT('h8)
	) name483 (
		_w963_,
		_w1015_,
		_w1016_
	);
	LUT4 #(
		.INIT('h0800)
	) name484 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w1017_
	);
	LUT4 #(
		.INIT('h1000)
	) name485 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w1018_
	);
	LUT4 #(
		.INIT('h0007)
	) name486 (
		_w973_,
		_w1014_,
		_w1017_,
		_w1018_,
		_w1019_
	);
	LUT4 #(
		.INIT('h5455)
	) name487 (
		\sa31_reg[1]/P0001 ,
		_w1013_,
		_w1016_,
		_w1019_,
		_w1020_
	);
	LUT2 #(
		.INIT('h8)
	) name488 (
		\sa31_reg[1]/P0001 ,
		\sa31_reg[2]/P0001 ,
		_w1021_
	);
	LUT4 #(
		.INIT('h0002)
	) name489 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w1022_
	);
	LUT4 #(
		.INIT('h0001)
	) name490 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w1023_
	);
	LUT4 #(
		.INIT('h0007)
	) name491 (
		\sa31_reg[3]/P0001 ,
		_w939_,
		_w1022_,
		_w1023_,
		_w1024_
	);
	LUT2 #(
		.INIT('h2)
	) name492 (
		_w1021_,
		_w1024_,
		_w1025_
	);
	LUT4 #(
		.INIT('h0001)
	) name493 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w1026_
	);
	LUT2 #(
		.INIT('h8)
	) name494 (
		\sa31_reg[2]/P0001 ,
		_w1026_,
		_w1027_
	);
	LUT2 #(
		.INIT('h8)
	) name495 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w1028_
	);
	LUT4 #(
		.INIT('h0020)
	) name496 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w1029_
	);
	LUT3 #(
		.INIT('h01)
	) name497 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w1030_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		_w1001_,
		_w1030_,
		_w1031_
	);
	LUT4 #(
		.INIT('h0777)
	) name499 (
		_w1028_,
		_w1029_,
		_w1001_,
		_w1030_,
		_w1032_
	);
	LUT2 #(
		.INIT('h8)
	) name500 (
		_w961_,
		_w982_,
		_w1033_
	);
	LUT2 #(
		.INIT('h2)
	) name501 (
		\sa31_reg[1]/P0001 ,
		\sa31_reg[2]/P0001 ,
		_w1034_
	);
	LUT3 #(
		.INIT('h02)
	) name502 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w1035_
	);
	LUT3 #(
		.INIT('h80)
	) name503 (
		_w947_,
		_w1034_,
		_w1035_,
		_w1036_
	);
	LUT4 #(
		.INIT('h0100)
	) name504 (
		_w1027_,
		_w1033_,
		_w1036_,
		_w1032_,
		_w1037_
	);
	LUT3 #(
		.INIT('h10)
	) name505 (
		_w1025_,
		_w1020_,
		_w1037_,
		_w1038_
	);
	LUT3 #(
		.INIT('h10)
	) name506 (
		_w980_,
		_w1009_,
		_w1038_,
		_w1039_
	);
	LUT4 #(
		.INIT('h5655)
	) name507 (
		\u0_w_reg[2][30]/P0001 ,
		_w980_,
		_w1009_,
		_w1038_,
		_w1040_
	);
	LUT4 #(
		.INIT('h4bb4)
	) name508 (
		_w775_,
		_w821_,
		_w933_,
		_w1040_,
		_w1041_
	);
	LUT3 #(
		.INIT('h82)
	) name509 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[62]/P0001 ,
		\u0_w_reg[2][30]/P0001 ,
		_w1042_
	);
	LUT4 #(
		.INIT('h00eb)
	) name510 (
		\ld_r_reg/P0001 ,
		_w746_,
		_w1041_,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('h2)
	) name511 (
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1044_
	);
	LUT3 #(
		.INIT('h08)
	) name512 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1045_
	);
	LUT4 #(
		.INIT('h0080)
	) name513 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1046_
	);
	LUT2 #(
		.INIT('h1)
	) name514 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1047_
	);
	LUT4 #(
		.INIT('h0020)
	) name515 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1048_
	);
	LUT4 #(
		.INIT('h2000)
	) name516 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1049_
	);
	LUT2 #(
		.INIT('h2)
	) name517 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1050_
	);
	LUT4 #(
		.INIT('hdfbb)
	) name518 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1051_
	);
	LUT4 #(
		.INIT('h5455)
	) name519 (
		\sa03_reg[2]/P0001 ,
		_w1046_,
		_w1048_,
		_w1051_,
		_w1052_
	);
	LUT2 #(
		.INIT('h4)
	) name520 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1053_
	);
	LUT3 #(
		.INIT('h80)
	) name521 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1054_
	);
	LUT2 #(
		.INIT('h8)
	) name522 (
		_w1053_,
		_w1054_,
		_w1055_
	);
	LUT4 #(
		.INIT('h0010)
	) name523 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1056_
	);
	LUT2 #(
		.INIT('h4)
	) name524 (
		\sa03_reg[5]/P0001 ,
		_w1056_,
		_w1057_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name525 (
		\sa03_reg[5]/P0001 ,
		_w1056_,
		_w1053_,
		_w1054_,
		_w1058_
	);
	LUT2 #(
		.INIT('h2)
	) name526 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1059_
	);
	LUT3 #(
		.INIT('h20)
	) name527 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		_w1060_
	);
	LUT2 #(
		.INIT('h8)
	) name528 (
		_w1044_,
		_w1060_,
		_w1061_
	);
	LUT4 #(
		.INIT('h000d)
	) name529 (
		\sa03_reg[2]/P0001 ,
		_w1058_,
		_w1052_,
		_w1061_,
		_w1062_
	);
	LUT3 #(
		.INIT('h10)
	) name530 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1063_
	);
	LUT2 #(
		.INIT('h8)
	) name531 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1064_
	);
	LUT4 #(
		.INIT('h0008)
	) name532 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1065_
	);
	LUT3 #(
		.INIT('ha8)
	) name533 (
		\sa03_reg[2]/P0001 ,
		_w1063_,
		_w1065_,
		_w1066_
	);
	LUT3 #(
		.INIT('h10)
	) name534 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1067_
	);
	LUT2 #(
		.INIT('h4)
	) name535 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1068_
	);
	LUT2 #(
		.INIT('h2)
	) name536 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1069_
	);
	LUT4 #(
		.INIT('h22bf)
	) name537 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1067_,
		_w1045_,
		_w1070_
	);
	LUT4 #(
		.INIT('h5455)
	) name538 (
		\sa03_reg[1]/P0001 ,
		_w1066_,
		_w1055_,
		_w1070_,
		_w1071_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1072_
	);
	LUT3 #(
		.INIT('h01)
	) name540 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1073_
	);
	LUT2 #(
		.INIT('h2)
	) name541 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1074_
	);
	LUT4 #(
		.INIT('hdfd3)
	) name542 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1075_
	);
	LUT3 #(
		.INIT('h45)
	) name543 (
		\sa03_reg[2]/P0001 ,
		_w1073_,
		_w1075_,
		_w1076_
	);
	LUT4 #(
		.INIT('h0200)
	) name544 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1077_
	);
	LUT3 #(
		.INIT('h07)
	) name545 (
		\sa03_reg[5]/P0001 ,
		_w1065_,
		_w1077_,
		_w1078_
	);
	LUT3 #(
		.INIT('h01)
	) name546 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1079_
	);
	LUT2 #(
		.INIT('h8)
	) name547 (
		_w1053_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h8)
	) name548 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1081_
	);
	LUT3 #(
		.INIT('h80)
	) name549 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1082_
	);
	LUT2 #(
		.INIT('h1)
	) name550 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1083_
	);
	LUT4 #(
		.INIT('h153f)
	) name551 (
		_w1053_,
		_w1082_,
		_w1083_,
		_w1079_,
		_w1084_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name552 (
		\sa03_reg[1]/P0001 ,
		_w1076_,
		_w1078_,
		_w1084_,
		_w1085_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name553 (
		\sa03_reg[0]/P0001 ,
		_w1071_,
		_w1085_,
		_w1062_,
		_w1086_
	);
	LUT4 #(
		.INIT('h0040)
	) name554 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1087_
	);
	LUT4 #(
		.INIT('h5155)
	) name555 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1088_
	);
	LUT3 #(
		.INIT('h10)
	) name556 (
		_w1056_,
		_w1087_,
		_w1088_,
		_w1089_
	);
	LUT4 #(
		.INIT('h0080)
	) name557 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1090_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name558 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1091_
	);
	LUT2 #(
		.INIT('h4)
	) name559 (
		_w1090_,
		_w1091_,
		_w1092_
	);
	LUT3 #(
		.INIT('h80)
	) name560 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1093_
	);
	LUT4 #(
		.INIT('h77ef)
	) name561 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1094_
	);
	LUT2 #(
		.INIT('h4)
	) name562 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1095_
	);
	LUT4 #(
		.INIT('h0400)
	) name563 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1096_
	);
	LUT4 #(
		.INIT('h0002)
	) name564 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1097_
	);
	LUT2 #(
		.INIT('h4)
	) name565 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1098_
	);
	LUT4 #(
		.INIT('h1000)
	) name566 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1099_
	);
	LUT4 #(
		.INIT('heffd)
	) name567 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1100_
	);
	LUT4 #(
		.INIT('h0d00)
	) name568 (
		\sa03_reg[5]/P0001 ,
		_w1094_,
		_w1096_,
		_w1100_,
		_w1101_
	);
	LUT4 #(
		.INIT('h02aa)
	) name569 (
		\sa03_reg[1]/P0001 ,
		_w1089_,
		_w1092_,
		_w1101_,
		_w1102_
	);
	LUT4 #(
		.INIT('h0100)
	) name570 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1103_
	);
	LUT2 #(
		.INIT('h8)
	) name571 (
		\sa03_reg[4]/P0001 ,
		_w1103_,
		_w1104_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1105_
	);
	LUT3 #(
		.INIT('h2a)
	) name573 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1106_
	);
	LUT4 #(
		.INIT('h0203)
	) name574 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1107_
	);
	LUT4 #(
		.INIT('h0777)
	) name575 (
		_w1105_,
		_w1054_,
		_w1106_,
		_w1107_,
		_w1108_
	);
	LUT3 #(
		.INIT('h45)
	) name576 (
		\sa03_reg[1]/P0001 ,
		_w1104_,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1110_
	);
	LUT2 #(
		.INIT('h4)
	) name578 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1111_
	);
	LUT4 #(
		.INIT('h1000)
	) name579 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1112_
	);
	LUT4 #(
		.INIT('h0008)
	) name580 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1113_
	);
	LUT3 #(
		.INIT('h54)
	) name581 (
		\sa03_reg[2]/P0001 ,
		_w1112_,
		_w1113_,
		_w1114_
	);
	LUT2 #(
		.INIT('h8)
	) name582 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1115_
	);
	LUT2 #(
		.INIT('h1)
	) name583 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1116_
	);
	LUT3 #(
		.INIT('h01)
	) name584 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1117_
	);
	LUT3 #(
		.INIT('h7e)
	) name585 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1118_
	);
	LUT2 #(
		.INIT('h2)
	) name586 (
		_w1115_,
		_w1118_,
		_w1119_
	);
	LUT3 #(
		.INIT('h08)
	) name587 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1120_
	);
	LUT4 #(
		.INIT('h0800)
	) name588 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1121_
	);
	LUT2 #(
		.INIT('h4)
	) name589 (
		\sa03_reg[2]/P0001 ,
		_w1121_,
		_w1122_
	);
	LUT3 #(
		.INIT('h04)
	) name590 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1123_
	);
	LUT3 #(
		.INIT('h20)
	) name591 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1124_
	);
	LUT2 #(
		.INIT('h2)
	) name592 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1125_
	);
	LUT3 #(
		.INIT('hf4)
	) name593 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1126_
	);
	LUT4 #(
		.INIT('h7707)
	) name594 (
		_w1123_,
		_w1124_,
		_w1047_,
		_w1126_,
		_w1127_
	);
	LUT4 #(
		.INIT('h0100)
	) name595 (
		_w1122_,
		_w1114_,
		_w1119_,
		_w1127_,
		_w1128_
	);
	LUT4 #(
		.INIT('h5455)
	) name596 (
		\sa03_reg[0]/P0001 ,
		_w1102_,
		_w1109_,
		_w1128_,
		_w1129_
	);
	LUT4 #(
		.INIT('h0080)
	) name597 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1130_
	);
	LUT4 #(
		.INIT('h1000)
	) name598 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1131_
	);
	LUT4 #(
		.INIT('h0103)
	) name599 (
		\sa03_reg[5]/P0001 ,
		_w1131_,
		_w1049_,
		_w1130_,
		_w1132_
	);
	LUT3 #(
		.INIT('h6b)
	) name600 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1133_
	);
	LUT2 #(
		.INIT('h2)
	) name601 (
		_w1124_,
		_w1133_,
		_w1134_
	);
	LUT4 #(
		.INIT('h0001)
	) name602 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1135_
	);
	LUT3 #(
		.INIT('h07)
	) name603 (
		_w1120_,
		_w1115_,
		_w1135_,
		_w1136_
	);
	LUT4 #(
		.INIT('h0e00)
	) name604 (
		\sa03_reg[2]/P0001 ,
		_w1132_,
		_w1134_,
		_w1136_,
		_w1137_
	);
	LUT4 #(
		.INIT('h4000)
	) name605 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1138_
	);
	LUT3 #(
		.INIT('h20)
	) name606 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1138_,
		_w1139_
	);
	LUT3 #(
		.INIT('h02)
	) name607 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1140_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name608 (
		\sa03_reg[2]/P0001 ,
		_w1121_,
		_w1116_,
		_w1140_,
		_w1141_
	);
	LUT2 #(
		.INIT('h4)
	) name609 (
		_w1139_,
		_w1141_,
		_w1142_
	);
	LUT4 #(
		.INIT('h0008)
	) name610 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1143_
	);
	LUT2 #(
		.INIT('h8)
	) name611 (
		_w1115_,
		_w1143_,
		_w1144_
	);
	LUT4 #(
		.INIT('h0004)
	) name612 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1145_
	);
	LUT4 #(
		.INIT('h5450)
	) name613 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1099_,
		_w1145_,
		_w1146_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		_w1144_,
		_w1146_,
		_w1147_
	);
	LUT4 #(
		.INIT('he400)
	) name615 (
		\sa03_reg[1]/P0001 ,
		_w1137_,
		_w1142_,
		_w1147_,
		_w1148_
	);
	LUT3 #(
		.INIT('h10)
	) name616 (
		_w1129_,
		_w1086_,
		_w1148_,
		_w1149_
	);
	LUT4 #(
		.INIT('h0004)
	) name617 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1150_
	);
	LUT3 #(
		.INIT('h23)
	) name618 (
		\sa03_reg[2]/P0001 ,
		_w1121_,
		_w1150_,
		_w1151_
	);
	LUT3 #(
		.INIT('h45)
	) name619 (
		\sa03_reg[1]/P0001 ,
		_w1114_,
		_w1151_,
		_w1152_
	);
	LUT4 #(
		.INIT('h2000)
	) name620 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1153_
	);
	LUT3 #(
		.INIT('h07)
	) name621 (
		\sa03_reg[5]/P0001 ,
		_w1065_,
		_w1153_,
		_w1154_
	);
	LUT3 #(
		.INIT('h08)
	) name622 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1155_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name623 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1156_
	);
	LUT4 #(
		.INIT('h20aa)
	) name624 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1099_,
		_w1156_,
		_w1157_
	);
	LUT3 #(
		.INIT('ha2)
	) name625 (
		\sa03_reg[1]/P0001 ,
		_w1154_,
		_w1157_,
		_w1158_
	);
	LUT4 #(
		.INIT('h0001)
	) name626 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1159_
	);
	LUT4 #(
		.INIT('h0007)
	) name627 (
		_w1053_,
		_w1054_,
		_w1130_,
		_w1159_,
		_w1160_
	);
	LUT2 #(
		.INIT('h2)
	) name628 (
		\sa03_reg[2]/P0001 ,
		_w1160_,
		_w1161_
	);
	LUT3 #(
		.INIT('h02)
	) name629 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		_w1162_
	);
	LUT4 #(
		.INIT('h0040)
	) name630 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1163_
	);
	LUT4 #(
		.INIT('h0405)
	) name631 (
		_w1087_,
		_w1111_,
		_w1163_,
		_w1162_,
		_w1164_
	);
	LUT2 #(
		.INIT('h4)
	) name632 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[2]/P0001 ,
		_w1165_
	);
	LUT3 #(
		.INIT('he0)
	) name633 (
		_w1093_,
		_w1123_,
		_w1165_,
		_w1166_
	);
	LUT2 #(
		.INIT('h8)
	) name634 (
		_w1115_,
		_w1067_,
		_w1167_
	);
	LUT4 #(
		.INIT('h0302)
	) name635 (
		\sa03_reg[2]/P0001 ,
		_w1166_,
		_w1167_,
		_w1164_,
		_w1168_
	);
	LUT4 #(
		.INIT('h0100)
	) name636 (
		_w1158_,
		_w1161_,
		_w1152_,
		_w1168_,
		_w1169_
	);
	LUT2 #(
		.INIT('h4)
	) name637 (
		_w1118_,
		_w1069_,
		_w1170_
	);
	LUT2 #(
		.INIT('h1)
	) name638 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1171_
	);
	LUT2 #(
		.INIT('h8)
	) name639 (
		_w1079_,
		_w1171_,
		_w1172_
	);
	LUT3 #(
		.INIT('h2a)
	) name640 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[5]/P0001 ,
		_w1130_,
		_w1173_
	);
	LUT3 #(
		.INIT('h10)
	) name641 (
		_w1172_,
		_w1170_,
		_w1173_,
		_w1174_
	);
	LUT3 #(
		.INIT('h08)
	) name642 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1175_
	);
	LUT4 #(
		.INIT('h0105)
	) name643 (
		\sa03_reg[1]/P0001 ,
		_w1050_,
		_w1163_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h8)
	) name644 (
		\sa03_reg[4]/P0001 ,
		_w1099_,
		_w1177_
	);
	LUT4 #(
		.INIT('h4000)
	) name645 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1178_
	);
	LUT3 #(
		.INIT('hd8)
	) name646 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1179_
	);
	LUT3 #(
		.INIT('h31)
	) name647 (
		_w1095_,
		_w1178_,
		_w1179_,
		_w1180_
	);
	LUT3 #(
		.INIT('h40)
	) name648 (
		_w1177_,
		_w1176_,
		_w1180_,
		_w1181_
	);
	LUT3 #(
		.INIT('h02)
	) name649 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1182_
	);
	LUT4 #(
		.INIT('h2220)
	) name650 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1183_
	);
	LUT3 #(
		.INIT('h54)
	) name651 (
		_w1064_,
		_w1182_,
		_w1183_,
		_w1184_
	);
	LUT4 #(
		.INIT('h2000)
	) name652 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1185_
	);
	LUT4 #(
		.INIT('h0045)
	) name653 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1138_,
		_w1185_,
		_w1186_
	);
	LUT4 #(
		.INIT('h0001)
	) name654 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1187_
	);
	LUT4 #(
		.INIT('h002a)
	) name655 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1099_,
		_w1187_,
		_w1188_
	);
	LUT3 #(
		.INIT('h0b)
	) name656 (
		_w1184_,
		_w1186_,
		_w1188_,
		_w1189_
	);
	LUT3 #(
		.INIT('h0e)
	) name657 (
		_w1174_,
		_w1181_,
		_w1189_,
		_w1190_
	);
	LUT4 #(
		.INIT('h4000)
	) name658 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1191_
	);
	LUT2 #(
		.INIT('h2)
	) name659 (
		\sa03_reg[2]/P0001 ,
		_w1191_,
		_w1192_
	);
	LUT4 #(
		.INIT('h0002)
	) name660 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1193_
	);
	LUT3 #(
		.INIT('h02)
	) name661 (
		\sa03_reg[2]/P0001 ,
		_w1191_,
		_w1193_,
		_w1194_
	);
	LUT4 #(
		.INIT('h0800)
	) name662 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1195_
	);
	LUT4 #(
		.INIT('h0020)
	) name663 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1196_
	);
	LUT4 #(
		.INIT('h0001)
	) name664 (
		\sa03_reg[2]/P0001 ,
		_w1121_,
		_w1195_,
		_w1196_,
		_w1197_
	);
	LUT4 #(
		.INIT('h1000)
	) name665 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1198_
	);
	LUT4 #(
		.INIT('h0800)
	) name666 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1199_
	);
	LUT2 #(
		.INIT('h1)
	) name667 (
		_w1198_,
		_w1199_,
		_w1200_
	);
	LUT4 #(
		.INIT('h0155)
	) name668 (
		\sa03_reg[1]/P0001 ,
		_w1194_,
		_w1197_,
		_w1200_,
		_w1201_
	);
	LUT4 #(
		.INIT('h0002)
	) name669 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1202_
	);
	LUT4 #(
		.INIT('h0023)
	) name670 (
		\sa03_reg[6]/NET0131 ,
		_w1135_,
		_w1153_,
		_w1202_,
		_w1203_
	);
	LUT2 #(
		.INIT('h8)
	) name671 (
		_w1064_,
		_w1123_,
		_w1204_
	);
	LUT4 #(
		.INIT('hcc08)
	) name672 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[2]/P0001 ,
		_w1203_,
		_w1204_,
		_w1205_
	);
	LUT2 #(
		.INIT('h8)
	) name673 (
		_w1121_,
		_w1068_,
		_w1206_
	);
	LUT2 #(
		.INIT('h4)
	) name674 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1207_
	);
	LUT4 #(
		.INIT('h0001)
	) name675 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1208_
	);
	LUT2 #(
		.INIT('h4)
	) name676 (
		_w1207_,
		_w1208_,
		_w1209_
	);
	LUT2 #(
		.INIT('h2)
	) name677 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[2]/P0001 ,
		_w1210_
	);
	LUT3 #(
		.INIT('h80)
	) name678 (
		\sa03_reg[3]/P0001 ,
		_w1145_,
		_w1210_,
		_w1211_
	);
	LUT3 #(
		.INIT('h01)
	) name679 (
		_w1209_,
		_w1211_,
		_w1206_,
		_w1212_
	);
	LUT3 #(
		.INIT('h10)
	) name680 (
		_w1205_,
		_w1201_,
		_w1212_,
		_w1213_
	);
	LUT4 #(
		.INIT('hd800)
	) name681 (
		\sa03_reg[0]/P0001 ,
		_w1169_,
		_w1190_,
		_w1213_,
		_w1214_
	);
	LUT2 #(
		.INIT('h4)
	) name682 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1215_
	);
	LUT2 #(
		.INIT('h4)
	) name683 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1216_
	);
	LUT4 #(
		.INIT('h1000)
	) name684 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1217_
	);
	LUT3 #(
		.INIT('h08)
	) name685 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1218_
	);
	LUT2 #(
		.INIT('h2)
	) name686 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1219_
	);
	LUT4 #(
		.INIT('h0400)
	) name687 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1220_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name688 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1221_
	);
	LUT4 #(
		.INIT('h20aa)
	) name689 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		_w1217_,
		_w1221_,
		_w1222_
	);
	LUT2 #(
		.INIT('h8)
	) name690 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1223_
	);
	LUT2 #(
		.INIT('h2)
	) name691 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1224_
	);
	LUT4 #(
		.INIT('h2000)
	) name692 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1225_
	);
	LUT2 #(
		.INIT('h2)
	) name693 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1226_
	);
	LUT2 #(
		.INIT('h8)
	) name694 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1227_
	);
	LUT3 #(
		.INIT('h08)
	) name695 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1228_
	);
	LUT3 #(
		.INIT('h15)
	) name696 (
		_w1225_,
		_w1226_,
		_w1228_,
		_w1229_
	);
	LUT2 #(
		.INIT('h1)
	) name697 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		_w1230_
	);
	LUT3 #(
		.INIT('h23)
	) name698 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1231_
	);
	LUT2 #(
		.INIT('h8)
	) name699 (
		_w1230_,
		_w1231_,
		_w1232_
	);
	LUT4 #(
		.INIT('haaa2)
	) name700 (
		\sa10_reg[1]/P0001 ,
		_w1229_,
		_w1232_,
		_w1222_,
		_w1233_
	);
	LUT2 #(
		.INIT('h1)
	) name701 (
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1234_
	);
	LUT3 #(
		.INIT('h02)
	) name702 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1235_
	);
	LUT4 #(
		.INIT('h0004)
	) name703 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1236_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		\sa10_reg[2]/P0001 ,
		_w1236_,
		_w1237_
	);
	LUT3 #(
		.INIT('h80)
	) name705 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1238_
	);
	LUT3 #(
		.INIT('h04)
	) name706 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1239_
	);
	LUT4 #(
		.INIT('heee4)
	) name707 (
		\sa10_reg[2]/P0001 ,
		_w1236_,
		_w1239_,
		_w1238_,
		_w1240_
	);
	LUT2 #(
		.INIT('h1)
	) name708 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1241_
	);
	LUT4 #(
		.INIT('h0008)
	) name709 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1242_
	);
	LUT3 #(
		.INIT('h54)
	) name710 (
		\sa10_reg[2]/P0001 ,
		_w1242_,
		_w1217_,
		_w1243_
	);
	LUT4 #(
		.INIT('h0800)
	) name711 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1244_
	);
	LUT4 #(
		.INIT('h00ab)
	) name712 (
		\sa10_reg[2]/P0001 ,
		_w1242_,
		_w1217_,
		_w1244_,
		_w1245_
	);
	LUT3 #(
		.INIT('h45)
	) name713 (
		\sa10_reg[1]/P0001 ,
		_w1240_,
		_w1245_,
		_w1246_
	);
	LUT4 #(
		.INIT('h0040)
	) name714 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1247_
	);
	LUT2 #(
		.INIT('h8)
	) name715 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1248_
	);
	LUT4 #(
		.INIT('h0040)
	) name716 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1249_
	);
	LUT3 #(
		.INIT('h54)
	) name717 (
		\sa10_reg[2]/P0001 ,
		_w1247_,
		_w1249_,
		_w1250_
	);
	LUT2 #(
		.INIT('h4)
	) name718 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1251_
	);
	LUT4 #(
		.INIT('h4000)
	) name719 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1252_
	);
	LUT4 #(
		.INIT('h0080)
	) name720 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1253_
	);
	LUT3 #(
		.INIT('h07)
	) name721 (
		\sa10_reg[4]/P0001 ,
		_w1252_,
		_w1253_,
		_w1254_
	);
	LUT2 #(
		.INIT('h2)
	) name722 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		_w1255_
	);
	LUT4 #(
		.INIT('h0200)
	) name723 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1256_
	);
	LUT3 #(
		.INIT('h01)
	) name724 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1257_
	);
	LUT4 #(
		.INIT('h0001)
	) name725 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1258_
	);
	LUT2 #(
		.INIT('h1)
	) name726 (
		_w1256_,
		_w1258_,
		_w1259_
	);
	LUT4 #(
		.INIT('h3111)
	) name727 (
		\sa10_reg[2]/P0001 ,
		_w1250_,
		_w1254_,
		_w1259_,
		_w1260_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name728 (
		\sa10_reg[0]/P0001 ,
		_w1246_,
		_w1233_,
		_w1260_,
		_w1261_
	);
	LUT2 #(
		.INIT('h4)
	) name729 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		_w1262_
	);
	LUT4 #(
		.INIT('h4000)
	) name730 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1263_
	);
	LUT4 #(
		.INIT('h0200)
	) name731 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1264_
	);
	LUT4 #(
		.INIT('h0001)
	) name732 (
		\sa10_reg[1]/P0001 ,
		_w1249_,
		_w1263_,
		_w1264_,
		_w1265_
	);
	LUT2 #(
		.INIT('h4)
	) name733 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1266_
	);
	LUT3 #(
		.INIT('h20)
	) name734 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1267_
	);
	LUT2 #(
		.INIT('h8)
	) name735 (
		_w1251_,
		_w1267_,
		_w1268_
	);
	LUT2 #(
		.INIT('h8)
	) name736 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		_w1269_
	);
	LUT2 #(
		.INIT('h1)
	) name737 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1270_
	);
	LUT3 #(
		.INIT('h10)
	) name738 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1271_
	);
	LUT4 #(
		.INIT('h0100)
	) name739 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1272_
	);
	LUT3 #(
		.INIT('h07)
	) name740 (
		_w1235_,
		_w1269_,
		_w1272_,
		_w1273_
	);
	LUT3 #(
		.INIT('h40)
	) name741 (
		_w1268_,
		_w1265_,
		_w1273_,
		_w1274_
	);
	LUT4 #(
		.INIT('h0001)
	) name742 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1275_
	);
	LUT2 #(
		.INIT('h4)
	) name743 (
		\sa10_reg[4]/P0001 ,
		_w1275_,
		_w1276_
	);
	LUT2 #(
		.INIT('h2)
	) name744 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		_w1277_
	);
	LUT3 #(
		.INIT('h80)
	) name745 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1278_
	);
	LUT3 #(
		.INIT('h7e)
	) name746 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1279_
	);
	LUT2 #(
		.INIT('h2)
	) name747 (
		_w1277_,
		_w1279_,
		_w1280_
	);
	LUT4 #(
		.INIT('h0080)
	) name748 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1281_
	);
	LUT3 #(
		.INIT('h2a)
	) name749 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1281_,
		_w1282_
	);
	LUT3 #(
		.INIT('h10)
	) name750 (
		_w1280_,
		_w1276_,
		_w1282_,
		_w1283_
	);
	LUT3 #(
		.INIT('h04)
	) name751 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1284_
	);
	LUT2 #(
		.INIT('h8)
	) name752 (
		_w1248_,
		_w1284_,
		_w1285_
	);
	LUT2 #(
		.INIT('h1)
	) name753 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1286_
	);
	LUT4 #(
		.INIT('h0004)
	) name754 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1287_
	);
	LUT3 #(
		.INIT('h2a)
	) name755 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1288_
	);
	LUT4 #(
		.INIT('h2220)
	) name756 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1289_
	);
	LUT3 #(
		.INIT('h45)
	) name757 (
		_w1287_,
		_w1288_,
		_w1289_,
		_w1290_
	);
	LUT3 #(
		.INIT('h20)
	) name758 (
		_w1231_,
		_w1288_,
		_w1277_,
		_w1291_
	);
	LUT4 #(
		.INIT('h00ba)
	) name759 (
		\sa10_reg[2]/P0001 ,
		_w1285_,
		_w1290_,
		_w1291_,
		_w1292_
	);
	LUT4 #(
		.INIT('h0155)
	) name760 (
		\sa10_reg[0]/P0001 ,
		_w1274_,
		_w1283_,
		_w1292_,
		_w1293_
	);
	LUT3 #(
		.INIT('h20)
	) name761 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1294_
	);
	LUT4 #(
		.INIT('h0020)
	) name762 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1295_
	);
	LUT4 #(
		.INIT('h5510)
	) name763 (
		\sa10_reg[2]/P0001 ,
		_w1270_,
		_w1294_,
		_w1295_,
		_w1296_
	);
	LUT4 #(
		.INIT('h1000)
	) name764 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1297_
	);
	LUT4 #(
		.INIT('h0800)
	) name765 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1298_
	);
	LUT2 #(
		.INIT('h1)
	) name766 (
		_w1297_,
		_w1298_,
		_w1299_
	);
	LUT4 #(
		.INIT('h4000)
	) name767 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1300_
	);
	LUT3 #(
		.INIT('h08)
	) name768 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1301_
	);
	LUT4 #(
		.INIT('h557f)
	) name769 (
		\sa10_reg[2]/P0001 ,
		_w1234_,
		_w1224_,
		_w1300_,
		_w1302_
	);
	LUT4 #(
		.INIT('h4555)
	) name770 (
		\sa10_reg[1]/P0001 ,
		_w1296_,
		_w1299_,
		_w1302_,
		_w1303_
	);
	LUT2 #(
		.INIT('h8)
	) name771 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[2]/P0001 ,
		_w1304_
	);
	LUT3 #(
		.INIT('h01)
	) name772 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1305_
	);
	LUT4 #(
		.INIT('h0800)
	) name773 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1306_
	);
	LUT4 #(
		.INIT('hf7fa)
	) name774 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1307_
	);
	LUT3 #(
		.INIT('h02)
	) name775 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1308_
	);
	LUT4 #(
		.INIT('h0002)
	) name776 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1309_
	);
	LUT4 #(
		.INIT('hcc04)
	) name777 (
		\sa10_reg[4]/P0001 ,
		_w1304_,
		_w1307_,
		_w1309_,
		_w1310_
	);
	LUT3 #(
		.INIT('h20)
	) name778 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		_w1311_
	);
	LUT2 #(
		.INIT('h8)
	) name779 (
		_w1234_,
		_w1311_,
		_w1312_
	);
	LUT3 #(
		.INIT('h40)
	) name780 (
		\sa10_reg[2]/P0001 ,
		_w1234_,
		_w1311_,
		_w1313_
	);
	LUT4 #(
		.INIT('h2000)
	) name781 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[2]/P0001 ,
		_w1234_,
		_w1311_,
		_w1314_
	);
	LUT2 #(
		.INIT('h2)
	) name782 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[5]/P0001 ,
		_w1315_
	);
	LUT4 #(
		.INIT('hff7a)
	) name783 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1316_
	);
	LUT2 #(
		.INIT('h2)
	) name784 (
		_w1315_,
		_w1316_,
		_w1317_
	);
	LUT4 #(
		.INIT('h0001)
	) name785 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1318_
	);
	LUT2 #(
		.INIT('h4)
	) name786 (
		\sa10_reg[5]/P0001 ,
		_w1318_,
		_w1319_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name787 (
		\sa10_reg[5]/P0001 ,
		_w1244_,
		_w1262_,
		_w1318_,
		_w1320_
	);
	LUT4 #(
		.INIT('h0100)
	) name788 (
		_w1310_,
		_w1317_,
		_w1314_,
		_w1320_,
		_w1321_
	);
	LUT2 #(
		.INIT('h4)
	) name789 (
		_w1303_,
		_w1321_,
		_w1322_
	);
	LUT3 #(
		.INIT('h10)
	) name790 (
		_w1261_,
		_w1293_,
		_w1322_,
		_w1323_
	);
	LUT2 #(
		.INIT('h6)
	) name791 (
		_w1214_,
		_w1323_,
		_w1324_
	);
	LUT3 #(
		.INIT('h96)
	) name792 (
		_w1149_,
		_w1214_,
		_w1323_,
		_w1325_
	);
	LUT2 #(
		.INIT('h2)
	) name793 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1326_
	);
	LUT2 #(
		.INIT('h1)
	) name794 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1327_
	);
	LUT4 #(
		.INIT('h0004)
	) name795 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1328_
	);
	LUT3 #(
		.INIT('h04)
	) name796 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1329_
	);
	LUT2 #(
		.INIT('h8)
	) name797 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w1330_
	);
	LUT3 #(
		.INIT('h80)
	) name798 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1331_
	);
	LUT4 #(
		.INIT('heee4)
	) name799 (
		\sa21_reg[2]/P0001 ,
		_w1328_,
		_w1331_,
		_w1329_,
		_w1332_
	);
	LUT2 #(
		.INIT('h4)
	) name800 (
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1333_
	);
	LUT3 #(
		.INIT('h20)
	) name801 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1334_
	);
	LUT4 #(
		.INIT('h0800)
	) name802 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1335_
	);
	LUT2 #(
		.INIT('h4)
	) name803 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1336_
	);
	LUT4 #(
		.INIT('h1000)
	) name804 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1337_
	);
	LUT2 #(
		.INIT('h1)
	) name805 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1338_
	);
	LUT4 #(
		.INIT('h0008)
	) name806 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1339_
	);
	LUT2 #(
		.INIT('h1)
	) name807 (
		_w1337_,
		_w1339_,
		_w1340_
	);
	LUT4 #(
		.INIT('h2223)
	) name808 (
		\sa21_reg[2]/P0001 ,
		_w1335_,
		_w1337_,
		_w1339_,
		_w1341_
	);
	LUT3 #(
		.INIT('h45)
	) name809 (
		\sa21_reg[1]/P0001 ,
		_w1332_,
		_w1341_,
		_w1342_
	);
	LUT4 #(
		.INIT('h0400)
	) name810 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1343_
	);
	LUT2 #(
		.INIT('h4)
	) name811 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1344_
	);
	LUT3 #(
		.INIT('h10)
	) name812 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1345_
	);
	LUT3 #(
		.INIT('h08)
	) name813 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1346_
	);
	LUT4 #(
		.INIT('h0007)
	) name814 (
		_w1344_,
		_w1345_,
		_w1346_,
		_w1343_,
		_w1347_
	);
	LUT2 #(
		.INIT('h2)
	) name815 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1348_
	);
	LUT2 #(
		.INIT('h2)
	) name816 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1349_
	);
	LUT3 #(
		.INIT('h08)
	) name817 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1350_
	);
	LUT2 #(
		.INIT('h8)
	) name818 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1351_
	);
	LUT3 #(
		.INIT('h80)
	) name819 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1352_
	);
	LUT4 #(
		.INIT('h2000)
	) name820 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1353_
	);
	LUT3 #(
		.INIT('h07)
	) name821 (
		_w1348_,
		_w1350_,
		_w1353_,
		_w1354_
	);
	LUT2 #(
		.INIT('h4)
	) name822 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1355_
	);
	LUT2 #(
		.INIT('h1)
	) name823 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		_w1356_
	);
	LUT3 #(
		.INIT('h01)
	) name824 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		_w1357_
	);
	LUT2 #(
		.INIT('h4)
	) name825 (
		_w1355_,
		_w1357_,
		_w1358_
	);
	LUT4 #(
		.INIT('h0c04)
	) name826 (
		\sa21_reg[2]/P0001 ,
		_w1354_,
		_w1358_,
		_w1347_,
		_w1359_
	);
	LUT2 #(
		.INIT('h4)
	) name827 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w1360_
	);
	LUT4 #(
		.INIT('h0040)
	) name828 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1361_
	);
	LUT4 #(
		.INIT('h0040)
	) name829 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1362_
	);
	LUT3 #(
		.INIT('h54)
	) name830 (
		\sa21_reg[2]/P0001 ,
		_w1361_,
		_w1362_,
		_w1363_
	);
	LUT4 #(
		.INIT('h0080)
	) name831 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1364_
	);
	LUT3 #(
		.INIT('h80)
	) name832 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1365_
	);
	LUT3 #(
		.INIT('h13)
	) name833 (
		_w1360_,
		_w1364_,
		_w1365_,
		_w1366_
	);
	LUT3 #(
		.INIT('h01)
	) name834 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1367_
	);
	LUT4 #(
		.INIT('h0001)
	) name835 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1368_
	);
	LUT2 #(
		.INIT('h2)
	) name836 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		_w1369_
	);
	LUT4 #(
		.INIT('h0200)
	) name837 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1370_
	);
	LUT2 #(
		.INIT('h1)
	) name838 (
		_w1368_,
		_w1370_,
		_w1371_
	);
	LUT4 #(
		.INIT('h3111)
	) name839 (
		\sa21_reg[2]/P0001 ,
		_w1363_,
		_w1366_,
		_w1371_,
		_w1372_
	);
	LUT4 #(
		.INIT('h0d00)
	) name840 (
		\sa21_reg[1]/P0001 ,
		_w1359_,
		_w1342_,
		_w1372_,
		_w1373_
	);
	LUT2 #(
		.INIT('h4)
	) name841 (
		\sa21_reg[2]/P0001 ,
		_w1368_,
		_w1374_
	);
	LUT2 #(
		.INIT('h2)
	) name842 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		_w1375_
	);
	LUT3 #(
		.INIT('h80)
	) name843 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1376_
	);
	LUT3 #(
		.INIT('h7e)
	) name844 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1377_
	);
	LUT2 #(
		.INIT('h8)
	) name845 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1378_
	);
	LUT3 #(
		.INIT('h80)
	) name846 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1379_
	);
	LUT2 #(
		.INIT('h2)
	) name847 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1380_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name848 (
		_w1375_,
		_w1377_,
		_w1379_,
		_w1380_,
		_w1381_
	);
	LUT3 #(
		.INIT('h8a)
	) name849 (
		\sa21_reg[1]/P0001 ,
		_w1374_,
		_w1381_,
		_w1382_
	);
	LUT4 #(
		.INIT('h0200)
	) name850 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1383_
	);
	LUT2 #(
		.INIT('h1)
	) name851 (
		_w1362_,
		_w1383_,
		_w1384_
	);
	LUT3 #(
		.INIT('h10)
	) name852 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1385_
	);
	LUT4 #(
		.INIT('h0100)
	) name853 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1386_
	);
	LUT3 #(
		.INIT('h08)
	) name854 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1387_
	);
	LUT3 #(
		.INIT('h13)
	) name855 (
		_w1349_,
		_w1386_,
		_w1387_,
		_w1388_
	);
	LUT4 #(
		.INIT('h4000)
	) name856 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1389_
	);
	LUT2 #(
		.INIT('h8)
	) name857 (
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1390_
	);
	LUT3 #(
		.INIT('h40)
	) name858 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1391_
	);
	LUT3 #(
		.INIT('h13)
	) name859 (
		_w1360_,
		_w1389_,
		_w1391_,
		_w1392_
	);
	LUT4 #(
		.INIT('h1555)
	) name860 (
		\sa21_reg[1]/P0001 ,
		_w1384_,
		_w1388_,
		_w1392_,
		_w1393_
	);
	LUT3 #(
		.INIT('h01)
	) name861 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1394_
	);
	LUT4 #(
		.INIT('h2000)
	) name862 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1395_
	);
	LUT4 #(
		.INIT('hdefe)
	) name863 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1396_
	);
	LUT2 #(
		.INIT('h2)
	) name864 (
		_w1375_,
		_w1396_,
		_w1397_
	);
	LUT3 #(
		.INIT('h02)
	) name865 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1398_
	);
	LUT4 #(
		.INIT('h0004)
	) name866 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1399_
	);
	LUT4 #(
		.INIT('h0040)
	) name867 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1400_
	);
	LUT2 #(
		.INIT('h1)
	) name868 (
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1401_
	);
	LUT4 #(
		.INIT('h2220)
	) name869 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1402_
	);
	LUT4 #(
		.INIT('h025f)
	) name870 (
		\sa21_reg[4]/P0001 ,
		_w1390_,
		_w1400_,
		_w1402_,
		_w1403_
	);
	LUT4 #(
		.INIT('h2322)
	) name871 (
		\sa21_reg[2]/P0001 ,
		_w1397_,
		_w1399_,
		_w1403_,
		_w1404_
	);
	LUT3 #(
		.INIT('h10)
	) name872 (
		_w1393_,
		_w1382_,
		_w1404_,
		_w1405_
	);
	LUT4 #(
		.INIT('h0800)
	) name873 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1406_
	);
	LUT4 #(
		.INIT('h0020)
	) name874 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1407_
	);
	LUT4 #(
		.INIT('hf7df)
	) name875 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1408_
	);
	LUT3 #(
		.INIT('h45)
	) name876 (
		\sa21_reg[2]/P0001 ,
		_w1406_,
		_w1408_,
		_w1409_
	);
	LUT4 #(
		.INIT('h0800)
	) name877 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1410_
	);
	LUT4 #(
		.INIT('h1000)
	) name878 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1411_
	);
	LUT2 #(
		.INIT('h1)
	) name879 (
		_w1410_,
		_w1411_,
		_w1412_
	);
	LUT4 #(
		.INIT('h4000)
	) name880 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1413_
	);
	LUT2 #(
		.INIT('h8)
	) name881 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		_w1414_
	);
	LUT3 #(
		.INIT('h08)
	) name882 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w1415_
	);
	LUT4 #(
		.INIT('h135f)
	) name883 (
		\sa21_reg[2]/P0001 ,
		_w1401_,
		_w1413_,
		_w1415_,
		_w1416_
	);
	LUT4 #(
		.INIT('h4555)
	) name884 (
		\sa21_reg[1]/P0001 ,
		_w1409_,
		_w1412_,
		_w1416_,
		_w1417_
	);
	LUT2 #(
		.INIT('h8)
	) name885 (
		\sa21_reg[1]/P0001 ,
		\sa21_reg[2]/P0001 ,
		_w1418_
	);
	LUT2 #(
		.INIT('h2)
	) name886 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w1419_
	);
	LUT3 #(
		.INIT('h20)
	) name887 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		_w1420_
	);
	LUT4 #(
		.INIT('h0002)
	) name888 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1421_
	);
	LUT4 #(
		.INIT('h0001)
	) name889 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1422_
	);
	LUT4 #(
		.INIT('h0103)
	) name890 (
		_w1333_,
		_w1421_,
		_w1422_,
		_w1420_,
		_w1423_
	);
	LUT2 #(
		.INIT('h2)
	) name891 (
		_w1418_,
		_w1423_,
		_w1424_
	);
	LUT2 #(
		.INIT('h4)
	) name892 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		_w1425_
	);
	LUT3 #(
		.INIT('h04)
	) name893 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1426_
	);
	LUT4 #(
		.INIT('h0004)
	) name894 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1427_
	);
	LUT2 #(
		.INIT('h8)
	) name895 (
		_w1425_,
		_w1427_,
		_w1428_
	);
	LUT3 #(
		.INIT('h80)
	) name896 (
		\sa21_reg[1]/P0001 ,
		_w1425_,
		_w1427_,
		_w1429_
	);
	LUT4 #(
		.INIT('h0001)
	) name897 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1430_
	);
	LUT4 #(
		.INIT('h0800)
	) name898 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1431_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name899 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1430_,
		_w1431_,
		_w1432_
	);
	LUT2 #(
		.INIT('h8)
	) name900 (
		_w1335_,
		_w1425_,
		_w1433_
	);
	LUT2 #(
		.INIT('h8)
	) name901 (
		_w1327_,
		_w1394_,
		_w1434_
	);
	LUT4 #(
		.INIT('h153f)
	) name902 (
		_w1335_,
		_w1327_,
		_w1394_,
		_w1425_,
		_w1435_
	);
	LUT3 #(
		.INIT('h10)
	) name903 (
		_w1432_,
		_w1429_,
		_w1435_,
		_w1436_
	);
	LUT3 #(
		.INIT('h10)
	) name904 (
		_w1424_,
		_w1417_,
		_w1436_,
		_w1437_
	);
	LUT4 #(
		.INIT('hd800)
	) name905 (
		\sa21_reg[0]/P0001 ,
		_w1373_,
		_w1405_,
		_w1437_,
		_w1438_
	);
	LUT2 #(
		.INIT('h2)
	) name906 (
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1439_
	);
	LUT3 #(
		.INIT('h04)
	) name907 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1440_
	);
	LUT4 #(
		.INIT('h0010)
	) name908 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1441_
	);
	LUT3 #(
		.INIT('h20)
	) name909 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1442_
	);
	LUT2 #(
		.INIT('h4)
	) name910 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w1443_
	);
	LUT2 #(
		.INIT('h2)
	) name911 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1444_
	);
	LUT4 #(
		.INIT('h0040)
	) name912 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1445_
	);
	LUT4 #(
		.INIT('h5554)
	) name913 (
		\sa32_reg[2]/P0001 ,
		_w1442_,
		_w1445_,
		_w1441_,
		_w1446_
	);
	LUT2 #(
		.INIT('h8)
	) name914 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1447_
	);
	LUT3 #(
		.INIT('h80)
	) name915 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1448_
	);
	LUT2 #(
		.INIT('h8)
	) name916 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1449_
	);
	LUT3 #(
		.INIT('h08)
	) name917 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1450_
	);
	LUT4 #(
		.INIT('h0080)
	) name918 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1451_
	);
	LUT3 #(
		.INIT('ha8)
	) name919 (
		\sa32_reg[2]/P0001 ,
		_w1448_,
		_w1451_,
		_w1452_
	);
	LUT3 #(
		.INIT('h40)
	) name920 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1453_
	);
	LUT4 #(
		.INIT('h1000)
	) name921 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1454_
	);
	LUT2 #(
		.INIT('h8)
	) name922 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w1455_
	);
	LUT4 #(
		.INIT('h8000)
	) name923 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1456_
	);
	LUT2 #(
		.INIT('h4)
	) name924 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		_w1457_
	);
	LUT4 #(
		.INIT('h0400)
	) name925 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1458_
	);
	LUT3 #(
		.INIT('h01)
	) name926 (
		_w1454_,
		_w1456_,
		_w1458_,
		_w1459_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1460_
	);
	LUT3 #(
		.INIT('h02)
	) name928 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1461_
	);
	LUT4 #(
		.INIT('h0002)
	) name929 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1462_
	);
	LUT2 #(
		.INIT('h1)
	) name930 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w1463_
	);
	LUT3 #(
		.INIT('h13)
	) name931 (
		_w1450_,
		_w1462_,
		_w1463_,
		_w1464_
	);
	LUT4 #(
		.INIT('h1000)
	) name932 (
		_w1452_,
		_w1446_,
		_w1459_,
		_w1464_,
		_w1465_
	);
	LUT2 #(
		.INIT('h2)
	) name933 (
		\sa32_reg[1]/P0001 ,
		_w1465_,
		_w1466_
	);
	LUT2 #(
		.INIT('h2)
	) name934 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w1467_
	);
	LUT3 #(
		.INIT('h02)
	) name935 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1468_
	);
	LUT4 #(
		.INIT('h0008)
	) name936 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1469_
	);
	LUT4 #(
		.INIT('h0400)
	) name937 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1470_
	);
	LUT3 #(
		.INIT('h54)
	) name938 (
		\sa32_reg[5]/P0001 ,
		_w1469_,
		_w1470_,
		_w1471_
	);
	LUT3 #(
		.INIT('h01)
	) name939 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1472_
	);
	LUT4 #(
		.INIT('h0001)
	) name940 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1473_
	);
	LUT2 #(
		.INIT('h8)
	) name941 (
		\sa32_reg[2]/P0001 ,
		_w1473_,
		_w1474_
	);
	LUT3 #(
		.INIT('h80)
	) name942 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1475_
	);
	LUT4 #(
		.INIT('h4000)
	) name943 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1476_
	);
	LUT2 #(
		.INIT('h4)
	) name944 (
		\sa32_reg[4]/P0001 ,
		_w1476_,
		_w1477_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name945 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w1473_,
		_w1476_,
		_w1478_
	);
	LUT3 #(
		.INIT('h45)
	) name946 (
		\sa32_reg[1]/P0001 ,
		_w1471_,
		_w1478_,
		_w1479_
	);
	LUT3 #(
		.INIT('h04)
	) name947 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1480_
	);
	LUT2 #(
		.INIT('h8)
	) name948 (
		_w1443_,
		_w1480_,
		_w1481_
	);
	LUT2 #(
		.INIT('h1)
	) name949 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1482_
	);
	LUT2 #(
		.INIT('h2)
	) name950 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		_w1483_
	);
	LUT3 #(
		.INIT('hd0)
	) name951 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1484_
	);
	LUT3 #(
		.INIT('h31)
	) name952 (
		_w1482_,
		_w1456_,
		_w1484_,
		_w1485_
	);
	LUT3 #(
		.INIT('h8a)
	) name953 (
		\sa32_reg[2]/P0001 ,
		_w1481_,
		_w1485_,
		_w1486_
	);
	LUT2 #(
		.INIT('h4)
	) name954 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		_w1487_
	);
	LUT3 #(
		.INIT('h02)
	) name955 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1488_
	);
	LUT2 #(
		.INIT('h1)
	) name956 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w1489_
	);
	LUT4 #(
		.INIT('h153f)
	) name957 (
		_w1453_,
		_w1487_,
		_w1488_,
		_w1489_,
		_w1490_
	);
	LUT2 #(
		.INIT('h8)
	) name958 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1491_
	);
	LUT4 #(
		.INIT('h0800)
	) name959 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1492_
	);
	LUT4 #(
		.INIT('h0001)
	) name960 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1493_
	);
	LUT3 #(
		.INIT('h0b)
	) name961 (
		\sa32_reg[2]/P0001 ,
		_w1492_,
		_w1493_,
		_w1494_
	);
	LUT2 #(
		.INIT('h8)
	) name962 (
		_w1490_,
		_w1494_,
		_w1495_
	);
	LUT3 #(
		.INIT('h10)
	) name963 (
		_w1479_,
		_w1486_,
		_w1495_,
		_w1496_
	);
	LUT3 #(
		.INIT('h45)
	) name964 (
		\sa32_reg[0]/P0002 ,
		_w1466_,
		_w1496_,
		_w1497_
	);
	LUT3 #(
		.INIT('h20)
	) name965 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		_w1498_
	);
	LUT2 #(
		.INIT('h4)
	) name966 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1499_
	);
	LUT3 #(
		.INIT('h23)
	) name967 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1500_
	);
	LUT4 #(
		.INIT('h0123)
	) name968 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1501_
	);
	LUT3 #(
		.INIT('ha8)
	) name969 (
		\sa32_reg[1]/P0001 ,
		_w1498_,
		_w1501_,
		_w1502_
	);
	LUT4 #(
		.INIT('h0080)
	) name970 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1503_
	);
	LUT2 #(
		.INIT('h8)
	) name971 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1504_
	);
	LUT4 #(
		.INIT('h0020)
	) name972 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1505_
	);
	LUT2 #(
		.INIT('h2)
	) name973 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1506_
	);
	LUT3 #(
		.INIT('h04)
	) name974 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1507_
	);
	LUT3 #(
		.INIT('h01)
	) name975 (
		_w1503_,
		_w1505_,
		_w1507_,
		_w1508_
	);
	LUT3 #(
		.INIT('h45)
	) name976 (
		\sa32_reg[2]/P0001 ,
		_w1502_,
		_w1508_,
		_w1509_
	);
	LUT4 #(
		.INIT('h4000)
	) name977 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1510_
	);
	LUT4 #(
		.INIT('h0105)
	) name978 (
		\sa32_reg[1]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1503_,
		_w1510_,
		_w1511_
	);
	LUT4 #(
		.INIT('h0008)
	) name979 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1512_
	);
	LUT3 #(
		.INIT('h10)
	) name980 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1513_
	);
	LUT4 #(
		.INIT('h0200)
	) name981 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1514_
	);
	LUT4 #(
		.INIT('hfd3f)
	) name982 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1515_
	);
	LUT4 #(
		.INIT('h5702)
	) name983 (
		\sa32_reg[2]/P0001 ,
		_w1512_,
		_w1513_,
		_w1515_,
		_w1516_
	);
	LUT2 #(
		.INIT('h8)
	) name984 (
		_w1511_,
		_w1516_,
		_w1517_
	);
	LUT4 #(
		.INIT('h0200)
	) name985 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1518_
	);
	LUT2 #(
		.INIT('h2)
	) name986 (
		\sa32_reg[1]/P0001 ,
		_w1518_,
		_w1519_
	);
	LUT2 #(
		.INIT('h8)
	) name987 (
		\sa32_reg[7]/P0001 ,
		_w1445_,
		_w1520_
	);
	LUT4 #(
		.INIT('h0080)
	) name988 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1521_
	);
	LUT4 #(
		.INIT('h23af)
	) name989 (
		\sa32_reg[6]/NET0131 ,
		_w1443_,
		_w1521_,
		_w1472_,
		_w1522_
	);
	LUT3 #(
		.INIT('h40)
	) name990 (
		_w1520_,
		_w1519_,
		_w1522_,
		_w1523_
	);
	LUT3 #(
		.INIT('h10)
	) name991 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1524_
	);
	LUT2 #(
		.INIT('h8)
	) name992 (
		_w1482_,
		_w1524_,
		_w1525_
	);
	LUT4 #(
		.INIT('h0777)
	) name993 (
		\sa32_reg[6]/NET0131 ,
		_w1510_,
		_w1482_,
		_w1524_,
		_w1526_
	);
	LUT4 #(
		.INIT('h2000)
	) name994 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1527_
	);
	LUT3 #(
		.INIT('h08)
	) name995 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1528_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name996 (
		\sa32_reg[2]/P0001 ,
		_w1527_,
		_w1528_,
		_w1457_,
		_w1529_
	);
	LUT3 #(
		.INIT('hd0)
	) name997 (
		\sa32_reg[2]/P0001 ,
		_w1526_,
		_w1529_,
		_w1530_
	);
	LUT4 #(
		.INIT('h0e00)
	) name998 (
		_w1517_,
		_w1523_,
		_w1509_,
		_w1530_,
		_w1531_
	);
	LUT3 #(
		.INIT('h10)
	) name999 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1532_
	);
	LUT4 #(
		.INIT('h1000)
	) name1000 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1533_
	);
	LUT4 #(
		.INIT('h0007)
	) name1001 (
		\sa32_reg[6]/NET0131 ,
		_w1521_,
		_w1527_,
		_w1533_,
		_w1534_
	);
	LUT4 #(
		.INIT('h0001)
	) name1002 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1535_
	);
	LUT3 #(
		.INIT('h10)
	) name1003 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1536_
	);
	LUT4 #(
		.INIT('h1445)
	) name1004 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1537_
	);
	LUT3 #(
		.INIT('ha2)
	) name1005 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1538_
	);
	LUT2 #(
		.INIT('h8)
	) name1006 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w1539_
	);
	LUT4 #(
		.INIT('h5455)
	) name1007 (
		_w1535_,
		_w1537_,
		_w1538_,
		_w1539_,
		_w1540_
	);
	LUT4 #(
		.INIT('h0155)
	) name1008 (
		\sa32_reg[1]/P0001 ,
		\sa32_reg[2]/P0001 ,
		_w1534_,
		_w1540_,
		_w1541_
	);
	LUT4 #(
		.INIT('h0080)
	) name1009 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1542_
	);
	LUT2 #(
		.INIT('h8)
	) name1010 (
		_w1443_,
		_w1542_,
		_w1543_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name1011 (
		\sa32_reg[2]/P0001 ,
		_w1472_,
		_w1467_,
		_w1492_,
		_w1544_
	);
	LUT3 #(
		.INIT('h8a)
	) name1012 (
		\sa32_reg[1]/P0001 ,
		_w1543_,
		_w1544_,
		_w1545_
	);
	LUT2 #(
		.INIT('h8)
	) name1013 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		_w1546_
	);
	LUT3 #(
		.INIT('h02)
	) name1014 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1547_
	);
	LUT3 #(
		.INIT('h80)
	) name1015 (
		\sa32_reg[4]/P0001 ,
		_w1546_,
		_w1547_,
		_w1548_
	);
	LUT4 #(
		.INIT('h5450)
	) name1016 (
		\sa32_reg[2]/P0001 ,
		_w1506_,
		_w1454_,
		_w1468_,
		_w1549_
	);
	LUT2 #(
		.INIT('h1)
	) name1017 (
		_w1548_,
		_w1549_,
		_w1550_
	);
	LUT3 #(
		.INIT('h10)
	) name1018 (
		_w1541_,
		_w1545_,
		_w1550_,
		_w1551_
	);
	LUT3 #(
		.INIT('hd0)
	) name1019 (
		\sa32_reg[0]/P0002 ,
		_w1531_,
		_w1551_,
		_w1552_
	);
	LUT4 #(
		.INIT('h9699)
	) name1020 (
		\u0_w_reg[3][6]/P0001 ,
		_w1438_,
		_w1497_,
		_w1552_,
		_w1553_
	);
	LUT3 #(
		.INIT('h82)
	) name1021 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[6]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w1554_
	);
	LUT4 #(
		.INIT('h00be)
	) name1022 (
		\ld_r_reg/P0001 ,
		_w1325_,
		_w1553_,
		_w1554_,
		_w1555_
	);
	LUT4 #(
		.INIT('h0400)
	) name1023 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1556_
	);
	LUT4 #(
		.INIT('h0020)
	) name1024 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1557_
	);
	LUT4 #(
		.INIT('hf5e4)
	) name1025 (
		\sa10_reg[2]/P0001 ,
		_w1228_,
		_w1556_,
		_w1557_,
		_w1558_
	);
	LUT3 #(
		.INIT('h07)
	) name1026 (
		_w1251_,
		_w1267_,
		_w1306_,
		_w1559_
	);
	LUT3 #(
		.INIT('h8a)
	) name1027 (
		\sa10_reg[1]/P0001 ,
		_w1558_,
		_w1559_,
		_w1560_
	);
	LUT4 #(
		.INIT('h0010)
	) name1028 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1561_
	);
	LUT2 #(
		.INIT('h1)
	) name1029 (
		_w1252_,
		_w1561_,
		_w1562_
	);
	LUT3 #(
		.INIT('h07)
	) name1030 (
		\sa10_reg[4]/P0001 ,
		_w1281_,
		_w1309_,
		_w1563_
	);
	LUT3 #(
		.INIT('h15)
	) name1031 (
		\sa10_reg[2]/P0001 ,
		_w1562_,
		_w1563_,
		_w1564_
	);
	LUT3 #(
		.INIT('h80)
	) name1032 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1565_
	);
	LUT2 #(
		.INIT('h8)
	) name1033 (
		_w1216_,
		_w1565_,
		_w1566_
	);
	LUT2 #(
		.INIT('h2)
	) name1034 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1567_
	);
	LUT4 #(
		.INIT('h0002)
	) name1035 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1568_
	);
	LUT3 #(
		.INIT('h10)
	) name1036 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1569_
	);
	LUT3 #(
		.INIT('h01)
	) name1037 (
		_w1225_,
		_w1569_,
		_w1568_,
		_w1570_
	);
	LUT4 #(
		.INIT('h0008)
	) name1038 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1571_
	);
	LUT4 #(
		.INIT('h8000)
	) name1039 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1572_
	);
	LUT4 #(
		.INIT('h7ff6)
	) name1040 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1573_
	);
	LUT2 #(
		.INIT('h2)
	) name1041 (
		_w1269_,
		_w1573_,
		_w1574_
	);
	LUT4 #(
		.INIT('h00ba)
	) name1042 (
		\sa10_reg[1]/P0001 ,
		_w1566_,
		_w1570_,
		_w1574_,
		_w1575_
	);
	LUT4 #(
		.INIT('h5455)
	) name1043 (
		\sa10_reg[0]/P0001 ,
		_w1564_,
		_w1560_,
		_w1575_,
		_w1576_
	);
	LUT4 #(
		.INIT('h0010)
	) name1044 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1577_
	);
	LUT4 #(
		.INIT('hbfef)
	) name1045 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1578_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name1046 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1579_
	);
	LUT2 #(
		.INIT('h2)
	) name1047 (
		_w1262_,
		_w1579_,
		_w1580_
	);
	LUT3 #(
		.INIT('had)
	) name1048 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1581_
	);
	LUT4 #(
		.INIT('h0004)
	) name1049 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1582_
	);
	LUT4 #(
		.INIT('hadfb)
	) name1050 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1583_
	);
	LUT4 #(
		.INIT('h0302)
	) name1051 (
		\sa10_reg[3]/P0001 ,
		_w1217_,
		_w1281_,
		_w1583_,
		_w1584_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1052 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[2]/P0001 ,
		_w1580_,
		_w1584_,
		_w1585_
	);
	LUT3 #(
		.INIT('h51)
	) name1053 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1586_
	);
	LUT4 #(
		.INIT('h7511)
	) name1054 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1587_
	);
	LUT2 #(
		.INIT('h2)
	) name1055 (
		_w1586_,
		_w1587_,
		_w1588_
	);
	LUT4 #(
		.INIT('h0040)
	) name1056 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1589_
	);
	LUT4 #(
		.INIT('h0020)
	) name1057 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1590_
	);
	LUT4 #(
		.INIT('h0010)
	) name1058 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1591_
	);
	LUT4 #(
		.INIT('h0007)
	) name1059 (
		_w1271_,
		_w1315_,
		_w1590_,
		_w1591_,
		_w1592_
	);
	LUT4 #(
		.INIT('h5455)
	) name1060 (
		\sa10_reg[1]/P0001 ,
		_w1588_,
		_w1589_,
		_w1592_,
		_w1593_
	);
	LUT4 #(
		.INIT('h0100)
	) name1061 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1594_
	);
	LUT4 #(
		.INIT('h8cbf)
	) name1062 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1238_,
		_w1594_,
		_w1595_
	);
	LUT2 #(
		.INIT('h8)
	) name1063 (
		\sa10_reg[4]/P0001 ,
		_w1591_,
		_w1596_
	);
	LUT4 #(
		.INIT('h0040)
	) name1064 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1597_
	);
	LUT3 #(
		.INIT('h07)
	) name1065 (
		_w1266_,
		_w1301_,
		_w1597_,
		_w1598_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1066 (
		\sa10_reg[1]/P0001 ,
		_w1595_,
		_w1596_,
		_w1598_,
		_w1599_
	);
	LUT3 #(
		.INIT('hf6)
	) name1067 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1600_
	);
	LUT3 #(
		.INIT('h2a)
	) name1068 (
		_w1304_,
		_w1581_,
		_w1600_,
		_w1601_
	);
	LUT4 #(
		.INIT('h0080)
	) name1069 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1602_
	);
	LUT4 #(
		.INIT('h1000)
	) name1070 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1603_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1071 (
		\sa10_reg[2]/P0001 ,
		_w1247_,
		_w1603_,
		_w1602_,
		_w1604_
	);
	LUT2 #(
		.INIT('h1)
	) name1072 (
		_w1601_,
		_w1604_,
		_w1605_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1073 (
		\sa10_reg[0]/P0001 ,
		_w1593_,
		_w1599_,
		_w1605_,
		_w1606_
	);
	LUT4 #(
		.INIT('h4000)
	) name1074 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1607_
	);
	LUT4 #(
		.INIT('hbdff)
	) name1075 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1608_
	);
	LUT3 #(
		.INIT('h10)
	) name1076 (
		_w1252_,
		_w1561_,
		_w1608_,
		_w1609_
	);
	LUT3 #(
		.INIT('h51)
	) name1077 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[2]/P0001 ,
		_w1607_,
		_w1610_
	);
	LUT2 #(
		.INIT('h4)
	) name1078 (
		_w1609_,
		_w1610_,
		_w1611_
	);
	LUT4 #(
		.INIT('h8caf)
	) name1079 (
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1242_,
		_w1297_,
		_w1612_
	);
	LUT2 #(
		.INIT('h4)
	) name1080 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[2]/P0001 ,
		_w1613_
	);
	LUT4 #(
		.INIT('h4000)
	) name1081 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1614_
	);
	LUT4 #(
		.INIT('h0002)
	) name1082 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1615_
	);
	LUT4 #(
		.INIT('h0007)
	) name1083 (
		_w1238_,
		_w1266_,
		_w1614_,
		_w1615_,
		_w1616_
	);
	LUT4 #(
		.INIT('hfcb8)
	) name1084 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[2]/P0001 ,
		_w1612_,
		_w1616_,
		_w1617_
	);
	LUT2 #(
		.INIT('h4)
	) name1085 (
		_w1611_,
		_w1617_,
		_w1618_
	);
	LUT4 #(
		.INIT('h0100)
	) name1086 (
		_w1585_,
		_w1576_,
		_w1606_,
		_w1618_,
		_w1619_
	);
	LUT3 #(
		.INIT('h08)
	) name1087 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1620_
	);
	LUT4 #(
		.INIT('h0020)
	) name1088 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1621_
	);
	LUT3 #(
		.INIT('h54)
	) name1089 (
		\sa03_reg[2]/P0001 ,
		_w1620_,
		_w1621_,
		_w1622_
	);
	LUT2 #(
		.INIT('h1)
	) name1090 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1623_
	);
	LUT4 #(
		.INIT('h0400)
	) name1091 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1624_
	);
	LUT3 #(
		.INIT('h45)
	) name1092 (
		_w1195_,
		_w1623_,
		_w1624_,
		_w1625_
	);
	LUT3 #(
		.INIT('h8a)
	) name1093 (
		\sa03_reg[1]/P0001 ,
		_w1622_,
		_w1625_,
		_w1626_
	);
	LUT4 #(
		.INIT('h0800)
	) name1094 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1627_
	);
	LUT3 #(
		.INIT('hc8)
	) name1095 (
		_w1079_,
		_w1165_,
		_w1627_,
		_w1628_
	);
	LUT3 #(
		.INIT('h8a)
	) name1096 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1629_
	);
	LUT2 #(
		.INIT('h1)
	) name1097 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1630_
	);
	LUT4 #(
		.INIT('h1101)
	) name1098 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1631_
	);
	LUT3 #(
		.INIT('h15)
	) name1099 (
		\sa03_reg[0]/P0001 ,
		_w1629_,
		_w1631_,
		_w1632_
	);
	LUT4 #(
		.INIT('hf2fa)
	) name1100 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		_w1633_
	);
	LUT2 #(
		.INIT('h4)
	) name1101 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1634_
	);
	LUT2 #(
		.INIT('h4)
	) name1102 (
		_w1633_,
		_w1634_,
		_w1635_
	);
	LUT3 #(
		.INIT('h80)
	) name1103 (
		\sa03_reg[2]/P0001 ,
		_w1116_,
		_w1140_,
		_w1636_
	);
	LUT4 #(
		.INIT('h0100)
	) name1104 (
		_w1628_,
		_w1635_,
		_w1636_,
		_w1632_,
		_w1637_
	);
	LUT4 #(
		.INIT('h8000)
	) name1105 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1638_
	);
	LUT4 #(
		.INIT('h7ff7)
	) name1106 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1639_
	);
	LUT2 #(
		.INIT('h2)
	) name1107 (
		_w1115_,
		_w1639_,
		_w1640_
	);
	LUT4 #(
		.INIT('h5540)
	) name1108 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[5]/P0001 ,
		_w1130_,
		_w1202_,
		_w1641_
	);
	LUT2 #(
		.INIT('h1)
	) name1109 (
		_w1640_,
		_w1641_,
		_w1642_
	);
	LUT3 #(
		.INIT('h40)
	) name1110 (
		_w1626_,
		_w1637_,
		_w1642_,
		_w1643_
	);
	LUT3 #(
		.INIT('h80)
	) name1111 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1644_
	);
	LUT4 #(
		.INIT('h7d5d)
	) name1112 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1645_
	);
	LUT2 #(
		.INIT('h1)
	) name1113 (
		\sa03_reg[2]/P0001 ,
		_w1645_,
		_w1646_
	);
	LUT3 #(
		.INIT('h8a)
	) name1114 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1647_
	);
	LUT4 #(
		.INIT('h00d0)
	) name1115 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1648_
	);
	LUT2 #(
		.INIT('h4)
	) name1116 (
		_w1647_,
		_w1648_,
		_w1649_
	);
	LUT3 #(
		.INIT('h10)
	) name1117 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1650_
	);
	LUT4 #(
		.INIT('h0020)
	) name1118 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1651_
	);
	LUT3 #(
		.INIT('h07)
	) name1119 (
		_w1069_,
		_w1650_,
		_w1651_,
		_w1652_
	);
	LUT4 #(
		.INIT('h5455)
	) name1120 (
		\sa03_reg[1]/P0001 ,
		_w1646_,
		_w1649_,
		_w1652_,
		_w1653_
	);
	LUT3 #(
		.INIT('h09)
	) name1121 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1654_
	);
	LUT3 #(
		.INIT('had)
	) name1122 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1655_
	);
	LUT3 #(
		.INIT('h8a)
	) name1123 (
		\sa03_reg[2]/P0001 ,
		_w1654_,
		_w1655_,
		_w1656_
	);
	LUT4 #(
		.INIT('h0800)
	) name1124 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1657_
	);
	LUT4 #(
		.INIT('h0100)
	) name1125 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1658_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name1126 (
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1657_,
		_w1658_,
		_w1659_
	);
	LUT3 #(
		.INIT('h8a)
	) name1127 (
		\sa03_reg[1]/P0001 ,
		_w1656_,
		_w1659_,
		_w1660_
	);
	LUT4 #(
		.INIT('ha7f7)
	) name1128 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1661_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name1129 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1090_,
		_w1661_,
		_w1662_
	);
	LUT2 #(
		.INIT('h8)
	) name1130 (
		_w1155_,
		_w1630_,
		_w1663_
	);
	LUT4 #(
		.INIT('h0040)
	) name1131 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1664_
	);
	LUT4 #(
		.INIT('h002a)
	) name1132 (
		\sa03_reg[0]/P0001 ,
		_w1115_,
		_w1063_,
		_w1664_,
		_w1665_
	);
	LUT3 #(
		.INIT('h10)
	) name1133 (
		_w1662_,
		_w1663_,
		_w1665_,
		_w1666_
	);
	LUT3 #(
		.INIT('h10)
	) name1134 (
		_w1660_,
		_w1653_,
		_w1666_,
		_w1667_
	);
	LUT4 #(
		.INIT('h0010)
	) name1135 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1668_
	);
	LUT4 #(
		.INIT('hbfef)
	) name1136 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1669_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name1137 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1670_
	);
	LUT2 #(
		.INIT('h2)
	) name1138 (
		_w1068_,
		_w1670_,
		_w1671_
	);
	LUT4 #(
		.INIT('h0200)
	) name1139 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1672_
	);
	LUT4 #(
		.INIT('hadfb)
	) name1140 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1673_
	);
	LUT4 #(
		.INIT('h1302)
	) name1141 (
		\sa03_reg[3]/P0001 ,
		_w1112_,
		_w1045_,
		_w1673_,
		_w1674_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1142 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[2]/P0001 ,
		_w1671_,
		_w1674_,
		_w1675_
	);
	LUT4 #(
		.INIT('h0040)
	) name1143 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1676_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name1144 (
		\sa03_reg[4]/P0001 ,
		_w1116_,
		_w1620_,
		_w1676_,
		_w1677_
	);
	LUT2 #(
		.INIT('h1)
	) name1145 (
		\sa03_reg[2]/P0001 ,
		_w1677_,
		_w1678_
	);
	LUT4 #(
		.INIT('h0103)
	) name1146 (
		\sa03_reg[7]/NET0131 ,
		_w1097_,
		_w1138_,
		_w1657_,
		_w1679_
	);
	LUT2 #(
		.INIT('h8)
	) name1147 (
		_w1068_,
		_w1650_,
		_w1680_
	);
	LUT4 #(
		.INIT('h4000)
	) name1148 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1681_
	);
	LUT3 #(
		.INIT('h07)
	) name1149 (
		_w1629_,
		_w1631_,
		_w1681_,
		_w1682_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1150 (
		\sa03_reg[2]/P0001 ,
		_w1679_,
		_w1680_,
		_w1682_,
		_w1683_
	);
	LUT4 #(
		.INIT('h0302)
	) name1151 (
		\sa03_reg[1]/P0001 ,
		_w1675_,
		_w1678_,
		_w1683_,
		_w1684_
	);
	LUT3 #(
		.INIT('he0)
	) name1152 (
		_w1643_,
		_w1667_,
		_w1684_,
		_w1685_
	);
	LUT3 #(
		.INIT('h69)
	) name1153 (
		_w1214_,
		_w1619_,
		_w1685_,
		_w1686_
	);
	LUT4 #(
		.INIT('h0004)
	) name1154 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1687_
	);
	LUT2 #(
		.INIT('h1)
	) name1155 (
		\sa32_reg[2]/P0001 ,
		_w1687_,
		_w1688_
	);
	LUT3 #(
		.INIT('h80)
	) name1156 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1689_
	);
	LUT4 #(
		.INIT('hfad8)
	) name1157 (
		\sa32_reg[2]/P0001 ,
		_w1480_,
		_w1687_,
		_w1689_,
		_w1690_
	);
	LUT4 #(
		.INIT('h5545)
	) name1158 (
		\sa32_reg[1]/P0001 ,
		_w1492_,
		_w1490_,
		_w1690_,
		_w1691_
	);
	LUT4 #(
		.INIT('h0100)
	) name1159 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1692_
	);
	LUT3 #(
		.INIT('h08)
	) name1160 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1693_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name1161 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1694_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1162 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1692_,
		_w1694_,
		_w1695_
	);
	LUT4 #(
		.INIT('h2000)
	) name1163 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1696_
	);
	LUT3 #(
		.INIT('h0b)
	) name1164 (
		\sa32_reg[6]/NET0131 ,
		_w1521_,
		_w1696_,
		_w1697_
	);
	LUT2 #(
		.INIT('h1)
	) name1165 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		_w1698_
	);
	LUT2 #(
		.INIT('h8)
	) name1166 (
		_w1500_,
		_w1698_,
		_w1699_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1167 (
		\sa32_reg[1]/P0001 ,
		_w1697_,
		_w1699_,
		_w1695_,
		_w1700_
	);
	LUT4 #(
		.INIT('h0040)
	) name1168 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1701_
	);
	LUT3 #(
		.INIT('h54)
	) name1169 (
		\sa32_reg[2]/P0001 ,
		_w1445_,
		_w1701_,
		_w1702_
	);
	LUT4 #(
		.INIT('h0080)
	) name1170 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1703_
	);
	LUT3 #(
		.INIT('h07)
	) name1171 (
		\sa32_reg[6]/NET0131 ,
		_w1510_,
		_w1703_,
		_w1704_
	);
	LUT2 #(
		.INIT('h1)
	) name1172 (
		_w1514_,
		_w1493_,
		_w1705_
	);
	LUT4 #(
		.INIT('h3111)
	) name1173 (
		\sa32_reg[2]/P0001 ,
		_w1702_,
		_w1704_,
		_w1705_,
		_w1706_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1174 (
		\sa32_reg[0]/P0002 ,
		_w1700_,
		_w1691_,
		_w1706_,
		_w1707_
	);
	LUT3 #(
		.INIT('he6)
	) name1175 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1708_
	);
	LUT2 #(
		.INIT('h2)
	) name1176 (
		_w1443_,
		_w1708_,
		_w1709_
	);
	LUT4 #(
		.INIT('h2220)
	) name1177 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1710_
	);
	LUT3 #(
		.INIT('h2a)
	) name1178 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1711_
	);
	LUT3 #(
		.INIT('h51)
	) name1179 (
		\sa32_reg[2]/P0001 ,
		_w1710_,
		_w1711_,
		_w1712_
	);
	LUT4 #(
		.INIT('h0001)
	) name1180 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1713_
	);
	LUT4 #(
		.INIT('h002a)
	) name1181 (
		\sa32_reg[2]/P0001 ,
		_w1491_,
		_w1524_,
		_w1713_,
		_w1714_
	);
	LUT3 #(
		.INIT('h0b)
	) name1182 (
		_w1709_,
		_w1712_,
		_w1714_,
		_w1715_
	);
	LUT4 #(
		.INIT('h0200)
	) name1183 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1716_
	);
	LUT3 #(
		.INIT('h01)
	) name1184 (
		\sa32_reg[1]/P0001 ,
		_w1701_,
		_w1716_,
		_w1717_
	);
	LUT4 #(
		.INIT('h4000)
	) name1185 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1718_
	);
	LUT3 #(
		.INIT('h07)
	) name1186 (
		_w1546_,
		_w1547_,
		_w1718_,
		_w1719_
	);
	LUT3 #(
		.INIT('h10)
	) name1187 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1720_
	);
	LUT4 #(
		.INIT('h0100)
	) name1188 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1721_
	);
	LUT3 #(
		.INIT('h07)
	) name1189 (
		_w1491_,
		_w1524_,
		_w1721_,
		_w1722_
	);
	LUT3 #(
		.INIT('h80)
	) name1190 (
		_w1717_,
		_w1719_,
		_w1722_,
		_w1723_
	);
	LUT2 #(
		.INIT('h2)
	) name1191 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		_w1724_
	);
	LUT3 #(
		.INIT('h80)
	) name1192 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1725_
	);
	LUT3 #(
		.INIT('h01)
	) name1193 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1726_
	);
	LUT3 #(
		.INIT('h7e)
	) name1194 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1727_
	);
	LUT2 #(
		.INIT('h2)
	) name1195 (
		_w1724_,
		_w1727_,
		_w1728_
	);
	LUT2 #(
		.INIT('h4)
	) name1196 (
		\sa32_reg[2]/P0001 ,
		_w1493_,
		_w1729_
	);
	LUT3 #(
		.INIT('h2a)
	) name1197 (
		\sa32_reg[1]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1521_,
		_w1730_
	);
	LUT3 #(
		.INIT('h10)
	) name1198 (
		_w1728_,
		_w1729_,
		_w1730_,
		_w1731_
	);
	LUT4 #(
		.INIT('h4445)
	) name1199 (
		\sa32_reg[0]/P0002 ,
		_w1715_,
		_w1723_,
		_w1731_,
		_w1732_
	);
	LUT4 #(
		.INIT('h0800)
	) name1200 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1733_
	);
	LUT4 #(
		.INIT('h0020)
	) name1201 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1734_
	);
	LUT4 #(
		.INIT('hf7df)
	) name1202 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1735_
	);
	LUT3 #(
		.INIT('h45)
	) name1203 (
		\sa32_reg[2]/P0001 ,
		_w1733_,
		_w1735_,
		_w1736_
	);
	LUT2 #(
		.INIT('h2)
	) name1204 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w1737_
	);
	LUT4 #(
		.INIT('h0002)
	) name1205 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1738_
	);
	LUT2 #(
		.INIT('h8)
	) name1206 (
		\sa32_reg[3]/P0001 ,
		_w1738_,
		_w1739_
	);
	LUT4 #(
		.INIT('h4000)
	) name1207 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1740_
	);
	LUT4 #(
		.INIT('h1000)
	) name1208 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1741_
	);
	LUT4 #(
		.INIT('h0800)
	) name1209 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1742_
	);
	LUT4 #(
		.INIT('h0013)
	) name1210 (
		\sa32_reg[2]/P0001 ,
		_w1741_,
		_w1740_,
		_w1742_,
		_w1743_
	);
	LUT4 #(
		.INIT('h5455)
	) name1211 (
		\sa32_reg[1]/P0001 ,
		_w1739_,
		_w1736_,
		_w1743_,
		_w1744_
	);
	LUT2 #(
		.INIT('h8)
	) name1212 (
		_w1444_,
		_w1718_,
		_w1745_
	);
	LUT3 #(
		.INIT('h01)
	) name1213 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1746_
	);
	LUT2 #(
		.INIT('h8)
	) name1214 (
		_w1460_,
		_w1746_,
		_w1747_
	);
	LUT4 #(
		.INIT('h0020)
	) name1215 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1748_
	);
	LUT4 #(
		.INIT('h135f)
	) name1216 (
		_w1460_,
		_w1539_,
		_w1746_,
		_w1748_,
		_w1749_
	);
	LUT3 #(
		.INIT('h10)
	) name1217 (
		_w1474_,
		_w1745_,
		_w1749_,
		_w1750_
	);
	LUT3 #(
		.INIT('h40)
	) name1218 (
		\sa32_reg[2]/P0001 ,
		_w1506_,
		_w1468_,
		_w1751_
	);
	LUT4 #(
		.INIT('h2000)
	) name1219 (
		\sa32_reg[1]/P0001 ,
		\sa32_reg[2]/P0001 ,
		_w1506_,
		_w1468_,
		_w1752_
	);
	LUT4 #(
		.INIT('hdfe2)
	) name1220 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1753_
	);
	LUT2 #(
		.INIT('h8)
	) name1221 (
		\sa32_reg[1]/P0001 ,
		\sa32_reg[2]/P0001 ,
		_w1754_
	);
	LUT3 #(
		.INIT('h08)
	) name1222 (
		\sa32_reg[1]/P0001 ,
		\sa32_reg[2]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1755_
	);
	LUT2 #(
		.INIT('h4)
	) name1223 (
		_w1753_,
		_w1755_,
		_w1756_
	);
	LUT2 #(
		.INIT('h1)
	) name1224 (
		_w1752_,
		_w1756_,
		_w1757_
	);
	LUT3 #(
		.INIT('h40)
	) name1225 (
		_w1744_,
		_w1750_,
		_w1757_,
		_w1758_
	);
	LUT3 #(
		.INIT('h10)
	) name1226 (
		_w1707_,
		_w1732_,
		_w1758_,
		_w1759_
	);
	LUT4 #(
		.INIT('h0020)
	) name1227 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1760_
	);
	LUT4 #(
		.INIT('h0010)
	) name1228 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1761_
	);
	LUT2 #(
		.INIT('h1)
	) name1229 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1762_
	);
	LUT4 #(
		.INIT('h0040)
	) name1230 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1763_
	);
	LUT3 #(
		.INIT('h01)
	) name1231 (
		_w1761_,
		_w1760_,
		_w1763_,
		_w1764_
	);
	LUT2 #(
		.INIT('h4)
	) name1232 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w1765_
	);
	LUT4 #(
		.INIT('h4404)
	) name1233 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1766_
	);
	LUT2 #(
		.INIT('h4)
	) name1234 (
		_w1391_,
		_w1766_,
		_w1767_
	);
	LUT4 #(
		.INIT('h0040)
	) name1235 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1768_
	);
	LUT2 #(
		.INIT('h4)
	) name1236 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1769_
	);
	LUT3 #(
		.INIT('h02)
	) name1237 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w1770_
	);
	LUT3 #(
		.INIT('h15)
	) name1238 (
		_w1768_,
		_w1769_,
		_w1770_,
		_w1771_
	);
	LUT4 #(
		.INIT('h4555)
	) name1239 (
		\sa21_reg[1]/P0001 ,
		_w1767_,
		_w1764_,
		_w1771_,
		_w1772_
	);
	LUT3 #(
		.INIT('h01)
	) name1240 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1773_
	);
	LUT3 #(
		.INIT('hf6)
	) name1241 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1774_
	);
	LUT3 #(
		.INIT('had)
	) name1242 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1775_
	);
	LUT3 #(
		.INIT('h2a)
	) name1243 (
		\sa21_reg[1]/P0001 ,
		_w1774_,
		_w1775_,
		_w1776_
	);
	LUT4 #(
		.INIT('h0080)
	) name1244 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1777_
	);
	LUT4 #(
		.INIT('h1000)
	) name1245 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1778_
	);
	LUT3 #(
		.INIT('h01)
	) name1246 (
		_w1361_,
		_w1778_,
		_w1777_,
		_w1779_
	);
	LUT3 #(
		.INIT('h8a)
	) name1247 (
		\sa21_reg[2]/P0001 ,
		_w1776_,
		_w1779_,
		_w1780_
	);
	LUT3 #(
		.INIT('h10)
	) name1248 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1781_
	);
	LUT4 #(
		.INIT('h153f)
	) name1249 (
		_w1356_,
		_w1330_,
		_w1391_,
		_w1781_,
		_w1782_
	);
	LUT2 #(
		.INIT('h8)
	) name1250 (
		_w1356_,
		_w1346_,
		_w1783_
	);
	LUT4 #(
		.INIT('h0040)
	) name1251 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1784_
	);
	LUT3 #(
		.INIT('h07)
	) name1252 (
		_w1345_,
		_w1414_,
		_w1784_,
		_w1785_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1253 (
		\sa21_reg[1]/P0001 ,
		_w1782_,
		_w1783_,
		_w1785_,
		_w1786_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1254 (
		\sa21_reg[0]/P0001 ,
		_w1780_,
		_w1772_,
		_w1786_,
		_w1787_
	);
	LUT4 #(
		.INIT('h0010)
	) name1255 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1788_
	);
	LUT4 #(
		.INIT('hbfef)
	) name1256 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1789_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name1257 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1790_
	);
	LUT2 #(
		.INIT('h2)
	) name1258 (
		_w1425_,
		_w1790_,
		_w1791_
	);
	LUT4 #(
		.INIT('h0200)
	) name1259 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1792_
	);
	LUT4 #(
		.INIT('hadfb)
	) name1260 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1793_
	);
	LUT4 #(
		.INIT('h0080)
	) name1261 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1794_
	);
	LUT4 #(
		.INIT('h0032)
	) name1262 (
		\sa21_reg[3]/P0001 ,
		_w1337_,
		_w1793_,
		_w1794_,
		_w1795_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1263 (
		\sa21_reg[1]/P0001 ,
		\sa21_reg[2]/P0001 ,
		_w1791_,
		_w1795_,
		_w1796_
	);
	LUT3 #(
		.INIT('h02)
	) name1264 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1797_
	);
	LUT4 #(
		.INIT('h0008)
	) name1265 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1798_
	);
	LUT4 #(
		.INIT('h8000)
	) name1266 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1799_
	);
	LUT3 #(
		.INIT('h20)
	) name1267 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1800_
	);
	LUT4 #(
		.INIT('h0400)
	) name1268 (
		\sa21_reg[1]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1801_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1269 (
		_w1414_,
		_w1799_,
		_w1801_,
		_w1798_,
		_w1802_
	);
	LUT3 #(
		.INIT('h01)
	) name1270 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1803_
	);
	LUT4 #(
		.INIT('h0002)
	) name1271 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1804_
	);
	LUT2 #(
		.INIT('h1)
	) name1272 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w1805_
	);
	LUT4 #(
		.INIT('hf2fa)
	) name1273 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		_w1806_
	);
	LUT4 #(
		.INIT('h5054)
	) name1274 (
		\sa21_reg[1]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1804_,
		_w1806_,
		_w1807_
	);
	LUT4 #(
		.INIT('h5540)
	) name1275 (
		\sa21_reg[2]/P0001 ,
		_w1379_,
		_w1380_,
		_w1421_,
		_w1808_
	);
	LUT4 #(
		.INIT('h3fbb)
	) name1276 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1809_
	);
	LUT2 #(
		.INIT('h2)
	) name1277 (
		_w1356_,
		_w1809_,
		_w1810_
	);
	LUT4 #(
		.INIT('h7f6e)
	) name1278 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		_w1368_,
		_w1809_,
		_w1811_
	);
	LUT4 #(
		.INIT('h0100)
	) name1279 (
		_w1807_,
		_w1808_,
		_w1802_,
		_w1811_,
		_w1812_
	);
	LUT2 #(
		.INIT('h1)
	) name1280 (
		\sa21_reg[0]/P0001 ,
		_w1812_,
		_w1813_
	);
	LUT4 #(
		.INIT('h4000)
	) name1281 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1814_
	);
	LUT4 #(
		.INIT('h0002)
	) name1282 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1815_
	);
	LUT4 #(
		.INIT('h0007)
	) name1283 (
		_w1330_,
		_w1391_,
		_w1815_,
		_w1814_,
		_w1816_
	);
	LUT4 #(
		.INIT('h4000)
	) name1284 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1817_
	);
	LUT3 #(
		.INIT('h0b)
	) name1285 (
		\sa21_reg[2]/P0001 ,
		_w1383_,
		_w1817_,
		_w1818_
	);
	LUT4 #(
		.INIT('h3100)
	) name1286 (
		\sa21_reg[2]/P0001 ,
		_w1810_,
		_w1816_,
		_w1818_,
		_w1819_
	);
	LUT4 #(
		.INIT('h0400)
	) name1287 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1820_
	);
	LUT2 #(
		.INIT('h4)
	) name1288 (
		_w1762_,
		_w1820_,
		_w1821_
	);
	LUT4 #(
		.INIT('h0020)
	) name1289 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w1822_
	);
	LUT4 #(
		.INIT('h0a0b)
	) name1290 (
		\sa21_reg[2]/P0001 ,
		_w1350_,
		_w1406_,
		_w1822_,
		_w1823_
	);
	LUT2 #(
		.INIT('h4)
	) name1291 (
		\sa21_reg[0]/P0001 ,
		\sa21_reg[1]/P0001 ,
		_w1824_
	);
	LUT4 #(
		.INIT('h0008)
	) name1292 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1825_
	);
	LUT4 #(
		.INIT('heff7)
	) name1293 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w1826_
	);
	LUT2 #(
		.INIT('h2)
	) name1294 (
		_w1762_,
		_w1826_,
		_w1827_
	);
	LUT4 #(
		.INIT('h004f)
	) name1295 (
		_w1821_,
		_w1823_,
		_w1824_,
		_w1827_,
		_w1828_
	);
	LUT3 #(
		.INIT('he0)
	) name1296 (
		\sa21_reg[1]/P0001 ,
		_w1819_,
		_w1828_,
		_w1829_
	);
	LUT4 #(
		.INIT('h0100)
	) name1297 (
		_w1796_,
		_w1787_,
		_w1813_,
		_w1829_,
		_w1830_
	);
	LUT3 #(
		.INIT('h69)
	) name1298 (
		\u0_w_reg[3][7]/P0001 ,
		_w1759_,
		_w1830_,
		_w1831_
	);
	LUT3 #(
		.INIT('h82)
	) name1299 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[7]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w1832_
	);
	LUT4 #(
		.INIT('h00eb)
	) name1300 (
		\ld_r_reg/P0001 ,
		_w1686_,
		_w1831_,
		_w1832_,
		_w1833_
	);
	LUT3 #(
		.INIT('h02)
	) name1301 (
		\sa10_reg[2]/P0001 ,
		_w1281_,
		_w1590_,
		_w1834_
	);
	LUT2 #(
		.INIT('h8)
	) name1302 (
		_w1238_,
		_w1286_,
		_w1835_
	);
	LUT4 #(
		.INIT('h0515)
	) name1303 (
		_w1236_,
		_w1238_,
		_w1286_,
		_w1271_,
		_w1836_
	);
	LUT4 #(
		.INIT('h2000)
	) name1304 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1837_
	);
	LUT2 #(
		.INIT('h8)
	) name1305 (
		\sa10_reg[5]/P0001 ,
		_w1837_,
		_w1838_
	);
	LUT4 #(
		.INIT('h1000)
	) name1306 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1839_
	);
	LUT3 #(
		.INIT('h01)
	) name1307 (
		\sa10_reg[2]/P0001 ,
		_w1556_,
		_w1839_,
		_w1840_
	);
	LUT4 #(
		.INIT('h7077)
	) name1308 (
		_w1834_,
		_w1836_,
		_w1838_,
		_w1840_,
		_w1841_
	);
	LUT2 #(
		.INIT('h4)
	) name1309 (
		\sa10_reg[4]/P0001 ,
		_w1236_,
		_w1842_
	);
	LUT4 #(
		.INIT('h0145)
	) name1310 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1236_,
		_w1281_,
		_w1843_
	);
	LUT4 #(
		.INIT('h0020)
	) name1311 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1844_
	);
	LUT2 #(
		.INIT('h8)
	) name1312 (
		\sa10_reg[4]/P0001 ,
		_w1844_,
		_w1845_
	);
	LUT3 #(
		.INIT('h2a)
	) name1313 (
		\sa10_reg[1]/P0001 ,
		_w1235_,
		_w1269_,
		_w1846_
	);
	LUT2 #(
		.INIT('h4)
	) name1314 (
		_w1845_,
		_w1846_,
		_w1847_
	);
	LUT3 #(
		.INIT('h0b)
	) name1315 (
		_w1841_,
		_w1843_,
		_w1847_,
		_w1848_
	);
	LUT3 #(
		.INIT('h80)
	) name1316 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1849_
	);
	LUT4 #(
		.INIT('h8000)
	) name1317 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1850_
	);
	LUT4 #(
		.INIT('hc840)
	) name1318 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		_w1577_,
		_w1849_,
		_w1851_
	);
	LUT2 #(
		.INIT('h4)
	) name1319 (
		\sa10_reg[4]/P0001 ,
		_w1252_,
		_w1852_
	);
	LUT3 #(
		.INIT('h23)
	) name1320 (
		\sa10_reg[5]/P0001 ,
		_w1289_,
		_w1318_,
		_w1853_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name1321 (
		\sa10_reg[4]/P0001 ,
		_w1256_,
		_w1238_,
		_w1266_,
		_w1854_
	);
	LUT4 #(
		.INIT('hba00)
	) name1322 (
		\sa10_reg[2]/P0001 ,
		_w1852_,
		_w1853_,
		_w1854_,
		_w1855_
	);
	LUT3 #(
		.INIT('h31)
	) name1323 (
		\sa10_reg[1]/P0001 ,
		_w1851_,
		_w1855_,
		_w1856_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name1324 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1857_
	);
	LUT2 #(
		.INIT('h1)
	) name1325 (
		\sa10_reg[2]/P0001 ,
		_w1857_,
		_w1858_
	);
	LUT2 #(
		.INIT('h4)
	) name1326 (
		\sa10_reg[7]/NET0131 ,
		_w1287_,
		_w1859_
	);
	LUT4 #(
		.INIT('h0200)
	) name1327 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1860_
	);
	LUT4 #(
		.INIT('h002a)
	) name1328 (
		\sa10_reg[1]/P0001 ,
		_w1234_,
		_w1311_,
		_w1860_,
		_w1861_
	);
	LUT3 #(
		.INIT('h10)
	) name1329 (
		_w1859_,
		_w1858_,
		_w1861_,
		_w1862_
	);
	LUT3 #(
		.INIT('h15)
	) name1330 (
		\sa10_reg[1]/P0001 ,
		_w1262_,
		_w1308_,
		_w1863_
	);
	LUT2 #(
		.INIT('h8)
	) name1331 (
		_w1278_,
		_w1567_,
		_w1864_
	);
	LUT4 #(
		.INIT('h1000)
	) name1332 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1865_
	);
	LUT3 #(
		.INIT('h80)
	) name1333 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1866_
	);
	LUT3 #(
		.INIT('h01)
	) name1334 (
		_w1837_,
		_w1866_,
		_w1865_,
		_w1867_
	);
	LUT3 #(
		.INIT('h20)
	) name1335 (
		_w1863_,
		_w1864_,
		_w1867_,
		_w1868_
	);
	LUT2 #(
		.INIT('h2)
	) name1336 (
		\sa10_reg[2]/P0001 ,
		_w1256_,
		_w1869_
	);
	LUT3 #(
		.INIT('h02)
	) name1337 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1870_
	);
	LUT3 #(
		.INIT('h01)
	) name1338 (
		_w1284_,
		_w1300_,
		_w1870_,
		_w1871_
	);
	LUT4 #(
		.INIT('h0020)
	) name1339 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1872_
	);
	LUT4 #(
		.INIT('h2000)
	) name1340 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1873_
	);
	LUT3 #(
		.INIT('h01)
	) name1341 (
		\sa10_reg[2]/P0001 ,
		_w1873_,
		_w1872_,
		_w1874_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name1342 (
		_w1319_,
		_w1869_,
		_w1871_,
		_w1874_,
		_w1875_
	);
	LUT4 #(
		.INIT('haa02)
	) name1343 (
		\sa10_reg[0]/P0001 ,
		_w1862_,
		_w1868_,
		_w1875_,
		_w1876_
	);
	LUT2 #(
		.INIT('h1)
	) name1344 (
		\sa10_reg[1]/P0001 ,
		_w1850_,
		_w1877_
	);
	LUT4 #(
		.INIT('hf351)
	) name1345 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		_w1878_
	);
	LUT4 #(
		.INIT('h5f13)
	) name1346 (
		\sa10_reg[5]/P0001 ,
		_w1234_,
		_w1591_,
		_w1878_,
		_w1879_
	);
	LUT2 #(
		.INIT('h8)
	) name1347 (
		_w1877_,
		_w1879_,
		_w1880_
	);
	LUT4 #(
		.INIT('h0100)
	) name1348 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1881_
	);
	LUT4 #(
		.INIT('h5510)
	) name1349 (
		\sa10_reg[2]/P0001 ,
		_w1224_,
		_w1294_,
		_w1881_,
		_w1882_
	);
	LUT3 #(
		.INIT('h20)
	) name1350 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1883_
	);
	LUT2 #(
		.INIT('h8)
	) name1351 (
		_w1277_,
		_w1883_,
		_w1884_
	);
	LUT3 #(
		.INIT('h08)
	) name1352 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1885_
	);
	LUT4 #(
		.INIT('h0080)
	) name1353 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1886_
	);
	LUT3 #(
		.INIT('h02)
	) name1354 (
		\sa10_reg[1]/P0001 ,
		_w1253_,
		_w1886_,
		_w1887_
	);
	LUT3 #(
		.INIT('h10)
	) name1355 (
		_w1884_,
		_w1882_,
		_w1887_,
		_w1888_
	);
	LUT4 #(
		.INIT('h2000)
	) name1356 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1889_
	);
	LUT4 #(
		.INIT('h0200)
	) name1357 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1890_
	);
	LUT4 #(
		.INIT('h0023)
	) name1358 (
		\sa10_reg[2]/P0001 ,
		_w1582_,
		_w1889_,
		_w1890_,
		_w1891_
	);
	LUT3 #(
		.INIT('h20)
	) name1359 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1242_,
		_w1892_
	);
	LUT3 #(
		.INIT('h0e)
	) name1360 (
		\sa10_reg[3]/P0001 ,
		_w1891_,
		_w1892_,
		_w1893_
	);
	LUT4 #(
		.INIT('h0155)
	) name1361 (
		\sa10_reg[0]/P0001 ,
		_w1880_,
		_w1888_,
		_w1893_,
		_w1894_
	);
	LUT4 #(
		.INIT('h0100)
	) name1362 (
		_w1848_,
		_w1876_,
		_w1894_,
		_w1856_,
		_w1895_
	);
	LUT3 #(
		.INIT('h20)
	) name1363 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1896_
	);
	LUT4 #(
		.INIT('h0100)
	) name1364 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1897_
	);
	LUT4 #(
		.INIT('h5510)
	) name1365 (
		\sa03_reg[2]/P0001 ,
		_w1059_,
		_w1896_,
		_w1897_,
		_w1898_
	);
	LUT2 #(
		.INIT('h8)
	) name1366 (
		_w1110_,
		_w1124_,
		_w1899_
	);
	LUT4 #(
		.INIT('h0080)
	) name1367 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1900_
	);
	LUT3 #(
		.INIT('h02)
	) name1368 (
		\sa03_reg[1]/P0001 ,
		_w1130_,
		_w1900_,
		_w1901_
	);
	LUT3 #(
		.INIT('h10)
	) name1369 (
		_w1898_,
		_w1899_,
		_w1901_,
		_w1902_
	);
	LUT4 #(
		.INIT('hfda8)
	) name1370 (
		\sa03_reg[2]/P0001 ,
		_w1079_,
		_w1644_,
		_w1676_,
		_w1903_
	);
	LUT2 #(
		.INIT('h1)
	) name1371 (
		\sa03_reg[1]/P0001 ,
		_w1193_,
		_w1904_
	);
	LUT2 #(
		.INIT('h4)
	) name1372 (
		_w1903_,
		_w1904_,
		_w1905_
	);
	LUT4 #(
		.INIT('h0100)
	) name1373 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w1906_
	);
	LUT4 #(
		.INIT('haa80)
	) name1374 (
		\sa03_reg[2]/P0001 ,
		_w1116_,
		_w1620_,
		_w1906_,
		_w1907_
	);
	LUT2 #(
		.INIT('h4)
	) name1375 (
		\sa03_reg[2]/P0001 ,
		_w1049_,
		_w1908_
	);
	LUT4 #(
		.INIT('h3310)
	) name1376 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1049_,
		_w1145_,
		_w1909_
	);
	LUT2 #(
		.INIT('h1)
	) name1377 (
		_w1907_,
		_w1909_,
		_w1910_
	);
	LUT4 #(
		.INIT('h0155)
	) name1378 (
		\sa03_reg[0]/P0001 ,
		_w1902_,
		_w1905_,
		_w1910_,
		_w1911_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name1379 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1912_
	);
	LUT2 #(
		.INIT('h1)
	) name1380 (
		\sa03_reg[2]/P0001 ,
		_w1912_,
		_w1913_
	);
	LUT4 #(
		.INIT('h0200)
	) name1381 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1914_
	);
	LUT4 #(
		.INIT('h002a)
	) name1382 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1145_,
		_w1914_,
		_w1915_
	);
	LUT3 #(
		.INIT('h10)
	) name1383 (
		_w1080_,
		_w1913_,
		_w1915_,
		_w1916_
	);
	LUT4 #(
		.INIT('h2000)
	) name1384 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1917_
	);
	LUT4 #(
		.INIT('h0015)
	) name1385 (
		\sa03_reg[1]/P0001 ,
		_w1623_,
		_w1620_,
		_w1917_,
		_w1918_
	);
	LUT2 #(
		.INIT('h8)
	) name1386 (
		_w1082_,
		_w1125_,
		_w1919_
	);
	LUT3 #(
		.INIT('h32)
	) name1387 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1920_
	);
	LUT4 #(
		.INIT('h7f33)
	) name1388 (
		\sa03_reg[4]/P0001 ,
		_w1081_,
		_w1125_,
		_w1920_,
		_w1921_
	);
	LUT2 #(
		.INIT('h8)
	) name1389 (
		_w1918_,
		_w1921_,
		_w1922_
	);
	LUT3 #(
		.INIT('h04)
	) name1390 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1923_
	);
	LUT4 #(
		.INIT('h0200)
	) name1391 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1924_
	);
	LUT3 #(
		.INIT('h01)
	) name1392 (
		_w1140_,
		_w1924_,
		_w1923_,
		_w1925_
	);
	LUT2 #(
		.INIT('h4)
	) name1393 (
		\sa03_reg[7]/NET0131 ,
		_w1187_,
		_w1926_
	);
	LUT3 #(
		.INIT('h01)
	) name1394 (
		\sa03_reg[2]/P0001 ,
		_w1048_,
		_w1185_,
		_w1927_
	);
	LUT4 #(
		.INIT('h7077)
	) name1395 (
		_w1192_,
		_w1925_,
		_w1926_,
		_w1927_,
		_w1928_
	);
	LUT4 #(
		.INIT('haa02)
	) name1396 (
		\sa03_reg[0]/P0001 ,
		_w1916_,
		_w1922_,
		_w1928_,
		_w1929_
	);
	LUT4 #(
		.INIT('h0084)
	) name1397 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1930_
	);
	LUT3 #(
		.INIT('h02)
	) name1398 (
		\sa03_reg[2]/P0001 ,
		_w1651_,
		_w1930_,
		_w1931_
	);
	LUT4 #(
		.INIT('h6fff)
	) name1399 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1072_,
		_w1932_
	);
	LUT2 #(
		.INIT('h8)
	) name1400 (
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1933_
	);
	LUT2 #(
		.INIT('h8)
	) name1401 (
		_w1060_,
		_w1933_,
		_w1934_
	);
	LUT3 #(
		.INIT('h01)
	) name1402 (
		\sa03_reg[2]/P0001 ,
		_w1099_,
		_w1624_,
		_w1935_
	);
	LUT4 #(
		.INIT('h7077)
	) name1403 (
		_w1931_,
		_w1932_,
		_w1934_,
		_w1935_,
		_w1936_
	);
	LUT2 #(
		.INIT('h4)
	) name1404 (
		\sa03_reg[3]/P0001 ,
		_w1145_,
		_w1937_
	);
	LUT3 #(
		.INIT('h15)
	) name1405 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[5]/P0001 ,
		_w1130_,
		_w1938_
	);
	LUT2 #(
		.INIT('h4)
	) name1406 (
		_w1937_,
		_w1938_,
		_w1939_
	);
	LUT3 #(
		.INIT('h07)
	) name1407 (
		_w1105_,
		_w1054_,
		_w1183_,
		_w1940_
	);
	LUT3 #(
		.INIT('h45)
	) name1408 (
		\sa03_reg[2]/P0001 ,
		_w1926_,
		_w1940_,
		_w1941_
	);
	LUT3 #(
		.INIT('h2a)
	) name1409 (
		\sa03_reg[1]/P0001 ,
		_w1050_,
		_w1175_,
		_w1942_
	);
	LUT2 #(
		.INIT('h8)
	) name1410 (
		_w1069_,
		_w1155_,
		_w1943_
	);
	LUT4 #(
		.INIT('h33bf)
	) name1411 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1140_,
		_w1657_,
		_w1944_
	);
	LUT3 #(
		.INIT('h40)
	) name1412 (
		_w1943_,
		_w1942_,
		_w1944_,
		_w1945_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1413 (
		_w1936_,
		_w1939_,
		_w1941_,
		_w1945_,
		_w1946_
	);
	LUT4 #(
		.INIT('hc840)
	) name1414 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1668_,
		_w1644_,
		_w1947_
	);
	LUT4 #(
		.INIT('h0001)
	) name1415 (
		_w1929_,
		_w1946_,
		_w1911_,
		_w1947_,
		_w1948_
	);
	LUT2 #(
		.INIT('h9)
	) name1416 (
		_w1895_,
		_w1948_,
		_w1949_
	);
	LUT3 #(
		.INIT('ha8)
	) name1417 (
		\sa10_reg[2]/P0001 ,
		_w1602_,
		_w1866_,
		_w1950_
	);
	LUT4 #(
		.INIT('h0010)
	) name1418 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1951_
	);
	LUT3 #(
		.INIT('h54)
	) name1419 (
		\sa10_reg[2]/P0001 ,
		_w1247_,
		_w1951_,
		_w1952_
	);
	LUT4 #(
		.INIT('h0400)
	) name1420 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1953_
	);
	LUT4 #(
		.INIT('h8000)
	) name1421 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1954_
	);
	LUT3 #(
		.INIT('h01)
	) name1422 (
		_w1839_,
		_w1954_,
		_w1953_,
		_w1955_
	);
	LUT4 #(
		.INIT('h0023)
	) name1423 (
		\sa10_reg[7]/NET0131 ,
		_w1220_,
		_w1297_,
		_w1615_,
		_w1956_
	);
	LUT4 #(
		.INIT('h1000)
	) name1424 (
		_w1950_,
		_w1952_,
		_w1955_,
		_w1956_,
		_w1957_
	);
	LUT4 #(
		.INIT('h0010)
	) name1425 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1958_
	);
	LUT3 #(
		.INIT('h32)
	) name1426 (
		_w1257_,
		_w1270_,
		_w1958_,
		_w1959_
	);
	LUT3 #(
		.INIT('h01)
	) name1427 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1960_
	);
	LUT2 #(
		.INIT('h1)
	) name1428 (
		_w1954_,
		_w1960_,
		_w1961_
	);
	LUT3 #(
		.INIT('h8a)
	) name1429 (
		\sa10_reg[2]/P0001 ,
		_w1959_,
		_w1961_,
		_w1962_
	);
	LUT4 #(
		.INIT('heffb)
	) name1430 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1963_
	);
	LUT4 #(
		.INIT('hfdf8)
	) name1431 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1964_
	);
	LUT4 #(
		.INIT('hf531)
	) name1432 (
		\sa10_reg[7]/NET0131 ,
		_w1315_,
		_w1963_,
		_w1964_,
		_w1965_
	);
	LUT3 #(
		.INIT('h23)
	) name1433 (
		\sa10_reg[2]/P0001 ,
		_w1258_,
		_w1244_,
		_w1966_
	);
	LUT4 #(
		.INIT('h3200)
	) name1434 (
		\sa10_reg[1]/P0001 ,
		_w1243_,
		_w1965_,
		_w1966_,
		_w1967_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1435 (
		\sa10_reg[1]/P0001 ,
		_w1957_,
		_w1962_,
		_w1967_,
		_w1968_
	);
	LUT4 #(
		.INIT('hfd3f)
	) name1436 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1969_
	);
	LUT2 #(
		.INIT('h1)
	) name1437 (
		\sa10_reg[2]/P0001 ,
		_w1969_,
		_w1970_
	);
	LUT2 #(
		.INIT('h8)
	) name1438 (
		_w1269_,
		_w1308_,
		_w1971_
	);
	LUT4 #(
		.INIT('h0007)
	) name1439 (
		\sa10_reg[4]/P0001 ,
		_w1252_,
		_w1281_,
		_w1890_,
		_w1972_
	);
	LUT4 #(
		.INIT('h5455)
	) name1440 (
		\sa10_reg[1]/P0001 ,
		_w1970_,
		_w1971_,
		_w1972_,
		_w1973_
	);
	LUT4 #(
		.INIT('h0123)
	) name1441 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1974_
	);
	LUT3 #(
		.INIT('ha8)
	) name1442 (
		\sa10_reg[1]/P0001 ,
		_w1311_,
		_w1974_,
		_w1975_
	);
	LUT3 #(
		.INIT('h04)
	) name1443 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1976_
	);
	LUT3 #(
		.INIT('h01)
	) name1444 (
		_w1281_,
		_w1872_,
		_w1976_,
		_w1977_
	);
	LUT3 #(
		.INIT('h45)
	) name1445 (
		\sa10_reg[2]/P0001 ,
		_w1975_,
		_w1977_,
		_w1978_
	);
	LUT4 #(
		.INIT('h0200)
	) name1446 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1979_
	);
	LUT3 #(
		.INIT('h07)
	) name1447 (
		_w1226_,
		_w1228_,
		_w1979_,
		_w1980_
	);
	LUT3 #(
		.INIT('h27)
	) name1448 (
		\sa10_reg[7]/NET0131 ,
		_w1247_,
		_w1287_,
		_w1981_
	);
	LUT3 #(
		.INIT('h2a)
	) name1449 (
		\sa10_reg[1]/P0001 ,
		_w1980_,
		_w1981_,
		_w1982_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name1450 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		_w1252_,
		_w1951_,
		_w1983_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name1451 (
		\sa10_reg[2]/P0001 ,
		_w1224_,
		_w1885_,
		_w1889_,
		_w1984_
	);
	LUT3 #(
		.INIT('hd0)
	) name1452 (
		\sa10_reg[2]/P0001 ,
		_w1983_,
		_w1984_,
		_w1985_
	);
	LUT4 #(
		.INIT('h0100)
	) name1453 (
		_w1978_,
		_w1982_,
		_w1973_,
		_w1985_,
		_w1986_
	);
	LUT3 #(
		.INIT('h6b)
	) name1454 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1987_
	);
	LUT3 #(
		.INIT('h20)
	) name1455 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1988_
	);
	LUT2 #(
		.INIT('h4)
	) name1456 (
		_w1987_,
		_w1988_,
		_w1989_
	);
	LUT3 #(
		.INIT('h13)
	) name1457 (
		_w1219_,
		_w1318_,
		_w1565_,
		_w1990_
	);
	LUT3 #(
		.INIT('h45)
	) name1458 (
		\sa10_reg[1]/P0001 ,
		_w1989_,
		_w1990_,
		_w1991_
	);
	LUT2 #(
		.INIT('h8)
	) name1459 (
		_w1277_,
		_w1602_,
		_w1992_
	);
	LUT4 #(
		.INIT('h23af)
	) name1460 (
		\sa10_reg[2]/P0001 ,
		_w1255_,
		_w1244_,
		_w1960_,
		_w1993_
	);
	LUT3 #(
		.INIT('h8a)
	) name1461 (
		\sa10_reg[1]/P0001 ,
		_w1992_,
		_w1993_,
		_w1994_
	);
	LUT2 #(
		.INIT('h1)
	) name1462 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[2]/P0001 ,
		_w1995_
	);
	LUT4 #(
		.INIT('h1000)
	) name1463 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1996_
	);
	LUT4 #(
		.INIT('h0007)
	) name1464 (
		\sa10_reg[4]/P0001 ,
		_w1281_,
		_w1889_,
		_w1996_,
		_w1997_
	);
	LUT3 #(
		.INIT('h80)
	) name1465 (
		\sa10_reg[5]/P0001 ,
		_w1269_,
		_w1308_,
		_w1998_
	);
	LUT4 #(
		.INIT('h5540)
	) name1466 (
		\sa10_reg[2]/P0001 ,
		_w1234_,
		_w1311_,
		_w1839_,
		_w1999_
	);
	LUT4 #(
		.INIT('h1101)
	) name1467 (
		_w1998_,
		_w1999_,
		_w1995_,
		_w1997_,
		_w2000_
	);
	LUT3 #(
		.INIT('h10)
	) name1468 (
		_w1991_,
		_w1994_,
		_w2000_,
		_w2001_
	);
	LUT4 #(
		.INIT('hd800)
	) name1469 (
		\sa10_reg[0]/P0001 ,
		_w1986_,
		_w1968_,
		_w2001_,
		_w2002_
	);
	LUT4 #(
		.INIT('h0008)
	) name1470 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2003_
	);
	LUT3 #(
		.INIT('ha8)
	) name1471 (
		\sa21_reg[2]/P0001 ,
		_w1345_,
		_w2003_,
		_w2004_
	);
	LUT2 #(
		.INIT('h8)
	) name1472 (
		_w1425_,
		_w1781_,
		_w2005_
	);
	LUT4 #(
		.INIT('h0007)
	) name1473 (
		_w1360_,
		_w1365_,
		_w1794_,
		_w1763_,
		_w2006_
	);
	LUT4 #(
		.INIT('h5455)
	) name1474 (
		\sa21_reg[1]/P0001 ,
		_w2004_,
		_w2005_,
		_w2006_,
		_w2007_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1475 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2008_
	);
	LUT3 #(
		.INIT('h8a)
	) name1476 (
		\sa21_reg[1]/P0001 ,
		_w1420_,
		_w2008_,
		_w2009_
	);
	LUT4 #(
		.INIT('h0020)
	) name1477 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2010_
	);
	LUT3 #(
		.INIT('h01)
	) name1478 (
		_w1426_,
		_w1794_,
		_w2010_,
		_w2011_
	);
	LUT3 #(
		.INIT('h45)
	) name1479 (
		\sa21_reg[2]/P0001 ,
		_w2009_,
		_w2011_,
		_w2012_
	);
	LUT4 #(
		.INIT('h0777)
	) name1480 (
		_w1348_,
		_w1350_,
		_w1334_,
		_w1360_,
		_w2013_
	);
	LUT3 #(
		.INIT('h20)
	) name1481 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2014_
	);
	LUT4 #(
		.INIT('h0200)
	) name1482 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2015_
	);
	LUT3 #(
		.INIT('h07)
	) name1483 (
		_w1327_,
		_w1398_,
		_w2015_,
		_w2016_
	);
	LUT3 #(
		.INIT('h2a)
	) name1484 (
		\sa21_reg[1]/P0001 ,
		_w2013_,
		_w2016_,
		_w2017_
	);
	LUT4 #(
		.INIT('h0010)
	) name1485 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2018_
	);
	LUT4 #(
		.INIT('h8cbf)
	) name1486 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w1365_,
		_w2018_,
		_w2019_
	);
	LUT3 #(
		.INIT('h02)
	) name1487 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w2020_
	);
	LUT4 #(
		.INIT('h135f)
	) name1488 (
		_w1391_,
		_w1378_,
		_w1765_,
		_w2020_,
		_w2021_
	);
	LUT3 #(
		.INIT('hd0)
	) name1489 (
		\sa21_reg[2]/P0001 ,
		_w2019_,
		_w2021_,
		_w2022_
	);
	LUT4 #(
		.INIT('h0100)
	) name1490 (
		_w2012_,
		_w2007_,
		_w2017_,
		_w2022_,
		_w2023_
	);
	LUT4 #(
		.INIT('h0010)
	) name1491 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2024_
	);
	LUT4 #(
		.INIT('h5554)
	) name1492 (
		\sa21_reg[2]/P0001 ,
		_w1361_,
		_w2014_,
		_w2024_,
		_w2025_
	);
	LUT3 #(
		.INIT('ha8)
	) name1493 (
		\sa21_reg[2]/P0001 ,
		_w1352_,
		_w1777_,
		_w2026_
	);
	LUT4 #(
		.INIT('hf3bf)
	) name1494 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2027_
	);
	LUT4 #(
		.INIT('h1000)
	) name1495 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2028_
	);
	LUT4 #(
		.INIT('heffd)
	) name1496 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2029_
	);
	LUT4 #(
		.INIT('h7200)
	) name1497 (
		\sa21_reg[4]/P0001 ,
		_w1352_,
		_w2027_,
		_w2029_,
		_w2030_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1498 (
		\sa21_reg[1]/P0001 ,
		_w2026_,
		_w2025_,
		_w2030_,
		_w2031_
	);
	LUT3 #(
		.INIT('h54)
	) name1499 (
		\sa21_reg[3]/P0001 ,
		_w1792_,
		_w1804_,
		_w2032_
	);
	LUT2 #(
		.INIT('h8)
	) name1500 (
		_w1385_,
		_w1378_,
		_w2033_
	);
	LUT2 #(
		.INIT('h2)
	) name1501 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w2034_
	);
	LUT3 #(
		.INIT('h02)
	) name1502 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w2035_
	);
	LUT4 #(
		.INIT('h0777)
	) name1503 (
		_w1385_,
		_w1378_,
		_w2034_,
		_w2035_,
		_w2036_
	);
	LUT3 #(
		.INIT('h45)
	) name1504 (
		\sa21_reg[1]/P0001 ,
		_w2032_,
		_w2036_,
		_w2037_
	);
	LUT4 #(
		.INIT('h8002)
	) name1505 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w2038_
	);
	LUT3 #(
		.INIT('h01)
	) name1506 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2039_
	);
	LUT3 #(
		.INIT('h04)
	) name1507 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w2040_
	);
	LUT4 #(
		.INIT('h0103)
	) name1508 (
		_w1336_,
		_w2039_,
		_w2038_,
		_w2040_,
		_w2041_
	);
	LUT3 #(
		.INIT('h13)
	) name1509 (
		_w1334_,
		_w1368_,
		_w1765_,
		_w2042_
	);
	LUT4 #(
		.INIT('he400)
	) name1510 (
		\sa21_reg[2]/P0001 ,
		_w1340_,
		_w2041_,
		_w2042_,
		_w2043_
	);
	LUT3 #(
		.INIT('h10)
	) name1511 (
		_w2031_,
		_w2037_,
		_w2043_,
		_w2044_
	);
	LUT4 #(
		.INIT('hee7f)
	) name1512 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2045_
	);
	LUT4 #(
		.INIT('h5054)
	) name1513 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[5]/P0001 ,
		_w1395_,
		_w2045_,
		_w2046_
	);
	LUT4 #(
		.INIT('h1445)
	) name1514 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2047_
	);
	LUT2 #(
		.INIT('h8)
	) name1515 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w2048_
	);
	LUT3 #(
		.INIT('ha2)
	) name1516 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w2049_
	);
	LUT4 #(
		.INIT('h5551)
	) name1517 (
		_w1422_,
		_w2048_,
		_w2049_,
		_w2047_,
		_w2050_
	);
	LUT3 #(
		.INIT('h45)
	) name1518 (
		\sa21_reg[1]/P0001 ,
		_w2046_,
		_w2050_,
		_w2051_
	);
	LUT2 #(
		.INIT('h8)
	) name1519 (
		_w1375_,
		_w1777_,
		_w2052_
	);
	LUT4 #(
		.INIT('h153f)
	) name1520 (
		_w1334_,
		_w1394_,
		_w1380_,
		_w1765_,
		_w2053_
	);
	LUT3 #(
		.INIT('h8a)
	) name1521 (
		\sa21_reg[1]/P0001 ,
		_w2052_,
		_w2053_,
		_w2054_
	);
	LUT2 #(
		.INIT('h8)
	) name1522 (
		_w1350_,
		_w1387_,
		_w2055_
	);
	LUT4 #(
		.INIT('h135f)
	) name1523 (
		_w1350_,
		_w1357_,
		_w1387_,
		_w1390_,
		_w2056_
	);
	LUT2 #(
		.INIT('h4)
	) name1524 (
		_w1428_,
		_w2056_,
		_w2057_
	);
	LUT3 #(
		.INIT('h10)
	) name1525 (
		_w2051_,
		_w2054_,
		_w2057_,
		_w2058_
	);
	LUT4 #(
		.INIT('he400)
	) name1526 (
		\sa21_reg[0]/P0001 ,
		_w2044_,
		_w2023_,
		_w2058_,
		_w2059_
	);
	LUT2 #(
		.INIT('h9)
	) name1527 (
		_w2002_,
		_w2059_,
		_w2060_
	);
	LUT3 #(
		.INIT('h65)
	) name1528 (
		\u0_w_reg[3][29]/P0001 ,
		_w1497_,
		_w1552_,
		_w2061_
	);
	LUT4 #(
		.INIT('h4114)
	) name1529 (
		\ld_r_reg/P0001 ,
		_w1949_,
		_w2060_,
		_w2061_,
		_w2062_
	);
	LUT3 #(
		.INIT('h28)
	) name1530 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[29]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		_w2063_
	);
	LUT2 #(
		.INIT('he)
	) name1531 (
		_w2062_,
		_w2063_,
		_w2064_
	);
	LUT2 #(
		.INIT('h9)
	) name1532 (
		_w1323_,
		_w1438_,
		_w2065_
	);
	LUT4 #(
		.INIT('h5655)
	) name1533 (
		\u0_w_reg[3][30]/P0001 ,
		_w1707_,
		_w1732_,
		_w1758_,
		_w2066_
	);
	LUT3 #(
		.INIT('h96)
	) name1534 (
		_w1149_,
		_w2002_,
		_w2066_,
		_w2067_
	);
	LUT3 #(
		.INIT('h82)
	) name1535 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[30]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w2068_
	);
	LUT4 #(
		.INIT('h00eb)
	) name1536 (
		\ld_r_reg/P0001 ,
		_w2065_,
		_w2067_,
		_w2068_,
		_w2069_
	);
	LUT2 #(
		.INIT('h4)
	) name1537 (
		\sa21_reg[2]/P0001 ,
		_w2003_,
		_w2070_
	);
	LUT2 #(
		.INIT('h8)
	) name1538 (
		_w1334_,
		_w2048_,
		_w2071_
	);
	LUT3 #(
		.INIT('h32)
	) name1539 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w2072_
	);
	LUT4 #(
		.INIT('h2000)
	) name1540 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2073_
	);
	LUT3 #(
		.INIT('h0d)
	) name1541 (
		_w1351_,
		_w2072_,
		_w2073_,
		_w2074_
	);
	LUT4 #(
		.INIT('h5455)
	) name1542 (
		\sa21_reg[1]/P0001 ,
		_w2070_,
		_w2071_,
		_w2074_,
		_w2075_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name1543 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2076_
	);
	LUT2 #(
		.INIT('h1)
	) name1544 (
		\sa21_reg[2]/P0001 ,
		_w2076_,
		_w2077_
	);
	LUT2 #(
		.INIT('h8)
	) name1545 (
		_w1401_,
		_w1420_,
		_w2078_
	);
	LUT4 #(
		.INIT('h0200)
	) name1546 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2079_
	);
	LUT3 #(
		.INIT('h07)
	) name1547 (
		_w1327_,
		_w1398_,
		_w2079_,
		_w2080_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1548 (
		\sa21_reg[1]/P0001 ,
		_w2077_,
		_w2078_,
		_w2080_,
		_w2081_
	);
	LUT4 #(
		.INIT('h35f5)
	) name1549 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2082_
	);
	LUT2 #(
		.INIT('h1)
	) name1550 (
		\sa21_reg[4]/P0001 ,
		_w2082_,
		_w2083_
	);
	LUT3 #(
		.INIT('h02)
	) name1551 (
		\sa21_reg[2]/P0001 ,
		_w1370_,
		_w2040_,
		_w2084_
	);
	LUT4 #(
		.INIT('h2000)
	) name1552 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2085_
	);
	LUT3 #(
		.INIT('h01)
	) name1553 (
		\sa21_reg[2]/P0001 ,
		_w2010_,
		_w2085_,
		_w2086_
	);
	LUT4 #(
		.INIT('h8acf)
	) name1554 (
		_w1434_,
		_w2083_,
		_w2084_,
		_w2086_,
		_w2087_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1555 (
		\sa21_reg[0]/P0001 ,
		_w2081_,
		_w2075_,
		_w2087_,
		_w2088_
	);
	LUT4 #(
		.INIT('h0100)
	) name1556 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2089_
	);
	LUT4 #(
		.INIT('h5504)
	) name1557 (
		\sa21_reg[2]/P0001 ,
		_w1334_,
		_w1419_,
		_w2089_,
		_w2090_
	);
	LUT4 #(
		.INIT('h0080)
	) name1558 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2091_
	);
	LUT4 #(
		.INIT('h0015)
	) name1559 (
		_w1364_,
		_w1375_,
		_w1800_,
		_w2091_,
		_w2092_
	);
	LUT3 #(
		.INIT('h8a)
	) name1560 (
		\sa21_reg[1]/P0001 ,
		_w2090_,
		_w2092_,
		_w2093_
	);
	LUT4 #(
		.INIT('h0200)
	) name1561 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w2094_
	);
	LUT4 #(
		.INIT('h0013)
	) name1562 (
		_w1391_,
		_w1427_,
		_w1765_,
		_w2094_,
		_w2095_
	);
	LUT2 #(
		.INIT('h1)
	) name1563 (
		\sa21_reg[3]/P0001 ,
		_w2095_,
		_w2096_
	);
	LUT4 #(
		.INIT('h0002)
	) name1564 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2097_
	);
	LUT4 #(
		.INIT('h5540)
	) name1565 (
		\sa21_reg[1]/P0001 ,
		\sa21_reg[5]/P0001 ,
		_w1761_,
		_w2097_,
		_w2098_
	);
	LUT4 #(
		.INIT('h22af)
	) name1566 (
		\sa21_reg[1]/P0001 ,
		_w1330_,
		_w1379_,
		_w1803_,
		_w2099_
	);
	LUT3 #(
		.INIT('h31)
	) name1567 (
		\sa21_reg[2]/P0001 ,
		_w2098_,
		_w2099_,
		_w2100_
	);
	LUT4 #(
		.INIT('h5455)
	) name1568 (
		\sa21_reg[0]/P0001 ,
		_w2096_,
		_w2093_,
		_w2100_,
		_w2101_
	);
	LUT4 #(
		.INIT('h0084)
	) name1569 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2102_
	);
	LUT2 #(
		.INIT('h8)
	) name1570 (
		_w1330_,
		_w1781_,
		_w2103_
	);
	LUT3 #(
		.INIT('h07)
	) name1571 (
		_w1344_,
		_w1394_,
		_w1760_,
		_w2104_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1572 (
		\sa21_reg[2]/P0001 ,
		_w2102_,
		_w2103_,
		_w2104_,
		_w2105_
	);
	LUT2 #(
		.INIT('h8)
	) name1573 (
		_w1390_,
		_w1420_,
		_w2106_
	);
	LUT4 #(
		.INIT('h0007)
	) name1574 (
		_w1390_,
		_w1420_,
		_w1820_,
		_w2028_,
		_w2107_
	);
	LUT3 #(
		.INIT('h01)
	) name1575 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w2108_
	);
	LUT2 #(
		.INIT('h8)
	) name1576 (
		_w1326_,
		_w2108_,
		_w2109_
	);
	LUT4 #(
		.INIT('h153f)
	) name1577 (
		_w1326_,
		_w1379_,
		_w1380_,
		_w2108_,
		_w2110_
	);
	LUT3 #(
		.INIT('he0)
	) name1578 (
		\sa21_reg[2]/P0001 ,
		_w2107_,
		_w2110_,
		_w2111_
	);
	LUT3 #(
		.INIT('h45)
	) name1579 (
		\sa21_reg[1]/P0001 ,
		_w2105_,
		_w2111_,
		_w2112_
	);
	LUT3 #(
		.INIT('h07)
	) name1580 (
		_w1327_,
		_w1394_,
		_w1402_,
		_w2113_
	);
	LUT3 #(
		.INIT('h45)
	) name1581 (
		\sa21_reg[2]/P0001 ,
		_w2033_,
		_w2113_,
		_w2114_
	);
	LUT2 #(
		.INIT('h4)
	) name1582 (
		\sa21_reg[5]/P0001 ,
		_w2015_,
		_w2115_
	);
	LUT2 #(
		.INIT('h8)
	) name1583 (
		_w1346_,
		_w1375_,
		_w2116_
	);
	LUT4 #(
		.INIT('h135f)
	) name1584 (
		_w1349_,
		_w1330_,
		_w1387_,
		_w1391_,
		_w2117_
	);
	LUT3 #(
		.INIT('h10)
	) name1585 (
		_w2116_,
		_w2115_,
		_w2117_,
		_w2118_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name1586 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		_w1379_,
		_w1788_,
		_w2119_
	);
	LUT4 #(
		.INIT('h7500)
	) name1587 (
		\sa21_reg[1]/P0001 ,
		_w2114_,
		_w2118_,
		_w2119_,
		_w2120_
	);
	LUT4 #(
		.INIT('h0100)
	) name1588 (
		_w2101_,
		_w2088_,
		_w2112_,
		_w2120_,
		_w2121_
	);
	LUT3 #(
		.INIT('h69)
	) name1589 (
		_w1149_,
		_w1895_,
		_w2121_,
		_w2122_
	);
	LUT4 #(
		.INIT('h9a65)
	) name1590 (
		\u0_w_reg[3][21]/P0001 ,
		_w1497_,
		_w1552_,
		_w2059_,
		_w2123_
	);
	LUT3 #(
		.INIT('h82)
	) name1591 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[21]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		_w2124_
	);
	LUT4 #(
		.INIT('h00eb)
	) name1592 (
		\ld_r_reg/P0001 ,
		_w2122_,
		_w2123_,
		_w2124_,
		_w2125_
	);
	LUT3 #(
		.INIT('h69)
	) name1593 (
		_w1214_,
		_w2002_,
		_w2059_,
		_w2126_
	);
	LUT4 #(
		.INIT('h5655)
	) name1594 (
		\u0_w_reg[3][22]/P0001 ,
		_w1707_,
		_w1732_,
		_w1758_,
		_w2127_
	);
	LUT2 #(
		.INIT('h6)
	) name1595 (
		_w1438_,
		_w2127_,
		_w2128_
	);
	LUT3 #(
		.INIT('h82)
	) name1596 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[22]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w2129_
	);
	LUT4 #(
		.INIT('h00eb)
	) name1597 (
		\ld_r_reg/P0001 ,
		_w2126_,
		_w2128_,
		_w2129_,
		_w2130_
	);
	LUT3 #(
		.INIT('h96)
	) name1598 (
		_w1149_,
		_w2002_,
		_w2121_,
		_w2131_
	);
	LUT4 #(
		.INIT('h0020)
	) name1599 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w2132_
	);
	LUT3 #(
		.INIT('h02)
	) name1600 (
		\sa32_reg[2]/P0001 ,
		_w1503_,
		_w2132_,
		_w2133_
	);
	LUT2 #(
		.INIT('h9)
	) name1601 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w2134_
	);
	LUT3 #(
		.INIT('h13)
	) name1602 (
		_w1536_,
		_w1687_,
		_w2134_,
		_w2135_
	);
	LUT2 #(
		.INIT('h4)
	) name1603 (
		_w1482_,
		_w1524_,
		_w2136_
	);
	LUT3 #(
		.INIT('h15)
	) name1604 (
		\sa32_reg[2]/P0001 ,
		_w1467_,
		_w1475_,
		_w2137_
	);
	LUT4 #(
		.INIT('h7077)
	) name1605 (
		_w2133_,
		_w2135_,
		_w2136_,
		_w2137_,
		_w2138_
	);
	LUT2 #(
		.INIT('h8)
	) name1606 (
		_w1444_,
		_w1746_,
		_w2139_
	);
	LUT4 #(
		.INIT('h1d3f)
	) name1607 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1521_,
		_w1746_,
		_w2140_
	);
	LUT3 #(
		.INIT('h45)
	) name1608 (
		\sa32_reg[1]/P0001 ,
		_w2138_,
		_w2140_,
		_w2141_
	);
	LUT3 #(
		.INIT('h07)
	) name1609 (
		_w1460_,
		_w1746_,
		_w1710_,
		_w2142_
	);
	LUT3 #(
		.INIT('h45)
	) name1610 (
		\sa32_reg[2]/P0001 ,
		_w1477_,
		_w2142_,
		_w2143_
	);
	LUT2 #(
		.INIT('h4)
	) name1611 (
		\sa32_reg[5]/P0001 ,
		_w1518_,
		_w2144_
	);
	LUT2 #(
		.INIT('h8)
	) name1612 (
		\sa32_reg[3]/P0001 ,
		_w1527_,
		_w2145_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name1613 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		_w1547_,
		_w1693_,
		_w2146_
	);
	LUT3 #(
		.INIT('h10)
	) name1614 (
		_w2144_,
		_w2145_,
		_w2146_,
		_w2147_
	);
	LUT3 #(
		.INIT('h80)
	) name1615 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w2148_
	);
	LUT4 #(
		.INIT('h135f)
	) name1616 (
		_w1489_,
		_w1546_,
		_w1748_,
		_w2148_,
		_w2149_
	);
	LUT4 #(
		.INIT('h7500)
	) name1617 (
		\sa32_reg[1]/P0001 ,
		_w2143_,
		_w2147_,
		_w2149_,
		_w2150_
	);
	LUT3 #(
		.INIT('h20)
	) name1618 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2151_
	);
	LUT3 #(
		.INIT('h10)
	) name1619 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w2152_
	);
	LUT4 #(
		.INIT('h0100)
	) name1620 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2153_
	);
	LUT4 #(
		.INIT('h5510)
	) name1621 (
		\sa32_reg[2]/P0001 ,
		_w1467_,
		_w2151_,
		_w2153_,
		_w2154_
	);
	LUT3 #(
		.INIT('h20)
	) name1622 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w2155_
	);
	LUT4 #(
		.INIT('h0111)
	) name1623 (
		_w1542_,
		_w1703_,
		_w1724_,
		_w2155_,
		_w2156_
	);
	LUT3 #(
		.INIT('h8a)
	) name1624 (
		\sa32_reg[1]/P0001 ,
		_w2154_,
		_w2156_,
		_w2157_
	);
	LUT4 #(
		.INIT('h1000)
	) name1625 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w2158_
	);
	LUT3 #(
		.INIT('h54)
	) name1626 (
		\sa32_reg[7]/P0001 ,
		_w1468_,
		_w2158_,
		_w2159_
	);
	LUT4 #(
		.INIT('h7f7c)
	) name1627 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2160_
	);
	LUT2 #(
		.INIT('h2)
	) name1628 (
		\sa32_reg[2]/P0001 ,
		_w2160_,
		_w2161_
	);
	LUT3 #(
		.INIT('h54)
	) name1629 (
		\sa32_reg[1]/P0001 ,
		_w2159_,
		_w2161_,
		_w2162_
	);
	LUT4 #(
		.INIT('haa20)
	) name1630 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[5]/P0001 ,
		_w1512_,
		_w1692_,
		_w2163_
	);
	LUT3 #(
		.INIT('h10)
	) name1631 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		_w1527_,
		_w2164_
	);
	LUT3 #(
		.INIT('h01)
	) name1632 (
		_w2139_,
		_w2164_,
		_w2163_,
		_w2165_
	);
	LUT4 #(
		.INIT('h5455)
	) name1633 (
		\sa32_reg[0]/P0002 ,
		_w2157_,
		_w2162_,
		_w2165_,
		_w2166_
	);
	LUT3 #(
		.INIT('h32)
	) name1634 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w2167_
	);
	LUT4 #(
		.INIT('h2000)
	) name1635 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2168_
	);
	LUT4 #(
		.INIT('h0051)
	) name1636 (
		\sa32_reg[1]/P0001 ,
		_w1447_,
		_w2167_,
		_w2168_,
		_w2169_
	);
	LUT3 #(
		.INIT('h1b)
	) name1637 (
		\sa32_reg[2]/P0001 ,
		_w1512_,
		_w1492_,
		_w2170_
	);
	LUT2 #(
		.INIT('h8)
	) name1638 (
		_w2169_,
		_w2170_,
		_w2171_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name1639 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2172_
	);
	LUT2 #(
		.INIT('h1)
	) name1640 (
		\sa32_reg[2]/P0001 ,
		_w2172_,
		_w2173_
	);
	LUT3 #(
		.INIT('h2a)
	) name1641 (
		\sa32_reg[1]/P0001 ,
		_w1506_,
		_w1468_,
		_w2174_
	);
	LUT4 #(
		.INIT('h0200)
	) name1642 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2175_
	);
	LUT3 #(
		.INIT('h07)
	) name1643 (
		_w1443_,
		_w1472_,
		_w2175_,
		_w2176_
	);
	LUT3 #(
		.INIT('h20)
	) name1644 (
		_w2174_,
		_w2173_,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h2)
	) name1645 (
		\sa32_reg[2]/P0001 ,
		_w1514_,
		_w2178_
	);
	LUT3 #(
		.INIT('h04)
	) name1646 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w2179_
	);
	LUT3 #(
		.INIT('h01)
	) name1647 (
		_w1468_,
		_w1740_,
		_w2179_,
		_w2180_
	);
	LUT4 #(
		.INIT('h2000)
	) name1648 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2181_
	);
	LUT3 #(
		.INIT('h01)
	) name1649 (
		\sa32_reg[2]/P0001 ,
		_w1505_,
		_w2181_,
		_w2182_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name1650 (
		_w1747_,
		_w2178_,
		_w2180_,
		_w2182_,
		_w2183_
	);
	LUT4 #(
		.INIT('haa02)
	) name1651 (
		\sa32_reg[0]/P0002 ,
		_w2171_,
		_w2177_,
		_w2183_,
		_w2184_
	);
	LUT4 #(
		.INIT('h0100)
	) name1652 (
		_w2141_,
		_w2166_,
		_w2184_,
		_w2150_,
		_w2185_
	);
	LUT4 #(
		.INIT('h9a65)
	) name1653 (
		\u0_w_reg[3][13]/P0001 ,
		_w1497_,
		_w1552_,
		_w2185_,
		_w2186_
	);
	LUT3 #(
		.INIT('h28)
	) name1654 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[13]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		_w2187_
	);
	LUT4 #(
		.INIT('hff14)
	) name1655 (
		\ld_r_reg/P0001 ,
		_w2131_,
		_w2186_,
		_w2187_,
		_w2188_
	);
	LUT3 #(
		.INIT('h96)
	) name1656 (
		_w1214_,
		_w1323_,
		_w2059_,
		_w2189_
	);
	LUT4 #(
		.INIT('h5655)
	) name1657 (
		\u0_w_reg[3][14]/P0001 ,
		_w1707_,
		_w1732_,
		_w1758_,
		_w2190_
	);
	LUT3 #(
		.INIT('hb4)
	) name1658 (
		_w1497_,
		_w1552_,
		_w2190_,
		_w2191_
	);
	LUT3 #(
		.INIT('h28)
	) name1659 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[14]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w2192_
	);
	LUT4 #(
		.INIT('hff14)
	) name1660 (
		\ld_r_reg/P0001 ,
		_w2189_,
		_w2191_,
		_w2192_,
		_w2193_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name1661 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2194_
	);
	LUT3 #(
		.INIT('h8a)
	) name1662 (
		\sa32_reg[2]/P0001 ,
		_w1473_,
		_w2194_,
		_w2195_
	);
	LUT3 #(
		.INIT('h80)
	) name1663 (
		\sa32_reg[4]/P0001 ,
		_w1536_,
		_w1698_,
		_w2196_
	);
	LUT3 #(
		.INIT('h8a)
	) name1664 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2197_
	);
	LUT4 #(
		.INIT('h0010)
	) name1665 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w2198_
	);
	LUT3 #(
		.INIT('h0d)
	) name1666 (
		_w1467_,
		_w2197_,
		_w2198_,
		_w2199_
	);
	LUT4 #(
		.INIT('h5455)
	) name1667 (
		\sa32_reg[1]/P0001 ,
		_w2196_,
		_w2195_,
		_w2199_,
		_w2200_
	);
	LUT3 #(
		.INIT('h07)
	) name1668 (
		\sa32_reg[7]/P0001 ,
		_w1445_,
		_w2153_,
		_w2201_
	);
	LUT3 #(
		.INIT('h2a)
	) name1669 (
		\sa32_reg[2]/P0001 ,
		_w1697_,
		_w2201_,
		_w2202_
	);
	LUT4 #(
		.INIT('h4041)
	) name1670 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2203_
	);
	LUT3 #(
		.INIT('ha8)
	) name1671 (
		\sa32_reg[1]/P0001 ,
		_w1734_,
		_w2203_,
		_w2204_
	);
	LUT4 #(
		.INIT('h8000)
	) name1672 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2205_
	);
	LUT4 #(
		.INIT('h0040)
	) name1673 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w2206_
	);
	LUT3 #(
		.INIT('h54)
	) name1674 (
		\sa32_reg[2]/P0001 ,
		_w2205_,
		_w2206_,
		_w2207_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name1675 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2208_
	);
	LUT4 #(
		.INIT('h0040)
	) name1676 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2209_
	);
	LUT3 #(
		.INIT('h0d)
	) name1677 (
		_w1487_,
		_w2208_,
		_w2209_,
		_w2210_
	);
	LUT4 #(
		.INIT('h0100)
	) name1678 (
		_w2144_,
		_w2204_,
		_w2207_,
		_w2210_,
		_w2211_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1679 (
		\sa32_reg[0]/P0002 ,
		_w2202_,
		_w2200_,
		_w2211_,
		_w2212_
	);
	LUT4 #(
		.INIT('h45cf)
	) name1680 (
		_w1444_,
		_w1457_,
		_w1440_,
		_w1746_,
		_w2213_
	);
	LUT2 #(
		.INIT('h1)
	) name1681 (
		\sa32_reg[2]/P0001 ,
		_w2213_,
		_w2214_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1682 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1741_,
		_w1713_,
		_w2215_
	);
	LUT4 #(
		.INIT('h0040)
	) name1683 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w2216_
	);
	LUT3 #(
		.INIT('h15)
	) name1684 (
		\sa32_reg[1]/P0001 ,
		_w1499_,
		_w2216_,
		_w2217_
	);
	LUT3 #(
		.INIT('h10)
	) name1685 (
		_w1548_,
		_w2215_,
		_w2217_,
		_w2218_
	);
	LUT4 #(
		.INIT('h5444)
	) name1686 (
		\sa32_reg[5]/P0001 ,
		_w1535_,
		_w1693_,
		_w1724_,
		_w2219_
	);
	LUT4 #(
		.INIT('h27af)
	) name1687 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		_w1510_,
		_w1536_,
		_w2220_
	);
	LUT3 #(
		.INIT('h20)
	) name1688 (
		_w2174_,
		_w2219_,
		_w2220_,
		_w2221_
	);
	LUT3 #(
		.INIT('h0b)
	) name1689 (
		_w2214_,
		_w2218_,
		_w2221_,
		_w2222_
	);
	LUT3 #(
		.INIT('hb9)
	) name1690 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2223_
	);
	LUT2 #(
		.INIT('h2)
	) name1691 (
		_w1467_,
		_w2223_,
		_w2224_
	);
	LUT3 #(
		.INIT('h40)
	) name1692 (
		\sa32_reg[1]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w2225_
	);
	LUT3 #(
		.INIT('h8a)
	) name1693 (
		\sa32_reg[2]/P0001 ,
		_w1504_,
		_w2225_,
		_w2226_
	);
	LUT3 #(
		.INIT('h80)
	) name1694 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2227_
	);
	LUT4 #(
		.INIT('h8000)
	) name1695 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2228_
	);
	LUT3 #(
		.INIT('h07)
	) name1696 (
		\sa32_reg[7]/P0001 ,
		_w1445_,
		_w2228_,
		_w2229_
	);
	LUT2 #(
		.INIT('h1)
	) name1697 (
		\sa32_reg[2]/P0001 ,
		_w1713_,
		_w2230_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name1698 (
		_w2224_,
		_w2226_,
		_w2229_,
		_w2230_,
		_w2231_
	);
	LUT2 #(
		.INIT('h8)
	) name1699 (
		\sa32_reg[3]/P0001 ,
		_w1542_,
		_w2232_
	);
	LUT4 #(
		.INIT('h8000)
	) name1700 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2233_
	);
	LUT4 #(
		.INIT('h0100)
	) name1701 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w2234_
	);
	LUT4 #(
		.INIT('h0007)
	) name1702 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2235_
	);
	LUT4 #(
		.INIT('h0002)
	) name1703 (
		\sa32_reg[1]/P0001 ,
		_w2233_,
		_w2234_,
		_w2235_,
		_w2236_
	);
	LUT4 #(
		.INIT('h0010)
	) name1704 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2237_
	);
	LUT4 #(
		.INIT('hbfef)
	) name1705 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2238_
	);
	LUT2 #(
		.INIT('h1)
	) name1706 (
		\sa32_reg[3]/P0001 ,
		_w2238_,
		_w2239_
	);
	LUT3 #(
		.INIT('h45)
	) name1707 (
		\sa32_reg[1]/P0001 ,
		\sa32_reg[2]/P0001 ,
		_w1512_,
		_w2240_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1708 (
		_w2232_,
		_w2236_,
		_w2239_,
		_w2240_,
		_w2241_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name1709 (
		\sa32_reg[2]/P0001 ,
		_w1463_,
		_w1542_,
		_w2233_,
		_w2242_
	);
	LUT4 #(
		.INIT('hab00)
	) name1710 (
		\sa32_reg[0]/P0002 ,
		_w2231_,
		_w2241_,
		_w2242_,
		_w2243_
	);
	LUT3 #(
		.INIT('h10)
	) name1711 (
		_w2212_,
		_w2222_,
		_w2243_,
		_w2244_
	);
	LUT3 #(
		.INIT('had)
	) name1712 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w2245_
	);
	LUT3 #(
		.INIT('hf6)
	) name1713 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2246_
	);
	LUT3 #(
		.INIT('h2a)
	) name1714 (
		\sa32_reg[2]/P0001 ,
		_w2245_,
		_w2246_,
		_w2247_
	);
	LUT4 #(
		.INIT('h2e3f)
	) name1715 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		_w1527_,
		_w1536_,
		_w2248_
	);
	LUT3 #(
		.INIT('h8a)
	) name1716 (
		\sa32_reg[1]/P0001 ,
		_w2247_,
		_w2248_,
		_w2249_
	);
	LUT3 #(
		.INIT('ha2)
	) name1717 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w2250_
	);
	LUT4 #(
		.INIT('h7d1d)
	) name1718 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2251_
	);
	LUT2 #(
		.INIT('h1)
	) name1719 (
		\sa32_reg[2]/P0001 ,
		_w2251_,
		_w2252_
	);
	LUT4 #(
		.INIT('h0100)
	) name1720 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w2253_
	);
	LUT2 #(
		.INIT('h8)
	) name1721 (
		\sa32_reg[2]/P0001 ,
		_w2253_,
		_w2254_
	);
	LUT3 #(
		.INIT('h0d)
	) name1722 (
		_w1440_,
		_w1737_,
		_w2132_,
		_w2255_
	);
	LUT4 #(
		.INIT('h5455)
	) name1723 (
		\sa32_reg[1]/P0001 ,
		_w2252_,
		_w2254_,
		_w2255_,
		_w2256_
	);
	LUT4 #(
		.INIT('hecfd)
	) name1724 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w2257_
	);
	LUT4 #(
		.INIT('h0301)
	) name1725 (
		\sa32_reg[6]/NET0131 ,
		_w1445_,
		_w1451_,
		_w2257_,
		_w2258_
	);
	LUT3 #(
		.INIT('h07)
	) name1726 (
		_w1698_,
		_w1693_,
		_w2206_,
		_w2259_
	);
	LUT3 #(
		.INIT('hd0)
	) name1727 (
		\sa32_reg[2]/P0001 ,
		_w2258_,
		_w2259_,
		_w2260_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1728 (
		\sa32_reg[0]/P0002 ,
		_w2256_,
		_w2249_,
		_w2260_,
		_w2261_
	);
	LUT3 #(
		.INIT('h08)
	) name1729 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w2262_
	);
	LUT3 #(
		.INIT('h54)
	) name1730 (
		\sa32_reg[2]/P0001 ,
		_w1748_,
		_w2262_,
		_w2263_
	);
	LUT3 #(
		.INIT('h20)
	) name1731 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w2264_
	);
	LUT2 #(
		.INIT('h8)
	) name1732 (
		_w1724_,
		_w2264_,
		_w2265_
	);
	LUT3 #(
		.INIT('h07)
	) name1733 (
		_w1491_,
		_w1524_,
		_w1733_,
		_w2266_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1734 (
		\sa32_reg[1]/P0001 ,
		_w2263_,
		_w2265_,
		_w2266_,
		_w2267_
	);
	LUT2 #(
		.INIT('h1)
	) name1735 (
		_w1476_,
		_w2198_,
		_w2268_
	);
	LUT4 #(
		.INIT('h0002)
	) name1736 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2269_
	);
	LUT3 #(
		.INIT('h07)
	) name1737 (
		\sa32_reg[6]/NET0131 ,
		_w1521_,
		_w2269_,
		_w2270_
	);
	LUT3 #(
		.INIT('h15)
	) name1738 (
		\sa32_reg[2]/P0001 ,
		_w2268_,
		_w2270_,
		_w2271_
	);
	LUT4 #(
		.INIT('hf2fa)
	) name1739 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		_w2272_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1740 (
		\sa32_reg[7]/P0001 ,
		_w1546_,
		_w2155_,
		_w2272_,
		_w2273_
	);
	LUT4 #(
		.INIT('h0008)
	) name1741 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2274_
	);
	LUT4 #(
		.INIT('h7ff7)
	) name1742 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2275_
	);
	LUT3 #(
		.INIT('ha2)
	) name1743 (
		\sa32_reg[1]/P0001 ,
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w2276_
	);
	LUT4 #(
		.INIT('h0002)
	) name1744 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2277_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name1745 (
		_w1546_,
		_w2275_,
		_w2276_,
		_w2277_,
		_w2278_
	);
	LUT3 #(
		.INIT('he0)
	) name1746 (
		\sa32_reg[1]/P0001 ,
		_w2273_,
		_w2278_,
		_w2279_
	);
	LUT4 #(
		.INIT('h5455)
	) name1747 (
		\sa32_reg[0]/P0002 ,
		_w2271_,
		_w2267_,
		_w2279_,
		_w2280_
	);
	LUT4 #(
		.INIT('h0004)
	) name1748 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2281_
	);
	LUT4 #(
		.INIT('hadfb)
	) name1749 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2282_
	);
	LUT4 #(
		.INIT('h1000)
	) name1750 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2283_
	);
	LUT4 #(
		.INIT('h0072)
	) name1751 (
		\sa32_reg[3]/P0001 ,
		_w1450_,
		_w2282_,
		_w2283_,
		_w2284_
	);
	LUT2 #(
		.INIT('h2)
	) name1752 (
		_w1754_,
		_w2284_,
		_w2285_
	);
	LUT2 #(
		.INIT('h2)
	) name1753 (
		\sa32_reg[2]/P0001 ,
		_w1510_,
		_w2286_
	);
	LUT4 #(
		.INIT('hbdff)
	) name1754 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w2287_
	);
	LUT3 #(
		.INIT('h10)
	) name1755 (
		_w1476_,
		_w2198_,
		_w2287_,
		_w2288_
	);
	LUT4 #(
		.INIT('h4000)
	) name1756 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w2289_
	);
	LUT4 #(
		.INIT('h0007)
	) name1757 (
		\sa32_reg[3]/P0001 ,
		_w1527_,
		_w1462_,
		_w2289_,
		_w2290_
	);
	LUT4 #(
		.INIT('hf250)
	) name1758 (
		\sa32_reg[2]/P0001 ,
		_w1510_,
		_w2288_,
		_w2290_,
		_w2291_
	);
	LUT4 #(
		.INIT('h23af)
	) name1759 (
		\sa32_reg[5]/P0001 ,
		_w1450_,
		_w1512_,
		_w1463_,
		_w2292_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name1760 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2293_
	);
	LUT3 #(
		.INIT('h20)
	) name1761 (
		\sa32_reg[1]/P0001 ,
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		_w2294_
	);
	LUT2 #(
		.INIT('h4)
	) name1762 (
		_w2293_,
		_w2294_,
		_w2295_
	);
	LUT3 #(
		.INIT('h0e)
	) name1763 (
		\sa32_reg[2]/P0001 ,
		_w2292_,
		_w2295_,
		_w2296_
	);
	LUT4 #(
		.INIT('h0e00)
	) name1764 (
		\sa32_reg[1]/P0001 ,
		_w2291_,
		_w2285_,
		_w2296_,
		_w2297_
	);
	LUT3 #(
		.INIT('h10)
	) name1765 (
		_w2280_,
		_w2261_,
		_w2297_,
		_w2298_
	);
	LUT4 #(
		.INIT('h5540)
	) name1766 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w1692_,
		_w1734_,
		_w2299_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name1767 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2300_
	);
	LUT2 #(
		.INIT('h2)
	) name1768 (
		\sa32_reg[2]/P0001 ,
		_w2300_,
		_w2301_
	);
	LUT4 #(
		.INIT('h153f)
	) name1769 (
		_w1483_,
		_w1467_,
		_w1475_,
		_w1693_,
		_w2302_
	);
	LUT4 #(
		.INIT('h5455)
	) name1770 (
		\sa32_reg[1]/P0001 ,
		_w2301_,
		_w2299_,
		_w2302_,
		_w2303_
	);
	LUT4 #(
		.INIT('h0800)
	) name1771 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w2304_
	);
	LUT3 #(
		.INIT('h01)
	) name1772 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w2305_
	);
	LUT4 #(
		.INIT('h5554)
	) name1773 (
		\sa32_reg[2]/P0001 ,
		_w1720_,
		_w2305_,
		_w2304_,
		_w2306_
	);
	LUT3 #(
		.INIT('ha8)
	) name1774 (
		\sa32_reg[2]/P0001 ,
		_w1476_,
		_w1725_,
		_w2307_
	);
	LUT3 #(
		.INIT('h01)
	) name1775 (
		_w1503_,
		_w1505_,
		_w1462_,
		_w2308_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1776 (
		\sa32_reg[1]/P0001 ,
		_w2307_,
		_w2306_,
		_w2308_,
		_w2309_
	);
	LUT4 #(
		.INIT('h575f)
	) name1777 (
		\sa32_reg[7]/P0001 ,
		_w1449_,
		_w1445_,
		_w1467_,
		_w2310_
	);
	LUT2 #(
		.INIT('h1)
	) name1778 (
		_w1473_,
		_w1746_,
		_w2311_
	);
	LUT4 #(
		.INIT('h1333)
	) name1779 (
		\sa32_reg[4]/P0001 ,
		_w1535_,
		_w1546_,
		_w1547_,
		_w2312_
	);
	LUT4 #(
		.INIT('hd800)
	) name1780 (
		\sa32_reg[2]/P0001 ,
		_w2311_,
		_w2310_,
		_w2312_,
		_w2313_
	);
	LUT4 #(
		.INIT('h5455)
	) name1781 (
		\sa32_reg[0]/P0002 ,
		_w2309_,
		_w2303_,
		_w2313_,
		_w2314_
	);
	LUT2 #(
		.INIT('h4)
	) name1782 (
		\sa32_reg[1]/P0001 ,
		_w1458_,
		_w2315_
	);
	LUT3 #(
		.INIT('h0d)
	) name1783 (
		_w1453_,
		_w1489_,
		_w2274_,
		_w2316_
	);
	LUT3 #(
		.INIT('h45)
	) name1784 (
		\sa32_reg[3]/P0001 ,
		_w2315_,
		_w2316_,
		_w2317_
	);
	LUT4 #(
		.INIT('h0001)
	) name1785 (
		_w1733_,
		_w2209_,
		_w2237_,
		_w2274_,
		_w2318_
	);
	LUT4 #(
		.INIT('h0031)
	) name1786 (
		_w1442_,
		_w1521_,
		_w1737_,
		_w2237_,
		_w2319_
	);
	LUT4 #(
		.INIT('hfca8)
	) name1787 (
		\sa32_reg[1]/P0001 ,
		\sa32_reg[2]/P0001 ,
		_w2318_,
		_w2319_,
		_w2320_
	);
	LUT3 #(
		.INIT('h8a)
	) name1788 (
		\sa32_reg[0]/P0002 ,
		_w2317_,
		_w2320_,
		_w2321_
	);
	LUT3 #(
		.INIT('h07)
	) name1789 (
		_w1449_,
		_w1689_,
		_w2283_,
		_w2322_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1790 (
		\sa32_reg[2]/P0001 ,
		_w2152_,
		_w2227_,
		_w2264_,
		_w2323_
	);
	LUT3 #(
		.INIT('ha2)
	) name1791 (
		\sa32_reg[0]/P0002 ,
		_w2322_,
		_w2323_,
		_w2324_
	);
	LUT3 #(
		.INIT('h04)
	) name1792 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w2325_
	);
	LUT3 #(
		.INIT('h54)
	) name1793 (
		_w1491_,
		_w1493_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h1)
	) name1794 (
		_w1462_,
		_w1701_,
		_w2327_
	);
	LUT3 #(
		.INIT('h45)
	) name1795 (
		\sa32_reg[2]/P0001 ,
		_w2326_,
		_w2327_,
		_w2328_
	);
	LUT3 #(
		.INIT('ha8)
	) name1796 (
		\sa32_reg[1]/P0001 ,
		_w2324_,
		_w2328_,
		_w2329_
	);
	LUT4 #(
		.INIT('h0100)
	) name1797 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2330_
	);
	LUT4 #(
		.INIT('h0007)
	) name1798 (
		\sa32_reg[6]/NET0131 ,
		_w1510_,
		_w1535_,
		_w2330_,
		_w2331_
	);
	LUT4 #(
		.INIT('h0007)
	) name1799 (
		_w1443_,
		_w1472_,
		_w1696_,
		_w1748_,
		_w2332_
	);
	LUT4 #(
		.INIT('hedff)
	) name1800 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w1455_,
		_w2333_
	);
	LUT4 #(
		.INIT('he400)
	) name1801 (
		\sa32_reg[2]/P0001 ,
		_w2332_,
		_w2331_,
		_w2333_,
		_w2334_
	);
	LUT4 #(
		.INIT('h8000)
	) name1802 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w2335_
	);
	LUT4 #(
		.INIT('hcc08)
	) name1803 (
		_w1453_,
		_w1754_,
		_w2134_,
		_w2335_,
		_w2336_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name1804 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2337_
	);
	LUT2 #(
		.INIT('h2)
	) name1805 (
		_w1546_,
		_w2337_,
		_w2338_
	);
	LUT2 #(
		.INIT('h1)
	) name1806 (
		_w2336_,
		_w2338_,
		_w2339_
	);
	LUT3 #(
		.INIT('he0)
	) name1807 (
		\sa32_reg[1]/P0001 ,
		_w2334_,
		_w2339_,
		_w2340_
	);
	LUT4 #(
		.INIT('h0100)
	) name1808 (
		_w2314_,
		_w2329_,
		_w2321_,
		_w2340_,
		_w2341_
	);
	LUT4 #(
		.INIT('h6996)
	) name1809 (
		\u0_w_reg[3][9]/P0001 ,
		_w2244_,
		_w2298_,
		_w2341_,
		_w2342_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1810 (
		\sa21_reg[2]/P0001 ,
		_w1395_,
		_w1430_,
		_w1777_,
		_w2343_
	);
	LUT3 #(
		.INIT('h10)
	) name1811 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2344_
	);
	LUT4 #(
		.INIT('h0100)
	) name1812 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2345_
	);
	LUT2 #(
		.INIT('h8)
	) name1813 (
		_w1765_,
		_w2345_,
		_w2346_
	);
	LUT3 #(
		.INIT('h8a)
	) name1814 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2347_
	);
	LUT4 #(
		.INIT('h0010)
	) name1815 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w2348_
	);
	LUT3 #(
		.INIT('h0d)
	) name1816 (
		_w1419_,
		_w2347_,
		_w2348_,
		_w2349_
	);
	LUT4 #(
		.INIT('h5455)
	) name1817 (
		\sa21_reg[1]/P0001 ,
		_w2343_,
		_w2346_,
		_w2349_,
		_w2350_
	);
	LUT4 #(
		.INIT('h5155)
	) name1818 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w2351_
	);
	LUT4 #(
		.INIT('hff9d)
	) name1819 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w2352_
	);
	LUT3 #(
		.INIT('h40)
	) name1820 (
		_w1799_,
		_w2351_,
		_w2352_,
		_w2353_
	);
	LUT4 #(
		.INIT('h002a)
	) name1821 (
		\sa21_reg[2]/P0001 ,
		_w1334_,
		_w1360_,
		_w2089_,
		_w2354_
	);
	LUT3 #(
		.INIT('h13)
	) name1822 (
		_w1354_,
		_w2353_,
		_w2354_,
		_w2355_
	);
	LUT4 #(
		.INIT('h4041)
	) name1823 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2356_
	);
	LUT3 #(
		.INIT('ha8)
	) name1824 (
		\sa21_reg[1]/P0001 ,
		_w1407_,
		_w2356_,
		_w2357_
	);
	LUT3 #(
		.INIT('h23)
	) name1825 (
		\sa21_reg[5]/P0001 ,
		_w1400_,
		_w2015_,
		_w2358_
	);
	LUT2 #(
		.INIT('h4)
	) name1826 (
		_w2357_,
		_w2358_,
		_w2359_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1827 (
		\sa21_reg[0]/P0001 ,
		_w2350_,
		_w2355_,
		_w2359_,
		_w2360_
	);
	LUT4 #(
		.INIT('h8000)
	) name1828 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2361_
	);
	LUT4 #(
		.INIT('h0001)
	) name1829 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w2362_
	);
	LUT4 #(
		.INIT('h0007)
	) name1830 (
		_w1334_,
		_w1360_,
		_w2361_,
		_w2362_,
		_w2363_
	);
	LUT3 #(
		.INIT('hb9)
	) name1831 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2364_
	);
	LUT3 #(
		.INIT('h8f)
	) name1832 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2365_
	);
	LUT2 #(
		.INIT('h4)
	) name1833 (
		\sa21_reg[1]/P0001 ,
		\sa21_reg[2]/P0001 ,
		_w2366_
	);
	LUT3 #(
		.INIT('h40)
	) name1834 (
		\sa21_reg[1]/P0001 ,
		\sa21_reg[2]/P0001 ,
		\sa21_reg[5]/P0001 ,
		_w2367_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name1835 (
		_w1415_,
		_w2364_,
		_w2365_,
		_w2367_,
		_w2368_
	);
	LUT3 #(
		.INIT('he0)
	) name1836 (
		\sa21_reg[2]/P0001 ,
		_w2363_,
		_w2368_,
		_w2369_
	);
	LUT4 #(
		.INIT('h0888)
	) name1837 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2370_
	);
	LUT4 #(
		.INIT('h8007)
	) name1838 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2371_
	);
	LUT4 #(
		.INIT('h0100)
	) name1839 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w2372_
	);
	LUT4 #(
		.INIT('h0007)
	) name1840 (
		\sa21_reg[2]/P0001 ,
		_w1794_,
		_w2372_,
		_w2371_,
		_w2373_
	);
	LUT4 #(
		.INIT('hb8fc)
	) name1841 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		_w1789_,
		_w1797_,
		_w2374_
	);
	LUT3 #(
		.INIT('hd8)
	) name1842 (
		\sa21_reg[1]/P0001 ,
		_w2373_,
		_w2374_,
		_w2375_
	);
	LUT3 #(
		.INIT('h15)
	) name1843 (
		\sa21_reg[0]/P0001 ,
		_w2369_,
		_w2375_,
		_w2376_
	);
	LUT3 #(
		.INIT('h01)
	) name1844 (
		\sa21_reg[2]/P0001 ,
		_w1768_,
		_w2018_,
		_w2377_
	);
	LUT4 #(
		.INIT('h002a)
	) name1845 (
		\sa21_reg[2]/P0001 ,
		_w1344_,
		_w1394_,
		_w1411_,
		_w2378_
	);
	LUT4 #(
		.INIT('h0040)
	) name1846 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w2379_
	);
	LUT4 #(
		.INIT('h135f)
	) name1847 (
		_w1350_,
		_w1355_,
		_w1387_,
		_w2379_,
		_w2380_
	);
	LUT4 #(
		.INIT('hf400)
	) name1848 (
		_w2109_,
		_w2377_,
		_w2378_,
		_w2380_,
		_w2381_
	);
	LUT4 #(
		.INIT('ha888)
	) name1849 (
		\sa21_reg[6]/NET0131 ,
		_w1389_,
		_w1375_,
		_w1426_,
		_w2382_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1850 (
		\sa21_reg[2]/P0001 ,
		_w1336_,
		_w1370_,
		_w2040_,
		_w2383_
	);
	LUT2 #(
		.INIT('h8)
	) name1851 (
		_w1356_,
		_w1376_,
		_w2384_
	);
	LUT4 #(
		.INIT('h0777)
	) name1852 (
		_w1327_,
		_w1394_,
		_w1401_,
		_w1420_,
		_w2385_
	);
	LUT3 #(
		.INIT('h10)
	) name1853 (
		_w2383_,
		_w2384_,
		_w2385_,
		_w2386_
	);
	LUT4 #(
		.INIT('h3210)
	) name1854 (
		\sa21_reg[1]/P0001 ,
		_w2382_,
		_w2381_,
		_w2386_,
		_w2387_
	);
	LUT3 #(
		.INIT('h10)
	) name1855 (
		_w2376_,
		_w2360_,
		_w2387_,
		_w2388_
	);
	LUT3 #(
		.INIT('h13)
	) name1856 (
		_w1248_,
		_w1217_,
		_w1238_,
		_w2389_
	);
	LUT3 #(
		.INIT('h4c)
	) name1857 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w2390_
	);
	LUT3 #(
		.INIT('h4c)
	) name1858 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w2391_
	);
	LUT4 #(
		.INIT('hb300)
	) name1859 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2392_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1860 (
		\sa10_reg[2]/P0001 ,
		_w1267_,
		_w2390_,
		_w2392_,
		_w2393_
	);
	LUT3 #(
		.INIT('ha2)
	) name1861 (
		\sa10_reg[1]/P0001 ,
		_w2389_,
		_w2393_,
		_w2394_
	);
	LUT4 #(
		.INIT('h0040)
	) name1862 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2395_
	);
	LUT4 #(
		.INIT('h0001)
	) name1863 (
		_w1306_,
		_w1577_,
		_w1571_,
		_w2395_,
		_w2396_
	);
	LUT2 #(
		.INIT('h1)
	) name1864 (
		\sa10_reg[2]/P0001 ,
		_w2396_,
		_w2397_
	);
	LUT4 #(
		.INIT('h0888)
	) name1865 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2398_
	);
	LUT2 #(
		.INIT('h4)
	) name1866 (
		_w1241_,
		_w2398_,
		_w2399_
	);
	LUT4 #(
		.INIT('h0203)
	) name1867 (
		\sa10_reg[6]/NET0131 ,
		_w1577_,
		_w1953_,
		_w1996_,
		_w2400_
	);
	LUT4 #(
		.INIT('h113f)
	) name1868 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1236_,
		_w1839_,
		_w2401_
	);
	LUT4 #(
		.INIT('hba00)
	) name1869 (
		\sa10_reg[1]/P0001 ,
		_w2399_,
		_w2400_,
		_w2401_,
		_w2402_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1870 (
		\sa10_reg[0]/P0001 ,
		_w2394_,
		_w2397_,
		_w2402_,
		_w2403_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name1871 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2404_
	);
	LUT2 #(
		.INIT('h2)
	) name1872 (
		\sa10_reg[2]/P0001 ,
		_w2404_,
		_w2405_
	);
	LUT4 #(
		.INIT('h5510)
	) name1873 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		_w1217_,
		_w1295_,
		_w2406_
	);
	LUT4 #(
		.INIT('h13df)
	) name1874 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		_w1218_,
		_w1837_,
		_w2407_
	);
	LUT4 #(
		.INIT('h5455)
	) name1875 (
		\sa10_reg[0]/P0001 ,
		_w2406_,
		_w2405_,
		_w2407_,
		_w2408_
	);
	LUT4 #(
		.INIT('h0023)
	) name1876 (
		\sa10_reg[7]/NET0131 ,
		_w1225_,
		_w1287_,
		_w1557_,
		_w2409_
	);
	LUT4 #(
		.INIT('hedff)
	) name1877 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w1227_,
		_w2410_
	);
	LUT3 #(
		.INIT('he0)
	) name1878 (
		\sa10_reg[2]/P0001 ,
		_w2409_,
		_w2410_,
		_w2411_
	);
	LUT3 #(
		.INIT('h45)
	) name1879 (
		\sa10_reg[1]/P0001 ,
		_w2408_,
		_w2411_,
		_w2412_
	);
	LUT3 #(
		.INIT('h10)
	) name1880 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2413_
	);
	LUT4 #(
		.INIT('h0803)
	) name1881 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w2414_
	);
	LUT3 #(
		.INIT('h54)
	) name1882 (
		\sa10_reg[2]/P0001 ,
		_w2413_,
		_w2414_,
		_w2415_
	);
	LUT3 #(
		.INIT('ha8)
	) name1883 (
		\sa10_reg[2]/P0001 ,
		_w1252_,
		_w1278_,
		_w2416_
	);
	LUT3 #(
		.INIT('h01)
	) name1884 (
		_w1281_,
		_w1615_,
		_w1872_,
		_w2417_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1885 (
		\sa10_reg[1]/P0001 ,
		_w2415_,
		_w2416_,
		_w2417_,
		_w2418_
	);
	LUT4 #(
		.INIT('h153f)
	) name1886 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1247_,
		_w1837_,
		_w2419_
	);
	LUT4 #(
		.INIT('hffa8)
	) name1887 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2420_
	);
	LUT2 #(
		.INIT('h2)
	) name1888 (
		_w1277_,
		_w2420_,
		_w2421_
	);
	LUT4 #(
		.INIT('h007f)
	) name1889 (
		\sa10_reg[5]/P0001 ,
		_w1269_,
		_w1308_,
		_w1318_,
		_w2422_
	);
	LUT4 #(
		.INIT('h3200)
	) name1890 (
		\sa10_reg[2]/P0001 ,
		_w2421_,
		_w2419_,
		_w2422_,
		_w2423_
	);
	LUT3 #(
		.INIT('h45)
	) name1891 (
		\sa10_reg[0]/P0001 ,
		_w2418_,
		_w2423_,
		_w2424_
	);
	LUT4 #(
		.INIT('h0010)
	) name1892 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w2425_
	);
	LUT3 #(
		.INIT('h01)
	) name1893 (
		_w1249_,
		_w1615_,
		_w2425_,
		_w2426_
	);
	LUT2 #(
		.INIT('h1)
	) name1894 (
		_w1258_,
		_w1236_,
		_w2427_
	);
	LUT4 #(
		.INIT('h3111)
	) name1895 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[2]/P0001 ,
		_w2426_,
		_w2427_,
		_w2428_
	);
	LUT4 #(
		.INIT('h0100)
	) name1896 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2429_
	);
	LUT4 #(
		.INIT('h0015)
	) name1897 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1252_,
		_w1318_,
		_w2430_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name1898 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2431_
	);
	LUT2 #(
		.INIT('h2)
	) name1899 (
		\sa10_reg[3]/P0001 ,
		_w2431_,
		_w2432_
	);
	LUT3 #(
		.INIT('h70)
	) name1900 (
		_w1251_,
		_w1267_,
		_w1304_,
		_w2433_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1901 (
		_w2429_,
		_w2430_,
		_w2432_,
		_w2433_,
		_w2434_
	);
	LUT4 #(
		.INIT('h153f)
	) name1902 (
		_w1255_,
		_w1238_,
		_w1286_,
		_w1960_,
		_w2435_
	);
	LUT3 #(
		.INIT('h45)
	) name1903 (
		_w2428_,
		_w2434_,
		_w2435_,
		_w2436_
	);
	LUT4 #(
		.INIT('h0001)
	) name1904 (
		_w2412_,
		_w2403_,
		_w2424_,
		_w2436_,
		_w2437_
	);
	LUT4 #(
		.INIT('h5510)
	) name1905 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1099_,
		_w1196_,
		_w2438_
	);
	LUT4 #(
		.INIT('h0777)
	) name1906 (
		_w1064_,
		_w1123_,
		_w1060_,
		_w1933_,
		_w2439_
	);
	LUT3 #(
		.INIT('h45)
	) name1907 (
		\sa03_reg[1]/P0001 ,
		_w2438_,
		_w2439_,
		_w2440_
	);
	LUT3 #(
		.INIT('h10)
	) name1908 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2441_
	);
	LUT4 #(
		.INIT('hf7fc)
	) name1909 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w2442_
	);
	LUT3 #(
		.INIT('h45)
	) name1910 (
		\sa03_reg[2]/P0001 ,
		_w2441_,
		_w2442_,
		_w2443_
	);
	LUT3 #(
		.INIT('h01)
	) name1911 (
		_w1097_,
		_w1046_,
		_w1048_,
		_w2444_
	);
	LUT3 #(
		.INIT('h8a)
	) name1912 (
		\sa03_reg[1]/P0001 ,
		_w2443_,
		_w2444_,
		_w2445_
	);
	LUT4 #(
		.INIT('hffa8)
	) name1913 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2446_
	);
	LUT2 #(
		.INIT('h2)
	) name1914 (
		_w1069_,
		_w2446_,
		_w2447_
	);
	LUT2 #(
		.INIT('h8)
	) name1915 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[2]/P0001 ,
		_w2448_
	);
	LUT4 #(
		.INIT('h4000)
	) name1916 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2449_
	);
	LUT3 #(
		.INIT('hc8)
	) name1917 (
		_w1082_,
		_w2448_,
		_w2449_,
		_w2450_
	);
	LUT3 #(
		.INIT('h13)
	) name1918 (
		_w1115_,
		_w1135_,
		_w1143_,
		_w2451_
	);
	LUT3 #(
		.INIT('h10)
	) name1919 (
		_w2450_,
		_w2447_,
		_w2451_,
		_w2452_
	);
	LUT4 #(
		.INIT('h0777)
	) name1920 (
		_w1082_,
		_w1083_,
		_w1060_,
		_w1933_,
		_w2453_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name1921 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2454_
	);
	LUT2 #(
		.INIT('h2)
	) name1922 (
		_w1165_,
		_w2454_,
		_w2455_
	);
	LUT3 #(
		.INIT('h0e)
	) name1923 (
		\sa03_reg[2]/P0001 ,
		_w2453_,
		_w2455_,
		_w2456_
	);
	LUT4 #(
		.INIT('h1000)
	) name1924 (
		_w2445_,
		_w2440_,
		_w2452_,
		_w2456_,
		_w2457_
	);
	LUT3 #(
		.INIT('h07)
	) name1925 (
		_w1064_,
		_w1054_,
		_w1112_,
		_w2458_
	);
	LUT3 #(
		.INIT('h80)
	) name1926 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2459_
	);
	LUT4 #(
		.INIT('hcedf)
	) name1927 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2460_
	);
	LUT3 #(
		.INIT('h8a)
	) name1928 (
		\sa03_reg[2]/P0001 ,
		_w2459_,
		_w2460_,
		_w2461_
	);
	LUT3 #(
		.INIT('ha2)
	) name1929 (
		\sa03_reg[1]/P0001 ,
		_w2458_,
		_w2461_,
		_w2462_
	);
	LUT4 #(
		.INIT('h5554)
	) name1930 (
		\sa03_reg[2]/P0001 ,
		_w1143_,
		_w1195_,
		_w1676_,
		_w2463_
	);
	LUT4 #(
		.INIT('h0888)
	) name1931 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2464_
	);
	LUT4 #(
		.INIT('h0400)
	) name1932 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2465_
	);
	LUT4 #(
		.INIT('h5510)
	) name1933 (
		\sa03_reg[1]/P0001 ,
		_w1116_,
		_w2464_,
		_w2465_,
		_w2466_
	);
	LUT3 #(
		.INIT('h04)
	) name1934 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w2467_
	);
	LUT3 #(
		.INIT('he3)
	) name1935 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w2468_
	);
	LUT2 #(
		.INIT('h2)
	) name1936 (
		_w2467_,
		_w2468_,
		_w2469_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1937 (
		_w1099_,
		_w1171_,
		_w1668_,
		_w2448_,
		_w2470_
	);
	LUT4 #(
		.INIT('h0100)
	) name1938 (
		_w2466_,
		_w2469_,
		_w2463_,
		_w2470_,
		_w2471_
	);
	LUT2 #(
		.INIT('h4)
	) name1939 (
		_w2462_,
		_w2471_,
		_w2472_
	);
	LUT4 #(
		.INIT('h0007)
	) name1940 (
		_w1053_,
		_w1054_,
		_w1103_,
		_w1135_,
		_w2473_
	);
	LUT4 #(
		.INIT('hedff)
	) name1941 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w1064_,
		_w2474_
	);
	LUT4 #(
		.INIT('h0455)
	) name1942 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[2]/P0001 ,
		_w2473_,
		_w2474_,
		_w2475_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name1943 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2476_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1944 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w1099_,
		_w2476_,
		_w2477_
	);
	LUT2 #(
		.INIT('h2)
	) name1945 (
		_w2448_,
		_w2477_,
		_w2478_
	);
	LUT4 #(
		.INIT('h000b)
	) name1946 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w2479_
	);
	LUT4 #(
		.INIT('hffa4)
	) name1947 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w2480_
	);
	LUT4 #(
		.INIT('h0010)
	) name1948 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w2481_
	);
	LUT4 #(
		.INIT('h0032)
	) name1949 (
		\sa03_reg[7]/NET0131 ,
		_w1163_,
		_w2480_,
		_w2481_,
		_w2482_
	);
	LUT2 #(
		.INIT('h2)
	) name1950 (
		_w1210_,
		_w2482_,
		_w2483_
	);
	LUT2 #(
		.INIT('h1)
	) name1951 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[2]/P0001 ,
		_w2484_
	);
	LUT4 #(
		.INIT('h0007)
	) name1952 (
		_w1053_,
		_w1079_,
		_w1153_,
		_w1621_,
		_w2485_
	);
	LUT2 #(
		.INIT('h8)
	) name1953 (
		_w1125_,
		_w1627_,
		_w2486_
	);
	LUT4 #(
		.INIT('h0051)
	) name1954 (
		_w1636_,
		_w2484_,
		_w2485_,
		_w2486_,
		_w2487_
	);
	LUT4 #(
		.INIT('h0100)
	) name1955 (
		_w2475_,
		_w2483_,
		_w2478_,
		_w2487_,
		_w2488_
	);
	LUT4 #(
		.INIT('he400)
	) name1956 (
		\sa03_reg[0]/P0001 ,
		_w2457_,
		_w2472_,
		_w2488_,
		_w2489_
	);
	LUT2 #(
		.INIT('h6)
	) name1957 (
		_w2437_,
		_w2489_,
		_w2490_
	);
	LUT4 #(
		.INIT('h9669)
	) name1958 (
		_w1830_,
		_w2388_,
		_w2437_,
		_w2489_,
		_w2491_
	);
	LUT3 #(
		.INIT('h28)
	) name1959 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[9]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w2492_
	);
	LUT4 #(
		.INIT('hff14)
	) name1960 (
		\ld_r_reg/P0001 ,
		_w2342_,
		_w2491_,
		_w2492_,
		_w2493_
	);
	LUT3 #(
		.INIT('h96)
	) name1961 (
		_w1149_,
		_w1948_,
		_w2002_,
		_w2494_
	);
	LUT3 #(
		.INIT('h69)
	) name1962 (
		\u0_w_reg[3][5]/P0001 ,
		_w2059_,
		_w2185_,
		_w2495_
	);
	LUT3 #(
		.INIT('h28)
	) name1963 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[5]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		_w2496_
	);
	LUT4 #(
		.INIT('hff14)
	) name1964 (
		\ld_r_reg/P0001 ,
		_w2494_,
		_w2495_,
		_w2496_,
		_w2497_
	);
	LUT4 #(
		.INIT('h6996)
	) name1965 (
		\u0_w_reg[3][28]/P0001 ,
		_w1895_,
		_w2121_,
		_w2185_,
		_w2498_
	);
	LUT3 #(
		.INIT('h53)
	) name1966 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w2499_
	);
	LUT4 #(
		.INIT('h0053)
	) name1967 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2500_
	);
	LUT2 #(
		.INIT('h1)
	) name1968 (
		\sa03_reg[2]/P0001 ,
		_w2500_,
		_w2501_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1969 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2502_
	);
	LUT3 #(
		.INIT('h20)
	) name1970 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w2503_
	);
	LUT3 #(
		.INIT('h10)
	) name1971 (
		_w2467_,
		_w2503_,
		_w2502_,
		_w2504_
	);
	LUT3 #(
		.INIT('h01)
	) name1972 (
		_w1121_,
		_w1185_,
		_w1681_,
		_w2505_
	);
	LUT4 #(
		.INIT('h02aa)
	) name1973 (
		\sa03_reg[1]/P0001 ,
		_w2501_,
		_w2504_,
		_w2505_,
		_w2506_
	);
	LUT4 #(
		.INIT('h0020)
	) name1974 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w2507_
	);
	LUT4 #(
		.INIT('h0007)
	) name1975 (
		_w1093_,
		_w1072_,
		_w1900_,
		_w2507_,
		_w2508_
	);
	LUT4 #(
		.INIT('hefdf)
	) name1976 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2509_
	);
	LUT2 #(
		.INIT('h1)
	) name1977 (
		\sa03_reg[2]/P0001 ,
		_w2509_,
		_w2510_
	);
	LUT4 #(
		.INIT('h0007)
	) name1978 (
		_w1115_,
		_w1067_,
		_w1135_,
		_w1198_,
		_w2511_
	);
	LUT4 #(
		.INIT('h4555)
	) name1979 (
		\sa03_reg[1]/P0001 ,
		_w2510_,
		_w2511_,
		_w2508_,
		_w2512_
	);
	LUT3 #(
		.INIT('h10)
	) name1980 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w2513_
	);
	LUT4 #(
		.INIT('h0100)
	) name1981 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w2514_
	);
	LUT4 #(
		.INIT('h8000)
	) name1982 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2515_
	);
	LUT4 #(
		.INIT('h0007)
	) name1983 (
		_w1082_,
		_w1083_,
		_w2514_,
		_w2515_,
		_w2516_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name1984 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2517_
	);
	LUT2 #(
		.INIT('h8)
	) name1985 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w2518_
	);
	LUT4 #(
		.INIT('h7077)
	) name1986 (
		_w1044_,
		_w1060_,
		_w2517_,
		_w2518_,
		_w2519_
	);
	LUT3 #(
		.INIT('he0)
	) name1987 (
		\sa03_reg[2]/P0001 ,
		_w2516_,
		_w2519_,
		_w2520_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1988 (
		\sa03_reg[0]/P0001 ,
		_w2512_,
		_w2506_,
		_w2520_,
		_w2521_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name1989 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1117_,
		_w1138_,
		_w2522_
	);
	LUT4 #(
		.INIT('h002a)
	) name1990 (
		\sa03_reg[1]/P0001 ,
		_w1105_,
		_w1054_,
		_w1924_,
		_w2523_
	);
	LUT4 #(
		.INIT('h23af)
	) name1991 (
		\sa03_reg[2]/P0001 ,
		_w1064_,
		_w1096_,
		_w1054_,
		_w2524_
	);
	LUT3 #(
		.INIT('h40)
	) name1992 (
		_w2522_,
		_w2523_,
		_w2524_,
		_w2525_
	);
	LUT2 #(
		.INIT('h1)
	) name1993 (
		\sa03_reg[1]/P0001 ,
		_w2514_,
		_w2526_
	);
	LUT3 #(
		.INIT('ha8)
	) name1994 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w2527_
	);
	LUT4 #(
		.INIT('h51f3)
	) name1995 (
		_w1098_,
		_w1074_,
		_w1126_,
		_w2527_,
		_w2528_
	);
	LUT3 #(
		.INIT('h40)
	) name1996 (
		_w1206_,
		_w2526_,
		_w2528_,
		_w2529_
	);
	LUT4 #(
		.INIT('h0015)
	) name1997 (
		\sa03_reg[2]/P0001 ,
		_w1053_,
		_w1054_,
		_w1130_,
		_w2530_
	);
	LUT4 #(
		.INIT('h0002)
	) name1998 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w2531_
	);
	LUT3 #(
		.INIT('h02)
	) name1999 (
		\sa03_reg[2]/P0001 ,
		_w1191_,
		_w2531_,
		_w2532_
	);
	LUT3 #(
		.INIT('h54)
	) name2000 (
		_w1057_,
		_w2530_,
		_w2532_,
		_w2533_
	);
	LUT4 #(
		.INIT('h0155)
	) name2001 (
		\sa03_reg[0]/P0001 ,
		_w2525_,
		_w2529_,
		_w2533_,
		_w2534_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name2002 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2535_
	);
	LUT2 #(
		.INIT('h2)
	) name2003 (
		_w1630_,
		_w2535_,
		_w2536_
	);
	LUT3 #(
		.INIT('h40)
	) name2004 (
		\sa03_reg[2]/P0001 ,
		_w1110_,
		_w1140_,
		_w2537_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2005 (
		\sa03_reg[1]/P0001 ,
		_w1919_,
		_w2537_,
		_w2536_,
		_w2538_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name2006 (
		\sa03_reg[5]/P0001 ,
		_w1056_,
		_w1053_,
		_w1079_,
		_w2539_
	);
	LUT2 #(
		.INIT('h2)
	) name2007 (
		_w1165_,
		_w2539_,
		_w2540_
	);
	LUT4 #(
		.INIT('h2000)
	) name2008 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w2541_
	);
	LUT3 #(
		.INIT('hc8)
	) name2009 (
		_w1185_,
		_w2448_,
		_w2541_,
		_w2542_
	);
	LUT4 #(
		.INIT('h575f)
	) name2010 (
		_w1064_,
		_w1110_,
		_w1123_,
		_w1125_,
		_w2543_
	);
	LUT4 #(
		.INIT('h0777)
	) name2011 (
		_w1112_,
		_w1115_,
		_w1917_,
		_w2484_,
		_w2544_
	);
	LUT3 #(
		.INIT('h40)
	) name2012 (
		_w2542_,
		_w2543_,
		_w2544_,
		_w2545_
	);
	LUT3 #(
		.INIT('h10)
	) name2013 (
		_w2538_,
		_w2540_,
		_w2545_,
		_w2546_
	);
	LUT3 #(
		.INIT('h10)
	) name2014 (
		_w2521_,
		_w2534_,
		_w2546_,
		_w2547_
	);
	LUT3 #(
		.INIT('h01)
	) name2015 (
		\sa10_reg[2]/P0001 ,
		_w1557_,
		_w1839_,
		_w2548_
	);
	LUT4 #(
		.INIT('hff3b)
	) name2016 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2549_
	);
	LUT3 #(
		.INIT('h20)
	) name2017 (
		\sa10_reg[2]/P0001 ,
		_w1256_,
		_w2549_,
		_w2550_
	);
	LUT4 #(
		.INIT('h0007)
	) name2018 (
		_w1238_,
		_w1286_,
		_w1297_,
		_w1318_,
		_w2551_
	);
	LUT4 #(
		.INIT('h0155)
	) name2019 (
		\sa10_reg[1]/P0001 ,
		_w2548_,
		_w2550_,
		_w2551_,
		_w2552_
	);
	LUT4 #(
		.INIT('h0c04)
	) name2020 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2553_
	);
	LUT3 #(
		.INIT('ha8)
	) name2021 (
		\sa10_reg[2]/P0001 ,
		_w1883_,
		_w2553_,
		_w2554_
	);
	LUT2 #(
		.INIT('h8)
	) name2022 (
		_w1223_,
		_w2390_,
		_w2555_
	);
	LUT3 #(
		.INIT('h01)
	) name2023 (
		_w1275_,
		_w1591_,
		_w1873_,
		_w2556_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2024 (
		\sa10_reg[1]/P0001 ,
		_w2555_,
		_w2554_,
		_w2556_,
		_w2557_
	);
	LUT4 #(
		.INIT('h0100)
	) name2025 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w2558_
	);
	LUT4 #(
		.INIT('h8000)
	) name2026 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2559_
	);
	LUT4 #(
		.INIT('h0007)
	) name2027 (
		\sa10_reg[7]/NET0131 ,
		_w1247_,
		_w2558_,
		_w2559_,
		_w2560_
	);
	LUT2 #(
		.INIT('h8)
	) name2028 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w2561_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name2029 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2562_
	);
	LUT4 #(
		.INIT('h7707)
	) name2030 (
		_w1224_,
		_w1885_,
		_w2561_,
		_w2562_,
		_w2563_
	);
	LUT3 #(
		.INIT('he0)
	) name2031 (
		\sa10_reg[2]/P0001 ,
		_w2560_,
		_w2563_,
		_w2564_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2032 (
		\sa10_reg[0]/P0001 ,
		_w2557_,
		_w2552_,
		_w2564_,
		_w2565_
	);
	LUT4 #(
		.INIT('h5400)
	) name2033 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2566_
	);
	LUT3 #(
		.INIT('ha8)
	) name2034 (
		\sa10_reg[2]/P0001 ,
		_w1308_,
		_w2566_,
		_w2567_
	);
	LUT4 #(
		.INIT('h0007)
	) name2035 (
		_w1244_,
		_w1262_,
		_w1309_,
		_w2558_,
		_w2568_
	);
	LUT3 #(
		.INIT('h45)
	) name2036 (
		\sa10_reg[1]/P0001 ,
		_w2567_,
		_w2568_,
		_w2569_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name2037 (
		\sa10_reg[2]/P0001 ,
		_w1248_,
		_w1257_,
		_w1284_,
		_w2570_
	);
	LUT3 #(
		.INIT('h0b)
	) name2038 (
		\sa10_reg[4]/P0001 ,
		_w1252_,
		_w1256_,
		_w2571_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name2039 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1238_,
		_w1569_,
		_w2572_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name2040 (
		\sa10_reg[1]/P0001 ,
		_w2570_,
		_w2571_,
		_w2572_,
		_w2573_
	);
	LUT4 #(
		.INIT('h5540)
	) name2041 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1252_,
		_w1253_,
		_w2574_
	);
	LUT2 #(
		.INIT('h8)
	) name2042 (
		_w1257_,
		_w1269_,
		_w2575_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name2043 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[5]/P0001 ,
		_w1300_,
		_w1951_,
		_w2576_
	);
	LUT3 #(
		.INIT('h10)
	) name2044 (
		_w2575_,
		_w2574_,
		_w2576_,
		_w2577_
	);
	LUT4 #(
		.INIT('h5455)
	) name2045 (
		\sa10_reg[0]/P0001 ,
		_w2573_,
		_w2569_,
		_w2577_,
		_w2578_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name2046 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2579_
	);
	LUT2 #(
		.INIT('h2)
	) name2047 (
		_w1230_,
		_w2579_,
		_w2580_
	);
	LUT3 #(
		.INIT('h02)
	) name2048 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w2581_
	);
	LUT4 #(
		.INIT('h135f)
	) name2049 (
		_w1278_,
		_w1569_,
		_w1567_,
		_w2581_,
		_w2582_
	);
	LUT3 #(
		.INIT('h8a)
	) name2050 (
		\sa10_reg[1]/P0001 ,
		_w2580_,
		_w2582_,
		_w2583_
	);
	LUT4 #(
		.INIT('h2000)
	) name2051 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w2584_
	);
	LUT3 #(
		.INIT('ha8)
	) name2052 (
		\sa10_reg[1]/P0001 ,
		_w1873_,
		_w2584_,
		_w2585_
	);
	LUT3 #(
		.INIT('ha8)
	) name2053 (
		\sa10_reg[2]/P0001 ,
		_w1835_,
		_w2585_,
		_w2586_
	);
	LUT4 #(
		.INIT('h8acf)
	) name2054 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1287_,
		_w1951_,
		_w2587_
	);
	LUT2 #(
		.INIT('h8)
	) name2055 (
		_w1837_,
		_w1995_,
		_w2588_
	);
	LUT4 #(
		.INIT('h135f)
	) name2056 (
		_w1255_,
		_w1217_,
		_w1218_,
		_w1269_,
		_w2589_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2057 (
		_w1613_,
		_w2587_,
		_w2588_,
		_w2589_,
		_w2590_
	);
	LUT3 #(
		.INIT('h10)
	) name2058 (
		_w2586_,
		_w2583_,
		_w2590_,
		_w2591_
	);
	LUT3 #(
		.INIT('h10)
	) name2059 (
		_w2578_,
		_w2565_,
		_w2591_,
		_w2592_
	);
	LUT4 #(
		.INIT('h9669)
	) name2060 (
		_w1619_,
		_w1685_,
		_w2547_,
		_w2592_,
		_w2593_
	);
	LUT3 #(
		.INIT('h82)
	) name2061 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[28]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w2594_
	);
	LUT4 #(
		.INIT('h00be)
	) name2062 (
		\ld_r_reg/P0001 ,
		_w2498_,
		_w2593_,
		_w2594_,
		_w2595_
	);
	LUT4 #(
		.INIT('h0c04)
	) name2063 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2596_
	);
	LUT3 #(
		.INIT('ha8)
	) name2064 (
		\sa21_reg[2]/P0001 ,
		_w1800_,
		_w2596_,
		_w2597_
	);
	LUT4 #(
		.INIT('h0001)
	) name2065 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2598_
	);
	LUT3 #(
		.INIT('h01)
	) name2066 (
		_w1817_,
		_w2085_,
		_w2598_,
		_w2599_
	);
	LUT3 #(
		.INIT('h02)
	) name2067 (
		\sa21_reg[1]/P0001 ,
		_w1335_,
		_w1761_,
		_w2600_
	);
	LUT3 #(
		.INIT('h40)
	) name2068 (
		_w2597_,
		_w2599_,
		_w2600_,
		_w2601_
	);
	LUT4 #(
		.INIT('h0001)
	) name2069 (
		\sa21_reg[1]/P0001 ,
		_w1422_,
		_w1411_,
		_w2091_,
		_w2602_
	);
	LUT4 #(
		.INIT('hefdf)
	) name2070 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2603_
	);
	LUT2 #(
		.INIT('h1)
	) name2071 (
		\sa21_reg[2]/P0001 ,
		_w2603_,
		_w2604_
	);
	LUT3 #(
		.INIT('h0e)
	) name2072 (
		_w1370_,
		_w1426_,
		_w1805_,
		_w2605_
	);
	LUT3 #(
		.INIT('h10)
	) name2073 (
		_w2604_,
		_w2605_,
		_w2602_,
		_w2606_
	);
	LUT4 #(
		.INIT('h0100)
	) name2074 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w2607_
	);
	LUT4 #(
		.INIT('h0007)
	) name2075 (
		_w1334_,
		_w1360_,
		_w2361_,
		_w2607_,
		_w2608_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name2076 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2609_
	);
	LUT4 #(
		.INIT('h7707)
	) name2077 (
		_w1378_,
		_w2020_,
		_w2048_,
		_w2609_,
		_w2610_
	);
	LUT3 #(
		.INIT('he0)
	) name2078 (
		\sa21_reg[2]/P0001 ,
		_w2608_,
		_w2610_,
		_w2611_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2079 (
		\sa21_reg[0]/P0001 ,
		_w2601_,
		_w2606_,
		_w2611_,
		_w2612_
	);
	LUT4 #(
		.INIT('ha820)
	) name2080 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w1338_,
		_w1400_,
		_w2613_
	);
	LUT4 #(
		.INIT('h0222)
	) name2081 (
		\sa21_reg[1]/P0001 ,
		_w1370_,
		_w1385_,
		_w1378_,
		_w2614_
	);
	LUT4 #(
		.INIT('h153f)
	) name2082 (
		_w1334_,
		_w1365_,
		_w1330_,
		_w1805_,
		_w2615_
	);
	LUT3 #(
		.INIT('h40)
	) name2083 (
		_w2613_,
		_w2614_,
		_w2615_,
		_w2616_
	);
	LUT3 #(
		.INIT('h01)
	) name2084 (
		\sa21_reg[1]/P0001 ,
		_w1421_,
		_w2607_,
		_w2617_
	);
	LUT4 #(
		.INIT('h5400)
	) name2085 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2618_
	);
	LUT3 #(
		.INIT('ha8)
	) name2086 (
		\sa21_reg[2]/P0001 ,
		_w1797_,
		_w2618_,
		_w2619_
	);
	LUT3 #(
		.INIT('h10)
	) name2087 (
		_w1433_,
		_w2619_,
		_w2617_,
		_w2620_
	);
	LUT4 #(
		.INIT('h5450)
	) name2088 (
		\sa21_reg[2]/P0001 ,
		_w1360_,
		_w1364_,
		_w1365_,
		_w2621_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name2089 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w2622_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2090 (
		\sa21_reg[2]/P0001 ,
		_w1338_,
		_w1413_,
		_w2622_,
		_w2623_
	);
	LUT2 #(
		.INIT('h4)
	) name2091 (
		_w2621_,
		_w2623_,
		_w2624_
	);
	LUT4 #(
		.INIT('h0155)
	) name2092 (
		\sa21_reg[0]/P0001 ,
		_w2616_,
		_w2620_,
		_w2624_,
		_w2625_
	);
	LUT4 #(
		.INIT('h2000)
	) name2093 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w2626_
	);
	LUT3 #(
		.INIT('ha8)
	) name2094 (
		\sa21_reg[2]/P0001 ,
		_w1335_,
		_w2626_,
		_w2627_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name2095 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2628_
	);
	LUT2 #(
		.INIT('h2)
	) name2096 (
		_w1356_,
		_w2628_,
		_w2629_
	);
	LUT2 #(
		.INIT('h8)
	) name2097 (
		_w1425_,
		_w2089_,
		_w2630_
	);
	LUT3 #(
		.INIT('h2a)
	) name2098 (
		\sa21_reg[1]/P0001 ,
		\sa21_reg[2]/P0001 ,
		_w2085_,
		_w2631_
	);
	LUT4 #(
		.INIT('h0100)
	) name2099 (
		_w2629_,
		_w2627_,
		_w2630_,
		_w2631_,
		_w2632_
	);
	LUT4 #(
		.INIT('hffed)
	) name2100 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2633_
	);
	LUT2 #(
		.INIT('h2)
	) name2101 (
		_w1375_,
		_w2633_,
		_w2634_
	);
	LUT3 #(
		.INIT('h80)
	) name2102 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2635_
	);
	LUT3 #(
		.INIT('h15)
	) name2103 (
		\sa21_reg[1]/P0001 ,
		_w1805_,
		_w2635_,
		_w2636_
	);
	LUT2 #(
		.INIT('h4)
	) name2104 (
		_w2634_,
		_w2636_,
		_w2637_
	);
	LUT4 #(
		.INIT('hedff)
	) name2105 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2638_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name2106 (
		\sa21_reg[7]/P0001 ,
		_w1431_,
		_w1414_,
		_w2638_,
		_w2639_
	);
	LUT3 #(
		.INIT('he0)
	) name2107 (
		_w2632_,
		_w2637_,
		_w2639_,
		_w2640_
	);
	LUT3 #(
		.INIT('h10)
	) name2108 (
		_w2625_,
		_w2612_,
		_w2640_,
		_w2641_
	);
	LUT4 #(
		.INIT('h6996)
	) name2109 (
		_w1619_,
		_w1948_,
		_w2592_,
		_w2641_,
		_w2642_
	);
	LUT4 #(
		.INIT('h9669)
	) name2110 (
		\u0_w_reg[3][20]/P0001 ,
		_w1830_,
		_w2121_,
		_w2185_,
		_w2643_
	);
	LUT3 #(
		.INIT('h82)
	) name2111 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[20]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w2644_
	);
	LUT4 #(
		.INIT('h00be)
	) name2112 (
		\ld_r_reg/P0001 ,
		_w2642_,
		_w2643_,
		_w2644_,
		_w2645_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2113 (
		\sa03_reg[2]/P0001 ,
		_w1090_,
		_w1049_,
		_w1208_,
		_w2646_
	);
	LUT2 #(
		.INIT('h8)
	) name2114 (
		_w1672_,
		_w1630_,
		_w2647_
	);
	LUT4 #(
		.INIT('h0010)
	) name2115 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w2648_
	);
	LUT3 #(
		.INIT('h0d)
	) name2116 (
		_w1059_,
		_w1629_,
		_w2648_,
		_w2649_
	);
	LUT4 #(
		.INIT('h5455)
	) name2117 (
		\sa03_reg[1]/P0001 ,
		_w2647_,
		_w2646_,
		_w2649_,
		_w2650_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name2118 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2651_
	);
	LUT4 #(
		.INIT('h0301)
	) name2119 (
		\sa03_reg[3]/P0001 ,
		_w1638_,
		_w1664_,
		_w2651_,
		_w2652_
	);
	LUT2 #(
		.INIT('h1)
	) name2120 (
		\sa03_reg[2]/P0001 ,
		_w2652_,
		_w2653_
	);
	LUT3 #(
		.INIT('h07)
	) name2121 (
		_w1082_,
		_w1083_,
		_w1897_,
		_w2654_
	);
	LUT3 #(
		.INIT('h2a)
	) name2122 (
		\sa03_reg[2]/P0001 ,
		_w1154_,
		_w2654_,
		_w2655_
	);
	LUT2 #(
		.INIT('h9)
	) name2123 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w2656_
	);
	LUT4 #(
		.INIT('h4041)
	) name2124 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2657_
	);
	LUT3 #(
		.INIT('ha8)
	) name2125 (
		\sa03_reg[1]/P0001 ,
		_w1196_,
		_w2657_,
		_w2658_
	);
	LUT3 #(
		.INIT('h07)
	) name2126 (
		_w1110_,
		_w1140_,
		_w1676_,
		_w2659_
	);
	LUT2 #(
		.INIT('h4)
	) name2127 (
		_w2658_,
		_w2659_,
		_w2660_
	);
	LUT4 #(
		.INIT('h0100)
	) name2128 (
		_w2655_,
		_w2653_,
		_w2650_,
		_w2660_,
		_w2661_
	);
	LUT4 #(
		.INIT('h0007)
	) name2129 (
		_w1082_,
		_w1083_,
		_w1187_,
		_w2515_,
		_w2662_
	);
	LUT3 #(
		.INIT('ha8)
	) name2130 (
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2663_
	);
	LUT3 #(
		.INIT('h08)
	) name2131 (
		_w1059_,
		_w2527_,
		_w2663_,
		_w2664_
	);
	LUT4 #(
		.INIT('h4c00)
	) name2132 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2665_
	);
	LUT2 #(
		.INIT('h8)
	) name2133 (
		_w1165_,
		_w2665_,
		_w2666_
	);
	LUT4 #(
		.INIT('h000e)
	) name2134 (
		\sa03_reg[2]/P0001 ,
		_w2662_,
		_w2664_,
		_w2666_,
		_w2667_
	);
	LUT4 #(
		.INIT('h0eee)
	) name2135 (
		\sa03_reg[3]/P0001 ,
		_w1669_,
		_w1623_,
		_w1620_,
		_w2668_
	);
	LUT4 #(
		.INIT('h8007)
	) name2136 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2669_
	);
	LUT4 #(
		.INIT('h0013)
	) name2137 (
		\sa03_reg[3]/P0001 ,
		_w1658_,
		_w1900_,
		_w2669_,
		_w2670_
	);
	LUT3 #(
		.INIT('he4)
	) name2138 (
		\sa03_reg[1]/P0001 ,
		_w2668_,
		_w2670_,
		_w2671_
	);
	LUT2 #(
		.INIT('h8)
	) name2139 (
		_w2667_,
		_w2671_,
		_w2672_
	);
	LUT4 #(
		.INIT('hff4b)
	) name2140 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2673_
	);
	LUT2 #(
		.INIT('h2)
	) name2141 (
		_w1630_,
		_w2673_,
		_w2674_
	);
	LUT2 #(
		.INIT('h8)
	) name2142 (
		_w1046_,
		_w1171_,
		_w2675_
	);
	LUT3 #(
		.INIT('h02)
	) name2143 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		_w2676_
	);
	LUT3 #(
		.INIT('h40)
	) name2144 (
		_w1116_,
		_w2656_,
		_w2676_,
		_w2677_
	);
	LUT4 #(
		.INIT('h0001)
	) name2145 (
		_w1144_,
		_w2677_,
		_w2675_,
		_w2674_,
		_w2678_
	);
	LUT2 #(
		.INIT('h8)
	) name2146 (
		_w1069_,
		_w1196_,
		_w2679_
	);
	LUT4 #(
		.INIT('h337f)
	) name2147 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1067_,
		_w1145_,
		_w2680_
	);
	LUT4 #(
		.INIT('h8acf)
	) name2148 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1187_,
		_w1681_,
		_w2681_
	);
	LUT3 #(
		.INIT('h40)
	) name2149 (
		_w2679_,
		_w2680_,
		_w2681_,
		_w2682_
	);
	LUT4 #(
		.INIT('h135f)
	) name2150 (
		\sa03_reg[6]/NET0131 ,
		_w1045_,
		_w1178_,
		_w2676_,
		_w2683_
	);
	LUT4 #(
		.INIT('he400)
	) name2151 (
		\sa03_reg[1]/P0001 ,
		_w2678_,
		_w2682_,
		_w2683_,
		_w2684_
	);
	LUT4 #(
		.INIT('hd800)
	) name2152 (
		\sa03_reg[0]/P0001 ,
		_w2661_,
		_w2672_,
		_w2684_,
		_w2685_
	);
	LUT4 #(
		.INIT('h9669)
	) name2153 (
		_w1685_,
		_w2437_,
		_w2489_,
		_w2685_,
		_w2686_
	);
	LUT2 #(
		.INIT('h4)
	) name2154 (
		_w1338_,
		_w2370_,
		_w2687_
	);
	LUT4 #(
		.INIT('h0400)
	) name2155 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2688_
	);
	LUT4 #(
		.INIT('h0007)
	) name2156 (
		_w1326_,
		_w1385_,
		_w1788_,
		_w2688_,
		_w2689_
	);
	LUT3 #(
		.INIT('h45)
	) name2157 (
		\sa21_reg[1]/P0001 ,
		_w2687_,
		_w2689_,
		_w2690_
	);
	LUT3 #(
		.INIT('h13)
	) name2158 (
		_w1365_,
		_w1337_,
		_w1330_,
		_w2691_
	);
	LUT3 #(
		.INIT('h10)
	) name2159 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w2692_
	);
	LUT3 #(
		.INIT('h20)
	) name2160 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w2693_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2161 (
		\sa21_reg[2]/P0001 ,
		_w2635_,
		_w2693_,
		_w2692_,
		_w2694_
	);
	LUT3 #(
		.INIT('ha2)
	) name2162 (
		\sa21_reg[1]/P0001 ,
		_w2691_,
		_w2694_,
		_w2695_
	);
	LUT4 #(
		.INIT('h5554)
	) name2163 (
		\sa21_reg[2]/P0001 ,
		_w1400_,
		_w1406_,
		_w1788_,
		_w2696_
	);
	LUT4 #(
		.INIT('h45cf)
	) name2164 (
		_w1391_,
		_w1414_,
		_w1798_,
		_w2072_,
		_w2697_
	);
	LUT2 #(
		.INIT('h4)
	) name2165 (
		_w2696_,
		_w2697_,
		_w2698_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2166 (
		\sa21_reg[0]/P0001 ,
		_w2695_,
		_w2690_,
		_w2698_,
		_w2699_
	);
	LUT4 #(
		.INIT('h5540)
	) name2167 (
		\sa21_reg[2]/P0001 ,
		_w1344_,
		_w1345_,
		_w1407_,
		_w2700_
	);
	LUT3 #(
		.INIT('h45)
	) name2168 (
		\sa21_reg[1]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w1431_,
		_w2701_
	);
	LUT2 #(
		.INIT('h8)
	) name2169 (
		\sa21_reg[2]/P0001 ,
		_w1400_,
		_w2702_
	);
	LUT4 #(
		.INIT('h0f7f)
	) name2170 (
		\sa21_reg[2]/P0001 ,
		_w1369_,
		_w1390_,
		_w1420_,
		_w2703_
	);
	LUT4 #(
		.INIT('h1000)
	) name2171 (
		_w2700_,
		_w2702_,
		_w2701_,
		_w2703_,
		_w2704_
	);
	LUT4 #(
		.INIT('h5554)
	) name2172 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w2705_
	);
	LUT3 #(
		.INIT('h10)
	) name2173 (
		_w1431_,
		_w2344_,
		_w2705_,
		_w2706_
	);
	LUT4 #(
		.INIT('h4000)
	) name2174 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2707_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2175 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w2708_
	);
	LUT2 #(
		.INIT('h4)
	) name2176 (
		_w2707_,
		_w2708_,
		_w2709_
	);
	LUT4 #(
		.INIT('h0002)
	) name2177 (
		\sa21_reg[1]/P0001 ,
		_w1794_,
		_w1815_,
		_w2010_,
		_w2710_
	);
	LUT3 #(
		.INIT('he0)
	) name2178 (
		_w2706_,
		_w2709_,
		_w2710_,
		_w2711_
	);
	LUT3 #(
		.INIT('h02)
	) name2179 (
		\sa21_reg[2]/P0001 ,
		_w1430_,
		_w2108_,
		_w2712_
	);
	LUT4 #(
		.INIT('h0015)
	) name2180 (
		\sa21_reg[2]/P0001 ,
		_w1334_,
		_w1360_,
		_w1422_,
		_w2713_
	);
	LUT4 #(
		.INIT('h5150)
	) name2181 (
		_w2055_,
		_w2106_,
		_w2712_,
		_w2713_,
		_w2714_
	);
	LUT4 #(
		.INIT('h0155)
	) name2182 (
		\sa21_reg[0]/P0001 ,
		_w2704_,
		_w2711_,
		_w2714_,
		_w2715_
	);
	LUT4 #(
		.INIT('h0015)
	) name2183 (
		_w1353_,
		_w1327_,
		_w1398_,
		_w1822_,
		_w2716_
	);
	LUT4 #(
		.INIT('h0777)
	) name2184 (
		_w1348_,
		_w1350_,
		_w1330_,
		_w1781_,
		_w2717_
	);
	LUT4 #(
		.INIT('h0155)
	) name2185 (
		\sa21_reg[1]/P0001 ,
		\sa21_reg[2]/P0001 ,
		_w2716_,
		_w2717_,
		_w2718_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name2186 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2719_
	);
	LUT4 #(
		.INIT('hbf15)
	) name2187 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		_w1391_,
		_w2719_,
		_w2720_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name2188 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2721_
	);
	LUT2 #(
		.INIT('h2)
	) name2189 (
		_w1414_,
		_w2721_,
		_w2722_
	);
	LUT3 #(
		.INIT('h0d)
	) name2190 (
		_w1418_,
		_w2720_,
		_w2722_,
		_w2723_
	);
	LUT4 #(
		.INIT('h0010)
	) name2191 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w2724_
	);
	LUT4 #(
		.INIT('hfff9)
	) name2192 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2725_
	);
	LUT4 #(
		.INIT('hffbe)
	) name2193 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2726_
	);
	LUT2 #(
		.INIT('h2)
	) name2194 (
		\sa21_reg[1]/P0001 ,
		\sa21_reg[2]/P0001 ,
		_w2727_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2195 (
		_w2724_,
		_w2725_,
		_w2726_,
		_w2727_,
		_w2728_
	);
	LUT4 #(
		.INIT('h0007)
	) name2196 (
		_w1360_,
		_w1365_,
		_w1422_,
		_w2345_,
		_w2729_
	);
	LUT3 #(
		.INIT('h31)
	) name2197 (
		_w2366_,
		_w2728_,
		_w2729_,
		_w2730_
	);
	LUT3 #(
		.INIT('h40)
	) name2198 (
		_w2718_,
		_w2723_,
		_w2730_,
		_w2731_
	);
	LUT3 #(
		.INIT('h10)
	) name2199 (
		_w2715_,
		_w2699_,
		_w2731_,
		_w2732_
	);
	LUT4 #(
		.INIT('h5655)
	) name2200 (
		\u0_w_reg[3][1]/P0001 ,
		_w2715_,
		_w2699_,
		_w2731_,
		_w2733_
	);
	LUT3 #(
		.INIT('h69)
	) name2201 (
		_w2244_,
		_w2298_,
		_w2733_,
		_w2734_
	);
	LUT3 #(
		.INIT('h28)
	) name2202 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[1]/P0001 ,
		\u0_w_reg[3][1]/P0001 ,
		_w2735_
	);
	LUT4 #(
		.INIT('hff14)
	) name2203 (
		\ld_r_reg/P0001 ,
		_w2686_,
		_w2734_,
		_w2735_,
		_w2736_
	);
	LUT4 #(
		.INIT('haa80)
	) name2204 (
		\sa32_reg[2]/P0001 ,
		_w1450_,
		_w1443_,
		_w1726_,
		_w2737_
	);
	LUT2 #(
		.INIT('h4)
	) name2205 (
		\sa32_reg[2]/P0001 ,
		_w1458_,
		_w2738_
	);
	LUT4 #(
		.INIT('h020a)
	) name2206 (
		\sa32_reg[1]/P0001 ,
		_w1449_,
		_w1514_,
		_w1689_,
		_w2739_
	);
	LUT4 #(
		.INIT('h0100)
	) name2207 (
		_w1477_,
		_w2738_,
		_w2737_,
		_w2739_,
		_w2740_
	);
	LUT4 #(
		.INIT('h0008)
	) name2208 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2741_
	);
	LUT3 #(
		.INIT('h01)
	) name2209 (
		\sa32_reg[1]/P0001 ,
		_w2269_,
		_w2741_,
		_w2742_
	);
	LUT3 #(
		.INIT('he0)
	) name2210 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2743_
	);
	LUT3 #(
		.INIT('h13)
	) name2211 (
		_w1724_,
		_w2253_,
		_w2743_,
		_w2744_
	);
	LUT3 #(
		.INIT('h40)
	) name2212 (
		_w1745_,
		_w2742_,
		_w2744_,
		_w2745_
	);
	LUT4 #(
		.INIT('h5540)
	) name2213 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w1510_,
		_w1703_,
		_w2746_
	);
	LUT2 #(
		.INIT('h8)
	) name2214 (
		_w1546_,
		_w1726_,
		_w2747_
	);
	LUT4 #(
		.INIT('h153f)
	) name2215 (
		\sa32_reg[2]/P0001 ,
		_w1482_,
		_w1524_,
		_w1740_,
		_w2748_
	);
	LUT3 #(
		.INIT('h10)
	) name2216 (
		_w2746_,
		_w2747_,
		_w2748_,
		_w2749_
	);
	LUT4 #(
		.INIT('h0155)
	) name2217 (
		\sa32_reg[0]/P0002 ,
		_w2740_,
		_w2745_,
		_w2749_,
		_w2750_
	);
	LUT3 #(
		.INIT('ha2)
	) name2218 (
		\sa32_reg[2]/P0001 ,
		_w1515_,
		_w1507_,
		_w2751_
	);
	LUT4 #(
		.INIT('hefdf)
	) name2219 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2752_
	);
	LUT2 #(
		.INIT('h1)
	) name2220 (
		\sa32_reg[2]/P0001 ,
		_w2752_,
		_w2753_
	);
	LUT4 #(
		.INIT('h0013)
	) name2221 (
		_w1460_,
		_w1535_,
		_w1689_,
		_w1741_,
		_w2754_
	);
	LUT4 #(
		.INIT('h5455)
	) name2222 (
		\sa32_reg[1]/P0001 ,
		_w2753_,
		_w2751_,
		_w2754_,
		_w2755_
	);
	LUT4 #(
		.INIT('hd1ff)
	) name2223 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2756_
	);
	LUT3 #(
		.INIT('h8a)
	) name2224 (
		\sa32_reg[2]/P0001 ,
		_w2325_,
		_w2756_,
		_w2757_
	);
	LUT4 #(
		.INIT('hffac)
	) name2225 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2758_
	);
	LUT2 #(
		.INIT('h1)
	) name2226 (
		\sa32_reg[2]/P0001 ,
		_w2758_,
		_w2759_
	);
	LUT3 #(
		.INIT('h01)
	) name2227 (
		_w1510_,
		_w1492_,
		_w2181_,
		_w2760_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2228 (
		\sa32_reg[1]/P0001 ,
		_w2757_,
		_w2759_,
		_w2760_,
		_w2761_
	);
	LUT4 #(
		.INIT('h0007)
	) name2229 (
		\sa32_reg[7]/P0001 ,
		_w1445_,
		_w2228_,
		_w2253_,
		_w2762_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name2230 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2763_
	);
	LUT4 #(
		.INIT('h7707)
	) name2231 (
		_w1528_,
		_w1457_,
		_w1539_,
		_w2763_,
		_w2764_
	);
	LUT3 #(
		.INIT('he0)
	) name2232 (
		\sa32_reg[2]/P0001 ,
		_w2762_,
		_w2764_,
		_w2765_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2233 (
		\sa32_reg[0]/P0002 ,
		_w2755_,
		_w2761_,
		_w2765_,
		_w2766_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name2234 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2767_
	);
	LUT2 #(
		.INIT('h2)
	) name2235 (
		_w1698_,
		_w2767_,
		_w2768_
	);
	LUT2 #(
		.INIT('h8)
	) name2236 (
		_w1514_,
		_w1489_,
		_w2769_
	);
	LUT4 #(
		.INIT('h2000)
	) name2237 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w2770_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2238 (
		\sa32_reg[2]/P0001 ,
		_w1492_,
		_w2181_,
		_w2770_,
		_w2771_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2239 (
		\sa32_reg[1]/P0001 ,
		_w2769_,
		_w2771_,
		_w2768_,
		_w2772_
	);
	LUT3 #(
		.INIT('h2a)
	) name2240 (
		\sa32_reg[2]/P0001 ,
		_w1443_,
		_w1472_,
		_w2773_
	);
	LUT3 #(
		.INIT('h54)
	) name2241 (
		\sa32_reg[1]/P0001 ,
		\sa32_reg[2]/P0001 ,
		_w2168_,
		_w2774_
	);
	LUT4 #(
		.INIT('hedff)
	) name2242 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2775_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2243 (
		_w1483_,
		_w1546_,
		_w1693_,
		_w2775_,
		_w2776_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2244 (
		_w1525_,
		_w2773_,
		_w2774_,
		_w2776_,
		_w2777_
	);
	LUT2 #(
		.INIT('h4)
	) name2245 (
		_w2772_,
		_w2777_,
		_w2778_
	);
	LUT3 #(
		.INIT('h10)
	) name2246 (
		_w2766_,
		_w2750_,
		_w2778_,
		_w2779_
	);
	LUT4 #(
		.INIT('h6996)
	) name2247 (
		\u0_w_reg[3][12]/P0001 ,
		_w2185_,
		_w2298_,
		_w2779_,
		_w2780_
	);
	LUT4 #(
		.INIT('h9669)
	) name2248 (
		_w1830_,
		_w1895_,
		_w1948_,
		_w2641_,
		_w2781_
	);
	LUT3 #(
		.INIT('h82)
	) name2249 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[12]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		_w2782_
	);
	LUT4 #(
		.INIT('h00be)
	) name2250 (
		\ld_r_reg/P0001 ,
		_w2780_,
		_w2781_,
		_w2782_,
		_w2783_
	);
	LUT4 #(
		.INIT('h0001)
	) name2251 (
		_w1561_,
		_w1837_,
		_w1844_,
		_w1860_,
		_w2784_
	);
	LUT2 #(
		.INIT('h1)
	) name2252 (
		_w1236_,
		_w1886_,
		_w2785_
	);
	LUT4 #(
		.INIT('haaef)
	) name2253 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[4]/P0001 ,
		_w1305_,
		_w1889_,
		_w2786_
	);
	LUT4 #(
		.INIT('h1555)
	) name2254 (
		\sa10_reg[1]/P0001 ,
		_w2784_,
		_w2785_,
		_w2786_,
		_w2787_
	);
	LUT4 #(
		.INIT('h0040)
	) name2255 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w2788_
	);
	LUT2 #(
		.INIT('h8)
	) name2256 (
		_w1215_,
		_w2788_,
		_w2789_
	);
	LUT4 #(
		.INIT('h0002)
	) name2257 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2790_
	);
	LUT3 #(
		.INIT('h07)
	) name2258 (
		_w1586_,
		_w2390_,
		_w2790_,
		_w2791_
	);
	LUT3 #(
		.INIT('h8a)
	) name2259 (
		\sa10_reg[1]/P0001 ,
		_w2789_,
		_w2791_,
		_w2792_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name2260 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2793_
	);
	LUT2 #(
		.INIT('h2)
	) name2261 (
		_w1269_,
		_w2793_,
		_w2794_
	);
	LUT4 #(
		.INIT('h45ef)
	) name2262 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1271_,
		_w1844_,
		_w2795_
	);
	LUT3 #(
		.INIT('h10)
	) name2263 (
		_w1842_,
		_w2794_,
		_w2795_,
		_w2796_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2264 (
		\sa10_reg[0]/P0001 ,
		_w2787_,
		_w2792_,
		_w2796_,
		_w2797_
	);
	LUT4 #(
		.INIT('hffda)
	) name2265 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2798_
	);
	LUT2 #(
		.INIT('h2)
	) name2266 (
		\sa10_reg[2]/P0001 ,
		_w2798_,
		_w2799_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name2267 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2800_
	);
	LUT3 #(
		.INIT('h51)
	) name2268 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w2801_
	);
	LUT3 #(
		.INIT('h45)
	) name2269 (
		_w1306_,
		_w2800_,
		_w2801_,
		_w2802_
	);
	LUT3 #(
		.INIT('h45)
	) name2270 (
		\sa10_reg[0]/P0001 ,
		_w2799_,
		_w2802_,
		_w2803_
	);
	LUT4 #(
		.INIT('h0400)
	) name2271 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2804_
	);
	LUT4 #(
		.INIT('h0013)
	) name2272 (
		_w1248_,
		_w1217_,
		_w1238_,
		_w2804_,
		_w2805_
	);
	LUT3 #(
		.INIT('h32)
	) name2273 (
		\sa10_reg[2]/P0001 ,
		_w1839_,
		_w2805_,
		_w2806_
	);
	LUT3 #(
		.INIT('h8a)
	) name2274 (
		\sa10_reg[1]/P0001 ,
		_w2803_,
		_w2806_,
		_w2807_
	);
	LUT3 #(
		.INIT('h02)
	) name2275 (
		\sa10_reg[2]/P0001 ,
		_w1607_,
		_w2581_,
		_w2808_
	);
	LUT4 #(
		.INIT('h0007)
	) name2276 (
		\sa10_reg[4]/P0001 ,
		_w1281_,
		_w1298_,
		_w1582_,
		_w2809_
	);
	LUT4 #(
		.INIT('h45cf)
	) name2277 (
		_w1237_,
		_w1838_,
		_w2808_,
		_w2809_,
		_w2810_
	);
	LUT3 #(
		.INIT('hb8)
	) name2278 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w2811_
	);
	LUT2 #(
		.INIT('h8)
	) name2279 (
		_w1286_,
		_w2811_,
		_w2812_
	);
	LUT3 #(
		.INIT('h54)
	) name2280 (
		\sa10_reg[1]/P0001 ,
		_w2810_,
		_w2812_,
		_w2813_
	);
	LUT3 #(
		.INIT('h54)
	) name2281 (
		\sa10_reg[1]/P0001 ,
		_w1607_,
		_w2788_,
		_w2814_
	);
	LUT3 #(
		.INIT('h15)
	) name2282 (
		_w1244_,
		_w1873_,
		_w2561_,
		_w2815_
	);
	LUT4 #(
		.INIT('h5455)
	) name2283 (
		\sa10_reg[0]/P0001 ,
		_w1313_,
		_w2814_,
		_w2815_,
		_w2816_
	);
	LUT3 #(
		.INIT('had)
	) name2284 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2817_
	);
	LUT2 #(
		.INIT('h2)
	) name2285 (
		_w1270_,
		_w2817_,
		_w2818_
	);
	LUT3 #(
		.INIT('ha8)
	) name2286 (
		\sa10_reg[1]/P0001 ,
		_w1271_,
		_w1889_,
		_w2819_
	);
	LUT3 #(
		.INIT('h80)
	) name2287 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[2]/P0001 ,
		\sa10_reg[3]/P0001 ,
		_w2820_
	);
	LUT4 #(
		.INIT('h153f)
	) name2288 (
		_w1577_,
		_w1569_,
		_w2581_,
		_w2820_,
		_w2821_
	);
	LUT4 #(
		.INIT('h5700)
	) name2289 (
		\sa10_reg[2]/P0001 ,
		_w2818_,
		_w2819_,
		_w2821_,
		_w2822_
	);
	LUT2 #(
		.INIT('h4)
	) name2290 (
		_w2816_,
		_w2822_,
		_w2823_
	);
	LUT4 #(
		.INIT('h0100)
	) name2291 (
		_w2797_,
		_w2813_,
		_w2807_,
		_w2823_,
		_w2824_
	);
	LUT4 #(
		.INIT('hffda)
	) name2292 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2825_
	);
	LUT2 #(
		.INIT('h2)
	) name2293 (
		\sa03_reg[2]/P0001 ,
		_w2825_,
		_w2826_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name2294 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2827_
	);
	LUT3 #(
		.INIT('h51)
	) name2295 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w2828_
	);
	LUT4 #(
		.INIT('h2022)
	) name2296 (
		\sa03_reg[1]/P0001 ,
		_w1195_,
		_w2827_,
		_w2828_,
		_w2829_
	);
	LUT4 #(
		.INIT('h0040)
	) name2297 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w2830_
	);
	LUT3 #(
		.INIT('h01)
	) name2298 (
		\sa03_reg[1]/P0001 ,
		_w1681_,
		_w2830_,
		_w2831_
	);
	LUT3 #(
		.INIT('h0b)
	) name2299 (
		_w2826_,
		_w2829_,
		_w2831_,
		_w2832_
	);
	LUT3 #(
		.INIT('h80)
	) name2300 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[7]/NET0131 ,
		_w1657_,
		_w2833_
	);
	LUT3 #(
		.INIT('h40)
	) name2301 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1145_,
		_w2834_
	);
	LUT2 #(
		.INIT('h1)
	) name2302 (
		\sa03_reg[0]/P0001 ,
		_w1121_,
		_w2835_
	);
	LUT3 #(
		.INIT('h10)
	) name2303 (
		_w2834_,
		_w2833_,
		_w2835_,
		_w2836_
	);
	LUT2 #(
		.INIT('h4)
	) name2304 (
		_w2832_,
		_w2836_,
		_w2837_
	);
	LUT2 #(
		.INIT('h4)
	) name2305 (
		\sa03_reg[2]/P0001 ,
		_w1135_,
		_w2838_
	);
	LUT3 #(
		.INIT('h01)
	) name2306 (
		\sa03_reg[1]/P0001 ,
		_w1917_,
		_w1900_,
		_w2839_
	);
	LUT4 #(
		.INIT('h0020)
	) name2307 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2840_
	);
	LUT4 #(
		.INIT('h0001)
	) name2308 (
		_w1150_,
		_w1914_,
		_w2648_,
		_w2840_,
		_w2841_
	);
	LUT4 #(
		.INIT('h1000)
	) name2309 (
		_w1908_,
		_w2838_,
		_w2841_,
		_w2839_,
		_w2842_
	);
	LUT4 #(
		.INIT('h0002)
	) name2310 (
		\sa03_reg[2]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2843_
	);
	LUT4 #(
		.INIT('h002a)
	) name2311 (
		\sa03_reg[1]/P0001 ,
		_w1207_,
		_w2499_,
		_w2843_,
		_w2844_
	);
	LUT2 #(
		.INIT('h4)
	) name2312 (
		_w2675_,
		_w2844_,
		_w2845_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name2313 (
		\sa03_reg[4]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2846_
	);
	LUT2 #(
		.INIT('h2)
	) name2314 (
		_w1115_,
		_w2846_,
		_w2847_
	);
	LUT3 #(
		.INIT('h8a)
	) name2315 (
		\sa03_reg[0]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w1145_,
		_w2848_
	);
	LUT4 #(
		.INIT('h153f)
	) name2316 (
		_w1098_,
		_w1045_,
		_w1069_,
		_w1073_,
		_w2849_
	);
	LUT3 #(
		.INIT('h40)
	) name2317 (
		_w2847_,
		_w2848_,
		_w2849_,
		_w2850_
	);
	LUT3 #(
		.INIT('he0)
	) name2318 (
		_w2842_,
		_w2845_,
		_w2850_,
		_w2851_
	);
	LUT4 #(
		.INIT('h0400)
	) name2319 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[4]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		\sa03_reg[7]/NET0131 ,
		_w2852_
	);
	LUT4 #(
		.INIT('h0007)
	) name2320 (
		_w1064_,
		_w1054_,
		_w1112_,
		_w2852_,
		_w2853_
	);
	LUT4 #(
		.INIT('h1113)
	) name2321 (
		\sa03_reg[2]/P0001 ,
		_w1099_,
		_w1049_,
		_w2513_,
		_w2854_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2322 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[2]/P0001 ,
		_w2853_,
		_w2854_,
		_w2855_
	);
	LUT2 #(
		.INIT('h4)
	) name2323 (
		_w1047_,
		_w2479_,
		_w2856_
	);
	LUT3 #(
		.INIT('h02)
	) name2324 (
		\sa03_reg[3]/P0001 ,
		\sa03_reg[5]/P0001 ,
		\sa03_reg[6]/NET0131 ,
		_w2857_
	);
	LUT3 #(
		.INIT('h02)
	) name2325 (
		\sa03_reg[2]/P0001 ,
		_w1681_,
		_w2857_,
		_w2858_
	);
	LUT3 #(
		.INIT('h01)
	) name2326 (
		\sa03_reg[2]/P0001 ,
		_w1145_,
		_w1150_,
		_w2859_
	);
	LUT3 #(
		.INIT('h07)
	) name2327 (
		\sa03_reg[5]/P0001 ,
		_w1130_,
		_w1199_,
		_w2860_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name2328 (
		_w1934_,
		_w2858_,
		_w2859_,
		_w2860_,
		_w2861_
	);
	LUT3 #(
		.INIT('h10)
	) name2329 (
		_w1116_,
		_w2663_,
		_w2676_,
		_w2862_
	);
	LUT3 #(
		.INIT('h80)
	) name2330 (
		\sa03_reg[1]/P0001 ,
		\sa03_reg[2]/P0001 ,
		\sa03_reg[3]/P0001 ,
		_w2863_
	);
	LUT2 #(
		.INIT('h8)
	) name2331 (
		_w1668_,
		_w2863_,
		_w2864_
	);
	LUT3 #(
		.INIT('h01)
	) name2332 (
		_w2537_,
		_w2864_,
		_w2862_,
		_w2865_
	);
	LUT4 #(
		.INIT('hab00)
	) name2333 (
		\sa03_reg[1]/P0001 ,
		_w2856_,
		_w2861_,
		_w2865_,
		_w2866_
	);
	LUT4 #(
		.INIT('h5400)
	) name2334 (
		_w2855_,
		_w2837_,
		_w2851_,
		_w2866_,
		_w2867_
	);
	LUT3 #(
		.INIT('h69)
	) name2335 (
		_w2489_,
		_w2824_,
		_w2867_,
		_w2868_
	);
	LUT4 #(
		.INIT('h0020)
	) name2336 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2869_
	);
	LUT4 #(
		.INIT('h0001)
	) name2337 (
		_w2079_,
		_w2073_,
		_w2348_,
		_w2869_,
		_w2870_
	);
	LUT4 #(
		.INIT('h0111)
	) name2338 (
		\sa21_reg[1]/P0001 ,
		_w1328_,
		_w1391_,
		_w1765_,
		_w2871_
	);
	LUT3 #(
		.INIT('h07)
	) name2339 (
		_w1773_,
		_w1805_,
		_w2091_,
		_w2872_
	);
	LUT3 #(
		.INIT('h80)
	) name2340 (
		_w2870_,
		_w2871_,
		_w2872_,
		_w2873_
	);
	LUT4 #(
		.INIT('hbbf3)
	) name2341 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		_w2874_
	);
	LUT2 #(
		.INIT('h1)
	) name2342 (
		\sa21_reg[2]/P0001 ,
		_w2874_,
		_w2875_
	);
	LUT4 #(
		.INIT('h0002)
	) name2343 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2876_
	);
	LUT4 #(
		.INIT('h002a)
	) name2344 (
		\sa21_reg[1]/P0001 ,
		_w1355_,
		_w2379_,
		_w2876_,
		_w2877_
	);
	LUT2 #(
		.INIT('h4)
	) name2345 (
		_w2875_,
		_w2877_,
		_w2878_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name2346 (
		\sa21_reg[4]/P0001 ,
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2879_
	);
	LUT2 #(
		.INIT('h2)
	) name2347 (
		_w1414_,
		_w2879_,
		_w2880_
	);
	LUT3 #(
		.INIT('h2a)
	) name2348 (
		\sa21_reg[0]/P0001 ,
		_w1326_,
		_w2108_,
		_w2881_
	);
	LUT4 #(
		.INIT('h153f)
	) name2349 (
		\sa21_reg[2]/P0001 ,
		_w1344_,
		_w1394_,
		_w1400_,
		_w2882_
	);
	LUT3 #(
		.INIT('h40)
	) name2350 (
		_w2880_,
		_w2881_,
		_w2882_,
		_w2883_
	);
	LUT3 #(
		.INIT('he0)
	) name2351 (
		_w2873_,
		_w2878_,
		_w2883_,
		_w2884_
	);
	LUT3 #(
		.INIT('h01)
	) name2352 (
		\sa21_reg[1]/P0001 ,
		_w1817_,
		_w2379_,
		_w2885_
	);
	LUT3 #(
		.INIT('h04)
	) name2353 (
		_w1367_,
		_w2351_,
		_w2635_,
		_w2886_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2354 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2887_
	);
	LUT2 #(
		.INIT('h4)
	) name2355 (
		_w2010_,
		_w2887_,
		_w2888_
	);
	LUT2 #(
		.INIT('h2)
	) name2356 (
		\sa21_reg[1]/P0001 ,
		_w1406_,
		_w2889_
	);
	LUT4 #(
		.INIT('h0155)
	) name2357 (
		_w2885_,
		_w2886_,
		_w2888_,
		_w2889_,
		_w2890_
	);
	LUT3 #(
		.INIT('h80)
	) name2358 (
		\sa21_reg[2]/P0001 ,
		_w1330_,
		_w1391_,
		_w2891_
	);
	LUT4 #(
		.INIT('h0111)
	) name2359 (
		\sa21_reg[0]/P0001 ,
		_w1335_,
		_w1425_,
		_w1427_,
		_w2892_
	);
	LUT2 #(
		.INIT('h4)
	) name2360 (
		_w2891_,
		_w2892_,
		_w2893_
	);
	LUT2 #(
		.INIT('h4)
	) name2361 (
		_w2890_,
		_w2893_,
		_w2894_
	);
	LUT4 #(
		.INIT('h0111)
	) name2362 (
		\sa21_reg[2]/P0001 ,
		_w1328_,
		_w1379_,
		_w1380_,
		_w2895_
	);
	LUT2 #(
		.INIT('h1)
	) name2363 (
		_w1427_,
		_w1410_,
		_w2896_
	);
	LUT3 #(
		.INIT('h02)
	) name2364 (
		\sa21_reg[2]/P0001 ,
		_w1817_,
		_w2035_,
		_w2897_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name2365 (
		_w2106_,
		_w2895_,
		_w2896_,
		_w2897_,
		_w2898_
	);
	LUT3 #(
		.INIT('h01)
	) name2366 (
		\sa21_reg[1]/P0001 ,
		_w1825_,
		_w2089_,
		_w2899_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2367 (
		\sa21_reg[2]/P0001 ,
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[7]/P0001 ,
		_w2900_
	);
	LUT4 #(
		.INIT('h1300)
	) name2368 (
		_w1345_,
		_w1395_,
		_w1380_,
		_w2900_,
		_w2901_
	);
	LUT4 #(
		.INIT('h0400)
	) name2369 (
		\sa21_reg[3]/P0001 ,
		\sa21_reg[4]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2902_
	);
	LUT2 #(
		.INIT('h1)
	) name2370 (
		\sa21_reg[2]/P0001 ,
		_w2902_,
		_w2903_
	);
	LUT2 #(
		.INIT('h2)
	) name2371 (
		\sa21_reg[1]/P0001 ,
		_w2028_,
		_w2904_
	);
	LUT4 #(
		.INIT('hec00)
	) name2372 (
		_w2691_,
		_w2901_,
		_w2903_,
		_w2904_,
		_w2905_
	);
	LUT3 #(
		.INIT('had)
	) name2373 (
		\sa21_reg[5]/P0001 ,
		\sa21_reg[6]/NET0131 ,
		\sa21_reg[7]/P0001 ,
		_w2906_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2374 (
		_w1425_,
		_w1770_,
		_w2089_,
		_w2906_,
		_w2907_
	);
	LUT4 #(
		.INIT('hf400)
	) name2375 (
		_w2898_,
		_w2899_,
		_w2905_,
		_w2907_,
		_w2908_
	);
	LUT3 #(
		.INIT('he0)
	) name2376 (
		_w2884_,
		_w2894_,
		_w2908_,
		_w2909_
	);
	LUT4 #(
		.INIT('ha955)
	) name2377 (
		\u0_w_reg[3][2]/P0001 ,
		_w2884_,
		_w2894_,
		_w2908_,
		_w2910_
	);
	LUT2 #(
		.INIT('h6)
	) name2378 (
		_w2341_,
		_w2910_,
		_w2911_
	);
	LUT3 #(
		.INIT('h28)
	) name2379 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[2]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		_w2912_
	);
	LUT4 #(
		.INIT('hff41)
	) name2380 (
		\ld_r_reg/P0001 ,
		_w2868_,
		_w2911_,
		_w2912_,
		_w2913_
	);
	LUT4 #(
		.INIT('h6996)
	) name2381 (
		\u0_w_reg[3][25]/P0001 ,
		_w2341_,
		_w2437_,
		_w2732_,
		_w2914_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name2382 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2915_
	);
	LUT2 #(
		.INIT('h2)
	) name2383 (
		\sa10_reg[2]/P0001 ,
		_w2915_,
		_w2916_
	);
	LUT3 #(
		.INIT('h54)
	) name2384 (
		\sa10_reg[3]/P0001 ,
		_w1568_,
		_w1976_,
		_w2917_
	);
	LUT3 #(
		.INIT('h20)
	) name2385 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w1594_,
		_w2918_
	);
	LUT3 #(
		.INIT('h8a)
	) name2386 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2919_
	);
	LUT2 #(
		.INIT('h2)
	) name2387 (
		_w1224_,
		_w2919_,
		_w2920_
	);
	LUT4 #(
		.INIT('h0001)
	) name2388 (
		_w2918_,
		_w2916_,
		_w2917_,
		_w2920_,
		_w2921_
	);
	LUT3 #(
		.INIT('h07)
	) name2389 (
		\sa10_reg[7]/NET0131 ,
		_w1247_,
		_w1881_,
		_w2922_
	);
	LUT3 #(
		.INIT('h2a)
	) name2390 (
		\sa10_reg[2]/P0001 ,
		_w1229_,
		_w2922_,
		_w2923_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name2391 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2924_
	);
	LUT4 #(
		.INIT('h0301)
	) name2392 (
		\sa10_reg[3]/P0001 ,
		_w1572_,
		_w1597_,
		_w2924_,
		_w2925_
	);
	LUT4 #(
		.INIT('h4041)
	) name2393 (
		\sa10_reg[2]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2926_
	);
	LUT3 #(
		.INIT('ha8)
	) name2394 (
		\sa10_reg[1]/P0001 ,
		_w1295_,
		_w2926_,
		_w2927_
	);
	LUT3 #(
		.INIT('h0b)
	) name2395 (
		\sa10_reg[4]/P0001 ,
		_w1256_,
		_w2395_,
		_w2928_
	);
	LUT4 #(
		.INIT('h3200)
	) name2396 (
		\sa10_reg[2]/P0001 ,
		_w2927_,
		_w2925_,
		_w2928_,
		_w2929_
	);
	LUT4 #(
		.INIT('h3200)
	) name2397 (
		\sa10_reg[1]/P0001 ,
		_w2923_,
		_w2921_,
		_w2929_,
		_w2930_
	);
	LUT4 #(
		.INIT('h0001)
	) name2398 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		_w2931_
	);
	LUT4 #(
		.INIT('h0007)
	) name2399 (
		\sa10_reg[7]/NET0131 ,
		_w1247_,
		_w2559_,
		_w2931_,
		_w2932_
	);
	LUT2 #(
		.INIT('h1)
	) name2400 (
		\sa10_reg[2]/P0001 ,
		_w2932_,
		_w2933_
	);
	LUT2 #(
		.INIT('h1)
	) name2401 (
		\sa10_reg[3]/P0001 ,
		_w1578_,
		_w2934_
	);
	LUT4 #(
		.INIT('h8007)
	) name2402 (
		\sa10_reg[3]/P0001 ,
		\sa10_reg[4]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2935_
	);
	LUT4 #(
		.INIT('h020a)
	) name2403 (
		\sa10_reg[1]/P0001 ,
		_w1269_,
		_w1594_,
		_w1885_,
		_w2936_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name2404 (
		_w1863_,
		_w2934_,
		_w2935_,
		_w2936_,
		_w2937_
	);
	LUT3 #(
		.INIT('hb9)
	) name2405 (
		\sa10_reg[5]/P0001 ,
		\sa10_reg[6]/NET0131 ,
		\sa10_reg[7]/NET0131 ,
		_w2938_
	);
	LUT3 #(
		.INIT('h40)
	) name2406 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[2]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w2939_
	);
	LUT4 #(
		.INIT('h31f5)
	) name2407 (
		_w1301_,
		_w2391_,
		_w2938_,
		_w2939_,
		_w2940_
	);
	LUT3 #(
		.INIT('h10)
	) name2408 (
		_w2937_,
		_w2933_,
		_w2940_,
		_w2941_
	);
	LUT4 #(
		.INIT('h000b)
	) name2409 (
		\sa10_reg[4]/P0001 ,
		_w1236_,
		_w1589_,
		_w1958_,
		_w2942_
	);
	LUT4 #(
		.INIT('h0302)
	) name2410 (
		\sa10_reg[2]/P0001 ,
		_w1998_,
		_w2789_,
		_w2942_,
		_w2943_
	);
	LUT4 #(
		.INIT('h3230)
	) name2411 (
		\sa10_reg[4]/P0001 ,
		\sa10_reg[5]/P0001 ,
		_w1318_,
		_w1844_,
		_w2944_
	);
	LUT3 #(
		.INIT('hd8)
	) name2412 (
		\sa10_reg[2]/P0001 ,
		_w1256_,
		_w1607_,
		_w2945_
	);
	LUT3 #(
		.INIT('h01)
	) name2413 (
		_w1312_,
		_w2944_,
		_w2945_,
		_w2946_
	);
	LUT2 #(
		.INIT('h8)
	) name2414 (
		\sa10_reg[6]/NET0131 ,
		_w1263_,
		_w2947_
	);
	LUT3 #(
		.INIT('h8a)
	) name2415 (
		\sa10_reg[1]/P0001 ,
		\sa10_reg[7]/NET0131 ,
		_w1297_,
		_w2948_
	);
	LUT4 #(
		.INIT('haa80)
	) name2416 (
		\sa10_reg[2]/P0001 ,
		_w1286_,
		_w1271_,
		_w1297_,
		_w2949_
	);
	LUT3 #(
		.INIT('h45)
	) name2417 (
		_w2947_,
		_w2948_,
		_w2949_,
		_w2950_
	);
	LUT4 #(
		.INIT('he400)
	) name2418 (
		\sa10_reg[1]/P0001 ,
		_w2943_,
		_w2946_,
		_w2950_,
		_w2951_
	);
	LUT4 #(
		.INIT('hd800)
	) name2419 (
		\sa10_reg[0]/P0001 ,
		_w2930_,
		_w2941_,
		_w2951_,
		_w2952_
	);
	LUT4 #(
		.INIT('h9669)
	) name2420 (
		_w1619_,
		_w1685_,
		_w2685_,
		_w2952_,
		_w2953_
	);
	LUT3 #(
		.INIT('h28)
	) name2421 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[25]/P0001 ,
		\u0_w_reg[3][25]/P0001 ,
		_w2954_
	);
	LUT4 #(
		.INIT('hff14)
	) name2422 (
		\ld_r_reg/P0001 ,
		_w2914_,
		_w2953_,
		_w2954_,
		_w2955_
	);
	LUT3 #(
		.INIT('h69)
	) name2423 (
		_w1438_,
		_w1619_,
		_w1685_,
		_w2956_
	);
	LUT4 #(
		.INIT('h5655)
	) name2424 (
		\u0_w_reg[3][15]/P0001 ,
		_w2280_,
		_w2261_,
		_w2297_,
		_w2957_
	);
	LUT2 #(
		.INIT('h6)
	) name2425 (
		_w1759_,
		_w2957_,
		_w2958_
	);
	LUT3 #(
		.INIT('h82)
	) name2426 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[15]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w2959_
	);
	LUT4 #(
		.INIT('h00eb)
	) name2427 (
		\ld_r_reg/P0001 ,
		_w2956_,
		_w2958_,
		_w2959_,
		_w2960_
	);
	LUT4 #(
		.INIT('h6996)
	) name2428 (
		_w1685_,
		_w1895_,
		_w1948_,
		_w2547_,
		_w2961_
	);
	LUT4 #(
		.INIT('h6996)
	) name2429 (
		\u0_w_reg[3][4]/P0001 ,
		_w2121_,
		_w2298_,
		_w2779_,
		_w2962_
	);
	LUT3 #(
		.INIT('h82)
	) name2430 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[4]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w2963_
	);
	LUT4 #(
		.INIT('h00eb)
	) name2431 (
		\ld_r_reg/P0001 ,
		_w2961_,
		_w2962_,
		_w2963_,
		_w2964_
	);
	LUT4 #(
		.INIT('h5655)
	) name2432 (
		\u0_w_reg[3][27]/P0001 ,
		_w2766_,
		_w2750_,
		_w2778_,
		_w2965_
	);
	LUT3 #(
		.INIT('h69)
	) name2433 (
		_w2592_,
		_w2641_,
		_w2965_,
		_w2966_
	);
	LUT4 #(
		.INIT('h9669)
	) name2434 (
		_w1619_,
		_w1685_,
		_w2824_,
		_w2867_,
		_w2967_
	);
	LUT3 #(
		.INIT('h82)
	) name2435 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[27]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w2968_
	);
	LUT4 #(
		.INIT('h00be)
	) name2436 (
		\ld_r_reg/P0001 ,
		_w2966_,
		_w2967_,
		_w2968_,
		_w2969_
	);
	LUT4 #(
		.INIT('h5655)
	) name2437 (
		\u0_w_reg[3][19]/P0001 ,
		_w2766_,
		_w2750_,
		_w2778_,
		_w2970_
	);
	LUT3 #(
		.INIT('h69)
	) name2438 (
		_w1830_,
		_w2641_,
		_w2970_,
		_w2971_
	);
	LUT4 #(
		.INIT('h6996)
	) name2439 (
		_w1619_,
		_w2547_,
		_w2824_,
		_w2909_,
		_w2972_
	);
	LUT3 #(
		.INIT('h82)
	) name2440 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[19]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w2973_
	);
	LUT4 #(
		.INIT('h00eb)
	) name2441 (
		\ld_r_reg/P0001 ,
		_w2971_,
		_w2972_,
		_w2973_,
		_w2974_
	);
	LUT4 #(
		.INIT('h6996)
	) name2442 (
		_w1619_,
		_w2388_,
		_w2489_,
		_w2952_,
		_w2975_
	);
	LUT4 #(
		.INIT('h5655)
	) name2443 (
		\u0_w_reg[3][17]/P0001 ,
		_w2715_,
		_w2699_,
		_w2731_,
		_w2976_
	);
	LUT3 #(
		.INIT('h96)
	) name2444 (
		_w1830_,
		_w2341_,
		_w2976_,
		_w2977_
	);
	LUT3 #(
		.INIT('h28)
	) name2445 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[17]/P0001 ,
		\u0_w_reg[3][17]/P0001 ,
		_w2978_
	);
	LUT4 #(
		.INIT('hff14)
	) name2446 (
		\ld_r_reg/P0001 ,
		_w2975_,
		_w2977_,
		_w2978_,
		_w2979_
	);
	LUT4 #(
		.INIT('h6996)
	) name2447 (
		_w1830_,
		_w2547_,
		_w2592_,
		_w2909_,
		_w2980_
	);
	LUT4 #(
		.INIT('h000b)
	) name2448 (
		\sa32_reg[2]/P0001 ,
		_w1527_,
		_w2175_,
		_w2198_,
		_w2981_
	);
	LUT3 #(
		.INIT('h01)
	) name2449 (
		\sa32_reg[1]/P0001 ,
		_w1687_,
		_w2168_,
		_w2982_
	);
	LUT4 #(
		.INIT('h8adf)
	) name2450 (
		\sa32_reg[2]/P0001 ,
		_w1483_,
		_w1439_,
		_w1535_,
		_w2983_
	);
	LUT3 #(
		.INIT('h80)
	) name2451 (
		_w2981_,
		_w2982_,
		_w2983_,
		_w2984_
	);
	LUT3 #(
		.INIT('h15)
	) name2452 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		_w2985_
	);
	LUT2 #(
		.INIT('h8)
	) name2453 (
		_w2250_,
		_w2985_,
		_w2986_
	);
	LUT4 #(
		.INIT('h020a)
	) name2454 (
		\sa32_reg[1]/P0001 ,
		_w1499_,
		_w1738_,
		_w2216_,
		_w2987_
	);
	LUT2 #(
		.INIT('h4)
	) name2455 (
		_w2986_,
		_w2987_,
		_w2988_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name2456 (
		\sa32_reg[4]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2989_
	);
	LUT2 #(
		.INIT('h2)
	) name2457 (
		_w1546_,
		_w2989_,
		_w2990_
	);
	LUT3 #(
		.INIT('h54)
	) name2458 (
		\sa32_reg[3]/P0001 ,
		_w1542_,
		_w2153_,
		_w2991_
	);
	LUT3 #(
		.INIT('h2a)
	) name2459 (
		\sa32_reg[0]/P0002 ,
		_w1444_,
		_w1746_,
		_w2992_
	);
	LUT3 #(
		.INIT('h10)
	) name2460 (
		_w2990_,
		_w2991_,
		_w2992_,
		_w2993_
	);
	LUT3 #(
		.INIT('he0)
	) name2461 (
		_w2984_,
		_w2988_,
		_w2993_,
		_w2994_
	);
	LUT4 #(
		.INIT('hffda)
	) name2462 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2995_
	);
	LUT2 #(
		.INIT('h2)
	) name2463 (
		\sa32_reg[2]/P0001 ,
		_w2995_,
		_w2996_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name2464 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w2997_
	);
	LUT3 #(
		.INIT('h51)
	) name2465 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[5]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w2998_
	);
	LUT4 #(
		.INIT('h2022)
	) name2466 (
		\sa32_reg[1]/P0001 ,
		_w1733_,
		_w2997_,
		_w2998_,
		_w2999_
	);
	LUT3 #(
		.INIT('h01)
	) name2467 (
		\sa32_reg[1]/P0001 ,
		_w1510_,
		_w2216_,
		_w3000_
	);
	LUT3 #(
		.INIT('h0b)
	) name2468 (
		_w2996_,
		_w2999_,
		_w3000_,
		_w3001_
	);
	LUT3 #(
		.INIT('h80)
	) name2469 (
		\sa32_reg[6]/NET0131 ,
		_w1546_,
		_w2155_,
		_w3002_
	);
	LUT2 #(
		.INIT('h1)
	) name2470 (
		\sa32_reg[0]/P0002 ,
		_w1492_,
		_w3003_
	);
	LUT3 #(
		.INIT('h10)
	) name2471 (
		_w1751_,
		_w3002_,
		_w3003_,
		_w3004_
	);
	LUT2 #(
		.INIT('h4)
	) name2472 (
		_w3001_,
		_w3004_,
		_w3005_
	);
	LUT4 #(
		.INIT('h0013)
	) name2473 (
		_w1449_,
		_w1470_,
		_w1689_,
		_w2283_,
		_w3006_
	);
	LUT4 #(
		.INIT('h0203)
	) name2474 (
		\sa32_reg[4]/P0001 ,
		_w1527_,
		_w1532_,
		_w1748_,
		_w3007_
	);
	LUT2 #(
		.INIT('h2)
	) name2475 (
		\sa32_reg[1]/P0001 ,
		_w1454_,
		_w3008_
	);
	LUT4 #(
		.INIT('hd800)
	) name2476 (
		\sa32_reg[2]/P0001 ,
		_w3007_,
		_w3006_,
		_w3008_,
		_w3009_
	);
	LUT4 #(
		.INIT('h0007)
	) name2477 (
		\sa32_reg[6]/NET0131 ,
		_w1521_,
		_w1742_,
		_w2281_,
		_w3010_
	);
	LUT3 #(
		.INIT('h13)
	) name2478 (
		_w1467_,
		_w1461_,
		_w1475_,
		_w3011_
	);
	LUT4 #(
		.INIT('h135f)
	) name2479 (
		_w1688_,
		_w2286_,
		_w3010_,
		_w3011_,
		_w3012_
	);
	LUT3 #(
		.INIT('hb8)
	) name2480 (
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		\sa32_reg[7]/P0001 ,
		_w3013_
	);
	LUT3 #(
		.INIT('h15)
	) name2481 (
		\sa32_reg[1]/P0001 ,
		_w1460_,
		_w3013_,
		_w3014_
	);
	LUT3 #(
		.INIT('had)
	) name2482 (
		\sa32_reg[5]/P0001 ,
		\sa32_reg[6]/NET0131 ,
		\sa32_reg[7]/P0001 ,
		_w3015_
	);
	LUT3 #(
		.INIT('h02)
	) name2483 (
		\sa32_reg[2]/P0001 ,
		\sa32_reg[3]/P0001 ,
		\sa32_reg[4]/P0001 ,
		_w3016_
	);
	LUT4 #(
		.INIT('h7077)
	) name2484 (
		_w1514_,
		_w1489_,
		_w3015_,
		_w3016_,
		_w3017_
	);
	LUT4 #(
		.INIT('hba00)
	) name2485 (
		_w3009_,
		_w3012_,
		_w3014_,
		_w3017_,
		_w3018_
	);
	LUT4 #(
		.INIT('ha955)
	) name2486 (
		\u0_w_reg[3][11]/P0001 ,
		_w2994_,
		_w3005_,
		_w3018_,
		_w3019_
	);
	LUT3 #(
		.INIT('h69)
	) name2487 (
		_w2298_,
		_w2779_,
		_w3019_,
		_w3020_
	);
	LUT3 #(
		.INIT('h82)
	) name2488 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[11]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w3021_
	);
	LUT4 #(
		.INIT('h00eb)
	) name2489 (
		\ld_r_reg/P0001 ,
		_w2980_,
		_w3020_,
		_w3021_,
		_w3022_
	);
	LUT4 #(
		.INIT('ha955)
	) name2490 (
		\u0_w_reg[3][26]/P0001 ,
		_w2994_,
		_w3005_,
		_w3018_,
		_w3023_
	);
	LUT3 #(
		.INIT('h69)
	) name2491 (
		_w2824_,
		_w2909_,
		_w3023_,
		_w3024_
	);
	LUT3 #(
		.INIT('h82)
	) name2492 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[26]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		_w3025_
	);
	LUT4 #(
		.INIT('h00eb)
	) name2493 (
		\ld_r_reg/P0001 ,
		_w2490_,
		_w3024_,
		_w3025_,
		_w3026_
	);
	LUT4 #(
		.INIT('h6996)
	) name2494 (
		_w1685_,
		_w2547_,
		_w2592_,
		_w2867_,
		_w3027_
	);
	LUT4 #(
		.INIT('ha955)
	) name2495 (
		\u0_w_reg[3][3]/P0001 ,
		_w2994_,
		_w3005_,
		_w3018_,
		_w3028_
	);
	LUT3 #(
		.INIT('h96)
	) name2496 (
		_w2298_,
		_w2641_,
		_w3028_,
		_w3029_
	);
	LUT3 #(
		.INIT('h82)
	) name2497 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[3]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w3030_
	);
	LUT4 #(
		.INIT('h00be)
	) name2498 (
		\ld_r_reg/P0001 ,
		_w3027_,
		_w3029_,
		_w3030_,
		_w3031_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name2499 (
		\u0_w_reg[3][24]/P0001 ,
		_w2212_,
		_w2222_,
		_w2243_,
		_w3032_
	);
	LUT4 #(
		.INIT('h9669)
	) name2500 (
		_w1619_,
		_w1685_,
		_w2388_,
		_w2952_,
		_w3033_
	);
	LUT3 #(
		.INIT('h28)
	) name2501 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[24]/P0001 ,
		\u0_w_reg[3][24]/P0001 ,
		_w3034_
	);
	LUT4 #(
		.INIT('hff14)
	) name2502 (
		\ld_r_reg/P0001 ,
		_w3032_,
		_w3033_,
		_w3034_,
		_w3035_
	);
	LUT4 #(
		.INIT('h6996)
	) name2503 (
		\u0_w_reg[3][31]/P0001 ,
		_w1619_,
		_w1830_,
		_w2298_,
		_w3036_
	);
	LUT3 #(
		.INIT('h28)
	) name2504 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[31]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w3037_
	);
	LUT4 #(
		.INIT('hff41)
	) name2505 (
		\ld_r_reg/P0001 ,
		_w1324_,
		_w3036_,
		_w3037_,
		_w3038_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name2506 (
		\u0_w_reg[3][16]/P0001 ,
		_w2212_,
		_w2222_,
		_w2243_,
		_w3039_
	);
	LUT4 #(
		.INIT('h6996)
	) name2507 (
		_w1619_,
		_w1830_,
		_w2388_,
		_w2685_,
		_w3040_
	);
	LUT3 #(
		.INIT('h28)
	) name2508 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[16]/P0001 ,
		\u0_w_reg[3][16]/P0001 ,
		_w3041_
	);
	LUT4 #(
		.INIT('hff41)
	) name2509 (
		\ld_r_reg/P0001 ,
		_w3039_,
		_w3040_,
		_w3041_,
		_w3042_
	);
	LUT3 #(
		.INIT('h69)
	) name2510 (
		_w2437_,
		_w2732_,
		_w2867_,
		_w3043_
	);
	LUT4 #(
		.INIT('ha955)
	) name2511 (
		\u0_w_reg[3][18]/P0001 ,
		_w2994_,
		_w3005_,
		_w3018_,
		_w3044_
	);
	LUT2 #(
		.INIT('h6)
	) name2512 (
		_w2909_,
		_w3044_,
		_w3045_
	);
	LUT3 #(
		.INIT('h82)
	) name2513 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[18]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		_w3046_
	);
	LUT4 #(
		.INIT('h00eb)
	) name2514 (
		\ld_r_reg/P0001 ,
		_w3043_,
		_w3045_,
		_w3046_,
		_w3047_
	);
	LUT3 #(
		.INIT('h69)
	) name2515 (
		_w1323_,
		_w1438_,
		_w1685_,
		_w3048_
	);
	LUT3 #(
		.INIT('h69)
	) name2516 (
		\u0_w_reg[3][23]/P0001 ,
		_w1830_,
		_w2298_,
		_w3049_
	);
	LUT3 #(
		.INIT('h82)
	) name2517 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[23]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w3050_
	);
	LUT4 #(
		.INIT('h00eb)
	) name2518 (
		\ld_r_reg/P0001 ,
		_w3048_,
		_w3049_,
		_w3050_,
		_w3051_
	);
	LUT3 #(
		.INIT('h69)
	) name2519 (
		_w2732_,
		_w2824_,
		_w2867_,
		_w3052_
	);
	LUT4 #(
		.INIT('ha955)
	) name2520 (
		\u0_w_reg[3][10]/P0001 ,
		_w2994_,
		_w3005_,
		_w3018_,
		_w3053_
	);
	LUT2 #(
		.INIT('h6)
	) name2521 (
		_w2341_,
		_w3053_,
		_w3054_
	);
	LUT3 #(
		.INIT('h82)
	) name2522 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[10]/P0001 ,
		\u0_w_reg[3][10]/P0001 ,
		_w3055_
	);
	LUT4 #(
		.INIT('h00eb)
	) name2523 (
		\ld_r_reg/P0001 ,
		_w3052_,
		_w3054_,
		_w3055_,
		_w3056_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name2524 (
		\u0_w_reg[3][8]/P0001 ,
		_w2212_,
		_w2222_,
		_w2243_,
		_w3057_
	);
	LUT4 #(
		.INIT('h9669)
	) name2525 (
		_w1830_,
		_w2298_,
		_w2685_,
		_w2952_,
		_w3058_
	);
	LUT3 #(
		.INIT('h82)
	) name2526 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[8]/P0001 ,
		\u0_w_reg[3][8]/P0001 ,
		_w3059_
	);
	LUT4 #(
		.INIT('h00be)
	) name2527 (
		\ld_r_reg/P0001 ,
		_w3057_,
		_w3058_,
		_w3059_,
		_w3060_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name2528 (
		\u0_w_reg[3][0]/P0001 ,
		_w2280_,
		_w2261_,
		_w2297_,
		_w3061_
	);
	LUT4 #(
		.INIT('h9669)
	) name2529 (
		_w1685_,
		_w2388_,
		_w2685_,
		_w2952_,
		_w3062_
	);
	LUT3 #(
		.INIT('h28)
	) name2530 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[0]/P0001 ,
		\u0_w_reg[3][0]/P0001 ,
		_w3063_
	);
	LUT4 #(
		.INIT('hff14)
	) name2531 (
		\ld_r_reg/P0001 ,
		_w3061_,
		_w3062_,
		_w3063_,
		_w3064_
	);
	LUT3 #(
		.INIT('h65)
	) name2532 (
		\u0_w_reg[3][5]/P0001 ,
		_w1497_,
		_w1552_,
		_w3065_
	);
	LUT4 #(
		.INIT('h5655)
	) name2533 (
		\u0_w_reg[3][6]/P0001 ,
		_w1707_,
		_w1732_,
		_w1758_,
		_w3066_
	);
	LUT2 #(
		.INIT('h9)
	) name2534 (
		\u0_w_reg[3][4]/P0001 ,
		_w2185_,
		_w3067_
	);
	LUT4 #(
		.INIT('h5655)
	) name2535 (
		\u0_w_reg[3][0]/P0001 ,
		_w2212_,
		_w2222_,
		_w2243_,
		_w3068_
	);
	LUT4 #(
		.INIT('h5655)
	) name2536 (
		\u0_w_reg[3][3]/P0001 ,
		_w2766_,
		_w2750_,
		_w2778_,
		_w3069_
	);
	LUT2 #(
		.INIT('h9)
	) name2537 (
		\u0_w_reg[3][1]/P0001 ,
		_w2341_,
		_w3070_
	);
	LUT4 #(
		.INIT('ha955)
	) name2538 (
		\u0_w_reg[3][2]/P0001 ,
		_w2994_,
		_w3005_,
		_w3018_,
		_w3071_
	);
	LUT4 #(
		.INIT('h5655)
	) name2539 (
		\u0_w_reg[3][7]/P0001 ,
		_w2280_,
		_w2261_,
		_w2297_,
		_w3072_
	);
	LUT4 #(
		.INIT('h0004)
	) name2540 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3073_
	);
	LUT4 #(
		.INIT('h5554)
	) name2541 (
		\sa02_reg[2]/P0001 ,
		_w895_,
		_w896_,
		_w3073_,
		_w3074_
	);
	LUT3 #(
		.INIT('h54)
	) name2542 (
		\sa02_reg[1]/P0001 ,
		_w904_,
		_w3074_,
		_w3075_
	);
	LUT4 #(
		.INIT('h0100)
	) name2543 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w3076_
	);
	LUT3 #(
		.INIT('h08)
	) name2544 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3077_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name2545 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3078_
	);
	LUT4 #(
		.INIT('h80aa)
	) name2546 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3076_,
		_w3078_,
		_w3079_
	);
	LUT4 #(
		.INIT('h0001)
	) name2547 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3080_
	);
	LUT4 #(
		.INIT('h0007)
	) name2548 (
		_w831_,
		_w832_,
		_w911_,
		_w3080_,
		_w3081_
	);
	LUT3 #(
		.INIT('h8a)
	) name2549 (
		\sa02_reg[2]/P0001 ,
		_w3079_,
		_w3081_,
		_w3082_
	);
	LUT4 #(
		.INIT('h2000)
	) name2550 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3083_
	);
	LUT3 #(
		.INIT('h0b)
	) name2551 (
		\sa02_reg[6]/NET0131 ,
		_w852_,
		_w3083_,
		_w3084_
	);
	LUT4 #(
		.INIT('haa20)
	) name2552 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w852_,
		_w3083_,
		_w3085_
	);
	LUT2 #(
		.INIT('h4)
	) name2553 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		_w3086_
	);
	LUT3 #(
		.INIT('he0)
	) name2554 (
		_w878_,
		_w915_,
		_w3086_,
		_w3087_
	);
	LUT4 #(
		.INIT('h0040)
	) name2555 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3088_
	);
	LUT3 #(
		.INIT('h54)
	) name2556 (
		\sa02_reg[2]/P0001 ,
		_w868_,
		_w3088_,
		_w3089_
	);
	LUT2 #(
		.INIT('h2)
	) name2557 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		_w3090_
	);
	LUT2 #(
		.INIT('h1)
	) name2558 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		_w3091_
	);
	LUT4 #(
		.INIT('h080a)
	) name2559 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w3092_
	);
	LUT4 #(
		.INIT('h0777)
	) name2560 (
		_w869_,
		_w3090_,
		_w3091_,
		_w3092_,
		_w3093_
	);
	LUT4 #(
		.INIT('h0100)
	) name2561 (
		_w3089_,
		_w3085_,
		_w3087_,
		_w3093_,
		_w3094_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2562 (
		\sa02_reg[0]/P0001 ,
		_w3082_,
		_w3075_,
		_w3094_,
		_w3095_
	);
	LUT2 #(
		.INIT('h2)
	) name2563 (
		_w833_,
		_w902_,
		_w3096_
	);
	LUT4 #(
		.INIT('h0001)
	) name2564 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3097_
	);
	LUT2 #(
		.INIT('h4)
	) name2565 (
		\sa02_reg[4]/P0001 ,
		_w3097_,
		_w3098_
	);
	LUT3 #(
		.INIT('h2a)
	) name2566 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w852_,
		_w3099_
	);
	LUT3 #(
		.INIT('h10)
	) name2567 (
		_w3098_,
		_w3096_,
		_w3099_,
		_w3100_
	);
	LUT2 #(
		.INIT('h8)
	) name2568 (
		\sa02_reg[4]/P0001 ,
		_w883_,
		_w3101_
	);
	LUT4 #(
		.INIT('h4000)
	) name2569 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3102_
	);
	LUT4 #(
		.INIT('h0100)
	) name2570 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3103_
	);
	LUT4 #(
		.INIT('h0200)
	) name2571 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3104_
	);
	LUT3 #(
		.INIT('h01)
	) name2572 (
		_w3103_,
		_w3104_,
		_w3102_,
		_w3105_
	);
	LUT3 #(
		.INIT('h08)
	) name2573 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3106_
	);
	LUT4 #(
		.INIT('h0105)
	) name2574 (
		\sa02_reg[1]/P0001 ,
		_w905_,
		_w3088_,
		_w3106_,
		_w3107_
	);
	LUT3 #(
		.INIT('h40)
	) name2575 (
		_w3101_,
		_w3105_,
		_w3107_,
		_w3108_
	);
	LUT4 #(
		.INIT('h2220)
	) name2576 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3109_
	);
	LUT3 #(
		.INIT('h2a)
	) name2577 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3110_
	);
	LUT2 #(
		.INIT('h2)
	) name2578 (
		_w3109_,
		_w3110_,
		_w3111_
	);
	LUT4 #(
		.INIT('h4000)
	) name2579 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w3112_
	);
	LUT4 #(
		.INIT('h0405)
	) name2580 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w855_,
		_w3112_,
		_w3113_
	);
	LUT4 #(
		.INIT('h0001)
	) name2581 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w3114_
	);
	LUT4 #(
		.INIT('h002a)
	) name2582 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w883_,
		_w3114_,
		_w3115_
	);
	LUT3 #(
		.INIT('h0b)
	) name2583 (
		_w3111_,
		_w3113_,
		_w3115_,
		_w3116_
	);
	LUT4 #(
		.INIT('h5501)
	) name2584 (
		\sa02_reg[0]/P0001 ,
		_w3100_,
		_w3108_,
		_w3116_,
		_w3117_
	);
	LUT4 #(
		.INIT('h0020)
	) name2585 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3118_
	);
	LUT4 #(
		.INIT('h0800)
	) name2586 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3119_
	);
	LUT4 #(
		.INIT('h5554)
	) name2587 (
		\sa02_reg[2]/P0001 ,
		_w904_,
		_w3119_,
		_w3118_,
		_w3120_
	);
	LUT4 #(
		.INIT('h4000)
	) name2588 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3121_
	);
	LUT2 #(
		.INIT('h8)
	) name2589 (
		\sa02_reg[2]/P0001 ,
		_w3121_,
		_w3122_
	);
	LUT2 #(
		.INIT('h2)
	) name2590 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w3123_
	);
	LUT4 #(
		.INIT('h0002)
	) name2591 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3124_
	);
	LUT4 #(
		.INIT('h0800)
	) name2592 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3125_
	);
	LUT4 #(
		.INIT('h1000)
	) name2593 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w3126_
	);
	LUT4 #(
		.INIT('h0013)
	) name2594 (
		\sa02_reg[3]/P0001 ,
		_w3125_,
		_w3124_,
		_w3126_,
		_w3127_
	);
	LUT4 #(
		.INIT('h5455)
	) name2595 (
		\sa02_reg[1]/P0001 ,
		_w3120_,
		_w3122_,
		_w3127_,
		_w3128_
	);
	LUT2 #(
		.INIT('h8)
	) name2596 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		_w3129_
	);
	LUT4 #(
		.INIT('hf7fa)
	) name2597 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3130_
	);
	LUT2 #(
		.INIT('h2)
	) name2598 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w3131_
	);
	LUT4 #(
		.INIT('h0002)
	) name2599 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3132_
	);
	LUT4 #(
		.INIT('hcc04)
	) name2600 (
		\sa02_reg[4]/P0001 ,
		_w3129_,
		_w3130_,
		_w3132_,
		_w3133_
	);
	LUT2 #(
		.INIT('h8)
	) name2601 (
		_w904_,
		_w829_,
		_w3134_
	);
	LUT2 #(
		.INIT('h4)
	) name2602 (
		\sa02_reg[7]/NET0131 ,
		_w3114_,
		_w3135_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name2603 (
		\sa02_reg[7]/NET0131 ,
		_w833_,
		_w889_,
		_w3114_,
		_w3136_
	);
	LUT2 #(
		.INIT('h2)
	) name2604 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		_w3137_
	);
	LUT3 #(
		.INIT('h80)
	) name2605 (
		_w847_,
		_w923_,
		_w3137_,
		_w3138_
	);
	LUT2 #(
		.INIT('h8)
	) name2606 (
		_w891_,
		_w3118_,
		_w3139_
	);
	LUT4 #(
		.INIT('h0100)
	) name2607 (
		_w3138_,
		_w3134_,
		_w3139_,
		_w3136_,
		_w3140_
	);
	LUT3 #(
		.INIT('h10)
	) name2608 (
		_w3133_,
		_w3128_,
		_w3140_,
		_w3141_
	);
	LUT3 #(
		.INIT('h10)
	) name2609 (
		_w3095_,
		_w3117_,
		_w3141_,
		_w3142_
	);
	LUT3 #(
		.INIT('h69)
	) name2610 (
		_w637_,
		_w933_,
		_w3142_,
		_w3143_
	);
	LUT4 #(
		.INIT('hf7a7)
	) name2611 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3144_
	);
	LUT4 #(
		.INIT('h4051)
	) name2612 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		_w937_,
		_w3144_,
		_w3145_
	);
	LUT4 #(
		.INIT('h0080)
	) name2613 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3146_
	);
	LUT3 #(
		.INIT('ha8)
	) name2614 (
		\sa31_reg[2]/P0001 ,
		_w945_,
		_w3146_,
		_w3147_
	);
	LUT4 #(
		.INIT('h0002)
	) name2615 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3148_
	);
	LUT2 #(
		.INIT('h1)
	) name2616 (
		_w939_,
		_w3148_,
		_w3149_
	);
	LUT4 #(
		.INIT('h8000)
	) name2617 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w3150_
	);
	LUT3 #(
		.INIT('h40)
	) name2618 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3151_
	);
	LUT4 #(
		.INIT('h1000)
	) name2619 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3152_
	);
	LUT4 #(
		.INIT('h0007)
	) name2620 (
		_w935_,
		_w967_,
		_w3152_,
		_w3150_,
		_w3153_
	);
	LUT4 #(
		.INIT('h1000)
	) name2621 (
		_w3145_,
		_w3147_,
		_w3149_,
		_w3153_,
		_w3154_
	);
	LUT4 #(
		.INIT('heffb)
	) name2622 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w3155_
	);
	LUT2 #(
		.INIT('h2)
	) name2623 (
		\sa31_reg[7]/P0001 ,
		_w3155_,
		_w3156_
	);
	LUT4 #(
		.INIT('h0777)
	) name2624 (
		\sa31_reg[2]/P0001 ,
		_w1026_,
		_w1001_,
		_w1015_,
		_w3157_
	);
	LUT2 #(
		.INIT('h4)
	) name2625 (
		_w3156_,
		_w3157_,
		_w3158_
	);
	LUT3 #(
		.INIT('h01)
	) name2626 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3159_
	);
	LUT4 #(
		.INIT('h00b1)
	) name2627 (
		\sa31_reg[3]/P0001 ,
		_w1011_,
		_w994_,
		_w3159_,
		_w3160_
	);
	LUT3 #(
		.INIT('h0b)
	) name2628 (
		\sa31_reg[2]/P0001 ,
		_w962_,
		_w976_,
		_w3161_
	);
	LUT4 #(
		.INIT('he400)
	) name2629 (
		\sa31_reg[2]/P0001 ,
		_w956_,
		_w3160_,
		_w3161_,
		_w3162_
	);
	LUT4 #(
		.INIT('hd800)
	) name2630 (
		\sa31_reg[1]/P0001 ,
		_w3154_,
		_w3158_,
		_w3162_,
		_w3163_
	);
	LUT3 #(
		.INIT('h20)
	) name2631 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		_w3164_
	);
	LUT4 #(
		.INIT('h0123)
	) name2632 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3165_
	);
	LUT3 #(
		.INIT('ha8)
	) name2633 (
		\sa31_reg[1]/P0001 ,
		_w3164_,
		_w3165_,
		_w3166_
	);
	LUT3 #(
		.INIT('h04)
	) name2634 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w3167_
	);
	LUT4 #(
		.INIT('h0080)
	) name2635 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3168_
	);
	LUT4 #(
		.INIT('h0020)
	) name2636 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3169_
	);
	LUT3 #(
		.INIT('h01)
	) name2637 (
		_w3167_,
		_w3168_,
		_w3169_,
		_w3170_
	);
	LUT3 #(
		.INIT('h45)
	) name2638 (
		\sa31_reg[2]/P0001 ,
		_w3166_,
		_w3170_,
		_w3171_
	);
	LUT3 #(
		.INIT('h10)
	) name2639 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w3172_
	);
	LUT4 #(
		.INIT('h0008)
	) name2640 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3173_
	);
	LUT3 #(
		.INIT('ha8)
	) name2641 (
		\sa31_reg[2]/P0001 ,
		_w3172_,
		_w3173_,
		_w3174_
	);
	LUT2 #(
		.INIT('h2)
	) name2642 (
		_w967_,
		_w992_,
		_w3175_
	);
	LUT2 #(
		.INIT('h4)
	) name2643 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		_w3176_
	);
	LUT3 #(
		.INIT('h10)
	) name2644 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3177_
	);
	LUT4 #(
		.INIT('h0777)
	) name2645 (
		_w969_,
		_w973_,
		_w3176_,
		_w3177_,
		_w3178_
	);
	LUT4 #(
		.INIT('h5455)
	) name2646 (
		\sa31_reg[1]/P0001 ,
		_w3174_,
		_w3175_,
		_w3178_,
		_w3179_
	);
	LUT2 #(
		.INIT('h8)
	) name2647 (
		\sa31_reg[7]/P0001 ,
		_w970_,
		_w3180_
	);
	LUT4 #(
		.INIT('h13df)
	) name2648 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w948_,
		_w970_,
		_w3181_
	);
	LUT3 #(
		.INIT('h04)
	) name2649 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w3182_
	);
	LUT2 #(
		.INIT('h8)
	) name2650 (
		_w1001_,
		_w3182_,
		_w3183_
	);
	LUT4 #(
		.INIT('h0200)
	) name2651 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3184_
	);
	LUT3 #(
		.INIT('h07)
	) name2652 (
		_w1001_,
		_w3182_,
		_w3184_,
		_w3185_
	);
	LUT3 #(
		.INIT('h2a)
	) name2653 (
		\sa31_reg[1]/P0001 ,
		_w3181_,
		_w3185_,
		_w3186_
	);
	LUT4 #(
		.INIT('h153f)
	) name2654 (
		_w934_,
		_w969_,
		_w973_,
		_w1030_,
		_w3187_
	);
	LUT4 #(
		.INIT('h2000)
	) name2655 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3188_
	);
	LUT4 #(
		.INIT('h23af)
	) name2656 (
		\sa31_reg[2]/P0001 ,
		_w940_,
		_w3188_,
		_w3164_,
		_w3189_
	);
	LUT3 #(
		.INIT('hd0)
	) name2657 (
		\sa31_reg[2]/P0001 ,
		_w3187_,
		_w3189_,
		_w3190_
	);
	LUT4 #(
		.INIT('h0100)
	) name2658 (
		_w3179_,
		_w3186_,
		_w3171_,
		_w3190_,
		_w3191_
	);
	LUT4 #(
		.INIT('hee7f)
	) name2659 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3192_
	);
	LUT4 #(
		.INIT('h5054)
	) name2660 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[5]/P0001 ,
		_w3188_,
		_w3192_,
		_w3193_
	);
	LUT4 #(
		.INIT('h1445)
	) name2661 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3194_
	);
	LUT3 #(
		.INIT('ha2)
	) name2662 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w3195_
	);
	LUT4 #(
		.INIT('h3331)
	) name2663 (
		_w1028_,
		_w1023_,
		_w3195_,
		_w3194_,
		_w3196_
	);
	LUT3 #(
		.INIT('h45)
	) name2664 (
		\sa31_reg[1]/P0001 ,
		_w3193_,
		_w3196_,
		_w3197_
	);
	LUT3 #(
		.INIT('h80)
	) name2665 (
		\sa31_reg[2]/P0001 ,
		_w947_,
		_w985_,
		_w3198_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2666 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w962_,
		_w3148_,
		_w3199_
	);
	LUT3 #(
		.INIT('h8a)
	) name2667 (
		\sa31_reg[1]/P0001 ,
		_w3198_,
		_w3199_,
		_w3200_
	);
	LUT3 #(
		.INIT('h80)
	) name2668 (
		\sa31_reg[4]/P0001 ,
		_w964_,
		_w981_,
		_w3201_
	);
	LUT4 #(
		.INIT('h5540)
	) name2669 (
		\sa31_reg[2]/P0001 ,
		_w947_,
		_w1035_,
		_w3152_,
		_w3202_
	);
	LUT2 #(
		.INIT('h1)
	) name2670 (
		_w3201_,
		_w3202_,
		_w3203_
	);
	LUT3 #(
		.INIT('h10)
	) name2671 (
		_w3197_,
		_w3200_,
		_w3203_,
		_w3204_
	);
	LUT4 #(
		.INIT('he400)
	) name2672 (
		\sa31_reg[0]/P0002 ,
		_w3163_,
		_w3191_,
		_w3204_,
		_w3205_
	);
	LUT3 #(
		.INIT('h69)
	) name2673 (
		\u0_w_reg[2][6]/P0001 ,
		_w745_,
		_w3205_,
		_w3206_
	);
	LUT3 #(
		.INIT('h28)
	) name2674 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[38]/P0001 ,
		\u0_w_reg[2][6]/P0001 ,
		_w3207_
	);
	LUT4 #(
		.INIT('hff41)
	) name2675 (
		\ld_r_reg/P0001 ,
		_w3143_,
		_w3206_,
		_w3207_,
		_w3208_
	);
	LUT4 #(
		.INIT('hbfef)
	) name2676 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3209_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name2677 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3210_
	);
	LUT2 #(
		.INIT('h2)
	) name2678 (
		_w829_,
		_w3210_,
		_w3211_
	);
	LUT3 #(
		.INIT('had)
	) name2679 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w3212_
	);
	LUT4 #(
		.INIT('h0004)
	) name2680 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3213_
	);
	LUT4 #(
		.INIT('hadfb)
	) name2681 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3214_
	);
	LUT4 #(
		.INIT('h0302)
	) name2682 (
		\sa02_reg[3]/P0001 ,
		_w895_,
		_w848_,
		_w3214_,
		_w3215_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2683 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		_w3211_,
		_w3215_,
		_w3216_
	);
	LUT3 #(
		.INIT('ha2)
	) name2684 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w3217_
	);
	LUT4 #(
		.INIT('h4555)
	) name2685 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3218_
	);
	LUT2 #(
		.INIT('h8)
	) name2686 (
		_w3217_,
		_w3218_,
		_w3219_
	);
	LUT3 #(
		.INIT('h8a)
	) name2687 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w3220_
	);
	LUT4 #(
		.INIT('h00d0)
	) name2688 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3221_
	);
	LUT2 #(
		.INIT('h4)
	) name2689 (
		_w3220_,
		_w3221_,
		_w3222_
	);
	LUT3 #(
		.INIT('h02)
	) name2690 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w3223_
	);
	LUT4 #(
		.INIT('h0020)
	) name2691 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w3224_
	);
	LUT3 #(
		.INIT('h07)
	) name2692 (
		_w894_,
		_w3223_,
		_w3224_,
		_w3225_
	);
	LUT4 #(
		.INIT('h5455)
	) name2693 (
		\sa02_reg[1]/P0001 ,
		_w3222_,
		_w3219_,
		_w3225_,
		_w3226_
	);
	LUT3 #(
		.INIT('hf6)
	) name2694 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3227_
	);
	LUT3 #(
		.INIT('h2a)
	) name2695 (
		\sa02_reg[1]/P0001 ,
		_w3212_,
		_w3227_,
		_w3228_
	);
	LUT4 #(
		.INIT('h1000)
	) name2696 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3229_
	);
	LUT3 #(
		.INIT('h01)
	) name2697 (
		_w868_,
		_w873_,
		_w3229_,
		_w3230_
	);
	LUT3 #(
		.INIT('h8a)
	) name2698 (
		\sa02_reg[2]/P0001 ,
		_w3228_,
		_w3230_,
		_w3231_
	);
	LUT4 #(
		.INIT('h0777)
	) name2699 (
		_w822_,
		_w878_,
		_w828_,
		_w3091_,
		_w3232_
	);
	LUT4 #(
		.INIT('hff23)
	) name2700 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3233_
	);
	LUT2 #(
		.INIT('h2)
	) name2701 (
		_w832_,
		_w3233_,
		_w3234_
	);
	LUT3 #(
		.INIT('h2a)
	) name2702 (
		\sa02_reg[0]/P0001 ,
		_w891_,
		_w823_,
		_w3235_
	);
	LUT4 #(
		.INIT('h3100)
	) name2703 (
		\sa02_reg[1]/P0001 ,
		_w3234_,
		_w3232_,
		_w3235_,
		_w3236_
	);
	LUT3 #(
		.INIT('h10)
	) name2704 (
		_w3231_,
		_w3226_,
		_w3236_,
		_w3237_
	);
	LUT4 #(
		.INIT('h77f0)
	) name2705 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3238_
	);
	LUT2 #(
		.INIT('h2)
	) name2706 (
		_w3090_,
		_w3238_,
		_w3239_
	);
	LUT3 #(
		.INIT('h10)
	) name2707 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3240_
	);
	LUT3 #(
		.INIT('h01)
	) name2708 (
		\sa02_reg[1]/P0001 ,
		_w3083_,
		_w3240_,
		_w3241_
	);
	LUT4 #(
		.INIT('h002a)
	) name2709 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		_w898_,
		_w3119_,
		_w3242_
	);
	LUT4 #(
		.INIT('hf5c5)
	) name2710 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3243_
	);
	LUT4 #(
		.INIT('h7707)
	) name2711 (
		\sa02_reg[4]/P0001 ,
		_w883_,
		_w829_,
		_w3243_,
		_w3244_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name2712 (
		_w3239_,
		_w3241_,
		_w3242_,
		_w3244_,
		_w3245_
	);
	LUT4 #(
		.INIT('h5540)
	) name2713 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w852_,
		_w3132_,
		_w3246_
	);
	LUT4 #(
		.INIT('h0008)
	) name2714 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3247_
	);
	LUT4 #(
		.INIT('h8000)
	) name2715 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3248_
	);
	LUT4 #(
		.INIT('h7ff7)
	) name2716 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3249_
	);
	LUT2 #(
		.INIT('h2)
	) name2717 (
		_w891_,
		_w3249_,
		_w3250_
	);
	LUT2 #(
		.INIT('h8)
	) name2718 (
		_w885_,
		_w3123_,
		_w3251_
	);
	LUT3 #(
		.INIT('h8a)
	) name2719 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3252_
	);
	LUT4 #(
		.INIT('h1101)
	) name2720 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3253_
	);
	LUT3 #(
		.INIT('h15)
	) name2721 (
		\sa02_reg[0]/P0001 ,
		_w3252_,
		_w3253_,
		_w3254_
	);
	LUT4 #(
		.INIT('h0100)
	) name2722 (
		_w3246_,
		_w3251_,
		_w3250_,
		_w3254_,
		_w3255_
	);
	LUT2 #(
		.INIT('h4)
	) name2723 (
		_w3245_,
		_w3255_,
		_w3256_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2724 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w825_,
		_w3126_,
		_w3257_
	);
	LUT2 #(
		.INIT('h1)
	) name2725 (
		\sa02_reg[2]/P0001 ,
		_w3257_,
		_w3258_
	);
	LUT4 #(
		.INIT('h0013)
	) name2726 (
		_w822_,
		_w885_,
		_w878_,
		_w3112_,
		_w3259_
	);
	LUT2 #(
		.INIT('h8)
	) name2727 (
		_w884_,
		_w3240_,
		_w3260_
	);
	LUT4 #(
		.INIT('h4000)
	) name2728 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3261_
	);
	LUT3 #(
		.INIT('h07)
	) name2729 (
		_w3252_,
		_w3253_,
		_w3261_,
		_w3262_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2730 (
		\sa02_reg[2]/P0001 ,
		_w3259_,
		_w3260_,
		_w3262_,
		_w3263_
	);
	LUT3 #(
		.INIT('h32)
	) name2731 (
		\sa02_reg[1]/P0001 ,
		_w3258_,
		_w3263_,
		_w3264_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2732 (
		_w3237_,
		_w3256_,
		_w3216_,
		_w3264_,
		_w3265_
	);
	LUT4 #(
		.INIT('hbfef)
	) name2733 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3266_
	);
	LUT2 #(
		.INIT('h4)
	) name2734 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w3267_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name2735 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3268_
	);
	LUT2 #(
		.INIT('h2)
	) name2736 (
		_w558_,
		_w3268_,
		_w3269_
	);
	LUT3 #(
		.INIT('had)
	) name2737 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w3270_
	);
	LUT4 #(
		.INIT('h0004)
	) name2738 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3271_
	);
	LUT4 #(
		.INIT('hadfb)
	) name2739 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3272_
	);
	LUT4 #(
		.INIT('h1302)
	) name2740 (
		\sa13_reg[3]/P0001 ,
		_w534_,
		_w747_,
		_w3272_,
		_w3273_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2741 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[2]/P0001 ,
		_w3269_,
		_w3273_,
		_w3274_
	);
	LUT3 #(
		.INIT('hf6)
	) name2742 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3275_
	);
	LUT3 #(
		.INIT('h2a)
	) name2743 (
		\sa13_reg[2]/P0001 ,
		_w3270_,
		_w3275_,
		_w3276_
	);
	LUT4 #(
		.INIT('h15bf)
	) name2744 (
		\sa13_reg[3]/P0001 ,
		_w537_,
		_w547_,
		_w798_,
		_w3277_
	);
	LUT3 #(
		.INIT('h8a)
	) name2745 (
		\sa13_reg[1]/P0001 ,
		_w3276_,
		_w3277_,
		_w3278_
	);
	LUT4 #(
		.INIT('h7d1d)
	) name2746 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3279_
	);
	LUT2 #(
		.INIT('h1)
	) name2747 (
		\sa13_reg[2]/P0001 ,
		_w3279_,
		_w3280_
	);
	LUT4 #(
		.INIT('h0100)
	) name2748 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w3281_
	);
	LUT2 #(
		.INIT('h8)
	) name2749 (
		\sa13_reg[2]/P0001 ,
		_w3281_,
		_w3282_
	);
	LUT4 #(
		.INIT('h0040)
	) name2750 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3283_
	);
	LUT4 #(
		.INIT('h0020)
	) name2751 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w3284_
	);
	LUT2 #(
		.INIT('h1)
	) name2752 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w3285_
	);
	LUT4 #(
		.INIT('h0010)
	) name2753 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3286_
	);
	LUT3 #(
		.INIT('h01)
	) name2754 (
		_w3283_,
		_w3284_,
		_w3286_,
		_w3287_
	);
	LUT4 #(
		.INIT('h5455)
	) name2755 (
		\sa13_reg[1]/P0001 ,
		_w3280_,
		_w3282_,
		_w3287_,
		_w3288_
	);
	LUT4 #(
		.INIT('h1000)
	) name2756 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3289_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2757 (
		\sa13_reg[2]/P0001 ,
		_w566_,
		_w754_,
		_w3289_,
		_w3290_
	);
	LUT2 #(
		.INIT('h4)
	) name2758 (
		\sa13_reg[2]/P0001 ,
		_w3283_,
		_w3291_
	);
	LUT4 #(
		.INIT('h0040)
	) name2759 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w3292_
	);
	LUT4 #(
		.INIT('h002a)
	) name2760 (
		\sa13_reg[0]/P0001 ,
		_w594_,
		_w779_,
		_w3292_,
		_w3293_
	);
	LUT3 #(
		.INIT('h10)
	) name2761 (
		_w3291_,
		_w3290_,
		_w3293_,
		_w3294_
	);
	LUT3 #(
		.INIT('h10)
	) name2762 (
		_w3288_,
		_w3278_,
		_w3294_,
		_w3295_
	);
	LUT3 #(
		.INIT('h54)
	) name2763 (
		\sa13_reg[2]/P0001 ,
		_w619_,
		_w804_,
		_w3296_
	);
	LUT4 #(
		.INIT('h0800)
	) name2764 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3297_
	);
	LUT3 #(
		.INIT('h0b)
	) name2765 (
		_w589_,
		_w600_,
		_w3297_,
		_w3298_
	);
	LUT3 #(
		.INIT('h8a)
	) name2766 (
		\sa13_reg[1]/P0001 ,
		_w3296_,
		_w3298_,
		_w3299_
	);
	LUT3 #(
		.INIT('h10)
	) name2767 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w3300_
	);
	LUT2 #(
		.INIT('h1)
	) name2768 (
		_w545_,
		_w3300_,
		_w3301_
	);
	LUT3 #(
		.INIT('h20)
	) name2769 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w3302_
	);
	LUT3 #(
		.INIT('h13)
	) name2770 (
		_w594_,
		_w764_,
		_w3302_,
		_w3303_
	);
	LUT3 #(
		.INIT('h15)
	) name2771 (
		\sa13_reg[1]/P0001 ,
		_w3301_,
		_w3303_,
		_w3304_
	);
	LUT4 #(
		.INIT('h3fbb)
	) name2772 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3305_
	);
	LUT2 #(
		.INIT('h2)
	) name2773 (
		_w3285_,
		_w3305_,
		_w3306_
	);
	LUT3 #(
		.INIT('h40)
	) name2774 (
		\sa13_reg[6]/NET0131 ,
		_w584_,
		_w594_,
		_w3307_
	);
	LUT4 #(
		.INIT('h4555)
	) name2775 (
		\sa13_reg[0]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w584_,
		_w594_,
		_w3308_
	);
	LUT4 #(
		.INIT('h0008)
	) name2776 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3309_
	);
	LUT4 #(
		.INIT('h7ff7)
	) name2777 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3310_
	);
	LUT2 #(
		.INIT('h2)
	) name2778 (
		_w594_,
		_w3310_,
		_w3311_
	);
	LUT4 #(
		.INIT('h5540)
	) name2779 (
		\sa13_reg[2]/P0001 ,
		_w535_,
		_w591_,
		_w615_,
		_w3312_
	);
	LUT4 #(
		.INIT('h0100)
	) name2780 (
		_w3311_,
		_w3306_,
		_w3312_,
		_w3308_,
		_w3313_
	);
	LUT3 #(
		.INIT('h10)
	) name2781 (
		_w3304_,
		_w3299_,
		_w3313_,
		_w3314_
	);
	LUT4 #(
		.INIT('h23af)
	) name2782 (
		\sa13_reg[4]/P0001 ,
		_w556_,
		_w748_,
		_w804_,
		_w3315_
	);
	LUT2 #(
		.INIT('h1)
	) name2783 (
		\sa13_reg[2]/P0001 ,
		_w3315_,
		_w3316_
	);
	LUT3 #(
		.INIT('h80)
	) name2784 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w3317_
	);
	LUT4 #(
		.INIT('h4000)
	) name2785 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w3318_
	);
	LUT4 #(
		.INIT('h0013)
	) name2786 (
		\sa13_reg[3]/P0001 ,
		_w750_,
		_w798_,
		_w3318_,
		_w3319_
	);
	LUT4 #(
		.INIT('h4000)
	) name2787 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w3320_
	);
	LUT3 #(
		.INIT('h07)
	) name2788 (
		_w578_,
		_w3300_,
		_w3320_,
		_w3321_
	);
	LUT4 #(
		.INIT('h3100)
	) name2789 (
		\sa13_reg[2]/P0001 ,
		_w3306_,
		_w3319_,
		_w3321_,
		_w3322_
	);
	LUT3 #(
		.INIT('h32)
	) name2790 (
		\sa13_reg[1]/P0001 ,
		_w3316_,
		_w3322_,
		_w3323_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2791 (
		_w3295_,
		_w3314_,
		_w3274_,
		_w3323_,
		_w3324_
	);
	LUT3 #(
		.INIT('h69)
	) name2792 (
		_w3142_,
		_w3265_,
		_w3324_,
		_w3325_
	);
	LUT4 #(
		.INIT('h0010)
	) name2793 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3326_
	);
	LUT4 #(
		.INIT('hbfef)
	) name2794 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3327_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name2795 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3328_
	);
	LUT2 #(
		.INIT('h2)
	) name2796 (
		_w686_,
		_w3328_,
		_w3329_
	);
	LUT3 #(
		.INIT('had)
	) name2797 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w3330_
	);
	LUT4 #(
		.INIT('h0004)
	) name2798 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3331_
	);
	LUT4 #(
		.INIT('hadfb)
	) name2799 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3332_
	);
	LUT4 #(
		.INIT('h0302)
	) name2800 (
		\sa20_reg[3]/P0001 ,
		_w661_,
		_w701_,
		_w3332_,
		_w3333_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2801 (
		\sa20_reg[1]/P0001 ,
		\sa20_reg[2]/P0001 ,
		_w3329_,
		_w3333_,
		_w3334_
	);
	LUT3 #(
		.INIT('hf6)
	) name2802 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3335_
	);
	LUT3 #(
		.INIT('h2a)
	) name2803 (
		\sa20_reg[1]/P0001 ,
		_w3330_,
		_w3335_,
		_w3336_
	);
	LUT4 #(
		.INIT('h0080)
	) name2804 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3337_
	);
	LUT4 #(
		.INIT('h1000)
	) name2805 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3338_
	);
	LUT3 #(
		.INIT('h01)
	) name2806 (
		_w672_,
		_w3338_,
		_w3337_,
		_w3339_
	);
	LUT3 #(
		.INIT('h8a)
	) name2807 (
		\sa20_reg[2]/P0001 ,
		_w3336_,
		_w3339_,
		_w3340_
	);
	LUT4 #(
		.INIT('h0100)
	) name2808 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w3341_
	);
	LUT3 #(
		.INIT('h7d)
	) name2809 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w3342_
	);
	LUT4 #(
		.INIT('he4f5)
	) name2810 (
		\sa20_reg[2]/P0001 ,
		_w641_,
		_w3341_,
		_w3342_,
		_w3343_
	);
	LUT2 #(
		.INIT('h2)
	) name2811 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w3344_
	);
	LUT3 #(
		.INIT('h04)
	) name2812 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3345_
	);
	LUT2 #(
		.INIT('h4)
	) name2813 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w3346_
	);
	LUT4 #(
		.INIT('h0040)
	) name2814 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3347_
	);
	LUT4 #(
		.INIT('h0020)
	) name2815 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w3348_
	);
	LUT4 #(
		.INIT('h1011)
	) name2816 (
		_w3347_,
		_w3348_,
		_w3344_,
		_w3345_,
		_w3349_
	);
	LUT3 #(
		.INIT('h45)
	) name2817 (
		\sa20_reg[1]/P0001 ,
		_w3343_,
		_w3349_,
		_w3350_
	);
	LUT3 #(
		.INIT('h10)
	) name2818 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3351_
	);
	LUT4 #(
		.INIT('h135f)
	) name2819 (
		\sa20_reg[4]/P0001 ,
		_w654_,
		_w708_,
		_w3351_,
		_w3352_
	);
	LUT2 #(
		.INIT('h8)
	) name2820 (
		_w641_,
		_w654_,
		_w3353_
	);
	LUT4 #(
		.INIT('h0200)
	) name2821 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w3354_
	);
	LUT4 #(
		.INIT('h0040)
	) name2822 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w3355_
	);
	LUT3 #(
		.INIT('h07)
	) name2823 (
		\sa20_reg[3]/P0001 ,
		_w3354_,
		_w3355_,
		_w3356_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2824 (
		\sa20_reg[1]/P0001 ,
		_w3352_,
		_w3353_,
		_w3356_,
		_w3357_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2825 (
		\sa20_reg[0]/P0001 ,
		_w3350_,
		_w3340_,
		_w3357_,
		_w3358_
	);
	LUT4 #(
		.INIT('hf2fa)
	) name2826 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		_w3359_
	);
	LUT2 #(
		.INIT('h2)
	) name2827 (
		\sa20_reg[7]/NET0131 ,
		_w3359_,
		_w3360_
	);
	LUT3 #(
		.INIT('h20)
	) name2828 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w3361_
	);
	LUT4 #(
		.INIT('h0002)
	) name2829 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3362_
	);
	LUT4 #(
		.INIT('h0105)
	) name2830 (
		\sa20_reg[1]/P0001 ,
		_w692_,
		_w3362_,
		_w3361_,
		_w3363_
	);
	LUT4 #(
		.INIT('h0020)
	) name2831 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3364_
	);
	LUT3 #(
		.INIT('h54)
	) name2832 (
		\sa20_reg[2]/P0001 ,
		_w648_,
		_w3364_,
		_w3365_
	);
	LUT3 #(
		.INIT('hcd)
	) name2833 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w3366_
	);
	LUT4 #(
		.INIT('h0a02)
	) name2834 (
		\sa20_reg[1]/P0001 ,
		_w693_,
		_w720_,
		_w3366_,
		_w3367_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2835 (
		_w3360_,
		_w3363_,
		_w3365_,
		_w3367_,
		_w3368_
	);
	LUT4 #(
		.INIT('h4000)
	) name2836 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3369_
	);
	LUT4 #(
		.INIT('h0010)
	) name2837 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w3370_
	);
	LUT2 #(
		.INIT('h1)
	) name2838 (
		_w3369_,
		_w3370_,
		_w3371_
	);
	LUT3 #(
		.INIT('h07)
	) name2839 (
		\sa20_reg[4]/P0001 ,
		_w701_,
		_w730_,
		_w3372_
	);
	LUT4 #(
		.INIT('h0008)
	) name2840 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3373_
	);
	LUT4 #(
		.INIT('h8000)
	) name2841 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3374_
	);
	LUT4 #(
		.INIT('h7ff6)
	) name2842 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3375_
	);
	LUT2 #(
		.INIT('h2)
	) name2843 (
		_w692_,
		_w3375_,
		_w3376_
	);
	LUT4 #(
		.INIT('h00ea)
	) name2844 (
		\sa20_reg[2]/P0001 ,
		_w3371_,
		_w3372_,
		_w3376_,
		_w3377_
	);
	LUT3 #(
		.INIT('h45)
	) name2845 (
		\sa20_reg[0]/P0001 ,
		_w3368_,
		_w3377_,
		_w3378_
	);
	LUT4 #(
		.INIT('h23af)
	) name2846 (
		\sa20_reg[6]/NET0131 ,
		_w642_,
		_w660_,
		_w3345_,
		_w3379_
	);
	LUT2 #(
		.INIT('h1)
	) name2847 (
		\sa20_reg[2]/P0001 ,
		_w3379_,
		_w3380_
	);
	LUT4 #(
		.INIT('h4000)
	) name2848 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w3381_
	);
	LUT3 #(
		.INIT('h2a)
	) name2849 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w708_,
		_w3382_
	);
	LUT3 #(
		.INIT('h02)
	) name2850 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w3383_
	);
	LUT4 #(
		.INIT('h0002)
	) name2851 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3384_
	);
	LUT2 #(
		.INIT('h1)
	) name2852 (
		_w678_,
		_w3384_,
		_w3385_
	);
	LUT4 #(
		.INIT('h0001)
	) name2853 (
		\sa20_reg[2]/P0001 ,
		_w688_,
		_w3369_,
		_w3370_,
		_w3386_
	);
	LUT4 #(
		.INIT('h5540)
	) name2854 (
		_w3381_,
		_w3382_,
		_w3385_,
		_w3386_,
		_w3387_
	);
	LUT3 #(
		.INIT('h32)
	) name2855 (
		\sa20_reg[1]/P0001 ,
		_w3380_,
		_w3387_,
		_w3388_
	);
	LUT4 #(
		.INIT('h0100)
	) name2856 (
		_w3358_,
		_w3334_,
		_w3378_,
		_w3388_,
		_w3389_
	);
	LUT3 #(
		.INIT('h69)
	) name2857 (
		\u0_w_reg[2][7]/P0001 ,
		_w1039_,
		_w3389_,
		_w3390_
	);
	LUT3 #(
		.INIT('h82)
	) name2858 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[39]/P0001 ,
		\u0_w_reg[2][7]/P0001 ,
		_w3391_
	);
	LUT4 #(
		.INIT('h00eb)
	) name2859 (
		\ld_r_reg/P0001 ,
		_w3325_,
		_w3390_,
		_w3391_,
		_w3392_
	);
	LUT4 #(
		.INIT('h1555)
	) name2860 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w3393_
	);
	LUT3 #(
		.INIT('h70)
	) name2861 (
		\sa13_reg[2]/P0001 ,
		_w563_,
		_w3393_,
		_w3394_
	);
	LUT3 #(
		.INIT('h80)
	) name2862 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3395_
	);
	LUT4 #(
		.INIT('h2000)
	) name2863 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3396_
	);
	LUT4 #(
		.INIT('h1000)
	) name2864 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w3397_
	);
	LUT4 #(
		.INIT('h0007)
	) name2865 (
		_w589_,
		_w804_,
		_w3397_,
		_w3396_,
		_w3398_
	);
	LUT2 #(
		.INIT('h8)
	) name2866 (
		_w3394_,
		_w3398_,
		_w3399_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name2867 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3400_
	);
	LUT2 #(
		.INIT('h1)
	) name2868 (
		\sa13_reg[2]/P0001 ,
		_w3400_,
		_w3401_
	);
	LUT3 #(
		.INIT('h2a)
	) name2869 (
		\sa13_reg[1]/P0001 ,
		_w543_,
		_w613_,
		_w3402_
	);
	LUT4 #(
		.INIT('h0200)
	) name2870 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3403_
	);
	LUT3 #(
		.INIT('h0b)
	) name2871 (
		\sa13_reg[3]/P0001 ,
		_w615_,
		_w3403_,
		_w3404_
	);
	LUT3 #(
		.INIT('h20)
	) name2872 (
		_w3402_,
		_w3401_,
		_w3404_,
		_w3405_
	);
	LUT4 #(
		.INIT('hd5dd)
	) name2873 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w3406_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2874 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w3407_
	);
	LUT4 #(
		.INIT('h3200)
	) name2875 (
		\sa13_reg[6]/NET0131 ,
		_w765_,
		_w3406_,
		_w3407_,
		_w3408_
	);
	LUT4 #(
		.INIT('h2000)
	) name2876 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3409_
	);
	LUT4 #(
		.INIT('h0045)
	) name2877 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[5]/P0001 ,
		_w617_,
		_w3409_,
		_w3410_
	);
	LUT3 #(
		.INIT('h23)
	) name2878 (
		_w790_,
		_w3408_,
		_w3410_,
		_w3411_
	);
	LUT4 #(
		.INIT('haa02)
	) name2879 (
		\sa13_reg[0]/P0001 ,
		_w3399_,
		_w3405_,
		_w3411_,
		_w3412_
	);
	LUT4 #(
		.INIT('h0100)
	) name2880 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3413_
	);
	LUT4 #(
		.INIT('h5504)
	) name2881 (
		\sa13_reg[2]/P0001 ,
		_w538_,
		_w613_,
		_w3413_,
		_w3414_
	);
	LUT4 #(
		.INIT('h0080)
	) name2882 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3415_
	);
	LUT4 #(
		.INIT('h0015)
	) name2883 (
		_w574_,
		_w583_,
		_w3302_,
		_w3415_,
		_w3416_
	);
	LUT3 #(
		.INIT('h8a)
	) name2884 (
		\sa13_reg[1]/P0001 ,
		_w3414_,
		_w3416_,
		_w3417_
	);
	LUT4 #(
		.INIT('h8000)
	) name2885 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w3418_
	);
	LUT2 #(
		.INIT('h1)
	) name2886 (
		_w764_,
		_w3418_,
		_w3419_
	);
	LUT4 #(
		.INIT('h0002)
	) name2887 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3420_
	);
	LUT3 #(
		.INIT('h07)
	) name2888 (
		_w747_,
		_w3285_,
		_w3420_,
		_w3421_
	);
	LUT3 #(
		.INIT('h15)
	) name2889 (
		\sa13_reg[1]/P0001 ,
		_w3419_,
		_w3421_,
		_w3422_
	);
	LUT4 #(
		.INIT('h3310)
	) name2890 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w798_,
		_w3271_,
		_w3423_
	);
	LUT4 #(
		.INIT('h0100)
	) name2891 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w3424_
	);
	LUT4 #(
		.INIT('haa80)
	) name2892 (
		\sa13_reg[2]/P0001 ,
		_w556_,
		_w804_,
		_w3424_,
		_w3425_
	);
	LUT2 #(
		.INIT('h1)
	) name2893 (
		_w3423_,
		_w3425_,
		_w3426_
	);
	LUT4 #(
		.INIT('h5455)
	) name2894 (
		\sa13_reg[0]/P0001 ,
		_w3422_,
		_w3417_,
		_w3426_,
		_w3427_
	);
	LUT4 #(
		.INIT('h0084)
	) name2895 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3428_
	);
	LUT2 #(
		.INIT('h8)
	) name2896 (
		_w576_,
		_w553_,
		_w3429_
	);
	LUT4 #(
		.INIT('h080a)
	) name2897 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w3284_,
		_w3413_,
		_w3430_
	);
	LUT3 #(
		.INIT('h10)
	) name2898 (
		_w3428_,
		_w3429_,
		_w3430_,
		_w3431_
	);
	LUT2 #(
		.INIT('h8)
	) name2899 (
		\sa13_reg[5]/P0001 ,
		_w3396_,
		_w3432_
	);
	LUT3 #(
		.INIT('h01)
	) name2900 (
		\sa13_reg[2]/P0001 ,
		_w600_,
		_w751_,
		_w3433_
	);
	LUT2 #(
		.INIT('h4)
	) name2901 (
		_w3432_,
		_w3433_,
		_w3434_
	);
	LUT4 #(
		.INIT('h135f)
	) name2902 (
		_w535_,
		_w543_,
		_w591_,
		_w616_,
		_w3435_
	);
	LUT4 #(
		.INIT('h0155)
	) name2903 (
		\sa13_reg[1]/P0001 ,
		_w3431_,
		_w3434_,
		_w3435_,
		_w3436_
	);
	LUT4 #(
		.INIT('hc840)
	) name2904 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w795_,
		_w3317_,
		_w3437_
	);
	LUT2 #(
		.INIT('h8)
	) name2905 (
		\sa13_reg[7]/NET0131 ,
		_w625_,
		_w3438_
	);
	LUT3 #(
		.INIT('h23)
	) name2906 (
		\sa13_reg[5]/P0001 ,
		_w605_,
		_w617_,
		_w3439_
	);
	LUT3 #(
		.INIT('h45)
	) name2907 (
		\sa13_reg[2]/P0001 ,
		_w3438_,
		_w3439_,
		_w3440_
	);
	LUT4 #(
		.INIT('h337f)
	) name2908 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w543_,
		_w798_,
		_w3441_
	);
	LUT4 #(
		.INIT('h0777)
	) name2909 (
		_w536_,
		_w583_,
		_w814_,
		_w3267_,
		_w3442_
	);
	LUT2 #(
		.INIT('h8)
	) name2910 (
		_w3441_,
		_w3442_,
		_w3443_
	);
	LUT4 #(
		.INIT('h1311)
	) name2911 (
		\sa13_reg[1]/P0001 ,
		_w3437_,
		_w3440_,
		_w3443_,
		_w3444_
	);
	LUT4 #(
		.INIT('h0100)
	) name2912 (
		_w3412_,
		_w3436_,
		_w3427_,
		_w3444_,
		_w3445_
	);
	LUT4 #(
		.INIT('h0100)
	) name2913 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3446_
	);
	LUT4 #(
		.INIT('h5504)
	) name2914 (
		\sa02_reg[2]/P0001 ,
		_w880_,
		_w837_,
		_w3446_,
		_w3447_
	);
	LUT3 #(
		.INIT('h20)
	) name2915 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3448_
	);
	LUT3 #(
		.INIT('h08)
	) name2916 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3449_
	);
	LUT4 #(
		.INIT('h0080)
	) name2917 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3450_
	);
	LUT4 #(
		.INIT('h0103)
	) name2918 (
		_w833_,
		_w911_,
		_w3450_,
		_w3448_,
		_w3451_
	);
	LUT3 #(
		.INIT('h8a)
	) name2919 (
		\sa02_reg[1]/P0001 ,
		_w3447_,
		_w3451_,
		_w3452_
	);
	LUT4 #(
		.INIT('h0040)
	) name2920 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3453_
	);
	LUT4 #(
		.INIT('h5150)
	) name2921 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		_w929_,
		_w3453_,
		_w3454_
	);
	LUT4 #(
		.INIT('h3310)
	) name2922 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		_w864_,
		_w3213_,
		_w3455_
	);
	LUT4 #(
		.INIT('haa20)
	) name2923 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		_w825_,
		_w3076_,
		_w3456_
	);
	LUT4 #(
		.INIT('h7f7c)
	) name2924 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3457_
	);
	LUT2 #(
		.INIT('h2)
	) name2925 (
		_w3086_,
		_w3457_,
		_w3458_
	);
	LUT4 #(
		.INIT('h0001)
	) name2926 (
		_w3454_,
		_w3456_,
		_w3458_,
		_w3455_,
		_w3459_
	);
	LUT3 #(
		.INIT('h45)
	) name2927 (
		\sa02_reg[0]/P0001 ,
		_w3452_,
		_w3459_,
		_w3460_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name2928 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3461_
	);
	LUT2 #(
		.INIT('h1)
	) name2929 (
		\sa02_reg[2]/P0001 ,
		_w3461_,
		_w3462_
	);
	LUT4 #(
		.INIT('h0200)
	) name2930 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3463_
	);
	LUT4 #(
		.INIT('h008a)
	) name2931 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w855_,
		_w3463_,
		_w3464_
	);
	LUT3 #(
		.INIT('h10)
	) name2932 (
		_w924_,
		_w3462_,
		_w3464_,
		_w3465_
	);
	LUT4 #(
		.INIT('h2000)
	) name2933 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3466_
	);
	LUT4 #(
		.INIT('h0015)
	) name2934 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		_w904_,
		_w3466_,
		_w3467_
	);
	LUT2 #(
		.INIT('h1)
	) name2935 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w3468_
	);
	LUT3 #(
		.INIT('h32)
	) name2936 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w3469_
	);
	LUT4 #(
		.INIT('haf23)
	) name2937 (
		\sa02_reg[2]/P0001 ,
		_w874_,
		_w825_,
		_w3469_,
		_w3470_
	);
	LUT2 #(
		.INIT('h8)
	) name2938 (
		_w3467_,
		_w3470_,
		_w3471_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2939 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w3472_
	);
	LUT4 #(
		.INIT('h0200)
	) name2940 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3473_
	);
	LUT3 #(
		.INIT('h04)
	) name2941 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3474_
	);
	LUT4 #(
		.INIT('h0100)
	) name2942 (
		_w3121_,
		_w3474_,
		_w3473_,
		_w3472_,
		_w3475_
	);
	LUT4 #(
		.INIT('h2000)
	) name2943 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3476_
	);
	LUT3 #(
		.INIT('h01)
	) name2944 (
		\sa02_reg[2]/P0001 ,
		_w846_,
		_w3476_,
		_w3477_
	);
	LUT3 #(
		.INIT('h23)
	) name2945 (
		_w3135_,
		_w3475_,
		_w3477_,
		_w3478_
	);
	LUT4 #(
		.INIT('haa02)
	) name2946 (
		\sa02_reg[0]/P0001 ,
		_w3465_,
		_w3471_,
		_w3478_,
		_w3479_
	);
	LUT3 #(
		.INIT('h07)
	) name2947 (
		_w870_,
		_w831_,
		_w3109_,
		_w3480_
	);
	LUT3 #(
		.INIT('h45)
	) name2948 (
		\sa02_reg[2]/P0001 ,
		_w3135_,
		_w3480_,
		_w3481_
	);
	LUT4 #(
		.INIT('h135f)
	) name2949 (
		\sa02_reg[4]/P0001 ,
		_w905_,
		_w927_,
		_w3106_,
		_w3482_
	);
	LUT4 #(
		.INIT('h0777)
	) name2950 (
		_w822_,
		_w878_,
		_w837_,
		_w828_,
		_w3483_
	);
	LUT2 #(
		.INIT('h8)
	) name2951 (
		_w3482_,
		_w3483_,
		_w3484_
	);
	LUT3 #(
		.INIT('h8a)
	) name2952 (
		\sa02_reg[1]/P0001 ,
		_w3481_,
		_w3484_,
		_w3485_
	);
	LUT4 #(
		.INIT('h0084)
	) name2953 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3486_
	);
	LUT2 #(
		.INIT('h9)
	) name2954 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w3487_
	);
	LUT4 #(
		.INIT('h020a)
	) name2955 (
		\sa02_reg[2]/P0001 ,
		_w828_,
		_w3224_,
		_w3487_,
		_w3488_
	);
	LUT3 #(
		.INIT('h13)
	) name2956 (
		_w861_,
		_w898_,
		_w875_,
		_w3489_
	);
	LUT4 #(
		.INIT('h45cf)
	) name2957 (
		_w922_,
		_w3486_,
		_w3488_,
		_w3489_,
		_w3490_
	);
	LUT4 #(
		.INIT('h0010)
	) name2958 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3491_
	);
	LUT3 #(
		.INIT('h27)
	) name2959 (
		\sa02_reg[6]/NET0131 ,
		_w852_,
		_w3491_,
		_w3492_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2960 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w3493_
	);
	LUT4 #(
		.INIT('h00c8)
	) name2961 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		_w862_,
		_w3493_,
		_w3494_
	);
	LUT4 #(
		.INIT('h00ba)
	) name2962 (
		\sa02_reg[1]/P0001 ,
		_w3490_,
		_w3492_,
		_w3494_,
		_w3495_
	);
	LUT4 #(
		.INIT('h0100)
	) name2963 (
		_w3460_,
		_w3479_,
		_w3485_,
		_w3495_,
		_w3496_
	);
	LUT2 #(
		.INIT('h9)
	) name2964 (
		_w3445_,
		_w3496_,
		_w3497_
	);
	LUT4 #(
		.INIT('h0010)
	) name2965 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3498_
	);
	LUT3 #(
		.INIT('h01)
	) name2966 (
		\sa20_reg[2]/P0001 ,
		_w672_,
		_w3498_,
		_w3499_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2967 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w3500_
	);
	LUT2 #(
		.INIT('h4)
	) name2968 (
		_w3337_,
		_w3500_,
		_w3501_
	);
	LUT2 #(
		.INIT('h1)
	) name2969 (
		_w3499_,
		_w3501_,
		_w3502_
	);
	LUT4 #(
		.INIT('h0400)
	) name2970 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3503_
	);
	LUT4 #(
		.INIT('h8000)
	) name2971 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w3504_
	);
	LUT3 #(
		.INIT('h01)
	) name2972 (
		_w644_,
		_w3504_,
		_w3503_,
		_w3505_
	);
	LUT4 #(
		.INIT('h020a)
	) name2973 (
		\sa20_reg[1]/P0001 ,
		_w642_,
		_w640_,
		_w3345_,
		_w3506_
	);
	LUT3 #(
		.INIT('h40)
	) name2974 (
		_w3384_,
		_w3505_,
		_w3506_,
		_w3507_
	);
	LUT3 #(
		.INIT('h15)
	) name2975 (
		\sa20_reg[1]/P0001 ,
		_w735_,
		_w736_,
		_w3508_
	);
	LUT2 #(
		.INIT('h8)
	) name2976 (
		_w3344_,
		_w3383_,
		_w3509_
	);
	LUT3 #(
		.INIT('h80)
	) name2977 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3510_
	);
	LUT2 #(
		.INIT('h8)
	) name2978 (
		_w710_,
		_w3510_,
		_w3511_
	);
	LUT4 #(
		.INIT('h0777)
	) name2979 (
		_w639_,
		_w704_,
		_w710_,
		_w3510_,
		_w3512_
	);
	LUT3 #(
		.INIT('h40)
	) name2980 (
		_w3509_,
		_w3508_,
		_w3512_,
		_w3513_
	);
	LUT4 #(
		.INIT('h0001)
	) name2981 (
		\sa20_reg[2]/P0001 ,
		_w666_,
		_w660_,
		_w661_,
		_w3514_
	);
	LUT3 #(
		.INIT('h2a)
	) name2982 (
		\sa20_reg[2]/P0001 ,
		_w671_,
		_w667_,
		_w3515_
	);
	LUT3 #(
		.INIT('hd0)
	) name2983 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w3516_
	);
	LUT3 #(
		.INIT('h0d)
	) name2984 (
		_w681_,
		_w3516_,
		_w3504_,
		_w3517_
	);
	LUT2 #(
		.INIT('h1)
	) name2985 (
		\sa20_reg[0]/P0001 ,
		_w682_,
		_w3518_
	);
	LUT4 #(
		.INIT('hea00)
	) name2986 (
		_w3514_,
		_w3515_,
		_w3517_,
		_w3518_,
		_w3519_
	);
	LUT4 #(
		.INIT('hf400)
	) name2987 (
		_w3502_,
		_w3507_,
		_w3513_,
		_w3519_,
		_w3520_
	);
	LUT3 #(
		.INIT('h10)
	) name2988 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w3521_
	);
	LUT4 #(
		.INIT('h0008)
	) name2989 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3522_
	);
	LUT3 #(
		.INIT('ha8)
	) name2990 (
		\sa20_reg[2]/P0001 ,
		_w3521_,
		_w3522_,
		_w3523_
	);
	LUT3 #(
		.INIT('h01)
	) name2991 (
		\sa20_reg[1]/P0001 ,
		_w701_,
		_w3347_,
		_w3524_
	);
	LUT4 #(
		.INIT('h0777)
	) name2992 (
		\sa20_reg[7]/NET0131 ,
		_w678_,
		_w686_,
		_w3351_,
		_w3525_
	);
	LUT3 #(
		.INIT('h40)
	) name2993 (
		_w3523_,
		_w3524_,
		_w3525_,
		_w3526_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2994 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w666_,
		_w649_,
		_w3527_
	);
	LUT2 #(
		.INIT('h8)
	) name2995 (
		_w671_,
		_w736_,
		_w3528_
	);
	LUT4 #(
		.INIT('h0200)
	) name2996 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3529_
	);
	LUT4 #(
		.INIT('h002a)
	) name2997 (
		\sa20_reg[1]/P0001 ,
		_w671_,
		_w736_,
		_w3529_,
		_w3530_
	);
	LUT2 #(
		.INIT('h8)
	) name2998 (
		_w3527_,
		_w3530_,
		_w3531_
	);
	LUT4 #(
		.INIT('h0123)
	) name2999 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3532_
	);
	LUT3 #(
		.INIT('ha8)
	) name3000 (
		\sa20_reg[1]/P0001 ,
		_w728_,
		_w3532_,
		_w3533_
	);
	LUT4 #(
		.INIT('h0020)
	) name3001 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3534_
	);
	LUT4 #(
		.INIT('h5545)
	) name3002 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w3535_
	);
	LUT3 #(
		.INIT('h10)
	) name3003 (
		_w701_,
		_w3534_,
		_w3535_,
		_w3536_
	);
	LUT2 #(
		.INIT('h8)
	) name3004 (
		_w667_,
		_w710_,
		_w3537_
	);
	LUT3 #(
		.INIT('h2a)
	) name3005 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w678_,
		_w3538_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3006 (
		_w3533_,
		_w3536_,
		_w3537_,
		_w3538_,
		_w3539_
	);
	LUT2 #(
		.INIT('h8)
	) name3007 (
		_w642_,
		_w675_,
		_w3540_
	);
	LUT3 #(
		.INIT('h2a)
	) name3008 (
		\sa20_reg[0]/P0001 ,
		_w3346_,
		_w3361_,
		_w3541_
	);
	LUT2 #(
		.INIT('h4)
	) name3009 (
		_w3540_,
		_w3541_,
		_w3542_
	);
	LUT4 #(
		.INIT('h5400)
	) name3010 (
		_w3539_,
		_w3526_,
		_w3531_,
		_w3542_,
		_w3543_
	);
	LUT4 #(
		.INIT('hd850)
	) name3011 (
		\sa20_reg[2]/P0001 ,
		_w677_,
		_w666_,
		_w707_,
		_w3544_
	);
	LUT3 #(
		.INIT('h2a)
	) name3012 (
		\sa20_reg[1]/P0001 ,
		\sa20_reg[3]/P0001 ,
		_w682_,
		_w3545_
	);
	LUT3 #(
		.INIT('h6b)
	) name3013 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3546_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3014 (
		\sa20_reg[2]/P0001 ,
		_w671_,
		_w649_,
		_w3546_,
		_w3547_
	);
	LUT2 #(
		.INIT('h1)
	) name3015 (
		\sa20_reg[1]/P0001 ,
		_w731_,
		_w3548_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3016 (
		_w3544_,
		_w3545_,
		_w3547_,
		_w3548_,
		_w3549_
	);
	LUT4 #(
		.INIT('h2000)
	) name3017 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3550_
	);
	LUT4 #(
		.INIT('h1000)
	) name3018 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w3551_
	);
	LUT4 #(
		.INIT('h0007)
	) name3019 (
		\sa20_reg[4]/P0001 ,
		_w701_,
		_w3550_,
		_w3551_,
		_w3552_
	);
	LUT3 #(
		.INIT('h15)
	) name3020 (
		_w640_,
		_w700_,
		_w740_,
		_w3553_
	);
	LUT4 #(
		.INIT('h0133)
	) name3021 (
		\sa20_reg[1]/P0001 ,
		\sa20_reg[2]/P0001 ,
		_w3552_,
		_w3553_,
		_w3554_
	);
	LUT2 #(
		.INIT('h8)
	) name3022 (
		_w692_,
		_w3373_,
		_w3555_
	);
	LUT3 #(
		.INIT('h01)
	) name3023 (
		_w3554_,
		_w3549_,
		_w3555_,
		_w3556_
	);
	LUT3 #(
		.INIT('he0)
	) name3024 (
		_w3520_,
		_w3543_,
		_w3556_,
		_w3557_
	);
	LUT3 #(
		.INIT('h4b)
	) name3025 (
		_w775_,
		_w821_,
		_w3557_,
		_w3558_
	);
	LUT2 #(
		.INIT('h9)
	) name3026 (
		\u0_w_reg[2][29]/P0001 ,
		_w3205_,
		_w3559_
	);
	LUT4 #(
		.INIT('h1441)
	) name3027 (
		\ld_r_reg/P0001 ,
		_w3497_,
		_w3558_,
		_w3559_,
		_w3560_
	);
	LUT3 #(
		.INIT('h82)
	) name3028 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[61]/P0001 ,
		\u0_w_reg[2][29]/P0001 ,
		_w3561_
	);
	LUT2 #(
		.INIT('h1)
	) name3029 (
		_w3560_,
		_w3561_,
		_w3562_
	);
	LUT4 #(
		.INIT('hb44b)
	) name3030 (
		_w775_,
		_w821_,
		_w3142_,
		_w3557_,
		_w3563_
	);
	LUT4 #(
		.INIT('h5655)
	) name3031 (
		\u0_w_reg[2][22]/P0001 ,
		_w980_,
		_w1009_,
		_w1038_,
		_w3564_
	);
	LUT2 #(
		.INIT('h6)
	) name3032 (
		_w745_,
		_w3564_,
		_w3565_
	);
	LUT3 #(
		.INIT('h82)
	) name3033 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[54]/P0001 ,
		\u0_w_reg[2][22]/P0001 ,
		_w3566_
	);
	LUT4 #(
		.INIT('h00eb)
	) name3034 (
		\ld_r_reg/P0001 ,
		_w3563_,
		_w3565_,
		_w3566_,
		_w3567_
	);
	LUT3 #(
		.INIT('h20)
	) name3035 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3568_
	);
	LUT4 #(
		.INIT('h0100)
	) name3036 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3569_
	);
	LUT4 #(
		.INIT('h5510)
	) name3037 (
		\sa20_reg[2]/P0001 ,
		_w652_,
		_w3568_,
		_w3569_,
		_w3570_
	);
	LUT4 #(
		.INIT('h0080)
	) name3038 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3571_
	);
	LUT4 #(
		.INIT('h0015)
	) name3039 (
		_w676_,
		_w735_,
		_w3361_,
		_w3571_,
		_w3572_
	);
	LUT3 #(
		.INIT('h8a)
	) name3040 (
		\sa20_reg[1]/P0001 ,
		_w3570_,
		_w3572_,
		_w3573_
	);
	LUT4 #(
		.INIT('h0040)
	) name3041 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3574_
	);
	LUT2 #(
		.INIT('h4)
	) name3042 (
		\sa20_reg[2]/P0001 ,
		_w3574_,
		_w3575_
	);
	LUT4 #(
		.INIT('h8000)
	) name3043 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w3576_
	);
	LUT3 #(
		.INIT('h01)
	) name3044 (
		_w718_,
		_w3362_,
		_w3576_,
		_w3577_
	);
	LUT3 #(
		.INIT('h45)
	) name3045 (
		\sa20_reg[1]/P0001 ,
		_w3575_,
		_w3577_,
		_w3578_
	);
	LUT4 #(
		.INIT('h5450)
	) name3046 (
		\sa20_reg[3]/P0001 ,
		_w3346_,
		_w3354_,
		_w3361_,
		_w3579_
	);
	LUT2 #(
		.INIT('h8)
	) name3047 (
		_w662_,
		_w710_,
		_w3580_
	);
	LUT4 #(
		.INIT('h67ef)
	) name3048 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w662_,
		_w3362_,
		_w3581_
	);
	LUT2 #(
		.INIT('h4)
	) name3049 (
		_w3579_,
		_w3581_,
		_w3582_
	);
	LUT4 #(
		.INIT('h5455)
	) name3050 (
		\sa20_reg[0]/P0001 ,
		_w3578_,
		_w3573_,
		_w3582_,
		_w3583_
	);
	LUT3 #(
		.INIT('h02)
	) name3051 (
		\sa20_reg[2]/P0001 ,
		_w701_,
		_w3348_,
		_w3584_
	);
	LUT2 #(
		.INIT('h8)
	) name3052 (
		\sa20_reg[7]/NET0131 ,
		_w711_,
		_w3585_
	);
	LUT3 #(
		.INIT('h13)
	) name3053 (
		_w665_,
		_w663_,
		_w3383_,
		_w3586_
	);
	LUT3 #(
		.INIT('h40)
	) name3054 (
		_w3585_,
		_w3584_,
		_w3586_,
		_w3587_
	);
	LUT3 #(
		.INIT('h15)
	) name3055 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w701_,
		_w3588_
	);
	LUT2 #(
		.INIT('h8)
	) name3056 (
		_w728_,
		_w715_,
		_w3589_
	);
	LUT3 #(
		.INIT('h54)
	) name3057 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w3590_
	);
	LUT4 #(
		.INIT('h153f)
	) name3058 (
		_w638_,
		_w728_,
		_w715_,
		_w3590_,
		_w3591_
	);
	LUT2 #(
		.INIT('h8)
	) name3059 (
		_w3588_,
		_w3591_,
		_w3592_
	);
	LUT4 #(
		.INIT('h4445)
	) name3060 (
		\sa20_reg[1]/P0001 ,
		_w3580_,
		_w3587_,
		_w3592_,
		_w3593_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name3061 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3594_
	);
	LUT2 #(
		.INIT('h1)
	) name3062 (
		\sa20_reg[2]/P0001 ,
		_w3594_,
		_w3595_
	);
	LUT3 #(
		.INIT('h2a)
	) name3063 (
		\sa20_reg[1]/P0001 ,
		_w700_,
		_w740_,
		_w3596_
	);
	LUT4 #(
		.INIT('h0200)
	) name3064 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3597_
	);
	LUT3 #(
		.INIT('h07)
	) name3065 (
		_w671_,
		_w736_,
		_w3597_,
		_w3598_
	);
	LUT3 #(
		.INIT('h20)
	) name3066 (
		_w3596_,
		_w3595_,
		_w3598_,
		_w3599_
	);
	LUT4 #(
		.INIT('h2000)
	) name3067 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3600_
	);
	LUT4 #(
		.INIT('h0015)
	) name3068 (
		\sa20_reg[1]/P0001 ,
		_w686_,
		_w729_,
		_w3600_,
		_w3601_
	);
	LUT3 #(
		.INIT('h32)
	) name3069 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w3602_
	);
	LUT4 #(
		.INIT('h7707)
	) name3070 (
		\sa20_reg[2]/P0001 ,
		_w666_,
		_w651_,
		_w3602_,
		_w3603_
	);
	LUT2 #(
		.INIT('h8)
	) name3071 (
		_w3601_,
		_w3603_,
		_w3604_
	);
	LUT3 #(
		.INIT('h01)
	) name3072 (
		\sa20_reg[2]/P0001 ,
		_w708_,
		_w3534_,
		_w3605_
	);
	LUT3 #(
		.INIT('h01)
	) name3073 (
		_w680_,
		_w707_,
		_w740_,
		_w3606_
	);
	LUT4 #(
		.INIT('h23af)
	) name3074 (
		_w737_,
		_w717_,
		_w3605_,
		_w3606_,
		_w3607_
	);
	LUT4 #(
		.INIT('haa02)
	) name3075 (
		\sa20_reg[0]/P0001 ,
		_w3599_,
		_w3604_,
		_w3607_,
		_w3608_
	);
	LUT4 #(
		.INIT('haa80)
	) name3076 (
		\sa20_reg[3]/P0001 ,
		_w697_,
		_w3346_,
		_w3576_,
		_w3609_
	);
	LUT3 #(
		.INIT('h23)
	) name3077 (
		\sa20_reg[7]/NET0131 ,
		_w705_,
		_w711_,
		_w3610_
	);
	LUT3 #(
		.INIT('h45)
	) name3078 (
		\sa20_reg[2]/P0001 ,
		_w3511_,
		_w3610_,
		_w3611_
	);
	LUT4 #(
		.INIT('h153f)
	) name3079 (
		\sa20_reg[4]/P0001 ,
		_w662_,
		_w692_,
		_w708_,
		_w3612_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name3080 (
		\sa20_reg[5]/P0001 ,
		_w641_,
		_w735_,
		_w3529_,
		_w3613_
	);
	LUT2 #(
		.INIT('h8)
	) name3081 (
		_w3612_,
		_w3613_,
		_w3614_
	);
	LUT4 #(
		.INIT('h1311)
	) name3082 (
		\sa20_reg[1]/P0001 ,
		_w3609_,
		_w3611_,
		_w3614_,
		_w3615_
	);
	LUT4 #(
		.INIT('h0100)
	) name3083 (
		_w3583_,
		_w3608_,
		_w3593_,
		_w3615_,
		_w3616_
	);
	LUT3 #(
		.INIT('h69)
	) name3084 (
		_w933_,
		_w3445_,
		_w3616_,
		_w3617_
	);
	LUT3 #(
		.INIT('h69)
	) name3085 (
		\u0_w_reg[2][21]/P0001 ,
		_w3205_,
		_w3557_,
		_w3618_
	);
	LUT3 #(
		.INIT('h82)
	) name3086 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[53]/P0001 ,
		\u0_w_reg[2][21]/P0001 ,
		_w3619_
	);
	LUT4 #(
		.INIT('h00eb)
	) name3087 (
		\ld_r_reg/P0001 ,
		_w3617_,
		_w3618_,
		_w3619_,
		_w3620_
	);
	LUT4 #(
		.INIT('h4bb4)
	) name3088 (
		_w775_,
		_w821_,
		_w933_,
		_w3616_,
		_w3621_
	);
	LUT4 #(
		.INIT('h4000)
	) name3089 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3622_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name3090 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3623_
	);
	LUT4 #(
		.INIT('h0200)
	) name3091 (
		\sa31_reg[2]/P0001 ,
		_w977_,
		_w3622_,
		_w3623_,
		_w3624_
	);
	LUT4 #(
		.INIT('h2000)
	) name3092 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3625_
	);
	LUT3 #(
		.INIT('h01)
	) name3093 (
		\sa31_reg[2]/P0001 ,
		_w3169_,
		_w3625_,
		_w3626_
	);
	LUT3 #(
		.INIT('h23)
	) name3094 (
		_w1031_,
		_w3624_,
		_w3626_,
		_w3627_
	);
	LUT3 #(
		.INIT('h20)
	) name3095 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w3628_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name3096 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3629_
	);
	LUT2 #(
		.INIT('h1)
	) name3097 (
		\sa31_reg[2]/P0001 ,
		_w3629_,
		_w3630_
	);
	LUT4 #(
		.INIT('h0200)
	) name3098 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3631_
	);
	LUT4 #(
		.INIT('h002a)
	) name3099 (
		\sa31_reg[1]/P0001 ,
		_w947_,
		_w1035_,
		_w3631_,
		_w3632_
	);
	LUT3 #(
		.INIT('h10)
	) name3100 (
		_w3183_,
		_w3630_,
		_w3632_,
		_w3633_
	);
	LUT3 #(
		.INIT('h45)
	) name3101 (
		\sa31_reg[1]/P0001 ,
		\sa31_reg[2]/P0001 ,
		_w3173_,
		_w3634_
	);
	LUT2 #(
		.INIT('h1)
	) name3102 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w3635_
	);
	LUT3 #(
		.INIT('h32)
	) name3103 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w3636_
	);
	LUT2 #(
		.INIT('h2)
	) name3104 (
		_w944_,
		_w3636_,
		_w3637_
	);
	LUT4 #(
		.INIT('h2000)
	) name3105 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3638_
	);
	LUT2 #(
		.INIT('h8)
	) name3106 (
		\sa31_reg[2]/P0001 ,
		_w962_,
		_w3639_
	);
	LUT3 #(
		.INIT('h07)
	) name3107 (
		\sa31_reg[2]/P0001 ,
		_w962_,
		_w3638_,
		_w3640_
	);
	LUT3 #(
		.INIT('h20)
	) name3108 (
		_w3634_,
		_w3637_,
		_w3640_,
		_w3641_
	);
	LUT4 #(
		.INIT('h888a)
	) name3109 (
		\sa31_reg[0]/P0002 ,
		_w3627_,
		_w3633_,
		_w3641_,
		_w3642_
	);
	LUT4 #(
		.INIT('h0100)
	) name3110 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3643_
	);
	LUT4 #(
		.INIT('h5504)
	) name3111 (
		\sa31_reg[2]/P0001 ,
		_w938_,
		_w984_,
		_w3643_,
		_w3644_
	);
	LUT2 #(
		.INIT('h2)
	) name3112 (
		\sa31_reg[1]/P0001 ,
		_w972_,
		_w3645_
	);
	LUT4 #(
		.INIT('h0080)
	) name3113 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3646_
	);
	LUT3 #(
		.INIT('h13)
	) name3114 (
		_w992_,
		_w3646_,
		_w3628_,
		_w3647_
	);
	LUT3 #(
		.INIT('h40)
	) name3115 (
		_w3644_,
		_w3645_,
		_w3647_,
		_w3648_
	);
	LUT4 #(
		.INIT('h1000)
	) name3116 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w3649_
	);
	LUT3 #(
		.INIT('h54)
	) name3117 (
		\sa31_reg[7]/P0001 ,
		_w1035_,
		_w3649_,
		_w3650_
	);
	LUT4 #(
		.INIT('h0002)
	) name3118 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3651_
	);
	LUT4 #(
		.INIT('h8000)
	) name3119 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w3652_
	);
	LUT3 #(
		.INIT('h01)
	) name3120 (
		\sa31_reg[1]/P0001 ,
		_w3651_,
		_w3652_,
		_w3653_
	);
	LUT2 #(
		.INIT('h4)
	) name3121 (
		_w3650_,
		_w3653_,
		_w3654_
	);
	LUT4 #(
		.INIT('h0100)
	) name3122 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w3655_
	);
	LUT4 #(
		.INIT('haa20)
	) name3123 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w953_,
		_w3655_,
		_w3656_
	);
	LUT4 #(
		.INIT('h0004)
	) name3124 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3657_
	);
	LUT4 #(
		.INIT('h3310)
	) name3125 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		_w3188_,
		_w3657_,
		_w3658_
	);
	LUT2 #(
		.INIT('h1)
	) name3126 (
		_w3656_,
		_w3658_,
		_w3659_
	);
	LUT4 #(
		.INIT('h0155)
	) name3127 (
		\sa31_reg[0]/P0002 ,
		_w3648_,
		_w3654_,
		_w3659_,
		_w3660_
	);
	LUT4 #(
		.INIT('h0010)
	) name3128 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3661_
	);
	LUT4 #(
		.INIT('hc480)
	) name3129 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		_w997_,
		_w3661_,
		_w3662_
	);
	LUT2 #(
		.INIT('h8)
	) name3130 (
		\sa31_reg[7]/P0001 ,
		_w1018_,
		_w3663_
	);
	LUT3 #(
		.INIT('h07)
	) name3131 (
		_w1001_,
		_w1030_,
		_w1005_,
		_w3664_
	);
	LUT3 #(
		.INIT('h45)
	) name3132 (
		\sa31_reg[2]/P0001 ,
		_w3663_,
		_w3664_,
		_w3665_
	);
	LUT3 #(
		.INIT('h2a)
	) name3133 (
		\sa31_reg[1]/P0001 ,
		_w964_,
		_w981_,
		_w3666_
	);
	LUT4 #(
		.INIT('h8000)
	) name3134 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3667_
	);
	LUT2 #(
		.INIT('h4)
	) name3135 (
		\sa31_reg[5]/P0001 ,
		_w3667_,
		_w3668_
	);
	LUT4 #(
		.INIT('h0020)
	) name3136 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3669_
	);
	LUT4 #(
		.INIT('h13df)
	) name3137 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w3177_,
		_w3669_,
		_w3670_
	);
	LUT3 #(
		.INIT('h40)
	) name3138 (
		_w3668_,
		_w3666_,
		_w3670_,
		_w3671_
	);
	LUT2 #(
		.INIT('h8)
	) name3139 (
		_w1003_,
		_w3164_,
		_w3672_
	);
	LUT3 #(
		.INIT('h15)
	) name3140 (
		\sa31_reg[2]/P0001 ,
		_w1003_,
		_w3164_,
		_w3673_
	);
	LUT4 #(
		.INIT('h0400)
	) name3141 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w3674_
	);
	LUT2 #(
		.INIT('h1)
	) name3142 (
		_w3152_,
		_w3674_,
		_w3675_
	);
	LUT2 #(
		.INIT('h9)
	) name3143 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w3676_
	);
	LUT4 #(
		.INIT('h020a)
	) name3144 (
		\sa31_reg[2]/P0001 ,
		_w3177_,
		_w3168_,
		_w3676_,
		_w3677_
	);
	LUT4 #(
		.INIT('h0020)
	) name3145 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w3678_
	);
	LUT4 #(
		.INIT('h0004)
	) name3146 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3679_
	);
	LUT2 #(
		.INIT('h1)
	) name3147 (
		_w3678_,
		_w3679_,
		_w3680_
	);
	LUT4 #(
		.INIT('h0777)
	) name3148 (
		_w3673_,
		_w3675_,
		_w3677_,
		_w3680_,
		_w3681_
	);
	LUT2 #(
		.INIT('h8)
	) name3149 (
		_w961_,
		_w1030_,
		_w3682_
	);
	LUT3 #(
		.INIT('h15)
	) name3150 (
		\sa31_reg[1]/P0001 ,
		_w996_,
		_w997_,
		_w3683_
	);
	LUT2 #(
		.INIT('h4)
	) name3151 (
		_w3682_,
		_w3683_,
		_w3684_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3152 (
		_w3665_,
		_w3671_,
		_w3681_,
		_w3684_,
		_w3685_
	);
	LUT4 #(
		.INIT('h0001)
	) name3153 (
		_w3660_,
		_w3662_,
		_w3642_,
		_w3685_,
		_w3686_
	);
	LUT3 #(
		.INIT('h69)
	) name3154 (
		\u0_w_reg[2][13]/P0001 ,
		_w3205_,
		_w3686_,
		_w3687_
	);
	LUT3 #(
		.INIT('h28)
	) name3155 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[45]/P0001 ,
		\u0_w_reg[2][13]/P0001 ,
		_w3688_
	);
	LUT4 #(
		.INIT('hff14)
	) name3156 (
		\ld_r_reg/P0001 ,
		_w3621_,
		_w3687_,
		_w3688_,
		_w3689_
	);
	LUT3 #(
		.INIT('h69)
	) name3157 (
		_w637_,
		_w3142_,
		_w3557_,
		_w3690_
	);
	LUT4 #(
		.INIT('h5655)
	) name3158 (
		\u0_w_reg[2][14]/P0001 ,
		_w980_,
		_w1009_,
		_w1038_,
		_w3691_
	);
	LUT2 #(
		.INIT('h6)
	) name3159 (
		_w3205_,
		_w3691_,
		_w3692_
	);
	LUT3 #(
		.INIT('h82)
	) name3160 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[46]/P0001 ,
		\u0_w_reg[2][14]/P0001 ,
		_w3693_
	);
	LUT4 #(
		.INIT('h00eb)
	) name3161 (
		\ld_r_reg/P0001 ,
		_w3690_,
		_w3692_,
		_w3693_,
		_w3694_
	);
	LUT4 #(
		.INIT('h0045)
	) name3162 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w534_,
		_w623_,
		_w3695_
	);
	LUT3 #(
		.INIT('h02)
	) name3163 (
		\sa13_reg[2]/P0001 ,
		_w748_,
		_w3409_,
		_w3696_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name3164 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		_w619_,
		_w3395_,
		_w3697_
	);
	LUT4 #(
		.INIT('h0155)
	) name3165 (
		\sa13_reg[1]/P0001 ,
		_w3695_,
		_w3696_,
		_w3697_,
		_w3698_
	);
	LUT4 #(
		.INIT('h0800)
	) name3166 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w3699_
	);
	LUT4 #(
		.INIT('h5554)
	) name3167 (
		\sa13_reg[2]/P0001 ,
		_w588_,
		_w598_,
		_w3699_,
		_w3700_
	);
	LUT3 #(
		.INIT('ha8)
	) name3168 (
		\sa13_reg[2]/P0001 ,
		_w572_,
		_w585_,
		_w3701_
	);
	LUT3 #(
		.INIT('h01)
	) name3169 (
		_w750_,
		_w776_,
		_w790_,
		_w3702_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3170 (
		\sa13_reg[1]/P0001 ,
		_w3701_,
		_w3700_,
		_w3702_,
		_w3703_
	);
	LUT4 #(
		.INIT('h153f)
	) name3171 (
		\sa13_reg[5]/P0001 ,
		_w562_,
		_w784_,
		_w3396_,
		_w3704_
	);
	LUT4 #(
		.INIT('hffa8)
	) name3172 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3705_
	);
	LUT2 #(
		.INIT('h2)
	) name3173 (
		_w583_,
		_w3705_,
		_w3706_
	);
	LUT4 #(
		.INIT('h007f)
	) name3174 (
		\sa13_reg[4]/P0001 ,
		_w543_,
		_w594_,
		_w617_,
		_w3707_
	);
	LUT4 #(
		.INIT('h3200)
	) name3175 (
		\sa13_reg[2]/P0001 ,
		_w3706_,
		_w3704_,
		_w3707_,
		_w3708_
	);
	LUT4 #(
		.INIT('h5455)
	) name3176 (
		\sa13_reg[0]/P0001 ,
		_w3703_,
		_w3698_,
		_w3708_,
		_w3709_
	);
	LUT3 #(
		.INIT('h07)
	) name3177 (
		_w571_,
		_w542_,
		_w534_,
		_w3710_
	);
	LUT3 #(
		.INIT('h10)
	) name3178 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w3711_
	);
	LUT3 #(
		.INIT('h20)
	) name3179 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w3712_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3180 (
		\sa13_reg[2]/P0001 ,
		_w3395_,
		_w3712_,
		_w3711_,
		_w3713_
	);
	LUT3 #(
		.INIT('ha2)
	) name3181 (
		\sa13_reg[1]/P0001 ,
		_w3710_,
		_w3713_,
		_w3714_
	);
	LUT4 #(
		.INIT('h2000)
	) name3182 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3715_
	);
	LUT4 #(
		.INIT('hdff7)
	) name3183 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3716_
	);
	LUT3 #(
		.INIT('h45)
	) name3184 (
		\sa13_reg[3]/P0001 ,
		_w3715_,
		_w3716_,
		_w3717_
	);
	LUT4 #(
		.INIT('h7c7f)
	) name3185 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w3718_
	);
	LUT2 #(
		.INIT('h1)
	) name3186 (
		\sa13_reg[7]/NET0131 ,
		_w3718_,
		_w3719_
	);
	LUT3 #(
		.INIT('h10)
	) name3187 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w3720_
	);
	LUT4 #(
		.INIT('h45cf)
	) name3188 (
		_w561_,
		_w628_,
		_w757_,
		_w3720_,
		_w3721_
	);
	LUT3 #(
		.INIT('h45)
	) name3189 (
		\sa13_reg[1]/P0001 ,
		_w3719_,
		_w3721_,
		_w3722_
	);
	LUT4 #(
		.INIT('h0001)
	) name3190 (
		_w748_,
		_w795_,
		_w3309_,
		_w3297_,
		_w3723_
	);
	LUT2 #(
		.INIT('h1)
	) name3191 (
		\sa13_reg[2]/P0001 ,
		_w3723_,
		_w3724_
	);
	LUT4 #(
		.INIT('h0001)
	) name3192 (
		_w3714_,
		_w3722_,
		_w3724_,
		_w3717_,
		_w3725_
	);
	LUT4 #(
		.INIT('h0203)
	) name3193 (
		\sa13_reg[3]/P0001 ,
		_w545_,
		_w619_,
		_w615_,
		_w3726_
	);
	LUT4 #(
		.INIT('hedff)
	) name3194 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w542_,
		_w3727_
	);
	LUT4 #(
		.INIT('h0155)
	) name3195 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[2]/P0001 ,
		_w3726_,
		_w3727_,
		_w3728_
	);
	LUT2 #(
		.INIT('h8)
	) name3196 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[2]/P0001 ,
		_w3729_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name3197 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3730_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3198 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w600_,
		_w3730_,
		_w3731_
	);
	LUT2 #(
		.INIT('h2)
	) name3199 (
		_w3729_,
		_w3731_,
		_w3732_
	);
	LUT2 #(
		.INIT('h4)
	) name3200 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[2]/P0001 ,
		_w3733_
	);
	LUT4 #(
		.INIT('h0100)
	) name3201 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3734_
	);
	LUT4 #(
		.INIT('h0007)
	) name3202 (
		\sa13_reg[4]/P0001 ,
		_w572_,
		_w617_,
		_w3734_,
		_w3735_
	);
	LUT2 #(
		.INIT('h2)
	) name3203 (
		_w3733_,
		_w3735_,
		_w3736_
	);
	LUT4 #(
		.INIT('hffbe)
	) name3204 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3737_
	);
	LUT4 #(
		.INIT('h40cc)
	) name3205 (
		_w562_,
		_w632_,
		_w784_,
		_w3737_,
		_w3738_
	);
	LUT2 #(
		.INIT('h8)
	) name3206 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w3739_
	);
	LUT2 #(
		.INIT('h8)
	) name3207 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w3740_
	);
	LUT4 #(
		.INIT('h0001)
	) name3208 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w3741_
	);
	LUT4 #(
		.INIT('h0777)
	) name3209 (
		_w579_,
		_w3739_,
		_w3740_,
		_w3741_,
		_w3742_
	);
	LUT3 #(
		.INIT('h10)
	) name3210 (
		_w3307_,
		_w3738_,
		_w3742_,
		_w3743_
	);
	LUT4 #(
		.INIT('h0100)
	) name3211 (
		_w3736_,
		_w3732_,
		_w3728_,
		_w3743_,
		_w3744_
	);
	LUT4 #(
		.INIT('h3100)
	) name3212 (
		\sa13_reg[0]/P0001 ,
		_w3709_,
		_w3725_,
		_w3744_,
		_w3745_
	);
	LUT3 #(
		.INIT('h13)
	) name3213 (
		_w831_,
		_w895_,
		_w824_,
		_w3746_
	);
	LUT3 #(
		.INIT('h32)
	) name3214 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3747_
	);
	LUT4 #(
		.INIT('h3120)
	) name3215 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3748_
	);
	LUT3 #(
		.INIT('h80)
	) name3216 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3749_
	);
	LUT3 #(
		.INIT('ha8)
	) name3217 (
		\sa02_reg[2]/P0001 ,
		_w3748_,
		_w3749_,
		_w3750_
	);
	LUT3 #(
		.INIT('ha2)
	) name3218 (
		\sa02_reg[1]/P0001 ,
		_w3746_,
		_w3750_,
		_w3751_
	);
	LUT2 #(
		.INIT('h2)
	) name3219 (
		_w869_,
		_w3123_,
		_w3752_
	);
	LUT4 #(
		.INIT('h0103)
	) name3220 (
		_w857_,
		_w852_,
		_w862_,
		_w910_,
		_w3753_
	);
	LUT3 #(
		.INIT('h45)
	) name3221 (
		\sa02_reg[1]/P0001 ,
		_w3752_,
		_w3753_,
		_w3754_
	);
	LUT4 #(
		.INIT('h5054)
	) name3222 (
		\sa02_reg[3]/P0001 ,
		_w882_,
		_w3247_,
		_w3468_,
		_w3755_
	);
	LUT4 #(
		.INIT('hffe7)
	) name3223 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3756_
	);
	LUT4 #(
		.INIT('h5455)
	) name3224 (
		\sa02_reg[2]/P0001 ,
		_w3119_,
		_w3453_,
		_w3756_,
		_w3757_
	);
	LUT2 #(
		.INIT('h1)
	) name3225 (
		_w3755_,
		_w3757_,
		_w3758_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3226 (
		\sa02_reg[0]/P0001 ,
		_w3751_,
		_w3754_,
		_w3758_,
		_w3759_
	);
	LUT4 #(
		.INIT('h5540)
	) name3227 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3076_,
		_w3118_,
		_w3760_
	);
	LUT2 #(
		.INIT('h8)
	) name3228 (
		_w884_,
		_w3077_,
		_w3761_
	);
	LUT3 #(
		.INIT('h15)
	) name3229 (
		\sa02_reg[1]/P0001 ,
		_w861_,
		_w875_,
		_w3762_
	);
	LUT3 #(
		.INIT('h10)
	) name3230 (
		_w3761_,
		_w3760_,
		_w3762_,
		_w3763_
	);
	LUT3 #(
		.INIT('h10)
	) name3231 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3764_
	);
	LUT4 #(
		.INIT('hf7fc)
	) name3232 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w3765_
	);
	LUT3 #(
		.INIT('h45)
	) name3233 (
		\sa02_reg[2]/P0001 ,
		_w3764_,
		_w3765_,
		_w3766_
	);
	LUT4 #(
		.INIT('h0002)
	) name3234 (
		\sa02_reg[1]/P0001 ,
		_w885_,
		_w846_,
		_w848_,
		_w3767_
	);
	LUT2 #(
		.INIT('h4)
	) name3235 (
		_w3766_,
		_w3767_,
		_w3768_
	);
	LUT4 #(
		.INIT('hffa8)
	) name3236 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3769_
	);
	LUT2 #(
		.INIT('h2)
	) name3237 (
		_w833_,
		_w3769_,
		_w3770_
	);
	LUT4 #(
		.INIT('h00df)
	) name3238 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w852_,
		_w914_,
		_w3771_
	);
	LUT2 #(
		.INIT('h4)
	) name3239 (
		_w3770_,
		_w3771_,
		_w3772_
	);
	LUT4 #(
		.INIT('h4000)
	) name3240 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3773_
	);
	LUT3 #(
		.INIT('hc8)
	) name3241 (
		_w900_,
		_w3129_,
		_w3773_,
		_w3774_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name3242 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3775_
	);
	LUT2 #(
		.INIT('h2)
	) name3243 (
		_w3086_,
		_w3775_,
		_w3776_
	);
	LUT4 #(
		.INIT('h153f)
	) name3244 (
		_w856_,
		_w861_,
		_w875_,
		_w858_,
		_w3777_
	);
	LUT4 #(
		.INIT('h0032)
	) name3245 (
		\sa02_reg[2]/P0001 ,
		_w3776_,
		_w3777_,
		_w3774_,
		_w3778_
	);
	LUT4 #(
		.INIT('he000)
	) name3246 (
		_w3763_,
		_w3768_,
		_w3772_,
		_w3778_,
		_w3779_
	);
	LUT4 #(
		.INIT('h0100)
	) name3247 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3780_
	);
	LUT4 #(
		.INIT('h0007)
	) name3248 (
		_w831_,
		_w832_,
		_w914_,
		_w3780_,
		_w3781_
	);
	LUT4 #(
		.INIT('hedff)
	) name3249 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w824_,
		_w3782_
	);
	LUT4 #(
		.INIT('h0455)
	) name3250 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		_w3781_,
		_w3782_,
		_w3783_
	);
	LUT4 #(
		.INIT('h8000)
	) name3251 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w3784_
	);
	LUT4 #(
		.INIT('haa08)
	) name3252 (
		\sa02_reg[1]/P0001 ,
		_w882_,
		_w3487_,
		_w3784_,
		_w3785_
	);
	LUT4 #(
		.INIT('haabf)
	) name3253 (
		\sa02_reg[5]/P0001 ,
		_w827_,
		_w824_,
		_w929_,
		_w3786_
	);
	LUT3 #(
		.INIT('h8a)
	) name3254 (
		\sa02_reg[2]/P0001 ,
		_w3785_,
		_w3786_,
		_w3787_
	);
	LUT2 #(
		.INIT('h1)
	) name3255 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		_w3788_
	);
	LUT4 #(
		.INIT('h0020)
	) name3256 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3789_
	);
	LUT4 #(
		.INIT('h000b)
	) name3257 (
		\sa02_reg[7]/NET0131 ,
		_w855_,
		_w3083_,
		_w3789_,
		_w3790_
	);
	LUT4 #(
		.INIT('hffbe)
	) name3258 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3791_
	);
	LUT4 #(
		.INIT('h2300)
	) name3259 (
		_w856_,
		_w885_,
		_w858_,
		_w3791_,
		_w3792_
	);
	LUT4 #(
		.INIT('hfedc)
	) name3260 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		_w3790_,
		_w3792_,
		_w3793_
	);
	LUT3 #(
		.INIT('h10)
	) name3261 (
		_w3787_,
		_w3783_,
		_w3793_,
		_w3794_
	);
	LUT4 #(
		.INIT('h0e00)
	) name3262 (
		\sa02_reg[0]/P0001 ,
		_w3779_,
		_w3759_,
		_w3794_,
		_w3795_
	);
	LUT2 #(
		.INIT('h6)
	) name3263 (
		_w3745_,
		_w3795_,
		_w3796_
	);
	LUT4 #(
		.INIT('h0001)
	) name3264 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3797_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name3265 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3798_
	);
	LUT3 #(
		.INIT('h8a)
	) name3266 (
		\sa02_reg[2]/P0001 ,
		_w3797_,
		_w3798_,
		_w3799_
	);
	LUT2 #(
		.INIT('h2)
	) name3267 (
		_w837_,
		_w3252_,
		_w3800_
	);
	LUT4 #(
		.INIT('h0100)
	) name3268 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3801_
	);
	LUT3 #(
		.INIT('h13)
	) name3269 (
		_w3131_,
		_w3491_,
		_w3801_,
		_w3802_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3270 (
		\sa02_reg[0]/P0001 ,
		_w3800_,
		_w3799_,
		_w3802_,
		_w3803_
	);
	LUT3 #(
		.INIT('h67)
	) name3271 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3804_
	);
	LUT2 #(
		.INIT('h2)
	) name3272 (
		_w870_,
		_w3804_,
		_w3805_
	);
	LUT4 #(
		.INIT('hff4b)
	) name3273 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3806_
	);
	LUT2 #(
		.INIT('h1)
	) name3274 (
		\sa02_reg[3]/P0001 ,
		_w3806_,
		_w3807_
	);
	LUT3 #(
		.INIT('h15)
	) name3275 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		_w846_,
		_w3808_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3276 (
		_w921_,
		_w3805_,
		_w3807_,
		_w3808_,
		_w3809_
	);
	LUT3 #(
		.INIT('h54)
	) name3277 (
		\sa02_reg[1]/P0001 ,
		_w3803_,
		_w3809_,
		_w3810_
	);
	LUT4 #(
		.INIT('h153f)
	) name3278 (
		_w869_,
		_w847_,
		_w923_,
		_w3090_,
		_w3811_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name3279 (
		\sa02_reg[7]/NET0131 ,
		_w900_,
		_w3091_,
		_w3114_,
		_w3812_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3280 (
		\sa02_reg[1]/P0001 ,
		_w899_,
		_w3811_,
		_w3812_,
		_w3813_
	);
	LUT4 #(
		.INIT('h0777)
	) name3281 (
		\sa02_reg[6]/NET0131 ,
		_w3102_,
		_w3123_,
		_w3453_,
		_w3814_
	);
	LUT2 #(
		.INIT('h4)
	) name3282 (
		_w3813_,
		_w3814_,
		_w3815_
	);
	LUT4 #(
		.INIT('h8000)
	) name3283 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3816_
	);
	LUT4 #(
		.INIT('h0007)
	) name3284 (
		_w856_,
		_w858_,
		_w3114_,
		_w3816_,
		_w3817_
	);
	LUT2 #(
		.INIT('h1)
	) name3285 (
		\sa02_reg[2]/P0001 ,
		_w3817_,
		_w3818_
	);
	LUT2 #(
		.INIT('h8)
	) name3286 (
		_w845_,
		_w3449_,
		_w3819_
	);
	LUT4 #(
		.INIT('h8000)
	) name3287 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3820_
	);
	LUT4 #(
		.INIT('h0007)
	) name3288 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3821_
	);
	LUT3 #(
		.INIT('h01)
	) name3289 (
		_w3801_,
		_w3820_,
		_w3821_,
		_w3822_
	);
	LUT3 #(
		.INIT('h8a)
	) name3290 (
		\sa02_reg[1]/P0001 ,
		_w3819_,
		_w3822_,
		_w3823_
	);
	LUT4 #(
		.INIT('haf8c)
	) name3291 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		_w825_,
		_w3209_,
		_w3824_
	);
	LUT3 #(
		.INIT('hb9)
	) name3292 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3825_
	);
	LUT3 #(
		.INIT('h40)
	) name3293 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3826_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3294 (
		_w837_,
		_w845_,
		_w3825_,
		_w3826_,
		_w3827_
	);
	LUT4 #(
		.INIT('hfa32)
	) name3295 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		_w3824_,
		_w3827_,
		_w3828_
	);
	LUT4 #(
		.INIT('h5455)
	) name3296 (
		\sa02_reg[0]/P0001 ,
		_w3818_,
		_w3823_,
		_w3828_,
		_w3829_
	);
	LUT4 #(
		.INIT('h4041)
	) name3297 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3830_
	);
	LUT3 #(
		.INIT('ha8)
	) name3298 (
		\sa02_reg[1]/P0001 ,
		_w3118_,
		_w3830_,
		_w3831_
	);
	LUT3 #(
		.INIT('h07)
	) name3299 (
		_w856_,
		_w858_,
		_w3446_,
		_w3832_
	);
	LUT3 #(
		.INIT('h2a)
	) name3300 (
		\sa02_reg[2]/P0001 ,
		_w3084_,
		_w3832_,
		_w3833_
	);
	LUT4 #(
		.INIT('h0040)
	) name3301 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w3834_
	);
	LUT3 #(
		.INIT('h54)
	) name3302 (
		\sa02_reg[2]/P0001 ,
		_w3248_,
		_w3834_,
		_w3835_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name3303 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w3836_
	);
	LUT2 #(
		.INIT('h2)
	) name3304 (
		_w829_,
		_w3836_,
		_w3837_
	);
	LUT3 #(
		.INIT('h07)
	) name3305 (
		_w837_,
		_w828_,
		_w3453_,
		_w3838_
	);
	LUT3 #(
		.INIT('h10)
	) name3306 (
		_w3835_,
		_w3837_,
		_w3838_,
		_w3839_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3307 (
		\sa02_reg[0]/P0001 ,
		_w3833_,
		_w3831_,
		_w3839_,
		_w3840_
	);
	LUT4 #(
		.INIT('h0100)
	) name3308 (
		_w3810_,
		_w3829_,
		_w3840_,
		_w3815_,
		_w3841_
	);
	LUT4 #(
		.INIT('h9669)
	) name3309 (
		_w3265_,
		_w3745_,
		_w3795_,
		_w3841_,
		_w3842_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3310 (
		\sa31_reg[2]/P0001 ,
		_w1026_,
		_w3146_,
		_w3188_,
		_w3843_
	);
	LUT3 #(
		.INIT('h80)
	) name3311 (
		\sa31_reg[4]/P0001 ,
		_w949_,
		_w3177_,
		_w3844_
	);
	LUT3 #(
		.INIT('h8a)
	) name3312 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3845_
	);
	LUT4 #(
		.INIT('h0010)
	) name3313 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w3846_
	);
	LUT3 #(
		.INIT('h0d)
	) name3314 (
		_w984_,
		_w3845_,
		_w3846_,
		_w3847_
	);
	LUT4 #(
		.INIT('h5455)
	) name3315 (
		\sa31_reg[1]/P0001 ,
		_w3844_,
		_w3843_,
		_w3847_,
		_w3848_
	);
	LUT2 #(
		.INIT('h1)
	) name3316 (
		_w946_,
		_w3643_,
		_w3849_
	);
	LUT3 #(
		.INIT('h2a)
	) name3317 (
		\sa31_reg[2]/P0001 ,
		_w3181_,
		_w3849_,
		_w3850_
	);
	LUT4 #(
		.INIT('h4041)
	) name3318 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3851_
	);
	LUT3 #(
		.INIT('ha8)
	) name3319 (
		\sa31_reg[1]/P0001 ,
		_w1011_,
		_w3851_,
		_w3852_
	);
	LUT4 #(
		.INIT('h0040)
	) name3320 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w3853_
	);
	LUT4 #(
		.INIT('h8000)
	) name3321 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3854_
	);
	LUT3 #(
		.INIT('h54)
	) name3322 (
		\sa31_reg[2]/P0001 ,
		_w3853_,
		_w3854_,
		_w3855_
	);
	LUT3 #(
		.INIT('h20)
	) name3323 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w3856_
	);
	LUT3 #(
		.INIT('h02)
	) name3324 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w3857_
	);
	LUT3 #(
		.INIT('h54)
	) name3325 (
		\sa31_reg[2]/P0001 ,
		_w3856_,
		_w3857_,
		_w3858_
	);
	LUT4 #(
		.INIT('h0040)
	) name3326 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3859_
	);
	LUT3 #(
		.INIT('h07)
	) name3327 (
		_w984_,
		_w3177_,
		_w3859_,
		_w3860_
	);
	LUT4 #(
		.INIT('h0100)
	) name3328 (
		_w3852_,
		_w3858_,
		_w3855_,
		_w3860_,
		_w3861_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3329 (
		\sa31_reg[0]/P0002 ,
		_w3850_,
		_w3848_,
		_w3861_,
		_w3862_
	);
	LUT4 #(
		.INIT('h0010)
	) name3330 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w3863_
	);
	LUT4 #(
		.INIT('hbbef)
	) name3331 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w3864_
	);
	LUT2 #(
		.INIT('h1)
	) name3332 (
		\sa31_reg[7]/P0001 ,
		_w3864_,
		_w3865_
	);
	LUT4 #(
		.INIT('h0010)
	) name3333 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3866_
	);
	LUT3 #(
		.INIT('h07)
	) name3334 (
		_w940_,
		_w3164_,
		_w3866_,
		_w3867_
	);
	LUT3 #(
		.INIT('h45)
	) name3335 (
		\sa31_reg[2]/P0001 ,
		_w3865_,
		_w3867_,
		_w3868_
	);
	LUT3 #(
		.INIT('h01)
	) name3336 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w3869_
	);
	LUT4 #(
		.INIT('h0001)
	) name3337 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w3870_
	);
	LUT2 #(
		.INIT('h8)
	) name3338 (
		\sa31_reg[7]/P0001 ,
		_w3870_,
		_w3871_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3339 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w1018_,
		_w3870_,
		_w3872_
	);
	LUT2 #(
		.INIT('h1)
	) name3340 (
		_w3201_,
		_w3872_,
		_w3873_
	);
	LUT3 #(
		.INIT('h45)
	) name3341 (
		\sa31_reg[1]/P0001 ,
		_w3868_,
		_w3873_,
		_w3874_
	);
	LUT4 #(
		.INIT('h8000)
	) name3342 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3875_
	);
	LUT4 #(
		.INIT('h0007)
	) name3343 (
		\sa31_reg[7]/P0001 ,
		_w970_,
		_w3875_,
		_w3870_,
		_w3876_
	);
	LUT2 #(
		.INIT('h1)
	) name3344 (
		\sa31_reg[2]/P0001 ,
		_w3876_,
		_w3877_
	);
	LUT4 #(
		.INIT('hbfef)
	) name3345 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3878_
	);
	LUT2 #(
		.INIT('h1)
	) name3346 (
		\sa31_reg[3]/P0001 ,
		_w3878_,
		_w3879_
	);
	LUT2 #(
		.INIT('h8)
	) name3347 (
		_w967_,
		_w981_,
		_w3880_
	);
	LUT4 #(
		.INIT('h0007)
	) name3348 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3881_
	);
	LUT4 #(
		.INIT('h0100)
	) name3349 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w3882_
	);
	LUT4 #(
		.INIT('h0002)
	) name3350 (
		\sa31_reg[1]/P0001 ,
		_w3667_,
		_w3881_,
		_w3882_,
		_w3883_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3351 (
		_w3634_,
		_w3879_,
		_w3880_,
		_w3883_,
		_w3884_
	);
	LUT2 #(
		.INIT('h4)
	) name3352 (
		\sa31_reg[1]/P0001 ,
		\sa31_reg[2]/P0001 ,
		_w3885_
	);
	LUT4 #(
		.INIT('h4c00)
	) name3353 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3886_
	);
	LUT3 #(
		.INIT('hb9)
	) name3354 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3887_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3355 (
		_w1015_,
		_w3885_,
		_w3886_,
		_w3887_,
		_w3888_
	);
	LUT4 #(
		.INIT('h5455)
	) name3356 (
		\sa31_reg[0]/P0002 ,
		_w3884_,
		_w3877_,
		_w3888_,
		_w3889_
	);
	LUT4 #(
		.INIT('h3320)
	) name3357 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w3674_,
		_w3678_,
		_w3890_
	);
	LUT4 #(
		.INIT('h4000)
	) name3358 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w3891_
	);
	LUT3 #(
		.INIT('hd8)
	) name3359 (
		\sa31_reg[2]/P0001 ,
		_w977_,
		_w3891_,
		_w3892_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3360 (
		\sa31_reg[1]/P0001 ,
		_w1031_,
		_w3890_,
		_w3892_,
		_w3893_
	);
	LUT4 #(
		.INIT('h135f)
	) name3361 (
		\sa31_reg[6]/NET0131 ,
		_w935_,
		_w982_,
		_w3646_,
		_w3894_
	);
	LUT2 #(
		.INIT('h4)
	) name3362 (
		_w3893_,
		_w3894_,
		_w3895_
	);
	LUT4 #(
		.INIT('h0100)
	) name3363 (
		_w3862_,
		_w3889_,
		_w3874_,
		_w3895_,
		_w3896_
	);
	LUT2 #(
		.INIT('h2)
	) name3364 (
		\sa31_reg[1]/P0001 ,
		_w1010_,
		_w3897_
	);
	LUT4 #(
		.INIT('h020a)
	) name3365 (
		\sa31_reg[1]/P0001 ,
		\sa31_reg[2]/P0001 ,
		_w1010_,
		_w3674_,
		_w3898_
	);
	LUT2 #(
		.INIT('h8)
	) name3366 (
		\sa31_reg[7]/P0001 ,
		_w3674_,
		_w3899_
	);
	LUT3 #(
		.INIT('h54)
	) name3367 (
		\sa31_reg[2]/P0001 ,
		_w948_,
		_w1029_,
		_w3900_
	);
	LUT3 #(
		.INIT('h10)
	) name3368 (
		_w3899_,
		_w3900_,
		_w3898_,
		_w3901_
	);
	LUT4 #(
		.INIT('hf2fa)
	) name3369 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		_w3902_
	);
	LUT2 #(
		.INIT('h2)
	) name3370 (
		\sa31_reg[7]/P0001 ,
		_w3902_,
		_w3903_
	);
	LUT4 #(
		.INIT('h0015)
	) name3371 (
		\sa31_reg[1]/P0001 ,
		_w981_,
		_w3628_,
		_w3651_,
		_w3904_
	);
	LUT2 #(
		.INIT('h4)
	) name3372 (
		_w3903_,
		_w3904_,
		_w3905_
	);
	LUT4 #(
		.INIT('h0008)
	) name3373 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3906_
	);
	LUT4 #(
		.INIT('h7ff7)
	) name3374 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3907_
	);
	LUT3 #(
		.INIT('ha2)
	) name3375 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		_w3907_,
		_w3908_
	);
	LUT3 #(
		.INIT('h15)
	) name3376 (
		\sa31_reg[2]/P0001 ,
		_w996_,
		_w997_,
		_w3909_
	);
	LUT4 #(
		.INIT('h4000)
	) name3377 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3910_
	);
	LUT3 #(
		.INIT('h01)
	) name3378 (
		_w1022_,
		_w3846_,
		_w3910_,
		_w3911_
	);
	LUT2 #(
		.INIT('h8)
	) name3379 (
		_w984_,
		_w3651_,
		_w3912_
	);
	LUT4 #(
		.INIT('h00ea)
	) name3380 (
		_w3908_,
		_w3909_,
		_w3911_,
		_w3912_,
		_w3913_
	);
	LUT4 #(
		.INIT('h0155)
	) name3381 (
		\sa31_reg[0]/P0002 ,
		_w3901_,
		_w3905_,
		_w3913_,
		_w3914_
	);
	LUT4 #(
		.INIT('ha7f7)
	) name3382 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3915_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name3383 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		_w3146_,
		_w3915_,
		_w3916_
	);
	LUT4 #(
		.INIT('h30b0)
	) name3384 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3917_
	);
	LUT3 #(
		.INIT('h02)
	) name3385 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w3918_
	);
	LUT3 #(
		.INIT('h01)
	) name3386 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3919_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3387 (
		_w1021_,
		_w3917_,
		_w3918_,
		_w3919_,
		_w3920_
	);
	LUT4 #(
		.INIT('haabf)
	) name3388 (
		\sa31_reg[5]/P0001 ,
		_w937_,
		_w949_,
		_w3667_,
		_w3921_
	);
	LUT2 #(
		.INIT('h8)
	) name3389 (
		_w941_,
		_w949_,
		_w3922_
	);
	LUT3 #(
		.INIT('h07)
	) name3390 (
		_w934_,
		_w1015_,
		_w3853_,
		_w3923_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3391 (
		\sa31_reg[1]/P0001 ,
		_w3921_,
		_w3922_,
		_w3923_,
		_w3924_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3392 (
		\sa31_reg[0]/P0002 ,
		_w3916_,
		_w3920_,
		_w3924_,
		_w3925_
	);
	LUT4 #(
		.INIT('h7d1d)
	) name3393 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3926_
	);
	LUT2 #(
		.INIT('h1)
	) name3394 (
		\sa31_reg[2]/P0001 ,
		_w3926_,
		_w3927_
	);
	LUT3 #(
		.INIT('h10)
	) name3395 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w3928_
	);
	LUT2 #(
		.INIT('h8)
	) name3396 (
		_w992_,
		_w3928_,
		_w3929_
	);
	LUT3 #(
		.INIT('h04)
	) name3397 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3930_
	);
	LUT3 #(
		.INIT('h23)
	) name3398 (
		_w1014_,
		_w3678_,
		_w3930_,
		_w3931_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3399 (
		\sa31_reg[0]/P0002 ,
		_w3929_,
		_w3927_,
		_w3931_,
		_w3932_
	);
	LUT3 #(
		.INIT('h54)
	) name3400 (
		\sa31_reg[2]/P0001 ,
		_w3846_,
		_w3910_,
		_w3933_
	);
	LUT3 #(
		.INIT('h13)
	) name3401 (
		_w3176_,
		_w3891_,
		_w3928_,
		_w3934_
	);
	LUT2 #(
		.INIT('h4)
	) name3402 (
		_w3933_,
		_w3934_,
		_w3935_
	);
	LUT3 #(
		.INIT('h45)
	) name3403 (
		\sa31_reg[1]/P0001 ,
		_w3932_,
		_w3935_,
		_w3936_
	);
	LUT4 #(
		.INIT('hadfb)
	) name3404 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3937_
	);
	LUT4 #(
		.INIT('h0302)
	) name3405 (
		\sa31_reg[3]/P0001 ,
		_w955_,
		_w3168_,
		_w3937_,
		_w3938_
	);
	LUT2 #(
		.INIT('h2)
	) name3406 (
		_w1021_,
		_w3938_,
		_w3939_
	);
	LUT4 #(
		.INIT('h4000)
	) name3407 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w3940_
	);
	LUT4 #(
		.INIT('h0023)
	) name3408 (
		\sa31_reg[5]/P0001 ,
		_w3148_,
		_w3667_,
		_w3940_,
		_w3941_
	);
	LUT2 #(
		.INIT('h2)
	) name3409 (
		_w3885_,
		_w3941_,
		_w3942_
	);
	LUT4 #(
		.INIT('h23af)
	) name3410 (
		\sa31_reg[6]/NET0131 ,
		_w935_,
		_w953_,
		_w967_,
		_w3943_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name3411 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w3944_
	);
	LUT3 #(
		.INIT('h20)
	) name3412 (
		\sa31_reg[1]/P0001 ,
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		_w3945_
	);
	LUT2 #(
		.INIT('h4)
	) name3413 (
		_w3944_,
		_w3945_,
		_w3946_
	);
	LUT3 #(
		.INIT('h0e)
	) name3414 (
		\sa31_reg[2]/P0001 ,
		_w3943_,
		_w3946_,
		_w3947_
	);
	LUT3 #(
		.INIT('h10)
	) name3415 (
		_w3939_,
		_w3942_,
		_w3947_,
		_w3948_
	);
	LUT4 #(
		.INIT('h0100)
	) name3416 (
		_w3936_,
		_w3925_,
		_w3914_,
		_w3948_,
		_w3949_
	);
	LUT3 #(
		.INIT('h13)
	) name3417 (
		_w647_,
		_w661_,
		_w3510_,
		_w3950_
	);
	LUT3 #(
		.INIT('h80)
	) name3418 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3951_
	);
	LUT4 #(
		.INIT('hcedf)
	) name3419 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3952_
	);
	LUT3 #(
		.INIT('h8a)
	) name3420 (
		\sa20_reg[2]/P0001 ,
		_w3951_,
		_w3952_,
		_w3953_
	);
	LUT3 #(
		.INIT('ha2)
	) name3421 (
		\sa20_reg[1]/P0001 ,
		_w3950_,
		_w3953_,
		_w3954_
	);
	LUT4 #(
		.INIT('h0001)
	) name3422 (
		_w720_,
		_w3326_,
		_w3373_,
		_w3574_,
		_w3955_
	);
	LUT2 #(
		.INIT('h1)
	) name3423 (
		\sa20_reg[2]/P0001 ,
		_w3955_,
		_w3956_
	);
	LUT2 #(
		.INIT('h4)
	) name3424 (
		\sa20_reg[6]/NET0131 ,
		_w3551_,
		_w3957_
	);
	LUT4 #(
		.INIT('h0888)
	) name3425 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3958_
	);
	LUT4 #(
		.INIT('h0207)
	) name3426 (
		_w659_,
		_w655_,
		_w3503_,
		_w3958_,
		_w3959_
	);
	LUT4 #(
		.INIT('h113f)
	) name3427 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w663_,
		_w640_,
		_w3960_
	);
	LUT4 #(
		.INIT('hba00)
	) name3428 (
		\sa20_reg[1]/P0001 ,
		_w3957_,
		_w3959_,
		_w3960_,
		_w3961_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3429 (
		\sa20_reg[0]/P0001 ,
		_w3954_,
		_w3956_,
		_w3961_,
		_w3962_
	);
	LUT4 #(
		.INIT('h5510)
	) name3430 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w640_,
		_w721_,
		_w3963_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name3431 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3964_
	);
	LUT2 #(
		.INIT('h2)
	) name3432 (
		\sa20_reg[2]/P0001 ,
		_w3964_,
		_w3965_
	);
	LUT4 #(
		.INIT('h0777)
	) name3433 (
		_w647_,
		_w667_,
		_w728_,
		_w715_,
		_w3966_
	);
	LUT4 #(
		.INIT('h5455)
	) name3434 (
		\sa20_reg[1]/P0001 ,
		_w3965_,
		_w3963_,
		_w3966_,
		_w3967_
	);
	LUT3 #(
		.INIT('h4c)
	) name3435 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w3968_
	);
	LUT4 #(
		.INIT('h0803)
	) name3436 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w3969_
	);
	LUT3 #(
		.INIT('h54)
	) name3437 (
		\sa20_reg[2]/P0001 ,
		_w690_,
		_w3969_,
		_w3970_
	);
	LUT3 #(
		.INIT('ha8)
	) name3438 (
		\sa20_reg[2]/P0001 ,
		_w696_,
		_w3369_,
		_w3971_
	);
	LUT3 #(
		.INIT('h01)
	) name3439 (
		_w701_,
		_w3384_,
		_w3534_,
		_w3972_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3440 (
		\sa20_reg[1]/P0001 ,
		_w3971_,
		_w3970_,
		_w3972_,
		_w3973_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name3441 (
		\sa20_reg[3]/P0001 ,
		_w666_,
		_w728_,
		_w715_,
		_w3974_
	);
	LUT4 #(
		.INIT('hffa8)
	) name3442 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3975_
	);
	LUT2 #(
		.INIT('h2)
	) name3443 (
		_w735_,
		_w3975_,
		_w3976_
	);
	LUT3 #(
		.INIT('h13)
	) name3444 (
		_w692_,
		_w731_,
		_w3373_,
		_w3977_
	);
	LUT4 #(
		.INIT('h0e00)
	) name3445 (
		\sa20_reg[2]/P0001 ,
		_w3974_,
		_w3976_,
		_w3977_,
		_w3978_
	);
	LUT4 #(
		.INIT('h5455)
	) name3446 (
		\sa20_reg[0]/P0001 ,
		_w3973_,
		_w3967_,
		_w3978_,
		_w3979_
	);
	LUT4 #(
		.INIT('h0013)
	) name3447 (
		_w671_,
		_w653_,
		_w736_,
		_w3364_,
		_w3980_
	);
	LUT4 #(
		.INIT('h47cf)
	) name3448 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w649_,
		_w3383_,
		_w3981_
	);
	LUT4 #(
		.INIT('h0155)
	) name3449 (
		\sa20_reg[1]/P0001 ,
		\sa20_reg[2]/P0001 ,
		_w3980_,
		_w3981_,
		_w3982_
	);
	LUT3 #(
		.INIT('h04)
	) name3450 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w3983_
	);
	LUT4 #(
		.INIT('h3332)
	) name3451 (
		_w682_,
		_w665_,
		_w3384_,
		_w3983_,
		_w3984_
	);
	LUT3 #(
		.INIT('hc8)
	) name3452 (
		_w673_,
		_w739_,
		_w3984_,
		_w3985_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name3453 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3986_
	);
	LUT4 #(
		.INIT('hbf15)
	) name3454 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w693_,
		_w3986_,
		_w3987_
	);
	LUT2 #(
		.INIT('h2)
	) name3455 (
		_w727_,
		_w3987_,
		_w3988_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name3456 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3989_
	);
	LUT2 #(
		.INIT('h2)
	) name3457 (
		_w692_,
		_w3989_,
		_w3990_
	);
	LUT2 #(
		.INIT('h4)
	) name3458 (
		\sa20_reg[1]/P0001 ,
		\sa20_reg[2]/P0001 ,
		_w3991_
	);
	LUT4 #(
		.INIT('h0100)
	) name3459 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w3992_
	);
	LUT4 #(
		.INIT('h0007)
	) name3460 (
		\sa20_reg[7]/NET0131 ,
		_w678_,
		_w731_,
		_w3992_,
		_w3993_
	);
	LUT3 #(
		.INIT('h51)
	) name3461 (
		_w3990_,
		_w3991_,
		_w3993_,
		_w3994_
	);
	LUT4 #(
		.INIT('h0100)
	) name3462 (
		_w3985_,
		_w3988_,
		_w3982_,
		_w3994_,
		_w3995_
	);
	LUT3 #(
		.INIT('h10)
	) name3463 (
		_w3979_,
		_w3962_,
		_w3995_,
		_w3996_
	);
	LUT4 #(
		.INIT('h5655)
	) name3464 (
		\u0_w_reg[2][1]/P0001 ,
		_w3979_,
		_w3962_,
		_w3995_,
		_w3997_
	);
	LUT3 #(
		.INIT('h69)
	) name3465 (
		_w3896_,
		_w3949_,
		_w3997_,
		_w3998_
	);
	LUT3 #(
		.INIT('h28)
	) name3466 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[33]/P0001 ,
		\u0_w_reg[2][1]/P0001 ,
		_w3999_
	);
	LUT4 #(
		.INIT('hff14)
	) name3467 (
		\ld_r_reg/P0001 ,
		_w3842_,
		_w3998_,
		_w3999_,
		_w4000_
	);
	LUT2 #(
		.INIT('h8)
	) name3468 (
		\sa31_reg[3]/P0001 ,
		_w3854_,
		_w4001_
	);
	LUT3 #(
		.INIT('h13)
	) name3469 (
		\sa31_reg[3]/P0001 ,
		_w955_,
		_w3854_,
		_w4002_
	);
	LUT3 #(
		.INIT('h80)
	) name3470 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4003_
	);
	LUT4 #(
		.INIT('hcedf)
	) name3471 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4004_
	);
	LUT3 #(
		.INIT('h8a)
	) name3472 (
		\sa31_reg[2]/P0001 ,
		_w4003_,
		_w4004_,
		_w4005_
	);
	LUT3 #(
		.INIT('ha2)
	) name3473 (
		\sa31_reg[1]/P0001 ,
		_w4002_,
		_w4005_,
		_w4006_
	);
	LUT2 #(
		.INIT('h8)
	) name3474 (
		_w936_,
		_w961_,
		_w4007_
	);
	LUT4 #(
		.INIT('h8880)
	) name3475 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w4008_
	);
	LUT4 #(
		.INIT('h0400)
	) name3476 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4009_
	);
	LUT4 #(
		.INIT('h0023)
	) name3477 (
		_w1003_,
		_w3661_,
		_w4008_,
		_w4009_,
		_w4010_
	);
	LUT3 #(
		.INIT('h45)
	) name3478 (
		\sa31_reg[1]/P0001 ,
		_w4007_,
		_w4010_,
		_w4011_
	);
	LUT4 #(
		.INIT('h5504)
	) name3479 (
		\sa31_reg[3]/P0001 ,
		_w3151_,
		_w3635_,
		_w3906_,
		_w4012_
	);
	LUT4 #(
		.INIT('h0001)
	) name3480 (
		_w1010_,
		_w3661_,
		_w3859_,
		_w3906_,
		_w4013_
	);
	LUT3 #(
		.INIT('h32)
	) name3481 (
		\sa31_reg[2]/P0001 ,
		_w4012_,
		_w4013_,
		_w4014_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3482 (
		\sa31_reg[0]/P0002 ,
		_w4006_,
		_w4011_,
		_w4014_,
		_w4015_
	);
	LUT3 #(
		.INIT('ha8)
	) name3483 (
		\sa31_reg[2]/P0001 ,
		_w993_,
		_w3910_,
		_w4016_
	);
	LUT4 #(
		.INIT('h0800)
	) name3484 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w4017_
	);
	LUT4 #(
		.INIT('h5554)
	) name3485 (
		\sa31_reg[2]/P0001 ,
		_w987_,
		_w3869_,
		_w4017_,
		_w4018_
	);
	LUT4 #(
		.INIT('h0002)
	) name3486 (
		\sa31_reg[1]/P0001 ,
		_w3148_,
		_w3168_,
		_w3169_,
		_w4019_
	);
	LUT3 #(
		.INIT('h10)
	) name3487 (
		_w4018_,
		_w4016_,
		_w4019_,
		_w4020_
	);
	LUT4 #(
		.INIT('h5540)
	) name3488 (
		\sa31_reg[2]/P0001 ,
		_w934_,
		_w936_,
		_w1011_,
		_w4021_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name3489 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4022_
	);
	LUT2 #(
		.INIT('h2)
	) name3490 (
		\sa31_reg[2]/P0001 ,
		_w4022_,
		_w4023_
	);
	LUT2 #(
		.INIT('h8)
	) name3491 (
		\sa31_reg[6]/NET0131 ,
		_w953_,
		_w4024_
	);
	LUT3 #(
		.INIT('h15)
	) name3492 (
		\sa31_reg[1]/P0001 ,
		_w1003_,
		_w3164_,
		_w4025_
	);
	LUT4 #(
		.INIT('h0100)
	) name3493 (
		_w4024_,
		_w4023_,
		_w4021_,
		_w4025_,
		_w4026_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3494 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w4027_
	);
	LUT2 #(
		.INIT('h4)
	) name3495 (
		_w1026_,
		_w4027_,
		_w4028_
	);
	LUT4 #(
		.INIT('h070f)
	) name3496 (
		\sa31_reg[4]/P0001 ,
		_w964_,
		_w1023_,
		_w981_,
		_w4029_
	);
	LUT4 #(
		.INIT('hf400)
	) name3497 (
		_w3180_,
		_w3673_,
		_w4028_,
		_w4029_,
		_w4030_
	);
	LUT4 #(
		.INIT('h0155)
	) name3498 (
		\sa31_reg[0]/P0002 ,
		_w4020_,
		_w4026_,
		_w4030_,
		_w4031_
	);
	LUT4 #(
		.INIT('h0111)
	) name3499 (
		_w946_,
		_w1029_,
		_w1001_,
		_w3182_,
		_w4032_
	);
	LUT3 #(
		.INIT('h9f)
	) name3500 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w948_,
		_w4033_
	);
	LUT4 #(
		.INIT('h0155)
	) name3501 (
		\sa31_reg[1]/P0001 ,
		\sa31_reg[2]/P0001 ,
		_w4032_,
		_w4033_,
		_w4034_
	);
	LUT4 #(
		.INIT('h0100)
	) name3502 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4035_
	);
	LUT4 #(
		.INIT('h0007)
	) name3503 (
		_w969_,
		_w973_,
		_w1023_,
		_w4035_,
		_w4036_
	);
	LUT3 #(
		.INIT('h40)
	) name3504 (
		\sa31_reg[6]/NET0131 ,
		_w981_,
		_w3628_,
		_w4037_
	);
	LUT4 #(
		.INIT('h0031)
	) name3505 (
		_w3885_,
		_w3912_,
		_w4036_,
		_w4037_,
		_w4038_
	);
	LUT3 #(
		.INIT('h01)
	) name3506 (
		_w968_,
		_w3148_,
		_w3863_,
		_w4039_
	);
	LUT2 #(
		.INIT('h1)
	) name3507 (
		_w976_,
		_w3679_,
		_w4040_
	);
	LUT3 #(
		.INIT('h2a)
	) name3508 (
		_w1034_,
		_w4039_,
		_w4040_,
		_w4041_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name3509 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4042_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3510 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w3674_,
		_w4042_,
		_w4043_
	);
	LUT2 #(
		.INIT('h2)
	) name3511 (
		_w1021_,
		_w4043_,
		_w4044_
	);
	LUT4 #(
		.INIT('h0100)
	) name3512 (
		_w4041_,
		_w4044_,
		_w4034_,
		_w4038_,
		_w4045_
	);
	LUT3 #(
		.INIT('h10)
	) name3513 (
		_w4031_,
		_w4015_,
		_w4045_,
		_w4046_
	);
	LUT4 #(
		.INIT('h5655)
	) name3514 (
		\u0_w_reg[2][9]/P0001 ,
		_w4031_,
		_w4015_,
		_w4045_,
		_w4047_
	);
	LUT3 #(
		.INIT('h69)
	) name3515 (
		_w3896_,
		_w3949_,
		_w4047_,
		_w4048_
	);
	LUT4 #(
		.INIT('h0001)
	) name3516 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4049_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name3517 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4050_
	);
	LUT3 #(
		.INIT('h8a)
	) name3518 (
		\sa20_reg[2]/P0001 ,
		_w4049_,
		_w4050_,
		_w4051_
	);
	LUT3 #(
		.INIT('h40)
	) name3519 (
		\sa20_reg[2]/P0001 ,
		_w639_,
		_w704_,
		_w4052_
	);
	LUT3 #(
		.INIT('h02)
	) name3520 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		_w4053_
	);
	LUT3 #(
		.INIT('h01)
	) name3521 (
		_w3370_,
		_w3529_,
		_w4053_,
		_w4054_
	);
	LUT4 #(
		.INIT('h5455)
	) name3522 (
		\sa20_reg[1]/P0001 ,
		_w4052_,
		_w4051_,
		_w4054_,
		_w4055_
	);
	LUT2 #(
		.INIT('h1)
	) name3523 (
		_w653_,
		_w3569_,
		_w4056_
	);
	LUT3 #(
		.INIT('h2a)
	) name3524 (
		\sa20_reg[2]/P0001 ,
		_w3527_,
		_w4056_,
		_w4057_
	);
	LUT3 #(
		.INIT('h51)
	) name3525 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w4058_
	);
	LUT4 #(
		.INIT('h4041)
	) name3526 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4059_
	);
	LUT3 #(
		.INIT('ha8)
	) name3527 (
		\sa20_reg[1]/P0001 ,
		_w721_,
		_w4059_,
		_w4060_
	);
	LUT3 #(
		.INIT('h54)
	) name3528 (
		\sa20_reg[2]/P0001 ,
		_w3355_,
		_w3374_,
		_w4061_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name3529 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4062_
	);
	LUT2 #(
		.INIT('h2)
	) name3530 (
		_w686_,
		_w4062_,
		_w4063_
	);
	LUT3 #(
		.INIT('h0b)
	) name3531 (
		\sa20_reg[5]/P0001 ,
		_w3529_,
		_w3574_,
		_w4064_
	);
	LUT4 #(
		.INIT('h0100)
	) name3532 (
		_w4061_,
		_w4063_,
		_w4060_,
		_w4064_,
		_w4065_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3533 (
		\sa20_reg[0]/P0001 ,
		_w4055_,
		_w4057_,
		_w4065_,
		_w4066_
	);
	LUT4 #(
		.INIT('h8000)
	) name3534 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4067_
	);
	LUT4 #(
		.INIT('h000b)
	) name3535 (
		\sa20_reg[3]/P0001 ,
		_w666_,
		_w711_,
		_w4067_,
		_w4068_
	);
	LUT3 #(
		.INIT('hb9)
	) name3536 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4069_
	);
	LUT3 #(
		.INIT('h08)
	) name3537 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w4070_
	);
	LUT4 #(
		.INIT('h4c00)
	) name3538 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4071_
	);
	LUT4 #(
		.INIT('h45cf)
	) name3539 (
		_w3991_,
		_w4069_,
		_w4070_,
		_w4071_,
		_w4072_
	);
	LUT3 #(
		.INIT('he0)
	) name3540 (
		\sa20_reg[2]/P0001 ,
		_w4068_,
		_w4072_,
		_w4073_
	);
	LUT4 #(
		.INIT('hbf8c)
	) name3541 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		_w729_,
		_w3327_,
		_w4074_
	);
	LUT3 #(
		.INIT('h80)
	) name3542 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w4075_
	);
	LUT4 #(
		.INIT('h0100)
	) name3543 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w4076_
	);
	LUT4 #(
		.INIT('h8007)
	) name3544 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4077_
	);
	LUT4 #(
		.INIT('h0103)
	) name3545 (
		_w700_,
		_w4076_,
		_w4077_,
		_w4075_,
		_w4078_
	);
	LUT3 #(
		.INIT('he4)
	) name3546 (
		\sa20_reg[1]/P0001 ,
		_w4074_,
		_w4078_,
		_w4079_
	);
	LUT3 #(
		.INIT('h15)
	) name3547 (
		\sa20_reg[0]/P0001 ,
		_w4073_,
		_w4079_,
		_w4080_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name3548 (
		_w642_,
		_w662_,
		_w710_,
		_w3345_,
		_w4081_
	);
	LUT2 #(
		.INIT('h1)
	) name3549 (
		\sa20_reg[2]/P0001 ,
		_w4081_,
		_w4082_
	);
	LUT3 #(
		.INIT('h02)
	) name3550 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		_w4083_
	);
	LUT3 #(
		.INIT('h67)
	) name3551 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4084_
	);
	LUT2 #(
		.INIT('h2)
	) name3552 (
		_w4083_,
		_w4084_,
		_w4085_
	);
	LUT3 #(
		.INIT('h15)
	) name3553 (
		\sa20_reg[1]/P0001 ,
		_w673_,
		_w686_,
		_w4086_
	);
	LUT3 #(
		.INIT('h10)
	) name3554 (
		_w3555_,
		_w4085_,
		_w4086_,
		_w4087_
	);
	LUT4 #(
		.INIT('hc480)
	) name3555 (
		\sa20_reg[2]/P0001 ,
		_w671_,
		_w667_,
		_w651_,
		_w4088_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name3556 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w680_,
		_w711_,
		_w4089_
	);
	LUT3 #(
		.INIT('h20)
	) name3557 (
		_w3596_,
		_w4088_,
		_w4089_,
		_w4090_
	);
	LUT4 #(
		.INIT('h0777)
	) name3558 (
		_w668_,
		_w3346_,
		_w3344_,
		_w3574_,
		_w4091_
	);
	LUT4 #(
		.INIT('hf400)
	) name3559 (
		_w4082_,
		_w4087_,
		_w4090_,
		_w4091_,
		_w4092_
	);
	LUT3 #(
		.INIT('h10)
	) name3560 (
		_w4066_,
		_w4080_,
		_w4092_,
		_w4093_
	);
	LUT4 #(
		.INIT('h9669)
	) name3561 (
		_w3389_,
		_w3745_,
		_w3795_,
		_w4093_,
		_w4094_
	);
	LUT3 #(
		.INIT('h28)
	) name3562 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[41]/P0001 ,
		\u0_w_reg[2][9]/P0001 ,
		_w4095_
	);
	LUT4 #(
		.INIT('hff14)
	) name3563 (
		\ld_r_reg/P0001 ,
		_w4048_,
		_w4094_,
		_w4095_,
		_w4096_
	);
	LUT4 #(
		.INIT('h4bb4)
	) name3564 (
		_w775_,
		_w821_,
		_w933_,
		_w3496_,
		_w4097_
	);
	LUT3 #(
		.INIT('h69)
	) name3565 (
		\u0_w_reg[2][5]/P0001 ,
		_w3557_,
		_w3686_,
		_w4098_
	);
	LUT3 #(
		.INIT('h28)
	) name3566 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[37]/P0001 ,
		\u0_w_reg[2][5]/P0001 ,
		_w4099_
	);
	LUT4 #(
		.INIT('hff14)
	) name3567 (
		\ld_r_reg/P0001 ,
		_w4097_,
		_w4098_,
		_w4099_,
		_w4100_
	);
	LUT4 #(
		.INIT('h6996)
	) name3568 (
		\u0_w_reg[2][28]/P0001 ,
		_w3445_,
		_w3616_,
		_w3686_,
		_w4101_
	);
	LUT4 #(
		.INIT('hf3fb)
	) name3569 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w4102_
	);
	LUT3 #(
		.INIT('h8a)
	) name3570 (
		\sa02_reg[2]/P0001 ,
		_w3448_,
		_w4102_,
		_w4103_
	);
	LUT2 #(
		.INIT('h2)
	) name3571 (
		_w900_,
		_w845_,
		_w4104_
	);
	LUT4 #(
		.INIT('h0010)
	) name3572 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w4105_
	);
	LUT3 #(
		.INIT('h01)
	) name3573 (
		_w3097_,
		_w3476_,
		_w4105_,
		_w4106_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3574 (
		\sa02_reg[1]/P0001 ,
		_w4103_,
		_w4104_,
		_w4106_,
		_w4107_
	);
	LUT4 #(
		.INIT('hefdf)
	) name3575 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w4108_
	);
	LUT2 #(
		.INIT('h1)
	) name3576 (
		\sa02_reg[2]/P0001 ,
		_w4108_,
		_w4109_
	);
	LUT4 #(
		.INIT('h0013)
	) name3577 (
		_w869_,
		_w914_,
		_w3090_,
		_w3126_,
		_w4110_
	);
	LUT4 #(
		.INIT('h7077)
	) name3578 (
		_w824_,
		_w828_,
		_w3131_,
		_w3449_,
		_w4111_
	);
	LUT4 #(
		.INIT('h4555)
	) name3579 (
		\sa02_reg[1]/P0001 ,
		_w4109_,
		_w4110_,
		_w4111_,
		_w4112_
	);
	LUT4 #(
		.INIT('h0100)
	) name3580 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w4113_
	);
	LUT4 #(
		.INIT('h0007)
	) name3581 (
		_w856_,
		_w858_,
		_w3816_,
		_w4113_,
		_w4114_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name3582 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w4115_
	);
	LUT4 #(
		.INIT('h7707)
	) name3583 (
		\sa02_reg[5]/P0001 ,
		_w846_,
		_w917_,
		_w4115_,
		_w4116_
	);
	LUT3 #(
		.INIT('he0)
	) name3584 (
		\sa02_reg[2]/P0001 ,
		_w4114_,
		_w4116_,
		_w4117_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3585 (
		\sa02_reg[0]/P0001 ,
		_w4112_,
		_w4107_,
		_w4117_,
		_w4118_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name3586 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w901_,
		_w3112_,
		_w4119_
	);
	LUT2 #(
		.INIT('h4)
	) name3587 (
		\sa02_reg[2]/P0001 ,
		_w881_,
		_w4120_
	);
	LUT4 #(
		.INIT('h006f)
	) name3588 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		_w831_,
		_w3473_,
		_w4121_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3589 (
		\sa02_reg[1]/P0001 ,
		_w4120_,
		_w4119_,
		_w4121_,
		_w4122_
	);
	LUT3 #(
		.INIT('h07)
	) name3590 (
		_w904_,
		_w829_,
		_w4113_,
		_w4123_
	);
	LUT3 #(
		.INIT('h20)
	) name3591 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w4124_
	);
	LUT4 #(
		.INIT('h2237)
	) name3592 (
		_w839_,
		_w841_,
		_w905_,
		_w4124_,
		_w4125_
	);
	LUT3 #(
		.INIT('h15)
	) name3593 (
		\sa02_reg[1]/P0001 ,
		_w4123_,
		_w4125_,
		_w4126_
	);
	LUT4 #(
		.INIT('h5540)
	) name3594 (
		\sa02_reg[2]/P0001 ,
		_w831_,
		_w832_,
		_w911_,
		_w4127_
	);
	LUT2 #(
		.INIT('h8)
	) name3595 (
		_w891_,
		_w901_,
		_w4128_
	);
	LUT4 #(
		.INIT('h45cf)
	) name3596 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		_w862_,
		_w3121_,
		_w4129_
	);
	LUT3 #(
		.INIT('h10)
	) name3597 (
		_w4127_,
		_w4128_,
		_w4129_,
		_w4130_
	);
	LUT4 #(
		.INIT('h5455)
	) name3598 (
		\sa02_reg[0]/P0001 ,
		_w4122_,
		_w4126_,
		_w4130_,
		_w4131_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name3599 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w4132_
	);
	LUT2 #(
		.INIT('h2)
	) name3600 (
		_w3091_,
		_w4132_,
		_w4133_
	);
	LUT3 #(
		.INIT('h40)
	) name3601 (
		\sa02_reg[2]/P0001 ,
		_w837_,
		_w828_,
		_w4134_
	);
	LUT4 #(
		.INIT('h2777)
	) name3602 (
		\sa02_reg[2]/P0001 ,
		_w904_,
		_w837_,
		_w828_,
		_w4135_
	);
	LUT3 #(
		.INIT('h8a)
	) name3603 (
		\sa02_reg[1]/P0001 ,
		_w4133_,
		_w4135_,
		_w4136_
	);
	LUT4 #(
		.INIT('h2000)
	) name3604 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w4137_
	);
	LUT3 #(
		.INIT('ha8)
	) name3605 (
		_w3129_,
		_w3476_,
		_w4137_,
		_w4138_
	);
	LUT4 #(
		.INIT('h8acf)
	) name3606 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w855_,
		_w862_,
		_w4139_
	);
	LUT4 #(
		.INIT('hedff)
	) name3607 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w4140_
	);
	LUT2 #(
		.INIT('h2)
	) name3608 (
		_w891_,
		_w4140_,
		_w4141_
	);
	LUT4 #(
		.INIT('h0777)
	) name3609 (
		_w884_,
		_w3077_,
		_w3466_,
		_w3788_,
		_w4142_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3610 (
		_w3086_,
		_w4139_,
		_w4141_,
		_w4142_,
		_w4143_
	);
	LUT3 #(
		.INIT('h10)
	) name3611 (
		_w4136_,
		_w4138_,
		_w4143_,
		_w4144_
	);
	LUT3 #(
		.INIT('h10)
	) name3612 (
		_w4131_,
		_w4118_,
		_w4144_,
		_w4145_
	);
	LUT4 #(
		.INIT('hefdf)
	) name3613 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4146_
	);
	LUT2 #(
		.INIT('h1)
	) name3614 (
		\sa13_reg[2]/P0001 ,
		_w4146_,
		_w4147_
	);
	LUT3 #(
		.INIT('h8a)
	) name3615 (
		\sa13_reg[2]/P0001 ,
		_w789_,
		_w778_,
		_w4148_
	);
	LUT4 #(
		.INIT('h0007)
	) name3616 (
		_w576_,
		_w553_,
		_w617_,
		_w625_,
		_w4149_
	);
	LUT4 #(
		.INIT('h5455)
	) name3617 (
		\sa13_reg[1]/P0001 ,
		_w4148_,
		_w4147_,
		_w4149_,
		_w4150_
	);
	LUT4 #(
		.INIT('hf3fb)
	) name3618 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4151_
	);
	LUT3 #(
		.INIT('h8a)
	) name3619 (
		\sa13_reg[2]/P0001 ,
		_w3302_,
		_w4151_,
		_w4152_
	);
	LUT2 #(
		.INIT('h1)
	) name3620 (
		_w563_,
		_w3286_,
		_w4153_
	);
	LUT3 #(
		.INIT('h01)
	) name3621 (
		_w3320_,
		_w3409_,
		_w3741_,
		_w4154_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3622 (
		\sa13_reg[1]/P0001 ,
		_w4152_,
		_w4153_,
		_w4154_,
		_w4155_
	);
	LUT4 #(
		.INIT('h8000)
	) name3623 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4156_
	);
	LUT4 #(
		.INIT('h0007)
	) name3624 (
		_w562_,
		_w784_,
		_w3281_,
		_w4156_,
		_w4157_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name3625 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4158_
	);
	LUT4 #(
		.INIT('h7707)
	) name3626 (
		\sa13_reg[3]/P0001 ,
		_w569_,
		_w3739_,
		_w4158_,
		_w4159_
	);
	LUT3 #(
		.INIT('he0)
	) name3627 (
		\sa13_reg[2]/P0001 ,
		_w4157_,
		_w4159_,
		_w4160_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3628 (
		\sa13_reg[0]/P0001 ,
		_w4150_,
		_w4155_,
		_w4160_,
		_w4161_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3629 (
		\sa13_reg[2]/P0001 ,
		_w567_,
		_w584_,
		_w607_,
		_w4162_
	);
	LUT3 #(
		.INIT('h13)
	) name3630 (
		\sa13_reg[7]/NET0131 ,
		_w579_,
		_w625_,
		_w4163_
	);
	LUT4 #(
		.INIT('h153f)
	) name3631 (
		_w561_,
		_w571_,
		_w542_,
		_w3300_,
		_w4164_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3632 (
		\sa13_reg[1]/P0001 ,
		_w4162_,
		_w4163_,
		_w4164_,
		_w4165_
	);
	LUT4 #(
		.INIT('h0008)
	) name3633 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4166_
	);
	LUT3 #(
		.INIT('h01)
	) name3634 (
		_w615_,
		_w3281_,
		_w4166_,
		_w4167_
	);
	LUT3 #(
		.INIT('he0)
	) name3635 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4168_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name3636 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w563_,
		_w4168_,
		_w4169_
	);
	LUT3 #(
		.INIT('h15)
	) name3637 (
		\sa13_reg[1]/P0001 ,
		_w4167_,
		_w4169_,
		_w4170_
	);
	LUT4 #(
		.INIT('h4440)
	) name3638 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w572_,
		_w573_,
		_w4171_
	);
	LUT2 #(
		.INIT('h8)
	) name3639 (
		_w554_,
		_w616_,
		_w4172_
	);
	LUT4 #(
		.INIT('h153f)
	) name3640 (
		_w571_,
		_w584_,
		_w594_,
		_w628_,
		_w4173_
	);
	LUT3 #(
		.INIT('h10)
	) name3641 (
		_w4171_,
		_w4172_,
		_w4173_,
		_w4174_
	);
	LUT4 #(
		.INIT('h5455)
	) name3642 (
		\sa13_reg[0]/P0001 ,
		_w4165_,
		_w4170_,
		_w4174_,
		_w4175_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name3643 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4176_
	);
	LUT2 #(
		.INIT('h2)
	) name3644 (
		_w3285_,
		_w4176_,
		_w4177_
	);
	LUT4 #(
		.INIT('h2777)
	) name3645 (
		\sa13_reg[2]/P0001 ,
		_w563_,
		_w814_,
		_w3267_,
		_w4178_
	);
	LUT3 #(
		.INIT('h8a)
	) name3646 (
		\sa13_reg[1]/P0001 ,
		_w4177_,
		_w4178_,
		_w4179_
	);
	LUT4 #(
		.INIT('haaef)
	) name3647 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w554_,
		_w615_,
		_w4180_
	);
	LUT2 #(
		.INIT('h2)
	) name3648 (
		_w3733_,
		_w4180_,
		_w4181_
	);
	LUT4 #(
		.INIT('h2000)
	) name3649 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w4182_
	);
	LUT3 #(
		.INIT('hc8)
	) name3650 (
		_w3409_,
		_w3729_,
		_w4182_,
		_w4183_
	);
	LUT2 #(
		.INIT('h8)
	) name3651 (
		_w809_,
		_w3396_,
		_w4184_
	);
	LUT2 #(
		.INIT('h8)
	) name3652 (
		_w534_,
		_w594_,
		_w4185_
	);
	LUT4 #(
		.INIT('h337f)
	) name3653 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w579_,
		_w619_,
		_w4186_
	);
	LUT4 #(
		.INIT('h0100)
	) name3654 (
		_w4185_,
		_w4183_,
		_w4184_,
		_w4186_,
		_w4187_
	);
	LUT3 #(
		.INIT('h10)
	) name3655 (
		_w4179_,
		_w4181_,
		_w4187_,
		_w4188_
	);
	LUT3 #(
		.INIT('h10)
	) name3656 (
		_w4175_,
		_w4161_,
		_w4188_,
		_w4189_
	);
	LUT4 #(
		.INIT('h9669)
	) name3657 (
		_w3265_,
		_w3324_,
		_w4145_,
		_w4189_,
		_w4190_
	);
	LUT3 #(
		.INIT('h82)
	) name3658 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[60]/P0001 ,
		\u0_w_reg[2][28]/P0001 ,
		_w4191_
	);
	LUT4 #(
		.INIT('h00be)
	) name3659 (
		\ld_r_reg/P0001 ,
		_w4101_,
		_w4190_,
		_w4191_,
		_w4192_
	);
	LUT4 #(
		.INIT('h5400)
	) name3660 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4193_
	);
	LUT3 #(
		.INIT('ha8)
	) name3661 (
		\sa20_reg[2]/P0001 ,
		_w729_,
		_w4193_,
		_w4194_
	);
	LUT4 #(
		.INIT('h0007)
	) name3662 (
		_w666_,
		_w686_,
		_w730_,
		_w3341_,
		_w4195_
	);
	LUT3 #(
		.INIT('h45)
	) name3663 (
		\sa20_reg[1]/P0001 ,
		_w4194_,
		_w4195_,
		_w4196_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3664 (
		\sa20_reg[2]/P0001 ,
		_w677_,
		_w697_,
		_w707_,
		_w4197_
	);
	LUT3 #(
		.INIT('h15)
	) name3665 (
		_w680_,
		_w710_,
		_w3510_,
		_w4198_
	);
	LUT4 #(
		.INIT('h23af)
	) name3666 (
		\sa20_reg[2]/P0001 ,
		_w647_,
		_w644_,
		_w3510_,
		_w4199_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3667 (
		\sa20_reg[1]/P0001 ,
		_w4197_,
		_w4198_,
		_w4199_,
		_w4200_
	);
	LUT4 #(
		.INIT('h0105)
	) name3668 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w676_,
		_w678_,
		_w4201_
	);
	LUT4 #(
		.INIT('h0002)
	) name3669 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w4202_
	);
	LUT3 #(
		.INIT('h02)
	) name3670 (
		\sa20_reg[2]/P0001 ,
		_w716_,
		_w4202_,
		_w4203_
	);
	LUT3 #(
		.INIT('h54)
	) name3671 (
		_w3537_,
		_w4201_,
		_w4203_,
		_w4204_
	);
	LUT4 #(
		.INIT('h5455)
	) name3672 (
		\sa20_reg[0]/P0001 ,
		_w4200_,
		_w4196_,
		_w4204_,
		_w4205_
	);
	LUT4 #(
		.INIT('hffac)
	) name3673 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4206_
	);
	LUT2 #(
		.INIT('h1)
	) name3674 (
		\sa20_reg[2]/P0001 ,
		_w4206_,
		_w4207_
	);
	LUT3 #(
		.INIT('h01)
	) name3675 (
		_w666_,
		_w708_,
		_w3381_,
		_w4208_
	);
	LUT3 #(
		.INIT('h8a)
	) name3676 (
		\sa20_reg[1]/P0001 ,
		_w4207_,
		_w4208_,
		_w4209_
	);
	LUT4 #(
		.INIT('h000b)
	) name3677 (
		\sa20_reg[3]/P0001 ,
		_w666_,
		_w3341_,
		_w4067_,
		_w4210_
	);
	LUT3 #(
		.INIT('h32)
	) name3678 (
		\sa20_reg[2]/P0001 ,
		_w3540_,
		_w4210_,
		_w4211_
	);
	LUT4 #(
		.INIT('hefdf)
	) name3679 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4212_
	);
	LUT2 #(
		.INIT('h1)
	) name3680 (
		\sa20_reg[2]/P0001 ,
		_w4212_,
		_w4213_
	);
	LUT4 #(
		.INIT('h0103)
	) name3681 (
		_w665_,
		_w731_,
		_w723_,
		_w3383_,
		_w4214_
	);
	LUT3 #(
		.INIT('h3b)
	) name3682 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w4215_
	);
	LUT4 #(
		.INIT('h5f5d)
	) name3683 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w680_,
		_w4215_,
		_w4216_
	);
	LUT4 #(
		.INIT('h4555)
	) name3684 (
		\sa20_reg[1]/P0001 ,
		_w4213_,
		_w4214_,
		_w4216_,
		_w4217_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name3685 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4218_
	);
	LUT2 #(
		.INIT('h2)
	) name3686 (
		\sa20_reg[4]/P0001 ,
		_w4218_,
		_w4219_
	);
	LUT4 #(
		.INIT('hd1ff)
	) name3687 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4220_
	);
	LUT3 #(
		.INIT('h8a)
	) name3688 (
		\sa20_reg[1]/P0001 ,
		_w3983_,
		_w4220_,
		_w4221_
	);
	LUT3 #(
		.INIT('ha8)
	) name3689 (
		\sa20_reg[2]/P0001 ,
		_w4219_,
		_w4221_,
		_w4222_
	);
	LUT4 #(
		.INIT('h0100)
	) name3690 (
		_w4209_,
		_w4217_,
		_w4222_,
		_w4211_,
		_w4223_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name3691 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4224_
	);
	LUT2 #(
		.INIT('h2)
	) name3692 (
		_w654_,
		_w4224_,
		_w4225_
	);
	LUT3 #(
		.INIT('h8b)
	) name3693 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w4226_
	);
	LUT2 #(
		.INIT('h2)
	) name3694 (
		_w4075_,
		_w4226_,
		_w4227_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name3695 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		_w666_,
		_w3569_,
		_w4228_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3696 (
		\sa20_reg[1]/P0001 ,
		_w4227_,
		_w4225_,
		_w4228_,
		_w4229_
	);
	LUT3 #(
		.INIT('h2a)
	) name3697 (
		\sa20_reg[2]/P0001 ,
		_w667_,
		_w710_,
		_w4230_
	);
	LUT3 #(
		.INIT('h54)
	) name3698 (
		\sa20_reg[1]/P0001 ,
		\sa20_reg[2]/P0001 ,
		_w3600_,
		_w4231_
	);
	LUT4 #(
		.INIT('hedff)
	) name3699 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4232_
	);
	LUT4 #(
		.INIT('h7707)
	) name3700 (
		_w647_,
		_w667_,
		_w692_,
		_w4232_,
		_w4233_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3701 (
		_w3528_,
		_w4230_,
		_w4231_,
		_w4233_,
		_w4234_
	);
	LUT2 #(
		.INIT('h4)
	) name3702 (
		_w4229_,
		_w4234_,
		_w4235_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3703 (
		\sa20_reg[0]/P0001 ,
		_w4223_,
		_w4205_,
		_w4235_,
		_w4236_
	);
	LUT4 #(
		.INIT('h6996)
	) name3704 (
		_w3324_,
		_w3496_,
		_w4189_,
		_w4236_,
		_w4237_
	);
	LUT4 #(
		.INIT('h9669)
	) name3705 (
		\u0_w_reg[2][20]/P0001 ,
		_w3389_,
		_w3616_,
		_w3686_,
		_w4238_
	);
	LUT3 #(
		.INIT('h82)
	) name3706 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[52]/P0001 ,
		\u0_w_reg[2][20]/P0001 ,
		_w4239_
	);
	LUT4 #(
		.INIT('h00be)
	) name3707 (
		\ld_r_reg/P0001 ,
		_w4237_,
		_w4238_,
		_w4239_,
		_w4240_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3708 (
		\sa31_reg[2]/P0001 ,
		_w947_,
		_w975_,
		_w985_,
		_w4241_
	);
	LUT2 #(
		.INIT('h8)
	) name3709 (
		_w938_,
		_w3635_,
		_w4242_
	);
	LUT3 #(
		.INIT('h13)
	) name3710 (
		\sa31_reg[7]/P0001 ,
		_w977_,
		_w1018_,
		_w4243_
	);
	LUT4 #(
		.INIT('h0100)
	) name3711 (
		_w4001_,
		_w4242_,
		_w4241_,
		_w4243_,
		_w4244_
	);
	LUT3 #(
		.INIT('he0)
	) name3712 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4245_
	);
	LUT2 #(
		.INIT('h8)
	) name3713 (
		_w992_,
		_w4245_,
		_w4246_
	);
	LUT4 #(
		.INIT('h0100)
	) name3714 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w4247_
	);
	LUT4 #(
		.INIT('h0008)
	) name3715 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4248_
	);
	LUT3 #(
		.INIT('h01)
	) name3716 (
		_w1022_,
		_w4247_,
		_w4248_,
		_w4249_
	);
	LUT3 #(
		.INIT('h10)
	) name3717 (
		_w1033_,
		_w4246_,
		_w4249_,
		_w4250_
	);
	LUT4 #(
		.INIT('h5450)
	) name3718 (
		\sa31_reg[2]/P0001 ,
		_w969_,
		_w972_,
		_w973_,
		_w4251_
	);
	LUT2 #(
		.INIT('h8)
	) name3719 (
		_w975_,
		_w981_,
		_w4252_
	);
	LUT4 #(
		.INIT('h135f)
	) name3720 (
		_w934_,
		_w973_,
		_w1030_,
		_w1014_,
		_w4253_
	);
	LUT3 #(
		.INIT('h10)
	) name3721 (
		_w4251_,
		_w4252_,
		_w4253_,
		_w4254_
	);
	LUT4 #(
		.INIT('hd800)
	) name3722 (
		\sa31_reg[1]/P0001 ,
		_w4244_,
		_w4250_,
		_w4254_,
		_w4255_
	);
	LUT4 #(
		.INIT('hff3b)
	) name3723 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4256_
	);
	LUT3 #(
		.INIT('h8a)
	) name3724 (
		\sa31_reg[2]/P0001 ,
		_w977_,
		_w4256_,
		_w4257_
	);
	LUT4 #(
		.INIT('hefdf)
	) name3725 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4258_
	);
	LUT2 #(
		.INIT('h1)
	) name3726 (
		\sa31_reg[2]/P0001 ,
		_w4258_,
		_w4259_
	);
	LUT4 #(
		.INIT('h0007)
	) name3727 (
		_w948_,
		_w954_,
		_w1023_,
		_w1018_,
		_w4260_
	);
	LUT4 #(
		.INIT('h5455)
	) name3728 (
		\sa31_reg[1]/P0001 ,
		_w4259_,
		_w4257_,
		_w4260_,
		_w4261_
	);
	LUT4 #(
		.INIT('hffac)
	) name3729 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4262_
	);
	LUT2 #(
		.INIT('h1)
	) name3730 (
		\sa31_reg[2]/P0001 ,
		_w4262_,
		_w4263_
	);
	LUT4 #(
		.INIT('h0c04)
	) name3731 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4264_
	);
	LUT3 #(
		.INIT('ha8)
	) name3732 (
		\sa31_reg[2]/P0001 ,
		_w3628_,
		_w4264_,
		_w4265_
	);
	LUT3 #(
		.INIT('h13)
	) name3733 (
		\sa31_reg[4]/P0001 ,
		_w3625_,
		_w3886_,
		_w4266_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3734 (
		\sa31_reg[1]/P0001 ,
		_w4265_,
		_w4263_,
		_w4266_,
		_w4267_
	);
	LUT4 #(
		.INIT('h0007)
	) name3735 (
		\sa31_reg[7]/P0001 ,
		_w970_,
		_w3875_,
		_w4247_,
		_w4268_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name3736 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4269_
	);
	LUT4 #(
		.INIT('h5f13)
	) name3737 (
		_w940_,
		_w1028_,
		_w3164_,
		_w4269_,
		_w4270_
	);
	LUT3 #(
		.INIT('he0)
	) name3738 (
		\sa31_reg[2]/P0001 ,
		_w4268_,
		_w4270_,
		_w4271_
	);
	LUT3 #(
		.INIT('h10)
	) name3739 (
		_w4261_,
		_w4267_,
		_w4271_,
		_w4272_
	);
	LUT4 #(
		.INIT('h2000)
	) name3740 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w4273_
	);
	LUT3 #(
		.INIT('ha8)
	) name3741 (
		\sa31_reg[2]/P0001 ,
		_w3625_,
		_w4273_,
		_w4274_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name3742 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4275_
	);
	LUT2 #(
		.INIT('h2)
	) name3743 (
		_w949_,
		_w4275_,
		_w4276_
	);
	LUT3 #(
		.INIT('h40)
	) name3744 (
		\sa31_reg[6]/NET0131 ,
		_w3176_,
		_w3928_,
		_w4277_
	);
	LUT4 #(
		.INIT('h0001)
	) name3745 (
		_w3639_,
		_w4276_,
		_w4274_,
		_w4277_,
		_w4278_
	);
	LUT4 #(
		.INIT('hffed)
	) name3746 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4279_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3747 (
		_w992_,
		_w3635_,
		_w4003_,
		_w4279_,
		_w4280_
	);
	LUT4 #(
		.INIT('hedff)
	) name3748 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4281_
	);
	LUT4 #(
		.INIT('h7707)
	) name3749 (
		\sa31_reg[6]/NET0131 ,
		_w953_,
		_w981_,
		_w4281_,
		_w4282_
	);
	LUT3 #(
		.INIT('he0)
	) name3750 (
		\sa31_reg[1]/P0001 ,
		_w4280_,
		_w4282_,
		_w4283_
	);
	LUT3 #(
		.INIT('hd0)
	) name3751 (
		\sa31_reg[1]/P0001 ,
		_w4278_,
		_w4283_,
		_w4284_
	);
	LUT4 #(
		.INIT('hd800)
	) name3752 (
		\sa31_reg[0]/P0002 ,
		_w4272_,
		_w4255_,
		_w4284_,
		_w4285_
	);
	LUT4 #(
		.INIT('h9669)
	) name3753 (
		\u0_w_reg[2][12]/P0001 ,
		_w3686_,
		_w3949_,
		_w4285_,
		_w4286_
	);
	LUT4 #(
		.INIT('h9669)
	) name3754 (
		_w3389_,
		_w3445_,
		_w3496_,
		_w4236_,
		_w4287_
	);
	LUT3 #(
		.INIT('h82)
	) name3755 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[44]/P0001 ,
		\u0_w_reg[2][12]/P0001 ,
		_w4288_
	);
	LUT4 #(
		.INIT('h00eb)
	) name3756 (
		\ld_r_reg/P0001 ,
		_w4286_,
		_w4287_,
		_w4288_,
		_w4289_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3757 (
		\sa13_reg[2]/P0001 ,
		_w620_,
		_w754_,
		_w798_,
		_w4290_
	);
	LUT3 #(
		.INIT('h80)
	) name3758 (
		\sa13_reg[4]/P0001 ,
		_w537_,
		_w548_,
		_w4291_
	);
	LUT3 #(
		.INIT('h8a)
	) name3759 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4292_
	);
	LUT4 #(
		.INIT('h0010)
	) name3760 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w4293_
	);
	LUT3 #(
		.INIT('h0d)
	) name3761 (
		_w613_,
		_w4292_,
		_w4293_,
		_w4294_
	);
	LUT4 #(
		.INIT('h5455)
	) name3762 (
		\sa13_reg[1]/P0001 ,
		_w4291_,
		_w4290_,
		_w4294_,
		_w4295_
	);
	LUT4 #(
		.INIT('h4041)
	) name3763 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4296_
	);
	LUT3 #(
		.INIT('ha8)
	) name3764 (
		\sa13_reg[1]/P0001 ,
		_w623_,
		_w4296_,
		_w4297_
	);
	LUT3 #(
		.INIT('h07)
	) name3765 (
		_w562_,
		_w784_,
		_w3413_,
		_w4298_
	);
	LUT3 #(
		.INIT('h2a)
	) name3766 (
		\sa13_reg[2]/P0001 ,
		_w546_,
		_w4298_,
		_w4299_
	);
	LUT3 #(
		.INIT('h54)
	) name3767 (
		\sa13_reg[2]/P0001 ,
		_w794_,
		_w3292_,
		_w4300_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name3768 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4301_
	);
	LUT2 #(
		.INIT('h2)
	) name3769 (
		_w558_,
		_w4301_,
		_w4302_
	);
	LUT3 #(
		.INIT('h15)
	) name3770 (
		_w748_,
		_w814_,
		_w3267_,
		_w4303_
	);
	LUT3 #(
		.INIT('h10)
	) name3771 (
		_w4300_,
		_w4302_,
		_w4303_,
		_w4304_
	);
	LUT4 #(
		.INIT('h0100)
	) name3772 (
		_w4295_,
		_w4299_,
		_w4297_,
		_w4304_,
		_w4305_
	);
	LUT4 #(
		.INIT('h0100)
	) name3773 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w4306_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3774 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[3]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4307_
	);
	LUT2 #(
		.INIT('h4)
	) name3775 (
		_w4306_,
		_w4307_,
		_w4308_
	);
	LUT4 #(
		.INIT('h8003)
	) name3776 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4309_
	);
	LUT3 #(
		.INIT('h07)
	) name3777 (
		_w594_,
		_w747_,
		_w4309_,
		_w4310_
	);
	LUT2 #(
		.INIT('h1)
	) name3778 (
		\sa13_reg[3]/P0001 ,
		_w3266_,
		_w4311_
	);
	LUT3 #(
		.INIT('h15)
	) name3779 (
		\sa13_reg[1]/P0001 ,
		_w589_,
		_w804_,
		_w4312_
	);
	LUT4 #(
		.INIT('h7077)
	) name3780 (
		_w4308_,
		_w4310_,
		_w4311_,
		_w4312_,
		_w4313_
	);
	LUT4 #(
		.INIT('h0013)
	) name3781 (
		_w562_,
		_w609_,
		_w784_,
		_w4156_,
		_w4314_
	);
	LUT3 #(
		.INIT('hb9)
	) name3782 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4315_
	);
	LUT4 #(
		.INIT('hb3ff)
	) name3783 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4316_
	);
	LUT4 #(
		.INIT('hf531)
	) name3784 (
		_w761_,
		_w3733_,
		_w4315_,
		_w4316_,
		_w4317_
	);
	LUT3 #(
		.INIT('he0)
	) name3785 (
		\sa13_reg[2]/P0001 ,
		_w4314_,
		_w4317_,
		_w4318_
	);
	LUT2 #(
		.INIT('h4)
	) name3786 (
		_w4313_,
		_w4318_,
		_w4319_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3787 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w579_,
		_w768_,
		_w4320_
	);
	LUT4 #(
		.INIT('h8acf)
	) name3788 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[5]/P0001 ,
		_w617_,
		_w3320_,
		_w4321_
	);
	LUT3 #(
		.INIT('h20)
	) name3789 (
		_w3402_,
		_w4320_,
		_w4321_,
		_w4322_
	);
	LUT3 #(
		.INIT('h07)
	) name3790 (
		\sa13_reg[3]/P0001 ,
		_w569_,
		_w768_,
		_w4323_
	);
	LUT3 #(
		.INIT('h07)
	) name3791 (
		_w543_,
		_w616_,
		_w3283_,
		_w4324_
	);
	LUT4 #(
		.INIT('h1555)
	) name3792 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w543_,
		_w594_,
		_w4325_
	);
	LUT4 #(
		.INIT('hea00)
	) name3793 (
		\sa13_reg[2]/P0001 ,
		_w4323_,
		_w4324_,
		_w4325_,
		_w4326_
	);
	LUT4 #(
		.INIT('hdc00)
	) name3794 (
		\sa13_reg[3]/P0001 ,
		_w625_,
		_w3413_,
		_w3733_,
		_w4327_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3795 (
		\sa13_reg[6]/NET0131 ,
		_w583_,
		_w596_,
		_w789_,
		_w4328_
	);
	LUT2 #(
		.INIT('h1)
	) name3796 (
		_w4327_,
		_w4328_,
		_w4329_
	);
	LUT3 #(
		.INIT('he0)
	) name3797 (
		_w4322_,
		_w4326_,
		_w4329_,
		_w4330_
	);
	LUT4 #(
		.INIT('hd800)
	) name3798 (
		\sa13_reg[0]/P0001 ,
		_w4305_,
		_w4319_,
		_w4330_,
		_w4331_
	);
	LUT4 #(
		.INIT('h6996)
	) name3799 (
		_w3324_,
		_w3795_,
		_w4093_,
		_w4331_,
		_w4332_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name3800 (
		\u0_w_reg[2][17]/P0001 ,
		_w4031_,
		_w4015_,
		_w4045_,
		_w4333_
	);
	LUT3 #(
		.INIT('h69)
	) name3801 (
		_w3389_,
		_w3996_,
		_w4333_,
		_w4334_
	);
	LUT3 #(
		.INIT('h28)
	) name3802 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[49]/P0001 ,
		\u0_w_reg[2][17]/P0001 ,
		_w4335_
	);
	LUT4 #(
		.INIT('hff14)
	) name3803 (
		\ld_r_reg/P0001 ,
		_w4332_,
		_w4334_,
		_w4335_,
		_w4336_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name3804 (
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4337_
	);
	LUT4 #(
		.INIT('h0002)
	) name3805 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4338_
	);
	LUT4 #(
		.INIT('h0b01)
	) name3806 (
		\sa13_reg[3]/P0001 ,
		_w747_,
		_w4338_,
		_w4337_,
		_w4339_
	);
	LUT2 #(
		.INIT('h2)
	) name3807 (
		\sa13_reg[2]/P0001 ,
		_w4339_,
		_w4340_
	);
	LUT3 #(
		.INIT('h01)
	) name3808 (
		_w551_,
		_w3396_,
		_w3415_,
		_w4341_
	);
	LUT3 #(
		.INIT('h54)
	) name3809 (
		\sa13_reg[2]/P0001 ,
		_w617_,
		_w798_,
		_w4342_
	);
	LUT4 #(
		.INIT('h0020)
	) name3810 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4343_
	);
	LUT3 #(
		.INIT('h01)
	) name3811 (
		_w3403_,
		_w4293_,
		_w4343_,
		_w4344_
	);
	LUT4 #(
		.INIT('h4555)
	) name3812 (
		\sa13_reg[1]/P0001 ,
		_w4342_,
		_w4344_,
		_w4341_,
		_w4345_
	);
	LUT4 #(
		.INIT('hbbf3)
	) name3813 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w4346_
	);
	LUT4 #(
		.INIT('h80f0)
	) name3814 (
		\sa13_reg[3]/P0001 ,
		_w569_,
		_w632_,
		_w4346_,
		_w4347_
	);
	LUT4 #(
		.INIT('haaef)
	) name3815 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		_w543_,
		_w3413_,
		_w4348_
	);
	LUT2 #(
		.INIT('h4)
	) name3816 (
		_w4347_,
		_w4348_,
		_w4349_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3817 (
		\sa13_reg[0]/P0001 ,
		_w4345_,
		_w4340_,
		_w4349_,
		_w4350_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3818 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4351_
	);
	LUT4 #(
		.INIT('h5554)
	) name3819 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w4352_
	);
	LUT4 #(
		.INIT('h5fdf)
	) name3820 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4353_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name3821 (
		_w790_,
		_w4351_,
		_w4352_,
		_w4353_,
		_w4354_
	);
	LUT3 #(
		.INIT('ha8)
	) name3822 (
		\sa13_reg[1]/P0001 ,
		_w3297_,
		_w4354_,
		_w4355_
	);
	LUT3 #(
		.INIT('h04)
	) name3823 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w4356_
	);
	LUT3 #(
		.INIT('ha8)
	) name3824 (
		_w558_,
		_w3271_,
		_w4356_,
		_w4357_
	);
	LUT2 #(
		.INIT('h4)
	) name3825 (
		\sa13_reg[1]/P0001 ,
		_w3320_,
		_w4358_
	);
	LUT3 #(
		.INIT('h15)
	) name3826 (
		_w563_,
		_w3409_,
		_w3739_,
		_w4359_
	);
	LUT3 #(
		.INIT('h10)
	) name3827 (
		_w4357_,
		_w4358_,
		_w4359_,
		_w4360_
	);
	LUT3 #(
		.INIT('h45)
	) name3828 (
		\sa13_reg[0]/P0001 ,
		_w4355_,
		_w4360_,
		_w4361_
	);
	LUT4 #(
		.INIT('h0007)
	) name3829 (
		_w535_,
		_w591_,
		_w626_,
		_w3271_,
		_w4362_
	);
	LUT4 #(
		.INIT('haaa2)
	) name3830 (
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		_w4363_
	);
	LUT4 #(
		.INIT('h1300)
	) name3831 (
		\sa13_reg[5]/P0001 ,
		_w3320_,
		_w3396_,
		_w4363_,
		_w4364_
	);
	LUT3 #(
		.INIT('hb8)
	) name3832 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[7]/NET0131 ,
		_w4365_
	);
	LUT2 #(
		.INIT('h8)
	) name3833 (
		_w576_,
		_w4365_,
		_w4366_
	);
	LUT4 #(
		.INIT('h00f8)
	) name3834 (
		_w552_,
		_w4362_,
		_w4364_,
		_w4366_,
		_w4367_
	);
	LUT4 #(
		.INIT('h0400)
	) name3835 (
		\sa13_reg[3]/P0001 ,
		\sa13_reg[4]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4368_
	);
	LUT4 #(
		.INIT('h0007)
	) name3836 (
		_w571_,
		_w542_,
		_w534_,
		_w4368_,
		_w4369_
	);
	LUT3 #(
		.INIT('h32)
	) name3837 (
		\sa13_reg[2]/P0001 ,
		_w751_,
		_w4369_,
		_w4370_
	);
	LUT3 #(
		.INIT('had)
	) name3838 (
		\sa13_reg[5]/P0001 ,
		\sa13_reg[6]/NET0131 ,
		\sa13_reg[7]/NET0131 ,
		_w4371_
	);
	LUT2 #(
		.INIT('h2)
	) name3839 (
		_w616_,
		_w4371_,
		_w4372_
	);
	LUT3 #(
		.INIT('ha8)
	) name3840 (
		\sa13_reg[1]/P0001 ,
		_w798_,
		_w3720_,
		_w4373_
	);
	LUT3 #(
		.INIT('h80)
	) name3841 (
		\sa13_reg[1]/P0001 ,
		\sa13_reg[2]/P0001 ,
		\sa13_reg[3]/P0001 ,
		_w4374_
	);
	LUT4 #(
		.INIT('h153f)
	) name3842 (
		_w795_,
		_w814_,
		_w3300_,
		_w4374_,
		_w4375_
	);
	LUT4 #(
		.INIT('h5700)
	) name3843 (
		\sa13_reg[2]/P0001 ,
		_w4372_,
		_w4373_,
		_w4375_,
		_w4376_
	);
	LUT4 #(
		.INIT('he400)
	) name3844 (
		\sa13_reg[1]/P0001 ,
		_w4367_,
		_w4370_,
		_w4376_,
		_w4377_
	);
	LUT3 #(
		.INIT('h10)
	) name3845 (
		_w4350_,
		_w4361_,
		_w4377_,
		_w4378_
	);
	LUT3 #(
		.INIT('h01)
	) name3846 (
		_w3073_,
		_w3450_,
		_w3491_,
		_w4379_
	);
	LUT3 #(
		.INIT('h54)
	) name3847 (
		\sa02_reg[2]/P0001 ,
		_w864_,
		_w914_,
		_w4380_
	);
	LUT3 #(
		.INIT('h01)
	) name3848 (
		_w927_,
		_w3463_,
		_w3466_,
		_w4381_
	);
	LUT4 #(
		.INIT('h4555)
	) name3849 (
		\sa02_reg[1]/P0001 ,
		_w4380_,
		_w4381_,
		_w4379_,
		_w4382_
	);
	LUT4 #(
		.INIT('h440c)
	) name3850 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w4383_
	);
	LUT4 #(
		.INIT('h5540)
	) name3851 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		_w846_,
		_w4383_,
		_w4384_
	);
	LUT3 #(
		.INIT('ha8)
	) name3852 (
		\sa02_reg[1]/P0001 ,
		_w3124_,
		_w4384_,
		_w4385_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name3853 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w4386_
	);
	LUT2 #(
		.INIT('h2)
	) name3854 (
		_w891_,
		_w4386_,
		_w4387_
	);
	LUT4 #(
		.INIT('hfefb)
	) name3855 (
		\sa02_reg[4]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w4388_
	);
	LUT3 #(
		.INIT('h45)
	) name3856 (
		\sa02_reg[3]/P0001 ,
		_w3450_,
		_w4388_,
		_w4389_
	);
	LUT2 #(
		.INIT('h1)
	) name3857 (
		_w4387_,
		_w4389_,
		_w4390_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3858 (
		\sa02_reg[0]/P0001 ,
		_w4385_,
		_w4382_,
		_w4390_,
		_w4391_
	);
	LUT3 #(
		.INIT('h01)
	) name3859 (
		\sa02_reg[2]/P0001 ,
		_w3073_,
		_w3125_,
		_w4392_
	);
	LUT3 #(
		.INIT('h07)
	) name3860 (
		\sa02_reg[6]/NET0131 ,
		_w852_,
		_w3213_,
		_w4393_
	);
	LUT4 #(
		.INIT('haaa2)
	) name3861 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w4394_
	);
	LUT4 #(
		.INIT('h0700)
	) name3862 (
		_w861_,
		_w875_,
		_w3261_,
		_w4394_,
		_w4395_
	);
	LUT3 #(
		.INIT('h0b)
	) name3863 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		_w4396_
	);
	LUT3 #(
		.INIT('h15)
	) name3864 (
		\sa02_reg[1]/P0001 ,
		_w3747_,
		_w4396_,
		_w4397_
	);
	LUT4 #(
		.INIT('hf800)
	) name3865 (
		_w4392_,
		_w4393_,
		_w4395_,
		_w4397_,
		_w4398_
	);
	LUT4 #(
		.INIT('h0400)
	) name3866 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w4399_
	);
	LUT4 #(
		.INIT('h0013)
	) name3867 (
		_w831_,
		_w895_,
		_w824_,
		_w4399_,
		_w4400_
	);
	LUT2 #(
		.INIT('h2)
	) name3868 (
		\sa02_reg[1]/P0001 ,
		_w883_,
		_w4401_
	);
	LUT3 #(
		.INIT('he0)
	) name3869 (
		\sa02_reg[2]/P0001 ,
		_w4400_,
		_w4401_,
		_w4402_
	);
	LUT2 #(
		.INIT('h1)
	) name3870 (
		_w4398_,
		_w4402_,
		_w4403_
	);
	LUT4 #(
		.INIT('hffda)
	) name3871 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w4404_
	);
	LUT2 #(
		.INIT('h2)
	) name3872 (
		\sa02_reg[2]/P0001 ,
		_w4404_,
		_w4405_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name3873 (
		\sa02_reg[3]/P0001 ,
		\sa02_reg[4]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w4406_
	);
	LUT3 #(
		.INIT('h51)
	) name3874 (
		\sa02_reg[2]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w4407_
	);
	LUT3 #(
		.INIT('h45)
	) name3875 (
		_w3119_,
		_w4406_,
		_w4407_,
		_w4408_
	);
	LUT3 #(
		.INIT('h8a)
	) name3876 (
		\sa02_reg[1]/P0001 ,
		_w4405_,
		_w4408_,
		_w4409_
	);
	LUT4 #(
		.INIT('h0040)
	) name3877 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[3]/P0001 ,
		\sa02_reg[5]/P0001 ,
		\sa02_reg[7]/NET0131 ,
		_w4410_
	);
	LUT4 #(
		.INIT('h5540)
	) name3878 (
		\sa02_reg[2]/P0001 ,
		_w847_,
		_w923_,
		_w4410_,
		_w4411_
	);
	LUT3 #(
		.INIT('h80)
	) name3879 (
		\sa02_reg[2]/P0001 ,
		_w822_,
		_w878_,
		_w4412_
	);
	LUT3 #(
		.INIT('h13)
	) name3880 (
		_w832_,
		_w904_,
		_w3826_,
		_w4413_
	);
	LUT3 #(
		.INIT('h10)
	) name3881 (
		_w4411_,
		_w4412_,
		_w4413_,
		_w4414_
	);
	LUT3 #(
		.INIT('h80)
	) name3882 (
		\sa02_reg[1]/P0001 ,
		\sa02_reg[2]/P0001 ,
		\sa02_reg[3]/P0001 ,
		_w4415_
	);
	LUT2 #(
		.INIT('h8)
	) name3883 (
		_w862_,
		_w4415_,
		_w4416_
	);
	LUT3 #(
		.INIT('he0)
	) name3884 (
		_w864_,
		_w910_,
		_w3129_,
		_w4417_
	);
	LUT3 #(
		.INIT('had)
	) name3885 (
		\sa02_reg[5]/P0001 ,
		\sa02_reg[6]/NET0131 ,
		\sa02_reg[7]/NET0131 ,
		_w4418_
	);
	LUT2 #(
		.INIT('h2)
	) name3886 (
		_w3223_,
		_w4418_,
		_w4419_
	);
	LUT4 #(
		.INIT('h0001)
	) name3887 (
		_w4134_,
		_w4417_,
		_w4416_,
		_w4419_,
		_w4420_
	);
	LUT4 #(
		.INIT('hba00)
	) name3888 (
		\sa02_reg[0]/P0001 ,
		_w4409_,
		_w4414_,
		_w4420_,
		_w4421_
	);
	LUT3 #(
		.INIT('h10)
	) name3889 (
		_w4391_,
		_w4403_,
		_w4421_,
		_w4422_
	);
	LUT3 #(
		.INIT('h69)
	) name3890 (
		_w3795_,
		_w4378_,
		_w4422_,
		_w4423_
	);
	LUT3 #(
		.INIT('h54)
	) name3891 (
		\sa20_reg[2]/P0001 ,
		_w731_,
		_w3550_,
		_w4424_
	);
	LUT4 #(
		.INIT('h0020)
	) name3892 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4425_
	);
	LUT4 #(
		.INIT('h0001)
	) name3893 (
		_w3370_,
		_w3571_,
		_w3597_,
		_w4425_,
		_w4426_
	);
	LUT3 #(
		.INIT('h01)
	) name3894 (
		\sa20_reg[1]/P0001 ,
		_w663_,
		_w3600_,
		_w4427_
	);
	LUT3 #(
		.INIT('h40)
	) name3895 (
		_w4424_,
		_w4426_,
		_w4427_,
		_w4428_
	);
	LUT2 #(
		.INIT('h8)
	) name3896 (
		_w3968_,
		_w4058_,
		_w4429_
	);
	LUT4 #(
		.INIT('h0002)
	) name3897 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4430_
	);
	LUT4 #(
		.INIT('h002a)
	) name3898 (
		\sa20_reg[1]/P0001 ,
		_w673_,
		_w686_,
		_w4430_,
		_w4431_
	);
	LUT2 #(
		.INIT('h4)
	) name3899 (
		_w4429_,
		_w4431_,
		_w4432_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name3900 (
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4433_
	);
	LUT2 #(
		.INIT('h2)
	) name3901 (
		_w692_,
		_w4433_,
		_w4434_
	);
	LUT3 #(
		.INIT('ha8)
	) name3902 (
		\sa20_reg[5]/P0001 ,
		_w731_,
		_w4425_,
		_w4435_
	);
	LUT3 #(
		.INIT('h2a)
	) name3903 (
		\sa20_reg[0]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w711_,
		_w4436_
	);
	LUT3 #(
		.INIT('h10)
	) name3904 (
		_w4434_,
		_w4435_,
		_w4436_,
		_w4437_
	);
	LUT3 #(
		.INIT('he0)
	) name3905 (
		_w4428_,
		_w4432_,
		_w4437_,
		_w4438_
	);
	LUT4 #(
		.INIT('hffda)
	) name3906 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4439_
	);
	LUT4 #(
		.INIT('h0a02)
	) name3907 (
		\sa20_reg[1]/P0001 ,
		\sa20_reg[2]/P0001 ,
		_w720_,
		_w4439_,
		_w4440_
	);
	LUT4 #(
		.INIT('h0040)
	) name3908 (
		\sa20_reg[2]/P0001 ,
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w4441_
	);
	LUT3 #(
		.INIT('h01)
	) name3909 (
		\sa20_reg[1]/P0001 ,
		_w3381_,
		_w4441_,
		_w4442_
	);
	LUT2 #(
		.INIT('h1)
	) name3910 (
		_w4440_,
		_w4442_,
		_w4443_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name3911 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4444_
	);
	LUT4 #(
		.INIT('h1131)
	) name3912 (
		\sa20_reg[1]/P0001 ,
		\sa20_reg[2]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[7]/NET0131 ,
		_w4445_
	);
	LUT4 #(
		.INIT('h7770)
	) name3913 (
		_w700_,
		_w740_,
		_w4444_,
		_w4445_,
		_w4446_
	);
	LUT2 #(
		.INIT('h1)
	) name3914 (
		\sa20_reg[0]/P0001 ,
		_w666_,
		_w4447_
	);
	LUT3 #(
		.INIT('he0)
	) name3915 (
		_w3382_,
		_w4446_,
		_w4447_,
		_w4448_
	);
	LUT2 #(
		.INIT('h4)
	) name3916 (
		_w4443_,
		_w4448_,
		_w4449_
	);
	LUT3 #(
		.INIT('h01)
	) name3917 (
		\sa20_reg[2]/P0001 ,
		_w724_,
		_w3331_,
		_w4450_
	);
	LUT3 #(
		.INIT('h13)
	) name3918 (
		\sa20_reg[4]/P0001 ,
		_w663_,
		_w701_,
		_w4451_
	);
	LUT3 #(
		.INIT('h02)
	) name3919 (
		\sa20_reg[2]/P0001 ,
		_w3381_,
		_w3383_,
		_w4452_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name3920 (
		_w3589_,
		_w4450_,
		_w4451_,
		_w4452_,
		_w4453_
	);
	LUT4 #(
		.INIT('h000b)
	) name3921 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		_w4454_
	);
	LUT2 #(
		.INIT('h4)
	) name3922 (
		_w681_,
		_w4454_,
		_w4455_
	);
	LUT3 #(
		.INIT('h54)
	) name3923 (
		\sa20_reg[1]/P0001 ,
		_w4453_,
		_w4455_,
		_w4456_
	);
	LUT4 #(
		.INIT('h0400)
	) name3924 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[4]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4457_
	);
	LUT4 #(
		.INIT('h0013)
	) name3925 (
		_w647_,
		_w661_,
		_w3510_,
		_w4457_,
		_w4458_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name3926 (
		\sa20_reg[1]/P0001 ,
		\sa20_reg[2]/P0001 ,
		_w640_,
		_w4458_,
		_w4459_
	);
	LUT4 #(
		.INIT('haadf)
	) name3927 (
		\sa20_reg[3]/P0001 ,
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4460_
	);
	LUT4 #(
		.INIT('hc0c4)
	) name3928 (
		\sa20_reg[4]/P0001 ,
		_w727_,
		_w3550_,
		_w4460_,
		_w4461_
	);
	LUT3 #(
		.INIT('had)
	) name3929 (
		\sa20_reg[5]/P0001 ,
		\sa20_reg[6]/NET0131 ,
		\sa20_reg[7]/NET0131 ,
		_w4462_
	);
	LUT4 #(
		.INIT('h7707)
	) name3930 (
		_w686_,
		_w3569_,
		_w4083_,
		_w4462_,
		_w4463_
	);
	LUT2 #(
		.INIT('h4)
	) name3931 (
		_w4461_,
		_w4463_,
		_w4464_
	);
	LUT2 #(
		.INIT('h4)
	) name3932 (
		_w4459_,
		_w4464_,
		_w4465_
	);
	LUT4 #(
		.INIT('h5400)
	) name3933 (
		_w4456_,
		_w4438_,
		_w4449_,
		_w4465_,
		_w4466_
	);
	LUT3 #(
		.INIT('h69)
	) name3934 (
		\u0_w_reg[2][2]/P0001 ,
		_w4046_,
		_w4466_,
		_w4467_
	);
	LUT3 #(
		.INIT('h28)
	) name3935 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[34]/P0001 ,
		\u0_w_reg[2][2]/P0001 ,
		_w4468_
	);
	LUT4 #(
		.INIT('hff41)
	) name3936 (
		\ld_r_reg/P0001 ,
		_w4423_,
		_w4467_,
		_w4468_,
		_w4469_
	);
	LUT4 #(
		.INIT('h5655)
	) name3937 (
		\u0_w_reg[2][25]/P0001 ,
		_w4031_,
		_w4015_,
		_w4045_,
		_w4470_
	);
	LUT3 #(
		.INIT('h69)
	) name3938 (
		_w3745_,
		_w3996_,
		_w4470_,
		_w4471_
	);
	LUT4 #(
		.INIT('h9669)
	) name3939 (
		_w3265_,
		_w3324_,
		_w3841_,
		_w4331_,
		_w4472_
	);
	LUT3 #(
		.INIT('h28)
	) name3940 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[57]/P0001 ,
		\u0_w_reg[2][25]/P0001 ,
		_w4473_
	);
	LUT4 #(
		.INIT('hff14)
	) name3941 (
		\ld_r_reg/P0001 ,
		_w4471_,
		_w4472_,
		_w4473_,
		_w4474_
	);
	LUT3 #(
		.INIT('h69)
	) name3942 (
		_w745_,
		_w3265_,
		_w3324_,
		_w4475_
	);
	LUT3 #(
		.INIT('h69)
	) name3943 (
		\u0_w_reg[2][15]/P0001 ,
		_w1039_,
		_w3949_,
		_w4476_
	);
	LUT3 #(
		.INIT('h82)
	) name3944 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[47]/P0001 ,
		\u0_w_reg[2][15]/P0001 ,
		_w4477_
	);
	LUT4 #(
		.INIT('h00eb)
	) name3945 (
		\ld_r_reg/P0001 ,
		_w4475_,
		_w4476_,
		_w4477_,
		_w4478_
	);
	LUT4 #(
		.INIT('h6996)
	) name3946 (
		_w3265_,
		_w3445_,
		_w3496_,
		_w4145_,
		_w4479_
	);
	LUT4 #(
		.INIT('h9669)
	) name3947 (
		\u0_w_reg[2][4]/P0001 ,
		_w3616_,
		_w3949_,
		_w4285_,
		_w4480_
	);
	LUT3 #(
		.INIT('h82)
	) name3948 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[36]/P0001 ,
		\u0_w_reg[2][4]/P0001 ,
		_w4481_
	);
	LUT4 #(
		.INIT('h00be)
	) name3949 (
		\ld_r_reg/P0001 ,
		_w4479_,
		_w4480_,
		_w4481_,
		_w4482_
	);
	LUT4 #(
		.INIT('h6996)
	) name3950 (
		\u0_w_reg[2][27]/P0001 ,
		_w4189_,
		_w4236_,
		_w4285_,
		_w4483_
	);
	LUT4 #(
		.INIT('h9669)
	) name3951 (
		_w3265_,
		_w3324_,
		_w4378_,
		_w4422_,
		_w4484_
	);
	LUT3 #(
		.INIT('h82)
	) name3952 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[59]/P0001 ,
		\u0_w_reg[2][27]/P0001 ,
		_w4485_
	);
	LUT4 #(
		.INIT('h00be)
	) name3953 (
		\ld_r_reg/P0001 ,
		_w4483_,
		_w4484_,
		_w4485_,
		_w4486_
	);
	LUT4 #(
		.INIT('h6996)
	) name3954 (
		\u0_w_reg[2][19]/P0001 ,
		_w3389_,
		_w4236_,
		_w4285_,
		_w4487_
	);
	LUT4 #(
		.INIT('h6996)
	) name3955 (
		_w3324_,
		_w4145_,
		_w4378_,
		_w4466_,
		_w4488_
	);
	LUT3 #(
		.INIT('h82)
	) name3956 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[51]/P0001 ,
		\u0_w_reg[2][19]/P0001 ,
		_w4489_
	);
	LUT4 #(
		.INIT('h00eb)
	) name3957 (
		\ld_r_reg/P0001 ,
		_w4487_,
		_w4488_,
		_w4489_,
		_w4490_
	);
	LUT4 #(
		.INIT('h6996)
	) name3958 (
		_w3389_,
		_w4145_,
		_w4189_,
		_w4466_,
		_w4491_
	);
	LUT4 #(
		.INIT('h0105)
	) name3959 (
		_w3646_,
		_w3635_,
		_w3679_,
		_w3919_,
		_w4492_
	);
	LUT3 #(
		.INIT('h01)
	) name3960 (
		_w3638_,
		_w3669_,
		_w3846_,
		_w4493_
	);
	LUT4 #(
		.INIT('h0045)
	) name3961 (
		\sa31_reg[1]/P0001 ,
		\sa31_reg[2]/P0001 ,
		_w3188_,
		_w3631_,
		_w4494_
	);
	LUT3 #(
		.INIT('h80)
	) name3962 (
		_w4493_,
		_w4494_,
		_w4492_,
		_w4495_
	);
	LUT4 #(
		.INIT('h440c)
	) name3963 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w4496_
	);
	LUT4 #(
		.INIT('h5540)
	) name3964 (
		\sa31_reg[2]/P0001 ,
		_w940_,
		_w3164_,
		_w4496_,
		_w4497_
	);
	LUT4 #(
		.INIT('h0002)
	) name3965 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4498_
	);
	LUT2 #(
		.INIT('h2)
	) name3966 (
		\sa31_reg[1]/P0001 ,
		_w4498_,
		_w4499_
	);
	LUT2 #(
		.INIT('h4)
	) name3967 (
		_w4497_,
		_w4499_,
		_w4500_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name3968 (
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4501_
	);
	LUT2 #(
		.INIT('h2)
	) name3969 (
		_w981_,
		_w4501_,
		_w4502_
	);
	LUT2 #(
		.INIT('h8)
	) name3970 (
		_w967_,
		_w992_,
		_w4503_
	);
	LUT3 #(
		.INIT('h2a)
	) name3971 (
		\sa31_reg[0]/P0002 ,
		_w961_,
		_w1030_,
		_w4504_
	);
	LUT4 #(
		.INIT('h0100)
	) name3972 (
		_w3871_,
		_w4502_,
		_w4503_,
		_w4504_,
		_w4505_
	);
	LUT3 #(
		.INIT('he0)
	) name3973 (
		_w4495_,
		_w4500_,
		_w4505_,
		_w4506_
	);
	LUT3 #(
		.INIT('h02)
	) name3974 (
		\sa31_reg[2]/P0001 ,
		_w3169_,
		_w3919_,
		_w4507_
	);
	LUT4 #(
		.INIT('ha020)
	) name3975 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4508_
	);
	LUT4 #(
		.INIT('h5554)
	) name3976 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w4509_
	);
	LUT2 #(
		.INIT('h4)
	) name3977 (
		_w4508_,
		_w4509_,
		_w4510_
	);
	LUT4 #(
		.INIT('h0040)
	) name3978 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w4511_
	);
	LUT3 #(
		.INIT('h01)
	) name3979 (
		\sa31_reg[1]/P0001 ,
		_w3891_,
		_w4511_,
		_w4512_
	);
	LUT4 #(
		.INIT('h0057)
	) name3980 (
		_w3897_,
		_w4507_,
		_w4510_,
		_w4512_,
		_w4513_
	);
	LUT3 #(
		.INIT('h40)
	) name3981 (
		\sa31_reg[2]/P0001 ,
		_w947_,
		_w1035_,
		_w4514_
	);
	LUT3 #(
		.INIT('h20)
	) name3982 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[5]/P0001 ,
		_w3667_,
		_w4515_
	);
	LUT2 #(
		.INIT('h1)
	) name3983 (
		\sa31_reg[0]/P0002 ,
		_w962_,
		_w4516_
	);
	LUT3 #(
		.INIT('h10)
	) name3984 (
		_w4515_,
		_w4514_,
		_w4516_,
		_w4517_
	);
	LUT2 #(
		.INIT('h4)
	) name3985 (
		_w4513_,
		_w4517_,
		_w4518_
	);
	LUT3 #(
		.INIT('h01)
	) name3986 (
		_w1017_,
		_w3657_,
		_w3679_,
		_w4519_
	);
	LUT3 #(
		.INIT('h02)
	) name3987 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w4520_
	);
	LUT3 #(
		.INIT('h02)
	) name3988 (
		\sa31_reg[2]/P0001 ,
		_w3891_,
		_w4520_,
		_w4521_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name3989 (
		_w3672_,
		_w3909_,
		_w4519_,
		_w4521_,
		_w4522_
	);
	LUT4 #(
		.INIT('h0008)
	) name3990 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		_w4523_
	);
	LUT3 #(
		.INIT('h01)
	) name3991 (
		\sa31_reg[1]/P0001 ,
		_w3643_,
		_w4523_,
		_w4524_
	);
	LUT4 #(
		.INIT('h0400)
	) name3992 (
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4525_
	);
	LUT2 #(
		.INIT('h1)
	) name3993 (
		\sa31_reg[2]/P0001 ,
		_w4525_,
		_w4526_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3994 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		\sa31_reg[7]/P0001 ,
		_w4527_
	);
	LUT4 #(
		.INIT('h0700)
	) name3995 (
		_w996_,
		_w3172_,
		_w3188_,
		_w4527_,
		_w4528_
	);
	LUT2 #(
		.INIT('h2)
	) name3996 (
		\sa31_reg[1]/P0001 ,
		_w3152_,
		_w4529_
	);
	LUT4 #(
		.INIT('hf800)
	) name3997 (
		_w4002_,
		_w4526_,
		_w4528_,
		_w4529_,
		_w4530_
	);
	LUT3 #(
		.INIT('had)
	) name3998 (
		\sa31_reg[5]/P0001 ,
		\sa31_reg[6]/NET0131 ,
		\sa31_reg[7]/P0001 ,
		_w4531_
	);
	LUT3 #(
		.INIT('h02)
	) name3999 (
		\sa31_reg[2]/P0001 ,
		\sa31_reg[3]/P0001 ,
		\sa31_reg[4]/P0001 ,
		_w4532_
	);
	LUT2 #(
		.INIT('h4)
	) name4000 (
		_w4531_,
		_w4532_,
		_w4533_
	);
	LUT2 #(
		.INIT('h1)
	) name4001 (
		_w4277_,
		_w4533_,
		_w4534_
	);
	LUT4 #(
		.INIT('hf400)
	) name4002 (
		_w4522_,
		_w4524_,
		_w4530_,
		_w4534_,
		_w4535_
	);
	LUT3 #(
		.INIT('he0)
	) name4003 (
		_w4506_,
		_w4518_,
		_w4535_,
		_w4536_
	);
	LUT4 #(
		.INIT('h6996)
	) name4004 (
		\u0_w_reg[2][11]/P0001 ,
		_w3949_,
		_w4285_,
		_w4536_,
		_w4537_
	);
	LUT3 #(
		.INIT('h82)
	) name4005 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[43]/P0001 ,
		\u0_w_reg[2][11]/P0001 ,
		_w4538_
	);
	LUT4 #(
		.INIT('h00eb)
	) name4006 (
		\ld_r_reg/P0001 ,
		_w4491_,
		_w4537_,
		_w4538_,
		_w4539_
	);
	LUT4 #(
		.INIT('ha955)
	) name4007 (
		\u0_w_reg[2][26]/P0001 ,
		_w4506_,
		_w4518_,
		_w4535_,
		_w4540_
	);
	LUT3 #(
		.INIT('h69)
	) name4008 (
		_w4378_,
		_w4466_,
		_w4540_,
		_w4541_
	);
	LUT3 #(
		.INIT('h28)
	) name4009 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[58]/P0001 ,
		\u0_w_reg[2][26]/P0001 ,
		_w4542_
	);
	LUT4 #(
		.INIT('hff41)
	) name4010 (
		\ld_r_reg/P0001 ,
		_w3796_,
		_w4541_,
		_w4542_,
		_w4543_
	);
	LUT4 #(
		.INIT('h6996)
	) name4011 (
		_w3265_,
		_w4145_,
		_w4189_,
		_w4422_,
		_w4544_
	);
	LUT4 #(
		.INIT('h6996)
	) name4012 (
		\u0_w_reg[2][3]/P0001 ,
		_w3949_,
		_w4236_,
		_w4536_,
		_w4545_
	);
	LUT3 #(
		.INIT('h82)
	) name4013 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[35]/P0001 ,
		\u0_w_reg[2][3]/P0001 ,
		_w4546_
	);
	LUT4 #(
		.INIT('h00eb)
	) name4014 (
		\ld_r_reg/P0001 ,
		_w4544_,
		_w4545_,
		_w4546_,
		_w4547_
	);
	LUT2 #(
		.INIT('h9)
	) name4015 (
		\u0_w_reg[2][31]/P0001 ,
		_w3324_,
		_w4548_
	);
	LUT4 #(
		.INIT('h6996)
	) name4016 (
		_w637_,
		_w3142_,
		_w3389_,
		_w3949_,
		_w4549_
	);
	LUT3 #(
		.INIT('h82)
	) name4017 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[63]/P0001 ,
		\u0_w_reg[2][31]/P0001 ,
		_w4550_
	);
	LUT4 #(
		.INIT('h00be)
	) name4018 (
		\ld_r_reg/P0001 ,
		_w4548_,
		_w4549_,
		_w4550_,
		_w4551_
	);
	LUT2 #(
		.INIT('h6)
	) name4019 (
		\u0_w_reg[2][24]/P0001 ,
		_w3896_,
		_w4552_
	);
	LUT4 #(
		.INIT('h9669)
	) name4020 (
		_w3265_,
		_w3324_,
		_w4093_,
		_w4331_,
		_w4553_
	);
	LUT3 #(
		.INIT('h28)
	) name4021 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[56]/P0001 ,
		\u0_w_reg[2][24]/P0001 ,
		_w4554_
	);
	LUT4 #(
		.INIT('hff14)
	) name4022 (
		\ld_r_reg/P0001 ,
		_w4552_,
		_w4553_,
		_w4554_,
		_w4555_
	);
	LUT2 #(
		.INIT('h6)
	) name4023 (
		\u0_w_reg[2][16]/P0001 ,
		_w3896_,
		_w4556_
	);
	LUT4 #(
		.INIT('h6996)
	) name4024 (
		_w3324_,
		_w3389_,
		_w3841_,
		_w4093_,
		_w4557_
	);
	LUT3 #(
		.INIT('h28)
	) name4025 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[48]/P0001 ,
		\u0_w_reg[2][16]/P0001 ,
		_w4558_
	);
	LUT4 #(
		.INIT('hff41)
	) name4026 (
		\ld_r_reg/P0001 ,
		_w4556_,
		_w4557_,
		_w4558_,
		_w4559_
	);
	LUT3 #(
		.INIT('h69)
	) name4027 (
		_w3745_,
		_w3996_,
		_w4422_,
		_w4560_
	);
	LUT4 #(
		.INIT('ha955)
	) name4028 (
		\u0_w_reg[2][18]/P0001 ,
		_w4506_,
		_w4518_,
		_w4535_,
		_w4561_
	);
	LUT2 #(
		.INIT('h6)
	) name4029 (
		_w4466_,
		_w4561_,
		_w4562_
	);
	LUT3 #(
		.INIT('h82)
	) name4030 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[50]/P0001 ,
		\u0_w_reg[2][18]/P0001 ,
		_w4563_
	);
	LUT4 #(
		.INIT('h00eb)
	) name4031 (
		\ld_r_reg/P0001 ,
		_w4560_,
		_w4562_,
		_w4563_,
		_w4564_
	);
	LUT3 #(
		.INIT('h69)
	) name4032 (
		_w637_,
		_w745_,
		_w3265_,
		_w4565_
	);
	LUT3 #(
		.INIT('h69)
	) name4033 (
		\u0_w_reg[2][23]/P0001 ,
		_w3389_,
		_w3949_,
		_w4566_
	);
	LUT3 #(
		.INIT('h82)
	) name4034 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[55]/P0001 ,
		\u0_w_reg[2][23]/P0001 ,
		_w4567_
	);
	LUT4 #(
		.INIT('h00eb)
	) name4035 (
		\ld_r_reg/P0001 ,
		_w4565_,
		_w4566_,
		_w4567_,
		_w4568_
	);
	LUT2 #(
		.INIT('h6)
	) name4036 (
		\u0_w_reg[2][8]/P0001 ,
		_w3896_,
		_w4569_
	);
	LUT4 #(
		.INIT('h6996)
	) name4037 (
		_w3389_,
		_w3841_,
		_w3949_,
		_w4331_,
		_w4570_
	);
	LUT3 #(
		.INIT('h82)
	) name4038 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[40]/P0001 ,
		\u0_w_reg[2][8]/P0001 ,
		_w4571_
	);
	LUT4 #(
		.INIT('h00eb)
	) name4039 (
		\ld_r_reg/P0001 ,
		_w4569_,
		_w4570_,
		_w4571_,
		_w4572_
	);
	LUT3 #(
		.INIT('h69)
	) name4040 (
		_w3996_,
		_w4378_,
		_w4422_,
		_w4573_
	);
	LUT4 #(
		.INIT('ha955)
	) name4041 (
		\u0_w_reg[2][10]/P0001 ,
		_w4506_,
		_w4518_,
		_w4535_,
		_w4574_
	);
	LUT2 #(
		.INIT('h6)
	) name4042 (
		_w4046_,
		_w4574_,
		_w4575_
	);
	LUT3 #(
		.INIT('h82)
	) name4043 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[42]/P0001 ,
		\u0_w_reg[2][10]/P0001 ,
		_w4576_
	);
	LUT4 #(
		.INIT('h00eb)
	) name4044 (
		\ld_r_reg/P0001 ,
		_w4573_,
		_w4575_,
		_w4576_,
		_w4577_
	);
	LUT2 #(
		.INIT('h9)
	) name4045 (
		\u0_w_reg[2][5]/P0001 ,
		_w3205_,
		_w4578_
	);
	LUT4 #(
		.INIT('h5655)
	) name4046 (
		\u0_w_reg[2][6]/P0001 ,
		_w980_,
		_w1009_,
		_w1038_,
		_w4579_
	);
	LUT2 #(
		.INIT('h9)
	) name4047 (
		\u0_w_reg[2][4]/P0001 ,
		_w3686_,
		_w4580_
	);
	LUT2 #(
		.INIT('h9)
	) name4048 (
		\u0_w_reg[2][0]/P0001 ,
		_w3896_,
		_w4581_
	);
	LUT2 #(
		.INIT('h9)
	) name4049 (
		\u0_w_reg[2][3]/P0001 ,
		_w4285_,
		_w4582_
	);
	LUT4 #(
		.INIT('h5655)
	) name4050 (
		\u0_w_reg[2][1]/P0001 ,
		_w4031_,
		_w4015_,
		_w4045_,
		_w4583_
	);
	LUT4 #(
		.INIT('ha955)
	) name4051 (
		\u0_w_reg[2][2]/P0001 ,
		_w4506_,
		_w4518_,
		_w4535_,
		_w4584_
	);
	LUT2 #(
		.INIT('h9)
	) name4052 (
		\u0_w_reg[2][7]/P0001 ,
		_w3949_,
		_w4585_
	);
	LUT2 #(
		.INIT('h8)
	) name4053 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4586_
	);
	LUT2 #(
		.INIT('h1)
	) name4054 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4587_
	);
	LUT4 #(
		.INIT('h0200)
	) name4055 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4588_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name4056 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4589_
	);
	LUT2 #(
		.INIT('h1)
	) name4057 (
		\sa12_reg[2]/P0001 ,
		_w4589_,
		_w4590_
	);
	LUT2 #(
		.INIT('h2)
	) name4058 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4591_
	);
	LUT2 #(
		.INIT('h2)
	) name4059 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4592_
	);
	LUT3 #(
		.INIT('h02)
	) name4060 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4593_
	);
	LUT2 #(
		.INIT('h8)
	) name4061 (
		_w4591_,
		_w4593_,
		_w4594_
	);
	LUT2 #(
		.INIT('h4)
	) name4062 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4595_
	);
	LUT3 #(
		.INIT('h01)
	) name4063 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4596_
	);
	LUT2 #(
		.INIT('h2)
	) name4064 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4597_
	);
	LUT4 #(
		.INIT('h0200)
	) name4065 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4598_
	);
	LUT4 #(
		.INIT('h002a)
	) name4066 (
		\sa12_reg[1]/P0001 ,
		_w4595_,
		_w4596_,
		_w4598_,
		_w4599_
	);
	LUT3 #(
		.INIT('h10)
	) name4067 (
		_w4590_,
		_w4594_,
		_w4599_,
		_w4600_
	);
	LUT2 #(
		.INIT('h8)
	) name4068 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4601_
	);
	LUT3 #(
		.INIT('h80)
	) name4069 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4602_
	);
	LUT4 #(
		.INIT('h0800)
	) name4070 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4603_
	);
	LUT2 #(
		.INIT('h8)
	) name4071 (
		\sa12_reg[2]/P0001 ,
		_w4603_,
		_w4604_
	);
	LUT2 #(
		.INIT('h4)
	) name4072 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		_w4605_
	);
	LUT3 #(
		.INIT('h02)
	) name4073 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4606_
	);
	LUT3 #(
		.INIT('h15)
	) name4074 (
		\sa12_reg[1]/P0001 ,
		_w4605_,
		_w4606_,
		_w4607_
	);
	LUT2 #(
		.INIT('h8)
	) name4075 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4608_
	);
	LUT3 #(
		.INIT('h80)
	) name4076 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4609_
	);
	LUT4 #(
		.INIT('h2000)
	) name4077 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4610_
	);
	LUT2 #(
		.INIT('h1)
	) name4078 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4611_
	);
	LUT3 #(
		.INIT('h32)
	) name4079 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4612_
	);
	LUT3 #(
		.INIT('h51)
	) name4080 (
		_w4610_,
		_w4601_,
		_w4612_,
		_w4613_
	);
	LUT3 #(
		.INIT('h20)
	) name4081 (
		_w4607_,
		_w4604_,
		_w4613_,
		_w4614_
	);
	LUT3 #(
		.INIT('h80)
	) name4082 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4615_
	);
	LUT3 #(
		.INIT('h54)
	) name4083 (
		_w4586_,
		_w4595_,
		_w4615_,
		_w4616_
	);
	LUT2 #(
		.INIT('h2)
	) name4084 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		_w4617_
	);
	LUT4 #(
		.INIT('h0200)
	) name4085 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4618_
	);
	LUT3 #(
		.INIT('h02)
	) name4086 (
		\sa12_reg[2]/P0001 ,
		_w4618_,
		_w4593_,
		_w4619_
	);
	LUT2 #(
		.INIT('h4)
	) name4087 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4620_
	);
	LUT4 #(
		.INIT('h2000)
	) name4088 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4621_
	);
	LUT2 #(
		.INIT('h1)
	) name4089 (
		\sa12_reg[2]/P0001 ,
		_w4621_,
		_w4622_
	);
	LUT2 #(
		.INIT('h1)
	) name4090 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4623_
	);
	LUT4 #(
		.INIT('h0001)
	) name4091 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4624_
	);
	LUT2 #(
		.INIT('h4)
	) name4092 (
		\sa12_reg[7]/NET0131 ,
		_w4624_,
		_w4625_
	);
	LUT4 #(
		.INIT('h0020)
	) name4093 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4626_
	);
	LUT3 #(
		.INIT('h0b)
	) name4094 (
		\sa12_reg[7]/NET0131 ,
		_w4624_,
		_w4626_,
		_w4627_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name4095 (
		_w4616_,
		_w4619_,
		_w4622_,
		_w4627_,
		_w4628_
	);
	LUT4 #(
		.INIT('h2220)
	) name4096 (
		\sa12_reg[0]/P0001 ,
		_w4628_,
		_w4600_,
		_w4614_,
		_w4629_
	);
	LUT4 #(
		.INIT('h0100)
	) name4097 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4630_
	);
	LUT3 #(
		.INIT('h20)
	) name4098 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4631_
	);
	LUT4 #(
		.INIT('h5150)
	) name4099 (
		\sa12_reg[2]/P0001 ,
		_w4592_,
		_w4630_,
		_w4631_,
		_w4632_
	);
	LUT3 #(
		.INIT('h08)
	) name4100 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4633_
	);
	LUT4 #(
		.INIT('h0080)
	) name4101 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4634_
	);
	LUT2 #(
		.INIT('h2)
	) name4102 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		_w4635_
	);
	LUT3 #(
		.INIT('h20)
	) name4103 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4636_
	);
	LUT2 #(
		.INIT('h8)
	) name4104 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4637_
	);
	LUT4 #(
		.INIT('h0080)
	) name4105 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4638_
	);
	LUT4 #(
		.INIT('h020a)
	) name4106 (
		\sa12_reg[1]/P0001 ,
		_w4635_,
		_w4638_,
		_w4636_,
		_w4639_
	);
	LUT4 #(
		.INIT('h0002)
	) name4107 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4640_
	);
	LUT4 #(
		.INIT('h0002)
	) name4108 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4641_
	);
	LUT2 #(
		.INIT('h8)
	) name4109 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4642_
	);
	LUT4 #(
		.INIT('h8000)
	) name4110 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4643_
	);
	LUT4 #(
		.INIT('h0001)
	) name4111 (
		\sa12_reg[1]/P0001 ,
		_w4643_,
		_w4641_,
		_w4640_,
		_w4644_
	);
	LUT4 #(
		.INIT('h00ef)
	) name4112 (
		_w4632_,
		_w4634_,
		_w4639_,
		_w4644_,
		_w4645_
	);
	LUT4 #(
		.INIT('h0040)
	) name4113 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4646_
	);
	LUT2 #(
		.INIT('h4)
	) name4114 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4647_
	);
	LUT4 #(
		.INIT('h0400)
	) name4115 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4648_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name4116 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4648_,
		_w4646_,
		_w4649_
	);
	LUT4 #(
		.INIT('h0008)
	) name4117 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4650_
	);
	LUT3 #(
		.INIT('h10)
	) name4118 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4651_
	);
	LUT4 #(
		.INIT('h0100)
	) name4119 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4652_
	);
	LUT3 #(
		.INIT('h0b)
	) name4120 (
		\sa12_reg[6]/NET0131 ,
		_w4650_,
		_w4652_,
		_w4653_
	);
	LUT3 #(
		.INIT('h02)
	) name4121 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4654_
	);
	LUT2 #(
		.INIT('h8)
	) name4122 (
		_w4654_,
		_w4623_,
		_w4655_
	);
	LUT3 #(
		.INIT('h15)
	) name4123 (
		\sa12_reg[0]/P0001 ,
		_w4654_,
		_w4623_,
		_w4656_
	);
	LUT4 #(
		.INIT('he400)
	) name4124 (
		\sa12_reg[2]/P0001 ,
		_w4649_,
		_w4653_,
		_w4656_,
		_w4657_
	);
	LUT2 #(
		.INIT('h4)
	) name4125 (
		_w4645_,
		_w4657_,
		_w4658_
	);
	LUT2 #(
		.INIT('h2)
	) name4126 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4659_
	);
	LUT4 #(
		.INIT('h0020)
	) name4127 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4660_
	);
	LUT4 #(
		.INIT('h0080)
	) name4128 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4661_
	);
	LUT3 #(
		.INIT('h02)
	) name4129 (
		\sa12_reg[2]/P0001 ,
		_w4661_,
		_w4660_,
		_w4662_
	);
	LUT4 #(
		.INIT('h0004)
	) name4130 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4663_
	);
	LUT3 #(
		.INIT('h80)
	) name4131 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4664_
	);
	LUT2 #(
		.INIT('h4)
	) name4132 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4665_
	);
	LUT3 #(
		.INIT('h10)
	) name4133 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4666_
	);
	LUT4 #(
		.INIT('h0037)
	) name4134 (
		_w4664_,
		_w4587_,
		_w4666_,
		_w4663_,
		_w4667_
	);
	LUT4 #(
		.INIT('h2000)
	) name4135 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4668_
	);
	LUT2 #(
		.INIT('h8)
	) name4136 (
		\sa12_reg[7]/NET0131 ,
		_w4668_,
		_w4669_
	);
	LUT4 #(
		.INIT('h1000)
	) name4137 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4670_
	);
	LUT3 #(
		.INIT('h01)
	) name4138 (
		\sa12_reg[2]/P0001 ,
		_w4648_,
		_w4670_,
		_w4671_
	);
	LUT4 #(
		.INIT('h7077)
	) name4139 (
		_w4662_,
		_w4667_,
		_w4669_,
		_w4671_,
		_w4672_
	);
	LUT3 #(
		.INIT('h15)
	) name4140 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4661_,
		_w4673_
	);
	LUT2 #(
		.INIT('h4)
	) name4141 (
		_w4655_,
		_w4673_,
		_w4674_
	);
	LUT4 #(
		.INIT('h4000)
	) name4142 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4675_
	);
	LUT4 #(
		.INIT('h2220)
	) name4143 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4676_
	);
	LUT3 #(
		.INIT('h0b)
	) name4144 (
		\sa12_reg[4]/P0001 ,
		_w4675_,
		_w4676_,
		_w4677_
	);
	LUT3 #(
		.INIT('h45)
	) name4145 (
		\sa12_reg[2]/P0001 ,
		_w4625_,
		_w4677_,
		_w4678_
	);
	LUT4 #(
		.INIT('h0200)
	) name4146 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4679_
	);
	LUT2 #(
		.INIT('h4)
	) name4147 (
		\sa12_reg[6]/NET0131 ,
		_w4679_,
		_w4680_
	);
	LUT3 #(
		.INIT('h2a)
	) name4148 (
		\sa12_reg[1]/P0001 ,
		_w4664_,
		_w4647_,
		_w4681_
	);
	LUT2 #(
		.INIT('h4)
	) name4149 (
		_w4680_,
		_w4681_,
		_w4682_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4150 (
		_w4672_,
		_w4674_,
		_w4678_,
		_w4682_,
		_w4683_
	);
	LUT2 #(
		.INIT('h8)
	) name4151 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		_w4684_
	);
	LUT3 #(
		.INIT('h08)
	) name4152 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4685_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name4153 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		_w4654_,
		_w4685_,
		_w4686_
	);
	LUT2 #(
		.INIT('h4)
	) name4154 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4687_
	);
	LUT4 #(
		.INIT('h0010)
	) name4155 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4688_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name4156 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		_w4643_,
		_w4688_,
		_w4689_
	);
	LUT3 #(
		.INIT('h0d)
	) name4157 (
		\sa12_reg[1]/P0001 ,
		_w4686_,
		_w4689_,
		_w4690_
	);
	LUT4 #(
		.INIT('h5400)
	) name4158 (
		_w4683_,
		_w4629_,
		_w4658_,
		_w4690_,
		_w4691_
	);
	LUT2 #(
		.INIT('h2)
	) name4159 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w4692_
	);
	LUT3 #(
		.INIT('h20)
	) name4160 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4693_
	);
	LUT3 #(
		.INIT('h10)
	) name4161 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w4694_
	);
	LUT4 #(
		.INIT('h0100)
	) name4162 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4695_
	);
	LUT4 #(
		.INIT('h5510)
	) name4163 (
		\sa01_reg[2]/P0001 ,
		_w4692_,
		_w4693_,
		_w4695_,
		_w4696_
	);
	LUT2 #(
		.INIT('h4)
	) name4164 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w4697_
	);
	LUT2 #(
		.INIT('h4)
	) name4165 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w4698_
	);
	LUT3 #(
		.INIT('h20)
	) name4166 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w4699_
	);
	LUT2 #(
		.INIT('h8)
	) name4167 (
		_w4697_,
		_w4699_,
		_w4700_
	);
	LUT2 #(
		.INIT('h2)
	) name4168 (
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4701_
	);
	LUT3 #(
		.INIT('h08)
	) name4169 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4702_
	);
	LUT4 #(
		.INIT('h0080)
	) name4170 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4703_
	);
	LUT2 #(
		.INIT('h8)
	) name4171 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w4704_
	);
	LUT4 #(
		.INIT('h0080)
	) name4172 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4705_
	);
	LUT3 #(
		.INIT('h02)
	) name4173 (
		\sa01_reg[1]/P0001 ,
		_w4703_,
		_w4705_,
		_w4706_
	);
	LUT3 #(
		.INIT('h10)
	) name4174 (
		_w4696_,
		_w4700_,
		_w4706_,
		_w4707_
	);
	LUT2 #(
		.INIT('h1)
	) name4175 (
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4708_
	);
	LUT3 #(
		.INIT('h01)
	) name4176 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4709_
	);
	LUT4 #(
		.INIT('h7f7c)
	) name4177 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4710_
	);
	LUT2 #(
		.INIT('h2)
	) name4178 (
		\sa01_reg[2]/P0001 ,
		_w4710_,
		_w4711_
	);
	LUT4 #(
		.INIT('h0040)
	) name4179 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4712_
	);
	LUT4 #(
		.INIT('h0002)
	) name4180 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4713_
	);
	LUT4 #(
		.INIT('h0045)
	) name4181 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[2]/P0001 ,
		_w4712_,
		_w4713_,
		_w4714_
	);
	LUT2 #(
		.INIT('h4)
	) name4182 (
		_w4711_,
		_w4714_,
		_w4715_
	);
	LUT2 #(
		.INIT('h2)
	) name4183 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[5]/P0001 ,
		_w4716_
	);
	LUT2 #(
		.INIT('h1)
	) name4184 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w4717_
	);
	LUT3 #(
		.INIT('h10)
	) name4185 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w4718_
	);
	LUT4 #(
		.INIT('h0008)
	) name4186 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4719_
	);
	LUT4 #(
		.INIT('hefe7)
	) name4187 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4720_
	);
	LUT2 #(
		.INIT('h2)
	) name4188 (
		_w4716_,
		_w4720_,
		_w4721_
	);
	LUT4 #(
		.INIT('h0004)
	) name4189 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4722_
	);
	LUT2 #(
		.INIT('h4)
	) name4190 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w4723_
	);
	LUT2 #(
		.INIT('h8)
	) name4191 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w4724_
	);
	LUT3 #(
		.INIT('h40)
	) name4192 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w4725_
	);
	LUT4 #(
		.INIT('h5444)
	) name4193 (
		\sa01_reg[3]/P0001 ,
		_w4722_,
		_w4723_,
		_w4725_,
		_w4726_
	);
	LUT2 #(
		.INIT('h1)
	) name4194 (
		_w4721_,
		_w4726_,
		_w4727_
	);
	LUT4 #(
		.INIT('h0155)
	) name4195 (
		\sa01_reg[0]/P0001 ,
		_w4707_,
		_w4715_,
		_w4727_,
		_w4728_
	);
	LUT3 #(
		.INIT('he0)
	) name4196 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4729_
	);
	LUT4 #(
		.INIT('h5410)
	) name4197 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4730_
	);
	LUT2 #(
		.INIT('h4)
	) name4198 (
		_w4729_,
		_w4730_,
		_w4731_
	);
	LUT3 #(
		.INIT('h02)
	) name4199 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4732_
	);
	LUT2 #(
		.INIT('h8)
	) name4200 (
		_w4692_,
		_w4732_,
		_w4733_
	);
	LUT2 #(
		.INIT('h2)
	) name4201 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w4734_
	);
	LUT4 #(
		.INIT('h0200)
	) name4202 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4735_
	);
	LUT4 #(
		.INIT('h002a)
	) name4203 (
		\sa01_reg[1]/P0001 ,
		_w4698_,
		_w4709_,
		_w4735_,
		_w4736_
	);
	LUT3 #(
		.INIT('h10)
	) name4204 (
		_w4733_,
		_w4731_,
		_w4736_,
		_w4737_
	);
	LUT2 #(
		.INIT('h8)
	) name4205 (
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4738_
	);
	LUT4 #(
		.INIT('h2000)
	) name4206 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4739_
	);
	LUT3 #(
		.INIT('h08)
	) name4207 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w4740_
	);
	LUT2 #(
		.INIT('h1)
	) name4208 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w4741_
	);
	LUT4 #(
		.INIT('h0111)
	) name4209 (
		\sa01_reg[1]/P0001 ,
		_w4739_,
		_w4740_,
		_w4741_,
		_w4742_
	);
	LUT4 #(
		.INIT('h0800)
	) name4210 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4743_
	);
	LUT2 #(
		.INIT('h8)
	) name4211 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w4744_
	);
	LUT2 #(
		.INIT('h1)
	) name4212 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w4745_
	);
	LUT3 #(
		.INIT('h32)
	) name4213 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w4746_
	);
	LUT4 #(
		.INIT('h7707)
	) name4214 (
		\sa01_reg[2]/P0001 ,
		_w4743_,
		_w4744_,
		_w4746_,
		_w4747_
	);
	LUT2 #(
		.INIT('h8)
	) name4215 (
		_w4742_,
		_w4747_,
		_w4748_
	);
	LUT3 #(
		.INIT('h80)
	) name4216 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4749_
	);
	LUT2 #(
		.INIT('h2)
	) name4217 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w4750_
	);
	LUT3 #(
		.INIT('h02)
	) name4218 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w4751_
	);
	LUT3 #(
		.INIT('hb9)
	) name4219 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w4752_
	);
	LUT3 #(
		.INIT('h45)
	) name4220 (
		_w4724_,
		_w4749_,
		_w4752_,
		_w4753_
	);
	LUT4 #(
		.INIT('h0200)
	) name4221 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4754_
	);
	LUT2 #(
		.INIT('h2)
	) name4222 (
		\sa01_reg[2]/P0001 ,
		_w4754_,
		_w4755_
	);
	LUT2 #(
		.INIT('h8)
	) name4223 (
		_w4709_,
		_w4717_,
		_w4756_
	);
	LUT2 #(
		.INIT('h8)
	) name4224 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w4757_
	);
	LUT4 #(
		.INIT('h2000)
	) name4225 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4758_
	);
	LUT2 #(
		.INIT('h1)
	) name4226 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w4759_
	);
	LUT4 #(
		.INIT('h0020)
	) name4227 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4760_
	);
	LUT3 #(
		.INIT('h01)
	) name4228 (
		\sa01_reg[2]/P0001 ,
		_w4760_,
		_w4758_,
		_w4761_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4229 (
		_w4753_,
		_w4755_,
		_w4756_,
		_w4761_,
		_w4762_
	);
	LUT4 #(
		.INIT('haa02)
	) name4230 (
		\sa01_reg[0]/P0001 ,
		_w4737_,
		_w4748_,
		_w4762_,
		_w4763_
	);
	LUT3 #(
		.INIT('h10)
	) name4231 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w4764_
	);
	LUT4 #(
		.INIT('h1000)
	) name4232 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w4765_
	);
	LUT2 #(
		.INIT('h8)
	) name4233 (
		\sa01_reg[6]/NET0131 ,
		_w4765_,
		_w4766_
	);
	LUT2 #(
		.INIT('h2)
	) name4234 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		_w4767_
	);
	LUT4 #(
		.INIT('h2220)
	) name4235 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4768_
	);
	LUT3 #(
		.INIT('h07)
	) name4236 (
		_w4709_,
		_w4717_,
		_w4768_,
		_w4769_
	);
	LUT3 #(
		.INIT('h45)
	) name4237 (
		\sa01_reg[2]/P0001 ,
		_w4766_,
		_w4769_,
		_w4770_
	);
	LUT3 #(
		.INIT('h04)
	) name4238 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4771_
	);
	LUT2 #(
		.INIT('h8)
	) name4239 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w4772_
	);
	LUT3 #(
		.INIT('h2a)
	) name4240 (
		\sa01_reg[1]/P0001 ,
		_w4771_,
		_w4772_,
		_w4773_
	);
	LUT2 #(
		.INIT('h8)
	) name4241 (
		_w4697_,
		_w4751_,
		_w4774_
	);
	LUT2 #(
		.INIT('h8)
	) name4242 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		_w4775_
	);
	LUT3 #(
		.INIT('h20)
	) name4243 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w4776_
	);
	LUT4 #(
		.INIT('h135f)
	) name4244 (
		_w4732_,
		_w4757_,
		_w4775_,
		_w4776_,
		_w4777_
	);
	LUT3 #(
		.INIT('h40)
	) name4245 (
		_w4774_,
		_w4773_,
		_w4777_,
		_w4778_
	);
	LUT4 #(
		.INIT('h0080)
	) name4246 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4779_
	);
	LUT4 #(
		.INIT('h0020)
	) name4247 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w4780_
	);
	LUT3 #(
		.INIT('h02)
	) name4248 (
		\sa01_reg[2]/P0001 ,
		_w4780_,
		_w4779_,
		_w4781_
	);
	LUT3 #(
		.INIT('h01)
	) name4249 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4782_
	);
	LUT4 #(
		.INIT('h0004)
	) name4250 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4783_
	);
	LUT3 #(
		.INIT('h10)
	) name4251 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4784_
	);
	LUT2 #(
		.INIT('h9)
	) name4252 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w4785_
	);
	LUT3 #(
		.INIT('h15)
	) name4253 (
		_w4783_,
		_w4784_,
		_w4785_,
		_w4786_
	);
	LUT3 #(
		.INIT('h20)
	) name4254 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		_w4787_
	);
	LUT2 #(
		.INIT('h8)
	) name4255 (
		_w4738_,
		_w4787_,
		_w4788_
	);
	LUT2 #(
		.INIT('h1)
	) name4256 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		_w4789_
	);
	LUT4 #(
		.INIT('h1000)
	) name4257 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4790_
	);
	LUT4 #(
		.INIT('h0400)
	) name4258 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w4791_
	);
	LUT3 #(
		.INIT('h01)
	) name4259 (
		\sa01_reg[2]/P0001 ,
		_w4790_,
		_w4791_,
		_w4792_
	);
	LUT4 #(
		.INIT('h7077)
	) name4260 (
		_w4781_,
		_w4786_,
		_w4788_,
		_w4792_,
		_w4793_
	);
	LUT4 #(
		.INIT('h0001)
	) name4261 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4794_
	);
	LUT2 #(
		.INIT('h8)
	) name4262 (
		\sa01_reg[5]/P0001 ,
		_w4794_,
		_w4795_
	);
	LUT4 #(
		.INIT('h0080)
	) name4263 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w4796_
	);
	LUT3 #(
		.INIT('h15)
	) name4264 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w4796_,
		_w4797_
	);
	LUT2 #(
		.INIT('h4)
	) name4265 (
		_w4795_,
		_w4797_,
		_w4798_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4266 (
		_w4770_,
		_w4778_,
		_w4793_,
		_w4798_,
		_w4799_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4267 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w4800_
	);
	LUT2 #(
		.INIT('h1)
	) name4268 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w4801_
	);
	LUT4 #(
		.INIT('h0010)
	) name4269 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4802_
	);
	LUT4 #(
		.INIT('h00c8)
	) name4270 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		_w4802_,
		_w4800_,
		_w4803_
	);
	LUT4 #(
		.INIT('h0001)
	) name4271 (
		_w4763_,
		_w4728_,
		_w4799_,
		_w4803_,
		_w4804_
	);
	LUT2 #(
		.INIT('h9)
	) name4272 (
		_w4691_,
		_w4804_,
		_w4805_
	);
	LUT4 #(
		.INIT('h0010)
	) name4273 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4806_
	);
	LUT4 #(
		.INIT('h0040)
	) name4274 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4807_
	);
	LUT3 #(
		.INIT('h20)
	) name4275 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4808_
	);
	LUT4 #(
		.INIT('h5554)
	) name4276 (
		\sa12_reg[2]/P0001 ,
		_w4807_,
		_w4808_,
		_w4806_,
		_w4809_
	);
	LUT3 #(
		.INIT('h80)
	) name4277 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4810_
	);
	LUT4 #(
		.INIT('h0080)
	) name4278 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4811_
	);
	LUT3 #(
		.INIT('ha8)
	) name4279 (
		\sa12_reg[2]/P0001 ,
		_w4810_,
		_w4811_,
		_w4812_
	);
	LUT4 #(
		.INIT('h1000)
	) name4280 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4813_
	);
	LUT2 #(
		.INIT('h4)
	) name4281 (
		\sa12_reg[7]/NET0131 ,
		_w4813_,
		_w4814_
	);
	LUT4 #(
		.INIT('h8000)
	) name4282 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4815_
	);
	LUT4 #(
		.INIT('h0002)
	) name4283 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4816_
	);
	LUT4 #(
		.INIT('h0400)
	) name4284 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4817_
	);
	LUT4 #(
		.INIT('h0001)
	) name4285 (
		_w4670_,
		_w4815_,
		_w4816_,
		_w4817_,
		_w4818_
	);
	LUT4 #(
		.INIT('h0100)
	) name4286 (
		_w4809_,
		_w4812_,
		_w4814_,
		_w4818_,
		_w4819_
	);
	LUT2 #(
		.INIT('h2)
	) name4287 (
		\sa12_reg[1]/P0001 ,
		_w4819_,
		_w4820_
	);
	LUT3 #(
		.INIT('h04)
	) name4288 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4821_
	);
	LUT4 #(
		.INIT('h0010)
	) name4289 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4822_
	);
	LUT3 #(
		.INIT('h01)
	) name4290 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4823_
	);
	LUT3 #(
		.INIT('h54)
	) name4291 (
		_w4623_,
		_w4822_,
		_w4823_,
		_w4824_
	);
	LUT3 #(
		.INIT('h01)
	) name4292 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4825_
	);
	LUT2 #(
		.INIT('h1)
	) name4293 (
		_w4815_,
		_w4825_,
		_w4826_
	);
	LUT3 #(
		.INIT('h8a)
	) name4294 (
		\sa12_reg[2]/P0001 ,
		_w4824_,
		_w4826_,
		_w4827_
	);
	LUT4 #(
		.INIT('h0008)
	) name4295 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4828_
	);
	LUT3 #(
		.INIT('h10)
	) name4296 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4829_
	);
	LUT4 #(
		.INIT('h0400)
	) name4297 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4830_
	);
	LUT3 #(
		.INIT('h54)
	) name4298 (
		\sa12_reg[5]/P0001 ,
		_w4828_,
		_w4830_,
		_w4831_
	);
	LUT2 #(
		.INIT('h4)
	) name4299 (
		\sa12_reg[3]/P0001 ,
		_w4641_,
		_w4832_
	);
	LUT4 #(
		.INIT('h8acf)
	) name4300 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4675_,
		_w4641_,
		_w4833_
	);
	LUT3 #(
		.INIT('h45)
	) name4301 (
		\sa12_reg[1]/P0001 ,
		_w4831_,
		_w4833_,
		_w4834_
	);
	LUT4 #(
		.INIT('h1000)
	) name4302 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4835_
	);
	LUT3 #(
		.INIT('h54)
	) name4303 (
		\sa12_reg[2]/P0001 ,
		_w4650_,
		_w4835_,
		_w4836_
	);
	LUT4 #(
		.INIT('h0001)
	) name4304 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4837_
	);
	LUT3 #(
		.INIT('h0b)
	) name4305 (
		\sa12_reg[2]/P0001 ,
		_w4603_,
		_w4837_,
		_w4838_
	);
	LUT2 #(
		.INIT('h4)
	) name4306 (
		_w4836_,
		_w4838_,
		_w4839_
	);
	LUT3 #(
		.INIT('h10)
	) name4307 (
		_w4834_,
		_w4827_,
		_w4839_,
		_w4840_
	);
	LUT3 #(
		.INIT('h45)
	) name4308 (
		\sa12_reg[0]/P0001 ,
		_w4820_,
		_w4840_,
		_w4841_
	);
	LUT4 #(
		.INIT('h0008)
	) name4309 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4842_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4310 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4843_
	);
	LUT2 #(
		.INIT('h4)
	) name4311 (
		_w4842_,
		_w4843_,
		_w4844_
	);
	LUT3 #(
		.INIT('h01)
	) name4312 (
		\sa12_reg[2]/P0001 ,
		_w4618_,
		_w4633_,
		_w4845_
	);
	LUT4 #(
		.INIT('h8000)
	) name4313 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4846_
	);
	LUT3 #(
		.INIT('h23)
	) name4314 (
		\sa12_reg[3]/P0001 ,
		_w4661_,
		_w4846_,
		_w4847_
	);
	LUT4 #(
		.INIT('h0155)
	) name4315 (
		\sa12_reg[1]/P0001 ,
		_w4844_,
		_w4845_,
		_w4847_,
		_w4848_
	);
	LUT3 #(
		.INIT('h08)
	) name4316 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4849_
	);
	LUT4 #(
		.INIT('h1d3f)
	) name4317 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4807_,
		_w4849_,
		_w4850_
	);
	LUT4 #(
		.INIT('h0200)
	) name4318 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4851_
	);
	LUT3 #(
		.INIT('h07)
	) name4319 (
		_w4595_,
		_w4596_,
		_w4851_,
		_w4852_
	);
	LUT3 #(
		.INIT('h2a)
	) name4320 (
		\sa12_reg[1]/P0001 ,
		_w4850_,
		_w4852_,
		_w4853_
	);
	LUT3 #(
		.INIT('h04)
	) name4321 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4854_
	);
	LUT4 #(
		.INIT('h5554)
	) name4322 (
		\sa12_reg[2]/P0001 ,
		_w4661_,
		_w4626_,
		_w4854_,
		_w4855_
	);
	LUT3 #(
		.INIT('hd0)
	) name4323 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		_w4856_
	);
	LUT2 #(
		.INIT('h2)
	) name4324 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[2]/P0001 ,
		_w4857_
	);
	LUT4 #(
		.INIT('h0222)
	) name4325 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4858_
	);
	LUT3 #(
		.INIT('h10)
	) name4326 (
		_w4651_,
		_w4856_,
		_w4858_,
		_w4859_
	);
	LUT3 #(
		.INIT('h02)
	) name4327 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4860_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name4328 (
		\sa12_reg[7]/NET0131 ,
		_w4668_,
		_w4821_,
		_w4860_,
		_w4861_
	);
	LUT3 #(
		.INIT('h20)
	) name4329 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4862_
	);
	LUT4 #(
		.INIT('h2000)
	) name4330 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4863_
	);
	LUT4 #(
		.INIT('h2a7f)
	) name4331 (
		\sa12_reg[2]/P0001 ,
		_w4595_,
		_w4615_,
		_w4863_,
		_w4864_
	);
	LUT4 #(
		.INIT('h1000)
	) name4332 (
		_w4855_,
		_w4859_,
		_w4861_,
		_w4864_,
		_w4865_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4333 (
		\sa12_reg[0]/P0001 ,
		_w4848_,
		_w4853_,
		_w4865_,
		_w4866_
	);
	LUT4 #(
		.INIT('hee7f)
	) name4334 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4867_
	);
	LUT4 #(
		.INIT('h5054)
	) name4335 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[5]/P0001 ,
		_w4863_,
		_w4867_,
		_w4868_
	);
	LUT3 #(
		.INIT('h6b)
	) name4336 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4869_
	);
	LUT2 #(
		.INIT('h2)
	) name4337 (
		_w4862_,
		_w4869_,
		_w4870_
	);
	LUT3 #(
		.INIT('h80)
	) name4338 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4871_
	);
	LUT4 #(
		.INIT('h0001)
	) name4339 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4872_
	);
	LUT3 #(
		.INIT('h07)
	) name4340 (
		_w4659_,
		_w4871_,
		_w4872_,
		_w4873_
	);
	LUT4 #(
		.INIT('h5455)
	) name4341 (
		\sa12_reg[1]/P0001 ,
		_w4868_,
		_w4870_,
		_w4873_,
		_w4874_
	);
	LUT4 #(
		.INIT('h0040)
	) name4342 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4875_
	);
	LUT3 #(
		.INIT('h80)
	) name4343 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4875_,
		_w4876_
	);
	LUT3 #(
		.INIT('h02)
	) name4344 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4877_
	);
	LUT2 #(
		.INIT('h1)
	) name4345 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4878_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name4346 (
		\sa12_reg[2]/P0001 ,
		_w4603_,
		_w4877_,
		_w4878_,
		_w4879_
	);
	LUT3 #(
		.INIT('h8a)
	) name4347 (
		\sa12_reg[1]/P0001 ,
		_w4876_,
		_w4879_,
		_w4880_
	);
	LUT4 #(
		.INIT('h0008)
	) name4348 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4881_
	);
	LUT2 #(
		.INIT('h8)
	) name4349 (
		_w4684_,
		_w4881_,
		_w4882_
	);
	LUT4 #(
		.INIT('h5450)
	) name4350 (
		\sa12_reg[2]/P0001 ,
		_w4591_,
		_w4670_,
		_w4593_,
		_w4883_
	);
	LUT2 #(
		.INIT('h1)
	) name4351 (
		_w4882_,
		_w4883_,
		_w4884_
	);
	LUT3 #(
		.INIT('h10)
	) name4352 (
		_w4874_,
		_w4880_,
		_w4884_,
		_w4885_
	);
	LUT2 #(
		.INIT('h4)
	) name4353 (
		_w4866_,
		_w4885_,
		_w4886_
	);
	LUT3 #(
		.INIT('h04)
	) name4354 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4887_
	);
	LUT4 #(
		.INIT('h0010)
	) name4355 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4888_
	);
	LUT2 #(
		.INIT('h2)
	) name4356 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4889_
	);
	LUT3 #(
		.INIT('h04)
	) name4357 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4890_
	);
	LUT4 #(
		.INIT('h0040)
	) name4358 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4891_
	);
	LUT3 #(
		.INIT('h20)
	) name4359 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4892_
	);
	LUT4 #(
		.INIT('h5554)
	) name4360 (
		\sa23_reg[2]/P0001 ,
		_w4891_,
		_w4892_,
		_w4888_,
		_w4893_
	);
	LUT2 #(
		.INIT('h8)
	) name4361 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4894_
	);
	LUT3 #(
		.INIT('h80)
	) name4362 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4895_
	);
	LUT2 #(
		.INIT('h8)
	) name4363 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4896_
	);
	LUT3 #(
		.INIT('h80)
	) name4364 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4897_
	);
	LUT4 #(
		.INIT('h0080)
	) name4365 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4898_
	);
	LUT3 #(
		.INIT('ha8)
	) name4366 (
		\sa23_reg[2]/P0001 ,
		_w4895_,
		_w4898_,
		_w4899_
	);
	LUT2 #(
		.INIT('h1)
	) name4367 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w4900_
	);
	LUT3 #(
		.INIT('h01)
	) name4368 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4901_
	);
	LUT2 #(
		.INIT('h8)
	) name4369 (
		_w4896_,
		_w4901_,
		_w4902_
	);
	LUT2 #(
		.INIT('h4)
	) name4370 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4903_
	);
	LUT4 #(
		.INIT('h0400)
	) name4371 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4904_
	);
	LUT2 #(
		.INIT('h4)
	) name4372 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4905_
	);
	LUT4 #(
		.INIT('h1000)
	) name4373 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4906_
	);
	LUT2 #(
		.INIT('h1)
	) name4374 (
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4907_
	);
	LUT2 #(
		.INIT('h2)
	) name4375 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		_w4908_
	);
	LUT4 #(
		.INIT('h0002)
	) name4376 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4909_
	);
	LUT2 #(
		.INIT('h8)
	) name4377 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w4910_
	);
	LUT4 #(
		.INIT('h8000)
	) name4378 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4911_
	);
	LUT4 #(
		.INIT('h0001)
	) name4379 (
		_w4904_,
		_w4906_,
		_w4909_,
		_w4911_,
		_w4912_
	);
	LUT4 #(
		.INIT('h0100)
	) name4380 (
		_w4893_,
		_w4902_,
		_w4899_,
		_w4912_,
		_w4913_
	);
	LUT3 #(
		.INIT('h10)
	) name4381 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4914_
	);
	LUT4 #(
		.INIT('h0400)
	) name4382 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4915_
	);
	LUT4 #(
		.INIT('h0002)
	) name4383 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4916_
	);
	LUT3 #(
		.INIT('h54)
	) name4384 (
		\sa23_reg[5]/P0001 ,
		_w4915_,
		_w4916_,
		_w4917_
	);
	LUT2 #(
		.INIT('h8)
	) name4385 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		_w4918_
	);
	LUT2 #(
		.INIT('h1)
	) name4386 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4919_
	);
	LUT3 #(
		.INIT('h01)
	) name4387 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4920_
	);
	LUT4 #(
		.INIT('h4000)
	) name4388 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4921_
	);
	LUT4 #(
		.INIT('h4c7f)
	) name4389 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		_w4920_,
		_w4921_,
		_w4922_
	);
	LUT2 #(
		.INIT('h4)
	) name4390 (
		_w4917_,
		_w4922_,
		_w4923_
	);
	LUT2 #(
		.INIT('h1)
	) name4391 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4924_
	);
	LUT2 #(
		.INIT('h2)
	) name4392 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w4925_
	);
	LUT2 #(
		.INIT('h4)
	) name4393 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w4926_
	);
	LUT3 #(
		.INIT('h40)
	) name4394 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4927_
	);
	LUT3 #(
		.INIT('h9d)
	) name4395 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4928_
	);
	LUT2 #(
		.INIT('h1)
	) name4396 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4929_
	);
	LUT3 #(
		.INIT('h01)
	) name4397 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4930_
	);
	LUT4 #(
		.INIT('h0051)
	) name4398 (
		_w4911_,
		_w4924_,
		_w4928_,
		_w4930_,
		_w4931_
	);
	LUT2 #(
		.INIT('h4)
	) name4399 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4932_
	);
	LUT4 #(
		.INIT('h1000)
	) name4400 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4933_
	);
	LUT4 #(
		.INIT('h0008)
	) name4401 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4934_
	);
	LUT2 #(
		.INIT('h1)
	) name4402 (
		_w4933_,
		_w4934_,
		_w4935_
	);
	LUT4 #(
		.INIT('h0001)
	) name4403 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4936_
	);
	LUT2 #(
		.INIT('h8)
	) name4404 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4937_
	);
	LUT4 #(
		.INIT('h0800)
	) name4405 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4938_
	);
	LUT3 #(
		.INIT('h23)
	) name4406 (
		\sa23_reg[2]/P0001 ,
		_w4936_,
		_w4938_,
		_w4939_
	);
	LUT4 #(
		.INIT('he400)
	) name4407 (
		\sa23_reg[2]/P0001 ,
		_w4935_,
		_w4931_,
		_w4939_,
		_w4940_
	);
	LUT4 #(
		.INIT('hd800)
	) name4408 (
		\sa23_reg[1]/P0001 ,
		_w4913_,
		_w4923_,
		_w4940_,
		_w4941_
	);
	LUT2 #(
		.INIT('h1)
	) name4409 (
		\sa23_reg[0]/P0001 ,
		_w4941_,
		_w4942_
	);
	LUT3 #(
		.INIT('h10)
	) name4410 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4943_
	);
	LUT2 #(
		.INIT('h2)
	) name4411 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4944_
	);
	LUT2 #(
		.INIT('h2)
	) name4412 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4945_
	);
	LUT4 #(
		.INIT('h0008)
	) name4413 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4946_
	);
	LUT3 #(
		.INIT('ha8)
	) name4414 (
		\sa23_reg[2]/P0001 ,
		_w4943_,
		_w4946_,
		_w4947_
	);
	LUT3 #(
		.INIT('h08)
	) name4415 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4948_
	);
	LUT4 #(
		.INIT('h0200)
	) name4416 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4949_
	);
	LUT4 #(
		.INIT('hfd3f)
	) name4417 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4950_
	);
	LUT2 #(
		.INIT('h2)
	) name4418 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4951_
	);
	LUT3 #(
		.INIT('h08)
	) name4419 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4952_
	);
	LUT4 #(
		.INIT('h4000)
	) name4420 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4953_
	);
	LUT4 #(
		.INIT('hbf5f)
	) name4421 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4954_
	);
	LUT4 #(
		.INIT('hfa32)
	) name4422 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4950_,
		_w4954_,
		_w4955_
	);
	LUT3 #(
		.INIT('h45)
	) name4423 (
		\sa23_reg[1]/P0001 ,
		_w4947_,
		_w4955_,
		_w4956_
	);
	LUT3 #(
		.INIT('h02)
	) name4424 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4957_
	);
	LUT4 #(
		.INIT('h135f)
	) name4425 (
		_w4890_,
		_w4910_,
		_w4937_,
		_w4957_,
		_w4958_
	);
	LUT3 #(
		.INIT('h04)
	) name4426 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4959_
	);
	LUT2 #(
		.INIT('h8)
	) name4427 (
		_w4919_,
		_w4959_,
		_w4960_
	);
	LUT4 #(
		.INIT('h0200)
	) name4428 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4961_
	);
	LUT3 #(
		.INIT('h07)
	) name4429 (
		_w4919_,
		_w4959_,
		_w4961_,
		_w4962_
	);
	LUT3 #(
		.INIT('h2a)
	) name4430 (
		\sa23_reg[1]/P0001 ,
		_w4958_,
		_w4962_,
		_w4963_
	);
	LUT3 #(
		.INIT('h10)
	) name4431 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4964_
	);
	LUT2 #(
		.INIT('h8)
	) name4432 (
		_w4929_,
		_w4964_,
		_w4965_
	);
	LUT4 #(
		.INIT('h0777)
	) name4433 (
		_w4894_,
		_w4927_,
		_w4929_,
		_w4964_,
		_w4966_
	);
	LUT4 #(
		.INIT('h2000)
	) name4434 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4967_
	);
	LUT4 #(
		.INIT('h23af)
	) name4435 (
		\sa23_reg[2]/P0001 ,
		_w4925_,
		_w4967_,
		_w4948_,
		_w4968_
	);
	LUT3 #(
		.INIT('hd0)
	) name4436 (
		\sa23_reg[2]/P0001 ,
		_w4966_,
		_w4968_,
		_w4969_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4437 (
		\sa23_reg[0]/P0001 ,
		_w4956_,
		_w4963_,
		_w4969_,
		_w4970_
	);
	LUT3 #(
		.INIT('h20)
	) name4438 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		_w4971_
	);
	LUT3 #(
		.INIT('h23)
	) name4439 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4972_
	);
	LUT4 #(
		.INIT('h0123)
	) name4440 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4973_
	);
	LUT3 #(
		.INIT('ha8)
	) name4441 (
		\sa23_reg[1]/P0001 ,
		_w4971_,
		_w4973_,
		_w4974_
	);
	LUT2 #(
		.INIT('h8)
	) name4442 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4975_
	);
	LUT4 #(
		.INIT('h0080)
	) name4443 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4976_
	);
	LUT4 #(
		.INIT('h0020)
	) name4444 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4977_
	);
	LUT3 #(
		.INIT('h04)
	) name4445 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4978_
	);
	LUT3 #(
		.INIT('h01)
	) name4446 (
		_w4976_,
		_w4977_,
		_w4978_,
		_w4979_
	);
	LUT3 #(
		.INIT('h8a)
	) name4447 (
		\sa23_reg[0]/P0001 ,
		_w4974_,
		_w4979_,
		_w4980_
	);
	LUT3 #(
		.INIT('h10)
	) name4448 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w4981_
	);
	LUT4 #(
		.INIT('h0080)
	) name4449 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4982_
	);
	LUT4 #(
		.INIT('hee7f)
	) name4450 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4983_
	);
	LUT4 #(
		.INIT('h5054)
	) name4451 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[5]/P0001 ,
		_w4967_,
		_w4983_,
		_w4984_
	);
	LUT3 #(
		.INIT('h15)
	) name4452 (
		_w4906_,
		_w4907_,
		_w4971_,
		_w4985_
	);
	LUT2 #(
		.INIT('h4)
	) name4453 (
		_w4984_,
		_w4985_,
		_w4986_
	);
	LUT3 #(
		.INIT('h45)
	) name4454 (
		\sa23_reg[2]/P0001 ,
		_w4980_,
		_w4986_,
		_w4987_
	);
	LUT3 #(
		.INIT('h04)
	) name4455 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4988_
	);
	LUT3 #(
		.INIT('h6b)
	) name4456 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4989_
	);
	LUT3 #(
		.INIT('h20)
	) name4457 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w4990_
	);
	LUT2 #(
		.INIT('h4)
	) name4458 (
		_w4989_,
		_w4990_,
		_w4991_
	);
	LUT2 #(
		.INIT('h2)
	) name4459 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4992_
	);
	LUT3 #(
		.INIT('h80)
	) name4460 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		_w4993_
	);
	LUT4 #(
		.INIT('h0001)
	) name4461 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4994_
	);
	LUT3 #(
		.INIT('h07)
	) name4462 (
		_w4992_,
		_w4993_,
		_w4994_,
		_w4995_
	);
	LUT3 #(
		.INIT('h45)
	) name4463 (
		\sa23_reg[1]/P0001 ,
		_w4991_,
		_w4995_,
		_w4996_
	);
	LUT4 #(
		.INIT('h0008)
	) name4464 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w4997_
	);
	LUT2 #(
		.INIT('h8)
	) name4465 (
		_w4918_,
		_w4997_,
		_w4998_
	);
	LUT2 #(
		.INIT('h8)
	) name4466 (
		_w4908_,
		_w4930_,
		_w4999_
	);
	LUT4 #(
		.INIT('h1bbb)
	) name4467 (
		\sa23_reg[2]/P0001 ,
		_w4938_,
		_w4926_,
		_w4948_,
		_w5000_
	);
	LUT4 #(
		.INIT('h1311)
	) name4468 (
		\sa23_reg[1]/P0001 ,
		_w4998_,
		_w4999_,
		_w5000_,
		_w5001_
	);
	LUT2 #(
		.INIT('h4)
	) name4469 (
		_w4996_,
		_w5001_,
		_w5002_
	);
	LUT3 #(
		.INIT('h10)
	) name4470 (
		_w4987_,
		_w4970_,
		_w5002_,
		_w5003_
	);
	LUT4 #(
		.INIT('hb4bb)
	) name4471 (
		_w4841_,
		_w4886_,
		_w4942_,
		_w5003_,
		_w5004_
	);
	LUT2 #(
		.INIT('h8)
	) name4472 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5005_
	);
	LUT3 #(
		.INIT('h08)
	) name4473 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5006_
	);
	LUT2 #(
		.INIT('h4)
	) name4474 (
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5007_
	);
	LUT4 #(
		.INIT('h0200)
	) name4475 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5008_
	);
	LUT4 #(
		.INIT('hfd3f)
	) name4476 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5009_
	);
	LUT2 #(
		.INIT('h1)
	) name4477 (
		\sa30_reg[2]/P0001 ,
		_w5009_,
		_w5010_
	);
	LUT2 #(
		.INIT('h8)
	) name4478 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w5011_
	);
	LUT2 #(
		.INIT('h1)
	) name4479 (
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5012_
	);
	LUT4 #(
		.INIT('h0008)
	) name4480 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5013_
	);
	LUT2 #(
		.INIT('h4)
	) name4481 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5014_
	);
	LUT3 #(
		.INIT('h10)
	) name4482 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5015_
	);
	LUT3 #(
		.INIT('ha8)
	) name4483 (
		\sa30_reg[2]/P0001 ,
		_w5013_,
		_w5015_,
		_w5016_
	);
	LUT2 #(
		.INIT('h2)
	) name4484 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5017_
	);
	LUT2 #(
		.INIT('h8)
	) name4485 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5018_
	);
	LUT4 #(
		.INIT('h0080)
	) name4486 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5019_
	);
	LUT2 #(
		.INIT('h8)
	) name4487 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5020_
	);
	LUT2 #(
		.INIT('h4)
	) name4488 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w5021_
	);
	LUT3 #(
		.INIT('h40)
	) name4489 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5022_
	);
	LUT3 #(
		.INIT('h07)
	) name4490 (
		_w5020_,
		_w5022_,
		_w5019_,
		_w5023_
	);
	LUT4 #(
		.INIT('h5455)
	) name4491 (
		\sa30_reg[1]/P0001 ,
		_w5016_,
		_w5010_,
		_w5023_,
		_w5024_
	);
	LUT4 #(
		.INIT('h0080)
	) name4492 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5025_
	);
	LUT3 #(
		.INIT('h20)
	) name4493 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5026_
	);
	LUT4 #(
		.INIT('h0200)
	) name4494 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5027_
	);
	LUT3 #(
		.INIT('h0b)
	) name4495 (
		\sa30_reg[6]/NET0131 ,
		_w5025_,
		_w5027_,
		_w5028_
	);
	LUT2 #(
		.INIT('h1)
	) name4496 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5029_
	);
	LUT3 #(
		.INIT('h04)
	) name4497 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5030_
	);
	LUT4 #(
		.INIT('h4000)
	) name4498 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5031_
	);
	LUT2 #(
		.INIT('h4)
	) name4499 (
		\sa30_reg[6]/NET0131 ,
		_w5031_,
		_w5032_
	);
	LUT4 #(
		.INIT('hdeff)
	) name4500 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5021_,
		_w5033_
	);
	LUT3 #(
		.INIT('h2a)
	) name4501 (
		\sa30_reg[1]/P0001 ,
		_w5028_,
		_w5033_,
		_w5034_
	);
	LUT3 #(
		.INIT('h04)
	) name4502 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5035_
	);
	LUT2 #(
		.INIT('h2)
	) name4503 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w5036_
	);
	LUT4 #(
		.INIT('h0020)
	) name4504 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5037_
	);
	LUT4 #(
		.INIT('h5554)
	) name4505 (
		\sa30_reg[2]/P0001 ,
		_w5035_,
		_w5019_,
		_w5037_,
		_w5038_
	);
	LUT2 #(
		.INIT('h8)
	) name4506 (
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5039_
	);
	LUT3 #(
		.INIT('h40)
	) name4507 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5040_
	);
	LUT2 #(
		.INIT('h4)
	) name4508 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w5041_
	);
	LUT4 #(
		.INIT('h135f)
	) name4509 (
		_w5006_,
		_w5040_,
		_w5036_,
		_w5041_,
		_w5042_
	);
	LUT2 #(
		.INIT('h4)
	) name4510 (
		_w5038_,
		_w5042_,
		_w5043_
	);
	LUT2 #(
		.INIT('h1)
	) name4511 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5044_
	);
	LUT2 #(
		.INIT('h4)
	) name4512 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5045_
	);
	LUT4 #(
		.INIT('h0010)
	) name4513 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5046_
	);
	LUT2 #(
		.INIT('h4)
	) name4514 (
		\sa30_reg[3]/P0001 ,
		_w5046_,
		_w5047_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name4515 (
		\sa30_reg[3]/P0001 ,
		_w5020_,
		_w5022_,
		_w5046_,
		_w5048_
	);
	LUT2 #(
		.INIT('h2)
	) name4516 (
		\sa30_reg[1]/P0001 ,
		\sa30_reg[2]/P0001 ,
		_w5049_
	);
	LUT3 #(
		.INIT('h01)
	) name4517 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5050_
	);
	LUT3 #(
		.INIT('h20)
	) name4518 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		_w5051_
	);
	LUT4 #(
		.INIT('hdfd3)
	) name4519 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5052_
	);
	LUT3 #(
		.INIT('h8a)
	) name4520 (
		_w5049_,
		_w5050_,
		_w5052_,
		_w5053_
	);
	LUT3 #(
		.INIT('h0d)
	) name4521 (
		\sa30_reg[2]/P0001 ,
		_w5048_,
		_w5053_,
		_w5054_
	);
	LUT4 #(
		.INIT('h1000)
	) name4522 (
		_w5034_,
		_w5024_,
		_w5043_,
		_w5054_,
		_w5055_
	);
	LUT2 #(
		.INIT('h2)
	) name4523 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5056_
	);
	LUT4 #(
		.INIT('hf7a7)
	) name4524 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5057_
	);
	LUT4 #(
		.INIT('h4051)
	) name4525 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		_w5007_,
		_w5057_,
		_w5058_
	);
	LUT3 #(
		.INIT('h80)
	) name4526 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5059_
	);
	LUT4 #(
		.INIT('h0080)
	) name4527 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5060_
	);
	LUT3 #(
		.INIT('ha8)
	) name4528 (
		\sa30_reg[2]/P0001 ,
		_w5059_,
		_w5060_,
		_w5061_
	);
	LUT3 #(
		.INIT('h20)
	) name4529 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5062_
	);
	LUT4 #(
		.INIT('h0400)
	) name4530 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5063_
	);
	LUT4 #(
		.INIT('h8000)
	) name4531 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5064_
	);
	LUT4 #(
		.INIT('h0002)
	) name4532 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5065_
	);
	LUT3 #(
		.INIT('h01)
	) name4533 (
		_w5063_,
		_w5064_,
		_w5065_,
		_w5066_
	);
	LUT2 #(
		.INIT('h1)
	) name4534 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w5067_
	);
	LUT4 #(
		.INIT('h1000)
	) name4535 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5068_
	);
	LUT4 #(
		.INIT('h1000)
	) name4536 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5069_
	);
	LUT3 #(
		.INIT('h0b)
	) name4537 (
		\sa30_reg[7]/P0001 ,
		_w5068_,
		_w5069_,
		_w5070_
	);
	LUT4 #(
		.INIT('h1000)
	) name4538 (
		_w5058_,
		_w5061_,
		_w5066_,
		_w5070_,
		_w5071_
	);
	LUT3 #(
		.INIT('h10)
	) name4539 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5072_
	);
	LUT2 #(
		.INIT('h8)
	) name4540 (
		_w5005_,
		_w5072_,
		_w5073_
	);
	LUT3 #(
		.INIT('h02)
	) name4541 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5074_
	);
	LUT4 #(
		.INIT('h0400)
	) name4542 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5075_
	);
	LUT3 #(
		.INIT('h01)
	) name4543 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5076_
	);
	LUT4 #(
		.INIT('hf9f8)
	) name4544 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5077_
	);
	LUT2 #(
		.INIT('h1)
	) name4545 (
		\sa30_reg[2]/P0001 ,
		_w5075_,
		_w5078_
	);
	LUT4 #(
		.INIT('h0032)
	) name4546 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[5]/P0001 ,
		_w5075_,
		_w5077_,
		_w5079_
	);
	LUT2 #(
		.INIT('h1)
	) name4547 (
		_w5073_,
		_w5079_,
		_w5080_
	);
	LUT3 #(
		.INIT('h9d)
	) name4548 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5081_
	);
	LUT3 #(
		.INIT('h01)
	) name4549 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5082_
	);
	LUT4 #(
		.INIT('h1101)
	) name4550 (
		_w5064_,
		_w5082_,
		_w5044_,
		_w5081_,
		_w5083_
	);
	LUT4 #(
		.INIT('h1000)
	) name4551 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5084_
	);
	LUT4 #(
		.INIT('h0008)
	) name4552 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5085_
	);
	LUT2 #(
		.INIT('h1)
	) name4553 (
		_w5084_,
		_w5085_,
		_w5086_
	);
	LUT3 #(
		.INIT('h54)
	) name4554 (
		\sa30_reg[2]/P0001 ,
		_w5084_,
		_w5085_,
		_w5087_
	);
	LUT2 #(
		.INIT('h8)
	) name4555 (
		_w5062_,
		_w5041_,
		_w5088_
	);
	LUT3 #(
		.INIT('h01)
	) name4556 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5089_
	);
	LUT4 #(
		.INIT('h0001)
	) name4557 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5090_
	);
	LUT3 #(
		.INIT('h07)
	) name4558 (
		_w5062_,
		_w5041_,
		_w5090_,
		_w5091_
	);
	LUT4 #(
		.INIT('hd800)
	) name4559 (
		\sa30_reg[2]/P0001 ,
		_w5083_,
		_w5086_,
		_w5091_,
		_w5092_
	);
	LUT4 #(
		.INIT('hd800)
	) name4560 (
		\sa30_reg[1]/P0001 ,
		_w5071_,
		_w5080_,
		_w5092_,
		_w5093_
	);
	LUT4 #(
		.INIT('h2000)
	) name4561 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5094_
	);
	LUT4 #(
		.INIT('h8000)
	) name4562 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5095_
	);
	LUT4 #(
		.INIT('h1000)
	) name4563 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5096_
	);
	LUT4 #(
		.INIT('h000b)
	) name4564 (
		\sa30_reg[7]/P0001 ,
		_w5095_,
		_w5094_,
		_w5096_,
		_w5097_
	);
	LUT4 #(
		.INIT('h0001)
	) name4565 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5098_
	);
	LUT3 #(
		.INIT('h10)
	) name4566 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5099_
	);
	LUT3 #(
		.INIT('h04)
	) name4567 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5100_
	);
	LUT4 #(
		.INIT('h1445)
	) name4568 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5101_
	);
	LUT2 #(
		.INIT('h8)
	) name4569 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w5102_
	);
	LUT3 #(
		.INIT('ha2)
	) name4570 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5103_
	);
	LUT4 #(
		.INIT('h5551)
	) name4571 (
		_w5098_,
		_w5102_,
		_w5103_,
		_w5101_,
		_w5104_
	);
	LUT4 #(
		.INIT('h0155)
	) name4572 (
		\sa30_reg[1]/P0001 ,
		\sa30_reg[2]/P0001 ,
		_w5097_,
		_w5104_,
		_w5105_
	);
	LUT3 #(
		.INIT('h02)
	) name4573 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5106_
	);
	LUT4 #(
		.INIT('h0002)
	) name4574 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5107_
	);
	LUT2 #(
		.INIT('h4)
	) name4575 (
		\sa30_reg[6]/NET0131 ,
		_w5107_,
		_w5108_
	);
	LUT3 #(
		.INIT('h04)
	) name4576 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5109_
	);
	LUT3 #(
		.INIT('h80)
	) name4577 (
		\sa30_reg[5]/P0001 ,
		_w5102_,
		_w5109_,
		_w5110_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4578 (
		\sa30_reg[1]/P0001 ,
		_w5088_,
		_w5110_,
		_w5108_,
		_w5111_
	);
	LUT2 #(
		.INIT('h8)
	) name4579 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		_w5112_
	);
	LUT3 #(
		.INIT('h02)
	) name4580 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5113_
	);
	LUT3 #(
		.INIT('h80)
	) name4581 (
		\sa30_reg[4]/P0001 ,
		_w5112_,
		_w5113_,
		_w5114_
	);
	LUT2 #(
		.INIT('h8)
	) name4582 (
		_w5074_,
		_w5017_,
		_w5115_
	);
	LUT3 #(
		.INIT('h40)
	) name4583 (
		\sa30_reg[2]/P0001 ,
		_w5074_,
		_w5017_,
		_w5116_
	);
	LUT2 #(
		.INIT('h1)
	) name4584 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		_w5117_
	);
	LUT2 #(
		.INIT('h8)
	) name4585 (
		_w5040_,
		_w5117_,
		_w5118_
	);
	LUT3 #(
		.INIT('h01)
	) name4586 (
		_w5116_,
		_w5118_,
		_w5114_,
		_w5119_
	);
	LUT3 #(
		.INIT('h10)
	) name4587 (
		_w5105_,
		_w5111_,
		_w5119_,
		_w5120_
	);
	LUT4 #(
		.INIT('he400)
	) name4588 (
		\sa30_reg[0]/P0002 ,
		_w5093_,
		_w5055_,
		_w5120_,
		_w5121_
	);
	LUT2 #(
		.INIT('h9)
	) name4589 (
		\u0_w_reg[1][29]/P0002 ,
		_w5121_,
		_w5122_
	);
	LUT4 #(
		.INIT('h1441)
	) name4590 (
		\ld_r_reg/P0001 ,
		_w4805_,
		_w5004_,
		_w5122_,
		_w5123_
	);
	LUT3 #(
		.INIT('h82)
	) name4591 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[93]/P0001 ,
		\u0_w_reg[1][29]/P0002 ,
		_w5124_
	);
	LUT2 #(
		.INIT('h1)
	) name4592 (
		_w5123_,
		_w5124_,
		_w5125_
	);
	LUT3 #(
		.INIT('h80)
	) name4593 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5126_
	);
	LUT3 #(
		.INIT('ha8)
	) name4594 (
		\sa30_reg[2]/P0001 ,
		_w5100_,
		_w5126_,
		_w5127_
	);
	LUT4 #(
		.INIT('h0004)
	) name4595 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5128_
	);
	LUT4 #(
		.INIT('h0800)
	) name4596 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5129_
	);
	LUT3 #(
		.INIT('h0b)
	) name4597 (
		\sa30_reg[2]/P0001 ,
		_w5128_,
		_w5129_,
		_w5130_
	);
	LUT4 #(
		.INIT('h5455)
	) name4598 (
		\sa30_reg[1]/P0001 ,
		_w5087_,
		_w5127_,
		_w5130_,
		_w5131_
	);
	LUT4 #(
		.INIT('h0100)
	) name4599 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5132_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name4600 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5133_
	);
	LUT4 #(
		.INIT('h80aa)
	) name4601 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5132_,
		_w5133_,
		_w5134_
	);
	LUT4 #(
		.INIT('h2000)
	) name4602 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5135_
	);
	LUT3 #(
		.INIT('h0b)
	) name4603 (
		\sa30_reg[6]/NET0131 ,
		_w5025_,
		_w5135_,
		_w5136_
	);
	LUT3 #(
		.INIT('h01)
	) name4604 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		_w5137_
	);
	LUT2 #(
		.INIT('h4)
	) name4605 (
		_w5045_,
		_w5137_,
		_w5138_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4606 (
		\sa30_reg[1]/P0001 ,
		_w5136_,
		_w5138_,
		_w5134_,
		_w5139_
	);
	LUT4 #(
		.INIT('h0040)
	) name4607 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5140_
	);
	LUT4 #(
		.INIT('h0040)
	) name4608 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5141_
	);
	LUT3 #(
		.INIT('h54)
	) name4609 (
		\sa30_reg[2]/P0001 ,
		_w5140_,
		_w5141_,
		_w5142_
	);
	LUT3 #(
		.INIT('h08)
	) name4610 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5143_
	);
	LUT4 #(
		.INIT('h0080)
	) name4611 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5144_
	);
	LUT3 #(
		.INIT('h07)
	) name4612 (
		_w5020_,
		_w5022_,
		_w5144_,
		_w5145_
	);
	LUT2 #(
		.INIT('h1)
	) name4613 (
		_w5090_,
		_w5008_,
		_w5146_
	);
	LUT4 #(
		.INIT('h3111)
	) name4614 (
		\sa30_reg[2]/P0001 ,
		_w5142_,
		_w5145_,
		_w5146_,
		_w5147_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4615 (
		\sa30_reg[0]/P0002 ,
		_w5139_,
		_w5131_,
		_w5147_,
		_w5148_
	);
	LUT3 #(
		.INIT('he6)
	) name4616 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5149_
	);
	LUT2 #(
		.INIT('h2)
	) name4617 (
		_w5021_,
		_w5149_,
		_w5150_
	);
	LUT3 #(
		.INIT('h2a)
	) name4618 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5151_
	);
	LUT4 #(
		.INIT('h2220)
	) name4619 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5152_
	);
	LUT3 #(
		.INIT('h45)
	) name4620 (
		\sa30_reg[2]/P0001 ,
		_w5151_,
		_w5152_,
		_w5153_
	);
	LUT4 #(
		.INIT('h0001)
	) name4621 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5154_
	);
	LUT4 #(
		.INIT('h002a)
	) name4622 (
		\sa30_reg[2]/P0001 ,
		_w5040_,
		_w5021_,
		_w5154_,
		_w5155_
	);
	LUT3 #(
		.INIT('h0b)
	) name4623 (
		_w5150_,
		_w5153_,
		_w5155_,
		_w5156_
	);
	LUT4 #(
		.INIT('h0100)
	) name4624 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5157_
	);
	LUT4 #(
		.INIT('h0200)
	) name4625 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5158_
	);
	LUT4 #(
		.INIT('h0001)
	) name4626 (
		\sa30_reg[1]/P0001 ,
		_w5140_,
		_w5157_,
		_w5158_,
		_w5159_
	);
	LUT4 #(
		.INIT('h4000)
	) name4627 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5160_
	);
	LUT4 #(
		.INIT('h0777)
	) name4628 (
		_w5040_,
		_w5021_,
		_w5112_,
		_w5113_,
		_w5161_
	);
	LUT3 #(
		.INIT('h40)
	) name4629 (
		_w5160_,
		_w5159_,
		_w5161_,
		_w5162_
	);
	LUT2 #(
		.INIT('h4)
	) name4630 (
		\sa30_reg[2]/P0001 ,
		_w5090_,
		_w5163_
	);
	LUT2 #(
		.INIT('h2)
	) name4631 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		_w5164_
	);
	LUT3 #(
		.INIT('h80)
	) name4632 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5165_
	);
	LUT3 #(
		.INIT('h7e)
	) name4633 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5166_
	);
	LUT2 #(
		.INIT('h2)
	) name4634 (
		_w5164_,
		_w5166_,
		_w5167_
	);
	LUT3 #(
		.INIT('h8a)
	) name4635 (
		\sa30_reg[1]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5095_,
		_w5168_
	);
	LUT3 #(
		.INIT('h10)
	) name4636 (
		_w5167_,
		_w5163_,
		_w5168_,
		_w5169_
	);
	LUT4 #(
		.INIT('h4445)
	) name4637 (
		\sa30_reg[0]/P0002 ,
		_w5156_,
		_w5162_,
		_w5169_,
		_w5170_
	);
	LUT4 #(
		.INIT('h0020)
	) name4638 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5171_
	);
	LUT4 #(
		.INIT('h5504)
	) name4639 (
		\sa30_reg[2]/P0001 ,
		_w5062_,
		_w5067_,
		_w5171_,
		_w5172_
	);
	LUT4 #(
		.INIT('h0800)
	) name4640 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5173_
	);
	LUT2 #(
		.INIT('h1)
	) name4641 (
		_w5068_,
		_w5173_,
		_w5174_
	);
	LUT3 #(
		.INIT('h45)
	) name4642 (
		\sa30_reg[1]/P0001 ,
		_w5172_,
		_w5174_,
		_w5175_
	);
	LUT4 #(
		.INIT('h4000)
	) name4643 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5176_
	);
	LUT4 #(
		.INIT('h0002)
	) name4644 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5177_
	);
	LUT3 #(
		.INIT('h54)
	) name4645 (
		\sa30_reg[1]/P0001 ,
		_w5176_,
		_w5177_,
		_w5178_
	);
	LUT4 #(
		.INIT('h0001)
	) name4646 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5179_
	);
	LUT3 #(
		.INIT('h07)
	) name4647 (
		_w5011_,
		_w5100_,
		_w5179_,
		_w5180_
	);
	LUT3 #(
		.INIT('h8a)
	) name4648 (
		\sa30_reg[2]/P0001 ,
		_w5178_,
		_w5180_,
		_w5181_
	);
	LUT3 #(
		.INIT('h01)
	) name4649 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5182_
	);
	LUT4 #(
		.INIT('hdfe2)
	) name4650 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5183_
	);
	LUT2 #(
		.INIT('h8)
	) name4651 (
		\sa30_reg[1]/P0001 ,
		\sa30_reg[2]/P0001 ,
		_w5184_
	);
	LUT3 #(
		.INIT('h08)
	) name4652 (
		\sa30_reg[1]/P0001 ,
		\sa30_reg[2]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5185_
	);
	LUT2 #(
		.INIT('h4)
	) name4653 (
		_w5183_,
		_w5185_,
		_w5186_
	);
	LUT3 #(
		.INIT('h80)
	) name4654 (
		_w5074_,
		_w5017_,
		_w5049_,
		_w5187_
	);
	LUT2 #(
		.INIT('h4)
	) name4655 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		_w5188_
	);
	LUT2 #(
		.INIT('h8)
	) name4656 (
		_w5129_,
		_w5188_,
		_w5189_
	);
	LUT2 #(
		.INIT('h8)
	) name4657 (
		_w5029_,
		_w5182_,
		_w5190_
	);
	LUT4 #(
		.INIT('h153f)
	) name4658 (
		_w5029_,
		_w5129_,
		_w5188_,
		_w5182_,
		_w5191_
	);
	LUT3 #(
		.INIT('h10)
	) name4659 (
		_w5187_,
		_w5186_,
		_w5191_,
		_w5192_
	);
	LUT3 #(
		.INIT('h10)
	) name4660 (
		_w5181_,
		_w5175_,
		_w5192_,
		_w5193_
	);
	LUT3 #(
		.INIT('h10)
	) name4661 (
		_w5148_,
		_w5170_,
		_w5193_,
		_w5194_
	);
	LUT4 #(
		.INIT('h5655)
	) name4662 (
		\u0_w_reg[1][30]/P0001 ,
		_w5148_,
		_w5170_,
		_w5193_,
		_w5195_
	);
	LUT2 #(
		.INIT('h1)
	) name4663 (
		\sa12_reg[2]/P0001 ,
		_w4663_,
		_w5196_
	);
	LUT4 #(
		.INIT('hfad8)
	) name4664 (
		\sa12_reg[2]/P0001 ,
		_w4664_,
		_w4663_,
		_w4821_,
		_w5197_
	);
	LUT4 #(
		.INIT('h2223)
	) name4665 (
		\sa12_reg[2]/P0001 ,
		_w4603_,
		_w4650_,
		_w4835_,
		_w5198_
	);
	LUT3 #(
		.INIT('h45)
	) name4666 (
		\sa12_reg[1]/P0001 ,
		_w5197_,
		_w5198_,
		_w5199_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name4667 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5200_
	);
	LUT4 #(
		.INIT('h80aa)
	) name4668 (
		\sa12_reg[2]/P0001 ,
		_w4665_,
		_w4651_,
		_w5200_,
		_w5201_
	);
	LUT2 #(
		.INIT('h1)
	) name4669 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		_w5202_
	);
	LUT3 #(
		.INIT('h23)
	) name4670 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w5203_
	);
	LUT2 #(
		.INIT('h8)
	) name4671 (
		_w5202_,
		_w5203_,
		_w5204_
	);
	LUT4 #(
		.INIT('h2000)
	) name4672 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w5205_
	);
	LUT3 #(
		.INIT('h07)
	) name4673 (
		_w4591_,
		_w4849_,
		_w5205_,
		_w5206_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4674 (
		\sa12_reg[1]/P0001 ,
		_w5204_,
		_w5201_,
		_w5206_,
		_w5207_
	);
	LUT4 #(
		.INIT('h0040)
	) name4675 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5208_
	);
	LUT3 #(
		.INIT('h54)
	) name4676 (
		\sa12_reg[2]/P0001 ,
		_w4807_,
		_w5208_,
		_w5209_
	);
	LUT3 #(
		.INIT('h23)
	) name4677 (
		\sa12_reg[3]/P0001 ,
		_w4638_,
		_w4846_,
		_w5210_
	);
	LUT2 #(
		.INIT('h1)
	) name4678 (
		_w4618_,
		_w4837_,
		_w5211_
	);
	LUT4 #(
		.INIT('h3111)
	) name4679 (
		\sa12_reg[2]/P0001 ,
		_w5209_,
		_w5210_,
		_w5211_,
		_w5212_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4680 (
		\sa12_reg[0]/P0001 ,
		_w5207_,
		_w5199_,
		_w5212_,
		_w5213_
	);
	LUT3 #(
		.INIT('h7e)
	) name4681 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w5214_
	);
	LUT2 #(
		.INIT('h2)
	) name4682 (
		_w4635_,
		_w5214_,
		_w5215_
	);
	LUT2 #(
		.INIT('h8)
	) name4683 (
		_w4596_,
		_w4611_,
		_w5216_
	);
	LUT3 #(
		.INIT('h2a)
	) name4684 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4661_,
		_w5217_
	);
	LUT3 #(
		.INIT('h10)
	) name4685 (
		_w5215_,
		_w5216_,
		_w5217_,
		_w5218_
	);
	LUT4 #(
		.INIT('h4000)
	) name4686 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w5219_
	);
	LUT4 #(
		.INIT('h0001)
	) name4687 (
		\sa12_reg[1]/P0001 ,
		_w4679_,
		_w5208_,
		_w5219_,
		_w5220_
	);
	LUT4 #(
		.INIT('h0100)
	) name4688 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5221_
	);
	LUT4 #(
		.INIT('h153f)
	) name4689 (
		\sa12_reg[7]/NET0131 ,
		_w4654_,
		_w4684_,
		_w4648_,
		_w5222_
	);
	LUT3 #(
		.INIT('h40)
	) name4690 (
		_w5221_,
		_w5220_,
		_w5222_,
		_w5223_
	);
	LUT4 #(
		.INIT('h002a)
	) name4691 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4648_,
		_w4624_,
		_w5224_
	);
	LUT3 #(
		.INIT('h02)
	) name4692 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w5225_
	);
	LUT3 #(
		.INIT('h32)
	) name4693 (
		_w4676_,
		_w4637_,
		_w5225_,
		_w5226_
	);
	LUT4 #(
		.INIT('h0105)
	) name4694 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4621_,
		_w4875_,
		_w5227_
	);
	LUT3 #(
		.INIT('h45)
	) name4695 (
		_w5224_,
		_w5226_,
		_w5227_,
		_w5228_
	);
	LUT4 #(
		.INIT('h5501)
	) name4696 (
		\sa12_reg[0]/P0001 ,
		_w5218_,
		_w5223_,
		_w5228_,
		_w5229_
	);
	LUT4 #(
		.INIT('h0020)
	) name4697 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5230_
	);
	LUT4 #(
		.INIT('h5510)
	) name4698 (
		\sa12_reg[2]/P0001 ,
		_w4623_,
		_w4631_,
		_w5230_,
		_w5231_
	);
	LUT4 #(
		.INIT('h4000)
	) name4699 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5232_
	);
	LUT3 #(
		.INIT('ha8)
	) name4700 (
		\sa12_reg[2]/P0001 ,
		_w4640_,
		_w5232_,
		_w5233_
	);
	LUT4 #(
		.INIT('h0800)
	) name4701 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5234_
	);
	LUT2 #(
		.INIT('h1)
	) name4702 (
		_w4813_,
		_w5234_,
		_w5235_
	);
	LUT4 #(
		.INIT('h5455)
	) name4703 (
		\sa12_reg[1]/P0001 ,
		_w5233_,
		_w5231_,
		_w5235_,
		_w5236_
	);
	LUT2 #(
		.INIT('h8)
	) name4704 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[2]/P0001 ,
		_w5237_
	);
	LUT4 #(
		.INIT('h0800)
	) name4705 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5238_
	);
	LUT4 #(
		.INIT('h0002)
	) name4706 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5239_
	);
	LUT4 #(
		.INIT('h0207)
	) name4707 (
		\sa12_reg[4]/P0001 ,
		_w4596_,
		_w4872_,
		_w5238_,
		_w5240_
	);
	LUT2 #(
		.INIT('h2)
	) name4708 (
		_w5237_,
		_w5240_,
		_w5241_
	);
	LUT4 #(
		.INIT('h0020)
	) name4709 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5242_
	);
	LUT4 #(
		.INIT('h23af)
	) name4710 (
		\sa12_reg[7]/NET0131 ,
		_w4642_,
		_w4624_,
		_w5242_,
		_w5243_
	);
	LUT3 #(
		.INIT('h80)
	) name4711 (
		_w4591_,
		_w4593_,
		_w4857_,
		_w5244_
	);
	LUT2 #(
		.INIT('h8)
	) name4712 (
		_w4605_,
		_w4603_,
		_w5245_
	);
	LUT4 #(
		.INIT('h0100)
	) name4713 (
		_w4832_,
		_w5244_,
		_w5245_,
		_w5243_,
		_w5246_
	);
	LUT3 #(
		.INIT('h10)
	) name4714 (
		_w5241_,
		_w5236_,
		_w5246_,
		_w5247_
	);
	LUT3 #(
		.INIT('h10)
	) name4715 (
		_w5213_,
		_w5229_,
		_w5247_,
		_w5248_
	);
	LUT3 #(
		.INIT('h08)
	) name4716 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5249_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name4717 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5250_
	);
	LUT4 #(
		.INIT('h80aa)
	) name4718 (
		\sa23_reg[2]/P0001 ,
		_w4905_,
		_w4981_,
		_w5250_,
		_w5251_
	);
	LUT2 #(
		.INIT('h1)
	) name4719 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		_w5252_
	);
	LUT2 #(
		.INIT('h8)
	) name4720 (
		_w4972_,
		_w5252_,
		_w5253_
	);
	LUT4 #(
		.INIT('h2000)
	) name4721 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5254_
	);
	LUT3 #(
		.INIT('h07)
	) name4722 (
		_w4910_,
		_w4957_,
		_w5254_,
		_w5255_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4723 (
		\sa23_reg[1]/P0001 ,
		_w5251_,
		_w5253_,
		_w5255_,
		_w5256_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4724 (
		\sa23_reg[2]/P0001 ,
		_w4933_,
		_w4934_,
		_w4938_,
		_w5257_
	);
	LUT4 #(
		.INIT('h0004)
	) name4725 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5258_
	);
	LUT3 #(
		.INIT('h80)
	) name4726 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5259_
	);
	LUT4 #(
		.INIT('h0527)
	) name4727 (
		\sa23_reg[2]/P0001 ,
		_w4988_,
		_w5258_,
		_w5259_,
		_w5260_
	);
	LUT3 #(
		.INIT('h15)
	) name4728 (
		\sa23_reg[1]/P0001 ,
		_w5257_,
		_w5260_,
		_w5261_
	);
	LUT4 #(
		.INIT('h0040)
	) name4729 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5262_
	);
	LUT3 #(
		.INIT('h54)
	) name4730 (
		\sa23_reg[2]/P0001 ,
		_w4891_,
		_w5262_,
		_w5263_
	);
	LUT3 #(
		.INIT('h07)
	) name4731 (
		_w4894_,
		_w4927_,
		_w4982_,
		_w5264_
	);
	LUT2 #(
		.INIT('h1)
	) name4732 (
		_w4936_,
		_w4949_,
		_w5265_
	);
	LUT4 #(
		.INIT('h3111)
	) name4733 (
		\sa23_reg[2]/P0001 ,
		_w5263_,
		_w5264_,
		_w5265_,
		_w5266_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4734 (
		\sa23_reg[0]/P0001 ,
		_w5261_,
		_w5256_,
		_w5266_,
		_w5267_
	);
	LUT4 #(
		.INIT('h0200)
	) name4735 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5268_
	);
	LUT4 #(
		.INIT('h0100)
	) name4736 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5269_
	);
	LUT3 #(
		.INIT('h01)
	) name4737 (
		_w5262_,
		_w5269_,
		_w5268_,
		_w5270_
	);
	LUT2 #(
		.INIT('h8)
	) name4738 (
		_w4952_,
		_w4992_,
		_w5271_
	);
	LUT4 #(
		.INIT('h4000)
	) name4739 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5272_
	);
	LUT3 #(
		.INIT('h0b)
	) name4740 (
		\sa23_reg[3]/P0001 ,
		_w4967_,
		_w5272_,
		_w5273_
	);
	LUT4 #(
		.INIT('h4555)
	) name4741 (
		\sa23_reg[0]/P0001 ,
		_w5271_,
		_w5270_,
		_w5273_,
		_w5274_
	);
	LUT4 #(
		.INIT('h0002)
	) name4742 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5275_
	);
	LUT3 #(
		.INIT('h02)
	) name4743 (
		\sa23_reg[2]/P0001 ,
		_w4921_,
		_w5275_,
		_w5276_
	);
	LUT3 #(
		.INIT('h20)
	) name4744 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w5277_
	);
	LUT4 #(
		.INIT('h0020)
	) name4745 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5278_
	);
	LUT4 #(
		.INIT('h0800)
	) name4746 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5279_
	);
	LUT4 #(
		.INIT('h0001)
	) name4747 (
		\sa23_reg[2]/P0001 ,
		_w4938_,
		_w5278_,
		_w5279_,
		_w5280_
	);
	LUT4 #(
		.INIT('h1000)
	) name4748 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w5281_
	);
	LUT4 #(
		.INIT('h0800)
	) name4749 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5282_
	);
	LUT2 #(
		.INIT('h1)
	) name4750 (
		_w5281_,
		_w5282_,
		_w5283_
	);
	LUT3 #(
		.INIT('he0)
	) name4751 (
		_w5276_,
		_w5280_,
		_w5283_,
		_w5284_
	);
	LUT3 #(
		.INIT('h45)
	) name4752 (
		\sa23_reg[1]/P0001 ,
		_w5274_,
		_w5284_,
		_w5285_
	);
	LUT3 #(
		.INIT('h80)
	) name4753 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5286_
	);
	LUT4 #(
		.INIT('h2000)
	) name4754 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5287_
	);
	LUT2 #(
		.INIT('h1)
	) name4755 (
		\sa23_reg[2]/P0001 ,
		_w5287_,
		_w5288_
	);
	LUT3 #(
		.INIT('h02)
	) name4756 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w5289_
	);
	LUT4 #(
		.INIT('h2220)
	) name4757 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5290_
	);
	LUT4 #(
		.INIT('h0007)
	) name4758 (
		_w4927_,
		_w4951_,
		_w5289_,
		_w5290_,
		_w5291_
	);
	LUT4 #(
		.INIT('h0001)
	) name4759 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w5292_
	);
	LUT4 #(
		.INIT('h008a)
	) name4760 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		_w4967_,
		_w5292_,
		_w5293_
	);
	LUT4 #(
		.INIT('h0037)
	) name4761 (
		_w4910_,
		_w5288_,
		_w5291_,
		_w5293_,
		_w5294_
	);
	LUT2 #(
		.INIT('h2)
	) name4762 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		_w5295_
	);
	LUT3 #(
		.INIT('h80)
	) name4763 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5296_
	);
	LUT3 #(
		.INIT('h01)
	) name4764 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5297_
	);
	LUT3 #(
		.INIT('h7e)
	) name4765 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5298_
	);
	LUT2 #(
		.INIT('h2)
	) name4766 (
		_w5295_,
		_w5298_,
		_w5299_
	);
	LUT4 #(
		.INIT('h23af)
	) name4767 (
		\sa23_reg[2]/P0001 ,
		_w4910_,
		_w4936_,
		_w4948_,
		_w5300_
	);
	LUT3 #(
		.INIT('h8a)
	) name4768 (
		\sa23_reg[1]/P0001 ,
		_w5299_,
		_w5300_,
		_w5301_
	);
	LUT3 #(
		.INIT('h54)
	) name4769 (
		\sa23_reg[0]/P0001 ,
		_w5294_,
		_w5301_,
		_w5302_
	);
	LUT4 #(
		.INIT('hdfee)
	) name4770 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5303_
	);
	LUT4 #(
		.INIT('h0002)
	) name4771 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5304_
	);
	LUT4 #(
		.INIT('haa02)
	) name4772 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w5303_,
		_w5304_,
		_w5305_
	);
	LUT4 #(
		.INIT('h0001)
	) name4773 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5306_
	);
	LUT4 #(
		.INIT('h0800)
	) name4774 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w5307_
	);
	LUT3 #(
		.INIT('h23)
	) name4775 (
		\sa23_reg[7]/NET0131 ,
		_w5306_,
		_w5307_,
		_w5308_
	);
	LUT3 #(
		.INIT('h8a)
	) name4776 (
		\sa23_reg[2]/P0001 ,
		_w5305_,
		_w5308_,
		_w5309_
	);
	LUT3 #(
		.INIT('h40)
	) name4777 (
		\sa23_reg[2]/P0001 ,
		_w4907_,
		_w4971_,
		_w5310_
	);
	LUT4 #(
		.INIT('h2000)
	) name4778 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[2]/P0001 ,
		_w4907_,
		_w4971_,
		_w5311_
	);
	LUT3 #(
		.INIT('h40)
	) name4779 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		_w4938_,
		_w5312_
	);
	LUT2 #(
		.INIT('h8)
	) name4780 (
		_w4901_,
		_w4919_,
		_w5313_
	);
	LUT3 #(
		.INIT('h01)
	) name4781 (
		_w5312_,
		_w5311_,
		_w5313_,
		_w5314_
	);
	LUT2 #(
		.INIT('h4)
	) name4782 (
		_w5309_,
		_w5314_,
		_w5315_
	);
	LUT4 #(
		.INIT('h0100)
	) name4783 (
		_w5267_,
		_w5302_,
		_w5285_,
		_w5315_,
		_w5316_
	);
	LUT2 #(
		.INIT('h9)
	) name4784 (
		_w5248_,
		_w5316_,
		_w5317_
	);
	LUT4 #(
		.INIT('h5515)
	) name4785 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5318_
	);
	LUT2 #(
		.INIT('h4)
	) name4786 (
		_w4754_,
		_w5318_,
		_w5319_
	);
	LUT3 #(
		.INIT('h10)
	) name4787 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w5320_
	);
	LUT3 #(
		.INIT('h02)
	) name4788 (
		\sa01_reg[2]/P0001 ,
		_w4719_,
		_w5320_,
		_w5321_
	);
	LUT3 #(
		.INIT('h07)
	) name4789 (
		_w4698_,
		_w4749_,
		_w4779_,
		_w5322_
	);
	LUT4 #(
		.INIT('h0155)
	) name4790 (
		\sa01_reg[1]/P0001 ,
		_w5319_,
		_w5321_,
		_w5322_,
		_w5323_
	);
	LUT4 #(
		.INIT('h0123)
	) name4791 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5324_
	);
	LUT3 #(
		.INIT('ha8)
	) name4792 (
		\sa01_reg[1]/P0001 ,
		_w4787_,
		_w5324_,
		_w5325_
	);
	LUT3 #(
		.INIT('h04)
	) name4793 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5326_
	);
	LUT3 #(
		.INIT('h01)
	) name4794 (
		_w4760_,
		_w4779_,
		_w5326_,
		_w5327_
	);
	LUT3 #(
		.INIT('h45)
	) name4795 (
		\sa01_reg[2]/P0001 ,
		_w5325_,
		_w5327_,
		_w5328_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name4796 (
		\sa01_reg[6]/NET0131 ,
		_w4698_,
		_w4709_,
		_w4796_,
		_w5329_
	);
	LUT4 #(
		.INIT('h0200)
	) name4797 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5330_
	);
	LUT3 #(
		.INIT('h07)
	) name4798 (
		_w4698_,
		_w4693_,
		_w5330_,
		_w5331_
	);
	LUT3 #(
		.INIT('h2a)
	) name4799 (
		\sa01_reg[1]/P0001 ,
		_w5329_,
		_w5331_,
		_w5332_
	);
	LUT4 #(
		.INIT('h0777)
	) name4800 (
		_w4698_,
		_w4749_,
		_w4718_,
		_w4801_,
		_w5333_
	);
	LUT4 #(
		.INIT('h153f)
	) name4801 (
		_w4701_,
		_w4723_,
		_w4725_,
		_w4787_,
		_w5334_
	);
	LUT3 #(
		.INIT('hd0)
	) name4802 (
		\sa01_reg[2]/P0001 ,
		_w5333_,
		_w5334_,
		_w5335_
	);
	LUT4 #(
		.INIT('h0100)
	) name4803 (
		_w5328_,
		_w5332_,
		_w5323_,
		_w5335_,
		_w5336_
	);
	LUT3 #(
		.INIT('h04)
	) name4804 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w5337_
	);
	LUT4 #(
		.INIT('h0040)
	) name4805 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w5338_
	);
	LUT3 #(
		.INIT('h20)
	) name4806 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5339_
	);
	LUT4 #(
		.INIT('hf5ef)
	) name4807 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5340_
	);
	LUT3 #(
		.INIT('h45)
	) name4808 (
		\sa01_reg[2]/P0001 ,
		_w5338_,
		_w5340_,
		_w5341_
	);
	LUT3 #(
		.INIT('h80)
	) name4809 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5342_
	);
	LUT4 #(
		.INIT('h0080)
	) name4810 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5343_
	);
	LUT3 #(
		.INIT('ha8)
	) name4811 (
		\sa01_reg[2]/P0001 ,
		_w5342_,
		_w5343_,
		_w5344_
	);
	LUT4 #(
		.INIT('h0400)
	) name4812 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5345_
	);
	LUT4 #(
		.INIT('h0002)
	) name4813 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5346_
	);
	LUT4 #(
		.INIT('heffd)
	) name4814 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5347_
	);
	LUT2 #(
		.INIT('h4)
	) name4815 (
		_w5345_,
		_w5347_,
		_w5348_
	);
	LUT4 #(
		.INIT('h8000)
	) name4816 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5349_
	);
	LUT3 #(
		.INIT('h07)
	) name4817 (
		_w4717_,
		_w4702_,
		_w5349_,
		_w5350_
	);
	LUT4 #(
		.INIT('h1000)
	) name4818 (
		_w5344_,
		_w5341_,
		_w5348_,
		_w5350_,
		_w5351_
	);
	LUT4 #(
		.INIT('h0400)
	) name4819 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5352_
	);
	LUT2 #(
		.INIT('h2)
	) name4820 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		_w5353_
	);
	LUT4 #(
		.INIT('h0002)
	) name4821 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5354_
	);
	LUT3 #(
		.INIT('h54)
	) name4822 (
		\sa01_reg[5]/P0001 ,
		_w5352_,
		_w5354_,
		_w5355_
	);
	LUT3 #(
		.INIT('h01)
	) name4823 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w5356_
	);
	LUT4 #(
		.INIT('h0777)
	) name4824 (
		\sa01_reg[6]/NET0131 ,
		_w4765_,
		_w4775_,
		_w5356_,
		_w5357_
	);
	LUT2 #(
		.INIT('h4)
	) name4825 (
		_w5355_,
		_w5357_,
		_w5358_
	);
	LUT2 #(
		.INIT('h4)
	) name4826 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w5359_
	);
	LUT2 #(
		.INIT('h8)
	) name4827 (
		_w4693_,
		_w5359_,
		_w5360_
	);
	LUT3 #(
		.INIT('h04)
	) name4828 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5361_
	);
	LUT4 #(
		.INIT('h0002)
	) name4829 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5362_
	);
	LUT4 #(
		.INIT('h0001)
	) name4830 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5363_
	);
	LUT4 #(
		.INIT('h0007)
	) name4831 (
		_w4699_,
		_w5361_,
		_w5362_,
		_w5363_,
		_w5364_
	);
	LUT4 #(
		.INIT('h0008)
	) name4832 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5365_
	);
	LUT4 #(
		.INIT('h1000)
	) name4833 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5366_
	);
	LUT3 #(
		.INIT('h54)
	) name4834 (
		\sa01_reg[2]/P0001 ,
		_w5365_,
		_w5366_,
		_w5367_
	);
	LUT3 #(
		.INIT('h80)
	) name4835 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5368_
	);
	LUT3 #(
		.INIT('h01)
	) name4836 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5369_
	);
	LUT3 #(
		.INIT('h7e)
	) name4837 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5370_
	);
	LUT2 #(
		.INIT('h2)
	) name4838 (
		_w4775_,
		_w5370_,
		_w5371_
	);
	LUT4 #(
		.INIT('h0100)
	) name4839 (
		_w5360_,
		_w5367_,
		_w5371_,
		_w5364_,
		_w5372_
	);
	LUT4 #(
		.INIT('hd800)
	) name4840 (
		\sa01_reg[1]/P0001 ,
		_w5351_,
		_w5358_,
		_w5372_,
		_w5373_
	);
	LUT4 #(
		.INIT('h2000)
	) name4841 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5374_
	);
	LUT4 #(
		.INIT('h0013)
	) name4842 (
		\sa01_reg[6]/NET0131 ,
		_w4765_,
		_w4796_,
		_w5374_,
		_w5375_
	);
	LUT3 #(
		.INIT('h6b)
	) name4843 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5376_
	);
	LUT2 #(
		.INIT('h2)
	) name4844 (
		_w4699_,
		_w5376_,
		_w5377_
	);
	LUT3 #(
		.INIT('h08)
	) name4845 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w5378_
	);
	LUT3 #(
		.INIT('h13)
	) name4846 (
		_w4772_,
		_w4794_,
		_w5378_,
		_w5379_
	);
	LUT4 #(
		.INIT('h3200)
	) name4847 (
		\sa01_reg[2]/P0001 ,
		_w5377_,
		_w5375_,
		_w5379_,
		_w5380_
	);
	LUT2 #(
		.INIT('h8)
	) name4848 (
		_w4750_,
		_w5369_,
		_w5381_
	);
	LUT4 #(
		.INIT('h135f)
	) name4849 (
		_w4702_,
		_w4693_,
		_w4699_,
		_w5359_,
		_w5382_
	);
	LUT2 #(
		.INIT('h4)
	) name4850 (
		_w5381_,
		_w5382_,
		_w5383_
	);
	LUT4 #(
		.INIT('h0008)
	) name4851 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5384_
	);
	LUT2 #(
		.INIT('h8)
	) name4852 (
		_w4775_,
		_w5384_,
		_w5385_
	);
	LUT4 #(
		.INIT('h5540)
	) name4853 (
		\sa01_reg[2]/P0001 ,
		_w4692_,
		_w4732_,
		_w4790_,
		_w5386_
	);
	LUT2 #(
		.INIT('h1)
	) name4854 (
		_w5385_,
		_w5386_,
		_w5387_
	);
	LUT4 #(
		.INIT('he400)
	) name4855 (
		\sa01_reg[1]/P0001 ,
		_w5380_,
		_w5383_,
		_w5387_,
		_w5388_
	);
	LUT4 #(
		.INIT('he400)
	) name4856 (
		\sa01_reg[0]/P0001 ,
		_w5373_,
		_w5336_,
		_w5388_,
		_w5389_
	);
	LUT3 #(
		.INIT('h4b)
	) name4857 (
		_w4841_,
		_w4886_,
		_w5389_,
		_w5390_
	);
	LUT4 #(
		.INIT('h1441)
	) name4858 (
		\ld_r_reg/P0001 ,
		_w5195_,
		_w5317_,
		_w5390_,
		_w5391_
	);
	LUT3 #(
		.INIT('h82)
	) name4859 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[94]/P0001 ,
		\u0_w_reg[1][30]/P0001 ,
		_w5392_
	);
	LUT2 #(
		.INIT('h1)
	) name4860 (
		_w5391_,
		_w5392_,
		_w5393_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name4861 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5394_
	);
	LUT4 #(
		.INIT('h80aa)
	) name4862 (
		\sa01_reg[1]/P0001 ,
		_w4697_,
		_w4718_,
		_w5394_,
		_w5395_
	);
	LUT4 #(
		.INIT('h0007)
	) name4863 (
		_w4698_,
		_w4749_,
		_w4705_,
		_w5363_,
		_w5396_
	);
	LUT3 #(
		.INIT('h8a)
	) name4864 (
		\sa01_reg[2]/P0001 ,
		_w5395_,
		_w5396_,
		_w5397_
	);
	LUT3 #(
		.INIT('h8a)
	) name4865 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w5398_
	);
	LUT4 #(
		.INIT('h0040)
	) name4866 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5399_
	);
	LUT4 #(
		.INIT('h0103)
	) name4867 (
		_w4789_,
		_w5338_,
		_w5399_,
		_w5398_,
		_w5400_
	);
	LUT2 #(
		.INIT('h1)
	) name4868 (
		\sa01_reg[2]/P0001 ,
		_w5400_,
		_w5401_
	);
	LUT3 #(
		.INIT('h13)
	) name4869 (
		_w4741_,
		_w4743_,
		_w5337_,
		_w5402_
	);
	LUT3 #(
		.INIT('h45)
	) name4870 (
		\sa01_reg[1]/P0001 ,
		_w5367_,
		_w5402_,
		_w5403_
	);
	LUT4 #(
		.INIT('h2000)
	) name4871 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5404_
	);
	LUT3 #(
		.INIT('h0b)
	) name4872 (
		\sa01_reg[6]/NET0131 ,
		_w4796_,
		_w5404_,
		_w5405_
	);
	LUT4 #(
		.INIT('haa20)
	) name4873 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w4796_,
		_w5404_,
		_w5406_
	);
	LUT2 #(
		.INIT('h4)
	) name4874 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[2]/P0001 ,
		_w5407_
	);
	LUT3 #(
		.INIT('h80)
	) name4875 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5408_
	);
	LUT3 #(
		.INIT('hc8)
	) name4876 (
		_w5361_,
		_w5407_,
		_w5408_,
		_w5409_
	);
	LUT2 #(
		.INIT('h8)
	) name4877 (
		_w4775_,
		_w4784_,
		_w5410_
	);
	LUT3 #(
		.INIT('h01)
	) name4878 (
		_w5406_,
		_w5409_,
		_w5410_,
		_w5411_
	);
	LUT4 #(
		.INIT('h0100)
	) name4879 (
		_w5403_,
		_w5401_,
		_w5397_,
		_w5411_,
		_w5412_
	);
	LUT4 #(
		.INIT('hb8ff)
	) name4880 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5413_
	);
	LUT2 #(
		.INIT('h2)
	) name4881 (
		\sa01_reg[3]/P0001 ,
		_w5413_,
		_w5414_
	);
	LUT4 #(
		.INIT('h0100)
	) name4882 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5415_
	);
	LUT3 #(
		.INIT('h01)
	) name4883 (
		\sa01_reg[1]/P0001 ,
		_w5399_,
		_w5415_,
		_w5416_
	);
	LUT4 #(
		.INIT('h153f)
	) name4884 (
		\sa01_reg[7]/NET0131 ,
		_w4732_,
		_w4775_,
		_w4791_,
		_w5417_
	);
	LUT3 #(
		.INIT('h40)
	) name4885 (
		_w5414_,
		_w5416_,
		_w5417_,
		_w5418_
	);
	LUT2 #(
		.INIT('h2)
	) name4886 (
		_w5353_,
		_w5370_,
		_w5419_
	);
	LUT2 #(
		.INIT('h4)
	) name4887 (
		\sa01_reg[2]/P0001 ,
		_w5363_,
		_w5420_
	);
	LUT3 #(
		.INIT('h2a)
	) name4888 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w4796_,
		_w5421_
	);
	LUT3 #(
		.INIT('h10)
	) name4889 (
		_w5419_,
		_w5420_,
		_w5421_,
		_w5422_
	);
	LUT4 #(
		.INIT('h0004)
	) name4890 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w5423_
	);
	LUT2 #(
		.INIT('h1)
	) name4891 (
		\sa01_reg[2]/P0001 ,
		_w5423_,
		_w5424_
	);
	LUT3 #(
		.INIT('h2a)
	) name4892 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5425_
	);
	LUT4 #(
		.INIT('h0040)
	) name4893 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5426_
	);
	LUT4 #(
		.INIT('h51f3)
	) name4894 (
		\sa01_reg[6]/NET0131 ,
		_w4768_,
		_w5425_,
		_w5426_,
		_w5427_
	);
	LUT4 #(
		.INIT('h0001)
	) name4895 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w5428_
	);
	LUT4 #(
		.INIT('h002a)
	) name4896 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w4791_,
		_w5428_,
		_w5429_
	);
	LUT3 #(
		.INIT('h07)
	) name4897 (
		_w5424_,
		_w5427_,
		_w5429_,
		_w5430_
	);
	LUT3 #(
		.INIT('h0e)
	) name4898 (
		_w5418_,
		_w5422_,
		_w5430_,
		_w5431_
	);
	LUT4 #(
		.INIT('h0800)
	) name4899 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5432_
	);
	LUT4 #(
		.INIT('h0020)
	) name4900 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5433_
	);
	LUT4 #(
		.INIT('hf7df)
	) name4901 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5434_
	);
	LUT3 #(
		.INIT('h45)
	) name4902 (
		\sa01_reg[2]/P0001 ,
		_w5432_,
		_w5434_,
		_w5435_
	);
	LUT4 #(
		.INIT('h4000)
	) name4903 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5436_
	);
	LUT2 #(
		.INIT('h8)
	) name4904 (
		\sa01_reg[2]/P0001 ,
		_w5436_,
		_w5437_
	);
	LUT4 #(
		.INIT('h0800)
	) name4905 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5438_
	);
	LUT4 #(
		.INIT('h1000)
	) name4906 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w5439_
	);
	LUT4 #(
		.INIT('h0007)
	) name4907 (
		\sa01_reg[3]/P0001 ,
		_w5362_,
		_w5438_,
		_w5439_,
		_w5440_
	);
	LUT4 #(
		.INIT('h5455)
	) name4908 (
		\sa01_reg[1]/P0001 ,
		_w5435_,
		_w5437_,
		_w5440_,
		_w5441_
	);
	LUT2 #(
		.INIT('h8)
	) name4909 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[2]/P0001 ,
		_w5442_
	);
	LUT4 #(
		.INIT('h0002)
	) name4910 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5443_
	);
	LUT4 #(
		.INIT('h0207)
	) name4911 (
		\sa01_reg[4]/P0001 ,
		_w4709_,
		_w4794_,
		_w5432_,
		_w5444_
	);
	LUT2 #(
		.INIT('h2)
	) name4912 (
		_w5442_,
		_w5444_,
		_w5445_
	);
	LUT4 #(
		.INIT('hff7a)
	) name4913 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5446_
	);
	LUT2 #(
		.INIT('h2)
	) name4914 (
		_w4716_,
		_w5446_,
		_w5447_
	);
	LUT2 #(
		.INIT('h2)
	) name4915 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[2]/P0001 ,
		_w5448_
	);
	LUT3 #(
		.INIT('h80)
	) name4916 (
		_w4692_,
		_w4732_,
		_w5448_,
		_w5449_
	);
	LUT2 #(
		.INIT('h4)
	) name4917 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		_w5450_
	);
	LUT4 #(
		.INIT('h135f)
	) name4918 (
		_w4709_,
		_w4743_,
		_w4717_,
		_w5450_,
		_w5451_
	);
	LUT3 #(
		.INIT('h10)
	) name4919 (
		_w5449_,
		_w5447_,
		_w5451_,
		_w5452_
	);
	LUT3 #(
		.INIT('h10)
	) name4920 (
		_w5441_,
		_w5445_,
		_w5452_,
		_w5453_
	);
	LUT4 #(
		.INIT('hd800)
	) name4921 (
		\sa01_reg[0]/P0001 ,
		_w5412_,
		_w5431_,
		_w5453_,
		_w5454_
	);
	LUT4 #(
		.INIT('h5655)
	) name4922 (
		\u0_w_reg[1][22]/P0001 ,
		_w5148_,
		_w5170_,
		_w5193_,
		_w5455_
	);
	LUT2 #(
		.INIT('h6)
	) name4923 (
		_w5316_,
		_w5455_,
		_w5456_
	);
	LUT4 #(
		.INIT('h4114)
	) name4924 (
		\ld_r_reg/P0001 ,
		_w5004_,
		_w5454_,
		_w5456_,
		_w5457_
	);
	LUT3 #(
		.INIT('h82)
	) name4925 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[86]/P0001 ,
		\u0_w_reg[1][22]/P0001 ,
		_w5458_
	);
	LUT2 #(
		.INIT('h1)
	) name4926 (
		_w5457_,
		_w5458_,
		_w5459_
	);
	LUT4 #(
		.INIT('haa2a)
	) name4927 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5460_
	);
	LUT3 #(
		.INIT('h20)
	) name4928 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5461_
	);
	LUT4 #(
		.INIT('h0100)
	) name4929 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5462_
	);
	LUT4 #(
		.INIT('h0405)
	) name4930 (
		\sa23_reg[2]/P0001 ,
		_w4925_,
		_w5462_,
		_w5461_,
		_w5463_
	);
	LUT3 #(
		.INIT('h13)
	) name4931 (
		_w4932_,
		_w4982_,
		_w4990_,
		_w5464_
	);
	LUT4 #(
		.INIT('h02aa)
	) name4932 (
		\sa23_reg[1]/P0001 ,
		_w5460_,
		_w5463_,
		_w5464_,
		_w5465_
	);
	LUT4 #(
		.INIT('h0040)
	) name4933 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5466_
	);
	LUT4 #(
		.INIT('h7f7c)
	) name4934 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5467_
	);
	LUT4 #(
		.INIT('h2031)
	) name4935 (
		\sa23_reg[2]/P0001 ,
		_w5275_,
		_w5467_,
		_w5466_,
		_w5468_
	);
	LUT4 #(
		.INIT('h0004)
	) name4936 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5469_
	);
	LUT4 #(
		.INIT('h3310)
	) name4937 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		_w4967_,
		_w5469_,
		_w5470_
	);
	LUT4 #(
		.INIT('h0100)
	) name4938 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w5471_
	);
	LUT4 #(
		.INIT('haa20)
	) name4939 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[5]/P0001 ,
		_w4946_,
		_w5471_,
		_w5472_
	);
	LUT4 #(
		.INIT('h0302)
	) name4940 (
		\sa23_reg[1]/P0001 ,
		_w5470_,
		_w5472_,
		_w5468_,
		_w5473_
	);
	LUT3 #(
		.INIT('h45)
	) name4941 (
		\sa23_reg[0]/P0001 ,
		_w5465_,
		_w5473_,
		_w5474_
	);
	LUT2 #(
		.INIT('h8)
	) name4942 (
		_w4889_,
		_w4901_,
		_w5475_
	);
	LUT4 #(
		.INIT('h0100)
	) name4943 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5476_
	);
	LUT2 #(
		.INIT('h4)
	) name4944 (
		\sa23_reg[6]/NET0131 ,
		_w5476_,
		_w5477_
	);
	LUT4 #(
		.INIT('h0020)
	) name4945 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w5478_
	);
	LUT2 #(
		.INIT('h1)
	) name4946 (
		_w5258_,
		_w5478_,
		_w5479_
	);
	LUT2 #(
		.INIT('h8)
	) name4947 (
		_w4919_,
		_w5259_,
		_w5480_
	);
	LUT4 #(
		.INIT('h020a)
	) name4948 (
		\sa23_reg[2]/P0001 ,
		_w4919_,
		_w4976_,
		_w5259_,
		_w5481_
	);
	LUT3 #(
		.INIT('h40)
	) name4949 (
		_w5477_,
		_w5479_,
		_w5481_,
		_w5482_
	);
	LUT3 #(
		.INIT('h15)
	) name4950 (
		\sa23_reg[2]/P0001 ,
		_w4910_,
		_w4948_,
		_w5483_
	);
	LUT2 #(
		.INIT('h8)
	) name4951 (
		\sa23_reg[6]/NET0131 ,
		_w5254_,
		_w5484_
	);
	LUT4 #(
		.INIT('h45cf)
	) name4952 (
		\sa23_reg[6]/NET0131 ,
		_w4929_,
		_w4964_,
		_w5254_,
		_w5485_
	);
	LUT2 #(
		.INIT('h8)
	) name4953 (
		_w5483_,
		_w5485_,
		_w5486_
	);
	LUT4 #(
		.INIT('h4445)
	) name4954 (
		\sa23_reg[1]/P0001 ,
		_w5475_,
		_w5482_,
		_w5486_,
		_w5487_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name4955 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5488_
	);
	LUT2 #(
		.INIT('h1)
	) name4956 (
		\sa23_reg[2]/P0001 ,
		_w5488_,
		_w5489_
	);
	LUT4 #(
		.INIT('h0200)
	) name4957 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5490_
	);
	LUT4 #(
		.INIT('h002a)
	) name4958 (
		\sa23_reg[1]/P0001 ,
		_w4907_,
		_w4971_,
		_w5490_,
		_w5491_
	);
	LUT3 #(
		.INIT('h10)
	) name4959 (
		_w4960_,
		_w5489_,
		_w5491_,
		_w5492_
	);
	LUT3 #(
		.INIT('h45)
	) name4960 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[2]/P0001 ,
		_w4946_,
		_w5493_
	);
	LUT2 #(
		.INIT('h8)
	) name4961 (
		\sa23_reg[2]/P0001 ,
		_w4938_,
		_w5494_
	);
	LUT2 #(
		.INIT('h1)
	) name4962 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w5495_
	);
	LUT3 #(
		.INIT('h32)
	) name4963 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w5496_
	);
	LUT4 #(
		.INIT('h2000)
	) name4964 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5497_
	);
	LUT3 #(
		.INIT('h0d)
	) name4965 (
		_w4894_,
		_w5496_,
		_w5497_,
		_w5498_
	);
	LUT3 #(
		.INIT('h20)
	) name4966 (
		_w5493_,
		_w5494_,
		_w5498_,
		_w5499_
	);
	LUT4 #(
		.INIT('h35f5)
	) name4967 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5500_
	);
	LUT2 #(
		.INIT('h1)
	) name4968 (
		\sa23_reg[4]/P0001 ,
		_w5500_,
		_w5501_
	);
	LUT3 #(
		.INIT('h02)
	) name4969 (
		\sa23_reg[2]/P0001 ,
		_w4949_,
		_w4959_,
		_w5502_
	);
	LUT3 #(
		.INIT('h07)
	) name4970 (
		_w4901_,
		_w4919_,
		_w4977_,
		_w5503_
	);
	LUT4 #(
		.INIT('h45cf)
	) name4971 (
		_w5288_,
		_w5501_,
		_w5502_,
		_w5503_,
		_w5504_
	);
	LUT4 #(
		.INIT('haa02)
	) name4972 (
		\sa23_reg[0]/P0001 ,
		_w5492_,
		_w5499_,
		_w5504_,
		_w5505_
	);
	LUT3 #(
		.INIT('h0b)
	) name4973 (
		\sa23_reg[3]/P0001 ,
		_w4921_,
		_w5290_,
		_w5506_
	);
	LUT3 #(
		.INIT('h45)
	) name4974 (
		\sa23_reg[2]/P0001 ,
		_w5313_,
		_w5506_,
		_w5507_
	);
	LUT4 #(
		.INIT('h0020)
	) name4975 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5508_
	);
	LUT4 #(
		.INIT('h153f)
	) name4976 (
		\sa23_reg[4]/P0001 ,
		_w4952_,
		_w4992_,
		_w5508_,
		_w5509_
	);
	LUT3 #(
		.INIT('h10)
	) name4977 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5510_
	);
	LUT4 #(
		.INIT('h135f)
	) name4978 (
		\sa23_reg[7]/NET0131 ,
		_w4945_,
		_w5307_,
		_w5510_,
		_w5511_
	);
	LUT2 #(
		.INIT('h8)
	) name4979 (
		_w5509_,
		_w5511_,
		_w5512_
	);
	LUT2 #(
		.INIT('h8)
	) name4980 (
		_w4897_,
		_w4918_,
		_w5513_
	);
	LUT3 #(
		.INIT('h40)
	) name4981 (
		\sa23_reg[2]/P0001 ,
		_w4887_,
		_w4908_,
		_w5514_
	);
	LUT2 #(
		.INIT('h1)
	) name4982 (
		_w5513_,
		_w5514_,
		_w5515_
	);
	LUT4 #(
		.INIT('h7500)
	) name4983 (
		\sa23_reg[1]/P0001 ,
		_w5507_,
		_w5512_,
		_w5515_,
		_w5516_
	);
	LUT4 #(
		.INIT('h0100)
	) name4984 (
		_w5505_,
		_w5487_,
		_w5474_,
		_w5516_,
		_w5517_
	);
	LUT3 #(
		.INIT('h69)
	) name4985 (
		_w4691_,
		_w5389_,
		_w5517_,
		_w5518_
	);
	LUT4 #(
		.INIT('h9a65)
	) name4986 (
		\u0_w_reg[1][21]/P0001 ,
		_w4942_,
		_w5003_,
		_w5121_,
		_w5519_
	);
	LUT3 #(
		.INIT('h82)
	) name4987 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[85]/P0001 ,
		\u0_w_reg[1][21]/P0001 ,
		_w5520_
	);
	LUT4 #(
		.INIT('h00eb)
	) name4988 (
		\ld_r_reg/P0001 ,
		_w5518_,
		_w5519_,
		_w5520_,
		_w5521_
	);
	LUT4 #(
		.INIT('hb44b)
	) name4989 (
		_w4841_,
		_w4886_,
		_w5389_,
		_w5517_,
		_w5522_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name4990 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5523_
	);
	LUT2 #(
		.INIT('h1)
	) name4991 (
		\sa30_reg[2]/P0001 ,
		_w5523_,
		_w5524_
	);
	LUT2 #(
		.INIT('h2)
	) name4992 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w5525_
	);
	LUT4 #(
		.INIT('h0200)
	) name4993 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5526_
	);
	LUT4 #(
		.INIT('h002a)
	) name4994 (
		\sa30_reg[1]/P0001 ,
		_w5029_,
		_w5030_,
		_w5526_,
		_w5527_
	);
	LUT3 #(
		.INIT('h10)
	) name4995 (
		_w5115_,
		_w5524_,
		_w5527_,
		_w5528_
	);
	LUT4 #(
		.INIT('h2000)
	) name4996 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5529_
	);
	LUT2 #(
		.INIT('h1)
	) name4997 (
		\sa30_reg[1]/P0001 ,
		_w5529_,
		_w5530_
	);
	LUT2 #(
		.INIT('h8)
	) name4998 (
		_w5062_,
		_w5102_,
		_w5531_
	);
	LUT2 #(
		.INIT('h1)
	) name4999 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w5532_
	);
	LUT3 #(
		.INIT('h32)
	) name5000 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w5533_
	);
	LUT4 #(
		.INIT('haf23)
	) name5001 (
		\sa30_reg[2]/P0001 ,
		_w5020_,
		_w5013_,
		_w5533_,
		_w5534_
	);
	LUT3 #(
		.INIT('h40)
	) name5002 (
		_w5531_,
		_w5530_,
		_w5534_,
		_w5535_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name5003 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5536_
	);
	LUT4 #(
		.INIT('h0200)
	) name5004 (
		\sa30_reg[2]/P0001 ,
		_w5008_,
		_w5176_,
		_w5536_,
		_w5537_
	);
	LUT4 #(
		.INIT('h2000)
	) name5005 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5538_
	);
	LUT3 #(
		.INIT('h01)
	) name5006 (
		\sa30_reg[2]/P0001 ,
		_w5037_,
		_w5538_,
		_w5539_
	);
	LUT3 #(
		.INIT('h23)
	) name5007 (
		_w5190_,
		_w5537_,
		_w5539_,
		_w5540_
	);
	LUT4 #(
		.INIT('haa02)
	) name5008 (
		\sa30_reg[0]/P0002 ,
		_w5528_,
		_w5535_,
		_w5540_,
		_w5541_
	);
	LUT4 #(
		.INIT('h0100)
	) name5009 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5542_
	);
	LUT4 #(
		.INIT('h5504)
	) name5010 (
		\sa30_reg[2]/P0001 ,
		_w5062_,
		_w5036_,
		_w5542_,
		_w5543_
	);
	LUT3 #(
		.INIT('h20)
	) name5011 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5544_
	);
	LUT4 #(
		.INIT('h0080)
	) name5012 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5545_
	);
	LUT4 #(
		.INIT('h0105)
	) name5013 (
		_w5144_,
		_w5164_,
		_w5545_,
		_w5544_,
		_w5546_
	);
	LUT3 #(
		.INIT('h8a)
	) name5014 (
		\sa30_reg[1]/P0001 ,
		_w5543_,
		_w5546_,
		_w5547_
	);
	LUT4 #(
		.INIT('h5f4e)
	) name5015 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5548_
	);
	LUT4 #(
		.INIT('h0002)
	) name5016 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5549_
	);
	LUT4 #(
		.INIT('h0301)
	) name5017 (
		_w5005_,
		_w5177_,
		_w5549_,
		_w5548_,
		_w5550_
	);
	LUT2 #(
		.INIT('h1)
	) name5018 (
		\sa30_reg[1]/P0001 ,
		_w5550_,
		_w5551_
	);
	LUT3 #(
		.INIT('h08)
	) name5019 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5552_
	);
	LUT4 #(
		.INIT('h0100)
	) name5020 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5553_
	);
	LUT4 #(
		.INIT('haa80)
	) name5021 (
		\sa30_reg[2]/P0001 ,
		_w5044_,
		_w5552_,
		_w5553_,
		_w5554_
	);
	LUT3 #(
		.INIT('h40)
	) name5022 (
		\sa30_reg[3]/P0001 ,
		_w5040_,
		_w5041_,
		_w5555_
	);
	LUT4 #(
		.INIT('h0010)
	) name5023 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5556_
	);
	LUT2 #(
		.INIT('h4)
	) name5024 (
		\sa30_reg[7]/P0001 ,
		_w5556_,
		_w5557_
	);
	LUT3 #(
		.INIT('h01)
	) name5025 (
		_w5555_,
		_w5554_,
		_w5557_,
		_w5558_
	);
	LUT4 #(
		.INIT('h5455)
	) name5026 (
		\sa30_reg[0]/P0002 ,
		_w5547_,
		_w5551_,
		_w5558_,
		_w5559_
	);
	LUT3 #(
		.INIT('h07)
	) name5027 (
		_w5005_,
		_w5072_,
		_w5152_,
		_w5560_
	);
	LUT3 #(
		.INIT('h45)
	) name5028 (
		\sa30_reg[2]/P0001 ,
		_w5190_,
		_w5560_,
		_w5561_
	);
	LUT3 #(
		.INIT('h2a)
	) name5029 (
		\sa30_reg[1]/P0001 ,
		_w5102_,
		_w5109_,
		_w5562_
	);
	LUT2 #(
		.INIT('h4)
	) name5030 (
		\sa30_reg[6]/NET0131 ,
		_w5158_,
		_w5563_
	);
	LUT4 #(
		.INIT('h8000)
	) name5031 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5564_
	);
	LUT4 #(
		.INIT('h2a7f)
	) name5032 (
		\sa30_reg[5]/P0001 ,
		_w5012_,
		_w5112_,
		_w5564_,
		_w5565_
	);
	LUT3 #(
		.INIT('h40)
	) name5033 (
		_w5563_,
		_w5562_,
		_w5565_,
		_w5566_
	);
	LUT3 #(
		.INIT('h20)
	) name5034 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5567_
	);
	LUT4 #(
		.INIT('hcfdf)
	) name5035 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5568_
	);
	LUT2 #(
		.INIT('h1)
	) name5036 (
		\sa30_reg[3]/P0001 ,
		_w5568_,
		_w5569_
	);
	LUT3 #(
		.INIT('h15)
	) name5037 (
		\sa30_reg[2]/P0001 ,
		_w5039_,
		_w5051_,
		_w5570_
	);
	LUT4 #(
		.INIT('h0020)
	) name5038 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5571_
	);
	LUT3 #(
		.INIT('h02)
	) name5039 (
		\sa30_reg[2]/P0001 ,
		_w5019_,
		_w5571_,
		_w5572_
	);
	LUT2 #(
		.INIT('h9)
	) name5040 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w5573_
	);
	LUT3 #(
		.INIT('h13)
	) name5041 (
		_w5099_,
		_w5128_,
		_w5573_,
		_w5574_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name5042 (
		_w5569_,
		_w5570_,
		_w5572_,
		_w5574_,
		_w5575_
	);
	LUT4 #(
		.INIT('h4445)
	) name5043 (
		\sa30_reg[1]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5095_,
		_w5556_,
		_w5576_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name5044 (
		_w5561_,
		_w5566_,
		_w5575_,
		_w5576_,
		_w5577_
	);
	LUT4 #(
		.INIT('h0020)
	) name5045 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5578_
	);
	LUT4 #(
		.INIT('hb1a0)
	) name5046 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w5095_,
		_w5578_,
		_w5579_
	);
	LUT4 #(
		.INIT('h0001)
	) name5047 (
		_w5559_,
		_w5541_,
		_w5577_,
		_w5579_,
		_w5580_
	);
	LUT3 #(
		.INIT('h69)
	) name5048 (
		\u0_w_reg[1][13]/P0001 ,
		_w5121_,
		_w5580_,
		_w5581_
	);
	LUT3 #(
		.INIT('h28)
	) name5049 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[77]/P0001 ,
		\u0_w_reg[1][13]/P0001 ,
		_w5582_
	);
	LUT4 #(
		.INIT('hff41)
	) name5050 (
		\ld_r_reg/P0001 ,
		_w5522_,
		_w5581_,
		_w5582_,
		_w5583_
	);
	LUT4 #(
		.INIT('hb44b)
	) name5051 (
		_w4942_,
		_w5003_,
		_w5248_,
		_w5454_,
		_w5584_
	);
	LUT4 #(
		.INIT('h5655)
	) name5052 (
		\u0_w_reg[1][14]/P0001 ,
		_w5148_,
		_w5170_,
		_w5193_,
		_w5585_
	);
	LUT2 #(
		.INIT('h6)
	) name5053 (
		_w5121_,
		_w5585_,
		_w5586_
	);
	LUT3 #(
		.INIT('h82)
	) name5054 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[78]/P0001 ,
		\u0_w_reg[1][14]/P0001 ,
		_w5587_
	);
	LUT4 #(
		.INIT('h00eb)
	) name5055 (
		\ld_r_reg/P0001 ,
		_w5584_,
		_w5586_,
		_w5587_,
		_w5588_
	);
	LUT3 #(
		.INIT('h69)
	) name5056 (
		_w5248_,
		_w5389_,
		_w5454_,
		_w5589_
	);
	LUT3 #(
		.INIT('h69)
	) name5057 (
		\u0_w_reg[1][6]/P0001 ,
		_w5121_,
		_w5316_,
		_w5590_
	);
	LUT3 #(
		.INIT('h28)
	) name5058 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[70]/P0001 ,
		\u0_w_reg[1][6]/P0001 ,
		_w5591_
	);
	LUT4 #(
		.INIT('hff41)
	) name5059 (
		\ld_r_reg/P0001 ,
		_w5589_,
		_w5590_,
		_w5591_,
		_w5592_
	);
	LUT4 #(
		.INIT('hbfef)
	) name5060 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5593_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name5061 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5594_
	);
	LUT2 #(
		.INIT('h2)
	) name5062 (
		_w5450_,
		_w5594_,
		_w5595_
	);
	LUT3 #(
		.INIT('had)
	) name5063 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w5596_
	);
	LUT4 #(
		.INIT('hadfb)
	) name5064 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5597_
	);
	LUT4 #(
		.INIT('h0302)
	) name5065 (
		\sa01_reg[3]/P0001 ,
		_w4779_,
		_w5366_,
		_w5597_,
		_w5598_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5066 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[2]/P0001 ,
		_w5595_,
		_w5598_,
		_w5599_
	);
	LUT4 #(
		.INIT('h7d5d)
	) name5067 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5600_
	);
	LUT2 #(
		.INIT('h1)
	) name5068 (
		\sa01_reg[2]/P0001 ,
		_w5600_,
		_w5601_
	);
	LUT4 #(
		.INIT('h0100)
	) name5069 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5602_
	);
	LUT3 #(
		.INIT('h31)
	) name5070 (
		\sa01_reg[2]/P0001 ,
		_w5318_,
		_w5602_,
		_w5603_
	);
	LUT3 #(
		.INIT('h0b)
	) name5071 (
		_w4734_,
		_w4771_,
		_w4780_,
		_w5604_
	);
	LUT4 #(
		.INIT('h5455)
	) name5072 (
		\sa01_reg[1]/P0001 ,
		_w5603_,
		_w5601_,
		_w5604_,
		_w5605_
	);
	LUT4 #(
		.INIT('h1000)
	) name5073 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5606_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5074 (
		\sa01_reg[2]/P0001 ,
		_w5343_,
		_w5338_,
		_w5606_,
		_w5607_
	);
	LUT3 #(
		.INIT('hf6)
	) name5075 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5608_
	);
	LUT3 #(
		.INIT('h2a)
	) name5076 (
		_w5442_,
		_w5596_,
		_w5608_,
		_w5609_
	);
	LUT2 #(
		.INIT('h1)
	) name5077 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		_w5610_
	);
	LUT4 #(
		.INIT('h0777)
	) name5078 (
		_w4757_,
		_w4776_,
		_w4784_,
		_w5610_,
		_w5611_
	);
	LUT2 #(
		.INIT('h8)
	) name5079 (
		_w4771_,
		_w5359_,
		_w5612_
	);
	LUT3 #(
		.INIT('h08)
	) name5080 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w5613_
	);
	LUT3 #(
		.INIT('h13)
	) name5081 (
		_w4723_,
		_w5426_,
		_w5613_,
		_w5614_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5082 (
		\sa01_reg[1]/P0001 ,
		_w5611_,
		_w5612_,
		_w5614_,
		_w5615_
	);
	LUT4 #(
		.INIT('h0100)
	) name5083 (
		_w5609_,
		_w5607_,
		_w5605_,
		_w5615_,
		_w5616_
	);
	LUT4 #(
		.INIT('h0020)
	) name5084 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5617_
	);
	LUT3 #(
		.INIT('h54)
	) name5085 (
		\sa01_reg[2]/P0001 ,
		_w4740_,
		_w5617_,
		_w5618_
	);
	LUT4 #(
		.INIT('h008a)
	) name5086 (
		\sa01_reg[1]/P0001 ,
		_w4741_,
		_w4791_,
		_w5432_,
		_w5619_
	);
	LUT4 #(
		.INIT('h77f0)
	) name5087 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5620_
	);
	LUT2 #(
		.INIT('h2)
	) name5088 (
		_w4716_,
		_w5620_,
		_w5621_
	);
	LUT3 #(
		.INIT('h10)
	) name5089 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5622_
	);
	LUT3 #(
		.INIT('h01)
	) name5090 (
		\sa01_reg[1]/P0001 ,
		_w5404_,
		_w5622_,
		_w5623_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name5091 (
		_w5618_,
		_w5619_,
		_w5621_,
		_w5623_,
		_w5624_
	);
	LUT4 #(
		.INIT('h5540)
	) name5092 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w4796_,
		_w5443_,
		_w5625_
	);
	LUT4 #(
		.INIT('h8000)
	) name5093 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5626_
	);
	LUT4 #(
		.INIT('h7ff7)
	) name5094 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5627_
	);
	LUT2 #(
		.INIT('h2)
	) name5095 (
		_w4775_,
		_w5627_,
		_w5628_
	);
	LUT4 #(
		.INIT('h3fbb)
	) name5096 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5629_
	);
	LUT2 #(
		.INIT('h2)
	) name5097 (
		_w5610_,
		_w5629_,
		_w5630_
	);
	LUT4 #(
		.INIT('h7f6e)
	) name5098 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		_w5363_,
		_w5629_,
		_w5631_
	);
	LUT3 #(
		.INIT('h10)
	) name5099 (
		_w5628_,
		_w5625_,
		_w5631_,
		_w5632_
	);
	LUT2 #(
		.INIT('h4)
	) name5100 (
		_w5624_,
		_w5632_,
		_w5633_
	);
	LUT4 #(
		.INIT('h2a7f)
	) name5101 (
		\sa01_reg[5]/P0001 ,
		_w4717_,
		_w4701_,
		_w4719_,
		_w5634_
	);
	LUT2 #(
		.INIT('h1)
	) name5102 (
		\sa01_reg[2]/P0001 ,
		_w5634_,
		_w5635_
	);
	LUT4 #(
		.INIT('h4000)
	) name5103 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w5636_
	);
	LUT4 #(
		.INIT('h0007)
	) name5104 (
		_w4757_,
		_w4776_,
		_w5346_,
		_w5636_,
		_w5637_
	);
	LUT4 #(
		.INIT('h4000)
	) name5105 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5638_
	);
	LUT3 #(
		.INIT('h07)
	) name5106 (
		_w4694_,
		_w5450_,
		_w5638_,
		_w5639_
	);
	LUT4 #(
		.INIT('h3100)
	) name5107 (
		\sa01_reg[2]/P0001 ,
		_w5630_,
		_w5637_,
		_w5639_,
		_w5640_
	);
	LUT3 #(
		.INIT('h32)
	) name5108 (
		\sa01_reg[1]/P0001 ,
		_w5635_,
		_w5640_,
		_w5641_
	);
	LUT4 #(
		.INIT('hd800)
	) name5109 (
		\sa01_reg[0]/P0001 ,
		_w5616_,
		_w5633_,
		_w5641_,
		_w5642_
	);
	LUT3 #(
		.INIT('had)
	) name5110 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w5643_
	);
	LUT3 #(
		.INIT('h01)
	) name5111 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5644_
	);
	LUT3 #(
		.INIT('hf6)
	) name5112 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5645_
	);
	LUT3 #(
		.INIT('h2a)
	) name5113 (
		\sa12_reg[2]/P0001 ,
		_w5643_,
		_w5645_,
		_w5646_
	);
	LUT4 #(
		.INIT('h0100)
	) name5114 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w5647_
	);
	LUT4 #(
		.INIT('h8cbf)
	) name5115 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4664_,
		_w5647_,
		_w5648_
	);
	LUT3 #(
		.INIT('h8a)
	) name5116 (
		\sa12_reg[1]/P0001 ,
		_w5646_,
		_w5648_,
		_w5649_
	);
	LUT4 #(
		.INIT('h7d5d)
	) name5117 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5650_
	);
	LUT2 #(
		.INIT('h1)
	) name5118 (
		\sa12_reg[2]/P0001 ,
		_w5650_,
		_w5651_
	);
	LUT3 #(
		.INIT('h8a)
	) name5119 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w5652_
	);
	LUT4 #(
		.INIT('h00d0)
	) name5120 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5653_
	);
	LUT2 #(
		.INIT('h4)
	) name5121 (
		_w5652_,
		_w5653_,
		_w5654_
	);
	LUT4 #(
		.INIT('h0100)
	) name5122 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w5655_
	);
	LUT3 #(
		.INIT('h13)
	) name5123 (
		\sa12_reg[2]/P0001 ,
		_w4660_,
		_w5655_,
		_w5656_
	);
	LUT4 #(
		.INIT('h5455)
	) name5124 (
		\sa12_reg[1]/P0001 ,
		_w5651_,
		_w5654_,
		_w5656_,
		_w5657_
	);
	LUT3 #(
		.INIT('h8d)
	) name5125 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w5658_
	);
	LUT4 #(
		.INIT('h0301)
	) name5126 (
		_w4687_,
		_w4807_,
		_w4811_,
		_w5658_,
		_w5659_
	);
	LUT3 #(
		.INIT('h13)
	) name5127 (
		_w4685_,
		_w4875_,
		_w5202_,
		_w5660_
	);
	LUT3 #(
		.INIT('hd0)
	) name5128 (
		\sa12_reg[2]/P0001 ,
		_w5659_,
		_w5660_,
		_w5661_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5129 (
		\sa12_reg[0]/P0001 ,
		_w5657_,
		_w5649_,
		_w5661_,
		_w5662_
	);
	LUT4 #(
		.INIT('hbfef)
	) name5130 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5663_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name5131 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5664_
	);
	LUT2 #(
		.INIT('h2)
	) name5132 (
		_w4605_,
		_w5664_,
		_w5665_
	);
	LUT4 #(
		.INIT('h0004)
	) name5133 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5666_
	);
	LUT4 #(
		.INIT('hadfb)
	) name5134 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5667_
	);
	LUT4 #(
		.INIT('h0302)
	) name5135 (
		\sa12_reg[3]/P0001 ,
		_w4661_,
		_w4835_,
		_w5667_,
		_w5668_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5136 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[2]/P0001 ,
		_w5665_,
		_w5668_,
		_w5669_
	);
	LUT4 #(
		.INIT('h4440)
	) name5137 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4661_,
		_w4596_,
		_w5670_
	);
	LUT4 #(
		.INIT('h7ff7)
	) name5138 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5671_
	);
	LUT2 #(
		.INIT('h2)
	) name5139 (
		_w4684_,
		_w5671_,
		_w5672_
	);
	LUT4 #(
		.INIT('h3fbb)
	) name5140 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5673_
	);
	LUT2 #(
		.INIT('h2)
	) name5141 (
		_w5202_,
		_w5673_,
		_w5674_
	);
	LUT4 #(
		.INIT('h0002)
	) name5142 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5675_
	);
	LUT4 #(
		.INIT('h51f3)
	) name5143 (
		_w4617_,
		_w5202_,
		_w5673_,
		_w5675_,
		_w5676_
	);
	LUT3 #(
		.INIT('h10)
	) name5144 (
		_w5672_,
		_w5670_,
		_w5676_,
		_w5677_
	);
	LUT3 #(
		.INIT('h54)
	) name5145 (
		\sa12_reg[2]/P0001 ,
		_w4849_,
		_w5242_,
		_w5678_
	);
	LUT2 #(
		.INIT('h1)
	) name5146 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w5679_
	);
	LUT3 #(
		.INIT('h31)
	) name5147 (
		_w4648_,
		_w5238_,
		_w5679_,
		_w5680_
	);
	LUT3 #(
		.INIT('h8a)
	) name5148 (
		\sa12_reg[1]/P0001 ,
		_w5678_,
		_w5680_,
		_w5681_
	);
	LUT2 #(
		.INIT('h8)
	) name5149 (
		_w4620_,
		_w4871_,
		_w5682_
	);
	LUT3 #(
		.INIT('h10)
	) name5150 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w5683_
	);
	LUT3 #(
		.INIT('h01)
	) name5151 (
		_w4641_,
		_w5205_,
		_w5683_,
		_w5684_
	);
	LUT3 #(
		.INIT('h45)
	) name5152 (
		\sa12_reg[1]/P0001 ,
		_w5682_,
		_w5684_,
		_w5685_
	);
	LUT4 #(
		.INIT('h5455)
	) name5153 (
		\sa12_reg[0]/P0001 ,
		_w5681_,
		_w5685_,
		_w5677_,
		_w5686_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5154 (
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w4650_,
		_w4813_,
		_w5687_
	);
	LUT2 #(
		.INIT('h1)
	) name5155 (
		\sa12_reg[2]/P0001 ,
		_w5687_,
		_w5688_
	);
	LUT4 #(
		.INIT('h4000)
	) name5156 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w5689_
	);
	LUT4 #(
		.INIT('h0007)
	) name5157 (
		_w4664_,
		_w4647_,
		_w4816_,
		_w5689_,
		_w5690_
	);
	LUT4 #(
		.INIT('h4000)
	) name5158 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w5691_
	);
	LUT3 #(
		.INIT('h07)
	) name5159 (
		_w4617_,
		_w5683_,
		_w5691_,
		_w5692_
	);
	LUT4 #(
		.INIT('h3100)
	) name5160 (
		\sa12_reg[2]/P0001 ,
		_w5674_,
		_w5690_,
		_w5692_,
		_w5693_
	);
	LUT3 #(
		.INIT('h32)
	) name5161 (
		\sa12_reg[1]/P0001 ,
		_w5688_,
		_w5693_,
		_w5694_
	);
	LUT4 #(
		.INIT('h0100)
	) name5162 (
		_w5669_,
		_w5662_,
		_w5686_,
		_w5694_,
		_w5695_
	);
	LUT3 #(
		.INIT('hb4)
	) name5163 (
		_w5599_,
		_w5642_,
		_w5695_,
		_w5696_
	);
	LUT4 #(
		.INIT('h659a)
	) name5164 (
		_w5454_,
		_w5599_,
		_w5642_,
		_w5695_,
		_w5697_
	);
	LUT4 #(
		.INIT('h7d1d)
	) name5165 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5698_
	);
	LUT2 #(
		.INIT('h1)
	) name5166 (
		\sa23_reg[2]/P0001 ,
		_w5698_,
		_w5699_
	);
	LUT2 #(
		.INIT('h2)
	) name5167 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w5700_
	);
	LUT4 #(
		.INIT('h00d0)
	) name5168 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5701_
	);
	LUT4 #(
		.INIT('h0200)
	) name5169 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5702_
	);
	LUT4 #(
		.INIT('h2223)
	) name5170 (
		\sa23_reg[3]/P0001 ,
		_w5478_,
		_w5701_,
		_w5702_,
		_w5703_
	);
	LUT3 #(
		.INIT('h45)
	) name5171 (
		\sa23_reg[1]/P0001 ,
		_w5699_,
		_w5703_,
		_w5704_
	);
	LUT4 #(
		.INIT('hcfca)
	) name5172 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5705_
	);
	LUT3 #(
		.INIT('h08)
	) name5173 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5706_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5174 (
		\sa23_reg[1]/P0001 ,
		_w5289_,
		_w5706_,
		_w5705_,
		_w5707_
	);
	LUT4 #(
		.INIT('h1000)
	) name5175 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5708_
	);
	LUT3 #(
		.INIT('h01)
	) name5176 (
		_w4891_,
		_w4898_,
		_w5708_,
		_w5709_
	);
	LUT3 #(
		.INIT('h8a)
	) name5177 (
		\sa23_reg[2]/P0001 ,
		_w5707_,
		_w5709_,
		_w5710_
	);
	LUT4 #(
		.INIT('h0100)
	) name5178 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5711_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name5179 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5307_,
		_w5711_,
		_w5712_
	);
	LUT4 #(
		.INIT('h0040)
	) name5180 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5713_
	);
	LUT3 #(
		.INIT('h08)
	) name5181 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w5714_
	);
	LUT4 #(
		.INIT('h153f)
	) name5182 (
		_w4905_,
		_w5249_,
		_w5252_,
		_w5714_,
		_w5715_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5183 (
		\sa23_reg[1]/P0001 ,
		_w5712_,
		_w5713_,
		_w5715_,
		_w5716_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5184 (
		\sa23_reg[0]/P0001 ,
		_w5710_,
		_w5704_,
		_w5716_,
		_w5717_
	);
	LUT3 #(
		.INIT('h20)
	) name5185 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5718_
	);
	LUT2 #(
		.INIT('h8)
	) name5186 (
		_w4918_,
		_w5718_,
		_w5719_
	);
	LUT4 #(
		.INIT('h0002)
	) name5187 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5720_
	);
	LUT3 #(
		.INIT('h10)
	) name5188 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5721_
	);
	LUT4 #(
		.INIT('h0001)
	) name5189 (
		\sa23_reg[1]/P0001 ,
		_w5254_,
		_w5720_,
		_w5721_,
		_w5722_
	);
	LUT4 #(
		.INIT('h0020)
	) name5190 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5723_
	);
	LUT3 #(
		.INIT('h08)
	) name5191 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w5724_
	);
	LUT3 #(
		.INIT('h54)
	) name5192 (
		\sa23_reg[2]/P0001 ,
		_w5723_,
		_w5724_,
		_w5725_
	);
	LUT2 #(
		.INIT('h8)
	) name5193 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w5726_
	);
	LUT3 #(
		.INIT('h37)
	) name5194 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5727_
	);
	LUT4 #(
		.INIT('h0a02)
	) name5195 (
		\sa23_reg[1]/P0001 ,
		_w4964_,
		_w5279_,
		_w5727_,
		_w5728_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name5196 (
		_w5719_,
		_w5722_,
		_w5725_,
		_w5728_,
		_w5729_
	);
	LUT2 #(
		.INIT('h8)
	) name5197 (
		_w4925_,
		_w5720_,
		_w5730_
	);
	LUT4 #(
		.INIT('h8000)
	) name5198 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5731_
	);
	LUT4 #(
		.INIT('h7ff7)
	) name5199 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5732_
	);
	LUT3 #(
		.INIT('ha2)
	) name5200 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		_w5732_,
		_w5733_
	);
	LUT4 #(
		.INIT('h4000)
	) name5201 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5734_
	);
	LUT4 #(
		.INIT('h0010)
	) name5202 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5735_
	);
	LUT3 #(
		.INIT('h01)
	) name5203 (
		_w5304_,
		_w5734_,
		_w5735_,
		_w5736_
	);
	LUT4 #(
		.INIT('h3230)
	) name5204 (
		_w5483_,
		_w5730_,
		_w5733_,
		_w5736_,
		_w5737_
	);
	LUT3 #(
		.INIT('h45)
	) name5205 (
		\sa23_reg[0]/P0001 ,
		_w5729_,
		_w5737_,
		_w5738_
	);
	LUT4 #(
		.INIT('hadfb)
	) name5206 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5739_
	);
	LUT2 #(
		.INIT('h1)
	) name5207 (
		\sa23_reg[3]/P0001 ,
		_w5739_,
		_w5740_
	);
	LUT3 #(
		.INIT('h02)
	) name5208 (
		\sa23_reg[2]/P0001 ,
		_w4933_,
		_w4976_,
		_w5741_
	);
	LUT4 #(
		.INIT('h0010)
	) name5209 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5742_
	);
	LUT4 #(
		.INIT('hbfef)
	) name5210 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5743_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name5211 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w5744_
	);
	LUT4 #(
		.INIT('h88a8)
	) name5212 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		_w5744_,
		_w5745_
	);
	LUT3 #(
		.INIT('hb0)
	) name5213 (
		_w5740_,
		_w5741_,
		_w5745_,
		_w5746_
	);
	LUT2 #(
		.INIT('h4)
	) name5214 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[2]/P0001 ,
		_w5747_
	);
	LUT4 #(
		.INIT('h4000)
	) name5215 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w5748_
	);
	LUT4 #(
		.INIT('h0013)
	) name5216 (
		\sa23_reg[7]/NET0131 ,
		_w4909_,
		_w5307_,
		_w5748_,
		_w5749_
	);
	LUT2 #(
		.INIT('h2)
	) name5217 (
		_w5747_,
		_w5749_,
		_w5750_
	);
	LUT4 #(
		.INIT('h2a7f)
	) name5218 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4901_,
		_w4946_,
		_w5751_
	);
	LUT2 #(
		.INIT('h2)
	) name5219 (
		\sa23_reg[2]/P0001 ,
		_w4953_,
		_w5752_
	);
	LUT3 #(
		.INIT('h51)
	) name5220 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[2]/P0001 ,
		_w4953_,
		_w5753_
	);
	LUT4 #(
		.INIT('hbdff)
	) name5221 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5754_
	);
	LUT3 #(
		.INIT('h10)
	) name5222 (
		_w5734_,
		_w5735_,
		_w5754_,
		_w5755_
	);
	LUT4 #(
		.INIT('hee0e)
	) name5223 (
		\sa23_reg[2]/P0001 ,
		_w5751_,
		_w5753_,
		_w5755_,
		_w5756_
	);
	LUT3 #(
		.INIT('h10)
	) name5224 (
		_w5750_,
		_w5746_,
		_w5756_,
		_w5757_
	);
	LUT3 #(
		.INIT('h10)
	) name5225 (
		_w5717_,
		_w5738_,
		_w5757_,
		_w5758_
	);
	LUT4 #(
		.INIT('h5655)
	) name5226 (
		\u0_w_reg[1][7]/P0001 ,
		_w5717_,
		_w5738_,
		_w5757_,
		_w5759_
	);
	LUT2 #(
		.INIT('h6)
	) name5227 (
		_w5194_,
		_w5759_,
		_w5760_
	);
	LUT3 #(
		.INIT('h82)
	) name5228 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[71]/P0001 ,
		\u0_w_reg[1][7]/P0001 ,
		_w5761_
	);
	LUT4 #(
		.INIT('h00be)
	) name5229 (
		\ld_r_reg/P0001 ,
		_w5697_,
		_w5760_,
		_w5761_,
		_w5762_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name5230 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5763_
	);
	LUT2 #(
		.INIT('h2)
	) name5231 (
		\sa12_reg[2]/P0001 ,
		_w5763_,
		_w5764_
	);
	LUT4 #(
		.INIT('h5540)
	) name5232 (
		\sa12_reg[2]/P0001 ,
		_w4665_,
		_w4651_,
		_w5230_,
		_w5765_
	);
	LUT2 #(
		.INIT('h8)
	) name5233 (
		\sa12_reg[4]/P0001 ,
		_w5242_,
		_w5766_
	);
	LUT4 #(
		.INIT('h153f)
	) name5234 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4668_,
		_w5242_,
		_w5767_
	);
	LUT4 #(
		.INIT('h5455)
	) name5235 (
		\sa12_reg[1]/P0001 ,
		_w5765_,
		_w5764_,
		_w5767_,
		_w5768_
	);
	LUT3 #(
		.INIT('h4c)
	) name5236 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w5769_
	);
	LUT4 #(
		.INIT('h0803)
	) name5237 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w5770_
	);
	LUT3 #(
		.INIT('h54)
	) name5238 (
		\sa12_reg[2]/P0001 ,
		_w4829_,
		_w5770_,
		_w5771_
	);
	LUT3 #(
		.INIT('ha8)
	) name5239 (
		\sa12_reg[2]/P0001 ,
		_w4675_,
		_w4602_,
		_w5772_
	);
	LUT3 #(
		.INIT('h01)
	) name5240 (
		_w4661_,
		_w4626_,
		_w4816_,
		_w5773_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5241 (
		\sa12_reg[1]/P0001 ,
		_w5771_,
		_w5772_,
		_w5773_,
		_w5774_
	);
	LUT4 #(
		.INIT('h4440)
	) name5242 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4668_,
		_w4807_,
		_w5775_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5243 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5776_
	);
	LUT2 #(
		.INIT('h2)
	) name5244 (
		_w4635_,
		_w5776_,
		_w5777_
	);
	LUT3 #(
		.INIT('h13)
	) name5245 (
		_w4684_,
		_w4872_,
		_w4881_,
		_w5778_
	);
	LUT3 #(
		.INIT('h10)
	) name5246 (
		_w5777_,
		_w5775_,
		_w5778_,
		_w5779_
	);
	LUT4 #(
		.INIT('h5455)
	) name5247 (
		\sa12_reg[0]/P0001 ,
		_w5768_,
		_w5774_,
		_w5779_,
		_w5780_
	);
	LUT3 #(
		.INIT('h07)
	) name5248 (
		_w4608_,
		_w4602_,
		_w4835_,
		_w5781_
	);
	LUT4 #(
		.INIT('h3120)
	) name5249 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5782_
	);
	LUT3 #(
		.INIT('ha8)
	) name5250 (
		\sa12_reg[2]/P0001 ,
		_w4609_,
		_w5782_,
		_w5783_
	);
	LUT3 #(
		.INIT('ha2)
	) name5251 (
		\sa12_reg[1]/P0001 ,
		_w5781_,
		_w5783_,
		_w5784_
	);
	LUT4 #(
		.INIT('h0001)
	) name5252 (
		_w4688_,
		_w4646_,
		_w4881_,
		_w5238_,
		_w5785_
	);
	LUT2 #(
		.INIT('h1)
	) name5253 (
		\sa12_reg[2]/P0001 ,
		_w5785_,
		_w5786_
	);
	LUT2 #(
		.INIT('h8)
	) name5254 (
		\sa12_reg[5]/P0001 ,
		_w5221_,
		_w5787_
	);
	LUT4 #(
		.INIT('h0080)
	) name5255 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w5788_
	);
	LUT4 #(
		.INIT('h0045)
	) name5256 (
		_w4688_,
		_w4597_,
		_w4808_,
		_w5788_,
		_w5789_
	);
	LUT4 #(
		.INIT('h113f)
	) name5257 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4663_,
		_w4670_,
		_w5790_
	);
	LUT4 #(
		.INIT('hba00)
	) name5258 (
		\sa12_reg[1]/P0001 ,
		_w5787_,
		_w5789_,
		_w5790_,
		_w5791_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5259 (
		\sa12_reg[0]/P0001 ,
		_w5784_,
		_w5786_,
		_w5791_,
		_w5792_
	);
	LUT4 #(
		.INIT('h0007)
	) name5260 (
		_w4595_,
		_w4596_,
		_w5205_,
		_w5242_,
		_w5793_
	);
	LUT4 #(
		.INIT('h153f)
	) name5261 (
		_w4591_,
		_w4664_,
		_w4587_,
		_w4849_,
		_w5794_
	);
	LUT4 #(
		.INIT('h0155)
	) name5262 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[2]/P0001 ,
		_w5793_,
		_w5794_,
		_w5795_
	);
	LUT3 #(
		.INIT('h04)
	) name5263 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w5796_
	);
	LUT4 #(
		.INIT('h0a0b)
	) name5264 (
		_w4586_,
		_w4837_,
		_w5208_,
		_w5796_,
		_w5797_
	);
	LUT2 #(
		.INIT('h2)
	) name5265 (
		_w4857_,
		_w5797_,
		_w5798_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name5266 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5799_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5267 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4648_,
		_w5799_,
		_w5800_
	);
	LUT2 #(
		.INIT('h2)
	) name5268 (
		_w5237_,
		_w5800_,
		_w5801_
	);
	LUT4 #(
		.INIT('h7cfa)
	) name5269 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w5802_
	);
	LUT2 #(
		.INIT('h4)
	) name5270 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[2]/P0001 ,
		_w5803_
	);
	LUT3 #(
		.INIT('h04)
	) name5271 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		_w5804_
	);
	LUT2 #(
		.INIT('h4)
	) name5272 (
		_w5802_,
		_w5804_,
		_w5805_
	);
	LUT3 #(
		.INIT('h2e)
	) name5273 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w5806_
	);
	LUT2 #(
		.INIT('h8)
	) name5274 (
		_w4816_,
		_w5806_,
		_w5807_
	);
	LUT3 #(
		.INIT('h80)
	) name5275 (
		\sa12_reg[2]/P0001 ,
		_w4664_,
		_w4587_,
		_w5808_
	);
	LUT3 #(
		.INIT('h01)
	) name5276 (
		_w5807_,
		_w5808_,
		_w5805_,
		_w5809_
	);
	LUT4 #(
		.INIT('h0100)
	) name5277 (
		_w5801_,
		_w5798_,
		_w5795_,
		_w5809_,
		_w5810_
	);
	LUT3 #(
		.INIT('h10)
	) name5278 (
		_w5792_,
		_w5780_,
		_w5810_,
		_w5811_
	);
	LUT3 #(
		.INIT('h20)
	) name5279 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w5812_
	);
	LUT4 #(
		.INIT('h0800)
	) name5280 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w5813_
	);
	LUT3 #(
		.INIT('h10)
	) name5281 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5814_
	);
	LUT4 #(
		.INIT('h5554)
	) name5282 (
		\sa01_reg[2]/P0001 ,
		_w5356_,
		_w5814_,
		_w5813_,
		_w5815_
	);
	LUT4 #(
		.INIT('h0002)
	) name5283 (
		\sa01_reg[1]/P0001 ,
		_w4760_,
		_w4779_,
		_w5346_,
		_w5816_
	);
	LUT2 #(
		.INIT('h4)
	) name5284 (
		_w5815_,
		_w5816_,
		_w5817_
	);
	LUT4 #(
		.INIT('h5540)
	) name5285 (
		\sa01_reg[2]/P0001 ,
		_w4697_,
		_w4718_,
		_w5433_,
		_w5818_
	);
	LUT2 #(
		.INIT('h8)
	) name5286 (
		_w4704_,
		_w5361_,
		_w5819_
	);
	LUT3 #(
		.INIT('h15)
	) name5287 (
		\sa01_reg[1]/P0001 ,
		_w4738_,
		_w4787_,
		_w5820_
	);
	LUT3 #(
		.INIT('h10)
	) name5288 (
		_w5819_,
		_w5818_,
		_w5820_,
		_w5821_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5289 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5822_
	);
	LUT2 #(
		.INIT('h2)
	) name5290 (
		_w5353_,
		_w5822_,
		_w5823_
	);
	LUT3 #(
		.INIT('h13)
	) name5291 (
		_w4775_,
		_w4794_,
		_w5384_,
		_w5824_
	);
	LUT2 #(
		.INIT('h4)
	) name5292 (
		_w5823_,
		_w5824_,
		_w5825_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name5293 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5826_
	);
	LUT2 #(
		.INIT('h2)
	) name5294 (
		_w5407_,
		_w5826_,
		_w5827_
	);
	LUT4 #(
		.INIT('h4000)
	) name5295 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5828_
	);
	LUT3 #(
		.INIT('hc8)
	) name5296 (
		_w5368_,
		_w5442_,
		_w5828_,
		_w5829_
	);
	LUT4 #(
		.INIT('h135f)
	) name5297 (
		_w4698_,
		_w4738_,
		_w4693_,
		_w4787_,
		_w5830_
	);
	LUT4 #(
		.INIT('h0032)
	) name5298 (
		\sa01_reg[2]/P0001 ,
		_w5829_,
		_w5830_,
		_w5827_,
		_w5831_
	);
	LUT4 #(
		.INIT('he000)
	) name5299 (
		_w5817_,
		_w5821_,
		_w5825_,
		_w5831_,
		_w5832_
	);
	LUT3 #(
		.INIT('h07)
	) name5300 (
		_w4704_,
		_w4749_,
		_w5366_,
		_w5833_
	);
	LUT3 #(
		.INIT('h80)
	) name5301 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5834_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5302 (
		\sa01_reg[2]/P0001 ,
		_w4694_,
		_w5834_,
		_w5812_,
		_w5835_
	);
	LUT3 #(
		.INIT('ha2)
	) name5303 (
		\sa01_reg[1]/P0001 ,
		_w5833_,
		_w5835_,
		_w5836_
	);
	LUT2 #(
		.INIT('h4)
	) name5304 (
		\sa01_reg[6]/NET0131 ,
		_w4765_,
		_w5837_
	);
	LUT4 #(
		.INIT('h0203)
	) name5305 (
		_w4734_,
		_w4796_,
		_w4802_,
		_w5339_,
		_w5838_
	);
	LUT3 #(
		.INIT('h45)
	) name5306 (
		\sa01_reg[1]/P0001 ,
		_w5837_,
		_w5838_,
		_w5839_
	);
	LUT2 #(
		.INIT('h4)
	) name5307 (
		_w4745_,
		_w4790_,
		_w5840_
	);
	LUT3 #(
		.INIT('h8a)
	) name5308 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		_w5384_,
		_w5841_
	);
	LUT4 #(
		.INIT('h0001)
	) name5309 (
		_w4712_,
		_w4802_,
		_w5384_,
		_w5432_,
		_w5842_
	);
	LUT3 #(
		.INIT('h54)
	) name5310 (
		_w5840_,
		_w5841_,
		_w5842_,
		_w5843_
	);
	LUT3 #(
		.INIT('h10)
	) name5311 (
		_w5836_,
		_w5839_,
		_w5843_,
		_w5844_
	);
	LUT4 #(
		.INIT('h0100)
	) name5312 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5845_
	);
	LUT4 #(
		.INIT('h0007)
	) name5313 (
		_w4698_,
		_w4749_,
		_w4794_,
		_w5845_,
		_w5846_
	);
	LUT2 #(
		.INIT('h8)
	) name5314 (
		_w4740_,
		_w4697_,
		_w5847_
	);
	LUT4 #(
		.INIT('hedff)
	) name5315 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w4704_,
		_w5848_
	);
	LUT4 #(
		.INIT('h0455)
	) name5316 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[2]/P0001 ,
		_w5846_,
		_w5848_,
		_w5849_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name5317 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5850_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5318 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w4791_,
		_w5850_,
		_w5851_
	);
	LUT2 #(
		.INIT('h2)
	) name5319 (
		_w5442_,
		_w5851_,
		_w5852_
	);
	LUT3 #(
		.INIT('h54)
	) name5320 (
		_w4724_,
		_w5337_,
		_w5363_,
		_w5853_
	);
	LUT2 #(
		.INIT('h1)
	) name5321 (
		_w5346_,
		_w5399_,
		_w5854_
	);
	LUT3 #(
		.INIT('h8a)
	) name5322 (
		_w5448_,
		_w5853_,
		_w5854_,
		_w5855_
	);
	LUT2 #(
		.INIT('h1)
	) name5323 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[2]/P0001 ,
		_w5856_
	);
	LUT4 #(
		.INIT('h0007)
	) name5324 (
		_w4698_,
		_w4709_,
		_w5404_,
		_w5617_,
		_w5857_
	);
	LUT4 #(
		.INIT('h153f)
	) name5325 (
		_w4716_,
		_w4775_,
		_w5363_,
		_w5438_,
		_w5858_
	);
	LUT3 #(
		.INIT('hd0)
	) name5326 (
		_w5856_,
		_w5857_,
		_w5858_,
		_w5859_
	);
	LUT4 #(
		.INIT('h0100)
	) name5327 (
		_w5855_,
		_w5852_,
		_w5849_,
		_w5859_,
		_w5860_
	);
	LUT4 #(
		.INIT('hd800)
	) name5328 (
		\sa01_reg[0]/P0001 ,
		_w5844_,
		_w5832_,
		_w5860_,
		_w5861_
	);
	LUT2 #(
		.INIT('h6)
	) name5329 (
		_w5811_,
		_w5861_,
		_w5862_
	);
	LUT4 #(
		.INIT('h0001)
	) name5330 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5863_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5331 (
		\sa01_reg[2]/P0001 ,
		_w5343_,
		_w5374_,
		_w5863_,
		_w5864_
	);
	LUT3 #(
		.INIT('h8a)
	) name5332 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5865_
	);
	LUT2 #(
		.INIT('h2)
	) name5333 (
		_w4692_,
		_w5865_,
		_w5866_
	);
	LUT4 #(
		.INIT('h0010)
	) name5334 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5867_
	);
	LUT3 #(
		.INIT('h07)
	) name5335 (
		_w5359_,
		_w5845_,
		_w5867_,
		_w5868_
	);
	LUT4 #(
		.INIT('h5455)
	) name5336 (
		\sa01_reg[1]/P0001 ,
		_w5866_,
		_w5864_,
		_w5868_,
		_w5869_
	);
	LUT3 #(
		.INIT('h07)
	) name5337 (
		_w4698_,
		_w4693_,
		_w4695_,
		_w5870_
	);
	LUT3 #(
		.INIT('h2a)
	) name5338 (
		\sa01_reg[2]/P0001 ,
		_w5405_,
		_w5870_,
		_w5871_
	);
	LUT4 #(
		.INIT('h4041)
	) name5339 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5872_
	);
	LUT3 #(
		.INIT('ha8)
	) name5340 (
		\sa01_reg[1]/P0001 ,
		_w5433_,
		_w5872_,
		_w5873_
	);
	LUT3 #(
		.INIT('h54)
	) name5341 (
		\sa01_reg[2]/P0001 ,
		_w5426_,
		_w5626_,
		_w5874_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name5342 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5875_
	);
	LUT2 #(
		.INIT('h2)
	) name5343 (
		_w5450_,
		_w5875_,
		_w5876_
	);
	LUT3 #(
		.INIT('h07)
	) name5344 (
		_w4697_,
		_w4751_,
		_w4712_,
		_w5877_
	);
	LUT4 #(
		.INIT('h0100)
	) name5345 (
		_w5873_,
		_w5876_,
		_w5874_,
		_w5877_,
		_w5878_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5346 (
		\sa01_reg[0]/P0001 ,
		_w5871_,
		_w5869_,
		_w5878_,
		_w5879_
	);
	LUT4 #(
		.INIT('h8000)
	) name5347 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5880_
	);
	LUT4 #(
		.INIT('h0007)
	) name5348 (
		_w4698_,
		_w4693_,
		_w5428_,
		_w5880_,
		_w5881_
	);
	LUT3 #(
		.INIT('hb9)
	) name5349 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5882_
	);
	LUT4 #(
		.INIT('h4c00)
	) name5350 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5883_
	);
	LUT4 #(
		.INIT('h51f3)
	) name5351 (
		_w5407_,
		_w5613_,
		_w5882_,
		_w5883_,
		_w5884_
	);
	LUT3 #(
		.INIT('he0)
	) name5352 (
		\sa01_reg[2]/P0001 ,
		_w5881_,
		_w5884_,
		_w5885_
	);
	LUT4 #(
		.INIT('h3f2a)
	) name5353 (
		\sa01_reg[3]/P0001 ,
		_w4740_,
		_w4741_,
		_w5593_,
		_w5886_
	);
	LUT2 #(
		.INIT('h8)
	) name5354 (
		_w4702_,
		_w4775_,
		_w5887_
	);
	LUT4 #(
		.INIT('h8000)
	) name5355 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5888_
	);
	LUT4 #(
		.INIT('h0100)
	) name5356 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w5889_
	);
	LUT4 #(
		.INIT('h0007)
	) name5357 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5890_
	);
	LUT3 #(
		.INIT('h01)
	) name5358 (
		_w5889_,
		_w5890_,
		_w5888_,
		_w5891_
	);
	LUT4 #(
		.INIT('h4e44)
	) name5359 (
		\sa01_reg[1]/P0001 ,
		_w5886_,
		_w5887_,
		_w5891_,
		_w5892_
	);
	LUT3 #(
		.INIT('h15)
	) name5360 (
		\sa01_reg[0]/P0001 ,
		_w5885_,
		_w5892_,
		_w5893_
	);
	LUT4 #(
		.INIT('h034f)
	) name5361 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		_w4771_,
		_w4794_,
		_w5894_
	);
	LUT2 #(
		.INIT('h1)
	) name5362 (
		\sa01_reg[2]/P0001 ,
		_w5894_,
		_w5895_
	);
	LUT3 #(
		.INIT('h02)
	) name5363 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		_w5896_
	);
	LUT3 #(
		.INIT('h67)
	) name5364 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w5897_
	);
	LUT2 #(
		.INIT('h2)
	) name5365 (
		_w5896_,
		_w5897_,
		_w5898_
	);
	LUT3 #(
		.INIT('h40)
	) name5366 (
		\sa01_reg[2]/P0001 ,
		_w4701_,
		_w4787_,
		_w5899_
	);
	LUT3 #(
		.INIT('h01)
	) name5367 (
		_w5385_,
		_w5899_,
		_w5898_,
		_w5900_
	);
	LUT3 #(
		.INIT('h45)
	) name5368 (
		\sa01_reg[1]/P0001 ,
		_w5895_,
		_w5900_,
		_w5901_
	);
	LUT4 #(
		.INIT('hdeff)
	) name5369 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		_w4708_,
		_w5902_
	);
	LUT4 #(
		.INIT('h153f)
	) name5370 (
		_w4699_,
		_w4775_,
		_w4784_,
		_w5361_,
		_w5903_
	);
	LUT3 #(
		.INIT('h2a)
	) name5371 (
		\sa01_reg[1]/P0001 ,
		_w5902_,
		_w5903_,
		_w5904_
	);
	LUT2 #(
		.INIT('h8)
	) name5372 (
		_w4734_,
		_w4712_,
		_w5905_
	);
	LUT4 #(
		.INIT('h3320)
	) name5373 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[2]/P0001 ,
		_w5638_,
		_w5888_,
		_w5906_
	);
	LUT2 #(
		.INIT('h1)
	) name5374 (
		_w5905_,
		_w5906_,
		_w5907_
	);
	LUT2 #(
		.INIT('h4)
	) name5375 (
		_w5904_,
		_w5907_,
		_w5908_
	);
	LUT4 #(
		.INIT('h0100)
	) name5376 (
		_w5879_,
		_w5893_,
		_w5901_,
		_w5908_,
		_w5909_
	);
	LUT3 #(
		.INIT('hb4)
	) name5377 (
		_w5599_,
		_w5642_,
		_w5909_,
		_w5910_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name5378 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5911_
	);
	LUT3 #(
		.INIT('h8a)
	) name5379 (
		\sa30_reg[2]/P0001 ,
		_w5179_,
		_w5911_,
		_w5912_
	);
	LUT3 #(
		.INIT('h10)
	) name5380 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5913_
	);
	LUT4 #(
		.INIT('h0100)
	) name5381 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5914_
	);
	LUT2 #(
		.INIT('h8)
	) name5382 (
		_w5041_,
		_w5914_,
		_w5915_
	);
	LUT3 #(
		.INIT('h8a)
	) name5383 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5916_
	);
	LUT4 #(
		.INIT('h0010)
	) name5384 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5917_
	);
	LUT3 #(
		.INIT('h0d)
	) name5385 (
		_w5036_,
		_w5916_,
		_w5917_,
		_w5918_
	);
	LUT4 #(
		.INIT('h5455)
	) name5386 (
		\sa30_reg[1]/P0001 ,
		_w5915_,
		_w5912_,
		_w5918_,
		_w5919_
	);
	LUT3 #(
		.INIT('h0b)
	) name5387 (
		\sa30_reg[6]/NET0131 ,
		_w5031_,
		_w5542_,
		_w5920_
	);
	LUT3 #(
		.INIT('h2a)
	) name5388 (
		\sa30_reg[2]/P0001 ,
		_w5136_,
		_w5920_,
		_w5921_
	);
	LUT4 #(
		.INIT('h4041)
	) name5389 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5922_
	);
	LUT3 #(
		.INIT('ha8)
	) name5390 (
		\sa30_reg[1]/P0001 ,
		_w5171_,
		_w5922_,
		_w5923_
	);
	LUT4 #(
		.INIT('h8000)
	) name5391 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5924_
	);
	LUT4 #(
		.INIT('h0040)
	) name5392 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5925_
	);
	LUT3 #(
		.INIT('h54)
	) name5393 (
		\sa30_reg[2]/P0001 ,
		_w5924_,
		_w5925_,
		_w5926_
	);
	LUT3 #(
		.INIT('h20)
	) name5394 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5927_
	);
	LUT3 #(
		.INIT('h54)
	) name5395 (
		\sa30_reg[2]/P0001 ,
		_w5106_,
		_w5927_,
		_w5928_
	);
	LUT4 #(
		.INIT('h0040)
	) name5396 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5929_
	);
	LUT3 #(
		.INIT('h0b)
	) name5397 (
		\sa30_reg[6]/NET0131 ,
		_w5158_,
		_w5929_,
		_w5930_
	);
	LUT4 #(
		.INIT('h0100)
	) name5398 (
		_w5923_,
		_w5928_,
		_w5926_,
		_w5930_,
		_w5931_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5399 (
		\sa30_reg[0]/P0002 ,
		_w5919_,
		_w5921_,
		_w5931_,
		_w5932_
	);
	LUT4 #(
		.INIT('h0027)
	) name5400 (
		\sa30_reg[6]/NET0131 ,
		_w5059_,
		_w5031_,
		_w5154_,
		_w5933_
	);
	LUT2 #(
		.INIT('h4)
	) name5401 (
		\sa30_reg[1]/P0001 ,
		\sa30_reg[2]/P0001 ,
		_w5934_
	);
	LUT4 #(
		.INIT('h4c00)
	) name5402 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5935_
	);
	LUT3 #(
		.INIT('h08)
	) name5403 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w5936_
	);
	LUT3 #(
		.INIT('hb9)
	) name5404 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5937_
	);
	LUT4 #(
		.INIT('h7707)
	) name5405 (
		_w5934_,
		_w5935_,
		_w5936_,
		_w5937_,
		_w5938_
	);
	LUT3 #(
		.INIT('he0)
	) name5406 (
		\sa30_reg[2]/P0001 ,
		_w5933_,
		_w5938_,
		_w5939_
	);
	LUT4 #(
		.INIT('hbfef)
	) name5407 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5940_
	);
	LUT4 #(
		.INIT('haf8c)
	) name5408 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		_w5013_,
		_w5940_,
		_w5941_
	);
	LUT2 #(
		.INIT('h8)
	) name5409 (
		_w5006_,
		_w5112_,
		_w5942_
	);
	LUT4 #(
		.INIT('hfff8)
	) name5410 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5943_
	);
	LUT4 #(
		.INIT('h0100)
	) name5411 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5944_
	);
	LUT3 #(
		.INIT('h10)
	) name5412 (
		_w5564_,
		_w5944_,
		_w5943_,
		_w5945_
	);
	LUT4 #(
		.INIT('h4e44)
	) name5413 (
		\sa30_reg[1]/P0001 ,
		_w5941_,
		_w5942_,
		_w5945_,
		_w5946_
	);
	LUT3 #(
		.INIT('h15)
	) name5414 (
		\sa30_reg[0]/P0002 ,
		_w5939_,
		_w5946_,
		_w5947_
	);
	LUT4 #(
		.INIT('hbbef)
	) name5415 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5948_
	);
	LUT4 #(
		.INIT('h0010)
	) name5416 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5949_
	);
	LUT4 #(
		.INIT('h5501)
	) name5417 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5948_,
		_w5949_,
		_w5950_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name5418 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5068_,
		_w5154_,
		_w5951_
	);
	LUT4 #(
		.INIT('h0040)
	) name5419 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5952_
	);
	LUT2 #(
		.INIT('h8)
	) name5420 (
		_w5036_,
		_w5952_,
		_w5953_
	);
	LUT4 #(
		.INIT('h0001)
	) name5421 (
		_w5114_,
		_w5950_,
		_w5953_,
		_w5951_,
		_w5954_
	);
	LUT3 #(
		.INIT('he4)
	) name5422 (
		\sa30_reg[2]/P0001 ,
		_w5031_,
		_w5008_,
		_w5955_
	);
	LUT4 #(
		.INIT('hffde)
	) name5423 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5956_
	);
	LUT4 #(
		.INIT('h4055)
	) name5424 (
		\sa30_reg[7]/P0001 ,
		_w5164_,
		_w5567_,
		_w5956_,
		_w5957_
	);
	LUT4 #(
		.INIT('h8daf)
	) name5425 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w5564_,
		_w5929_,
		_w5958_
	);
	LUT4 #(
		.INIT('h5700)
	) name5426 (
		\sa30_reg[1]/P0001 ,
		_w5955_,
		_w5957_,
		_w5958_,
		_w5959_
	);
	LUT3 #(
		.INIT('he0)
	) name5427 (
		\sa30_reg[1]/P0001 ,
		_w5954_,
		_w5959_,
		_w5960_
	);
	LUT3 #(
		.INIT('h10)
	) name5428 (
		_w5932_,
		_w5947_,
		_w5960_,
		_w5961_
	);
	LUT2 #(
		.INIT('h1)
	) name5429 (
		_w5571_,
		_w5952_,
		_w5962_
	);
	LUT3 #(
		.INIT('h10)
	) name5430 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5963_
	);
	LUT2 #(
		.INIT('h8)
	) name5431 (
		_w5164_,
		_w5963_,
		_w5964_
	);
	LUT4 #(
		.INIT('h4404)
	) name5432 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5965_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name5433 (
		_w5040_,
		_w5109_,
		_w5525_,
		_w5965_,
		_w5966_
	);
	LUT4 #(
		.INIT('h4555)
	) name5434 (
		\sa30_reg[1]/P0001 ,
		_w5964_,
		_w5962_,
		_w5966_,
		_w5967_
	);
	LUT4 #(
		.INIT('ha7f7)
	) name5435 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5968_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name5436 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		_w5060_,
		_w5968_,
		_w5969_
	);
	LUT4 #(
		.INIT('hcfca)
	) name5437 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5970_
	);
	LUT3 #(
		.INIT('h02)
	) name5438 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5971_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name5439 (
		_w5143_,
		_w5184_,
		_w5971_,
		_w5970_,
		_w5972_
	);
	LUT4 #(
		.INIT('haabf)
	) name5440 (
		\sa30_reg[5]/P0001 ,
		_w5007_,
		_w5117_,
		_w5564_,
		_w5973_
	);
	LUT2 #(
		.INIT('h8)
	) name5441 (
		_w5041_,
		_w5109_,
		_w5974_
	);
	LUT3 #(
		.INIT('h13)
	) name5442 (
		_w5014_,
		_w5925_,
		_w5936_,
		_w5975_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5443 (
		\sa30_reg[1]/P0001 ,
		_w5973_,
		_w5974_,
		_w5975_,
		_w5976_
	);
	LUT4 #(
		.INIT('h0100)
	) name5444 (
		_w5967_,
		_w5969_,
		_w5972_,
		_w5976_,
		_w5977_
	);
	LUT3 #(
		.INIT('h54)
	) name5445 (
		\sa30_reg[2]/P0001 ,
		_w5552_,
		_w5578_,
		_w5978_
	);
	LUT4 #(
		.INIT('h0800)
	) name5446 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5979_
	);
	LUT4 #(
		.INIT('h0777)
	) name5447 (
		_w5040_,
		_w5021_,
		_w5164_,
		_w5567_,
		_w5980_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5448 (
		\sa30_reg[1]/P0001 ,
		_w5978_,
		_w5979_,
		_w5980_,
		_w5981_
	);
	LUT4 #(
		.INIT('h4000)
	) name5449 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5982_
	);
	LUT2 #(
		.INIT('h1)
	) name5450 (
		_w5917_,
		_w5982_,
		_w5983_
	);
	LUT4 #(
		.INIT('h0002)
	) name5451 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5984_
	);
	LUT3 #(
		.INIT('h0b)
	) name5452 (
		\sa30_reg[7]/P0001 ,
		_w5095_,
		_w5984_,
		_w5985_
	);
	LUT3 #(
		.INIT('h15)
	) name5453 (
		\sa30_reg[2]/P0001 ,
		_w5983_,
		_w5985_,
		_w5986_
	);
	LUT4 #(
		.INIT('hf2fa)
	) name5454 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		_w5987_
	);
	LUT2 #(
		.INIT('h2)
	) name5455 (
		\sa30_reg[7]/P0001 ,
		_w5987_,
		_w5988_
	);
	LUT3 #(
		.INIT('h07)
	) name5456 (
		_w5112_,
		_w5544_,
		_w5549_,
		_w5989_
	);
	LUT4 #(
		.INIT('h0008)
	) name5457 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5990_
	);
	LUT4 #(
		.INIT('h7ff6)
	) name5458 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5991_
	);
	LUT2 #(
		.INIT('h2)
	) name5459 (
		_w5112_,
		_w5991_,
		_w5992_
	);
	LUT4 #(
		.INIT('h00ba)
	) name5460 (
		\sa30_reg[1]/P0001 ,
		_w5988_,
		_w5989_,
		_w5992_,
		_w5993_
	);
	LUT3 #(
		.INIT('h10)
	) name5461 (
		_w5986_,
		_w5981_,
		_w5993_,
		_w5994_
	);
	LUT4 #(
		.INIT('h0004)
	) name5462 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5995_
	);
	LUT4 #(
		.INIT('hadfb)
	) name5463 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5996_
	);
	LUT4 #(
		.INIT('h0302)
	) name5464 (
		\sa30_reg[3]/P0001 ,
		_w5084_,
		_w5019_,
		_w5996_,
		_w5997_
	);
	LUT2 #(
		.INIT('h2)
	) name5465 (
		_w5184_,
		_w5997_,
		_w5998_
	);
	LUT4 #(
		.INIT('hbdff)
	) name5466 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5999_
	);
	LUT3 #(
		.INIT('h10)
	) name5467 (
		_w5917_,
		_w5982_,
		_w5999_,
		_w6000_
	);
	LUT3 #(
		.INIT('h51)
	) name5468 (
		\sa30_reg[1]/P0001 ,
		\sa30_reg[2]/P0001 ,
		_w5031_,
		_w6001_
	);
	LUT2 #(
		.INIT('h4)
	) name5469 (
		_w6000_,
		_w6001_,
		_w6002_
	);
	LUT4 #(
		.INIT('h4000)
	) name5470 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w6003_
	);
	LUT4 #(
		.INIT('h0023)
	) name5471 (
		\sa30_reg[5]/P0001 ,
		_w5065_,
		_w5564_,
		_w6003_,
		_w6004_
	);
	LUT2 #(
		.INIT('h2)
	) name5472 (
		_w5934_,
		_w6004_,
		_w6005_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name5473 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6006_
	);
	LUT3 #(
		.INIT('h20)
	) name5474 (
		\sa30_reg[1]/P0001 ,
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		_w6007_
	);
	LUT2 #(
		.INIT('h4)
	) name5475 (
		_w6006_,
		_w6007_,
		_w6008_
	);
	LUT4 #(
		.INIT('hcecf)
	) name5476 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5068_,
		_w5552_,
		_w6009_
	);
	LUT3 #(
		.INIT('h32)
	) name5477 (
		\sa30_reg[2]/P0001 ,
		_w6008_,
		_w6009_,
		_w6010_
	);
	LUT4 #(
		.INIT('h0100)
	) name5478 (
		_w6005_,
		_w6002_,
		_w5998_,
		_w6010_,
		_w6011_
	);
	LUT4 #(
		.INIT('he400)
	) name5479 (
		\sa30_reg[0]/P0002 ,
		_w5994_,
		_w5977_,
		_w6011_,
		_w6012_
	);
	LUT4 #(
		.INIT('h0015)
	) name5480 (
		\sa23_reg[1]/P0001 ,
		_w4890_,
		_w4903_,
		_w5742_,
		_w6013_
	);
	LUT4 #(
		.INIT('h0080)
	) name5481 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w6014_
	);
	LUT3 #(
		.INIT('h0d)
	) name5482 (
		_w4892_,
		_w5700_,
		_w6014_,
		_w6015_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5483 (
		\sa23_reg[2]/P0001 ,
		_w5286_,
		_w5277_,
		_w5510_,
		_w6016_
	);
	LUT4 #(
		.INIT('h020a)
	) name5484 (
		\sa23_reg[1]/P0001 ,
		_w4896_,
		_w4933_,
		_w5259_,
		_w6017_
	);
	LUT4 #(
		.INIT('h7077)
	) name5485 (
		_w6013_,
		_w6015_,
		_w6016_,
		_w6017_,
		_w6018_
	);
	LUT4 #(
		.INIT('h5554)
	) name5486 (
		\sa23_reg[2]/P0001 ,
		_w5279_,
		_w5466_,
		_w5742_,
		_w6019_
	);
	LUT2 #(
		.INIT('h2)
	) name5487 (
		_w4906_,
		_w5495_,
		_w6020_
	);
	LUT3 #(
		.INIT('h8a)
	) name5488 (
		\sa23_reg[0]/P0001 ,
		_w4918_,
		_w4997_,
		_w6021_
	);
	LUT3 #(
		.INIT('h10)
	) name5489 (
		_w6019_,
		_w6020_,
		_w6021_,
		_w6022_
	);
	LUT2 #(
		.INIT('h4)
	) name5490 (
		_w6018_,
		_w6022_,
		_w6023_
	);
	LUT4 #(
		.INIT('h0015)
	) name5491 (
		\sa23_reg[2]/P0001 ,
		_w4905_,
		_w4981_,
		_w5278_,
		_w6024_
	);
	LUT3 #(
		.INIT('h02)
	) name5492 (
		\sa23_reg[2]/P0001 ,
		_w5287_,
		_w5466_,
		_w6025_
	);
	LUT3 #(
		.INIT('h45)
	) name5493 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w5307_,
		_w6026_
	);
	LUT4 #(
		.INIT('h5400)
	) name5494 (
		_w5484_,
		_w6024_,
		_w6025_,
		_w6026_,
		_w6027_
	);
	LUT4 #(
		.INIT('h5554)
	) name5495 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w6028_
	);
	LUT3 #(
		.INIT('h10)
	) name5496 (
		_w4914_,
		_w5307_,
		_w6028_,
		_w6029_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name5497 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w6030_
	);
	LUT2 #(
		.INIT('h4)
	) name5498 (
		_w5734_,
		_w6030_,
		_w6031_
	);
	LUT4 #(
		.INIT('h0002)
	) name5499 (
		\sa23_reg[1]/P0001 ,
		_w4909_,
		_w4976_,
		_w4977_,
		_w6032_
	);
	LUT3 #(
		.INIT('he0)
	) name5500 (
		_w6029_,
		_w6031_,
		_w6032_,
		_w6033_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5501 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w6034_
	);
	LUT2 #(
		.INIT('h4)
	) name5502 (
		_w5306_,
		_w6034_,
		_w6035_
	);
	LUT2 #(
		.INIT('h1)
	) name5503 (
		\sa23_reg[2]/P0001 ,
		_w4994_,
		_w6036_
	);
	LUT4 #(
		.INIT('h153f)
	) name5504 (
		\sa23_reg[6]/NET0131 ,
		_w4890_,
		_w4937_,
		_w5254_,
		_w6037_
	);
	LUT3 #(
		.INIT('h15)
	) name5505 (
		\sa23_reg[0]/P0001 ,
		_w4918_,
		_w4997_,
		_w6038_
	);
	LUT4 #(
		.INIT('hea00)
	) name5506 (
		_w6035_,
		_w6036_,
		_w6037_,
		_w6038_,
		_w6039_
	);
	LUT3 #(
		.INIT('he0)
	) name5507 (
		_w6027_,
		_w6033_,
		_w6039_,
		_w6040_
	);
	LUT3 #(
		.INIT('h15)
	) name5508 (
		\sa23_reg[1]/P0001 ,
		_w4910_,
		_w4957_,
		_w6041_
	);
	LUT4 #(
		.INIT('h0007)
	) name5509 (
		_w4894_,
		_w4927_,
		_w4994_,
		_w5711_,
		_w6042_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name5510 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6043_
	);
	LUT4 #(
		.INIT('h8a02)
	) name5511 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[3]/P0001 ,
		_w4967_,
		_w6043_,
		_w6044_
	);
	LUT4 #(
		.INIT('h135f)
	) name5512 (
		_w4908_,
		_w4919_,
		_w4930_,
		_w5259_,
		_w6045_
	);
	LUT4 #(
		.INIT('hf800)
	) name5513 (
		_w6041_,
		_w6042_,
		_w6044_,
		_w6045_,
		_w6046_
	);
	LUT4 #(
		.INIT('h0007)
	) name5514 (
		_w4919_,
		_w4959_,
		_w5254_,
		_w5723_,
		_w6047_
	);
	LUT3 #(
		.INIT('h40)
	) name5515 (
		_w5480_,
		_w6041_,
		_w6047_,
		_w6048_
	);
	LUT3 #(
		.INIT('h0e)
	) name5516 (
		_w4890_,
		_w4936_,
		_w4937_,
		_w6049_
	);
	LUT3 #(
		.INIT('h02)
	) name5517 (
		\sa23_reg[1]/P0001 ,
		_w4909_,
		_w5262_,
		_w6050_
	);
	LUT2 #(
		.INIT('h4)
	) name5518 (
		_w6049_,
		_w6050_,
		_w6051_
	);
	LUT4 #(
		.INIT('hddd8)
	) name5519 (
		\sa23_reg[2]/P0001 ,
		_w6046_,
		_w6051_,
		_w6048_,
		_w6052_
	);
	LUT3 #(
		.INIT('he0)
	) name5520 (
		_w6023_,
		_w6040_,
		_w6052_,
		_w6053_
	);
	LUT4 #(
		.INIT('ha955)
	) name5521 (
		\u0_w_reg[1][1]/P0001 ,
		_w6023_,
		_w6040_,
		_w6052_,
		_w6054_
	);
	LUT3 #(
		.INIT('h69)
	) name5522 (
		_w5961_,
		_w6012_,
		_w6054_,
		_w6055_
	);
	LUT4 #(
		.INIT('h1441)
	) name5523 (
		\ld_r_reg/P0001 ,
		_w5862_,
		_w5910_,
		_w6055_,
		_w6056_
	);
	LUT3 #(
		.INIT('h28)
	) name5524 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[65]/P0001 ,
		\u0_w_reg[1][1]/P0001 ,
		_w6057_
	);
	LUT2 #(
		.INIT('he)
	) name5525 (
		_w6056_,
		_w6057_,
		_w6058_
	);
	LUT4 #(
		.INIT('h6996)
	) name5526 (
		\u0_w_reg[1][28]/P0001 ,
		_w4691_,
		_w5517_,
		_w5580_,
		_w6059_
	);
	LUT4 #(
		.INIT('hd1ff)
	) name5527 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w6060_
	);
	LUT3 #(
		.INIT('h8a)
	) name5528 (
		\sa01_reg[2]/P0001 ,
		_w5337_,
		_w6060_,
		_w6061_
	);
	LUT4 #(
		.INIT('h0051)
	) name5529 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w6062_
	);
	LUT4 #(
		.INIT('h2223)
	) name5530 (
		_w4757_,
		_w4758_,
		_w5368_,
		_w6062_,
		_w6063_
	);
	LUT3 #(
		.INIT('h8a)
	) name5531 (
		\sa01_reg[1]/P0001 ,
		_w6061_,
		_w6063_,
		_w6064_
	);
	LUT3 #(
		.INIT('h01)
	) name5532 (
		\sa01_reg[2]/P0001 ,
		_w4790_,
		_w5617_,
		_w6065_
	);
	LUT4 #(
		.INIT('haa2a)
	) name5533 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w6066_
	);
	LUT2 #(
		.INIT('h4)
	) name5534 (
		_w5326_,
		_w6066_,
		_w6067_
	);
	LUT4 #(
		.INIT('h0007)
	) name5535 (
		_w4775_,
		_w4784_,
		_w4794_,
		_w5439_,
		_w6068_
	);
	LUT4 #(
		.INIT('h5400)
	) name5536 (
		_w5847_,
		_w6065_,
		_w6067_,
		_w6068_,
		_w6069_
	);
	LUT4 #(
		.INIT('h0007)
	) name5537 (
		_w4698_,
		_w4693_,
		_w5602_,
		_w5880_,
		_w6070_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name5538 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w6071_
	);
	LUT4 #(
		.INIT('h5f13)
	) name5539 (
		_w4701_,
		_w4772_,
		_w4787_,
		_w6071_,
		_w6072_
	);
	LUT3 #(
		.INIT('he0)
	) name5540 (
		\sa01_reg[2]/P0001 ,
		_w6070_,
		_w6072_,
		_w6073_
	);
	LUT4 #(
		.INIT('h0e00)
	) name5541 (
		\sa01_reg[1]/P0001 ,
		_w6069_,
		_w6064_,
		_w6073_,
		_w6074_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name5542 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w5369_,
		_w5426_,
		_w6075_
	);
	LUT2 #(
		.INIT('h8)
	) name5543 (
		_w4745_,
		_w4693_,
		_w6076_
	);
	LUT3 #(
		.INIT('h13)
	) name5544 (
		_w4704_,
		_w4754_,
		_w4749_,
		_w6077_
	);
	LUT4 #(
		.INIT('h0100)
	) name5545 (
		_w4766_,
		_w6075_,
		_w6076_,
		_w6077_,
		_w6078_
	);
	LUT4 #(
		.INIT('h0008)
	) name5546 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w6079_
	);
	LUT4 #(
		.INIT('h0007)
	) name5547 (
		_w4743_,
		_w5450_,
		_w5602_,
		_w6079_,
		_w6080_
	);
	LUT3 #(
		.INIT('h07)
	) name5548 (
		_w4729_,
		_w5353_,
		_w5443_,
		_w6081_
	);
	LUT2 #(
		.INIT('h8)
	) name5549 (
		_w6080_,
		_w6081_,
		_w6082_
	);
	LUT4 #(
		.INIT('h5540)
	) name5550 (
		\sa01_reg[2]/P0001 ,
		_w4698_,
		_w4749_,
		_w4705_,
		_w6083_
	);
	LUT2 #(
		.INIT('h8)
	) name5551 (
		_w4775_,
		_w5369_,
		_w6084_
	);
	LUT4 #(
		.INIT('h153f)
	) name5552 (
		\sa01_reg[2]/P0001 ,
		_w4718_,
		_w4801_,
		_w5436_,
		_w6085_
	);
	LUT3 #(
		.INIT('h10)
	) name5553 (
		_w6083_,
		_w6084_,
		_w6085_,
		_w6086_
	);
	LUT4 #(
		.INIT('he400)
	) name5554 (
		\sa01_reg[1]/P0001 ,
		_w6082_,
		_w6078_,
		_w6086_,
		_w6087_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name5555 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w6088_
	);
	LUT2 #(
		.INIT('h2)
	) name5556 (
		_w5610_,
		_w6088_,
		_w6089_
	);
	LUT3 #(
		.INIT('h40)
	) name5557 (
		\sa01_reg[2]/P0001 ,
		_w4697_,
		_w4751_,
		_w6090_
	);
	LUT4 #(
		.INIT('h2777)
	) name5558 (
		\sa01_reg[2]/P0001 ,
		_w4743_,
		_w4697_,
		_w4751_,
		_w6091_
	);
	LUT3 #(
		.INIT('h8a)
	) name5559 (
		\sa01_reg[1]/P0001 ,
		_w6089_,
		_w6091_,
		_w6092_
	);
	LUT4 #(
		.INIT('h0777)
	) name5560 (
		_w4698_,
		_w4709_,
		_w4718_,
		_w4801_,
		_w6093_
	);
	LUT2 #(
		.INIT('h2)
	) name5561 (
		_w5407_,
		_w6093_,
		_w6094_
	);
	LUT2 #(
		.INIT('h8)
	) name5562 (
		_w4739_,
		_w5856_,
		_w6095_
	);
	LUT4 #(
		.INIT('h135f)
	) name5563 (
		_w4704_,
		_w4716_,
		_w5361_,
		_w5438_,
		_w6096_
	);
	LUT4 #(
		.INIT('h2000)
	) name5564 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w6097_
	);
	LUT3 #(
		.INIT('hc8)
	) name5565 (
		_w4758_,
		_w5442_,
		_w6097_,
		_w6098_
	);
	LUT3 #(
		.INIT('h80)
	) name5566 (
		\sa01_reg[7]/NET0131 ,
		_w4723_,
		_w5613_,
		_w6099_
	);
	LUT4 #(
		.INIT('h0100)
	) name5567 (
		_w6095_,
		_w6098_,
		_w6099_,
		_w6096_,
		_w6100_
	);
	LUT3 #(
		.INIT('h10)
	) name5568 (
		_w6092_,
		_w6094_,
		_w6100_,
		_w6101_
	);
	LUT4 #(
		.INIT('he400)
	) name5569 (
		\sa01_reg[0]/P0001 ,
		_w6087_,
		_w6074_,
		_w6101_,
		_w6102_
	);
	LUT3 #(
		.INIT('h4b)
	) name5570 (
		_w5599_,
		_w5642_,
		_w6102_,
		_w6103_
	);
	LUT3 #(
		.INIT('h32)
	) name5571 (
		_w4618_,
		_w4611_,
		_w4854_,
		_w6104_
	);
	LUT4 #(
		.INIT('hefdf)
	) name5572 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6105_
	);
	LUT2 #(
		.INIT('h1)
	) name5573 (
		\sa12_reg[2]/P0001 ,
		_w6105_,
		_w6106_
	);
	LUT3 #(
		.INIT('h01)
	) name5574 (
		_w4634_,
		_w4813_,
		_w4872_,
		_w6107_
	);
	LUT4 #(
		.INIT('h5455)
	) name5575 (
		\sa12_reg[1]/P0001 ,
		_w6106_,
		_w6104_,
		_w6107_,
		_w6108_
	);
	LUT4 #(
		.INIT('hd1ff)
	) name5576 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6109_
	);
	LUT3 #(
		.INIT('h8a)
	) name5577 (
		\sa12_reg[2]/P0001 ,
		_w5796_,
		_w6109_,
		_w6110_
	);
	LUT4 #(
		.INIT('h0051)
	) name5578 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6111_
	);
	LUT4 #(
		.INIT('h2223)
	) name5579 (
		_w4608_,
		_w4621_,
		_w4602_,
		_w6111_,
		_w6112_
	);
	LUT3 #(
		.INIT('h8a)
	) name5580 (
		\sa12_reg[1]/P0001 ,
		_w6110_,
		_w6112_,
		_w6113_
	);
	LUT4 #(
		.INIT('h8000)
	) name5581 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6114_
	);
	LUT3 #(
		.INIT('h07)
	) name5582 (
		\sa12_reg[7]/NET0131 ,
		_w4807_,
		_w6114_,
		_w6115_
	);
	LUT4 #(
		.INIT('h0007)
	) name5583 (
		\sa12_reg[7]/NET0131 ,
		_w4807_,
		_w5655_,
		_w6114_,
		_w6116_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name5584 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6117_
	);
	LUT4 #(
		.INIT('haf23)
	) name5585 (
		\sa12_reg[7]/NET0131 ,
		_w4642_,
		_w4668_,
		_w6117_,
		_w6118_
	);
	LUT3 #(
		.INIT('he0)
	) name5586 (
		\sa12_reg[2]/P0001 ,
		_w6116_,
		_w6118_,
		_w6119_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5587 (
		\sa12_reg[0]/P0001 ,
		_w6113_,
		_w6108_,
		_w6119_,
		_w6120_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name5588 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4823_,
		_w4875_,
		_w6121_
	);
	LUT4 #(
		.INIT('h008a)
	) name5589 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4675_,
		_w4618_,
		_w6122_
	);
	LUT4 #(
		.INIT('h135f)
	) name5590 (
		_w4608_,
		_w4659_,
		_w4602_,
		_w5683_,
		_w6123_
	);
	LUT3 #(
		.INIT('h40)
	) name5591 (
		_w6121_,
		_w6122_,
		_w6123_,
		_w6124_
	);
	LUT4 #(
		.INIT('h5400)
	) name5592 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6125_
	);
	LUT3 #(
		.INIT('ha8)
	) name5593 (
		\sa12_reg[2]/P0001 ,
		_w4606_,
		_w6125_,
		_w6126_
	);
	LUT3 #(
		.INIT('h01)
	) name5594 (
		\sa12_reg[1]/P0001 ,
		_w5239_,
		_w5655_,
		_w6127_
	);
	LUT3 #(
		.INIT('h10)
	) name5595 (
		_w5245_,
		_w6126_,
		_w6127_,
		_w6128_
	);
	LUT4 #(
		.INIT('h5150)
	) name5596 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		_w4638_,
		_w4846_,
		_w6129_
	);
	LUT2 #(
		.INIT('h4)
	) name5597 (
		\sa12_reg[4]/P0001 ,
		_w4822_,
		_w6130_
	);
	LUT4 #(
		.INIT('h0002)
	) name5598 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w6131_
	);
	LUT3 #(
		.INIT('ha8)
	) name5599 (
		\sa12_reg[2]/P0001 ,
		_w5232_,
		_w6131_,
		_w6132_
	);
	LUT3 #(
		.INIT('h01)
	) name5600 (
		_w6130_,
		_w6129_,
		_w6132_,
		_w6133_
	);
	LUT4 #(
		.INIT('h0155)
	) name5601 (
		\sa12_reg[0]/P0001 ,
		_w6124_,
		_w6128_,
		_w6133_,
		_w6134_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name5602 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6135_
	);
	LUT2 #(
		.INIT('h2)
	) name5603 (
		_w5202_,
		_w6135_,
		_w6136_
	);
	LUT3 #(
		.INIT('h10)
	) name5604 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4679_,
		_w6137_
	);
	LUT4 #(
		.INIT('hcdef)
	) name5605 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w4679_,
		_w4602_,
		_w6138_
	);
	LUT3 #(
		.INIT('h8a)
	) name5606 (
		\sa12_reg[1]/P0001 ,
		_w6136_,
		_w6138_,
		_w6139_
	);
	LUT4 #(
		.INIT('h153f)
	) name5607 (
		_w4635_,
		_w4821_,
		_w4860_,
		_w5239_,
		_w6140_
	);
	LUT2 #(
		.INIT('h1)
	) name5608 (
		\sa12_reg[1]/P0001 ,
		_w6140_,
		_w6141_
	);
	LUT4 #(
		.INIT('h2e3f)
	) name5609 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[2]/P0001 ,
		_w4621_,
		_w4609_,
		_w6142_
	);
	LUT2 #(
		.INIT('h1)
	) name5610 (
		\sa12_reg[4]/P0001 ,
		_w6142_,
		_w6143_
	);
	LUT3 #(
		.INIT('he0)
	) name5611 (
		_w4668_,
		_w4621_,
		_w5237_,
		_w6144_
	);
	LUT3 #(
		.INIT('h01)
	) name5612 (
		_w5766_,
		_w5808_,
		_w6144_,
		_w6145_
	);
	LUT4 #(
		.INIT('h0100)
	) name5613 (
		_w6143_,
		_w6141_,
		_w6139_,
		_w6145_,
		_w6146_
	);
	LUT3 #(
		.INIT('h10)
	) name5614 (
		_w6134_,
		_w6120_,
		_w6146_,
		_w6147_
	);
	LUT2 #(
		.INIT('h9)
	) name5615 (
		_w5695_,
		_w6147_,
		_w6148_
	);
	LUT4 #(
		.INIT('h4114)
	) name5616 (
		\ld_r_reg/P0001 ,
		_w6059_,
		_w6103_,
		_w6148_,
		_w6149_
	);
	LUT3 #(
		.INIT('h82)
	) name5617 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[92]/P0001 ,
		\u0_w_reg[1][28]/P0001 ,
		_w6150_
	);
	LUT2 #(
		.INIT('h1)
	) name5618 (
		_w6149_,
		_w6150_,
		_w6151_
	);
	LUT2 #(
		.INIT('h1)
	) name5619 (
		\sa23_reg[1]/P0001 ,
		_w5476_,
		_w6152_
	);
	LUT3 #(
		.INIT('h20)
	) name5620 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w6153_
	);
	LUT4 #(
		.INIT('h2237)
	) name5621 (
		_w4919_,
		_w4944_,
		_w4992_,
		_w6153_,
		_w6154_
	);
	LUT3 #(
		.INIT('h40)
	) name5622 (
		_w5312_,
		_w6152_,
		_w6154_,
		_w6155_
	);
	LUT4 #(
		.INIT('h008a)
	) name5623 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[3]/P0001 ,
		_w4921_,
		_w4949_,
		_w6156_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name5624 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w5259_,
		_w5721_,
		_w6157_
	);
	LUT2 #(
		.INIT('h8)
	) name5625 (
		_w6156_,
		_w6157_,
		_w6158_
	);
	LUT4 #(
		.INIT('h0015)
	) name5626 (
		\sa23_reg[2]/P0001 ,
		_w4894_,
		_w4927_,
		_w4982_,
		_w6159_
	);
	LUT4 #(
		.INIT('haa80)
	) name5627 (
		\sa23_reg[1]/P0001 ,
		_w4927_,
		_w4951_,
		_w5297_,
		_w6160_
	);
	LUT4 #(
		.INIT('h0002)
	) name5628 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w6161_
	);
	LUT3 #(
		.INIT('h02)
	) name5629 (
		\sa23_reg[2]/P0001 ,
		_w4921_,
		_w6161_,
		_w6162_
	);
	LUT4 #(
		.INIT('h4544)
	) name5630 (
		_w4965_,
		_w6159_,
		_w6160_,
		_w6162_,
		_w6163_
	);
	LUT4 #(
		.INIT('h0155)
	) name5631 (
		\sa23_reg[0]/P0001 ,
		_w6155_,
		_w6158_,
		_w6163_,
		_w6164_
	);
	LUT3 #(
		.INIT('h10)
	) name5632 (
		_w4978_,
		_w4949_,
		_w5460_,
		_w6165_
	);
	LUT3 #(
		.INIT('h01)
	) name5633 (
		\sa23_reg[2]/P0001 ,
		_w4906_,
		_w5723_,
		_w6166_
	);
	LUT4 #(
		.INIT('h0013)
	) name5634 (
		_w4919_,
		_w4994_,
		_w5259_,
		_w5281_,
		_w6167_
	);
	LUT4 #(
		.INIT('h0155)
	) name5635 (
		\sa23_reg[1]/P0001 ,
		_w6165_,
		_w6166_,
		_w6167_,
		_w6168_
	);
	LUT4 #(
		.INIT('hf3fb)
	) name5636 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6169_
	);
	LUT3 #(
		.INIT('h8a)
	) name5637 (
		\sa23_reg[2]/P0001 ,
		_w5718_,
		_w6169_,
		_w6170_
	);
	LUT4 #(
		.INIT('h0010)
	) name5638 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6171_
	);
	LUT2 #(
		.INIT('h1)
	) name5639 (
		_w5287_,
		_w6171_,
		_w6172_
	);
	LUT4 #(
		.INIT('h0001)
	) name5640 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6173_
	);
	LUT3 #(
		.INIT('h0b)
	) name5641 (
		_w4975_,
		_w5296_,
		_w6173_,
		_w6174_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5642 (
		\sa23_reg[1]/P0001 ,
		_w6170_,
		_w6172_,
		_w6174_,
		_w6175_
	);
	LUT4 #(
		.INIT('h8000)
	) name5643 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6176_
	);
	LUT4 #(
		.INIT('h0007)
	) name5644 (
		_w4890_,
		_w4937_,
		_w5476_,
		_w6176_,
		_w6177_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name5645 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6178_
	);
	LUT4 #(
		.INIT('h7707)
	) name5646 (
		_w4925_,
		_w4948_,
		_w5726_,
		_w6178_,
		_w6179_
	);
	LUT3 #(
		.INIT('he0)
	) name5647 (
		\sa23_reg[2]/P0001 ,
		_w6177_,
		_w6179_,
		_w6180_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5648 (
		\sa23_reg[0]/P0001 ,
		_w6175_,
		_w6168_,
		_w6180_,
		_w6181_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name5649 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6182_
	);
	LUT2 #(
		.INIT('h2)
	) name5650 (
		_w5252_,
		_w6182_,
		_w6183_
	);
	LUT4 #(
		.INIT('h2000)
	) name5651 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w6184_
	);
	LUT3 #(
		.INIT('ha8)
	) name5652 (
		\sa23_reg[2]/P0001 ,
		_w5287_,
		_w6184_,
		_w6185_
	);
	LUT3 #(
		.INIT('h40)
	) name5653 (
		\sa23_reg[2]/P0001 ,
		_w4945_,
		_w5510_,
		_w6186_
	);
	LUT4 #(
		.INIT('h2777)
	) name5654 (
		\sa23_reg[2]/P0001 ,
		_w4938_,
		_w4945_,
		_w5510_,
		_w6187_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5655 (
		\sa23_reg[1]/P0001 ,
		_w6185_,
		_w6183_,
		_w6187_,
		_w6188_
	);
	LUT4 #(
		.INIT('hffed)
	) name5656 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6189_
	);
	LUT4 #(
		.INIT('h5f13)
	) name5657 (
		_w4975_,
		_w5295_,
		_w5721_,
		_w6189_,
		_w6190_
	);
	LUT4 #(
		.INIT('hedff)
	) name5658 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6191_
	);
	LUT4 #(
		.INIT('haf23)
	) name5659 (
		\sa23_reg[7]/NET0131 ,
		_w4918_,
		_w5307_,
		_w6191_,
		_w6192_
	);
	LUT3 #(
		.INIT('he0)
	) name5660 (
		\sa23_reg[1]/P0001 ,
		_w6190_,
		_w6192_,
		_w6193_
	);
	LUT2 #(
		.INIT('h4)
	) name5661 (
		_w6188_,
		_w6193_,
		_w6194_
	);
	LUT3 #(
		.INIT('h10)
	) name5662 (
		_w6181_,
		_w6164_,
		_w6194_,
		_w6195_
	);
	LUT4 #(
		.INIT('h6996)
	) name5663 (
		_w4804_,
		_w5695_,
		_w6147_,
		_w6195_,
		_w6196_
	);
	LUT4 #(
		.INIT('h5655)
	) name5664 (
		\u0_w_reg[1][20]/P0001 ,
		_w5717_,
		_w5738_,
		_w5757_,
		_w6197_
	);
	LUT3 #(
		.INIT('h96)
	) name5665 (
		_w5517_,
		_w5580_,
		_w6197_,
		_w6198_
	);
	LUT3 #(
		.INIT('h82)
	) name5666 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[84]/P0001 ,
		\u0_w_reg[1][20]/P0001 ,
		_w6199_
	);
	LUT4 #(
		.INIT('h00be)
	) name5667 (
		\ld_r_reg/P0001 ,
		_w6196_,
		_w6198_,
		_w6199_,
		_w6200_
	);
	LUT4 #(
		.INIT('h9a65)
	) name5668 (
		_w4804_,
		_w4841_,
		_w4886_,
		_w5389_,
		_w6201_
	);
	LUT4 #(
		.INIT('h9a65)
	) name5669 (
		\u0_w_reg[1][5]/P0001 ,
		_w4942_,
		_w5003_,
		_w5580_,
		_w6202_
	);
	LUT3 #(
		.INIT('h28)
	) name5670 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[69]/P0001 ,
		\u0_w_reg[1][5]/P0001 ,
		_w6203_
	);
	LUT4 #(
		.INIT('hff41)
	) name5671 (
		\ld_r_reg/P0001 ,
		_w6201_,
		_w6202_,
		_w6203_,
		_w6204_
	);
	LUT4 #(
		.INIT('hff3b)
	) name5672 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6205_
	);
	LUT4 #(
		.INIT('hd8fa)
	) name5673 (
		\sa30_reg[2]/P0001 ,
		_w5008_,
		_w5578_,
		_w6205_,
		_w6206_
	);
	LUT2 #(
		.INIT('h8)
	) name5674 (
		_w5029_,
		_w5126_,
		_w6207_
	);
	LUT4 #(
		.INIT('h0105)
	) name5675 (
		_w5068_,
		_w5040_,
		_w5098_,
		_w5117_,
		_w6208_
	);
	LUT4 #(
		.INIT('h5455)
	) name5676 (
		\sa30_reg[1]/P0001 ,
		_w6206_,
		_w6207_,
		_w6208_,
		_w6209_
	);
	LUT4 #(
		.INIT('hf3fb)
	) name5677 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6210_
	);
	LUT3 #(
		.INIT('h8a)
	) name5678 (
		\sa30_reg[2]/P0001 ,
		_w5544_,
		_w6210_,
		_w6211_
	);
	LUT4 #(
		.INIT('hffac)
	) name5679 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6212_
	);
	LUT2 #(
		.INIT('h1)
	) name5680 (
		\sa30_reg[2]/P0001 ,
		_w6212_,
		_w6213_
	);
	LUT3 #(
		.INIT('h13)
	) name5681 (
		\sa30_reg[4]/P0001 ,
		_w5538_,
		_w5935_,
		_w6214_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5682 (
		\sa30_reg[1]/P0001 ,
		_w6213_,
		_w6211_,
		_w6214_,
		_w6215_
	);
	LUT4 #(
		.INIT('h0027)
	) name5683 (
		\sa30_reg[6]/NET0131 ,
		_w5059_,
		_w5031_,
		_w5132_,
		_w6216_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name5684 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6217_
	);
	LUT4 #(
		.INIT('h7707)
	) name5685 (
		_w5006_,
		_w5036_,
		_w5102_,
		_w6217_,
		_w6218_
	);
	LUT3 #(
		.INIT('he0)
	) name5686 (
		\sa30_reg[2]/P0001 ,
		_w6216_,
		_w6218_,
		_w6219_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5687 (
		\sa30_reg[0]/P0002 ,
		_w6215_,
		_w6209_,
		_w6219_,
		_w6220_
	);
	LUT4 #(
		.INIT('haa20)
	) name5688 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		_w5060_,
		_w5089_,
		_w6221_
	);
	LUT4 #(
		.INIT('h002a)
	) name5689 (
		\sa30_reg[1]/P0001 ,
		_w5005_,
		_w5072_,
		_w5008_,
		_w6222_
	);
	LUT4 #(
		.INIT('h575f)
	) name5690 (
		\sa30_reg[7]/P0001 ,
		_w5056_,
		_w5095_,
		_w5532_,
		_w6223_
	);
	LUT3 #(
		.INIT('h40)
	) name5691 (
		_w6221_,
		_w6222_,
		_w6223_,
		_w6224_
	);
	LUT4 #(
		.INIT('h0008)
	) name5692 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6225_
	);
	LUT3 #(
		.INIT('h01)
	) name5693 (
		\sa30_reg[1]/P0001 ,
		_w5132_,
		_w6225_,
		_w6226_
	);
	LUT3 #(
		.INIT('he0)
	) name5694 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6227_
	);
	LUT3 #(
		.INIT('h13)
	) name5695 (
		_w5164_,
		_w5984_,
		_w6227_,
		_w6228_
	);
	LUT3 #(
		.INIT('h40)
	) name5696 (
		_w5189_,
		_w6226_,
		_w6228_,
		_w6229_
	);
	LUT3 #(
		.INIT('ha8)
	) name5697 (
		\sa30_reg[2]/P0001 ,
		_w5107_,
		_w5176_,
		_w6230_
	);
	LUT4 #(
		.INIT('h5540)
	) name5698 (
		\sa30_reg[2]/P0001 ,
		_w5020_,
		_w5022_,
		_w5144_,
		_w6231_
	);
	LUT3 #(
		.INIT('h01)
	) name5699 (
		_w5047_,
		_w6231_,
		_w6230_,
		_w6232_
	);
	LUT4 #(
		.INIT('h0155)
	) name5700 (
		\sa30_reg[0]/P0002 ,
		_w6224_,
		_w6229_,
		_w6232_,
		_w6233_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name5701 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6234_
	);
	LUT2 #(
		.INIT('h2)
	) name5702 (
		_w5117_,
		_w6234_,
		_w6235_
	);
	LUT3 #(
		.INIT('h10)
	) name5703 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5158_,
		_w6236_
	);
	LUT2 #(
		.INIT('h8)
	) name5704 (
		_w5005_,
		_w5936_,
		_w6237_
	);
	LUT4 #(
		.INIT('h135f)
	) name5705 (
		_w5062_,
		_w5040_,
		_w5102_,
		_w5112_,
		_w6238_
	);
	LUT4 #(
		.INIT('h0100)
	) name5706 (
		_w6236_,
		_w6235_,
		_w6237_,
		_w6238_,
		_w6239_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name5707 (
		\sa30_reg[3]/P0001 ,
		_w5046_,
		_w5029_,
		_w5030_,
		_w6240_
	);
	LUT3 #(
		.INIT('h80)
	) name5708 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6241_
	);
	LUT2 #(
		.INIT('h8)
	) name5709 (
		_w5532_,
		_w6241_,
		_w6242_
	);
	LUT3 #(
		.INIT('h0d)
	) name5710 (
		\sa30_reg[2]/P0001 ,
		_w6240_,
		_w6242_,
		_w6243_
	);
	LUT4 #(
		.INIT('hedff)
	) name5711 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6244_
	);
	LUT4 #(
		.INIT('h7707)
	) name5712 (
		_w5011_,
		_w5100_,
		_w5112_,
		_w6244_,
		_w6245_
	);
	LUT4 #(
		.INIT('hd800)
	) name5713 (
		\sa30_reg[1]/P0001 ,
		_w6239_,
		_w6243_,
		_w6245_,
		_w6246_
	);
	LUT4 #(
		.INIT('h5655)
	) name5714 (
		\u0_w_reg[1][12]/P0001 ,
		_w6233_,
		_w6220_,
		_w6246_,
		_w6247_
	);
	LUT3 #(
		.INIT('h96)
	) name5715 (
		_w5580_,
		_w6012_,
		_w6247_,
		_w6248_
	);
	LUT4 #(
		.INIT('h9669)
	) name5716 (
		_w4691_,
		_w4804_,
		_w5758_,
		_w6195_,
		_w6249_
	);
	LUT3 #(
		.INIT('h82)
	) name5717 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[76]/P0001 ,
		\u0_w_reg[1][12]/P0001 ,
		_w6250_
	);
	LUT4 #(
		.INIT('h00eb)
	) name5718 (
		\ld_r_reg/P0001 ,
		_w6248_,
		_w6249_,
		_w6250_,
		_w6251_
	);
	LUT4 #(
		.INIT('h0001)
	) name5719 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6252_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name5720 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6253_
	);
	LUT3 #(
		.INIT('h8a)
	) name5721 (
		\sa12_reg[2]/P0001 ,
		_w6252_,
		_w6253_,
		_w6254_
	);
	LUT3 #(
		.INIT('h8a)
	) name5722 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6255_
	);
	LUT2 #(
		.INIT('h2)
	) name5723 (
		_w4592_,
		_w6255_,
		_w6256_
	);
	LUT4 #(
		.INIT('h0010)
	) name5724 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w6257_
	);
	LUT3 #(
		.INIT('h07)
	) name5725 (
		_w4588_,
		_w5202_,
		_w6257_,
		_w6258_
	);
	LUT4 #(
		.INIT('h5455)
	) name5726 (
		\sa12_reg[1]/P0001 ,
		_w6256_,
		_w6254_,
		_w6258_,
		_w6259_
	);
	LUT2 #(
		.INIT('h1)
	) name5727 (
		_w4630_,
		_w5205_,
		_w6260_
	);
	LUT3 #(
		.INIT('h2a)
	) name5728 (
		\sa12_reg[2]/P0001 ,
		_w4850_,
		_w6260_,
		_w6261_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name5729 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6262_
	);
	LUT4 #(
		.INIT('h0301)
	) name5730 (
		\sa12_reg[3]/P0001 ,
		_w4846_,
		_w4875_,
		_w6262_,
		_w6263_
	);
	LUT3 #(
		.INIT('h51)
	) name5731 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w6264_
	);
	LUT4 #(
		.INIT('h4041)
	) name5732 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6265_
	);
	LUT3 #(
		.INIT('ha8)
	) name5733 (
		\sa12_reg[1]/P0001 ,
		_w5230_,
		_w6265_,
		_w6266_
	);
	LUT3 #(
		.INIT('h0b)
	) name5734 (
		\sa12_reg[6]/NET0131 ,
		_w4679_,
		_w4646_,
		_w6267_
	);
	LUT4 #(
		.INIT('h3200)
	) name5735 (
		\sa12_reg[2]/P0001 ,
		_w6266_,
		_w6263_,
		_w6267_,
		_w6268_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5736 (
		\sa12_reg[0]/P0001 ,
		_w6261_,
		_w6259_,
		_w6268_,
		_w6269_
	);
	LUT4 #(
		.INIT('h8000)
	) name5737 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6270_
	);
	LUT3 #(
		.INIT('h01)
	) name5738 (
		_w5644_,
		_w5647_,
		_w6270_,
		_w6271_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5739 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6272_
	);
	LUT3 #(
		.INIT('h70)
	) name5740 (
		\sa12_reg[2]/P0001 ,
		_w4661_,
		_w6272_,
		_w6273_
	);
	LUT2 #(
		.INIT('h8)
	) name5741 (
		_w6271_,
		_w6273_,
		_w6274_
	);
	LUT2 #(
		.INIT('h1)
	) name5742 (
		\sa12_reg[3]/P0001 ,
		_w5663_,
		_w6275_
	);
	LUT3 #(
		.INIT('h2a)
	) name5743 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w6276_
	);
	LUT2 #(
		.INIT('h8)
	) name5744 (
		_w4601_,
		_w6276_,
		_w6277_
	);
	LUT3 #(
		.INIT('h02)
	) name5745 (
		_w4607_,
		_w6277_,
		_w6275_,
		_w6278_
	);
	LUT3 #(
		.INIT('hb9)
	) name5746 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6279_
	);
	LUT3 #(
		.INIT('ha2)
	) name5747 (
		\sa12_reg[2]/P0001 ,
		_w4592_,
		_w6279_,
		_w6280_
	);
	LUT2 #(
		.INIT('h1)
	) name5748 (
		\sa12_reg[2]/P0001 ,
		_w4624_,
		_w6281_
	);
	LUT3 #(
		.INIT('h13)
	) name5749 (
		_w6115_,
		_w6280_,
		_w6281_,
		_w6282_
	);
	LUT4 #(
		.INIT('h5501)
	) name5750 (
		\sa12_reg[0]/P0001 ,
		_w6274_,
		_w6278_,
		_w6282_,
		_w6283_
	);
	LUT4 #(
		.INIT('hff4b)
	) name5751 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6284_
	);
	LUT2 #(
		.INIT('h2)
	) name5752 (
		_w5202_,
		_w6284_,
		_w6285_
	);
	LUT4 #(
		.INIT('h0040)
	) name5753 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w6286_
	);
	LUT4 #(
		.INIT('h135f)
	) name5754 (
		_w4684_,
		_w4687_,
		_w4881_,
		_w6286_,
		_w6287_
	);
	LUT3 #(
		.INIT('h45)
	) name5755 (
		\sa12_reg[1]/P0001 ,
		_w6285_,
		_w6287_,
		_w6288_
	);
	LUT2 #(
		.INIT('h8)
	) name5756 (
		_w4642_,
		_w4822_,
		_w6289_
	);
	LUT3 #(
		.INIT('hd8)
	) name5757 (
		\sa12_reg[2]/P0001 ,
		_w4618_,
		_w5691_,
		_w6290_
	);
	LUT4 #(
		.INIT('hcdcf)
	) name5758 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[7]/NET0131 ,
		_w4624_,
		_w4593_,
		_w6291_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5759 (
		\sa12_reg[1]/P0001 ,
		_w6290_,
		_w6289_,
		_w6291_,
		_w6292_
	);
	LUT4 #(
		.INIT('hf800)
	) name5760 (
		_w4587_,
		_w4666_,
		_w4813_,
		_w5803_,
		_w6293_
	);
	LUT2 #(
		.INIT('h8)
	) name5761 (
		_w4635_,
		_w4633_,
		_w6294_
	);
	LUT4 #(
		.INIT('h3320)
	) name5762 (
		_w4635_,
		_w4642_,
		_w4633_,
		_w6270_,
		_w6295_
	);
	LUT2 #(
		.INIT('h1)
	) name5763 (
		_w6293_,
		_w6295_,
		_w6296_
	);
	LUT3 #(
		.INIT('h10)
	) name5764 (
		_w6292_,
		_w6288_,
		_w6296_,
		_w6297_
	);
	LUT3 #(
		.INIT('h10)
	) name5765 (
		_w6269_,
		_w6283_,
		_w6297_,
		_w6298_
	);
	LUT2 #(
		.INIT('h9)
	) name5766 (
		_w5695_,
		_w6298_,
		_w6299_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name5767 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6300_
	);
	LUT3 #(
		.INIT('h8a)
	) name5768 (
		\sa23_reg[2]/P0001 ,
		_w5306_,
		_w6300_,
		_w6301_
	);
	LUT3 #(
		.INIT('h40)
	) name5769 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w5711_,
		_w6302_
	);
	LUT3 #(
		.INIT('h8a)
	) name5770 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6303_
	);
	LUT3 #(
		.INIT('h31)
	) name5771 (
		_w4925_,
		_w5735_,
		_w6303_,
		_w6304_
	);
	LUT4 #(
		.INIT('h5455)
	) name5772 (
		\sa23_reg[1]/P0001 ,
		_w6302_,
		_w6301_,
		_w6304_,
		_w6305_
	);
	LUT4 #(
		.INIT('h8082)
	) name5773 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6306_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name5774 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6307_
	);
	LUT4 #(
		.INIT('h0301)
	) name5775 (
		\sa23_reg[3]/P0001 ,
		_w5713_,
		_w5731_,
		_w6307_,
		_w6308_
	);
	LUT3 #(
		.INIT('h45)
	) name5776 (
		\sa23_reg[2]/P0001 ,
		_w6306_,
		_w6308_,
		_w6309_
	);
	LUT2 #(
		.INIT('h1)
	) name5777 (
		_w5254_,
		_w5462_,
		_w6310_
	);
	LUT3 #(
		.INIT('h2a)
	) name5778 (
		\sa23_reg[2]/P0001 ,
		_w4958_,
		_w6310_,
		_w6311_
	);
	LUT2 #(
		.INIT('h8)
	) name5779 (
		\sa23_reg[1]/P0001 ,
		_w5278_,
		_w6312_
	);
	LUT3 #(
		.INIT('h07)
	) name5780 (
		_w4945_,
		_w5510_,
		_w5466_,
		_w6313_
	);
	LUT2 #(
		.INIT('h4)
	) name5781 (
		_w6312_,
		_w6313_,
		_w6314_
	);
	LUT4 #(
		.INIT('h0100)
	) name5782 (
		_w6309_,
		_w6311_,
		_w6305_,
		_w6314_,
		_w6315_
	);
	LUT2 #(
		.INIT('h2)
	) name5783 (
		\sa23_reg[0]/P0001 ,
		_w6315_,
		_w6316_
	);
	LUT4 #(
		.INIT('h9aff)
	) name5784 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w6317_
	);
	LUT4 #(
		.INIT('hbfaa)
	) name5785 (
		\sa23_reg[7]/NET0131 ,
		_w4889_,
		_w4900_,
		_w6317_,
		_w6318_
	);
	LUT3 #(
		.INIT('h67)
	) name5786 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6319_
	);
	LUT3 #(
		.INIT('h02)
	) name5787 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		_w6320_
	);
	LUT4 #(
		.INIT('h7077)
	) name5788 (
		_w4918_,
		_w4997_,
		_w6319_,
		_w6320_,
		_w6321_
	);
	LUT4 #(
		.INIT('h0155)
	) name5789 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[2]/P0001 ,
		_w6318_,
		_w6321_,
		_w6322_
	);
	LUT2 #(
		.INIT('h1)
	) name5790 (
		\sa23_reg[3]/P0001 ,
		_w5743_,
		_w6323_
	);
	LUT2 #(
		.INIT('h8)
	) name5791 (
		_w4918_,
		_w4948_,
		_w6324_
	);
	LUT4 #(
		.INIT('h0100)
	) name5792 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w6325_
	);
	LUT4 #(
		.INIT('h8000)
	) name5793 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6326_
	);
	LUT4 #(
		.INIT('h7ff8)
	) name5794 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6327_
	);
	LUT3 #(
		.INIT('h20)
	) name5795 (
		\sa23_reg[1]/P0001 ,
		_w6325_,
		_w6327_,
		_w6328_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name5796 (
		_w5493_,
		_w6323_,
		_w6324_,
		_w6328_,
		_w6329_
	);
	LUT4 #(
		.INIT('h0007)
	) name5797 (
		_w4890_,
		_w4937_,
		_w5292_,
		_w6176_,
		_w6330_
	);
	LUT3 #(
		.INIT('hb9)
	) name5798 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6331_
	);
	LUT4 #(
		.INIT('h4c00)
	) name5799 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6332_
	);
	LUT4 #(
		.INIT('h31f5)
	) name5800 (
		_w5714_,
		_w5747_,
		_w6331_,
		_w6332_,
		_w6333_
	);
	LUT3 #(
		.INIT('he0)
	) name5801 (
		\sa23_reg[2]/P0001 ,
		_w6330_,
		_w6333_,
		_w6334_
	);
	LUT3 #(
		.INIT('h45)
	) name5802 (
		\sa23_reg[0]/P0001 ,
		_w6329_,
		_w6334_,
		_w6335_
	);
	LUT3 #(
		.INIT('hd8)
	) name5803 (
		\sa23_reg[2]/P0001 ,
		_w4949_,
		_w4953_,
		_w6336_
	);
	LUT2 #(
		.INIT('h8)
	) name5804 (
		_w5295_,
		_w5278_,
		_w6337_
	);
	LUT4 #(
		.INIT('h135f)
	) name5805 (
		_w4901_,
		_w4907_,
		_w4919_,
		_w4971_,
		_w6338_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5806 (
		\sa23_reg[1]/P0001 ,
		_w6337_,
		_w6336_,
		_w6338_,
		_w6339_
	);
	LUT4 #(
		.INIT('h2a7f)
	) name5807 (
		\sa23_reg[2]/P0001 ,
		_w4896_,
		_w4901_,
		_w6326_,
		_w6340_
	);
	LUT2 #(
		.INIT('h4)
	) name5808 (
		_w6339_,
		_w6340_,
		_w6341_
	);
	LUT3 #(
		.INIT('h10)
	) name5809 (
		_w6335_,
		_w6322_,
		_w6341_,
		_w6342_
	);
	LUT3 #(
		.INIT('h65)
	) name5810 (
		_w5861_,
		_w6316_,
		_w6342_,
		_w6343_
	);
	LUT3 #(
		.INIT('ha8)
	) name5811 (
		\sa30_reg[2]/P0001 ,
		_w5165_,
		_w5982_,
		_w6344_
	);
	LUT4 #(
		.INIT('h0800)
	) name5812 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w6345_
	);
	LUT4 #(
		.INIT('h5554)
	) name5813 (
		\sa30_reg[2]/P0001 ,
		_w5050_,
		_w5913_,
		_w6345_,
		_w6346_
	);
	LUT4 #(
		.INIT('h0002)
	) name5814 (
		\sa30_reg[1]/P0001 ,
		_w5065_,
		_w5019_,
		_w5037_,
		_w6347_
	);
	LUT3 #(
		.INIT('h10)
	) name5815 (
		_w6346_,
		_w6344_,
		_w6347_,
		_w6348_
	);
	LUT4 #(
		.INIT('h5540)
	) name5816 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w5132_,
		_w5171_,
		_w6349_
	);
	LUT3 #(
		.INIT('h15)
	) name5817 (
		\sa30_reg[1]/P0001 ,
		_w5011_,
		_w5100_,
		_w6350_
	);
	LUT4 #(
		.INIT('h0020)
	) name5818 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6351_
	);
	LUT2 #(
		.INIT('h8)
	) name5819 (
		\sa30_reg[5]/P0001 ,
		_w6351_,
		_w6352_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name5820 (
		\sa30_reg[5]/P0001 ,
		_w5039_,
		_w5036_,
		_w5112_,
		_w6353_
	);
	LUT4 #(
		.INIT('h1000)
	) name5821 (
		_w6352_,
		_w6349_,
		_w6350_,
		_w6353_,
		_w6354_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5822 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w6355_
	);
	LUT2 #(
		.INIT('h4)
	) name5823 (
		_w5179_,
		_w6355_,
		_w6356_
	);
	LUT4 #(
		.INIT('h1333)
	) name5824 (
		\sa30_reg[4]/P0001 ,
		_w5098_,
		_w5112_,
		_w5113_,
		_w6357_
	);
	LUT4 #(
		.INIT('hf400)
	) name5825 (
		_w5032_,
		_w5570_,
		_w6356_,
		_w6357_,
		_w6358_
	);
	LUT4 #(
		.INIT('h0155)
	) name5826 (
		\sa30_reg[0]/P0002 ,
		_w6348_,
		_w6354_,
		_w6358_,
		_w6359_
	);
	LUT3 #(
		.INIT('h13)
	) name5827 (
		\sa30_reg[7]/P0001 ,
		_w5084_,
		_w5095_,
		_w6360_
	);
	LUT4 #(
		.INIT('hcedf)
	) name5828 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6361_
	);
	LUT3 #(
		.INIT('h8a)
	) name5829 (
		\sa30_reg[2]/P0001 ,
		_w6241_,
		_w6361_,
		_w6362_
	);
	LUT3 #(
		.INIT('ha2)
	) name5830 (
		\sa30_reg[1]/P0001 ,
		_w6360_,
		_w6362_,
		_w6363_
	);
	LUT2 #(
		.INIT('h8)
	) name5831 (
		_w5062_,
		_w5067_,
		_w6364_
	);
	LUT4 #(
		.INIT('h0301)
	) name5832 (
		_w5026_,
		_w5046_,
		_w5025_,
		_w5525_,
		_w6365_
	);
	LUT3 #(
		.INIT('h45)
	) name5833 (
		\sa30_reg[1]/P0001 ,
		_w6364_,
		_w6365_,
		_w6366_
	);
	LUT4 #(
		.INIT('h5504)
	) name5834 (
		\sa30_reg[3]/P0001 ,
		_w5040_,
		_w5532_,
		_w5990_,
		_w6367_
	);
	LUT4 #(
		.INIT('h0001)
	) name5835 (
		_w5046_,
		_w5929_,
		_w5990_,
		_w5979_,
		_w6368_
	);
	LUT3 #(
		.INIT('h32)
	) name5836 (
		\sa30_reg[2]/P0001 ,
		_w6367_,
		_w6368_,
		_w6369_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5837 (
		\sa30_reg[0]/P0002 ,
		_w6363_,
		_w6366_,
		_w6369_,
		_w6370_
	);
	LUT4 #(
		.INIT('h0007)
	) name5838 (
		_w5029_,
		_w5030_,
		_w5135_,
		_w5578_,
		_w6371_
	);
	LUT4 #(
		.INIT('hedff)
	) name5839 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w5011_,
		_w6372_
	);
	LUT4 #(
		.INIT('h0155)
	) name5840 (
		\sa30_reg[1]/P0001 ,
		\sa30_reg[2]/P0001 ,
		_w6371_,
		_w6372_,
		_w6373_
	);
	LUT3 #(
		.INIT('h01)
	) name5841 (
		_w5065_,
		_w5140_,
		_w5556_,
		_w6374_
	);
	LUT2 #(
		.INIT('h1)
	) name5842 (
		_w5090_,
		_w5128_,
		_w6375_
	);
	LUT3 #(
		.INIT('h2a)
	) name5843 (
		_w5049_,
		_w6374_,
		_w6375_,
		_w6376_
	);
	LUT4 #(
		.INIT('h0007)
	) name5844 (
		_w5020_,
		_w5022_,
		_w5098_,
		_w5914_,
		_w6377_
	);
	LUT4 #(
		.INIT('hc0e0)
	) name5845 (
		_w5040_,
		_w5095_,
		_w5184_,
		_w5573_,
		_w6378_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name5846 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6379_
	);
	LUT2 #(
		.INIT('h2)
	) name5847 (
		_w5112_,
		_w6379_,
		_w6380_
	);
	LUT4 #(
		.INIT('h0301)
	) name5848 (
		_w5934_,
		_w6378_,
		_w6380_,
		_w6377_,
		_w6381_
	);
	LUT3 #(
		.INIT('h10)
	) name5849 (
		_w6376_,
		_w6373_,
		_w6381_,
		_w6382_
	);
	LUT3 #(
		.INIT('h10)
	) name5850 (
		_w6370_,
		_w6359_,
		_w6382_,
		_w6383_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name5851 (
		\u0_w_reg[1][17]/P0001 ,
		_w6370_,
		_w6359_,
		_w6382_,
		_w6384_
	);
	LUT3 #(
		.INIT('h69)
	) name5852 (
		_w5758_,
		_w6053_,
		_w6384_,
		_w6385_
	);
	LUT4 #(
		.INIT('h4114)
	) name5853 (
		\ld_r_reg/P0001 ,
		_w6299_,
		_w6343_,
		_w6385_,
		_w6386_
	);
	LUT3 #(
		.INIT('h28)
	) name5854 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[81]/P0001 ,
		\u0_w_reg[1][17]/P0001 ,
		_w6387_
	);
	LUT2 #(
		.INIT('he)
	) name5855 (
		_w6386_,
		_w6387_,
		_w6388_
	);
	LUT4 #(
		.INIT('hffda)
	) name5856 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6389_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5857 (
		\sa12_reg[1]/P0001 ,
		\sa12_reg[2]/P0001 ,
		_w5238_,
		_w6389_,
		_w6390_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name5858 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6391_
	);
	LUT4 #(
		.INIT('h3f1d)
	) name5859 (
		\sa12_reg[1]/P0001 ,
		_w4591_,
		_w4593_,
		_w6391_,
		_w6392_
	);
	LUT3 #(
		.INIT('h54)
	) name5860 (
		\sa12_reg[1]/P0001 ,
		_w5691_,
		_w6286_,
		_w6393_
	);
	LUT4 #(
		.INIT('hcc80)
	) name5861 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4621_,
		_w4631_,
		_w6394_
	);
	LUT4 #(
		.INIT('h0302)
	) name5862 (
		\sa12_reg[2]/P0001 ,
		_w6393_,
		_w6394_,
		_w6392_,
		_w6395_
	);
	LUT3 #(
		.INIT('h45)
	) name5863 (
		\sa12_reg[0]/P0001 ,
		_w6390_,
		_w6395_,
		_w6396_
	);
	LUT2 #(
		.INIT('h8)
	) name5864 (
		_w5769_,
		_w6264_,
		_w6397_
	);
	LUT4 #(
		.INIT('h020a)
	) name5865 (
		\sa12_reg[1]/P0001 ,
		_w4687_,
		_w5675_,
		_w6286_,
		_w6398_
	);
	LUT2 #(
		.INIT('h4)
	) name5866 (
		_w6397_,
		_w6398_,
		_w6399_
	);
	LUT2 #(
		.INIT('h8)
	) name5867 (
		_w4611_,
		_w5644_,
		_w6400_
	);
	LUT3 #(
		.INIT('h23)
	) name5868 (
		\sa12_reg[2]/P0001 ,
		_w4634_,
		_w4863_,
		_w6401_
	);
	LUT4 #(
		.INIT('h0020)
	) name5869 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6402_
	);
	LUT4 #(
		.INIT('h0001)
	) name5870 (
		\sa12_reg[1]/P0001 ,
		_w4598_,
		_w6257_,
		_w6402_,
		_w6403_
	);
	LUT2 #(
		.INIT('h1)
	) name5871 (
		_w4663_,
		_w4610_,
		_w6404_
	);
	LUT4 #(
		.INIT('h4000)
	) name5872 (
		_w6400_,
		_w6403_,
		_w6404_,
		_w6401_,
		_w6405_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name5873 (
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6406_
	);
	LUT2 #(
		.INIT('h2)
	) name5874 (
		_w4684_,
		_w6406_,
		_w6407_
	);
	LUT4 #(
		.INIT('h153f)
	) name5875 (
		_w4654_,
		_w4587_,
		_w4666_,
		_w4623_,
		_w6408_
	);
	LUT3 #(
		.INIT('h10)
	) name5876 (
		_w6294_,
		_w6407_,
		_w6408_,
		_w6409_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5877 (
		\sa12_reg[0]/P0001 ,
		_w6399_,
		_w6405_,
		_w6409_,
		_w6410_
	);
	LUT4 #(
		.INIT('h0007)
	) name5878 (
		\sa12_reg[4]/P0001 ,
		_w4661_,
		_w5234_,
		_w5666_,
		_w6411_
	);
	LUT4 #(
		.INIT('haaa2)
	) name5879 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w6412_
	);
	LUT4 #(
		.INIT('h0700)
	) name5880 (
		\sa12_reg[7]/NET0131 ,
		_w4668_,
		_w5691_,
		_w6412_,
		_w6413_
	);
	LUT4 #(
		.INIT('h000b)
	) name5881 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[4]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		_w6414_
	);
	LUT3 #(
		.INIT('h45)
	) name5882 (
		\sa12_reg[1]/P0001 ,
		_w4878_,
		_w6414_,
		_w6415_
	);
	LUT4 #(
		.INIT('hf800)
	) name5883 (
		_w5196_,
		_w6411_,
		_w6413_,
		_w6415_,
		_w6416_
	);
	LUT4 #(
		.INIT('haadf)
	) name5884 (
		\sa12_reg[3]/P0001 ,
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6417_
	);
	LUT4 #(
		.INIT('h0a08)
	) name5885 (
		\sa12_reg[2]/P0001 ,
		\sa12_reg[4]/P0001 ,
		_w4863_,
		_w6417_,
		_w6418_
	);
	LUT2 #(
		.INIT('h1)
	) name5886 (
		\sa12_reg[2]/P0001 ,
		_w4830_,
		_w6419_
	);
	LUT2 #(
		.INIT('h2)
	) name5887 (
		\sa12_reg[1]/P0001 ,
		_w4670_,
		_w6420_
	);
	LUT4 #(
		.INIT('hec00)
	) name5888 (
		_w5781_,
		_w6418_,
		_w6419_,
		_w6420_,
		_w6421_
	);
	LUT3 #(
		.INIT('had)
	) name5889 (
		\sa12_reg[5]/P0001 ,
		\sa12_reg[6]/NET0131 ,
		\sa12_reg[7]/NET0131 ,
		_w6422_
	);
	LUT2 #(
		.INIT('h2)
	) name5890 (
		_w4860_,
		_w6422_,
		_w6423_
	);
	LUT2 #(
		.INIT('h1)
	) name5891 (
		_w6137_,
		_w6423_,
		_w6424_
	);
	LUT3 #(
		.INIT('he0)
	) name5892 (
		_w6416_,
		_w6421_,
		_w6424_,
		_w6425_
	);
	LUT3 #(
		.INIT('h10)
	) name5893 (
		_w6410_,
		_w6396_,
		_w6425_,
		_w6426_
	);
	LUT4 #(
		.INIT('h0001)
	) name5894 (
		\sa01_reg[1]/P0001 ,
		_w4735_,
		_w4739_,
		_w5867_,
		_w6427_
	);
	LUT3 #(
		.INIT('h0e)
	) name5895 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		_w6428_
	);
	LUT2 #(
		.INIT('h2)
	) name5896 (
		_w4782_,
		_w6428_,
		_w6429_
	);
	LUT3 #(
		.INIT('h08)
	) name5897 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w6430_
	);
	LUT4 #(
		.INIT('h7077)
	) name5898 (
		_w4723_,
		_w4725_,
		_w4767_,
		_w6430_,
		_w6431_
	);
	LUT3 #(
		.INIT('h40)
	) name5899 (
		_w6429_,
		_w6427_,
		_w6431_,
		_w6432_
	);
	LUT3 #(
		.INIT('h53)
	) name5900 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w6433_
	);
	LUT4 #(
		.INIT('h0222)
	) name5901 (
		\sa01_reg[1]/P0001 ,
		_w5362_,
		_w5359_,
		_w6433_,
		_w6434_
	);
	LUT2 #(
		.INIT('h4)
	) name5902 (
		_w5899_,
		_w6434_,
		_w6435_
	);
	LUT4 #(
		.INIT('h5554)
	) name5903 (
		\sa01_reg[3]/P0001 ,
		_w4703_,
		_w4695_,
		_w4722_,
		_w6436_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name5904 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w6437_
	);
	LUT2 #(
		.INIT('h2)
	) name5905 (
		_w4775_,
		_w6437_,
		_w6438_
	);
	LUT2 #(
		.INIT('h1)
	) name5906 (
		_w6436_,
		_w6438_,
		_w6439_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5907 (
		\sa01_reg[0]/P0001 ,
		_w6432_,
		_w6435_,
		_w6439_,
		_w6440_
	);
	LUT4 #(
		.INIT('h0007)
	) name5908 (
		_w4704_,
		_w4749_,
		_w5352_,
		_w5366_,
		_w6441_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name5909 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[2]/P0001 ,
		_w4790_,
		_w6441_,
		_w6442_
	);
	LUT3 #(
		.INIT('he0)
	) name5910 (
		_w4764_,
		_w5374_,
		_w5442_,
		_w6443_
	);
	LUT3 #(
		.INIT('had)
	) name5911 (
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w6444_
	);
	LUT2 #(
		.INIT('h2)
	) name5912 (
		_w5896_,
		_w6444_,
		_w6445_
	);
	LUT3 #(
		.INIT('h80)
	) name5913 (
		\sa01_reg[1]/P0001 ,
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		_w6446_
	);
	LUT2 #(
		.INIT('h8)
	) name5914 (
		_w4802_,
		_w6446_,
		_w6447_
	);
	LUT4 #(
		.INIT('h0001)
	) name5915 (
		_w6090_,
		_w6443_,
		_w6447_,
		_w6445_,
		_w6448_
	);
	LUT2 #(
		.INIT('h4)
	) name5916 (
		_w6442_,
		_w6448_,
		_w6449_
	);
	LUT4 #(
		.INIT('hbcfc)
	) name5917 (
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w6450_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5918 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		_w5638_,
		_w6450_,
		_w6451_
	);
	LUT4 #(
		.INIT('h0013)
	) name5919 (
		\sa01_reg[6]/NET0131 ,
		_w4722_,
		_w4796_,
		_w5438_,
		_w6452_
	);
	LUT4 #(
		.INIT('h000b)
	) name5920 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		_w6453_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name5921 (
		_w4741_,
		_w4759_,
		_w5337_,
		_w6453_,
		_w6454_
	);
	LUT4 #(
		.INIT('h3200)
	) name5922 (
		\sa01_reg[2]/P0001 ,
		_w6451_,
		_w6452_,
		_w6454_,
		_w6455_
	);
	LUT2 #(
		.INIT('h1)
	) name5923 (
		\sa01_reg[1]/P0001 ,
		_w6455_,
		_w6456_
	);
	LUT4 #(
		.INIT('hffda)
	) name5924 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w6457_
	);
	LUT2 #(
		.INIT('h2)
	) name5925 (
		\sa01_reg[2]/P0001 ,
		_w6457_,
		_w6458_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name5926 (
		\sa01_reg[3]/P0001 ,
		\sa01_reg[4]/P0001 ,
		\sa01_reg[6]/NET0131 ,
		\sa01_reg[7]/NET0131 ,
		_w6459_
	);
	LUT3 #(
		.INIT('h51)
	) name5927 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w6460_
	);
	LUT3 #(
		.INIT('h45)
	) name5928 (
		_w5432_,
		_w6459_,
		_w6460_,
		_w6461_
	);
	LUT3 #(
		.INIT('h8a)
	) name5929 (
		\sa01_reg[1]/P0001 ,
		_w6458_,
		_w6461_,
		_w6462_
	);
	LUT4 #(
		.INIT('h1333)
	) name5930 (
		\sa01_reg[2]/P0001 ,
		_w4743_,
		_w4757_,
		_w4776_,
		_w6463_
	);
	LUT4 #(
		.INIT('h0040)
	) name5931 (
		\sa01_reg[2]/P0001 ,
		\sa01_reg[3]/P0001 ,
		\sa01_reg[5]/P0001 ,
		\sa01_reg[7]/NET0131 ,
		_w6464_
	);
	LUT3 #(
		.INIT('h54)
	) name5932 (
		\sa01_reg[1]/P0001 ,
		_w5638_,
		_w6464_,
		_w6465_
	);
	LUT3 #(
		.INIT('h40)
	) name5933 (
		\sa01_reg[2]/P0001 ,
		_w4692_,
		_w4732_,
		_w6466_
	);
	LUT3 #(
		.INIT('h10)
	) name5934 (
		_w6465_,
		_w6466_,
		_w6463_,
		_w6467_
	);
	LUT3 #(
		.INIT('h45)
	) name5935 (
		\sa01_reg[0]/P0001 ,
		_w6462_,
		_w6467_,
		_w6468_
	);
	LUT4 #(
		.INIT('h0100)
	) name5936 (
		_w6440_,
		_w6456_,
		_w6468_,
		_w6449_,
		_w6469_
	);
	LUT3 #(
		.INIT('h69)
	) name5937 (
		_w5861_,
		_w6426_,
		_w6469_,
		_w6470_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name5938 (
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6471_
	);
	LUT4 #(
		.INIT('h20a8)
	) name5939 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		_w4948_,
		_w6471_,
		_w6472_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5940 (
		\sa23_reg[2]/P0001 ,
		_w4967_,
		_w4994_,
		_w5460_,
		_w6473_
	);
	LUT4 #(
		.INIT('h0001)
	) name5941 (
		_w5490_,
		_w5497_,
		_w5508_,
		_w5735_,
		_w6474_
	);
	LUT4 #(
		.INIT('h5455)
	) name5942 (
		\sa23_reg[1]/P0001 ,
		_w5258_,
		_w6473_,
		_w6474_,
		_w6475_
	);
	LUT4 #(
		.INIT('h4555)
	) name5943 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w6476_
	);
	LUT4 #(
		.INIT('h0700)
	) name5944 (
		_w4925_,
		_w4948_,
		_w5289_,
		_w6476_,
		_w6477_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5945 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6478_
	);
	LUT2 #(
		.INIT('h2)
	) name5946 (
		\sa23_reg[1]/P0001 ,
		_w6478_,
		_w6479_
	);
	LUT4 #(
		.INIT('hcedf)
	) name5947 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w4901_,
		_w4981_,
		_w6480_
	);
	LUT3 #(
		.INIT('hb0)
	) name5948 (
		_w6477_,
		_w6479_,
		_w6480_,
		_w6481_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5949 (
		\sa23_reg[0]/P0001 ,
		_w6475_,
		_w6472_,
		_w6481_,
		_w6482_
	);
	LUT3 #(
		.INIT('h01)
	) name5950 (
		_w5258_,
		_w5282_,
		_w5469_,
		_w6483_
	);
	LUT3 #(
		.INIT('h02)
	) name5951 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w6484_
	);
	LUT3 #(
		.INIT('h07)
	) name5952 (
		\sa23_reg[6]/NET0131 ,
		_w5254_,
		_w6484_,
		_w6485_
	);
	LUT4 #(
		.INIT('h135f)
	) name5953 (
		_w5483_,
		_w5752_,
		_w6483_,
		_w6485_,
		_w6486_
	);
	LUT4 #(
		.INIT('h000b)
	) name5954 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		_w6487_
	);
	LUT2 #(
		.INIT('h4)
	) name5955 (
		_w4929_,
		_w6487_,
		_w6488_
	);
	LUT3 #(
		.INIT('h54)
	) name5956 (
		\sa23_reg[1]/P0001 ,
		_w6486_,
		_w6488_,
		_w6489_
	);
	LUT3 #(
		.INIT('had)
	) name5957 (
		\sa23_reg[5]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6490_
	);
	LUT2 #(
		.INIT('h2)
	) name5958 (
		_w4900_,
		_w6490_,
		_w6491_
	);
	LUT4 #(
		.INIT('h0007)
	) name5959 (
		_w4887_,
		_w4908_,
		_w4967_,
		_w4981_,
		_w6492_
	);
	LUT4 #(
		.INIT('hc0c8)
	) name5960 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[2]/P0001 ,
		_w6491_,
		_w6492_,
		_w6493_
	);
	LUT2 #(
		.INIT('h1)
	) name5961 (
		_w6186_,
		_w6493_,
		_w6494_
	);
	LUT4 #(
		.INIT('hffda)
	) name5962 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6495_
	);
	LUT2 #(
		.INIT('h2)
	) name5963 (
		\sa23_reg[2]/P0001 ,
		_w6495_,
		_w6496_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name5964 (
		\sa23_reg[3]/P0001 ,
		\sa23_reg[4]/P0001 ,
		\sa23_reg[6]/NET0131 ,
		\sa23_reg[7]/NET0131 ,
		_w6497_
	);
	LUT3 #(
		.INIT('h51)
	) name5965 (
		\sa23_reg[2]/P0001 ,
		\sa23_reg[5]/P0001 ,
		\sa23_reg[7]/NET0131 ,
		_w6498_
	);
	LUT3 #(
		.INIT('h45)
	) name5966 (
		_w5279_,
		_w6497_,
		_w6498_,
		_w6499_
	);
	LUT3 #(
		.INIT('h8a)
	) name5967 (
		\sa23_reg[1]/P0001 ,
		_w6496_,
		_w6499_,
		_w6500_
	);
	LUT4 #(
		.INIT('h0051)
	) name5968 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[2]/P0001 ,
		_w4953_,
		_w4954_,
		_w6501_
	);
	LUT3 #(
		.INIT('h13)
	) name5969 (
		_w4918_,
		_w4938_,
		_w4967_,
		_w6502_
	);
	LUT3 #(
		.INIT('h10)
	) name5970 (
		_w5310_,
		_w6501_,
		_w6502_,
		_w6503_
	);
	LUT4 #(
		.INIT('h0103)
	) name5971 (
		_w4896_,
		_w4915_,
		_w4933_,
		_w5259_,
		_w6504_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name5972 (
		\sa23_reg[1]/P0001 ,
		\sa23_reg[2]/P0001 ,
		_w4906_,
		_w6504_,
		_w6505_
	);
	LUT4 #(
		.INIT('h00ba)
	) name5973 (
		\sa23_reg[0]/P0001 ,
		_w6500_,
		_w6503_,
		_w6505_,
		_w6506_
	);
	LUT4 #(
		.INIT('h1000)
	) name5974 (
		_w6482_,
		_w6489_,
		_w6494_,
		_w6506_,
		_w6507_
	);
	LUT3 #(
		.INIT('h69)
	) name5975 (
		\u0_w_reg[1][2]/P0001 ,
		_w6383_,
		_w6507_,
		_w6508_
	);
	LUT3 #(
		.INIT('h28)
	) name5976 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[66]/P0001 ,
		\u0_w_reg[1][2]/P0001 ,
		_w6509_
	);
	LUT4 #(
		.INIT('hff41)
	) name5977 (
		\ld_r_reg/P0001 ,
		_w6470_,
		_w6508_,
		_w6509_,
		_w6510_
	);
	LUT4 #(
		.INIT('h5655)
	) name5978 (
		\u0_w_reg[1][25]/P0001 ,
		_w6370_,
		_w6359_,
		_w6382_,
		_w6511_
	);
	LUT3 #(
		.INIT('h69)
	) name5979 (
		_w5811_,
		_w6053_,
		_w6511_,
		_w6512_
	);
	LUT4 #(
		.INIT('h4114)
	) name5980 (
		\ld_r_reg/P0001 ,
		_w5910_,
		_w6299_,
		_w6512_,
		_w6513_
	);
	LUT3 #(
		.INIT('h28)
	) name5981 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[89]/P0001 ,
		\u0_w_reg[1][25]/P0001 ,
		_w6514_
	);
	LUT2 #(
		.INIT('he)
	) name5982 (
		_w6513_,
		_w6514_,
		_w6515_
	);
	LUT4 #(
		.INIT('h659a)
	) name5983 (
		_w5316_,
		_w5599_,
		_w5642_,
		_w5695_,
		_w6516_
	);
	LUT3 #(
		.INIT('h69)
	) name5984 (
		\u0_w_reg[1][15]/P0001 ,
		_w5194_,
		_w6012_,
		_w6517_
	);
	LUT3 #(
		.INIT('h82)
	) name5985 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[79]/P0001 ,
		\u0_w_reg[1][15]/P0001 ,
		_w6518_
	);
	LUT4 #(
		.INIT('h00be)
	) name5986 (
		\ld_r_reg/P0001 ,
		_w6516_,
		_w6517_,
		_w6518_,
		_w6519_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name5987 (
		\u0_w_reg[1][27]/P0001 ,
		_w6233_,
		_w6220_,
		_w6246_,
		_w6520_
	);
	LUT3 #(
		.INIT('h69)
	) name5988 (
		_w6147_,
		_w6195_,
		_w6520_,
		_w6521_
	);
	LUT3 #(
		.INIT('h4b)
	) name5989 (
		_w5599_,
		_w5642_,
		_w6469_,
		_w6522_
	);
	LUT2 #(
		.INIT('h9)
	) name5990 (
		_w5695_,
		_w6426_,
		_w6523_
	);
	LUT4 #(
		.INIT('h1441)
	) name5991 (
		\ld_r_reg/P0001 ,
		_w6521_,
		_w6522_,
		_w6523_,
		_w6524_
	);
	LUT3 #(
		.INIT('h82)
	) name5992 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[91]/P0001 ,
		\u0_w_reg[1][27]/P0001 ,
		_w6525_
	);
	LUT2 #(
		.INIT('h1)
	) name5993 (
		_w6524_,
		_w6525_,
		_w6526_
	);
	LUT4 #(
		.INIT('h5655)
	) name5994 (
		\u0_w_reg[1][19]/P0001 ,
		_w6233_,
		_w6220_,
		_w6246_,
		_w6527_
	);
	LUT3 #(
		.INIT('h69)
	) name5995 (
		_w5758_,
		_w6195_,
		_w6527_,
		_w6528_
	);
	LUT4 #(
		.INIT('h6996)
	) name5996 (
		_w5695_,
		_w6102_,
		_w6426_,
		_w6507_,
		_w6529_
	);
	LUT3 #(
		.INIT('h82)
	) name5997 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[83]/P0001 ,
		\u0_w_reg[1][19]/P0001 ,
		_w6530_
	);
	LUT4 #(
		.INIT('h00eb)
	) name5998 (
		\ld_r_reg/P0001 ,
		_w6528_,
		_w6529_,
		_w6530_,
		_w6531_
	);
	LUT2 #(
		.INIT('h9)
	) name5999 (
		_w6102_,
		_w6147_,
		_w6532_
	);
	LUT4 #(
		.INIT('h6996)
	) name6000 (
		_w5758_,
		_w6102_,
		_w6147_,
		_w6507_,
		_w6533_
	);
	LUT4 #(
		.INIT('h0002)
	) name6001 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6534_
	);
	LUT4 #(
		.INIT('h008a)
	) name6002 (
		\sa30_reg[1]/P0001 ,
		_w5018_,
		_w5965_,
		_w6534_,
		_w6535_
	);
	LUT2 #(
		.INIT('h4)
	) name6003 (
		_w5953_,
		_w6535_,
		_w6536_
	);
	LUT3 #(
		.INIT('h07)
	) name6004 (
		_w5040_,
		_w5041_,
		_w5128_,
		_w6537_
	);
	LUT3 #(
		.INIT('h13)
	) name6005 (
		_w5076_,
		_w5545_,
		_w5532_,
		_w6538_
	);
	LUT3 #(
		.INIT('h01)
	) name6006 (
		_w5526_,
		_w5917_,
		_w6351_,
		_w6539_
	);
	LUT4 #(
		.INIT('h8000)
	) name6007 (
		_w5530_,
		_w6539_,
		_w6537_,
		_w6538_,
		_w6540_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name6008 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6541_
	);
	LUT2 #(
		.INIT('h2)
	) name6009 (
		_w5112_,
		_w6541_,
		_w6542_
	);
	LUT3 #(
		.INIT('h8a)
	) name6010 (
		\sa30_reg[0]/P0002 ,
		\sa30_reg[7]/P0001 ,
		_w5556_,
		_w6543_
	);
	LUT4 #(
		.INIT('h153f)
	) name6011 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5154_,
		_w6351_,
		_w6544_
	);
	LUT3 #(
		.INIT('h40)
	) name6012 (
		_w6542_,
		_w6543_,
		_w6544_,
		_w6545_
	);
	LUT3 #(
		.INIT('he0)
	) name6013 (
		_w6536_,
		_w6540_,
		_w6545_,
		_w6546_
	);
	LUT4 #(
		.INIT('h0040)
	) name6014 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w6547_
	);
	LUT3 #(
		.INIT('h01)
	) name6015 (
		\sa30_reg[1]/P0001 ,
		_w5031_,
		_w6547_,
		_w6548_
	);
	LUT4 #(
		.INIT('haaa8)
	) name6016 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6549_
	);
	LUT4 #(
		.INIT('ha020)
	) name6017 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6550_
	);
	LUT4 #(
		.INIT('h5554)
	) name6018 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w6551_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name6019 (
		_w5037_,
		_w6549_,
		_w6550_,
		_w6551_,
		_w6552_
	);
	LUT2 #(
		.INIT('h2)
	) name6020 (
		\sa30_reg[1]/P0001 ,
		_w5979_,
		_w6553_
	);
	LUT3 #(
		.INIT('h45)
	) name6021 (
		_w6548_,
		_w6552_,
		_w6553_,
		_w6554_
	);
	LUT4 #(
		.INIT('h0105)
	) name6022 (
		\sa30_reg[0]/P0002 ,
		_w5102_,
		_w5129_,
		_w5538_,
		_w6555_
	);
	LUT2 #(
		.INIT('h4)
	) name6023 (
		_w5116_,
		_w6555_,
		_w6556_
	);
	LUT2 #(
		.INIT('h4)
	) name6024 (
		_w6554_,
		_w6556_,
		_w6557_
	);
	LUT4 #(
		.INIT('hbcfc)
	) name6025 (
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6558_
	);
	LUT4 #(
		.INIT('h0a02)
	) name6026 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		_w5031_,
		_w6558_,
		_w6559_
	);
	LUT4 #(
		.INIT('h0045)
	) name6027 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w5095_,
		_w5173_,
		_w6560_
	);
	LUT2 #(
		.INIT('h1)
	) name6028 (
		_w5128_,
		_w5995_,
		_w6561_
	);
	LUT4 #(
		.INIT('h0008)
	) name6029 (
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		_w6562_
	);
	LUT3 #(
		.INIT('h01)
	) name6030 (
		\sa30_reg[1]/P0001 ,
		_w5542_,
		_w6562_,
		_w6563_
	);
	LUT4 #(
		.INIT('hea00)
	) name6031 (
		_w6559_,
		_w6560_,
		_w6561_,
		_w6563_,
		_w6564_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6032 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		\sa30_reg[7]/P0001 ,
		_w6565_
	);
	LUT4 #(
		.INIT('h1300)
	) name6033 (
		_w5014_,
		_w5094_,
		_w5106_,
		_w6565_,
		_w6566_
	);
	LUT2 #(
		.INIT('h2)
	) name6034 (
		\sa30_reg[1]/P0001 ,
		_w5069_,
		_w6567_
	);
	LUT4 #(
		.INIT('hf800)
	) name6035 (
		_w5078_,
		_w6360_,
		_w6566_,
		_w6567_,
		_w6568_
	);
	LUT3 #(
		.INIT('had)
	) name6036 (
		\sa30_reg[5]/P0001 ,
		\sa30_reg[6]/NET0131 ,
		\sa30_reg[7]/P0001 ,
		_w6569_
	);
	LUT3 #(
		.INIT('h02)
	) name6037 (
		\sa30_reg[2]/P0001 ,
		\sa30_reg[3]/P0001 ,
		\sa30_reg[4]/P0001 ,
		_w6570_
	);
	LUT2 #(
		.INIT('h4)
	) name6038 (
		_w6569_,
		_w6570_,
		_w6571_
	);
	LUT2 #(
		.INIT('h1)
	) name6039 (
		_w6236_,
		_w6571_,
		_w6572_
	);
	LUT3 #(
		.INIT('he0)
	) name6040 (
		_w6564_,
		_w6568_,
		_w6572_,
		_w6573_
	);
	LUT3 #(
		.INIT('he0)
	) name6041 (
		_w6546_,
		_w6557_,
		_w6573_,
		_w6574_
	);
	LUT4 #(
		.INIT('h5655)
	) name6042 (
		\u0_w_reg[1][11]/P0001 ,
		_w6233_,
		_w6220_,
		_w6246_,
		_w6575_
	);
	LUT3 #(
		.INIT('h69)
	) name6043 (
		_w6012_,
		_w6574_,
		_w6575_,
		_w6576_
	);
	LUT3 #(
		.INIT('h82)
	) name6044 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[75]/P0001 ,
		\u0_w_reg[1][11]/P0001 ,
		_w6577_
	);
	LUT4 #(
		.INIT('h00eb)
	) name6045 (
		\ld_r_reg/P0001 ,
		_w6533_,
		_w6576_,
		_w6577_,
		_w6578_
	);
	LUT4 #(
		.INIT('h5655)
	) name6046 (
		\u0_w_reg[1][4]/P0001 ,
		_w6233_,
		_w6220_,
		_w6246_,
		_w6579_
	);
	LUT3 #(
		.INIT('h96)
	) name6047 (
		_w5517_,
		_w6012_,
		_w6579_,
		_w6580_
	);
	LUT4 #(
		.INIT('h1441)
	) name6048 (
		\ld_r_reg/P0001 ,
		_w4805_,
		_w6103_,
		_w6580_,
		_w6581_
	);
	LUT3 #(
		.INIT('h82)
	) name6049 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[68]/P0001 ,
		\u0_w_reg[1][4]/P0001 ,
		_w6582_
	);
	LUT2 #(
		.INIT('h1)
	) name6050 (
		_w6581_,
		_w6582_,
		_w6583_
	);
	LUT4 #(
		.INIT('h56aa)
	) name6051 (
		\u0_w_reg[1][26]/P0001 ,
		_w6546_,
		_w6557_,
		_w6573_,
		_w6584_
	);
	LUT3 #(
		.INIT('h69)
	) name6052 (
		_w6426_,
		_w6507_,
		_w6584_,
		_w6585_
	);
	LUT3 #(
		.INIT('h28)
	) name6053 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[90]/P0001 ,
		\u0_w_reg[1][26]/P0001 ,
		_w6586_
	);
	LUT4 #(
		.INIT('hff14)
	) name6054 (
		\ld_r_reg/P0001 ,
		_w5862_,
		_w6585_,
		_w6586_,
		_w6587_
	);
	LUT2 #(
		.INIT('h9)
	) name6055 (
		\u0_w_reg[1][31]/P0001 ,
		_w6012_,
		_w6588_
	);
	LUT4 #(
		.INIT('h6996)
	) name6056 (
		_w5248_,
		_w5454_,
		_w5695_,
		_w5758_,
		_w6589_
	);
	LUT3 #(
		.INIT('h82)
	) name6057 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[95]/P0001 ,
		\u0_w_reg[1][31]/P0001 ,
		_w6590_
	);
	LUT4 #(
		.INIT('h00be)
	) name6058 (
		\ld_r_reg/P0001 ,
		_w6588_,
		_w6589_,
		_w6590_,
		_w6591_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name6059 (
		\u0_w_reg[1][16]/P0001 ,
		_w5932_,
		_w5947_,
		_w5960_,
		_w6592_
	);
	LUT3 #(
		.INIT('h65)
	) name6060 (
		_w5758_,
		_w6316_,
		_w6342_,
		_w6593_
	);
	LUT2 #(
		.INIT('h9)
	) name6061 (
		_w5695_,
		_w5909_,
		_w6594_
	);
	LUT4 #(
		.INIT('h1441)
	) name6062 (
		\ld_r_reg/P0001 ,
		_w6592_,
		_w6593_,
		_w6594_,
		_w6595_
	);
	LUT3 #(
		.INIT('h28)
	) name6063 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[80]/P0001 ,
		\u0_w_reg[1][16]/P0001 ,
		_w6596_
	);
	LUT2 #(
		.INIT('he)
	) name6064 (
		_w6595_,
		_w6596_,
		_w6597_
	);
	LUT3 #(
		.INIT('h69)
	) name6065 (
		_w5811_,
		_w6053_,
		_w6469_,
		_w6598_
	);
	LUT4 #(
		.INIT('ha955)
	) name6066 (
		\u0_w_reg[1][18]/P0001 ,
		_w6546_,
		_w6557_,
		_w6573_,
		_w6599_
	);
	LUT2 #(
		.INIT('h6)
	) name6067 (
		_w6507_,
		_w6599_,
		_w6600_
	);
	LUT3 #(
		.INIT('h82)
	) name6068 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[82]/P0001 ,
		\u0_w_reg[1][18]/P0001 ,
		_w6601_
	);
	LUT4 #(
		.INIT('h00eb)
	) name6069 (
		\ld_r_reg/P0001 ,
		_w6598_,
		_w6600_,
		_w6601_,
		_w6602_
	);
	LUT4 #(
		.INIT('h9699)
	) name6070 (
		_w5248_,
		_w5316_,
		_w5599_,
		_w5642_,
		_w6603_
	);
	LUT3 #(
		.INIT('h69)
	) name6071 (
		\u0_w_reg[1][23]/P0001 ,
		_w5758_,
		_w6012_,
		_w6604_
	);
	LUT3 #(
		.INIT('h82)
	) name6072 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[87]/P0001 ,
		\u0_w_reg[1][23]/P0001 ,
		_w6605_
	);
	LUT4 #(
		.INIT('h00eb)
	) name6073 (
		\ld_r_reg/P0001 ,
		_w6603_,
		_w6604_,
		_w6605_,
		_w6606_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name6074 (
		\u0_w_reg[1][24]/P0002 ,
		_w5932_,
		_w5947_,
		_w5960_,
		_w6607_
	);
	LUT3 #(
		.INIT('h65)
	) name6075 (
		_w6298_,
		_w6316_,
		_w6342_,
		_w6608_
	);
	LUT4 #(
		.INIT('h4114)
	) name6076 (
		\ld_r_reg/P0001 ,
		_w5696_,
		_w6607_,
		_w6608_,
		_w6609_
	);
	LUT3 #(
		.INIT('h28)
	) name6077 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[88]/P0001 ,
		\u0_w_reg[1][24]/P0002 ,
		_w6610_
	);
	LUT2 #(
		.INIT('he)
	) name6078 (
		_w6609_,
		_w6610_,
		_w6611_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name6079 (
		\u0_w_reg[1][8]/P0001 ,
		_w5932_,
		_w5947_,
		_w5960_,
		_w6612_
	);
	LUT4 #(
		.INIT('h6996)
	) name6080 (
		_w5758_,
		_w5909_,
		_w6012_,
		_w6298_,
		_w6613_
	);
	LUT3 #(
		.INIT('h82)
	) name6081 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[72]/P0001 ,
		\u0_w_reg[1][8]/P0001 ,
		_w6614_
	);
	LUT4 #(
		.INIT('h00eb)
	) name6082 (
		\ld_r_reg/P0001 ,
		_w6612_,
		_w6613_,
		_w6614_,
		_w6615_
	);
	LUT3 #(
		.INIT('h69)
	) name6083 (
		_w6053_,
		_w6426_,
		_w6469_,
		_w6616_
	);
	LUT4 #(
		.INIT('ha955)
	) name6084 (
		\u0_w_reg[1][10]/P0001 ,
		_w6546_,
		_w6557_,
		_w6573_,
		_w6617_
	);
	LUT2 #(
		.INIT('h6)
	) name6085 (
		_w6383_,
		_w6617_,
		_w6618_
	);
	LUT3 #(
		.INIT('h82)
	) name6086 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[74]/P0001 ,
		\u0_w_reg[1][10]/P0001 ,
		_w6619_
	);
	LUT4 #(
		.INIT('h00eb)
	) name6087 (
		\ld_r_reg/P0001 ,
		_w6616_,
		_w6618_,
		_w6619_,
		_w6620_
	);
	LUT4 #(
		.INIT('h5655)
	) name6088 (
		\u0_w_reg[1][3]/P0001 ,
		_w6181_,
		_w6164_,
		_w6194_,
		_w6621_
	);
	LUT3 #(
		.INIT('h69)
	) name6089 (
		_w6012_,
		_w6574_,
		_w6621_,
		_w6622_
	);
	LUT4 #(
		.INIT('h4114)
	) name6090 (
		\ld_r_reg/P0001 ,
		_w6522_,
		_w6532_,
		_w6622_,
		_w6623_
	);
	LUT3 #(
		.INIT('h82)
	) name6091 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[67]/P0001 ,
		\u0_w_reg[1][3]/P0001 ,
		_w6624_
	);
	LUT2 #(
		.INIT('h1)
	) name6092 (
		_w6623_,
		_w6624_,
		_w6625_
	);
	LUT2 #(
		.INIT('h9)
	) name6093 (
		\u0_w_reg[1][5]/P0001 ,
		_w5121_,
		_w6626_
	);
	LUT4 #(
		.INIT('h5655)
	) name6094 (
		\u0_w_reg[1][6]/P0001 ,
		_w5148_,
		_w5170_,
		_w5193_,
		_w6627_
	);
	LUT2 #(
		.INIT('h9)
	) name6095 (
		\u0_w_reg[1][4]/P0001 ,
		_w5580_,
		_w6628_
	);
	LUT4 #(
		.INIT('h5655)
	) name6096 (
		\u0_w_reg[1][0]/P0001 ,
		_w5932_,
		_w5947_,
		_w5960_,
		_w6629_
	);
	LUT4 #(
		.INIT('h5655)
	) name6097 (
		\u0_w_reg[1][3]/P0001 ,
		_w6233_,
		_w6220_,
		_w6246_,
		_w6630_
	);
	LUT4 #(
		.INIT('h5655)
	) name6098 (
		\u0_w_reg[1][1]/P0001 ,
		_w6370_,
		_w6359_,
		_w6382_,
		_w6631_
	);
	LUT4 #(
		.INIT('ha955)
	) name6099 (
		\u0_w_reg[1][2]/P0001 ,
		_w6546_,
		_w6557_,
		_w6573_,
		_w6632_
	);
	LUT2 #(
		.INIT('h9)
	) name6100 (
		\u0_w_reg[1][7]/P0001 ,
		_w6012_,
		_w6633_
	);
	LUT2 #(
		.INIT('h2)
	) name6101 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w6634_
	);
	LUT2 #(
		.INIT('h2)
	) name6102 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6635_
	);
	LUT3 #(
		.INIT('h20)
	) name6103 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6636_
	);
	LUT2 #(
		.INIT('h4)
	) name6104 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6637_
	);
	LUT4 #(
		.INIT('h0100)
	) name6105 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6638_
	);
	LUT4 #(
		.INIT('h5510)
	) name6106 (
		\sa11_reg[2]/P0001 ,
		_w6634_,
		_w6636_,
		_w6638_,
		_w6639_
	);
	LUT2 #(
		.INIT('h2)
	) name6107 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w6640_
	);
	LUT3 #(
		.INIT('h20)
	) name6108 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6641_
	);
	LUT3 #(
		.INIT('h08)
	) name6109 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6642_
	);
	LUT4 #(
		.INIT('h0080)
	) name6110 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6643_
	);
	LUT2 #(
		.INIT('h8)
	) name6111 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w6644_
	);
	LUT4 #(
		.INIT('h0080)
	) name6112 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6645_
	);
	LUT4 #(
		.INIT('h0111)
	) name6113 (
		_w6643_,
		_w6645_,
		_w6640_,
		_w6641_,
		_w6646_
	);
	LUT3 #(
		.INIT('h8a)
	) name6114 (
		\sa11_reg[1]/P0001 ,
		_w6639_,
		_w6646_,
		_w6647_
	);
	LUT4 #(
		.INIT('h0040)
	) name6115 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6648_
	);
	LUT2 #(
		.INIT('h4)
	) name6116 (
		\sa11_reg[2]/P0001 ,
		_w6648_,
		_w6649_
	);
	LUT2 #(
		.INIT('h8)
	) name6117 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6650_
	);
	LUT2 #(
		.INIT('h8)
	) name6118 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w6651_
	);
	LUT4 #(
		.INIT('h8000)
	) name6119 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6652_
	);
	LUT4 #(
		.INIT('h0002)
	) name6120 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6653_
	);
	LUT2 #(
		.INIT('h2)
	) name6121 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6654_
	);
	LUT4 #(
		.INIT('h0002)
	) name6122 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6655_
	);
	LUT3 #(
		.INIT('h01)
	) name6123 (
		_w6653_,
		_w6655_,
		_w6652_,
		_w6656_
	);
	LUT3 #(
		.INIT('h45)
	) name6124 (
		\sa11_reg[1]/P0001 ,
		_w6649_,
		_w6656_,
		_w6657_
	);
	LUT3 #(
		.INIT('h02)
	) name6125 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6658_
	);
	LUT4 #(
		.INIT('h0008)
	) name6126 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6659_
	);
	LUT3 #(
		.INIT('h10)
	) name6127 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6660_
	);
	LUT4 #(
		.INIT('h0100)
	) name6128 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6661_
	);
	LUT4 #(
		.INIT('haa20)
	) name6129 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6659_,
		_w6661_,
		_w6662_
	);
	LUT2 #(
		.INIT('h8)
	) name6130 (
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6663_
	);
	LUT3 #(
		.INIT('h40)
	) name6131 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6664_
	);
	LUT2 #(
		.INIT('h4)
	) name6132 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w6665_
	);
	LUT2 #(
		.INIT('h2)
	) name6133 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6666_
	);
	LUT4 #(
		.INIT('h0004)
	) name6134 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6667_
	);
	LUT4 #(
		.INIT('h5540)
	) name6135 (
		\sa11_reg[3]/P0001 ,
		_w6664_,
		_w6665_,
		_w6667_,
		_w6668_
	);
	LUT2 #(
		.INIT('h1)
	) name6136 (
		_w6662_,
		_w6668_,
		_w6669_
	);
	LUT4 #(
		.INIT('h5455)
	) name6137 (
		\sa11_reg[0]/P0001 ,
		_w6647_,
		_w6657_,
		_w6669_,
		_w6670_
	);
	LUT2 #(
		.INIT('h8)
	) name6138 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6671_
	);
	LUT4 #(
		.INIT('h0080)
	) name6139 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6672_
	);
	LUT4 #(
		.INIT('h008a)
	) name6140 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w6638_,
		_w6672_,
		_w6673_
	);
	LUT2 #(
		.INIT('h1)
	) name6141 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6674_
	);
	LUT3 #(
		.INIT('h80)
	) name6142 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6675_
	);
	LUT3 #(
		.INIT('h02)
	) name6143 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6676_
	);
	LUT4 #(
		.INIT('h0004)
	) name6144 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6677_
	);
	LUT4 #(
		.INIT('h0020)
	) name6145 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6678_
	);
	LUT4 #(
		.INIT('h0103)
	) name6146 (
		_w6674_,
		_w6677_,
		_w6678_,
		_w6675_,
		_w6679_
	);
	LUT4 #(
		.INIT('h1000)
	) name6147 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6680_
	);
	LUT3 #(
		.INIT('h80)
	) name6148 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6681_
	);
	LUT2 #(
		.INIT('h4)
	) name6149 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w6682_
	);
	LUT4 #(
		.INIT('h0400)
	) name6150 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6683_
	);
	LUT4 #(
		.INIT('h0015)
	) name6151 (
		\sa11_reg[2]/P0001 ,
		_w6634_,
		_w6681_,
		_w6683_,
		_w6684_
	);
	LUT4 #(
		.INIT('h7077)
	) name6152 (
		_w6673_,
		_w6679_,
		_w6680_,
		_w6684_,
		_w6685_
	);
	LUT2 #(
		.INIT('h1)
	) name6153 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w6686_
	);
	LUT4 #(
		.INIT('h0010)
	) name6154 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6687_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name6155 (
		\sa11_reg[6]/NET0131 ,
		_w6642_,
		_w6644_,
		_w6687_,
		_w6688_
	);
	LUT3 #(
		.INIT('h45)
	) name6156 (
		\sa11_reg[1]/P0001 ,
		_w6685_,
		_w6688_,
		_w6689_
	);
	LUT2 #(
		.INIT('h4)
	) name6157 (
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6690_
	);
	LUT3 #(
		.INIT('h10)
	) name6158 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6691_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name6159 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6692_
	);
	LUT2 #(
		.INIT('h1)
	) name6160 (
		\sa11_reg[2]/P0001 ,
		_w6692_,
		_w6693_
	);
	LUT3 #(
		.INIT('h02)
	) name6161 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6694_
	);
	LUT2 #(
		.INIT('h8)
	) name6162 (
		_w6666_,
		_w6694_,
		_w6695_
	);
	LUT3 #(
		.INIT('h04)
	) name6163 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6696_
	);
	LUT2 #(
		.INIT('h4)
	) name6164 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6697_
	);
	LUT4 #(
		.INIT('h0200)
	) name6165 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6698_
	);
	LUT4 #(
		.INIT('h002a)
	) name6166 (
		\sa11_reg[1]/P0001 ,
		_w6674_,
		_w6696_,
		_w6698_,
		_w6699_
	);
	LUT3 #(
		.INIT('h10)
	) name6167 (
		_w6695_,
		_w6693_,
		_w6699_,
		_w6700_
	);
	LUT3 #(
		.INIT('h08)
	) name6168 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6701_
	);
	LUT4 #(
		.INIT('h0008)
	) name6169 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6702_
	);
	LUT2 #(
		.INIT('h4)
	) name6170 (
		\sa11_reg[2]/P0001 ,
		_w6702_,
		_w6703_
	);
	LUT4 #(
		.INIT('h0800)
	) name6171 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6704_
	);
	LUT2 #(
		.INIT('h8)
	) name6172 (
		\sa11_reg[2]/P0001 ,
		_w6704_,
		_w6705_
	);
	LUT2 #(
		.INIT('h8)
	) name6173 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6706_
	);
	LUT2 #(
		.INIT('h1)
	) name6174 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w6707_
	);
	LUT3 #(
		.INIT('h32)
	) name6175 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w6708_
	);
	LUT4 #(
		.INIT('h2000)
	) name6176 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6709_
	);
	LUT4 #(
		.INIT('h0051)
	) name6177 (
		\sa11_reg[1]/P0001 ,
		_w6706_,
		_w6708_,
		_w6709_,
		_w6710_
	);
	LUT3 #(
		.INIT('h10)
	) name6178 (
		_w6705_,
		_w6703_,
		_w6710_,
		_w6711_
	);
	LUT2 #(
		.INIT('h4)
	) name6179 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6712_
	);
	LUT4 #(
		.INIT('h4000)
	) name6180 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6713_
	);
	LUT4 #(
		.INIT('h0200)
	) name6181 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6714_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name6182 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6715_
	);
	LUT4 #(
		.INIT('h0200)
	) name6183 (
		\sa11_reg[2]/P0001 ,
		_w6713_,
		_w6714_,
		_w6715_,
		_w6716_
	);
	LUT4 #(
		.INIT('h2000)
	) name6184 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6717_
	);
	LUT2 #(
		.INIT('h1)
	) name6185 (
		\sa11_reg[2]/P0001 ,
		_w6717_,
		_w6718_
	);
	LUT4 #(
		.INIT('h0001)
	) name6186 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6719_
	);
	LUT2 #(
		.INIT('h4)
	) name6187 (
		\sa11_reg[5]/P0001 ,
		_w6719_,
		_w6720_
	);
	LUT4 #(
		.INIT('h0020)
	) name6188 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6721_
	);
	LUT3 #(
		.INIT('h0b)
	) name6189 (
		\sa11_reg[5]/P0001 ,
		_w6719_,
		_w6721_,
		_w6722_
	);
	LUT3 #(
		.INIT('h15)
	) name6190 (
		_w6716_,
		_w6718_,
		_w6722_,
		_w6723_
	);
	LUT4 #(
		.INIT('haa02)
	) name6191 (
		\sa11_reg[0]/P0001 ,
		_w6700_,
		_w6711_,
		_w6723_,
		_w6724_
	);
	LUT3 #(
		.INIT('h10)
	) name6192 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6725_
	);
	LUT4 #(
		.INIT('h2220)
	) name6193 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6726_
	);
	LUT3 #(
		.INIT('h07)
	) name6194 (
		_w6650_,
		_w6725_,
		_w6726_,
		_w6727_
	);
	LUT4 #(
		.INIT('h153f)
	) name6195 (
		_w6634_,
		_w6641_,
		_w6671_,
		_w6691_,
		_w6728_
	);
	LUT4 #(
		.INIT('hba00)
	) name6196 (
		\sa11_reg[2]/P0001 ,
		_w6720_,
		_w6727_,
		_w6728_,
		_w6729_
	);
	LUT2 #(
		.INIT('h8)
	) name6197 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w6730_
	);
	LUT4 #(
		.INIT('h0020)
	) name6198 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6731_
	);
	LUT4 #(
		.INIT('h153f)
	) name6199 (
		\sa11_reg[4]/P0001 ,
		_w6730_,
		_w6676_,
		_w6731_,
		_w6732_
	);
	LUT4 #(
		.INIT('h0010)
	) name6200 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6733_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name6201 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w6652_,
		_w6733_,
		_w6734_
	);
	LUT3 #(
		.INIT('h0d)
	) name6202 (
		\sa11_reg[1]/P0001 ,
		_w6732_,
		_w6734_,
		_w6735_
	);
	LUT3 #(
		.INIT('hd0)
	) name6203 (
		\sa11_reg[1]/P0001 ,
		_w6729_,
		_w6735_,
		_w6736_
	);
	LUT4 #(
		.INIT('h0100)
	) name6204 (
		_w6670_,
		_w6724_,
		_w6689_,
		_w6736_,
		_w6737_
	);
	LUT2 #(
		.INIT('h2)
	) name6205 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w6738_
	);
	LUT2 #(
		.INIT('h4)
	) name6206 (
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6739_
	);
	LUT3 #(
		.INIT('h20)
	) name6207 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6740_
	);
	LUT3 #(
		.INIT('h10)
	) name6208 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w6741_
	);
	LUT4 #(
		.INIT('h0100)
	) name6209 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6742_
	);
	LUT4 #(
		.INIT('h5510)
	) name6210 (
		\sa00_reg[2]/P0001 ,
		_w6738_,
		_w6740_,
		_w6742_,
		_w6743_
	);
	LUT2 #(
		.INIT('h4)
	) name6211 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w6744_
	);
	LUT2 #(
		.INIT('h4)
	) name6212 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w6745_
	);
	LUT3 #(
		.INIT('h20)
	) name6213 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w6746_
	);
	LUT2 #(
		.INIT('h2)
	) name6214 (
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6747_
	);
	LUT2 #(
		.INIT('h8)
	) name6215 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w6748_
	);
	LUT4 #(
		.INIT('h0080)
	) name6216 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6749_
	);
	LUT2 #(
		.INIT('h8)
	) name6217 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w6750_
	);
	LUT4 #(
		.INIT('h0080)
	) name6218 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6751_
	);
	LUT4 #(
		.INIT('h0111)
	) name6219 (
		_w6749_,
		_w6751_,
		_w6744_,
		_w6746_,
		_w6752_
	);
	LUT3 #(
		.INIT('h8a)
	) name6220 (
		\sa00_reg[1]/P0001 ,
		_w6743_,
		_w6752_,
		_w6753_
	);
	LUT3 #(
		.INIT('h02)
	) name6221 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w6754_
	);
	LUT3 #(
		.INIT('h40)
	) name6222 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w6755_
	);
	LUT4 #(
		.INIT('h1000)
	) name6223 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w6756_
	);
	LUT3 #(
		.INIT('h54)
	) name6224 (
		\sa00_reg[7]/NET0131 ,
		_w6754_,
		_w6756_,
		_w6757_
	);
	LUT2 #(
		.INIT('h1)
	) name6225 (
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6758_
	);
	LUT3 #(
		.INIT('h01)
	) name6226 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6759_
	);
	LUT4 #(
		.INIT('h7f7c)
	) name6227 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6760_
	);
	LUT2 #(
		.INIT('h2)
	) name6228 (
		\sa00_reg[2]/P0001 ,
		_w6760_,
		_w6761_
	);
	LUT3 #(
		.INIT('h54)
	) name6229 (
		\sa00_reg[1]/P0001 ,
		_w6757_,
		_w6761_,
		_w6762_
	);
	LUT2 #(
		.INIT('h2)
	) name6230 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w6763_
	);
	LUT3 #(
		.INIT('h02)
	) name6231 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6764_
	);
	LUT2 #(
		.INIT('h4)
	) name6232 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w6765_
	);
	LUT3 #(
		.INIT('h10)
	) name6233 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w6766_
	);
	LUT4 #(
		.INIT('h0100)
	) name6234 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w6767_
	);
	LUT4 #(
		.INIT('haa80)
	) name6235 (
		\sa00_reg[2]/P0001 ,
		_w6763_,
		_w6764_,
		_w6767_,
		_w6768_
	);
	LUT2 #(
		.INIT('h4)
	) name6236 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w6769_
	);
	LUT3 #(
		.INIT('h01)
	) name6237 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6770_
	);
	LUT4 #(
		.INIT('h1000)
	) name6238 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6771_
	);
	LUT2 #(
		.INIT('h4)
	) name6239 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w6772_
	);
	LUT4 #(
		.INIT('h0777)
	) name6240 (
		_w6769_,
		_w6770_,
		_w6771_,
		_w6772_,
		_w6773_
	);
	LUT2 #(
		.INIT('h4)
	) name6241 (
		_w6768_,
		_w6773_,
		_w6774_
	);
	LUT4 #(
		.INIT('h5455)
	) name6242 (
		\sa00_reg[0]/P0001 ,
		_w6762_,
		_w6753_,
		_w6774_,
		_w6775_
	);
	LUT2 #(
		.INIT('h2)
	) name6243 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w6776_
	);
	LUT4 #(
		.INIT('h0080)
	) name6244 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6777_
	);
	LUT4 #(
		.INIT('h0020)
	) name6245 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w6778_
	);
	LUT3 #(
		.INIT('h02)
	) name6246 (
		\sa00_reg[2]/P0001 ,
		_w6778_,
		_w6777_,
		_w6779_
	);
	LUT2 #(
		.INIT('h8)
	) name6247 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w6780_
	);
	LUT3 #(
		.INIT('h02)
	) name6248 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w6781_
	);
	LUT2 #(
		.INIT('h8)
	) name6249 (
		_w6780_,
		_w6781_,
		_w6782_
	);
	LUT4 #(
		.INIT('h0100)
	) name6250 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w6783_
	);
	LUT3 #(
		.INIT('h02)
	) name6251 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6784_
	);
	LUT4 #(
		.INIT('h0004)
	) name6252 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6785_
	);
	LUT3 #(
		.INIT('h0b)
	) name6253 (
		\sa00_reg[6]/NET0131 ,
		_w6783_,
		_w6785_,
		_w6786_
	);
	LUT3 #(
		.INIT('h40)
	) name6254 (
		_w6782_,
		_w6779_,
		_w6786_,
		_w6787_
	);
	LUT3 #(
		.INIT('h80)
	) name6255 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6788_
	);
	LUT2 #(
		.INIT('h8)
	) name6256 (
		_w6738_,
		_w6788_,
		_w6789_
	);
	LUT4 #(
		.INIT('h0400)
	) name6257 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w6790_
	);
	LUT3 #(
		.INIT('h01)
	) name6258 (
		\sa00_reg[2]/P0001 ,
		_w6771_,
		_w6790_,
		_w6791_
	);
	LUT2 #(
		.INIT('h4)
	) name6259 (
		_w6789_,
		_w6791_,
		_w6792_
	);
	LUT4 #(
		.INIT('h33bf)
	) name6260 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w6770_,
		_w6749_,
		_w6793_
	);
	LUT4 #(
		.INIT('h0155)
	) name6261 (
		\sa00_reg[1]/P0001 ,
		_w6787_,
		_w6792_,
		_w6793_,
		_w6794_
	);
	LUT4 #(
		.INIT('h0200)
	) name6262 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6795_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name6263 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6796_
	);
	LUT2 #(
		.INIT('h1)
	) name6264 (
		\sa00_reg[2]/P0001 ,
		_w6796_,
		_w6797_
	);
	LUT2 #(
		.INIT('h8)
	) name6265 (
		_w6738_,
		_w6784_,
		_w6798_
	);
	LUT4 #(
		.INIT('h0200)
	) name6266 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6799_
	);
	LUT4 #(
		.INIT('h0222)
	) name6267 (
		\sa00_reg[1]/P0001 ,
		_w6799_,
		_w6745_,
		_w6759_,
		_w6800_
	);
	LUT3 #(
		.INIT('h10)
	) name6268 (
		_w6797_,
		_w6798_,
		_w6800_,
		_w6801_
	);
	LUT4 #(
		.INIT('h0800)
	) name6269 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6802_
	);
	LUT2 #(
		.INIT('h8)
	) name6270 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w6803_
	);
	LUT3 #(
		.INIT('h80)
	) name6271 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w6804_
	);
	LUT2 #(
		.INIT('h4)
	) name6272 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w6805_
	);
	LUT4 #(
		.INIT('h1000)
	) name6273 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w6806_
	);
	LUT4 #(
		.INIT('h0013)
	) name6274 (
		\sa00_reg[2]/P0001 ,
		_w6804_,
		_w6802_,
		_w6806_,
		_w6807_
	);
	LUT4 #(
		.INIT('h2000)
	) name6275 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6808_
	);
	LUT4 #(
		.INIT('h0008)
	) name6276 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6809_
	);
	LUT4 #(
		.INIT('h0405)
	) name6277 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[2]/P0001 ,
		_w6808_,
		_w6809_,
		_w6810_
	);
	LUT2 #(
		.INIT('h8)
	) name6278 (
		_w6807_,
		_w6810_,
		_w6811_
	);
	LUT3 #(
		.INIT('h32)
	) name6279 (
		_w6745_,
		_w6780_,
		_w6788_,
		_w6812_
	);
	LUT4 #(
		.INIT('h0200)
	) name6280 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6813_
	);
	LUT3 #(
		.INIT('h02)
	) name6281 (
		\sa00_reg[2]/P0001 ,
		_w6813_,
		_w6754_,
		_w6814_
	);
	LUT2 #(
		.INIT('h1)
	) name6282 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w6815_
	);
	LUT2 #(
		.INIT('h8)
	) name6283 (
		_w6759_,
		_w6815_,
		_w6816_
	);
	LUT4 #(
		.INIT('h2000)
	) name6284 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6817_
	);
	LUT2 #(
		.INIT('h1)
	) name6285 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w6818_
	);
	LUT4 #(
		.INIT('h0020)
	) name6286 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6819_
	);
	LUT3 #(
		.INIT('h01)
	) name6287 (
		\sa00_reg[2]/P0001 ,
		_w6817_,
		_w6819_,
		_w6820_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name6288 (
		_w6812_,
		_w6814_,
		_w6816_,
		_w6820_,
		_w6821_
	);
	LUT4 #(
		.INIT('haa02)
	) name6289 (
		\sa00_reg[0]/P0001 ,
		_w6801_,
		_w6811_,
		_w6821_,
		_w6822_
	);
	LUT4 #(
		.INIT('h1000)
	) name6290 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6823_
	);
	LUT2 #(
		.INIT('h8)
	) name6291 (
		\sa00_reg[5]/P0001 ,
		_w6823_,
		_w6824_
	);
	LUT4 #(
		.INIT('h2220)
	) name6292 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6825_
	);
	LUT3 #(
		.INIT('h07)
	) name6293 (
		_w6759_,
		_w6815_,
		_w6825_,
		_w6826_
	);
	LUT3 #(
		.INIT('h45)
	) name6294 (
		\sa00_reg[2]/P0001 ,
		_w6824_,
		_w6826_,
		_w6827_
	);
	LUT3 #(
		.INIT('h80)
	) name6295 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w6828_
	);
	LUT4 #(
		.INIT('h0200)
	) name6296 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w6829_
	);
	LUT4 #(
		.INIT('h8cbf)
	) name6297 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w6828_,
		_w6829_,
		_w6830_
	);
	LUT2 #(
		.INIT('h8)
	) name6298 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		_w6831_
	);
	LUT2 #(
		.INIT('h2)
	) name6299 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		_w6832_
	);
	LUT3 #(
		.INIT('h08)
	) name6300 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6833_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name6301 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		_w6784_,
		_w6833_,
		_w6834_
	);
	LUT2 #(
		.INIT('h8)
	) name6302 (
		_w6830_,
		_w6834_,
		_w6835_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6303 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w6836_
	);
	LUT2 #(
		.INIT('h1)
	) name6304 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w6837_
	);
	LUT2 #(
		.INIT('h4)
	) name6305 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w6838_
	);
	LUT4 #(
		.INIT('h0010)
	) name6306 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6839_
	);
	LUT4 #(
		.INIT('h00c8)
	) name6307 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		_w6839_,
		_w6836_,
		_w6840_
	);
	LUT4 #(
		.INIT('h0075)
	) name6308 (
		\sa00_reg[1]/P0001 ,
		_w6827_,
		_w6835_,
		_w6840_,
		_w6841_
	);
	LUT4 #(
		.INIT('h0100)
	) name6309 (
		_w6822_,
		_w6794_,
		_w6775_,
		_w6841_,
		_w6842_
	);
	LUT2 #(
		.INIT('h9)
	) name6310 (
		_w6737_,
		_w6842_,
		_w6843_
	);
	LUT3 #(
		.INIT('ha8)
	) name6311 (
		\sa11_reg[2]/P0001 ,
		_w6660_,
		_w6702_,
		_w6844_
	);
	LUT2 #(
		.INIT('h4)
	) name6312 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w6845_
	);
	LUT2 #(
		.INIT('h8)
	) name6313 (
		_w6691_,
		_w6845_,
		_w6846_
	);
	LUT2 #(
		.INIT('h8)
	) name6314 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6847_
	);
	LUT4 #(
		.INIT('h8000)
	) name6315 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6848_
	);
	LUT4 #(
		.INIT('h0c2f)
	) name6316 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w6642_,
		_w6848_,
		_w6849_
	);
	LUT4 #(
		.INIT('h5455)
	) name6317 (
		\sa11_reg[1]/P0001 ,
		_w6844_,
		_w6846_,
		_w6849_,
		_w6850_
	);
	LUT3 #(
		.INIT('h01)
	) name6318 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6851_
	);
	LUT4 #(
		.INIT('hdfd3)
	) name6319 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6852_
	);
	LUT3 #(
		.INIT('h8a)
	) name6320 (
		\sa11_reg[1]/P0001 ,
		_w6851_,
		_w6852_,
		_w6853_
	);
	LUT3 #(
		.INIT('h04)
	) name6321 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6854_
	);
	LUT3 #(
		.INIT('h01)
	) name6322 (
		_w6721_,
		_w6672_,
		_w6854_,
		_w6855_
	);
	LUT3 #(
		.INIT('h45)
	) name6323 (
		\sa11_reg[2]/P0001 ,
		_w6853_,
		_w6855_,
		_w6856_
	);
	LUT4 #(
		.INIT('h37bf)
	) name6324 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w6636_,
		_w6676_,
		_w6857_
	);
	LUT4 #(
		.INIT('h0200)
	) name6325 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6858_
	);
	LUT3 #(
		.INIT('h07)
	) name6326 (
		_w6674_,
		_w6696_,
		_w6858_,
		_w6859_
	);
	LUT3 #(
		.INIT('h2a)
	) name6327 (
		\sa11_reg[1]/P0001 ,
		_w6857_,
		_w6859_,
		_w6860_
	);
	LUT3 #(
		.INIT('h04)
	) name6328 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6861_
	);
	LUT2 #(
		.INIT('h8)
	) name6329 (
		_w6686_,
		_w6861_,
		_w6862_
	);
	LUT4 #(
		.INIT('haeaf)
	) name6330 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w6848_,
		_w6861_,
		_w6863_
	);
	LUT4 #(
		.INIT('h0777)
	) name6331 (
		_w6642_,
		_w6634_,
		_w6664_,
		_w6665_,
		_w6864_
	);
	LUT3 #(
		.INIT('hd0)
	) name6332 (
		\sa11_reg[2]/P0001 ,
		_w6863_,
		_w6864_,
		_w6865_
	);
	LUT4 #(
		.INIT('h0100)
	) name6333 (
		_w6856_,
		_w6860_,
		_w6850_,
		_w6865_,
		_w6866_
	);
	LUT2 #(
		.INIT('h2)
	) name6334 (
		\sa11_reg[0]/P0001 ,
		_w6866_,
		_w6867_
	);
	LUT4 #(
		.INIT('h0002)
	) name6335 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6868_
	);
	LUT4 #(
		.INIT('heffd)
	) name6336 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6869_
	);
	LUT4 #(
		.INIT('h1000)
	) name6337 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6870_
	);
	LUT2 #(
		.INIT('h4)
	) name6338 (
		\sa11_reg[7]/NET0131 ,
		_w6870_,
		_w6871_
	);
	LUT4 #(
		.INIT('h0400)
	) name6339 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6872_
	);
	LUT3 #(
		.INIT('h8b)
	) name6340 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6873_
	);
	LUT3 #(
		.INIT('h13)
	) name6341 (
		_w6706_,
		_w6872_,
		_w6873_,
		_w6874_
	);
	LUT3 #(
		.INIT('h40)
	) name6342 (
		_w6871_,
		_w6869_,
		_w6874_,
		_w6875_
	);
	LUT4 #(
		.INIT('h0040)
	) name6343 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6876_
	);
	LUT4 #(
		.INIT('h0010)
	) name6344 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6877_
	);
	LUT3 #(
		.INIT('h54)
	) name6345 (
		\sa11_reg[2]/P0001 ,
		_w6876_,
		_w6877_,
		_w6878_
	);
	LUT3 #(
		.INIT('h80)
	) name6346 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6879_
	);
	LUT4 #(
		.INIT('h0080)
	) name6347 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6880_
	);
	LUT3 #(
		.INIT('ha8)
	) name6348 (
		\sa11_reg[2]/P0001 ,
		_w6879_,
		_w6880_,
		_w6881_
	);
	LUT2 #(
		.INIT('h1)
	) name6349 (
		_w6878_,
		_w6881_,
		_w6882_
	);
	LUT3 #(
		.INIT('h2a)
	) name6350 (
		\sa11_reg[1]/P0001 ,
		_w6875_,
		_w6882_,
		_w6883_
	);
	LUT3 #(
		.INIT('h80)
	) name6351 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6884_
	);
	LUT3 #(
		.INIT('h01)
	) name6352 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6885_
	);
	LUT3 #(
		.INIT('h7e)
	) name6353 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6886_
	);
	LUT4 #(
		.INIT('h8002)
	) name6354 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6887_
	);
	LUT4 #(
		.INIT('hfbcc)
	) name6355 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6888_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name6356 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6887_,
		_w6888_,
		_w6889_
	);
	LUT4 #(
		.INIT('h0004)
	) name6357 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6890_
	);
	LUT4 #(
		.INIT('heffb)
	) name6358 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6891_
	);
	LUT2 #(
		.INIT('h2)
	) name6359 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[5]/P0001 ,
		_w6892_
	);
	LUT3 #(
		.INIT('h01)
	) name6360 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6893_
	);
	LUT4 #(
		.INIT('hfdf8)
	) name6361 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6894_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name6362 (
		\sa11_reg[7]/NET0131 ,
		_w6891_,
		_w6892_,
		_w6894_,
		_w6895_
	);
	LUT4 #(
		.INIT('h1000)
	) name6363 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6896_
	);
	LUT3 #(
		.INIT('h54)
	) name6364 (
		\sa11_reg[2]/P0001 ,
		_w6659_,
		_w6896_,
		_w6897_
	);
	LUT4 #(
		.INIT('h0001)
	) name6365 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6898_
	);
	LUT3 #(
		.INIT('h07)
	) name6366 (
		_w6636_,
		_w6665_,
		_w6898_,
		_w6899_
	);
	LUT4 #(
		.INIT('h3200)
	) name6367 (
		\sa11_reg[1]/P0001 ,
		_w6897_,
		_w6895_,
		_w6899_,
		_w6900_
	);
	LUT2 #(
		.INIT('h4)
	) name6368 (
		_w6889_,
		_w6900_,
		_w6901_
	);
	LUT3 #(
		.INIT('h20)
	) name6369 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w6902_
	);
	LUT3 #(
		.INIT('h6b)
	) name6370 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6903_
	);
	LUT2 #(
		.INIT('h2)
	) name6371 (
		_w6902_,
		_w6903_,
		_w6904_
	);
	LUT3 #(
		.INIT('h80)
	) name6372 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		_w6905_
	);
	LUT3 #(
		.INIT('h13)
	) name6373 (
		_w6654_,
		_w6719_,
		_w6905_,
		_w6906_
	);
	LUT3 #(
		.INIT('h45)
	) name6374 (
		\sa11_reg[1]/P0001 ,
		_w6904_,
		_w6906_,
		_w6907_
	);
	LUT2 #(
		.INIT('h1)
	) name6375 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[2]/P0001 ,
		_w6908_
	);
	LUT4 #(
		.INIT('h1000)
	) name6376 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6909_
	);
	LUT4 #(
		.INIT('h2000)
	) name6377 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6910_
	);
	LUT4 #(
		.INIT('h0007)
	) name6378 (
		_w6642_,
		_w6644_,
		_w6910_,
		_w6909_,
		_w6911_
	);
	LUT2 #(
		.INIT('h2)
	) name6379 (
		_w6908_,
		_w6911_,
		_w6912_
	);
	LUT2 #(
		.INIT('h8)
	) name6380 (
		_w6642_,
		_w6902_,
		_w6913_
	);
	LUT4 #(
		.INIT('h153f)
	) name6381 (
		\sa11_reg[3]/P0001 ,
		_w6636_,
		_w6665_,
		_w6898_,
		_w6914_
	);
	LUT3 #(
		.INIT('h8a)
	) name6382 (
		\sa11_reg[1]/P0001 ,
		_w6913_,
		_w6914_,
		_w6915_
	);
	LUT3 #(
		.INIT('h80)
	) name6383 (
		\sa11_reg[4]/P0001 ,
		_w6730_,
		_w6676_,
		_w6916_
	);
	LUT4 #(
		.INIT('h5540)
	) name6384 (
		\sa11_reg[2]/P0001 ,
		_w6666_,
		_w6694_,
		_w6680_,
		_w6917_
	);
	LUT2 #(
		.INIT('h1)
	) name6385 (
		_w6916_,
		_w6917_,
		_w6918_
	);
	LUT4 #(
		.INIT('h0100)
	) name6386 (
		_w6907_,
		_w6915_,
		_w6912_,
		_w6918_,
		_w6919_
	);
	LUT4 #(
		.INIT('hba00)
	) name6387 (
		\sa11_reg[0]/P0001 ,
		_w6883_,
		_w6901_,
		_w6919_,
		_w6920_
	);
	LUT2 #(
		.INIT('h2)
	) name6388 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w6921_
	);
	LUT3 #(
		.INIT('h20)
	) name6389 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		_w6922_
	);
	LUT2 #(
		.INIT('h8)
	) name6390 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w6923_
	);
	LUT3 #(
		.INIT('h23)
	) name6391 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w6924_
	);
	LUT4 #(
		.INIT('h0123)
	) name6392 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6925_
	);
	LUT3 #(
		.INIT('ha8)
	) name6393 (
		\sa22_reg[1]/P0001 ,
		_w6922_,
		_w6925_,
		_w6926_
	);
	LUT3 #(
		.INIT('h08)
	) name6394 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w6927_
	);
	LUT4 #(
		.INIT('h0080)
	) name6395 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6928_
	);
	LUT2 #(
		.INIT('h2)
	) name6396 (
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6929_
	);
	LUT4 #(
		.INIT('h0020)
	) name6397 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6930_
	);
	LUT3 #(
		.INIT('h04)
	) name6398 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w6931_
	);
	LUT3 #(
		.INIT('h01)
	) name6399 (
		_w6928_,
		_w6930_,
		_w6931_,
		_w6932_
	);
	LUT3 #(
		.INIT('h45)
	) name6400 (
		\sa22_reg[2]/P0001 ,
		_w6926_,
		_w6932_,
		_w6933_
	);
	LUT2 #(
		.INIT('h4)
	) name6401 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w6934_
	);
	LUT3 #(
		.INIT('h10)
	) name6402 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w6935_
	);
	LUT2 #(
		.INIT('h8)
	) name6403 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w6936_
	);
	LUT3 #(
		.INIT('h08)
	) name6404 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w6937_
	);
	LUT4 #(
		.INIT('h0008)
	) name6405 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6938_
	);
	LUT3 #(
		.INIT('ha8)
	) name6406 (
		\sa22_reg[2]/P0001 ,
		_w6935_,
		_w6938_,
		_w6939_
	);
	LUT2 #(
		.INIT('h2)
	) name6407 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w6940_
	);
	LUT4 #(
		.INIT('h0200)
	) name6408 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6941_
	);
	LUT2 #(
		.INIT('h4)
	) name6409 (
		\sa22_reg[2]/P0001 ,
		_w6941_,
		_w6942_
	);
	LUT2 #(
		.INIT('h4)
	) name6410 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w6943_
	);
	LUT2 #(
		.INIT('h8)
	) name6411 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w6944_
	);
	LUT3 #(
		.INIT('h80)
	) name6412 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6945_
	);
	LUT3 #(
		.INIT('h08)
	) name6413 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6946_
	);
	LUT2 #(
		.INIT('h2)
	) name6414 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		_w6947_
	);
	LUT4 #(
		.INIT('h7707)
	) name6415 (
		_w6943_,
		_w6945_,
		_w6946_,
		_w6947_,
		_w6948_
	);
	LUT4 #(
		.INIT('h5455)
	) name6416 (
		\sa22_reg[1]/P0001 ,
		_w6939_,
		_w6942_,
		_w6948_,
		_w6949_
	);
	LUT3 #(
		.INIT('h04)
	) name6417 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w6950_
	);
	LUT3 #(
		.INIT('h02)
	) name6418 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6951_
	);
	LUT4 #(
		.INIT('h153f)
	) name6419 (
		_w6936_,
		_w6923_,
		_w6950_,
		_w6951_,
		_w6952_
	);
	LUT2 #(
		.INIT('h1)
	) name6420 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w6953_
	);
	LUT3 #(
		.INIT('h04)
	) name6421 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w6954_
	);
	LUT4 #(
		.INIT('h0200)
	) name6422 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6955_
	);
	LUT3 #(
		.INIT('h07)
	) name6423 (
		_w6953_,
		_w6954_,
		_w6955_,
		_w6956_
	);
	LUT3 #(
		.INIT('h2a)
	) name6424 (
		\sa22_reg[1]/P0001 ,
		_w6952_,
		_w6956_,
		_w6957_
	);
	LUT3 #(
		.INIT('h20)
	) name6425 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w6958_
	);
	LUT4 #(
		.INIT('h2000)
	) name6426 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6959_
	);
	LUT2 #(
		.INIT('h4)
	) name6427 (
		\sa22_reg[2]/P0001 ,
		_w6959_,
		_w6960_
	);
	LUT3 #(
		.INIT('h80)
	) name6428 (
		\sa22_reg[2]/P0001 ,
		_w6943_,
		_w6945_,
		_w6961_
	);
	LUT2 #(
		.INIT('h1)
	) name6429 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w6962_
	);
	LUT4 #(
		.INIT('h0010)
	) name6430 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6963_
	);
	LUT4 #(
		.INIT('h0777)
	) name6431 (
		_w6921_,
		_w6946_,
		_w6947_,
		_w6963_,
		_w6964_
	);
	LUT3 #(
		.INIT('h10)
	) name6432 (
		_w6961_,
		_w6960_,
		_w6964_,
		_w6965_
	);
	LUT4 #(
		.INIT('h0100)
	) name6433 (
		_w6949_,
		_w6957_,
		_w6933_,
		_w6965_,
		_w6966_
	);
	LUT2 #(
		.INIT('h1)
	) name6434 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w6967_
	);
	LUT4 #(
		.INIT('h0010)
	) name6435 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6968_
	);
	LUT4 #(
		.INIT('h0040)
	) name6436 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w6969_
	);
	LUT3 #(
		.INIT('h01)
	) name6437 (
		\sa22_reg[2]/P0001 ,
		_w6968_,
		_w6969_,
		_w6970_
	);
	LUT3 #(
		.INIT('h08)
	) name6438 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6971_
	);
	LUT4 #(
		.INIT('h0080)
	) name6439 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6972_
	);
	LUT2 #(
		.INIT('h8)
	) name6440 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w6973_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6441 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w6974_
	);
	LUT2 #(
		.INIT('h4)
	) name6442 (
		_w6972_,
		_w6974_,
		_w6975_
	);
	LUT2 #(
		.INIT('h1)
	) name6443 (
		_w6970_,
		_w6975_,
		_w6976_
	);
	LUT3 #(
		.INIT('h02)
	) name6444 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w6977_
	);
	LUT4 #(
		.INIT('h0002)
	) name6445 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6978_
	);
	LUT2 #(
		.INIT('h2)
	) name6446 (
		\sa22_reg[1]/P0001 ,
		_w6978_,
		_w6979_
	);
	LUT4 #(
		.INIT('h1000)
	) name6447 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w6980_
	);
	LUT4 #(
		.INIT('h1000)
	) name6448 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6981_
	);
	LUT2 #(
		.INIT('h4)
	) name6449 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		_w6982_
	);
	LUT4 #(
		.INIT('h0400)
	) name6450 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6983_
	);
	LUT4 #(
		.INIT('h000b)
	) name6451 (
		\sa22_reg[7]/NET0131 ,
		_w6980_,
		_w6981_,
		_w6983_,
		_w6984_
	);
	LUT3 #(
		.INIT('h80)
	) name6452 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		_w6985_
	);
	LUT4 #(
		.INIT('h8000)
	) name6453 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w6986_
	);
	LUT3 #(
		.INIT('h20)
	) name6454 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6987_
	);
	LUT4 #(
		.INIT('h0400)
	) name6455 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6988_
	);
	LUT2 #(
		.INIT('h1)
	) name6456 (
		_w6986_,
		_w6988_,
		_w6989_
	);
	LUT3 #(
		.INIT('h80)
	) name6457 (
		_w6979_,
		_w6984_,
		_w6989_,
		_w6990_
	);
	LUT4 #(
		.INIT('h0100)
	) name6458 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6991_
	);
	LUT3 #(
		.INIT('h15)
	) name6459 (
		\sa22_reg[1]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w6991_,
		_w6992_
	);
	LUT2 #(
		.INIT('h2)
	) name6460 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w6993_
	);
	LUT2 #(
		.INIT('h8)
	) name6461 (
		_w6977_,
		_w6993_,
		_w6994_
	);
	LUT2 #(
		.INIT('h2)
	) name6462 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w6995_
	);
	LUT4 #(
		.INIT('h0002)
	) name6463 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6996_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name6464 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w6980_,
		_w6996_,
		_w6997_
	);
	LUT3 #(
		.INIT('h40)
	) name6465 (
		_w6994_,
		_w6992_,
		_w6997_,
		_w6998_
	);
	LUT3 #(
		.INIT('h9d)
	) name6466 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w6999_
	);
	LUT3 #(
		.INIT('h01)
	) name6467 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7000_
	);
	LUT4 #(
		.INIT('h0501)
	) name6468 (
		_w6986_,
		_w6962_,
		_w7000_,
		_w6999_,
		_w7001_
	);
	LUT4 #(
		.INIT('h0008)
	) name6469 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7002_
	);
	LUT4 #(
		.INIT('h1000)
	) name6470 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7003_
	);
	LUT2 #(
		.INIT('h1)
	) name6471 (
		_w7002_,
		_w7003_,
		_w7004_
	);
	LUT3 #(
		.INIT('h54)
	) name6472 (
		\sa22_reg[2]/P0001 ,
		_w7002_,
		_w7003_,
		_w7005_
	);
	LUT3 #(
		.INIT('h01)
	) name6473 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7006_
	);
	LUT4 #(
		.INIT('h0001)
	) name6474 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7007_
	);
	LUT4 #(
		.INIT('h0800)
	) name6475 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7008_
	);
	LUT3 #(
		.INIT('h23)
	) name6476 (
		\sa22_reg[2]/P0001 ,
		_w7007_,
		_w7008_,
		_w7009_
	);
	LUT4 #(
		.INIT('he400)
	) name6477 (
		\sa22_reg[2]/P0001 ,
		_w7004_,
		_w7001_,
		_w7009_,
		_w7010_
	);
	LUT4 #(
		.INIT('hf400)
	) name6478 (
		_w6976_,
		_w6990_,
		_w6998_,
		_w7010_,
		_w7011_
	);
	LUT3 #(
		.INIT('h6b)
	) name6479 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7012_
	);
	LUT3 #(
		.INIT('h20)
	) name6480 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w7013_
	);
	LUT2 #(
		.INIT('h4)
	) name6481 (
		_w7012_,
		_w7013_,
		_w7014_
	);
	LUT4 #(
		.INIT('h0001)
	) name6482 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7015_
	);
	LUT3 #(
		.INIT('h07)
	) name6483 (
		_w6985_,
		_w6995_,
		_w7015_,
		_w7016_
	);
	LUT3 #(
		.INIT('h45)
	) name6484 (
		\sa22_reg[1]/P0001 ,
		_w7014_,
		_w7016_,
		_w7017_
	);
	LUT3 #(
		.INIT('h80)
	) name6485 (
		\sa22_reg[2]/P0001 ,
		_w6944_,
		_w6954_,
		_w7018_
	);
	LUT3 #(
		.INIT('h01)
	) name6486 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7019_
	);
	LUT4 #(
		.INIT('h23af)
	) name6487 (
		\sa22_reg[2]/P0001 ,
		_w6940_,
		_w7008_,
		_w7019_,
		_w7020_
	);
	LUT3 #(
		.INIT('h8a)
	) name6488 (
		\sa22_reg[1]/P0001 ,
		_w7018_,
		_w7020_,
		_w7021_
	);
	LUT2 #(
		.INIT('h1)
	) name6489 (
		\sa22_reg[1]/P0001 ,
		\sa22_reg[2]/P0001 ,
		_w7022_
	);
	LUT3 #(
		.INIT('h10)
	) name6490 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7023_
	);
	LUT4 #(
		.INIT('h1000)
	) name6491 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7024_
	);
	LUT4 #(
		.INIT('h0007)
	) name6492 (
		_w6929_,
		_w6985_,
		_w6959_,
		_w7024_,
		_w7025_
	);
	LUT4 #(
		.INIT('h0080)
	) name6493 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7026_
	);
	LUT2 #(
		.INIT('h8)
	) name6494 (
		_w6995_,
		_w7026_,
		_w7027_
	);
	LUT4 #(
		.INIT('h5444)
	) name6495 (
		\sa22_reg[2]/P0001 ,
		_w6981_,
		_w6921_,
		_w6951_,
		_w7028_
	);
	LUT4 #(
		.INIT('h0051)
	) name6496 (
		_w7027_,
		_w7022_,
		_w7025_,
		_w7028_,
		_w7029_
	);
	LUT3 #(
		.INIT('h10)
	) name6497 (
		_w7017_,
		_w7021_,
		_w7029_,
		_w7030_
	);
	LUT4 #(
		.INIT('he400)
	) name6498 (
		\sa22_reg[0]/P0001 ,
		_w7011_,
		_w6966_,
		_w7030_,
		_w7031_
	);
	LUT3 #(
		.INIT('h4b)
	) name6499 (
		_w6867_,
		_w6920_,
		_w7031_,
		_w7032_
	);
	LUT2 #(
		.INIT('h2)
	) name6500 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7033_
	);
	LUT3 #(
		.INIT('h20)
	) name6501 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		_w7034_
	);
	LUT2 #(
		.INIT('h8)
	) name6502 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7035_
	);
	LUT4 #(
		.INIT('h0123)
	) name6503 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7036_
	);
	LUT3 #(
		.INIT('ha8)
	) name6504 (
		\sa33_reg[1]/P0001 ,
		_w7034_,
		_w7036_,
		_w7037_
	);
	LUT3 #(
		.INIT('h04)
	) name6505 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7038_
	);
	LUT2 #(
		.INIT('h2)
	) name6506 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		_w7039_
	);
	LUT3 #(
		.INIT('h08)
	) name6507 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7040_
	);
	LUT3 #(
		.INIT('h23)
	) name6508 (
		_w7039_,
		_w7038_,
		_w7040_,
		_w7041_
	);
	LUT3 #(
		.INIT('h45)
	) name6509 (
		\sa33_reg[2]/P0001 ,
		_w7037_,
		_w7041_,
		_w7042_
	);
	LUT2 #(
		.INIT('h8)
	) name6510 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7043_
	);
	LUT2 #(
		.INIT('h1)
	) name6511 (
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7044_
	);
	LUT4 #(
		.INIT('h0008)
	) name6512 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7045_
	);
	LUT3 #(
		.INIT('h10)
	) name6513 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7046_
	);
	LUT3 #(
		.INIT('ha8)
	) name6514 (
		\sa33_reg[2]/P0001 ,
		_w7045_,
		_w7046_,
		_w7047_
	);
	LUT2 #(
		.INIT('h8)
	) name6515 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7048_
	);
	LUT2 #(
		.INIT('h4)
	) name6516 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7049_
	);
	LUT3 #(
		.INIT('h40)
	) name6517 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7050_
	);
	LUT2 #(
		.INIT('h8)
	) name6518 (
		_w7048_,
		_w7050_,
		_w7051_
	);
	LUT2 #(
		.INIT('h4)
	) name6519 (
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7052_
	);
	LUT2 #(
		.INIT('h2)
	) name6520 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		_w7053_
	);
	LUT4 #(
		.INIT('h0200)
	) name6521 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7054_
	);
	LUT2 #(
		.INIT('h2)
	) name6522 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		_w7055_
	);
	LUT3 #(
		.INIT('h08)
	) name6523 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7056_
	);
	LUT4 #(
		.INIT('h22af)
	) name6524 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		_w7054_,
		_w7056_,
		_w7057_
	);
	LUT4 #(
		.INIT('h5455)
	) name6525 (
		\sa33_reg[1]/P0001 ,
		_w7047_,
		_w7051_,
		_w7057_,
		_w7058_
	);
	LUT4 #(
		.INIT('h4000)
	) name6526 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7059_
	);
	LUT4 #(
		.INIT('h0200)
	) name6527 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7060_
	);
	LUT3 #(
		.INIT('h0b)
	) name6528 (
		\sa33_reg[6]/P0001 ,
		_w7059_,
		_w7060_,
		_w7061_
	);
	LUT3 #(
		.INIT('h01)
	) name6529 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7062_
	);
	LUT4 #(
		.INIT('h0080)
	) name6530 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7063_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name6531 (
		\sa33_reg[6]/P0001 ,
		_w7049_,
		_w7062_,
		_w7063_,
		_w7064_
	);
	LUT3 #(
		.INIT('h2a)
	) name6532 (
		\sa33_reg[1]/P0001 ,
		_w7061_,
		_w7064_,
		_w7065_
	);
	LUT2 #(
		.INIT('h1)
	) name6533 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7066_
	);
	LUT3 #(
		.INIT('h04)
	) name6534 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7067_
	);
	LUT4 #(
		.INIT('h0777)
	) name6535 (
		_w7048_,
		_w7050_,
		_w7066_,
		_w7067_,
		_w7068_
	);
	LUT2 #(
		.INIT('h4)
	) name6536 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7069_
	);
	LUT4 #(
		.INIT('h2000)
	) name6537 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7070_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name6538 (
		\sa33_reg[2]/P0001 ,
		_w7033_,
		_w7056_,
		_w7070_,
		_w7071_
	);
	LUT3 #(
		.INIT('hd0)
	) name6539 (
		\sa33_reg[2]/P0001 ,
		_w7068_,
		_w7071_,
		_w7072_
	);
	LUT4 #(
		.INIT('h0100)
	) name6540 (
		_w7058_,
		_w7065_,
		_w7042_,
		_w7072_,
		_w7073_
	);
	LUT2 #(
		.INIT('h2)
	) name6541 (
		\sa33_reg[0]/P0001 ,
		_w7073_,
		_w7074_
	);
	LUT3 #(
		.INIT('h04)
	) name6542 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7075_
	);
	LUT4 #(
		.INIT('h0010)
	) name6543 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7076_
	);
	LUT2 #(
		.INIT('h2)
	) name6544 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7077_
	);
	LUT3 #(
		.INIT('h04)
	) name6545 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7078_
	);
	LUT4 #(
		.INIT('h0040)
	) name6546 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7079_
	);
	LUT3 #(
		.INIT('h20)
	) name6547 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7080_
	);
	LUT4 #(
		.INIT('h5554)
	) name6548 (
		\sa33_reg[2]/P0001 ,
		_w7079_,
		_w7080_,
		_w7076_,
		_w7081_
	);
	LUT3 #(
		.INIT('h80)
	) name6549 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7082_
	);
	LUT3 #(
		.INIT('h08)
	) name6550 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7083_
	);
	LUT4 #(
		.INIT('h0080)
	) name6551 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7084_
	);
	LUT3 #(
		.INIT('ha8)
	) name6552 (
		\sa33_reg[2]/P0001 ,
		_w7082_,
		_w7084_,
		_w7085_
	);
	LUT3 #(
		.INIT('h40)
	) name6553 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7086_
	);
	LUT2 #(
		.INIT('h4)
	) name6554 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		_w7087_
	);
	LUT4 #(
		.INIT('h0040)
	) name6555 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7088_
	);
	LUT4 #(
		.INIT('hcfbf)
	) name6556 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7089_
	);
	LUT2 #(
		.INIT('h1)
	) name6557 (
		\sa33_reg[3]/P0001 ,
		_w7089_,
		_w7090_
	);
	LUT3 #(
		.INIT('h02)
	) name6558 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7091_
	);
	LUT4 #(
		.INIT('h0002)
	) name6559 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7092_
	);
	LUT4 #(
		.INIT('h0400)
	) name6560 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7093_
	);
	LUT4 #(
		.INIT('h8000)
	) name6561 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7094_
	);
	LUT3 #(
		.INIT('h01)
	) name6562 (
		_w7093_,
		_w7094_,
		_w7092_,
		_w7095_
	);
	LUT4 #(
		.INIT('h0100)
	) name6563 (
		_w7090_,
		_w7085_,
		_w7081_,
		_w7095_,
		_w7096_
	);
	LUT2 #(
		.INIT('h2)
	) name6564 (
		\sa33_reg[1]/P0001 ,
		_w7096_,
		_w7097_
	);
	LUT3 #(
		.INIT('h02)
	) name6565 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		_w7098_
	);
	LUT4 #(
		.INIT('h0400)
	) name6566 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7099_
	);
	LUT4 #(
		.INIT('hf9fd)
	) name6567 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7100_
	);
	LUT2 #(
		.INIT('h1)
	) name6568 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7101_
	);
	LUT3 #(
		.INIT('h01)
	) name6569 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7102_
	);
	LUT4 #(
		.INIT('h0302)
	) name6570 (
		\sa33_reg[7]/NET0131 ,
		_w7094_,
		_w7102_,
		_w7100_,
		_w7103_
	);
	LUT2 #(
		.INIT('h2)
	) name6571 (
		\sa33_reg[2]/P0001 ,
		_w7103_,
		_w7104_
	);
	LUT3 #(
		.INIT('h10)
	) name6572 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7105_
	);
	LUT4 #(
		.INIT('h0777)
	) name6573 (
		_w7039_,
		_w7105_,
		_w7055_,
		_w7062_,
		_w7106_
	);
	LUT2 #(
		.INIT('h1)
	) name6574 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7107_
	);
	LUT3 #(
		.INIT('h08)
	) name6575 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7108_
	);
	LUT2 #(
		.INIT('h8)
	) name6576 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7109_
	);
	LUT3 #(
		.INIT('h80)
	) name6577 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7110_
	);
	LUT4 #(
		.INIT('h0777)
	) name6578 (
		_w7107_,
		_w7108_,
		_w7066_,
		_w7110_,
		_w7111_
	);
	LUT3 #(
		.INIT('h15)
	) name6579 (
		\sa33_reg[1]/P0001 ,
		_w7106_,
		_w7111_,
		_w7112_
	);
	LUT2 #(
		.INIT('h4)
	) name6580 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		_w7113_
	);
	LUT3 #(
		.INIT('h02)
	) name6581 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7114_
	);
	LUT2 #(
		.INIT('h4)
	) name6582 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7115_
	);
	LUT4 #(
		.INIT('h1000)
	) name6583 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7116_
	);
	LUT4 #(
		.INIT('haabf)
	) name6584 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		_w7114_,
		_w7116_,
		_w7117_
	);
	LUT4 #(
		.INIT('h0001)
	) name6585 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7118_
	);
	LUT4 #(
		.INIT('h0800)
	) name6586 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7119_
	);
	LUT3 #(
		.INIT('h23)
	) name6587 (
		\sa33_reg[2]/P0001 ,
		_w7118_,
		_w7119_,
		_w7120_
	);
	LUT2 #(
		.INIT('h8)
	) name6588 (
		_w7117_,
		_w7120_,
		_w7121_
	);
	LUT3 #(
		.INIT('h10)
	) name6589 (
		_w7104_,
		_w7112_,
		_w7121_,
		_w7122_
	);
	LUT3 #(
		.INIT('h10)
	) name6590 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7123_
	);
	LUT4 #(
		.INIT('h1000)
	) name6591 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7124_
	);
	LUT4 #(
		.INIT('h0007)
	) name6592 (
		\sa33_reg[6]/P0001 ,
		_w7063_,
		_w7070_,
		_w7124_,
		_w7125_
	);
	LUT3 #(
		.INIT('h10)
	) name6593 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7126_
	);
	LUT3 #(
		.INIT('h6b)
	) name6594 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7127_
	);
	LUT3 #(
		.INIT('h20)
	) name6595 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7128_
	);
	LUT2 #(
		.INIT('h4)
	) name6596 (
		_w7127_,
		_w7128_,
		_w7129_
	);
	LUT3 #(
		.INIT('h80)
	) name6597 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7130_
	);
	LUT4 #(
		.INIT('h0001)
	) name6598 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7131_
	);
	LUT3 #(
		.INIT('h07)
	) name6599 (
		_w7077_,
		_w7130_,
		_w7131_,
		_w7132_
	);
	LUT4 #(
		.INIT('h3200)
	) name6600 (
		\sa33_reg[2]/P0001 ,
		_w7129_,
		_w7125_,
		_w7132_,
		_w7133_
	);
	LUT4 #(
		.INIT('h0040)
	) name6601 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7134_
	);
	LUT3 #(
		.INIT('h80)
	) name6602 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7134_,
		_w7135_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name6603 (
		\sa33_reg[2]/P0001 ,
		_w7091_,
		_w7101_,
		_w7119_,
		_w7136_
	);
	LUT2 #(
		.INIT('h4)
	) name6604 (
		_w7135_,
		_w7136_,
		_w7137_
	);
	LUT2 #(
		.INIT('h8)
	) name6605 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		_w7138_
	);
	LUT3 #(
		.INIT('h02)
	) name6606 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7139_
	);
	LUT3 #(
		.INIT('h80)
	) name6607 (
		\sa33_reg[4]/P0001 ,
		_w7138_,
		_w7139_,
		_w7140_
	);
	LUT4 #(
		.INIT('h1000)
	) name6608 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7141_
	);
	LUT4 #(
		.INIT('h0020)
	) name6609 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7142_
	);
	LUT4 #(
		.INIT('h5150)
	) name6610 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7141_,
		_w7142_,
		_w7143_
	);
	LUT2 #(
		.INIT('h1)
	) name6611 (
		_w7140_,
		_w7143_,
		_w7144_
	);
	LUT4 #(
		.INIT('he400)
	) name6612 (
		\sa33_reg[1]/P0001 ,
		_w7133_,
		_w7137_,
		_w7144_,
		_w7145_
	);
	LUT4 #(
		.INIT('hba00)
	) name6613 (
		\sa33_reg[0]/P0001 ,
		_w7097_,
		_w7122_,
		_w7145_,
		_w7146_
	);
	LUT3 #(
		.INIT('h65)
	) name6614 (
		\u0_w_reg[0][29]/P0001 ,
		_w7074_,
		_w7146_,
		_w7147_
	);
	LUT4 #(
		.INIT('h4114)
	) name6615 (
		\ld_r_reg/P0001 ,
		_w6843_,
		_w7032_,
		_w7147_,
		_w7148_
	);
	LUT3 #(
		.INIT('h28)
	) name6616 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[125]/P0001 ,
		\u0_w_reg[0][29]/P0001 ,
		_w7149_
	);
	LUT2 #(
		.INIT('he)
	) name6617 (
		_w7148_,
		_w7149_,
		_w7150_
	);
	LUT4 #(
		.INIT('h0040)
	) name6618 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w7151_
	);
	LUT4 #(
		.INIT('h0010)
	) name6619 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7152_
	);
	LUT3 #(
		.INIT('h20)
	) name6620 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7153_
	);
	LUT4 #(
		.INIT('hf5ef)
	) name6621 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7154_
	);
	LUT3 #(
		.INIT('h45)
	) name6622 (
		\sa00_reg[2]/P0001 ,
		_w7151_,
		_w7154_,
		_w7155_
	);
	LUT4 #(
		.INIT('h0080)
	) name6623 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7156_
	);
	LUT3 #(
		.INIT('ha8)
	) name6624 (
		\sa00_reg[2]/P0001 ,
		_w6804_,
		_w7156_,
		_w7157_
	);
	LUT4 #(
		.INIT('h77ef)
	) name6625 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7158_
	);
	LUT4 #(
		.INIT('h0400)
	) name6626 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7159_
	);
	LUT4 #(
		.INIT('h0002)
	) name6627 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7160_
	);
	LUT4 #(
		.INIT('heffd)
	) name6628 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7161_
	);
	LUT4 #(
		.INIT('h0d00)
	) name6629 (
		\sa00_reg[5]/P0001 ,
		_w7158_,
		_w7159_,
		_w7161_,
		_w7162_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6630 (
		\sa00_reg[1]/P0001 ,
		_w7157_,
		_w7155_,
		_w7162_,
		_w7163_
	);
	LUT3 #(
		.INIT('h08)
	) name6631 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w7164_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name6632 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w7165_
	);
	LUT4 #(
		.INIT('h0400)
	) name6633 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7166_
	);
	LUT4 #(
		.INIT('h5501)
	) name6634 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w7165_,
		_w7166_,
		_w7167_
	);
	LUT3 #(
		.INIT('h54)
	) name6635 (
		\sa00_reg[1]/P0001 ,
		_w6824_,
		_w7167_,
		_w7168_
	);
	LUT3 #(
		.INIT('h80)
	) name6636 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w7169_
	);
	LUT3 #(
		.INIT('h01)
	) name6637 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w7170_
	);
	LUT3 #(
		.INIT('h7e)
	) name6638 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w7171_
	);
	LUT4 #(
		.INIT('h8002)
	) name6639 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w7172_
	);
	LUT3 #(
		.INIT('h01)
	) name6640 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7173_
	);
	LUT4 #(
		.INIT('h000b)
	) name6641 (
		\sa00_reg[7]/NET0131 ,
		_w6790_,
		_w7172_,
		_w7173_,
		_w7174_
	);
	LUT4 #(
		.INIT('h1000)
	) name6642 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7175_
	);
	LUT4 #(
		.INIT('h0008)
	) name6643 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w7176_
	);
	LUT2 #(
		.INIT('h1)
	) name6644 (
		_w7175_,
		_w7176_,
		_w7177_
	);
	LUT3 #(
		.INIT('h54)
	) name6645 (
		\sa00_reg[2]/P0001 ,
		_w7175_,
		_w7176_,
		_w7178_
	);
	LUT3 #(
		.INIT('h01)
	) name6646 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w7179_
	);
	LUT4 #(
		.INIT('h0001)
	) name6647 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7180_
	);
	LUT3 #(
		.INIT('h07)
	) name6648 (
		_w6772_,
		_w6740_,
		_w7180_,
		_w7181_
	);
	LUT4 #(
		.INIT('he400)
	) name6649 (
		\sa00_reg[2]/P0001 ,
		_w7177_,
		_w7174_,
		_w7181_,
		_w7182_
	);
	LUT4 #(
		.INIT('h5455)
	) name6650 (
		\sa00_reg[0]/P0001 ,
		_w7168_,
		_w7163_,
		_w7182_,
		_w7183_
	);
	LUT3 #(
		.INIT('ha8)
	) name6651 (
		\sa00_reg[2]/P0001 ,
		_w6809_,
		_w6766_,
		_w7184_
	);
	LUT2 #(
		.INIT('h4)
	) name6652 (
		\sa00_reg[2]/P0001 ,
		_w6813_,
		_w7185_
	);
	LUT3 #(
		.INIT('h08)
	) name6653 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7186_
	);
	LUT4 #(
		.INIT('h7077)
	) name6654 (
		_w6745_,
		_w6788_,
		_w6832_,
		_w7186_,
		_w7187_
	);
	LUT4 #(
		.INIT('h5455)
	) name6655 (
		\sa00_reg[1]/P0001 ,
		_w7185_,
		_w7184_,
		_w7187_,
		_w7188_
	);
	LUT4 #(
		.INIT('hff9d)
	) name6656 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w7189_
	);
	LUT2 #(
		.INIT('h2)
	) name6657 (
		\sa00_reg[7]/NET0131 ,
		_w7189_,
		_w7190_
	);
	LUT3 #(
		.INIT('h08)
	) name6658 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w7191_
	);
	LUT4 #(
		.INIT('h0777)
	) name6659 (
		_w6745_,
		_w6759_,
		_w6776_,
		_w7191_,
		_w7192_
	);
	LUT3 #(
		.INIT('h8a)
	) name6660 (
		\sa00_reg[1]/P0001 ,
		_w7190_,
		_w7192_,
		_w7193_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name6661 (
		\sa00_reg[5]/P0001 ,
		_w6745_,
		_w6788_,
		_w7152_,
		_w7194_
	);
	LUT2 #(
		.INIT('h8)
	) name6662 (
		_w6738_,
		_w7186_,
		_w7195_
	);
	LUT3 #(
		.INIT('h0d)
	) name6663 (
		\sa00_reg[2]/P0001 ,
		_w7194_,
		_w7195_,
		_w7196_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name6664 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7197_
	);
	LUT4 #(
		.INIT('h2044)
	) name6665 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7198_
	);
	LUT4 #(
		.INIT('h5554)
	) name6666 (
		\sa00_reg[2]/P0001 ,
		_w6819_,
		_w6777_,
		_w7198_,
		_w7199_
	);
	LUT2 #(
		.INIT('h2)
	) name6667 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[2]/P0001 ,
		_w7200_
	);
	LUT3 #(
		.INIT('h20)
	) name6668 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w7201_
	);
	LUT4 #(
		.INIT('hfedc)
	) name6669 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7202_
	);
	LUT3 #(
		.INIT('h8a)
	) name6670 (
		_w7200_,
		_w7201_,
		_w7202_,
		_w7203_
	);
	LUT2 #(
		.INIT('h1)
	) name6671 (
		_w7199_,
		_w7203_,
		_w7204_
	);
	LUT4 #(
		.INIT('h1000)
	) name6672 (
		_w7193_,
		_w7188_,
		_w7196_,
		_w7204_,
		_w7205_
	);
	LUT3 #(
		.INIT('h10)
	) name6673 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w7206_
	);
	LUT4 #(
		.INIT('h1000)
	) name6674 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w7207_
	);
	LUT4 #(
		.INIT('h2000)
	) name6675 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7208_
	);
	LUT4 #(
		.INIT('h0007)
	) name6676 (
		\sa00_reg[5]/P0001 ,
		_w6749_,
		_w7208_,
		_w7207_,
		_w7209_
	);
	LUT3 #(
		.INIT('h10)
	) name6677 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7210_
	);
	LUT3 #(
		.INIT('h04)
	) name6678 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7211_
	);
	LUT3 #(
		.INIT('h6b)
	) name6679 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7212_
	);
	LUT2 #(
		.INIT('h2)
	) name6680 (
		_w6746_,
		_w7212_,
		_w7213_
	);
	LUT4 #(
		.INIT('h0001)
	) name6681 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7214_
	);
	LUT3 #(
		.INIT('h07)
	) name6682 (
		_w6750_,
		_w7191_,
		_w7214_,
		_w7215_
	);
	LUT4 #(
		.INIT('h3200)
	) name6683 (
		\sa00_reg[2]/P0001 ,
		_w7213_,
		_w7209_,
		_w7215_,
		_w7216_
	);
	LUT2 #(
		.INIT('h8)
	) name6684 (
		_w6832_,
		_w7156_,
		_w7217_
	);
	LUT4 #(
		.INIT('h0777)
	) name6685 (
		_w6754_,
		_w6837_,
		_w6772_,
		_w6740_,
		_w7218_
	);
	LUT2 #(
		.INIT('h4)
	) name6686 (
		_w7217_,
		_w7218_,
		_w7219_
	);
	LUT3 #(
		.INIT('h40)
	) name6687 (
		\sa00_reg[7]/NET0131 ,
		_w6750_,
		_w7191_,
		_w7220_
	);
	LUT4 #(
		.INIT('h5540)
	) name6688 (
		\sa00_reg[2]/P0001 ,
		_w6738_,
		_w6784_,
		_w6771_,
		_w7221_
	);
	LUT2 #(
		.INIT('h1)
	) name6689 (
		_w7220_,
		_w7221_,
		_w7222_
	);
	LUT4 #(
		.INIT('he400)
	) name6690 (
		\sa00_reg[1]/P0001 ,
		_w7216_,
		_w7219_,
		_w7222_,
		_w7223_
	);
	LUT4 #(
		.INIT('h3100)
	) name6691 (
		\sa00_reg[0]/P0001 ,
		_w7183_,
		_w7205_,
		_w7223_,
		_w7224_
	);
	LUT3 #(
		.INIT('h20)
	) name6692 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7225_
	);
	LUT2 #(
		.INIT('h4)
	) name6693 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7226_
	);
	LUT4 #(
		.INIT('h0100)
	) name6694 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7227_
	);
	LUT4 #(
		.INIT('h5510)
	) name6695 (
		\sa22_reg[2]/P0001 ,
		_w6921_,
		_w7225_,
		_w7227_,
		_w7228_
	);
	LUT4 #(
		.INIT('h0080)
	) name6696 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7229_
	);
	LUT4 #(
		.INIT('h0080)
	) name6697 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7230_
	);
	LUT4 #(
		.INIT('h0007)
	) name6698 (
		_w6947_,
		_w6958_,
		_w7229_,
		_w7230_,
		_w7231_
	);
	LUT3 #(
		.INIT('h8a)
	) name6699 (
		\sa22_reg[1]/P0001 ,
		_w7228_,
		_w7231_,
		_w7232_
	);
	LUT4 #(
		.INIT('h0040)
	) name6700 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7233_
	);
	LUT2 #(
		.INIT('h4)
	) name6701 (
		\sa22_reg[2]/P0001 ,
		_w7233_,
		_w7234_
	);
	LUT3 #(
		.INIT('h80)
	) name6702 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7235_
	);
	LUT4 #(
		.INIT('h8000)
	) name6703 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7236_
	);
	LUT4 #(
		.INIT('h0002)
	) name6704 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7237_
	);
	LUT3 #(
		.INIT('h01)
	) name6705 (
		_w6996_,
		_w7237_,
		_w7236_,
		_w7238_
	);
	LUT3 #(
		.INIT('h45)
	) name6706 (
		\sa22_reg[1]/P0001 ,
		_w7234_,
		_w7238_,
		_w7239_
	);
	LUT4 #(
		.INIT('h0004)
	) name6707 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7240_
	);
	LUT4 #(
		.INIT('h3310)
	) name6708 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		_w6959_,
		_w7240_,
		_w7241_
	);
	LUT4 #(
		.INIT('h0100)
	) name6709 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7242_
	);
	LUT4 #(
		.INIT('haa20)
	) name6710 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7002_,
		_w7242_,
		_w7243_
	);
	LUT2 #(
		.INIT('h1)
	) name6711 (
		_w7241_,
		_w7243_,
		_w7244_
	);
	LUT4 #(
		.INIT('h5455)
	) name6712 (
		\sa22_reg[0]/P0001 ,
		_w7239_,
		_w7232_,
		_w7244_,
		_w7245_
	);
	LUT3 #(
		.INIT('hab)
	) name6713 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7246_
	);
	LUT2 #(
		.INIT('h2)
	) name6714 (
		_w6934_,
		_w7246_,
		_w7247_
	);
	LUT2 #(
		.INIT('h8)
	) name6715 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7248_
	);
	LUT3 #(
		.INIT('h80)
	) name6716 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7249_
	);
	LUT3 #(
		.INIT('h15)
	) name6717 (
		\sa22_reg[2]/P0001 ,
		_w6982_,
		_w7249_,
		_w7250_
	);
	LUT2 #(
		.INIT('h4)
	) name6718 (
		_w7247_,
		_w7250_,
		_w7251_
	);
	LUT3 #(
		.INIT('h2a)
	) name6719 (
		\sa22_reg[2]/P0001 ,
		_w6953_,
		_w7023_,
		_w7252_
	);
	LUT4 #(
		.INIT('h0020)
	) name6720 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7253_
	);
	LUT2 #(
		.INIT('h1)
	) name6721 (
		_w6928_,
		_w7253_,
		_w7254_
	);
	LUT3 #(
		.INIT('h80)
	) name6722 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7255_
	);
	LUT4 #(
		.INIT('h0004)
	) name6723 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7256_
	);
	LUT3 #(
		.INIT('h07)
	) name6724 (
		_w6953_,
		_w7255_,
		_w7256_,
		_w7257_
	);
	LUT3 #(
		.INIT('h80)
	) name6725 (
		_w7252_,
		_w7254_,
		_w7257_,
		_w7258_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name6726 (
		\sa22_reg[3]/P0001 ,
		_w6929_,
		_w6985_,
		_w7240_,
		_w7259_
	);
	LUT4 #(
		.INIT('h0155)
	) name6727 (
		\sa22_reg[1]/P0001 ,
		_w7251_,
		_w7258_,
		_w7259_,
		_w7260_
	);
	LUT4 #(
		.INIT('h0200)
	) name6728 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7261_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name6729 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7262_
	);
	LUT2 #(
		.INIT('h1)
	) name6730 (
		\sa22_reg[2]/P0001 ,
		_w7262_,
		_w7263_
	);
	LUT3 #(
		.INIT('h2a)
	) name6731 (
		\sa22_reg[1]/P0001 ,
		_w6921_,
		_w6951_,
		_w7264_
	);
	LUT4 #(
		.INIT('h0200)
	) name6732 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7265_
	);
	LUT3 #(
		.INIT('h07)
	) name6733 (
		_w6953_,
		_w6954_,
		_w7265_,
		_w7266_
	);
	LUT3 #(
		.INIT('h20)
	) name6734 (
		_w7264_,
		_w7263_,
		_w7266_,
		_w7267_
	);
	LUT2 #(
		.INIT('h1)
	) name6735 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7268_
	);
	LUT3 #(
		.INIT('h15)
	) name6736 (
		\sa22_reg[1]/P0001 ,
		_w6937_,
		_w7268_,
		_w7269_
	);
	LUT2 #(
		.INIT('h8)
	) name6737 (
		\sa22_reg[2]/P0001 ,
		_w7008_,
		_w7270_
	);
	LUT4 #(
		.INIT('h2000)
	) name6738 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7271_
	);
	LUT2 #(
		.INIT('h1)
	) name6739 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w7272_
	);
	LUT3 #(
		.INIT('h32)
	) name6740 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w7273_
	);
	LUT3 #(
		.INIT('h31)
	) name6741 (
		_w6973_,
		_w7271_,
		_w7273_,
		_w7274_
	);
	LUT3 #(
		.INIT('h20)
	) name6742 (
		_w7269_,
		_w7270_,
		_w7274_,
		_w7275_
	);
	LUT2 #(
		.INIT('h4)
	) name6743 (
		\sa22_reg[3]/P0001 ,
		_w7007_,
		_w7276_
	);
	LUT4 #(
		.INIT('h2000)
	) name6744 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7277_
	);
	LUT3 #(
		.INIT('h01)
	) name6745 (
		\sa22_reg[2]/P0001 ,
		_w6930_,
		_w7277_,
		_w7278_
	);
	LUT4 #(
		.INIT('h4000)
	) name6746 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7279_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name6747 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7280_
	);
	LUT4 #(
		.INIT('h0200)
	) name6748 (
		\sa22_reg[2]/P0001 ,
		_w6941_,
		_w7279_,
		_w7280_,
		_w7281_
	);
	LUT3 #(
		.INIT('h0b)
	) name6749 (
		_w7276_,
		_w7278_,
		_w7281_,
		_w7282_
	);
	LUT4 #(
		.INIT('haa02)
	) name6750 (
		\sa22_reg[0]/P0001 ,
		_w7267_,
		_w7275_,
		_w7282_,
		_w7283_
	);
	LUT4 #(
		.INIT('h2220)
	) name6751 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7284_
	);
	LUT3 #(
		.INIT('h07)
	) name6752 (
		\sa22_reg[7]/NET0131 ,
		_w6980_,
		_w7284_,
		_w7285_
	);
	LUT3 #(
		.INIT('h45)
	) name6753 (
		\sa22_reg[2]/P0001 ,
		_w7276_,
		_w7285_,
		_w7286_
	);
	LUT3 #(
		.INIT('h20)
	) name6754 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7287_
	);
	LUT4 #(
		.INIT('h135f)
	) name6755 (
		_w6995_,
		_w6923_,
		_w6927_,
		_w7287_,
		_w7288_
	);
	LUT4 #(
		.INIT('h2a7f)
	) name6756 (
		\sa22_reg[4]/P0001 ,
		_w6929_,
		_w6947_,
		_w6941_,
		_w7289_
	);
	LUT2 #(
		.INIT('h8)
	) name6757 (
		_w7288_,
		_w7289_,
		_w7290_
	);
	LUT4 #(
		.INIT('h0020)
	) name6758 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7291_
	);
	LUT2 #(
		.INIT('h8)
	) name6759 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		_w7292_
	);
	LUT4 #(
		.INIT('h0777)
	) name6760 (
		_w7272_,
		_w7291_,
		_w7292_,
		_w7235_,
		_w7293_
	);
	LUT4 #(
		.INIT('h7500)
	) name6761 (
		\sa22_reg[1]/P0001 ,
		_w7286_,
		_w7290_,
		_w7293_,
		_w7294_
	);
	LUT4 #(
		.INIT('h0100)
	) name6762 (
		_w7245_,
		_w7283_,
		_w7260_,
		_w7294_,
		_w7295_
	);
	LUT3 #(
		.INIT('h69)
	) name6763 (
		_w6737_,
		_w7224_,
		_w7295_,
		_w7296_
	);
	LUT4 #(
		.INIT('h9699)
	) name6764 (
		\u0_w_reg[0][21]/P0001 ,
		_w7031_,
		_w7074_,
		_w7146_,
		_w7297_
	);
	LUT3 #(
		.INIT('h82)
	) name6765 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[117]/P0001 ,
		\u0_w_reg[0][21]/P0001 ,
		_w7298_
	);
	LUT4 #(
		.INIT('h00eb)
	) name6766 (
		\ld_r_reg/P0001 ,
		_w7296_,
		_w7297_,
		_w7298_,
		_w7299_
	);
	LUT3 #(
		.INIT('h4b)
	) name6767 (
		_w6867_,
		_w6920_,
		_w7224_,
		_w7300_
	);
	LUT4 #(
		.INIT('hb44b)
	) name6768 (
		_w6867_,
		_w6920_,
		_w7224_,
		_w7295_,
		_w7301_
	);
	LUT3 #(
		.INIT('h10)
	) name6769 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7302_
	);
	LUT3 #(
		.INIT('hd3)
	) name6770 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		_w7303_
	);
	LUT2 #(
		.INIT('h8)
	) name6771 (
		_w7302_,
		_w7303_,
		_w7304_
	);
	LUT4 #(
		.INIT('h0080)
	) name6772 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7305_
	);
	LUT2 #(
		.INIT('h8)
	) name6773 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7306_
	);
	LUT4 #(
		.INIT('h0080)
	) name6774 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7307_
	);
	LUT4 #(
		.INIT('h0007)
	) name6775 (
		_w7115_,
		_w7128_,
		_w7307_,
		_w7305_,
		_w7308_
	);
	LUT3 #(
		.INIT('h8a)
	) name6776 (
		\sa33_reg[1]/P0001 ,
		_w7304_,
		_w7308_,
		_w7309_
	);
	LUT4 #(
		.INIT('h7f7c)
	) name6777 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7310_
	);
	LUT4 #(
		.INIT('h0002)
	) name6778 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7311_
	);
	LUT4 #(
		.INIT('h5504)
	) name6779 (
		\sa33_reg[1]/P0001 ,
		\sa33_reg[2]/P0001 ,
		_w7310_,
		_w7311_,
		_w7312_
	);
	LUT4 #(
		.INIT('h0040)
	) name6780 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7313_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name6781 (
		\sa33_reg[1]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7141_,
		_w7313_,
		_w7314_
	);
	LUT2 #(
		.INIT('h8)
	) name6782 (
		_w7066_,
		_w7139_,
		_w7315_
	);
	LUT4 #(
		.INIT('h0100)
	) name6783 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7316_
	);
	LUT3 #(
		.INIT('h07)
	) name6784 (
		_w7043_,
		_w7062_,
		_w7316_,
		_w7317_
	);
	LUT4 #(
		.INIT('h3210)
	) name6785 (
		\sa33_reg[2]/P0001 ,
		_w7315_,
		_w7314_,
		_w7317_,
		_w7318_
	);
	LUT4 #(
		.INIT('h5455)
	) name6786 (
		\sa33_reg[0]/P0001 ,
		_w7312_,
		_w7309_,
		_w7318_,
		_w7319_
	);
	LUT3 #(
		.INIT('h2a)
	) name6787 (
		\sa33_reg[2]/P0001 ,
		_w7107_,
		_w7123_,
		_w7320_
	);
	LUT4 #(
		.INIT('h0004)
	) name6788 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7321_
	);
	LUT2 #(
		.INIT('h1)
	) name6789 (
		_w7142_,
		_w7321_,
		_w7322_
	);
	LUT4 #(
		.INIT('h0080)
	) name6790 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7323_
	);
	LUT3 #(
		.INIT('h07)
	) name6791 (
		_w7080_,
		_w7039_,
		_w7323_,
		_w7324_
	);
	LUT3 #(
		.INIT('h80)
	) name6792 (
		_w7320_,
		_w7322_,
		_w7324_,
		_w7325_
	);
	LUT2 #(
		.INIT('h1)
	) name6793 (
		\sa33_reg[2]/P0001 ,
		_w7099_,
		_w7326_
	);
	LUT3 #(
		.INIT('h07)
	) name6794 (
		_w7033_,
		_w7110_,
		_w7141_,
		_w7327_
	);
	LUT2 #(
		.INIT('h8)
	) name6795 (
		_w7326_,
		_w7327_,
		_w7328_
	);
	LUT4 #(
		.INIT('h135f)
	) name6796 (
		\sa33_reg[6]/P0001 ,
		_w7066_,
		_w7063_,
		_w7139_,
		_w7329_
	);
	LUT4 #(
		.INIT('h0155)
	) name6797 (
		\sa33_reg[1]/P0001 ,
		_w7325_,
		_w7328_,
		_w7329_,
		_w7330_
	);
	LUT3 #(
		.INIT('h8a)
	) name6798 (
		\sa33_reg[1]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7142_,
		_w7331_
	);
	LUT3 #(
		.INIT('he0)
	) name6799 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7332_
	);
	LUT4 #(
		.INIT('h5410)
	) name6800 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7333_
	);
	LUT2 #(
		.INIT('h4)
	) name6801 (
		_w7332_,
		_w7333_,
		_w7334_
	);
	LUT2 #(
		.INIT('h2)
	) name6802 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7335_
	);
	LUT4 #(
		.INIT('h0200)
	) name6803 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7336_
	);
	LUT3 #(
		.INIT('h07)
	) name6804 (
		_w7049_,
		_w7062_,
		_w7336_,
		_w7337_
	);
	LUT3 #(
		.INIT('h40)
	) name6805 (
		_w7334_,
		_w7331_,
		_w7337_,
		_w7338_
	);
	LUT2 #(
		.INIT('h8)
	) name6806 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7339_
	);
	LUT4 #(
		.INIT('h2000)
	) name6807 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7340_
	);
	LUT3 #(
		.INIT('h08)
	) name6808 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7341_
	);
	LUT2 #(
		.INIT('h1)
	) name6809 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7342_
	);
	LUT4 #(
		.INIT('h0111)
	) name6810 (
		\sa33_reg[1]/P0001 ,
		_w7340_,
		_w7341_,
		_w7342_,
		_w7343_
	);
	LUT2 #(
		.INIT('h1)
	) name6811 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7344_
	);
	LUT3 #(
		.INIT('h32)
	) name6812 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7345_
	);
	LUT4 #(
		.INIT('h5f13)
	) name6813 (
		\sa33_reg[2]/P0001 ,
		_w7048_,
		_w7119_,
		_w7345_,
		_w7346_
	);
	LUT2 #(
		.INIT('h8)
	) name6814 (
		_w7343_,
		_w7346_,
		_w7347_
	);
	LUT2 #(
		.INIT('h8)
	) name6815 (
		_w7110_,
		_w7335_,
		_w7348_
	);
	LUT2 #(
		.INIT('h6)
	) name6816 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7349_
	);
	LUT4 #(
		.INIT('h0246)
	) name6817 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7350_
	);
	LUT3 #(
		.INIT('h02)
	) name6818 (
		\sa33_reg[2]/P0001 ,
		_w7054_,
		_w7350_,
		_w7351_
	);
	LUT2 #(
		.INIT('h4)
	) name6819 (
		\sa33_reg[5]/P0001 ,
		_w7131_,
		_w7352_
	);
	LUT4 #(
		.INIT('h2000)
	) name6820 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7353_
	);
	LUT4 #(
		.INIT('h0020)
	) name6821 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7354_
	);
	LUT3 #(
		.INIT('h01)
	) name6822 (
		\sa33_reg[2]/P0001 ,
		_w7353_,
		_w7354_,
		_w7355_
	);
	LUT4 #(
		.INIT('h4544)
	) name6823 (
		_w7348_,
		_w7351_,
		_w7352_,
		_w7355_,
		_w7356_
	);
	LUT4 #(
		.INIT('h02aa)
	) name6824 (
		\sa33_reg[0]/P0001 ,
		_w7338_,
		_w7347_,
		_w7356_,
		_w7357_
	);
	LUT4 #(
		.INIT('h2220)
	) name6825 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7358_
	);
	LUT3 #(
		.INIT('h07)
	) name6826 (
		_w7066_,
		_w7110_,
		_w7358_,
		_w7359_
	);
	LUT3 #(
		.INIT('h45)
	) name6827 (
		\sa33_reg[2]/P0001 ,
		_w7352_,
		_w7359_,
		_w7360_
	);
	LUT4 #(
		.INIT('h57df)
	) name6828 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		_w7083_,
		_w7139_,
		_w7361_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name6829 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7086_,
		_w7126_,
		_w7362_
	);
	LUT2 #(
		.INIT('h8)
	) name6830 (
		_w7361_,
		_w7362_,
		_w7363_
	);
	LUT4 #(
		.INIT('h0010)
	) name6831 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7364_
	);
	LUT4 #(
		.INIT('h153f)
	) name6832 (
		_w7113_,
		_w7109_,
		_w7130_,
		_w7364_,
		_w7365_
	);
	LUT4 #(
		.INIT('h7500)
	) name6833 (
		\sa33_reg[1]/P0001 ,
		_w7360_,
		_w7363_,
		_w7365_,
		_w7366_
	);
	LUT4 #(
		.INIT('h0100)
	) name6834 (
		_w7357_,
		_w7330_,
		_w7319_,
		_w7366_,
		_w7367_
	);
	LUT4 #(
		.INIT('h9a65)
	) name6835 (
		\u0_w_reg[0][13]/P0001 ,
		_w7074_,
		_w7146_,
		_w7367_,
		_w7368_
	);
	LUT3 #(
		.INIT('h28)
	) name6836 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[109]/P0001 ,
		\u0_w_reg[0][13]/P0001 ,
		_w7369_
	);
	LUT4 #(
		.INIT('hff41)
	) name6837 (
		\ld_r_reg/P0001 ,
		_w7301_,
		_w7368_,
		_w7369_,
		_w7370_
	);
	LUT4 #(
		.INIT('h9a65)
	) name6838 (
		_w6842_,
		_w6867_,
		_w6920_,
		_w7224_,
		_w7371_
	);
	LUT3 #(
		.INIT('h69)
	) name6839 (
		\u0_w_reg[0][5]/P0001 ,
		_w7031_,
		_w7367_,
		_w7372_
	);
	LUT3 #(
		.INIT('h28)
	) name6840 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[101]/P0001 ,
		\u0_w_reg[0][5]/P0001 ,
		_w7373_
	);
	LUT4 #(
		.INIT('hff41)
	) name6841 (
		\ld_r_reg/P0001 ,
		_w7371_,
		_w7372_,
		_w7373_,
		_w7374_
	);
	LUT3 #(
		.INIT('h15)
	) name6842 (
		_w6802_,
		_w6805_,
		_w6770_,
		_w7375_
	);
	LUT3 #(
		.INIT('h45)
	) name6843 (
		\sa00_reg[1]/P0001 ,
		_w7178_,
		_w7375_,
		_w7376_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name6844 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7377_
	);
	LUT4 #(
		.INIT('h20aa)
	) name6845 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w6771_,
		_w7377_,
		_w7378_
	);
	LUT4 #(
		.INIT('h0007)
	) name6846 (
		_w6745_,
		_w6788_,
		_w6749_,
		_w7180_,
		_w7379_
	);
	LUT3 #(
		.INIT('h8a)
	) name6847 (
		\sa00_reg[2]/P0001 ,
		_w7378_,
		_w7379_,
		_w7380_
	);
	LUT4 #(
		.INIT('h2000)
	) name6848 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w7381_
	);
	LUT3 #(
		.INIT('h07)
	) name6849 (
		_w6776_,
		_w7191_,
		_w7381_,
		_w7382_
	);
	LUT4 #(
		.INIT('haa80)
	) name6850 (
		\sa00_reg[1]/P0001 ,
		_w6776_,
		_w7191_,
		_w7381_,
		_w7383_
	);
	LUT3 #(
		.INIT('h02)
	) name6851 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w7384_
	);
	LUT4 #(
		.INIT('h0040)
	) name6852 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7385_
	);
	LUT4 #(
		.INIT('h0203)
	) name6853 (
		_w6838_,
		_w7151_,
		_w7385_,
		_w7384_,
		_w7386_
	);
	LUT2 #(
		.INIT('h2)
	) name6854 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w7387_
	);
	LUT2 #(
		.INIT('h8)
	) name6855 (
		_w7153_,
		_w7387_,
		_w7388_
	);
	LUT2 #(
		.INIT('h4)
	) name6856 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[2]/P0001 ,
		_w7389_
	);
	LUT3 #(
		.INIT('he0)
	) name6857 (
		_w6828_,
		_w7211_,
		_w7389_,
		_w7390_
	);
	LUT4 #(
		.INIT('h0032)
	) name6858 (
		\sa00_reg[2]/P0001 ,
		_w7388_,
		_w7386_,
		_w7390_,
		_w7391_
	);
	LUT4 #(
		.INIT('h0100)
	) name6859 (
		_w7380_,
		_w7383_,
		_w7376_,
		_w7391_,
		_w7392_
	);
	LUT3 #(
		.INIT('h02)
	) name6860 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w7393_
	);
	LUT4 #(
		.INIT('h0004)
	) name6861 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w7394_
	);
	LUT3 #(
		.INIT('h01)
	) name6862 (
		\sa00_reg[2]/P0001 ,
		_w6817_,
		_w7394_,
		_w7395_
	);
	LUT4 #(
		.INIT('h0040)
	) name6863 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w7396_
	);
	LUT4 #(
		.INIT('h23af)
	) name6864 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w6825_,
		_w7396_,
		_w7397_
	);
	LUT4 #(
		.INIT('h0001)
	) name6865 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w7398_
	);
	LUT3 #(
		.INIT('h40)
	) name6866 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w7399_
	);
	LUT4 #(
		.INIT('h002a)
	) name6867 (
		\sa00_reg[2]/P0001 ,
		_w6744_,
		_w7399_,
		_w7398_,
		_w7400_
	);
	LUT3 #(
		.INIT('h07)
	) name6868 (
		_w7395_,
		_w7397_,
		_w7400_,
		_w7401_
	);
	LUT2 #(
		.INIT('h4)
	) name6869 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		_w7402_
	);
	LUT4 #(
		.INIT('h4000)
	) name6870 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w7403_
	);
	LUT4 #(
		.INIT('h0001)
	) name6871 (
		\sa00_reg[1]/P0001 ,
		_w6829_,
		_w7385_,
		_w7403_,
		_w7404_
	);
	LUT3 #(
		.INIT('h10)
	) name6872 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7405_
	);
	LUT4 #(
		.INIT('h0100)
	) name6873 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7406_
	);
	LUT4 #(
		.INIT('h0777)
	) name6874 (
		_w6784_,
		_w6831_,
		_w6744_,
		_w7399_,
		_w7407_
	);
	LUT3 #(
		.INIT('h40)
	) name6875 (
		_w7406_,
		_w7404_,
		_w7407_,
		_w7408_
	);
	LUT2 #(
		.INIT('h4)
	) name6876 (
		\sa00_reg[2]/P0001 ,
		_w7180_,
		_w7409_
	);
	LUT2 #(
		.INIT('h2)
	) name6877 (
		_w6832_,
		_w7171_,
		_w7410_
	);
	LUT3 #(
		.INIT('h2a)
	) name6878 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w6749_,
		_w7411_
	);
	LUT3 #(
		.INIT('h10)
	) name6879 (
		_w7410_,
		_w7409_,
		_w7411_,
		_w7412_
	);
	LUT3 #(
		.INIT('h54)
	) name6880 (
		_w7401_,
		_w7408_,
		_w7412_,
		_w7413_
	);
	LUT4 #(
		.INIT('h0800)
	) name6881 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7414_
	);
	LUT4 #(
		.INIT('h0020)
	) name6882 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7415_
	);
	LUT4 #(
		.INIT('hf7df)
	) name6883 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7416_
	);
	LUT3 #(
		.INIT('h45)
	) name6884 (
		\sa00_reg[2]/P0001 ,
		_w7414_,
		_w7416_,
		_w7417_
	);
	LUT4 #(
		.INIT('h1000)
	) name6885 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w7418_
	);
	LUT3 #(
		.INIT('h40)
	) name6886 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7419_
	);
	LUT3 #(
		.INIT('h13)
	) name6887 (
		_w6750_,
		_w7418_,
		_w7419_,
		_w7420_
	);
	LUT4 #(
		.INIT('h0800)
	) name6888 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7421_
	);
	LUT3 #(
		.INIT('h07)
	) name6889 (
		_w6831_,
		_w7173_,
		_w7421_,
		_w7422_
	);
	LUT4 #(
		.INIT('h4555)
	) name6890 (
		\sa00_reg[1]/P0001 ,
		_w7417_,
		_w7420_,
		_w7422_,
		_w7423_
	);
	LUT3 #(
		.INIT('h40)
	) name6891 (
		\sa00_reg[2]/P0001 ,
		_w6738_,
		_w6784_,
		_w7424_
	);
	LUT4 #(
		.INIT('h0002)
	) name6892 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7425_
	);
	LUT4 #(
		.INIT('h0007)
	) name6893 (
		_w6803_,
		_w6754_,
		_w7214_,
		_w7425_,
		_w7426_
	);
	LUT4 #(
		.INIT('h20a8)
	) name6894 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[2]/P0001 ,
		_w6798_,
		_w7426_,
		_w7427_
	);
	LUT4 #(
		.INIT('hff7a)
	) name6895 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7428_
	);
	LUT2 #(
		.INIT('h2)
	) name6896 (
		_w7387_,
		_w7428_,
		_w7429_
	);
	LUT4 #(
		.INIT('h135f)
	) name6897 (
		_w6759_,
		_w6802_,
		_w6815_,
		_w7402_,
		_w7430_
	);
	LUT2 #(
		.INIT('h4)
	) name6898 (
		_w7429_,
		_w7430_,
		_w7431_
	);
	LUT3 #(
		.INIT('h10)
	) name6899 (
		_w7427_,
		_w7423_,
		_w7431_,
		_w7432_
	);
	LUT4 #(
		.INIT('hd800)
	) name6900 (
		\sa00_reg[0]/P0001 ,
		_w7392_,
		_w7413_,
		_w7432_,
		_w7433_
	);
	LUT2 #(
		.INIT('h4)
	) name6901 (
		\sa11_reg[2]/P0001 ,
		_w6677_,
		_w7434_
	);
	LUT4 #(
		.INIT('h1113)
	) name6902 (
		\sa11_reg[2]/P0001 ,
		_w6704_,
		_w6675_,
		_w6861_,
		_w7435_
	);
	LUT4 #(
		.INIT('h5455)
	) name6903 (
		\sa11_reg[1]/P0001 ,
		_w6897_,
		_w7434_,
		_w7435_,
		_w7436_
	);
	LUT3 #(
		.INIT('h08)
	) name6904 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7437_
	);
	LUT4 #(
		.INIT('h0400)
	) name6905 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7438_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name6906 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7439_
	);
	LUT4 #(
		.INIT('h20aa)
	) name6907 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w6896_,
		_w7439_,
		_w7440_
	);
	LUT2 #(
		.INIT('h1)
	) name6908 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w7441_
	);
	LUT3 #(
		.INIT('h01)
	) name6909 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		_w7442_
	);
	LUT2 #(
		.INIT('h4)
	) name6910 (
		_w6712_,
		_w7442_,
		_w7443_
	);
	LUT4 #(
		.INIT('h2000)
	) name6911 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w7444_
	);
	LUT3 #(
		.INIT('h07)
	) name6912 (
		_w6644_,
		_w6676_,
		_w7444_,
		_w7445_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6913 (
		\sa11_reg[1]/P0001 ,
		_w7440_,
		_w7443_,
		_w7445_,
		_w7446_
	);
	LUT2 #(
		.INIT('h1)
	) name6914 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w7447_
	);
	LUT4 #(
		.INIT('h0040)
	) name6915 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7448_
	);
	LUT3 #(
		.INIT('h54)
	) name6916 (
		\sa11_reg[2]/P0001 ,
		_w6876_,
		_w7448_,
		_w7449_
	);
	LUT3 #(
		.INIT('h23)
	) name6917 (
		\sa11_reg[3]/P0001 ,
		_w6645_,
		_w6848_,
		_w7450_
	);
	LUT2 #(
		.INIT('h1)
	) name6918 (
		_w6714_,
		_w6898_,
		_w7451_
	);
	LUT4 #(
		.INIT('h3111)
	) name6919 (
		\sa11_reg[2]/P0001 ,
		_w7449_,
		_w7450_,
		_w7451_,
		_w7452_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6920 (
		\sa11_reg[0]/P0001 ,
		_w7446_,
		_w7436_,
		_w7452_,
		_w7453_
	);
	LUT3 #(
		.INIT('h01)
	) name6921 (
		\sa11_reg[2]/P0001 ,
		_w6717_,
		_w6890_,
		_w7454_
	);
	LUT4 #(
		.INIT('h0040)
	) name6922 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w7455_
	);
	LUT4 #(
		.INIT('h23af)
	) name6923 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6726_,
		_w7455_,
		_w7456_
	);
	LUT3 #(
		.INIT('h40)
	) name6924 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w7457_
	);
	LUT4 #(
		.INIT('h0001)
	) name6925 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w7458_
	);
	LUT4 #(
		.INIT('h002a)
	) name6926 (
		\sa11_reg[2]/P0001 ,
		_w6637_,
		_w7457_,
		_w7458_,
		_w7459_
	);
	LUT3 #(
		.INIT('h07)
	) name6927 (
		_w7454_,
		_w7456_,
		_w7459_,
		_w7460_
	);
	LUT4 #(
		.INIT('h0200)
	) name6928 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w7461_
	);
	LUT3 #(
		.INIT('h01)
	) name6929 (
		\sa11_reg[1]/P0001 ,
		_w7448_,
		_w7461_,
		_w7462_
	);
	LUT4 #(
		.INIT('h153f)
	) name6930 (
		_w6637_,
		_w6730_,
		_w6676_,
		_w7457_,
		_w7463_
	);
	LUT4 #(
		.INIT('h4000)
	) name6931 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w7464_
	);
	LUT3 #(
		.INIT('h10)
	) name6932 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7465_
	);
	LUT4 #(
		.INIT('h0100)
	) name6933 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7466_
	);
	LUT2 #(
		.INIT('h1)
	) name6934 (
		_w7464_,
		_w7466_,
		_w7467_
	);
	LUT3 #(
		.INIT('h80)
	) name6935 (
		_w7462_,
		_w7463_,
		_w7467_,
		_w7468_
	);
	LUT2 #(
		.INIT('h2)
	) name6936 (
		_w6640_,
		_w6886_,
		_w7469_
	);
	LUT2 #(
		.INIT('h4)
	) name6937 (
		\sa11_reg[2]/P0001 ,
		_w6898_,
		_w7470_
	);
	LUT3 #(
		.INIT('h2a)
	) name6938 (
		\sa11_reg[1]/P0001 ,
		_w6642_,
		_w6644_,
		_w7471_
	);
	LUT3 #(
		.INIT('h10)
	) name6939 (
		_w7469_,
		_w7470_,
		_w7471_,
		_w7472_
	);
	LUT4 #(
		.INIT('h4445)
	) name6940 (
		\sa11_reg[0]/P0001 ,
		_w7460_,
		_w7468_,
		_w7472_,
		_w7473_
	);
	LUT4 #(
		.INIT('h0020)
	) name6941 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7474_
	);
	LUT4 #(
		.INIT('h5504)
	) name6942 (
		\sa11_reg[2]/P0001 ,
		_w6636_,
		_w6686_,
		_w7474_,
		_w7475_
	);
	LUT3 #(
		.INIT('ha8)
	) name6943 (
		\sa11_reg[2]/P0001 ,
		_w6653_,
		_w6713_,
		_w7476_
	);
	LUT4 #(
		.INIT('h0800)
	) name6944 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7477_
	);
	LUT2 #(
		.INIT('h1)
	) name6945 (
		_w6870_,
		_w7477_,
		_w7478_
	);
	LUT4 #(
		.INIT('h5455)
	) name6946 (
		\sa11_reg[1]/P0001 ,
		_w7476_,
		_w7475_,
		_w7478_,
		_w7479_
	);
	LUT2 #(
		.INIT('h8)
	) name6947 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[2]/P0001 ,
		_w7480_
	);
	LUT4 #(
		.INIT('h0002)
	) name6948 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7481_
	);
	LUT4 #(
		.INIT('h0013)
	) name6949 (
		\sa11_reg[3]/P0001 ,
		_w6719_,
		_w7438_,
		_w7481_,
		_w7482_
	);
	LUT2 #(
		.INIT('h2)
	) name6950 (
		_w7480_,
		_w7482_,
		_w7483_
	);
	LUT2 #(
		.INIT('h2)
	) name6951 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[2]/P0001 ,
		_w7484_
	);
	LUT3 #(
		.INIT('h80)
	) name6952 (
		_w6666_,
		_w6694_,
		_w7484_,
		_w7485_
	);
	LUT4 #(
		.INIT('hff7a)
	) name6953 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7486_
	);
	LUT2 #(
		.INIT('h2)
	) name6954 (
		_w6892_,
		_w7486_,
		_w7487_
	);
	LUT3 #(
		.INIT('h80)
	) name6955 (
		\sa11_reg[3]/P0001 ,
		_w6636_,
		_w6665_,
		_w7488_
	);
	LUT4 #(
		.INIT('h0001)
	) name6956 (
		_w6720_,
		_w7485_,
		_w7487_,
		_w7488_,
		_w7489_
	);
	LUT3 #(
		.INIT('h10)
	) name6957 (
		_w7479_,
		_w7483_,
		_w7489_,
		_w7490_
	);
	LUT3 #(
		.INIT('h10)
	) name6958 (
		_w7453_,
		_w7473_,
		_w7490_,
		_w7491_
	);
	LUT3 #(
		.INIT('h69)
	) name6959 (
		_w7224_,
		_w7433_,
		_w7491_,
		_w7492_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name6960 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7493_
	);
	LUT4 #(
		.INIT('h80aa)
	) name6961 (
		\sa22_reg[2]/P0001 ,
		_w6934_,
		_w7023_,
		_w7493_,
		_w7494_
	);
	LUT4 #(
		.INIT('h2000)
	) name6962 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7495_
	);
	LUT3 #(
		.INIT('h07)
	) name6963 (
		_w6936_,
		_w6951_,
		_w7495_,
		_w7496_
	);
	LUT2 #(
		.INIT('h1)
	) name6964 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		_w7497_
	);
	LUT2 #(
		.INIT('h8)
	) name6965 (
		_w6924_,
		_w7497_,
		_w7498_
	);
	LUT4 #(
		.INIT('haaa2)
	) name6966 (
		\sa22_reg[1]/P0001 ,
		_w7496_,
		_w7498_,
		_w7494_,
		_w7499_
	);
	LUT3 #(
		.INIT('h04)
	) name6967 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7500_
	);
	LUT3 #(
		.INIT('ha8)
	) name6968 (
		\sa22_reg[2]/P0001 ,
		_w7255_,
		_w7500_,
		_w7501_
	);
	LUT3 #(
		.INIT('h15)
	) name6969 (
		_w7008_,
		_w6951_,
		_w7497_,
		_w7502_
	);
	LUT4 #(
		.INIT('h5455)
	) name6970 (
		\sa22_reg[1]/P0001 ,
		_w7005_,
		_w7501_,
		_w7502_,
		_w7503_
	);
	LUT4 #(
		.INIT('h0040)
	) name6971 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7504_
	);
	LUT3 #(
		.INIT('h54)
	) name6972 (
		\sa22_reg[2]/P0001 ,
		_w6969_,
		_w7504_,
		_w7505_
	);
	LUT3 #(
		.INIT('h07)
	) name6973 (
		_w6943_,
		_w6945_,
		_w7229_,
		_w7506_
	);
	LUT2 #(
		.INIT('h1)
	) name6974 (
		_w7007_,
		_w6941_,
		_w7507_
	);
	LUT4 #(
		.INIT('h3111)
	) name6975 (
		\sa22_reg[2]/P0001 ,
		_w7505_,
		_w7506_,
		_w7507_,
		_w7508_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6976 (
		\sa22_reg[0]/P0001 ,
		_w7503_,
		_w7499_,
		_w7508_,
		_w7509_
	);
	LUT3 #(
		.INIT('h80)
	) name6977 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7510_
	);
	LUT3 #(
		.INIT('h7e)
	) name6978 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7511_
	);
	LUT2 #(
		.INIT('h2)
	) name6979 (
		_w6947_,
		_w7511_,
		_w7512_
	);
	LUT2 #(
		.INIT('h8)
	) name6980 (
		_w7006_,
		_w7268_,
		_w7513_
	);
	LUT3 #(
		.INIT('h2a)
	) name6981 (
		\sa22_reg[1]/P0001 ,
		_w6929_,
		_w6985_,
		_w7514_
	);
	LUT3 #(
		.INIT('h10)
	) name6982 (
		_w7512_,
		_w7513_,
		_w7514_,
		_w7515_
	);
	LUT3 #(
		.INIT('h10)
	) name6983 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7516_
	);
	LUT4 #(
		.INIT('hfa3f)
	) name6984 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7517_
	);
	LUT2 #(
		.INIT('h1)
	) name6985 (
		\sa22_reg[4]/P0001 ,
		_w7517_,
		_w7518_
	);
	LUT4 #(
		.INIT('h0200)
	) name6986 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7519_
	);
	LUT2 #(
		.INIT('h4)
	) name6987 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		_w7520_
	);
	LUT4 #(
		.INIT('h4000)
	) name6988 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7521_
	);
	LUT3 #(
		.INIT('h01)
	) name6989 (
		\sa22_reg[1]/P0001 ,
		_w7521_,
		_w7519_,
		_w7522_
	);
	LUT4 #(
		.INIT('h0777)
	) name6990 (
		\sa22_reg[4]/P0001 ,
		_w6981_,
		_w6995_,
		_w6927_,
		_w7523_
	);
	LUT3 #(
		.INIT('h40)
	) name6991 (
		_w7518_,
		_w7522_,
		_w7523_,
		_w7524_
	);
	LUT3 #(
		.INIT('h02)
	) name6992 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7525_
	);
	LUT3 #(
		.INIT('h54)
	) name6993 (
		_w6936_,
		_w7284_,
		_w7525_,
		_w7526_
	);
	LUT4 #(
		.INIT('h0015)
	) name6994 (
		\sa22_reg[2]/P0001 ,
		_w6944_,
		_w6954_,
		_w7277_,
		_w7527_
	);
	LUT4 #(
		.INIT('h0001)
	) name6995 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7528_
	);
	LUT4 #(
		.INIT('h002a)
	) name6996 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w6981_,
		_w7528_,
		_w7529_
	);
	LUT3 #(
		.INIT('h0b)
	) name6997 (
		_w7526_,
		_w7527_,
		_w7529_,
		_w7530_
	);
	LUT4 #(
		.INIT('h5501)
	) name6998 (
		\sa22_reg[0]/P0001 ,
		_w7515_,
		_w7524_,
		_w7530_,
		_w7531_
	);
	LUT4 #(
		.INIT('h0800)
	) name6999 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7532_
	);
	LUT4 #(
		.INIT('h0020)
	) name7000 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7533_
	);
	LUT4 #(
		.INIT('hf7df)
	) name7001 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7534_
	);
	LUT3 #(
		.INIT('h45)
	) name7002 (
		\sa22_reg[2]/P0001 ,
		_w7532_,
		_w7534_,
		_w7535_
	);
	LUT2 #(
		.INIT('h8)
	) name7003 (
		_w6993_,
		_w6945_,
		_w7536_
	);
	LUT4 #(
		.INIT('h0800)
	) name7004 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7537_
	);
	LUT4 #(
		.INIT('h0015)
	) name7005 (
		_w6980_,
		_w7000_,
		_w7292_,
		_w7537_,
		_w7538_
	);
	LUT4 #(
		.INIT('h5455)
	) name7006 (
		\sa22_reg[1]/P0001 ,
		_w7535_,
		_w7536_,
		_w7538_,
		_w7539_
	);
	LUT2 #(
		.INIT('h8)
	) name7007 (
		\sa22_reg[1]/P0001 ,
		\sa22_reg[2]/P0001 ,
		_w7540_
	);
	LUT3 #(
		.INIT('h01)
	) name7008 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7541_
	);
	LUT4 #(
		.INIT('hf7fa)
	) name7009 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7542_
	);
	LUT3 #(
		.INIT('h02)
	) name7010 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7543_
	);
	LUT4 #(
		.INIT('h0002)
	) name7011 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7544_
	);
	LUT4 #(
		.INIT('hcc04)
	) name7012 (
		\sa22_reg[4]/P0001 ,
		_w7540_,
		_w7542_,
		_w7544_,
		_w7545_
	);
	LUT4 #(
		.INIT('h8bcf)
	) name7013 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		_w6996_,
		_w7008_,
		_w7546_
	);
	LUT3 #(
		.INIT('h80)
	) name7014 (
		\sa22_reg[1]/P0001 ,
		_w7240_,
		_w7520_,
		_w7547_
	);
	LUT3 #(
		.INIT('h80)
	) name7015 (
		\sa22_reg[2]/P0001 ,
		_w6936_,
		_w7500_,
		_w7548_
	);
	LUT4 #(
		.INIT('h0100)
	) name7016 (
		_w7276_,
		_w7547_,
		_w7548_,
		_w7546_,
		_w7549_
	);
	LUT3 #(
		.INIT('h10)
	) name7017 (
		_w7539_,
		_w7545_,
		_w7549_,
		_w7550_
	);
	LUT3 #(
		.INIT('h10)
	) name7018 (
		_w7509_,
		_w7531_,
		_w7550_,
		_w7551_
	);
	LUT4 #(
		.INIT('h5655)
	) name7019 (
		\u0_w_reg[0][6]/P0001 ,
		_w7509_,
		_w7531_,
		_w7550_,
		_w7552_
	);
	LUT3 #(
		.INIT('hb4)
	) name7020 (
		_w7074_,
		_w7146_,
		_w7552_,
		_w7553_
	);
	LUT3 #(
		.INIT('h28)
	) name7021 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[102]/P0001 ,
		\u0_w_reg[0][6]/P0001 ,
		_w7554_
	);
	LUT4 #(
		.INIT('hff41)
	) name7022 (
		\ld_r_reg/P0001 ,
		_w7492_,
		_w7553_,
		_w7554_,
		_w7555_
	);
	LUT4 #(
		.INIT('h0001)
	) name7023 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7556_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name7024 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7557_
	);
	LUT3 #(
		.INIT('h8a)
	) name7025 (
		\sa22_reg[2]/P0001 ,
		_w7556_,
		_w7557_,
		_w7558_
	);
	LUT2 #(
		.INIT('h8)
	) name7026 (
		_w7261_,
		_w7497_,
		_w7559_
	);
	LUT3 #(
		.INIT('h8a)
	) name7027 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7560_
	);
	LUT4 #(
		.INIT('h0010)
	) name7028 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7561_
	);
	LUT3 #(
		.INIT('h0d)
	) name7029 (
		_w6921_,
		_w7560_,
		_w7561_,
		_w7562_
	);
	LUT4 #(
		.INIT('h5455)
	) name7030 (
		\sa22_reg[1]/P0001 ,
		_w7559_,
		_w7558_,
		_w7562_,
		_w7563_
	);
	LUT3 #(
		.INIT('h0e)
	) name7031 (
		_w6921_,
		_w6945_,
		_w7226_,
		_w7564_
	);
	LUT4 #(
		.INIT('h0040)
	) name7032 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7565_
	);
	LUT4 #(
		.INIT('h5155)
	) name7033 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7566_
	);
	LUT2 #(
		.INIT('h4)
	) name7034 (
		_w7565_,
		_w7566_,
		_w7567_
	);
	LUT4 #(
		.INIT('h002a)
	) name7035 (
		\sa22_reg[2]/P0001 ,
		_w6923_,
		_w6950_,
		_w7227_,
		_w7568_
	);
	LUT4 #(
		.INIT('h45cf)
	) name7036 (
		_w7496_,
		_w7564_,
		_w7567_,
		_w7568_,
		_w7569_
	);
	LUT4 #(
		.INIT('h4041)
	) name7037 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7570_
	);
	LUT3 #(
		.INIT('ha8)
	) name7038 (
		\sa22_reg[1]/P0001 ,
		_w7533_,
		_w7570_,
		_w7571_
	);
	LUT3 #(
		.INIT('h0b)
	) name7039 (
		\sa22_reg[4]/P0001 ,
		_w6941_,
		_w7233_,
		_w7572_
	);
	LUT2 #(
		.INIT('h4)
	) name7040 (
		_w7571_,
		_w7572_,
		_w7573_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7041 (
		\sa22_reg[0]/P0001 ,
		_w7563_,
		_w7569_,
		_w7573_,
		_w7574_
	);
	LUT4 #(
		.INIT('hbfef)
	) name7042 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7575_
	);
	LUT2 #(
		.INIT('h1)
	) name7043 (
		\sa22_reg[3]/P0001 ,
		_w7575_,
		_w7576_
	);
	LUT4 #(
		.INIT('h8005)
	) name7044 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7577_
	);
	LUT4 #(
		.INIT('h0100)
	) name7045 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7578_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7046 (
		\sa22_reg[1]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7579_
	);
	LUT4 #(
		.INIT('h0700)
	) name7047 (
		_w6946_,
		_w7292_,
		_w7578_,
		_w7579_,
		_w7580_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name7048 (
		_w7269_,
		_w7576_,
		_w7577_,
		_w7580_,
		_w7581_
	);
	LUT3 #(
		.INIT('hb9)
	) name7049 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7582_
	);
	LUT2 #(
		.INIT('h2)
	) name7050 (
		_w6921_,
		_w7582_,
		_w7583_
	);
	LUT3 #(
		.INIT('h40)
	) name7051 (
		\sa22_reg[1]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7584_
	);
	LUT3 #(
		.INIT('h8a)
	) name7052 (
		\sa22_reg[2]/P0001 ,
		_w7248_,
		_w7584_,
		_w7585_
	);
	LUT4 #(
		.INIT('h8000)
	) name7053 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7586_
	);
	LUT3 #(
		.INIT('h07)
	) name7054 (
		_w6923_,
		_w6950_,
		_w7586_,
		_w7587_
	);
	LUT2 #(
		.INIT('h1)
	) name7055 (
		\sa22_reg[2]/P0001 ,
		_w7528_,
		_w7588_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7056 (
		_w7583_,
		_w7585_,
		_w7587_,
		_w7588_,
		_w7589_
	);
	LUT3 #(
		.INIT('h54)
	) name7057 (
		\sa22_reg[0]/P0001 ,
		_w7581_,
		_w7589_,
		_w7590_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name7058 (
		\sa22_reg[2]/P0001 ,
		_w6943_,
		_w6941_,
		_w7500_,
		_w7591_
	);
	LUT4 #(
		.INIT('h4000)
	) name7059 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7592_
	);
	LUT4 #(
		.INIT('h8acf)
	) name7060 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		_w7007_,
		_w7592_,
		_w7593_
	);
	LUT3 #(
		.INIT('h20)
	) name7061 (
		_w7264_,
		_w7591_,
		_w7593_,
		_w7594_
	);
	LUT4 #(
		.INIT('h020a)
	) name7062 (
		\sa22_reg[2]/P0001 ,
		_w6953_,
		_w6980_,
		_w7023_,
		_w7595_
	);
	LUT3 #(
		.INIT('h15)
	) name7063 (
		\sa22_reg[2]/P0001 ,
		_w6921_,
		_w6946_,
		_w7596_
	);
	LUT3 #(
		.INIT('h04)
	) name7064 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7597_
	);
	LUT4 #(
		.INIT('hfefb)
	) name7065 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w6982_,
		_w7598_
	);
	LUT3 #(
		.INIT('h15)
	) name7066 (
		\sa22_reg[1]/P0001 ,
		_w6995_,
		_w7026_,
		_w7599_
	);
	LUT4 #(
		.INIT('hea00)
	) name7067 (
		_w7595_,
		_w7596_,
		_w7598_,
		_w7599_,
		_w7600_
	);
	LUT4 #(
		.INIT('h153f)
	) name7068 (
		\sa22_reg[6]/NET0131 ,
		_w6993_,
		_w7233_,
		_w7521_,
		_w7601_
	);
	LUT3 #(
		.INIT('he0)
	) name7069 (
		_w7594_,
		_w7600_,
		_w7601_,
		_w7602_
	);
	LUT3 #(
		.INIT('h10)
	) name7070 (
		_w7574_,
		_w7590_,
		_w7602_,
		_w7603_
	);
	LUT3 #(
		.INIT('h80)
	) name7071 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w7604_
	);
	LUT3 #(
		.INIT('ha8)
	) name7072 (
		\sa11_reg[7]/NET0131 ,
		_w7442_,
		_w7604_,
		_w7605_
	);
	LUT4 #(
		.INIT('h0007)
	) name7073 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7606_
	);
	LUT3 #(
		.INIT('h07)
	) name7074 (
		\sa11_reg[3]/P0001 ,
		_w6643_,
		_w7606_,
		_w7607_
	);
	LUT3 #(
		.INIT('h8a)
	) name7075 (
		\sa11_reg[1]/P0001 ,
		_w7605_,
		_w7607_,
		_w7608_
	);
	LUT4 #(
		.INIT('hbfef)
	) name7076 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7609_
	);
	LUT4 #(
		.INIT('haf8c)
	) name7077 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w6702_,
		_w7609_,
		_w7610_
	);
	LUT2 #(
		.INIT('h1)
	) name7078 (
		\sa11_reg[1]/P0001 ,
		_w7610_,
		_w7611_
	);
	LUT4 #(
		.INIT('h8000)
	) name7079 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7612_
	);
	LUT4 #(
		.INIT('h0007)
	) name7080 (
		_w6636_,
		_w6682_,
		_w7458_,
		_w7612_,
		_w7613_
	);
	LUT3 #(
		.INIT('hb9)
	) name7081 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7614_
	);
	LUT3 #(
		.INIT('h15)
	) name7082 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[3]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w7615_
	);
	LUT4 #(
		.INIT('h31f5)
	) name7083 (
		_w6634_,
		_w6706_,
		_w7614_,
		_w7615_,
		_w7616_
	);
	LUT3 #(
		.INIT('he4)
	) name7084 (
		\sa11_reg[2]/P0001 ,
		_w7613_,
		_w7616_,
		_w7617_
	);
	LUT4 #(
		.INIT('h5455)
	) name7085 (
		\sa11_reg[0]/P0001 ,
		_w7608_,
		_w7611_,
		_w7617_,
		_w7618_
	);
	LUT4 #(
		.INIT('h0001)
	) name7086 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7619_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name7087 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7620_
	);
	LUT3 #(
		.INIT('h8a)
	) name7088 (
		\sa11_reg[2]/P0001 ,
		_w7619_,
		_w7620_,
		_w7621_
	);
	LUT4 #(
		.INIT('h0100)
	) name7089 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7622_
	);
	LUT2 #(
		.INIT('h8)
	) name7090 (
		_w6665_,
		_w7622_,
		_w7623_
	);
	LUT3 #(
		.INIT('h8a)
	) name7091 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7624_
	);
	LUT3 #(
		.INIT('h31)
	) name7092 (
		_w6634_,
		_w6687_,
		_w7624_,
		_w7625_
	);
	LUT4 #(
		.INIT('h5455)
	) name7093 (
		\sa11_reg[1]/P0001 ,
		_w7623_,
		_w7621_,
		_w7625_,
		_w7626_
	);
	LUT4 #(
		.INIT('h0001)
	) name7094 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7627_
	);
	LUT3 #(
		.INIT('h40)
	) name7095 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w7628_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7096 (
		\sa11_reg[1]/P0001 ,
		_w7474_,
		_w7628_,
		_w7627_,
		_w7629_
	);
	LUT2 #(
		.INIT('h1)
	) name7097 (
		_w6638_,
		_w7444_,
		_w7630_
	);
	LUT3 #(
		.INIT('h2a)
	) name7098 (
		\sa11_reg[2]/P0001 ,
		_w6857_,
		_w7630_,
		_w7631_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name7099 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7632_
	);
	LUT4 #(
		.INIT('h0301)
	) name7100 (
		\sa11_reg[3]/P0001 ,
		_w6848_,
		_w7455_,
		_w7632_,
		_w7633_
	);
	LUT3 #(
		.INIT('h13)
	) name7101 (
		_w6634_,
		_w6648_,
		_w6691_,
		_w7634_
	);
	LUT3 #(
		.INIT('he0)
	) name7102 (
		\sa11_reg[2]/P0001 ,
		_w7633_,
		_w7634_,
		_w7635_
	);
	LUT4 #(
		.INIT('h0100)
	) name7103 (
		_w7631_,
		_w7629_,
		_w7626_,
		_w7635_,
		_w7636_
	);
	LUT4 #(
		.INIT('h4000)
	) name7104 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w7637_
	);
	LUT2 #(
		.INIT('h4)
	) name7105 (
		\sa11_reg[2]/P0001 ,
		_w7637_,
		_w7638_
	);
	LUT4 #(
		.INIT('h8daf)
	) name7106 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6719_,
		_w6694_,
		_w7639_
	);
	LUT2 #(
		.INIT('h8)
	) name7107 (
		_w6730_,
		_w6691_,
		_w7640_
	);
	LUT4 #(
		.INIT('h0777)
	) name7108 (
		_w6730_,
		_w6691_,
		_w6861_,
		_w6902_,
		_w7641_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name7109 (
		\sa11_reg[1]/P0001 ,
		_w7638_,
		_w7639_,
		_w7641_,
		_w7642_
	);
	LUT4 #(
		.INIT('hff4b)
	) name7110 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7643_
	);
	LUT2 #(
		.INIT('h2)
	) name7111 (
		_w7441_,
		_w7643_,
		_w7644_
	);
	LUT4 #(
		.INIT('h0040)
	) name7112 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w7645_
	);
	LUT2 #(
		.INIT('h8)
	) name7113 (
		_w6712_,
		_w7645_,
		_w7646_
	);
	LUT4 #(
		.INIT('h5554)
	) name7114 (
		\sa11_reg[1]/P0001 ,
		_w6916_,
		_w7646_,
		_w7644_,
		_w7647_
	);
	LUT2 #(
		.INIT('h8)
	) name7115 (
		\sa11_reg[6]/NET0131 ,
		_w7464_,
		_w7648_
	);
	LUT3 #(
		.INIT('h8a)
	) name7116 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w6870_,
		_w7649_
	);
	LUT3 #(
		.INIT('h02)
	) name7117 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w7650_
	);
	LUT3 #(
		.INIT('h67)
	) name7118 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7651_
	);
	LUT2 #(
		.INIT('h2)
	) name7119 (
		_w7650_,
		_w7651_,
		_w7652_
	);
	LUT3 #(
		.INIT('h45)
	) name7120 (
		_w7648_,
		_w7649_,
		_w7652_,
		_w7653_
	);
	LUT3 #(
		.INIT('h10)
	) name7121 (
		_w7647_,
		_w7642_,
		_w7653_,
		_w7654_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7122 (
		\sa11_reg[0]/P0001 ,
		_w7636_,
		_w7618_,
		_w7654_,
		_w7655_
	);
	LUT2 #(
		.INIT('h9)
	) name7123 (
		_w7603_,
		_w7655_,
		_w7656_
	);
	LUT4 #(
		.INIT('hcfca)
	) name7124 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7657_
	);
	LUT3 #(
		.INIT('h08)
	) name7125 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7658_
	);
	LUT3 #(
		.INIT('h02)
	) name7126 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w7659_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7127 (
		\sa11_reg[2]/P0001 ,
		_w7658_,
		_w7659_,
		_w7657_,
		_w7660_
	);
	LUT4 #(
		.INIT('h0777)
	) name7128 (
		_w6641_,
		_w6671_,
		_w6690_,
		_w7442_,
		_w7661_
	);
	LUT3 #(
		.INIT('h8a)
	) name7129 (
		\sa11_reg[1]/P0001 ,
		_w7660_,
		_w7661_,
		_w7662_
	);
	LUT3 #(
		.INIT('h54)
	) name7130 (
		\sa11_reg[7]/NET0131 ,
		_w7457_,
		_w7628_,
		_w7663_
	);
	LUT4 #(
		.INIT('h0010)
	) name7131 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7664_
	);
	LUT2 #(
		.INIT('h1)
	) name7132 (
		_w6678_,
		_w7664_,
		_w7665_
	);
	LUT4 #(
		.INIT('h4404)
	) name7133 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w7666_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name7134 (
		_w6637_,
		_w6664_,
		_w7650_,
		_w7666_,
		_w7667_
	);
	LUT4 #(
		.INIT('h4555)
	) name7135 (
		\sa11_reg[1]/P0001 ,
		_w7663_,
		_w7665_,
		_w7667_,
		_w7668_
	);
	LUT4 #(
		.INIT('hecfd)
	) name7136 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w7669_
	);
	LUT4 #(
		.INIT('h0301)
	) name7137 (
		\sa11_reg[6]/NET0131 ,
		_w6876_,
		_w6880_,
		_w7669_,
		_w7670_
	);
	LUT3 #(
		.INIT('h07)
	) name7138 (
		_w7437_,
		_w7441_,
		_w7455_,
		_w7671_
	);
	LUT3 #(
		.INIT('hd0)
	) name7139 (
		\sa11_reg[2]/P0001 ,
		_w7670_,
		_w7671_,
		_w7672_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7140 (
		\sa11_reg[0]/P0001 ,
		_w7668_,
		_w7662_,
		_w7672_,
		_w7673_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name7141 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7674_
	);
	LUT2 #(
		.INIT('h2)
	) name7142 (
		_w6845_,
		_w7674_,
		_w7675_
	);
	LUT4 #(
		.INIT('hadfb)
	) name7143 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7676_
	);
	LUT4 #(
		.INIT('h0302)
	) name7144 (
		\sa11_reg[3]/P0001 ,
		_w6672_,
		_w6896_,
		_w7676_,
		_w7677_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7145 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[2]/P0001 ,
		_w7675_,
		_w7677_,
		_w7678_
	);
	LUT2 #(
		.INIT('h8)
	) name7146 (
		_w6641_,
		_w6730_,
		_w7679_
	);
	LUT3 #(
		.INIT('h10)
	) name7147 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w7680_
	);
	LUT4 #(
		.INIT('h0001)
	) name7148 (
		\sa11_reg[1]/P0001 ,
		_w6655_,
		_w7444_,
		_w7680_,
		_w7681_
	);
	LUT4 #(
		.INIT('h0020)
	) name7149 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7682_
	);
	LUT4 #(
		.INIT('hf5e4)
	) name7150 (
		\sa11_reg[2]/P0001 ,
		_w6701_,
		_w6683_,
		_w7682_,
		_w7683_
	);
	LUT4 #(
		.INIT('h0800)
	) name7151 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7684_
	);
	LUT4 #(
		.INIT('h002a)
	) name7152 (
		\sa11_reg[1]/P0001 ,
		_w6637_,
		_w7457_,
		_w7684_,
		_w7685_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name7153 (
		_w7679_,
		_w7681_,
		_w7683_,
		_w7685_,
		_w7686_
	);
	LUT4 #(
		.INIT('h8808)
	) name7154 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7687_
	);
	LUT2 #(
		.INIT('h8)
	) name7155 (
		_w7624_,
		_w7687_,
		_w7688_
	);
	LUT3 #(
		.INIT('h2a)
	) name7156 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w6898_,
		_w7689_
	);
	LUT3 #(
		.INIT('h15)
	) name7157 (
		\sa11_reg[2]/P0001 ,
		_w6642_,
		_w6644_,
		_w7690_
	);
	LUT4 #(
		.INIT('h4000)
	) name7158 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w7691_
	);
	LUT3 #(
		.INIT('h01)
	) name7159 (
		_w6687_,
		_w7481_,
		_w7691_,
		_w7692_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7160 (
		_w7688_,
		_w7689_,
		_w7690_,
		_w7692_,
		_w7693_
	);
	LUT3 #(
		.INIT('h54)
	) name7161 (
		\sa11_reg[0]/P0001 ,
		_w7686_,
		_w7693_,
		_w7694_
	);
	LUT4 #(
		.INIT('hbdff)
	) name7162 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w7695_
	);
	LUT3 #(
		.INIT('h10)
	) name7163 (
		_w6687_,
		_w7691_,
		_w7695_,
		_w7696_
	);
	LUT2 #(
		.INIT('h2)
	) name7164 (
		\sa11_reg[2]/P0001 ,
		_w7637_,
		_w7697_
	);
	LUT3 #(
		.INIT('h51)
	) name7165 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[2]/P0001 ,
		_w7637_,
		_w7698_
	);
	LUT2 #(
		.INIT('h4)
	) name7166 (
		_w7696_,
		_w7698_,
		_w7699_
	);
	LUT4 #(
		.INIT('h8caf)
	) name7167 (
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6659_,
		_w6870_,
		_w7700_
	);
	LUT2 #(
		.INIT('h4)
	) name7168 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[2]/P0001 ,
		_w7701_
	);
	LUT4 #(
		.INIT('h4000)
	) name7169 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w7702_
	);
	LUT4 #(
		.INIT('h0007)
	) name7170 (
		_w6641_,
		_w6671_,
		_w6868_,
		_w7702_,
		_w7703_
	);
	LUT4 #(
		.INIT('hfcb8)
	) name7171 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[2]/P0001 ,
		_w7700_,
		_w7703_,
		_w7704_
	);
	LUT2 #(
		.INIT('h4)
	) name7172 (
		_w7699_,
		_w7704_,
		_w7705_
	);
	LUT4 #(
		.INIT('h0100)
	) name7173 (
		_w7673_,
		_w7694_,
		_w7678_,
		_w7705_,
		_w7706_
	);
	LUT3 #(
		.INIT('h07)
	) name7174 (
		_w6748_,
		_w6788_,
		_w7175_,
		_w7707_
	);
	LUT3 #(
		.INIT('h80)
	) name7175 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7708_
	);
	LUT4 #(
		.INIT('hcedf)
	) name7176 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7709_
	);
	LUT3 #(
		.INIT('h8a)
	) name7177 (
		\sa00_reg[2]/P0001 ,
		_w7708_,
		_w7709_,
		_w7710_
	);
	LUT3 #(
		.INIT('ha2)
	) name7178 (
		\sa00_reg[1]/P0001 ,
		_w7707_,
		_w7710_,
		_w7711_
	);
	LUT4 #(
		.INIT('h0040)
	) name7179 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7712_
	);
	LUT4 #(
		.INIT('h0008)
	) name7180 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7713_
	);
	LUT4 #(
		.INIT('h0001)
	) name7181 (
		_w6839_,
		_w7414_,
		_w7712_,
		_w7713_,
		_w7714_
	);
	LUT2 #(
		.INIT('h1)
	) name7182 (
		\sa00_reg[2]/P0001 ,
		_w7714_,
		_w7715_
	);
	LUT4 #(
		.INIT('hb8bb)
	) name7183 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w7716_
	);
	LUT2 #(
		.INIT('h2)
	) name7184 (
		_w6739_,
		_w7716_,
		_w7717_
	);
	LUT4 #(
		.INIT('h0888)
	) name7185 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7718_
	);
	LUT3 #(
		.INIT('h23)
	) name7186 (
		_w6837_,
		_w6839_,
		_w7718_,
		_w7719_
	);
	LUT3 #(
		.INIT('h45)
	) name7187 (
		\sa00_reg[1]/P0001 ,
		_w7717_,
		_w7719_,
		_w7720_
	);
	LUT2 #(
		.INIT('h8)
	) name7188 (
		\sa00_reg[2]/P0001 ,
		_w6771_,
		_w7721_
	);
	LUT4 #(
		.INIT('hbdff)
	) name7189 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w6745_,
		_w7722_
	);
	LUT2 #(
		.INIT('h4)
	) name7190 (
		_w7721_,
		_w7722_,
		_w7723_
	);
	LUT4 #(
		.INIT('h0100)
	) name7191 (
		_w7711_,
		_w7720_,
		_w7715_,
		_w7723_,
		_w7724_
	);
	LUT2 #(
		.INIT('h2)
	) name7192 (
		\sa00_reg[0]/P0001 ,
		_w7724_,
		_w7725_
	);
	LUT4 #(
		.INIT('h5510)
	) name7193 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w6771_,
		_w7415_,
		_w7726_
	);
	LUT4 #(
		.INIT('h0020)
	) name7194 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7727_
	);
	LUT4 #(
		.INIT('h13df)
	) name7195 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w6788_,
		_w7727_,
		_w7728_
	);
	LUT3 #(
		.INIT('h45)
	) name7196 (
		\sa00_reg[1]/P0001 ,
		_w7726_,
		_w7728_,
		_w7729_
	);
	LUT4 #(
		.INIT('h0800)
	) name7197 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w7730_
	);
	LUT4 #(
		.INIT('h5554)
	) name7198 (
		\sa00_reg[2]/P0001 ,
		_w7179_,
		_w7405_,
		_w7730_,
		_w7731_
	);
	LUT3 #(
		.INIT('h01)
	) name7199 (
		_w6819_,
		_w6777_,
		_w7160_,
		_w7732_
	);
	LUT3 #(
		.INIT('h8a)
	) name7200 (
		\sa00_reg[1]/P0001 ,
		_w7731_,
		_w7732_,
		_w7733_
	);
	LUT4 #(
		.INIT('h00bf)
	) name7201 (
		\sa00_reg[7]/NET0131 ,
		_w6750_,
		_w7191_,
		_w7214_,
		_w7734_
	);
	LUT4 #(
		.INIT('hffa8)
	) name7202 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7735_
	);
	LUT4 #(
		.INIT('hdbff)
	) name7203 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7736_
	);
	LUT4 #(
		.INIT('hf351)
	) name7204 (
		_w6805_,
		_w6832_,
		_w7735_,
		_w7736_,
		_w7737_
	);
	LUT2 #(
		.INIT('h8)
	) name7205 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[2]/P0001 ,
		_w7738_
	);
	LUT4 #(
		.INIT('h4000)
	) name7206 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7739_
	);
	LUT3 #(
		.INIT('hc8)
	) name7207 (
		_w7169_,
		_w7738_,
		_w7739_,
		_w7740_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name7208 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7741_
	);
	LUT2 #(
		.INIT('h2)
	) name7209 (
		_w7389_,
		_w7741_,
		_w7742_
	);
	LUT4 #(
		.INIT('h1000)
	) name7210 (
		_w7740_,
		_w7742_,
		_w7734_,
		_w7737_,
		_w7743_
	);
	LUT4 #(
		.INIT('h5455)
	) name7211 (
		\sa00_reg[0]/P0001 ,
		_w7733_,
		_w7729_,
		_w7743_,
		_w7744_
	);
	LUT4 #(
		.INIT('h0100)
	) name7212 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7745_
	);
	LUT4 #(
		.INIT('h002a)
	) name7213 (
		\sa00_reg[2]/P0001 ,
		_w6745_,
		_w6788_,
		_w7214_,
		_w7746_
	);
	LUT2 #(
		.INIT('h1)
	) name7214 (
		\sa00_reg[2]/P0001 ,
		_w7727_,
		_w7747_
	);
	LUT3 #(
		.INIT('h07)
	) name7215 (
		_w6745_,
		_w6759_,
		_w7381_,
		_w7748_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7216 (
		_w7745_,
		_w7746_,
		_w7747_,
		_w7748_,
		_w7749_
	);
	LUT4 #(
		.INIT('h0777)
	) name7217 (
		_w6780_,
		_w6781_,
		_w6776_,
		_w7191_,
		_w7750_
	);
	LUT3 #(
		.INIT('h45)
	) name7218 (
		\sa00_reg[1]/P0001 ,
		_w7749_,
		_w7750_,
		_w7751_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name7219 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w7752_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7220 (
		\sa00_reg[3]/P0001 ,
		_w6744_,
		_w7399_,
		_w7752_,
		_w7753_
	);
	LUT2 #(
		.INIT('h2)
	) name7221 (
		_w7738_,
		_w7753_,
		_w7754_
	);
	LUT3 #(
		.INIT('h80)
	) name7222 (
		\sa00_reg[2]/P0001 ,
		_w6780_,
		_w6781_,
		_w7755_
	);
	LUT4 #(
		.INIT('h007f)
	) name7223 (
		\sa00_reg[2]/P0001 ,
		_w6780_,
		_w6781_,
		_w7180_,
		_w7756_
	);
	LUT3 #(
		.INIT('h04)
	) name7224 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w7757_
	);
	LUT4 #(
		.INIT('h0203)
	) name7225 (
		_w6780_,
		_w7160_,
		_w7385_,
		_w7757_,
		_w7758_
	);
	LUT4 #(
		.INIT('h0ece)
	) name7226 (
		_w6831_,
		_w7200_,
		_w7756_,
		_w7758_,
		_w7759_
	);
	LUT2 #(
		.INIT('h1)
	) name7227 (
		_w7754_,
		_w7759_,
		_w7760_
	);
	LUT3 #(
		.INIT('h10)
	) name7228 (
		_w7744_,
		_w7751_,
		_w7760_,
		_w7761_
	);
	LUT3 #(
		.INIT('h65)
	) name7229 (
		_w7706_,
		_w7725_,
		_w7761_,
		_w7762_
	);
	LUT3 #(
		.INIT('h23)
	) name7230 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7763_
	);
	LUT3 #(
		.INIT('h4c)
	) name7231 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7764_
	);
	LUT4 #(
		.INIT('h0803)
	) name7232 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7765_
	);
	LUT3 #(
		.INIT('h54)
	) name7233 (
		\sa33_reg[2]/P0001 ,
		_w7105_,
		_w7765_,
		_w7766_
	);
	LUT3 #(
		.INIT('h80)
	) name7234 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7767_
	);
	LUT4 #(
		.INIT('h4000)
	) name7235 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7768_
	);
	LUT3 #(
		.INIT('ha8)
	) name7236 (
		\sa33_reg[2]/P0001 ,
		_w7767_,
		_w7768_,
		_w7769_
	);
	LUT3 #(
		.INIT('h45)
	) name7237 (
		_w7092_,
		_w7039_,
		_w7040_,
		_w7770_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7238 (
		\sa33_reg[1]/P0001 ,
		_w7769_,
		_w7766_,
		_w7770_,
		_w7771_
	);
	LUT4 #(
		.INIT('h0020)
	) name7239 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7772_
	);
	LUT4 #(
		.INIT('h5540)
	) name7240 (
		\sa33_reg[2]/P0001 ,
		_w7069_,
		_w7123_,
		_w7772_,
		_w7773_
	);
	LUT4 #(
		.INIT('h153f)
	) name7241 (
		_w7055_,
		_w7033_,
		_w7110_,
		_w7056_,
		_w7774_
	);
	LUT4 #(
		.INIT('h135f)
	) name7242 (
		_w7086_,
		_w7114_,
		_w7138_,
		_w7339_,
		_w7775_
	);
	LUT4 #(
		.INIT('h4555)
	) name7243 (
		\sa33_reg[1]/P0001 ,
		_w7773_,
		_w7774_,
		_w7775_,
		_w7776_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name7244 (
		\sa33_reg[6]/P0001 ,
		_w7033_,
		_w7110_,
		_w7059_,
		_w7777_
	);
	LUT4 #(
		.INIT('hffa8)
	) name7245 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7778_
	);
	LUT2 #(
		.INIT('h2)
	) name7246 (
		_w7055_,
		_w7778_,
		_w7779_
	);
	LUT4 #(
		.INIT('h1333)
	) name7247 (
		\sa33_reg[4]/P0001 ,
		_w7131_,
		_w7138_,
		_w7139_,
		_w7780_
	);
	LUT4 #(
		.INIT('h3200)
	) name7248 (
		\sa33_reg[2]/P0001 ,
		_w7779_,
		_w7777_,
		_w7780_,
		_w7781_
	);
	LUT4 #(
		.INIT('h5455)
	) name7249 (
		\sa33_reg[0]/P0001 ,
		_w7771_,
		_w7776_,
		_w7781_,
		_w7782_
	);
	LUT3 #(
		.INIT('h20)
	) name7250 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7783_
	);
	LUT4 #(
		.INIT('h54fc)
	) name7251 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7784_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7252 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7783_,
		_w7784_,
		_w7785_
	);
	LUT4 #(
		.INIT('h8000)
	) name7253 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7786_
	);
	LUT3 #(
		.INIT('h13)
	) name7254 (
		\sa33_reg[4]/P0001 ,
		_w7116_,
		_w7786_,
		_w7787_
	);
	LUT3 #(
		.INIT('h8a)
	) name7255 (
		\sa33_reg[1]/P0001 ,
		_w7785_,
		_w7787_,
		_w7788_
	);
	LUT2 #(
		.INIT('h8)
	) name7256 (
		_w7087_,
		_w7105_,
		_w7789_
	);
	LUT4 #(
		.INIT('h0031)
	) name7257 (
		_w7080_,
		_w7063_,
		_w7335_,
		_w7364_,
		_w7790_
	);
	LUT3 #(
		.INIT('h45)
	) name7258 (
		\sa33_reg[1]/P0001 ,
		_w7789_,
		_w7790_,
		_w7791_
	);
	LUT4 #(
		.INIT('h0008)
	) name7259 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7792_
	);
	LUT4 #(
		.INIT('h0800)
	) name7260 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7793_
	);
	LUT4 #(
		.INIT('h0001)
	) name7261 (
		_w7364_,
		_w7313_,
		_w7792_,
		_w7793_,
		_w7794_
	);
	LUT4 #(
		.INIT('h7707)
	) name7262 (
		_w7049_,
		_w7139_,
		_w7141_,
		_w7344_,
		_w7795_
	);
	LUT3 #(
		.INIT('he0)
	) name7263 (
		\sa33_reg[2]/P0001 ,
		_w7794_,
		_w7795_,
		_w7796_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7264 (
		\sa33_reg[0]/P0001 ,
		_w7788_,
		_w7791_,
		_w7796_,
		_w7797_
	);
	LUT4 #(
		.INIT('h2000)
	) name7265 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7798_
	);
	LUT4 #(
		.INIT('h0020)
	) name7266 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7799_
	);
	LUT4 #(
		.INIT('h0007)
	) name7267 (
		_w7049_,
		_w7062_,
		_w7799_,
		_w7798_,
		_w7800_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name7268 (
		\sa33_reg[6]/P0001 ,
		_w7080_,
		_w7039_,
		_w7063_,
		_w7801_
	);
	LUT4 #(
		.INIT('h0155)
	) name7269 (
		\sa33_reg[1]/P0001 ,
		\sa33_reg[2]/P0001 ,
		_w7800_,
		_w7801_,
		_w7802_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name7270 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7803_
	);
	LUT2 #(
		.INIT('h2)
	) name7271 (
		\sa33_reg[3]/P0001 ,
		_w7803_,
		_w7804_
	);
	LUT3 #(
		.INIT('h2a)
	) name7272 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7141_,
		_w7805_
	);
	LUT2 #(
		.INIT('h4)
	) name7273 (
		_w7804_,
		_w7805_,
		_w7806_
	);
	LUT2 #(
		.INIT('h4)
	) name7274 (
		_w7049_,
		_w7062_,
		_w7807_
	);
	LUT4 #(
		.INIT('h1101)
	) name7275 (
		\sa33_reg[2]/P0001 ,
		_w7088_,
		_w7078_,
		_w7035_,
		_w7808_
	);
	LUT3 #(
		.INIT('h8a)
	) name7276 (
		\sa33_reg[1]/P0001 ,
		_w7807_,
		_w7808_,
		_w7809_
	);
	LUT2 #(
		.INIT('h4)
	) name7277 (
		\sa33_reg[1]/P0001 ,
		\sa33_reg[2]/P0001 ,
		_w7810_
	);
	LUT4 #(
		.INIT('hfcfa)
	) name7278 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7811_
	);
	LUT4 #(
		.INIT('h3f2a)
	) name7279 (
		\sa33_reg[3]/P0001 ,
		_w7048_,
		_w7050_,
		_w7811_,
		_w7812_
	);
	LUT3 #(
		.INIT('h80)
	) name7280 (
		\sa33_reg[4]/P0001 ,
		_w7126_,
		_w7138_,
		_w7813_
	);
	LUT3 #(
		.INIT('h40)
	) name7281 (
		\sa33_reg[7]/NET0131 ,
		_w7107_,
		_w7108_,
		_w7814_
	);
	LUT4 #(
		.INIT('h0051)
	) name7282 (
		_w7813_,
		_w7810_,
		_w7812_,
		_w7814_,
		_w7815_
	);
	LUT4 #(
		.INIT('h4500)
	) name7283 (
		_w7802_,
		_w7806_,
		_w7809_,
		_w7815_,
		_w7816_
	);
	LUT3 #(
		.INIT('h10)
	) name7284 (
		_w7797_,
		_w7782_,
		_w7816_,
		_w7817_
	);
	LUT4 #(
		.INIT('h5540)
	) name7285 (
		\sa22_reg[2]/P0001 ,
		_w6934_,
		_w7023_,
		_w7533_,
		_w7818_
	);
	LUT2 #(
		.INIT('h4)
	) name7286 (
		\sa22_reg[3]/P0001 ,
		_w7230_,
		_w7819_
	);
	LUT3 #(
		.INIT('h15)
	) name7287 (
		\sa22_reg[1]/P0001 ,
		_w6982_,
		_w7249_,
		_w7820_
	);
	LUT4 #(
		.INIT('h135f)
	) name7288 (
		\sa22_reg[2]/P0001 ,
		_w6936_,
		_w7277_,
		_w7500_,
		_w7821_
	);
	LUT4 #(
		.INIT('h1000)
	) name7289 (
		_w7819_,
		_w7818_,
		_w7820_,
		_w7821_,
		_w7822_
	);
	LUT4 #(
		.INIT('h4000)
	) name7290 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7823_
	);
	LUT3 #(
		.INIT('ha8)
	) name7291 (
		\sa22_reg[2]/P0001 ,
		_w7510_,
		_w7823_,
		_w7824_
	);
	LUT4 #(
		.INIT('h0800)
	) name7292 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7825_
	);
	LUT4 #(
		.INIT('h5554)
	) name7293 (
		\sa22_reg[2]/P0001 ,
		_w7006_,
		_w7516_,
		_w7825_,
		_w7826_
	);
	LUT4 #(
		.INIT('h0002)
	) name7294 (
		\sa22_reg[1]/P0001 ,
		_w6978_,
		_w6928_,
		_w6930_,
		_w7827_
	);
	LUT3 #(
		.INIT('h10)
	) name7295 (
		_w7826_,
		_w7824_,
		_w7827_,
		_w7828_
	);
	LUT3 #(
		.INIT('h07)
	) name7296 (
		_w6923_,
		_w6950_,
		_w7015_,
		_w7829_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7297 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7830_
	);
	LUT2 #(
		.INIT('h4)
	) name7298 (
		_w7556_,
		_w7830_,
		_w7831_
	);
	LUT4 #(
		.INIT('h5540)
	) name7299 (
		_w7027_,
		_w7250_,
		_w7829_,
		_w7831_,
		_w7832_
	);
	LUT4 #(
		.INIT('h0155)
	) name7300 (
		\sa22_reg[0]/P0001 ,
		_w7822_,
		_w7828_,
		_w7832_,
		_w7833_
	);
	LUT3 #(
		.INIT('h32)
	) name7301 (
		_w7007_,
		_w6923_,
		_w6950_,
		_w7834_
	);
	LUT2 #(
		.INIT('h1)
	) name7302 (
		_w6978_,
		_w7504_,
		_w7835_
	);
	LUT3 #(
		.INIT('h45)
	) name7303 (
		\sa22_reg[2]/P0001 ,
		_w7834_,
		_w7835_,
		_w7836_
	);
	LUT2 #(
		.INIT('h8)
	) name7304 (
		\sa22_reg[6]/NET0131 ,
		_w6986_,
		_w7837_
	);
	LUT3 #(
		.INIT('h07)
	) name7305 (
		\sa22_reg[6]/NET0131 ,
		_w6986_,
		_w7003_,
		_w7838_
	);
	LUT3 #(
		.INIT('h20)
	) name7306 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7839_
	);
	LUT3 #(
		.INIT('h10)
	) name7307 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7840_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7308 (
		\sa22_reg[2]/P0001 ,
		_w7249_,
		_w7840_,
		_w7839_,
		_w7841_
	);
	LUT3 #(
		.INIT('ha2)
	) name7309 (
		\sa22_reg[0]/P0001 ,
		_w7838_,
		_w7841_,
		_w7842_
	);
	LUT3 #(
		.INIT('ha8)
	) name7310 (
		\sa22_reg[1]/P0001 ,
		_w7836_,
		_w7842_,
		_w7843_
	);
	LUT2 #(
		.INIT('h2)
	) name7311 (
		_w6987_,
		_w6993_,
		_w7844_
	);
	LUT3 #(
		.INIT('h13)
	) name7312 (
		_w6967_,
		_w7026_,
		_w7225_,
		_w7845_
	);
	LUT3 #(
		.INIT('h45)
	) name7313 (
		\sa22_reg[1]/P0001 ,
		_w7844_,
		_w7845_,
		_w7846_
	);
	LUT4 #(
		.INIT('h0008)
	) name7314 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7847_
	);
	LUT4 #(
		.INIT('hf7bf)
	) name7315 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7848_
	);
	LUT3 #(
		.INIT('h45)
	) name7316 (
		\sa22_reg[2]/P0001 ,
		_w7847_,
		_w7848_,
		_w7849_
	);
	LUT2 #(
		.INIT('h8)
	) name7317 (
		\sa22_reg[4]/P0001 ,
		_w7256_,
		_w7850_
	);
	LUT4 #(
		.INIT('hf531)
	) name7318 (
		_w6981_,
		_w6963_,
		_w7272_,
		_w7540_,
		_w7851_
	);
	LUT3 #(
		.INIT('h10)
	) name7319 (
		_w7850_,
		_w7849_,
		_w7851_,
		_w7852_
	);
	LUT3 #(
		.INIT('h8a)
	) name7320 (
		\sa22_reg[0]/P0001 ,
		_w7846_,
		_w7852_,
		_w7853_
	);
	LUT4 #(
		.INIT('h0007)
	) name7321 (
		_w6953_,
		_w6954_,
		_w7291_,
		_w7495_,
		_w7854_
	);
	LUT4 #(
		.INIT('h153f)
	) name7322 (
		_w6953_,
		_w6936_,
		_w6951_,
		_w7255_,
		_w7855_
	);
	LUT4 #(
		.INIT('h0155)
	) name7323 (
		\sa22_reg[1]/P0001 ,
		\sa22_reg[2]/P0001 ,
		_w7854_,
		_w7855_,
		_w7856_
	);
	LUT2 #(
		.INIT('h4)
	) name7324 (
		\sa22_reg[1]/P0001 ,
		\sa22_reg[2]/P0001 ,
		_w7857_
	);
	LUT4 #(
		.INIT('h0013)
	) name7325 (
		_w6943_,
		_w6991_,
		_w6945_,
		_w7015_,
		_w7858_
	);
	LUT2 #(
		.INIT('h2)
	) name7326 (
		_w7857_,
		_w7858_,
		_w7859_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name7327 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7860_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7328 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w6981_,
		_w7860_,
		_w7861_
	);
	LUT4 #(
		.INIT('h153f)
	) name7329 (
		_w6953_,
		_w6940_,
		_w7019_,
		_w7255_,
		_w7862_
	);
	LUT4 #(
		.INIT('hf733)
	) name7330 (
		\sa22_reg[1]/P0001 ,
		\sa22_reg[2]/P0001 ,
		_w7861_,
		_w7862_,
		_w7863_
	);
	LUT3 #(
		.INIT('h10)
	) name7331 (
		_w7859_,
		_w7856_,
		_w7863_,
		_w7864_
	);
	LUT4 #(
		.INIT('h0100)
	) name7332 (
		_w7833_,
		_w7853_,
		_w7843_,
		_w7864_,
		_w7865_
	);
	LUT4 #(
		.INIT('hcf4f)
	) name7333 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7866_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7334 (
		\sa22_reg[2]/P0001 ,
		_w7525_,
		_w7541_,
		_w7866_,
		_w7867_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7335 (
		\sa22_reg[2]/P0001 ,
		_w6991_,
		_w6923_,
		_w7287_,
		_w7868_
	);
	LUT3 #(
		.INIT('h8a)
	) name7336 (
		\sa22_reg[1]/P0001 ,
		_w7867_,
		_w7868_,
		_w7869_
	);
	LUT4 #(
		.INIT('h7d1d)
	) name7337 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7870_
	);
	LUT2 #(
		.INIT('h1)
	) name7338 (
		\sa22_reg[2]/P0001 ,
		_w7870_,
		_w7871_
	);
	LUT2 #(
		.INIT('h4)
	) name7339 (
		_w6993_,
		_w7597_,
		_w7872_
	);
	LUT3 #(
		.INIT('h13)
	) name7340 (
		_w6947_,
		_w7253_,
		_w7840_,
		_w7873_
	);
	LUT4 #(
		.INIT('h5455)
	) name7341 (
		\sa22_reg[1]/P0001 ,
		_w7871_,
		_w7872_,
		_w7873_,
		_w7874_
	);
	LUT4 #(
		.INIT('h1000)
	) name7342 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7875_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name7343 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7876_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7344 (
		\sa22_reg[2]/P0001 ,
		_w6972_,
		_w7875_,
		_w7876_,
		_w7877_
	);
	LUT3 #(
		.INIT('h07)
	) name7345 (
		_w6971_,
		_w7497_,
		_w7565_,
		_w7878_
	);
	LUT2 #(
		.INIT('h4)
	) name7346 (
		_w7877_,
		_w7878_,
		_w7879_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7347 (
		\sa22_reg[0]/P0001 ,
		_w7874_,
		_w7869_,
		_w7879_,
		_w7880_
	);
	LUT3 #(
		.INIT('h54)
	) name7348 (
		\sa22_reg[2]/P0001 ,
		_w6937_,
		_w7291_,
		_w7881_
	);
	LUT4 #(
		.INIT('h0400)
	) name7349 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7882_
	);
	LUT4 #(
		.INIT('h080a)
	) name7350 (
		\sa22_reg[1]/P0001 ,
		_w7268_,
		_w7532_,
		_w7882_,
		_w7883_
	);
	LUT2 #(
		.INIT('h8)
	) name7351 (
		_w6958_,
		_w7292_,
		_w7884_
	);
	LUT3 #(
		.INIT('h10)
	) name7352 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w7885_
	);
	LUT4 #(
		.INIT('h0001)
	) name7353 (
		\sa22_reg[1]/P0001 ,
		_w6996_,
		_w7495_,
		_w7885_,
		_w7886_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name7354 (
		_w7881_,
		_w7883_,
		_w7884_,
		_w7886_,
		_w7887_
	);
	LUT4 #(
		.INIT('h7ff7)
	) name7355 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7888_
	);
	LUT4 #(
		.INIT('hdf55)
	) name7356 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7019_,
		_w7888_,
		_w7889_
	);
	LUT2 #(
		.INIT('h1)
	) name7357 (
		_w7561_,
		_w7823_,
		_w7890_
	);
	LUT3 #(
		.INIT('h07)
	) name7358 (
		_w6929_,
		_w6985_,
		_w7544_,
		_w7891_
	);
	LUT4 #(
		.INIT('hd888)
	) name7359 (
		\sa22_reg[2]/P0001 ,
		_w7889_,
		_w7890_,
		_w7891_,
		_w7892_
	);
	LUT3 #(
		.INIT('h45)
	) name7360 (
		\sa22_reg[0]/P0001 ,
		_w7887_,
		_w7892_,
		_w7893_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name7361 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7894_
	);
	LUT2 #(
		.INIT('h2)
	) name7362 (
		_w7520_,
		_w7894_,
		_w7895_
	);
	LUT4 #(
		.INIT('hadfb)
	) name7363 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w7896_
	);
	LUT4 #(
		.INIT('h0302)
	) name7364 (
		\sa22_reg[3]/P0001 ,
		_w7003_,
		_w6928_,
		_w7896_,
		_w7897_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7365 (
		\sa22_reg[1]/P0001 ,
		\sa22_reg[2]/P0001 ,
		_w7895_,
		_w7897_,
		_w7898_
	);
	LUT4 #(
		.INIT('h5554)
	) name7366 (
		\sa22_reg[2]/P0001 ,
		_w7519_,
		_w7561_,
		_w7823_,
		_w7899_
	);
	LUT3 #(
		.INIT('h54)
	) name7367 (
		\sa22_reg[1]/P0001 ,
		_w7592_,
		_w7899_,
		_w7900_
	);
	LUT4 #(
		.INIT('h0008)
	) name7368 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7901_
	);
	LUT4 #(
		.INIT('heff7)
	) name7369 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7902_
	);
	LUT2 #(
		.INIT('h2)
	) name7370 (
		_w7268_,
		_w7902_,
		_w7903_
	);
	LUT4 #(
		.INIT('h4000)
	) name7371 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w7904_
	);
	LUT4 #(
		.INIT('h0015)
	) name7372 (
		_w6978_,
		_w6923_,
		_w7287_,
		_w7904_,
		_w7905_
	);
	LUT3 #(
		.INIT('h31)
	) name7373 (
		_w7857_,
		_w7903_,
		_w7905_,
		_w7906_
	);
	LUT3 #(
		.INIT('h10)
	) name7374 (
		_w7898_,
		_w7900_,
		_w7906_,
		_w7907_
	);
	LUT3 #(
		.INIT('h10)
	) name7375 (
		_w7893_,
		_w7880_,
		_w7907_,
		_w7908_
	);
	LUT4 #(
		.INIT('h5655)
	) name7376 (
		\u0_w_reg[0][17]/P0001 ,
		_w7893_,
		_w7880_,
		_w7907_,
		_w7909_
	);
	LUT3 #(
		.INIT('h69)
	) name7377 (
		_w7817_,
		_w7865_,
		_w7909_,
		_w7910_
	);
	LUT4 #(
		.INIT('h1441)
	) name7378 (
		\ld_r_reg/P0001 ,
		_w7656_,
		_w7762_,
		_w7910_,
		_w7911_
	);
	LUT3 #(
		.INIT('h28)
	) name7379 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[113]/P0001 ,
		\u0_w_reg[0][17]/P0001 ,
		_w7912_
	);
	LUT2 #(
		.INIT('he)
	) name7380 (
		_w7911_,
		_w7912_,
		_w7913_
	);
	LUT3 #(
		.INIT('h02)
	) name7381 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7914_
	);
	LUT3 #(
		.INIT('had)
	) name7382 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7915_
	);
	LUT3 #(
		.INIT('h01)
	) name7383 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7916_
	);
	LUT3 #(
		.INIT('hf6)
	) name7384 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7917_
	);
	LUT3 #(
		.INIT('h2a)
	) name7385 (
		\sa33_reg[1]/P0001 ,
		_w7915_,
		_w7917_,
		_w7918_
	);
	LUT4 #(
		.INIT('h1000)
	) name7386 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7919_
	);
	LUT3 #(
		.INIT('h01)
	) name7387 (
		_w7084_,
		_w7079_,
		_w7919_,
		_w7920_
	);
	LUT3 #(
		.INIT('h8a)
	) name7388 (
		\sa33_reg[2]/P0001 ,
		_w7918_,
		_w7920_,
		_w7921_
	);
	LUT4 #(
		.INIT('h7d1d)
	) name7389 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7922_
	);
	LUT2 #(
		.INIT('h1)
	) name7390 (
		\sa33_reg[2]/P0001 ,
		_w7922_,
		_w7923_
	);
	LUT2 #(
		.INIT('h2)
	) name7391 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[5]/P0001 ,
		_w7924_
	);
	LUT2 #(
		.INIT('h8)
	) name7392 (
		_w7123_,
		_w7924_,
		_w7925_
	);
	LUT3 #(
		.INIT('h31)
	) name7393 (
		_w7075_,
		_w7142_,
		_w7335_,
		_w7926_
	);
	LUT4 #(
		.INIT('h5455)
	) name7394 (
		\sa33_reg[1]/P0001 ,
		_w7925_,
		_w7923_,
		_w7926_,
		_w7927_
	);
	LUT2 #(
		.INIT('h1)
	) name7395 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		_w7928_
	);
	LUT4 #(
		.INIT('h0100)
	) name7396 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7929_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name7397 (
		\sa33_reg[6]/P0001 ,
		_w7086_,
		_w7043_,
		_w7929_,
		_w7930_
	);
	LUT2 #(
		.INIT('h8)
	) name7398 (
		_w7108_,
		_w7069_,
		_w7931_
	);
	LUT3 #(
		.INIT('h13)
	) name7399 (
		_w7083_,
		_w7134_,
		_w7928_,
		_w7932_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7400 (
		\sa33_reg[1]/P0001 ,
		_w7930_,
		_w7931_,
		_w7932_,
		_w7933_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7401 (
		\sa33_reg[0]/P0001 ,
		_w7927_,
		_w7921_,
		_w7933_,
		_w7934_
	);
	LUT3 #(
		.INIT('h54)
	) name7402 (
		\sa33_reg[2]/P0001 ,
		_w7341_,
		_w7799_,
		_w7935_
	);
	LUT3 #(
		.INIT('h0d)
	) name7403 (
		_w7099_,
		_w7342_,
		_w7793_,
		_w7936_
	);
	LUT3 #(
		.INIT('h8a)
	) name7404 (
		\sa33_reg[1]/P0001 ,
		_w7935_,
		_w7936_,
		_w7937_
	);
	LUT3 #(
		.INIT('h80)
	) name7405 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7938_
	);
	LUT4 #(
		.INIT('h77f0)
	) name7406 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7939_
	);
	LUT4 #(
		.INIT('h4454)
	) name7407 (
		\sa33_reg[1]/P0001 ,
		_w7798_,
		_w7924_,
		_w7939_,
		_w7940_
	);
	LUT4 #(
		.INIT('h3fbb)
	) name7408 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7941_
	);
	LUT2 #(
		.INIT('h2)
	) name7409 (
		_w7928_,
		_w7941_,
		_w7942_
	);
	LUT4 #(
		.INIT('h0100)
	) name7410 (
		\sa33_reg[1]/P0001 ,
		\sa33_reg[2]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7943_
	);
	LUT4 #(
		.INIT('h00bf)
	) name7411 (
		\sa33_reg[7]/NET0131 ,
		_w7107_,
		_w7108_,
		_w7943_,
		_w7944_
	);
	LUT4 #(
		.INIT('h8000)
	) name7412 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7945_
	);
	LUT4 #(
		.INIT('h7ff7)
	) name7413 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7946_
	);
	LUT2 #(
		.INIT('h2)
	) name7414 (
		_w7138_,
		_w7946_,
		_w7947_
	);
	LUT4 #(
		.INIT('h0002)
	) name7415 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7948_
	);
	LUT4 #(
		.INIT('h5540)
	) name7416 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7063_,
		_w7948_,
		_w7949_
	);
	LUT4 #(
		.INIT('h0100)
	) name7417 (
		_w7947_,
		_w7949_,
		_w7942_,
		_w7944_,
		_w7950_
	);
	LUT4 #(
		.INIT('h5455)
	) name7418 (
		\sa33_reg[0]/P0001 ,
		_w7940_,
		_w7937_,
		_w7950_,
		_w7951_
	);
	LUT2 #(
		.INIT('h8)
	) name7419 (
		\sa33_reg[1]/P0001 ,
		\sa33_reg[2]/P0001 ,
		_w7952_
	);
	LUT4 #(
		.INIT('h0004)
	) name7420 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7953_
	);
	LUT4 #(
		.INIT('hadfb)
	) name7421 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7954_
	);
	LUT4 #(
		.INIT('h0302)
	) name7422 (
		\sa33_reg[3]/P0001 ,
		_w7116_,
		_w7323_,
		_w7954_,
		_w7955_
	);
	LUT2 #(
		.INIT('h2)
	) name7423 (
		_w7952_,
		_w7955_,
		_w7956_
	);
	LUT4 #(
		.INIT('h4000)
	) name7424 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7957_
	);
	LUT4 #(
		.INIT('h0007)
	) name7425 (
		_w7086_,
		_w7043_,
		_w7092_,
		_w7957_,
		_w7958_
	);
	LUT3 #(
		.INIT('h20)
	) name7426 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7959_
	);
	LUT3 #(
		.INIT('h15)
	) name7427 (
		_w7059_,
		_w7344_,
		_w7959_,
		_w7960_
	);
	LUT4 #(
		.INIT('h3100)
	) name7428 (
		\sa33_reg[2]/P0001 ,
		_w7942_,
		_w7958_,
		_w7960_,
		_w7961_
	);
	LUT4 #(
		.INIT('h1000)
	) name7429 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7962_
	);
	LUT4 #(
		.INIT('h0008)
	) name7430 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7963_
	);
	LUT4 #(
		.INIT('heff7)
	) name7431 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7964_
	);
	LUT4 #(
		.INIT('h4000)
	) name7432 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7965_
	);
	LUT4 #(
		.INIT('hbfef)
	) name7433 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7966_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name7434 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7967_
	);
	LUT3 #(
		.INIT('h20)
	) name7435 (
		\sa33_reg[1]/P0001 ,
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		_w7968_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name7436 (
		_w7342_,
		_w7964_,
		_w7967_,
		_w7968_,
		_w7969_
	);
	LUT4 #(
		.INIT('h0e00)
	) name7437 (
		\sa33_reg[1]/P0001 ,
		_w7961_,
		_w7956_,
		_w7969_,
		_w7970_
	);
	LUT3 #(
		.INIT('h10)
	) name7438 (
		_w7951_,
		_w7934_,
		_w7970_,
		_w7971_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name7439 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7972_
	);
	LUT2 #(
		.INIT('h2)
	) name7440 (
		\sa33_reg[2]/P0001 ,
		_w7972_,
		_w7973_
	);
	LUT4 #(
		.INIT('h0002)
	) name7441 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7974_
	);
	LUT4 #(
		.INIT('h5540)
	) name7442 (
		\sa33_reg[5]/P0001 ,
		_w7049_,
		_w7302_,
		_w7974_,
		_w7975_
	);
	LUT4 #(
		.INIT('h0010)
	) name7443 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7976_
	);
	LUT3 #(
		.INIT('h01)
	) name7444 (
		_w7098_,
		_w7060_,
		_w7976_,
		_w7977_
	);
	LUT4 #(
		.INIT('h5455)
	) name7445 (
		\sa33_reg[1]/P0001 ,
		_w7975_,
		_w7973_,
		_w7977_,
		_w7978_
	);
	LUT3 #(
		.INIT('h0b)
	) name7446 (
		\sa33_reg[6]/P0001 ,
		_w7063_,
		_w7798_,
		_w7979_
	);
	LUT4 #(
		.INIT('h0100)
	) name7447 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7980_
	);
	LUT3 #(
		.INIT('h0b)
	) name7448 (
		\sa33_reg[6]/P0001 ,
		_w7059_,
		_w7980_,
		_w7981_
	);
	LUT3 #(
		.INIT('h2a)
	) name7449 (
		\sa33_reg[2]/P0001 ,
		_w7979_,
		_w7981_,
		_w7982_
	);
	LUT3 #(
		.INIT('h54)
	) name7450 (
		\sa33_reg[2]/P0001 ,
		_w7134_,
		_w7945_,
		_w7983_
	);
	LUT3 #(
		.INIT('h51)
	) name7451 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7984_
	);
	LUT4 #(
		.INIT('h4041)
	) name7452 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7985_
	);
	LUT3 #(
		.INIT('ha8)
	) name7453 (
		\sa33_reg[1]/P0001 ,
		_w7772_,
		_w7985_,
		_w7986_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name7454 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7987_
	);
	LUT2 #(
		.INIT('h2)
	) name7455 (
		_w7113_,
		_w7987_,
		_w7988_
	);
	LUT3 #(
		.INIT('h07)
	) name7456 (
		_w7033_,
		_w7126_,
		_w7313_,
		_w7989_
	);
	LUT4 #(
		.INIT('h0100)
	) name7457 (
		_w7986_,
		_w7988_,
		_w7983_,
		_w7989_,
		_w7990_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7458 (
		\sa33_reg[0]/P0001 ,
		_w7982_,
		_w7978_,
		_w7990_,
		_w7991_
	);
	LUT2 #(
		.INIT('h8)
	) name7459 (
		\sa33_reg[2]/P0001 ,
		_w7323_,
		_w7992_
	);
	LUT4 #(
		.INIT('h7ff8)
	) name7460 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7993_
	);
	LUT3 #(
		.INIT('h20)
	) name7461 (
		\sa33_reg[1]/P0001 ,
		_w7929_,
		_w7993_,
		_w7994_
	);
	LUT2 #(
		.INIT('h1)
	) name7462 (
		\sa33_reg[3]/P0001 ,
		_w7966_,
		_w7995_
	);
	LUT3 #(
		.INIT('h15)
	) name7463 (
		\sa33_reg[1]/P0001 ,
		_w7341_,
		_w7342_,
		_w7996_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name7464 (
		_w7992_,
		_w7994_,
		_w7995_,
		_w7996_,
		_w7997_
	);
	LUT3 #(
		.INIT('hb9)
	) name7465 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7998_
	);
	LUT3 #(
		.INIT('h40)
	) name7466 (
		\sa33_reg[1]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w7999_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name7467 (
		_w7033_,
		_w7339_,
		_w7998_,
		_w7999_,
		_w8000_
	);
	LUT4 #(
		.INIT('h0001)
	) name7468 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w8001_
	);
	LUT4 #(
		.INIT('h000b)
	) name7469 (
		\sa33_reg[6]/P0001 ,
		_w7059_,
		_w7786_,
		_w8001_,
		_w8002_
	);
	LUT3 #(
		.INIT('hd8)
	) name7470 (
		\sa33_reg[2]/P0001 ,
		_w8000_,
		_w8002_,
		_w8003_
	);
	LUT3 #(
		.INIT('h45)
	) name7471 (
		\sa33_reg[0]/P0001 ,
		_w7997_,
		_w8003_,
		_w8004_
	);
	LUT4 #(
		.INIT('h4000)
	) name7472 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8005_
	);
	LUT4 #(
		.INIT('haa80)
	) name7473 (
		\sa33_reg[6]/P0001 ,
		_w7055_,
		_w7038_,
		_w8005_,
		_w8006_
	);
	LUT2 #(
		.INIT('h8)
	) name7474 (
		_w7767_,
		_w7928_,
		_w8007_
	);
	LUT4 #(
		.INIT('habaf)
	) name7475 (
		\sa33_reg[5]/P0001 ,
		_w7052_,
		_w7131_,
		_w7138_,
		_w8008_
	);
	LUT3 #(
		.INIT('h40)
	) name7476 (
		\sa33_reg[5]/P0001 ,
		_w7083_,
		_w7055_,
		_w8009_
	);
	LUT4 #(
		.INIT('h0200)
	) name7477 (
		_w7331_,
		_w8007_,
		_w8009_,
		_w8008_,
		_w8010_
	);
	LUT4 #(
		.INIT('h002a)
	) name7478 (
		\sa33_reg[2]/P0001 ,
		_w7107_,
		_w7123_,
		_w7962_,
		_w8011_
	);
	LUT2 #(
		.INIT('h4)
	) name7479 (
		_w7087_,
		_w7075_,
		_w8012_
	);
	LUT3 #(
		.INIT('h15)
	) name7480 (
		\sa33_reg[2]/P0001 ,
		_w7066_,
		_w7139_,
		_w8013_
	);
	LUT3 #(
		.INIT('h45)
	) name7481 (
		_w8011_,
		_w8012_,
		_w8013_,
		_w8014_
	);
	LUT3 #(
		.INIT('h15)
	) name7482 (
		\sa33_reg[1]/P0001 ,
		_w7088_,
		_w7113_,
		_w8015_
	);
	LUT2 #(
		.INIT('h4)
	) name7483 (
		_w7140_,
		_w8015_,
		_w8016_
	);
	LUT4 #(
		.INIT('h4544)
	) name7484 (
		_w8006_,
		_w8010_,
		_w8014_,
		_w8016_,
		_w8017_
	);
	LUT3 #(
		.INIT('h10)
	) name7485 (
		_w7991_,
		_w8004_,
		_w8017_,
		_w8018_
	);
	LUT4 #(
		.INIT('h5655)
	) name7486 (
		\u0_w_reg[0][9]/P0001 ,
		_w7797_,
		_w7782_,
		_w7816_,
		_w8019_
	);
	LUT3 #(
		.INIT('h69)
	) name7487 (
		_w7971_,
		_w8018_,
		_w8019_,
		_w8020_
	);
	LUT2 #(
		.INIT('h9)
	) name7488 (
		_w7603_,
		_w7908_,
		_w8021_
	);
	LUT4 #(
		.INIT('h5510)
	) name7489 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w6896_,
		_w7474_,
		_w8022_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name7490 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8023_
	);
	LUT2 #(
		.INIT('h2)
	) name7491 (
		\sa11_reg[2]/P0001 ,
		_w8023_,
		_w8024_
	);
	LUT4 #(
		.INIT('h153f)
	) name7492 (
		_w6634_,
		_w6658_,
		_w6671_,
		_w6681_,
		_w8025_
	);
	LUT4 #(
		.INIT('h5455)
	) name7493 (
		\sa11_reg[1]/P0001 ,
		_w8024_,
		_w8022_,
		_w8025_,
		_w8026_
	);
	LUT4 #(
		.INIT('h0800)
	) name7494 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w8027_
	);
	LUT4 #(
		.INIT('h5554)
	) name7495 (
		\sa11_reg[2]/P0001 ,
		_w6851_,
		_w7465_,
		_w8027_,
		_w8028_
	);
	LUT3 #(
		.INIT('ha8)
	) name7496 (
		\sa11_reg[2]/P0001 ,
		_w6884_,
		_w7691_,
		_w8029_
	);
	LUT3 #(
		.INIT('h01)
	) name7497 (
		_w6721_,
		_w6672_,
		_w6868_,
		_w8030_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7498 (
		\sa11_reg[1]/P0001 ,
		_w8029_,
		_w8028_,
		_w8030_,
		_w8031_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name7499 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w6636_,
		_w6681_,
		_w8032_
	);
	LUT4 #(
		.INIT('hffa8)
	) name7500 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8033_
	);
	LUT2 #(
		.INIT('h2)
	) name7501 (
		_w6640_,
		_w8033_,
		_w8034_
	);
	LUT4 #(
		.INIT('h007f)
	) name7502 (
		\sa11_reg[4]/P0001 ,
		_w6730_,
		_w6676_,
		_w6719_,
		_w8035_
	);
	LUT4 #(
		.INIT('h0e00)
	) name7503 (
		\sa11_reg[2]/P0001 ,
		_w8032_,
		_w8034_,
		_w8035_,
		_w8036_
	);
	LUT4 #(
		.INIT('h5455)
	) name7504 (
		\sa11_reg[0]/P0001 ,
		_w8031_,
		_w8026_,
		_w8036_,
		_w8037_
	);
	LUT3 #(
		.INIT('h07)
	) name7505 (
		_w6879_,
		_w6847_,
		_w6896_,
		_w8038_
	);
	LUT4 #(
		.INIT('h3120)
	) name7506 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8039_
	);
	LUT3 #(
		.INIT('h80)
	) name7507 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8040_
	);
	LUT3 #(
		.INIT('ha8)
	) name7508 (
		\sa11_reg[2]/P0001 ,
		_w8039_,
		_w8040_,
		_w8041_
	);
	LUT3 #(
		.INIT('ha2)
	) name7509 (
		\sa11_reg[1]/P0001 ,
		_w8038_,
		_w8041_,
		_w8042_
	);
	LUT4 #(
		.INIT('h8880)
	) name7510 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w8043_
	);
	LUT4 #(
		.INIT('h0203)
	) name7511 (
		_w6663_,
		_w6733_,
		_w6872_,
		_w8043_,
		_w8044_
	);
	LUT2 #(
		.INIT('h1)
	) name7512 (
		\sa11_reg[1]/P0001 ,
		_w8044_,
		_w8045_
	);
	LUT4 #(
		.INIT('h0008)
	) name7513 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8046_
	);
	LUT4 #(
		.INIT('h0001)
	) name7514 (
		_w6648_,
		_w6733_,
		_w7684_,
		_w8046_,
		_w8047_
	);
	LUT2 #(
		.INIT('h1)
	) name7515 (
		\sa11_reg[2]/P0001 ,
		_w8047_,
		_w8048_
	);
	LUT2 #(
		.INIT('h4)
	) name7516 (
		\sa11_reg[1]/P0001 ,
		_w7438_,
		_w8049_
	);
	LUT3 #(
		.INIT('h0d)
	) name7517 (
		_w6664_,
		_w6707_,
		_w8046_,
		_w8050_
	);
	LUT3 #(
		.INIT('h45)
	) name7518 (
		\sa11_reg[3]/P0001 ,
		_w8049_,
		_w8050_,
		_w8051_
	);
	LUT4 #(
		.INIT('h0001)
	) name7519 (
		_w8042_,
		_w8048_,
		_w8051_,
		_w8045_,
		_w8052_
	);
	LUT4 #(
		.INIT('h0007)
	) name7520 (
		_w6674_,
		_w6696_,
		_w7444_,
		_w7682_,
		_w8053_
	);
	LUT4 #(
		.INIT('hedff)
	) name7521 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w6644_,
		_w8054_
	);
	LUT4 #(
		.INIT('h0155)
	) name7522 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[2]/P0001 ,
		_w8053_,
		_w8054_,
		_w8055_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name7523 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8056_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7524 (
		\sa11_reg[3]/P0001 ,
		_w6637_,
		_w7457_,
		_w8056_,
		_w8057_
	);
	LUT3 #(
		.INIT('h80)
	) name7525 (
		\sa11_reg[4]/P0001 ,
		_w6730_,
		_w6691_,
		_w8058_
	);
	LUT3 #(
		.INIT('h2e)
	) name7526 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[2]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w8059_
	);
	LUT2 #(
		.INIT('h8)
	) name7527 (
		_w6868_,
		_w8059_,
		_w8060_
	);
	LUT4 #(
		.INIT('h0031)
	) name7528 (
		_w7480_,
		_w8058_,
		_w8057_,
		_w8060_,
		_w8061_
	);
	LUT4 #(
		.INIT('h0010)
	) name7529 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w8062_
	);
	LUT4 #(
		.INIT('hffbe)
	) name7530 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8063_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name7531 (
		_w6677_,
		_w7484_,
		_w8062_,
		_w8063_,
		_w8064_
	);
	LUT4 #(
		.INIT('h0023)
	) name7532 (
		\sa11_reg[3]/P0001 ,
		_w6719_,
		_w6848_,
		_w7622_,
		_w8065_
	);
	LUT3 #(
		.INIT('h31)
	) name7533 (
		_w7701_,
		_w8064_,
		_w8065_,
		_w8066_
	);
	LUT3 #(
		.INIT('h40)
	) name7534 (
		_w8055_,
		_w8061_,
		_w8066_,
		_w8067_
	);
	LUT4 #(
		.INIT('h3100)
	) name7535 (
		\sa11_reg[0]/P0001 ,
		_w8037_,
		_w8052_,
		_w8067_,
		_w8068_
	);
	LUT3 #(
		.INIT('h4b)
	) name7536 (
		_w7725_,
		_w7761_,
		_w8068_,
		_w8069_
	);
	LUT4 #(
		.INIT('h1441)
	) name7537 (
		\ld_r_reg/P0001 ,
		_w8020_,
		_w8021_,
		_w8069_,
		_w8070_
	);
	LUT3 #(
		.INIT('h28)
	) name7538 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[105]/P0001 ,
		\u0_w_reg[0][9]/P0001 ,
		_w8071_
	);
	LUT2 #(
		.INIT('he)
	) name7539 (
		_w8070_,
		_w8071_,
		_w8072_
	);
	LUT4 #(
		.INIT('h6996)
	) name7540 (
		\u0_w_reg[0][1]/P0001 ,
		_w7865_,
		_w7971_,
		_w8018_,
		_w8073_
	);
	LUT4 #(
		.INIT('hbfef)
	) name7541 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8074_
	);
	LUT4 #(
		.INIT('haf8c)
	) name7542 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		_w6809_,
		_w8074_,
		_w8075_
	);
	LUT2 #(
		.INIT('h1)
	) name7543 (
		\sa00_reg[1]/P0001 ,
		_w8075_,
		_w8076_
	);
	LUT2 #(
		.INIT('h8)
	) name7544 (
		\sa00_reg[3]/P0001 ,
		_w6751_,
		_w8077_
	);
	LUT4 #(
		.INIT('hfff8)
	) name7545 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8078_
	);
	LUT2 #(
		.INIT('h1)
	) name7546 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		_w8079_
	);
	LUT4 #(
		.INIT('h0100)
	) name7547 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w8080_
	);
	LUT4 #(
		.INIT('h8000)
	) name7548 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8081_
	);
	LUT3 #(
		.INIT('h10)
	) name7549 (
		_w8080_,
		_w8081_,
		_w8078_,
		_w8082_
	);
	LUT3 #(
		.INIT('h8a)
	) name7550 (
		\sa00_reg[1]/P0001 ,
		_w8077_,
		_w8082_,
		_w8083_
	);
	LUT4 #(
		.INIT('h8000)
	) name7551 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8084_
	);
	LUT4 #(
		.INIT('h0013)
	) name7552 (
		_w6780_,
		_w7398_,
		_w7757_,
		_w8084_,
		_w8085_
	);
	LUT3 #(
		.INIT('hb9)
	) name7553 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8086_
	);
	LUT4 #(
		.INIT('h4c00)
	) name7554 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8087_
	);
	LUT4 #(
		.INIT('h31f5)
	) name7555 (
		_w7164_,
		_w7389_,
		_w8086_,
		_w8087_,
		_w8088_
	);
	LUT3 #(
		.INIT('he0)
	) name7556 (
		\sa00_reg[2]/P0001 ,
		_w8085_,
		_w8088_,
		_w8089_
	);
	LUT4 #(
		.INIT('h5455)
	) name7557 (
		\sa00_reg[0]/P0001 ,
		_w8076_,
		_w8083_,
		_w8089_,
		_w8090_
	);
	LUT4 #(
		.INIT('h0001)
	) name7558 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8091_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name7559 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8092_
	);
	LUT3 #(
		.INIT('h8a)
	) name7560 (
		\sa00_reg[2]/P0001 ,
		_w8091_,
		_w8092_,
		_w8093_
	);
	LUT2 #(
		.INIT('h8)
	) name7561 (
		_w6795_,
		_w8079_,
		_w8094_
	);
	LUT3 #(
		.INIT('h8a)
	) name7562 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8095_
	);
	LUT4 #(
		.INIT('h0010)
	) name7563 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w8096_
	);
	LUT3 #(
		.INIT('h0d)
	) name7564 (
		_w6738_,
		_w8095_,
		_w8096_,
		_w8097_
	);
	LUT4 #(
		.INIT('h5455)
	) name7565 (
		\sa00_reg[1]/P0001 ,
		_w8094_,
		_w8093_,
		_w8097_,
		_w8098_
	);
	LUT3 #(
		.INIT('h13)
	) name7566 (
		_w6780_,
		_w6742_,
		_w7757_,
		_w8099_
	);
	LUT3 #(
		.INIT('h2a)
	) name7567 (
		\sa00_reg[2]/P0001 ,
		_w7382_,
		_w8099_,
		_w8100_
	);
	LUT4 #(
		.INIT('h0001)
	) name7568 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8101_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7569 (
		\sa00_reg[1]/P0001 ,
		_w6755_,
		_w7415_,
		_w8101_,
		_w8102_
	);
	LUT4 #(
		.INIT('h8000)
	) name7570 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8103_
	);
	LUT3 #(
		.INIT('h54)
	) name7571 (
		\sa00_reg[2]/P0001 ,
		_w7396_,
		_w8103_,
		_w8104_
	);
	LUT2 #(
		.INIT('h4)
	) name7572 (
		_w7197_,
		_w7402_,
		_w8105_
	);
	LUT3 #(
		.INIT('h0b)
	) name7573 (
		\sa00_reg[6]/NET0131 ,
		_w6829_,
		_w7712_,
		_w8106_
	);
	LUT4 #(
		.INIT('h0100)
	) name7574 (
		_w8102_,
		_w8105_,
		_w8104_,
		_w8106_,
		_w8107_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7575 (
		\sa00_reg[0]/P0001 ,
		_w8100_,
		_w8098_,
		_w8107_,
		_w8108_
	);
	LUT3 #(
		.INIT('h04)
	) name7576 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8109_
	);
	LUT4 #(
		.INIT('h5140)
	) name7577 (
		\sa00_reg[2]/P0001 ,
		_w6769_,
		_w6770_,
		_w8109_,
		_w8110_
	);
	LUT3 #(
		.INIT('h02)
	) name7578 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w8111_
	);
	LUT3 #(
		.INIT('h67)
	) name7579 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8112_
	);
	LUT2 #(
		.INIT('h2)
	) name7580 (
		_w8111_,
		_w8112_,
		_w8113_
	);
	LUT2 #(
		.INIT('h8)
	) name7581 (
		_w7385_,
		_w7402_,
		_w8114_
	);
	LUT4 #(
		.INIT('h0001)
	) name7582 (
		_w7220_,
		_w8110_,
		_w8113_,
		_w8114_,
		_w8115_
	);
	LUT3 #(
		.INIT('h04)
	) name7583 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w8116_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name7584 (
		\sa00_reg[6]/NET0131 ,
		_w6832_,
		_w7403_,
		_w8116_,
		_w8117_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name7585 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w6813_,
		_w6790_,
		_w8118_
	);
	LUT2 #(
		.INIT('h8)
	) name7586 (
		_w7169_,
		_w8079_,
		_w8119_
	);
	LUT4 #(
		.INIT('hdeff)
	) name7587 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w6758_,
		_w8120_
	);
	LUT3 #(
		.INIT('h10)
	) name7588 (
		_w8118_,
		_w8119_,
		_w8120_,
		_w8121_
	);
	LUT4 #(
		.INIT('h3120)
	) name7589 (
		\sa00_reg[1]/P0001 ,
		_w8117_,
		_w8121_,
		_w8115_,
		_w8122_
	);
	LUT3 #(
		.INIT('h10)
	) name7590 (
		_w8108_,
		_w8090_,
		_w8122_,
		_w8123_
	);
	LUT4 #(
		.INIT('h7f5f)
	) name7591 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8124_
	);
	LUT4 #(
		.INIT('h5455)
	) name7592 (
		\sa00_reg[2]/P0001 ,
		_w7393_,
		_w8109_,
		_w8124_,
		_w8125_
	);
	LUT3 #(
		.INIT('h54)
	) name7593 (
		\sa00_reg[7]/NET0131 ,
		_w6755_,
		_w7399_,
		_w8126_
	);
	LUT3 #(
		.INIT('h15)
	) name7594 (
		_w6778_,
		_w6832_,
		_w6741_,
		_w8127_
	);
	LUT4 #(
		.INIT('h5455)
	) name7595 (
		\sa00_reg[1]/P0001 ,
		_w8125_,
		_w8126_,
		_w8127_,
		_w8128_
	);
	LUT4 #(
		.INIT('hcfca)
	) name7596 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8129_
	);
	LUT3 #(
		.INIT('h08)
	) name7597 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8130_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7598 (
		\sa00_reg[1]/P0001 ,
		_w7393_,
		_w8130_,
		_w8129_,
		_w8131_
	);
	LUT3 #(
		.INIT('h01)
	) name7599 (
		_w6823_,
		_w7156_,
		_w7151_,
		_w8132_
	);
	LUT3 #(
		.INIT('h8a)
	) name7600 (
		\sa00_reg[2]/P0001 ,
		_w8131_,
		_w8132_,
		_w8133_
	);
	LUT4 #(
		.INIT('h0777)
	) name7601 (
		_w6765_,
		_w6828_,
		_w7210_,
		_w8079_,
		_w8134_
	);
	LUT2 #(
		.INIT('h8)
	) name7602 (
		_w6772_,
		_w8109_,
		_w8135_
	);
	LUT3 #(
		.INIT('h07)
	) name7603 (
		_w6831_,
		_w6766_,
		_w7396_,
		_w8136_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7604 (
		\sa00_reg[1]/P0001 ,
		_w8134_,
		_w8135_,
		_w8136_,
		_w8137_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7605 (
		\sa00_reg[0]/P0001 ,
		_w8133_,
		_w8128_,
		_w8137_,
		_w8138_
	);
	LUT4 #(
		.INIT('hddd8)
	) name7606 (
		\sa00_reg[2]/P0001 ,
		_w6790_,
		_w7191_,
		_w7727_,
		_w8139_
	);
	LUT3 #(
		.INIT('h07)
	) name7607 (
		_w6744_,
		_w7399_,
		_w7414_,
		_w8140_
	);
	LUT3 #(
		.INIT('h8a)
	) name7608 (
		\sa00_reg[1]/P0001 ,
		_w8139_,
		_w8140_,
		_w8141_
	);
	LUT2 #(
		.INIT('h1)
	) name7609 (
		_w7739_,
		_w8096_,
		_w8142_
	);
	LUT3 #(
		.INIT('h07)
	) name7610 (
		\sa00_reg[5]/P0001 ,
		_w6749_,
		_w7425_,
		_w8143_
	);
	LUT3 #(
		.INIT('h15)
	) name7611 (
		\sa00_reg[2]/P0001 ,
		_w8142_,
		_w8143_,
		_w8144_
	);
	LUT4 #(
		.INIT('h7ff6)
	) name7612 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8145_
	);
	LUT2 #(
		.INIT('h2)
	) name7613 (
		_w6831_,
		_w8145_,
		_w8146_
	);
	LUT4 #(
		.INIT('h77f0)
	) name7614 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8147_
	);
	LUT3 #(
		.INIT('h10)
	) name7615 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w8148_
	);
	LUT4 #(
		.INIT('h0031)
	) name7616 (
		_w7387_,
		_w7381_,
		_w8147_,
		_w8148_,
		_w8149_
	);
	LUT3 #(
		.INIT('h32)
	) name7617 (
		\sa00_reg[1]/P0001 ,
		_w8146_,
		_w8149_,
		_w8150_
	);
	LUT4 #(
		.INIT('h5455)
	) name7618 (
		\sa00_reg[0]/P0001 ,
		_w8144_,
		_w8141_,
		_w8150_,
		_w8151_
	);
	LUT4 #(
		.INIT('h0004)
	) name7619 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8152_
	);
	LUT4 #(
		.INIT('hadfb)
	) name7620 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8153_
	);
	LUT4 #(
		.INIT('h0302)
	) name7621 (
		\sa00_reg[3]/P0001 ,
		_w6777_,
		_w7175_,
		_w8153_,
		_w8154_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name7622 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8155_
	);
	LUT2 #(
		.INIT('h2)
	) name7623 (
		_w7402_,
		_w8155_,
		_w8156_
	);
	LUT4 #(
		.INIT('haa08)
	) name7624 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[2]/P0001 ,
		_w8154_,
		_w8156_,
		_w8157_
	);
	LUT4 #(
		.INIT('h4000)
	) name7625 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w8158_
	);
	LUT4 #(
		.INIT('hbdff)
	) name7626 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w8159_
	);
	LUT3 #(
		.INIT('h10)
	) name7627 (
		_w7739_,
		_w8096_,
		_w8159_,
		_w8160_
	);
	LUT2 #(
		.INIT('h2)
	) name7628 (
		\sa00_reg[2]/P0001 ,
		_w8158_,
		_w8161_
	);
	LUT3 #(
		.INIT('h51)
	) name7629 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[2]/P0001 ,
		_w8158_,
		_w8162_
	);
	LUT2 #(
		.INIT('h4)
	) name7630 (
		_w8160_,
		_w8162_,
		_w8163_
	);
	LUT4 #(
		.INIT('h153f)
	) name7631 (
		_w6747_,
		_w6763_,
		_w6764_,
		_w7206_,
		_w8164_
	);
	LUT4 #(
		.INIT('h4000)
	) name7632 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w8165_
	);
	LUT4 #(
		.INIT('h0007)
	) name7633 (
		_w6765_,
		_w6828_,
		_w7160_,
		_w8165_,
		_w8166_
	);
	LUT4 #(
		.INIT('hfcb8)
	) name7634 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[2]/P0001 ,
		_w8164_,
		_w8166_,
		_w8167_
	);
	LUT3 #(
		.INIT('h10)
	) name7635 (
		_w8157_,
		_w8163_,
		_w8167_,
		_w8168_
	);
	LUT3 #(
		.INIT('h10)
	) name7636 (
		_w8151_,
		_w8138_,
		_w8168_,
		_w8169_
	);
	LUT2 #(
		.INIT('h9)
	) name7637 (
		_w8123_,
		_w8169_,
		_w8170_
	);
	LUT4 #(
		.INIT('h1441)
	) name7638 (
		\ld_r_reg/P0001 ,
		_w8069_,
		_w8073_,
		_w8170_,
		_w8171_
	);
	LUT3 #(
		.INIT('h28)
	) name7639 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[97]/P0001 ,
		\u0_w_reg[0][1]/P0001 ,
		_w8172_
	);
	LUT2 #(
		.INIT('he)
	) name7640 (
		_w8171_,
		_w8172_,
		_w8173_
	);
	LUT4 #(
		.INIT('hefdf)
	) name7641 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8174_
	);
	LUT2 #(
		.INIT('h1)
	) name7642 (
		\sa11_reg[2]/P0001 ,
		_w8174_,
		_w8175_
	);
	LUT4 #(
		.INIT('hff3b)
	) name7643 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8176_
	);
	LUT2 #(
		.INIT('h2)
	) name7644 (
		\sa11_reg[2]/P0001 ,
		_w8176_,
		_w8177_
	);
	LUT4 #(
		.INIT('h0015)
	) name7645 (
		_w6719_,
		_w6674_,
		_w6675_,
		_w6870_,
		_w8178_
	);
	LUT4 #(
		.INIT('h0100)
	) name7646 (
		_w7640_,
		_w8175_,
		_w8177_,
		_w8178_,
		_w8179_
	);
	LUT4 #(
		.INIT('h0c04)
	) name7647 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8180_
	);
	LUT3 #(
		.INIT('ha8)
	) name7648 (
		\sa11_reg[2]/P0001 ,
		_w6641_,
		_w8180_,
		_w8181_
	);
	LUT3 #(
		.INIT('h01)
	) name7649 (
		_w6704_,
		_w6717_,
		_w7664_,
		_w8182_
	);
	LUT2 #(
		.INIT('h1)
	) name7650 (
		_w7627_,
		_w7637_,
		_w8183_
	);
	LUT3 #(
		.INIT('h40)
	) name7651 (
		_w8181_,
		_w8182_,
		_w8183_,
		_w8184_
	);
	LUT4 #(
		.INIT('h0100)
	) name7652 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w8185_
	);
	LUT4 #(
		.INIT('h0007)
	) name7653 (
		_w6636_,
		_w6682_,
		_w7612_,
		_w8185_,
		_w8186_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name7654 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8187_
	);
	LUT4 #(
		.INIT('h7707)
	) name7655 (
		_w6642_,
		_w6634_,
		_w6651_,
		_w8187_,
		_w8188_
	);
	LUT3 #(
		.INIT('he0)
	) name7656 (
		\sa11_reg[2]/P0001 ,
		_w8186_,
		_w8188_,
		_w8189_
	);
	LUT4 #(
		.INIT('he400)
	) name7657 (
		\sa11_reg[1]/P0001 ,
		_w8179_,
		_w8184_,
		_w8189_,
		_w8190_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name7658 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w6885_,
		_w7455_,
		_w8191_
	);
	LUT4 #(
		.INIT('h002a)
	) name7659 (
		\sa11_reg[1]/P0001 ,
		_w6650_,
		_w6725_,
		_w6714_,
		_w8192_
	);
	LUT4 #(
		.INIT('h153f)
	) name7660 (
		_w6635_,
		_w6879_,
		_w6847_,
		_w7680_,
		_w8193_
	);
	LUT3 #(
		.INIT('h40)
	) name7661 (
		_w8191_,
		_w8192_,
		_w8193_,
		_w8194_
	);
	LUT4 #(
		.INIT('h0008)
	) name7662 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8195_
	);
	LUT3 #(
		.INIT('h01)
	) name7663 (
		\sa11_reg[1]/P0001 ,
		_w8185_,
		_w8195_,
		_w8196_
	);
	LUT3 #(
		.INIT('h20)
	) name7664 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w8197_
	);
	LUT3 #(
		.INIT('h23)
	) name7665 (
		_w6674_,
		_w7481_,
		_w8197_,
		_w8198_
	);
	LUT3 #(
		.INIT('h40)
	) name7666 (
		_w7488_,
		_w8196_,
		_w8198_,
		_w8199_
	);
	LUT4 #(
		.INIT('h0405)
	) name7667 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w6645_,
		_w6848_,
		_w8200_
	);
	LUT4 #(
		.INIT('h0002)
	) name7668 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[7]/NET0131 ,
		_w8201_
	);
	LUT3 #(
		.INIT('h02)
	) name7669 (
		\sa11_reg[2]/P0001 ,
		_w6713_,
		_w8201_,
		_w8202_
	);
	LUT3 #(
		.INIT('h54)
	) name7670 (
		_w6862_,
		_w8200_,
		_w8202_,
		_w8203_
	);
	LUT3 #(
		.INIT('he0)
	) name7671 (
		_w8194_,
		_w8199_,
		_w8203_,
		_w8204_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name7672 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8205_
	);
	LUT2 #(
		.INIT('h2)
	) name7673 (
		_w7441_,
		_w8205_,
		_w8206_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name7674 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[4]/P0001 ,
		_w6636_,
		_w6714_,
		_w8207_
	);
	LUT3 #(
		.INIT('h8a)
	) name7675 (
		\sa11_reg[1]/P0001 ,
		_w8206_,
		_w8207_,
		_w8208_
	);
	LUT4 #(
		.INIT('h153f)
	) name7676 (
		_w6686_,
		_w6674_,
		_w6696_,
		_w6861_,
		_w8209_
	);
	LUT4 #(
		.INIT('h3777)
	) name7677 (
		_w6658_,
		_w6671_,
		_w6697_,
		_w6908_,
		_w8210_
	);
	LUT3 #(
		.INIT('hd0)
	) name7678 (
		_w7701_,
		_w8209_,
		_w8210_,
		_w8211_
	);
	LUT4 #(
		.INIT('hedff)
	) name7679 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8212_
	);
	LUT2 #(
		.INIT('h2)
	) name7680 (
		_w6730_,
		_w8212_,
		_w8213_
	);
	LUT4 #(
		.INIT('h2000)
	) name7681 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w8214_
	);
	LUT3 #(
		.INIT('hc8)
	) name7682 (
		_w6717_,
		_w7480_,
		_w8214_,
		_w8215_
	);
	LUT2 #(
		.INIT('h1)
	) name7683 (
		_w8213_,
		_w8215_,
		_w8216_
	);
	LUT3 #(
		.INIT('h40)
	) name7684 (
		_w8208_,
		_w8211_,
		_w8216_,
		_w8217_
	);
	LUT4 #(
		.INIT('hd800)
	) name7685 (
		\sa11_reg[0]/P0001 ,
		_w8190_,
		_w8204_,
		_w8217_,
		_w8218_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7686 (
		\sa22_reg[2]/P0001 ,
		_w6950_,
		_w6958_,
		_w7225_,
		_w8219_
	);
	LUT2 #(
		.INIT('h1)
	) name7687 (
		_w7008_,
		_w7277_,
		_w8220_
	);
	LUT4 #(
		.INIT('h0010)
	) name7688 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w8221_
	);
	LUT4 #(
		.INIT('h0001)
	) name7689 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w8222_
	);
	LUT3 #(
		.INIT('h01)
	) name7690 (
		_w7592_,
		_w8222_,
		_w8221_,
		_w8223_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name7691 (
		\sa22_reg[1]/P0001 ,
		_w8219_,
		_w8220_,
		_w8223_,
		_w8224_
	);
	LUT4 #(
		.INIT('hff3b)
	) name7692 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w8225_
	);
	LUT3 #(
		.INIT('h20)
	) name7693 (
		\sa22_reg[2]/P0001 ,
		_w6941_,
		_w8225_,
		_w8226_
	);
	LUT3 #(
		.INIT('h01)
	) name7694 (
		\sa22_reg[2]/P0001 ,
		_w6981_,
		_w7291_,
		_w8227_
	);
	LUT4 #(
		.INIT('h0103)
	) name7695 (
		_w6953_,
		_w6980_,
		_w7015_,
		_w7255_,
		_w8228_
	);
	LUT4 #(
		.INIT('h0155)
	) name7696 (
		\sa22_reg[1]/P0001 ,
		_w8226_,
		_w8227_,
		_w8228_,
		_w8229_
	);
	LUT4 #(
		.INIT('h0100)
	) name7697 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w8230_
	);
	LUT4 #(
		.INIT('h0007)
	) name7698 (
		_w6923_,
		_w6950_,
		_w7586_,
		_w8230_,
		_w8231_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name7699 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w8232_
	);
	LUT2 #(
		.INIT('h8)
	) name7700 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w8233_
	);
	LUT4 #(
		.INIT('h7077)
	) name7701 (
		_w6921_,
		_w6946_,
		_w8232_,
		_w8233_,
		_w8234_
	);
	LUT3 #(
		.INIT('he0)
	) name7702 (
		\sa22_reg[2]/P0001 ,
		_w8231_,
		_w8234_,
		_w8235_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7703 (
		\sa22_reg[0]/P0001 ,
		_w8229_,
		_w8224_,
		_w8235_,
		_w8236_
	);
	LUT4 #(
		.INIT('haa80)
	) name7704 (
		\sa22_reg[2]/P0001 ,
		_w6944_,
		_w6954_,
		_w7019_,
		_w8237_
	);
	LUT2 #(
		.INIT('h4)
	) name7705 (
		\sa22_reg[2]/P0001 ,
		_w6983_,
		_w8238_
	);
	LUT3 #(
		.INIT('h07)
	) name7706 (
		\sa22_reg[7]/NET0131 ,
		_w6980_,
		_w6941_,
		_w8239_
	);
	LUT4 #(
		.INIT('h0100)
	) name7707 (
		_w7837_,
		_w8238_,
		_w8237_,
		_w8239_,
		_w8240_
	);
	LUT4 #(
		.INIT('h5400)
	) name7708 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w8241_
	);
	LUT3 #(
		.INIT('ha8)
	) name7709 (
		\sa22_reg[2]/P0001 ,
		_w7543_,
		_w8241_,
		_w8242_
	);
	LUT4 #(
		.INIT('h0007)
	) name7710 (
		_w7008_,
		_w7520_,
		_w7544_,
		_w8230_,
		_w8243_
	);
	LUT2 #(
		.INIT('h4)
	) name7711 (
		_w8242_,
		_w8243_,
		_w8244_
	);
	LUT4 #(
		.INIT('h5540)
	) name7712 (
		\sa22_reg[2]/P0001 ,
		_w6943_,
		_w6945_,
		_w7229_,
		_w8245_
	);
	LUT2 #(
		.INIT('h8)
	) name7713 (
		_w7019_,
		_w7292_,
		_w8246_
	);
	LUT4 #(
		.INIT('h153f)
	) name7714 (
		_w6967_,
		_w6993_,
		_w6945_,
		_w7500_,
		_w8247_
	);
	LUT3 #(
		.INIT('h10)
	) name7715 (
		_w8245_,
		_w8246_,
		_w8247_,
		_w8248_
	);
	LUT4 #(
		.INIT('he400)
	) name7716 (
		\sa22_reg[1]/P0001 ,
		_w8244_,
		_w8240_,
		_w8248_,
		_w8249_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name7717 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w8250_
	);
	LUT2 #(
		.INIT('h2)
	) name7718 (
		_w7497_,
		_w8250_,
		_w8251_
	);
	LUT2 #(
		.INIT('h8)
	) name7719 (
		_w7227_,
		_w7520_,
		_w8252_
	);
	LUT4 #(
		.INIT('h2000)
	) name7720 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w8253_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7721 (
		\sa22_reg[2]/P0001 ,
		_w7008_,
		_w7277_,
		_w8253_,
		_w8254_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7722 (
		\sa22_reg[1]/P0001 ,
		_w8252_,
		_w8254_,
		_w8251_,
		_w8255_
	);
	LUT4 #(
		.INIT('h135f)
	) name7723 (
		_w6953_,
		_w6967_,
		_w6954_,
		_w7500_,
		_w8256_
	);
	LUT4 #(
		.INIT('hedff)
	) name7724 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w8257_
	);
	LUT2 #(
		.INIT('h2)
	) name7725 (
		_w7292_,
		_w8257_,
		_w8258_
	);
	LUT4 #(
		.INIT('h153f)
	) name7726 (
		_w6936_,
		_w7022_,
		_w7271_,
		_w7500_,
		_w8259_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7727 (
		_w7857_,
		_w8256_,
		_w8258_,
		_w8259_,
		_w8260_
	);
	LUT2 #(
		.INIT('h4)
	) name7728 (
		_w8255_,
		_w8260_,
		_w8261_
	);
	LUT4 #(
		.INIT('h0e00)
	) name7729 (
		\sa22_reg[0]/P0001 ,
		_w8249_,
		_w8236_,
		_w8261_,
		_w8262_
	);
	LUT4 #(
		.INIT('hefdf)
	) name7730 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8263_
	);
	LUT2 #(
		.INIT('h1)
	) name7731 (
		\sa33_reg[2]/P0001 ,
		_w8263_,
		_w8264_
	);
	LUT3 #(
		.INIT('h01)
	) name7732 (
		_w7131_,
		_w7307_,
		_w7962_,
		_w8265_
	);
	LUT4 #(
		.INIT('h0020)
	) name7733 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8266_
	);
	LUT4 #(
		.INIT('h0777)
	) name7734 (
		_w7080_,
		_w7039_,
		_w7126_,
		_w7138_,
		_w8267_
	);
	LUT4 #(
		.INIT('h1000)
	) name7735 (
		_w8266_,
		_w8264_,
		_w8265_,
		_w8267_,
		_w8268_
	);
	LUT4 #(
		.INIT('h2e00)
	) name7736 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8269_
	);
	LUT3 #(
		.INIT('ha8)
	) name7737 (
		\sa33_reg[2]/P0001 ,
		_w7078_,
		_w8269_,
		_w8270_
	);
	LUT4 #(
		.INIT('hffac)
	) name7738 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8271_
	);
	LUT2 #(
		.INIT('h1)
	) name7739 (
		\sa33_reg[2]/P0001 ,
		_w8271_,
		_w8272_
	);
	LUT3 #(
		.INIT('h13)
	) name7740 (
		_w7048_,
		_w7353_,
		_w7764_,
		_w8273_
	);
	LUT3 #(
		.INIT('h10)
	) name7741 (
		_w8270_,
		_w8272_,
		_w8273_,
		_w8274_
	);
	LUT4 #(
		.INIT('h0100)
	) name7742 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8275_
	);
	LUT4 #(
		.INIT('h000b)
	) name7743 (
		\sa33_reg[6]/P0001 ,
		_w7059_,
		_w7786_,
		_w8275_,
		_w8276_
	);
	LUT2 #(
		.INIT('h8)
	) name7744 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w8277_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name7745 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8278_
	);
	LUT4 #(
		.INIT('h7707)
	) name7746 (
		_w7033_,
		_w7056_,
		_w8277_,
		_w8278_,
		_w8279_
	);
	LUT3 #(
		.INIT('he0)
	) name7747 (
		\sa33_reg[2]/P0001 ,
		_w8276_,
		_w8279_,
		_w8280_
	);
	LUT4 #(
		.INIT('he400)
	) name7748 (
		\sa33_reg[1]/P0001 ,
		_w8268_,
		_w8274_,
		_w8280_,
		_w8281_
	);
	LUT3 #(
		.INIT('h01)
	) name7749 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8282_
	);
	LUT4 #(
		.INIT('haa80)
	) name7750 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7134_,
		_w8282_,
		_w8283_
	);
	LUT2 #(
		.INIT('h4)
	) name7751 (
		\sa33_reg[2]/P0001 ,
		_w7093_,
		_w8284_
	);
	LUT4 #(
		.INIT('h0a02)
	) name7752 (
		\sa33_reg[1]/P0001 ,
		_w7110_,
		_w7054_,
		_w7349_,
		_w8285_
	);
	LUT3 #(
		.INIT('h10)
	) name7753 (
		_w8283_,
		_w8284_,
		_w8285_,
		_w8286_
	);
	LUT4 #(
		.INIT('h0015)
	) name7754 (
		\sa33_reg[1]/P0001 ,
		_w7113_,
		_w7119_,
		_w8275_,
		_w8287_
	);
	LUT3 #(
		.INIT('h73)
	) name7755 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		_w8288_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7756 (
		_w7044_,
		_w7055_,
		_w7332_,
		_w8288_,
		_w8289_
	);
	LUT2 #(
		.INIT('h8)
	) name7757 (
		_w8287_,
		_w8289_,
		_w8290_
	);
	LUT3 #(
		.INIT('h07)
	) name7758 (
		_w7048_,
		_w7050_,
		_w7305_,
		_w8291_
	);
	LUT4 #(
		.INIT('h5540)
	) name7759 (
		\sa33_reg[2]/P0001 ,
		_w7048_,
		_w7050_,
		_w7305_,
		_w8292_
	);
	LUT3 #(
		.INIT('h02)
	) name7760 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8293_
	);
	LUT2 #(
		.INIT('h8)
	) name7761 (
		_w7924_,
		_w8293_,
		_w8294_
	);
	LUT4 #(
		.INIT('h135f)
	) name7762 (
		_w7066_,
		_w7110_,
		_w7067_,
		_w7335_,
		_w8295_
	);
	LUT3 #(
		.INIT('h10)
	) name7763 (
		_w8292_,
		_w8294_,
		_w8295_,
		_w8296_
	);
	LUT3 #(
		.INIT('he0)
	) name7764 (
		_w8286_,
		_w8290_,
		_w8296_,
		_w8297_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name7765 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8298_
	);
	LUT2 #(
		.INIT('h2)
	) name7766 (
		_w7928_,
		_w8298_,
		_w8299_
	);
	LUT4 #(
		.INIT('hd5df)
	) name7767 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8300_
	);
	LUT2 #(
		.INIT('h2)
	) name7768 (
		_w7306_,
		_w8300_,
		_w8301_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name7769 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		_w7119_,
		_w7980_,
		_w8302_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7770 (
		\sa33_reg[1]/P0001 ,
		_w8301_,
		_w8299_,
		_w8302_,
		_w8303_
	);
	LUT4 #(
		.INIT('haebf)
	) name7771 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7062_,
		_w7067_,
		_w8304_
	);
	LUT3 #(
		.INIT('hc8)
	) name7772 (
		_w7114_,
		_w7339_,
		_w7943_,
		_w8305_
	);
	LUT4 #(
		.INIT('h13ff)
	) name7773 (
		\sa33_reg[4]/P0001 ,
		_w7116_,
		_w7126_,
		_w7138_,
		_w8306_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7774 (
		_w7810_,
		_w8304_,
		_w8305_,
		_w8306_,
		_w8307_
	);
	LUT2 #(
		.INIT('h4)
	) name7775 (
		_w8303_,
		_w8307_,
		_w8308_
	);
	LUT4 #(
		.INIT('hd800)
	) name7776 (
		\sa33_reg[0]/P0001 ,
		_w8281_,
		_w8297_,
		_w8308_,
		_w8309_
	);
	LUT4 #(
		.INIT('h6996)
	) name7777 (
		\u0_w_reg[0][27]/P0001 ,
		_w8218_,
		_w8262_,
		_w8309_,
		_w8310_
	);
	LUT3 #(
		.INIT('h01)
	) name7778 (
		_w6731_,
		_w6698_,
		_w6687_,
		_w8311_
	);
	LUT3 #(
		.INIT('h15)
	) name7779 (
		_w6643_,
		_w6664_,
		_w6665_,
		_w8312_
	);
	LUT3 #(
		.INIT('h0e)
	) name7780 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		_w8313_
	);
	LUT4 #(
		.INIT('h1101)
	) name7781 (
		\sa11_reg[1]/P0001 ,
		_w6709_,
		_w6893_,
		_w8313_,
		_w8314_
	);
	LUT3 #(
		.INIT('h80)
	) name7782 (
		_w8311_,
		_w8312_,
		_w8314_,
		_w8315_
	);
	LUT4 #(
		.INIT('hbbf3)
	) name7783 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w8316_
	);
	LUT2 #(
		.INIT('h1)
	) name7784 (
		\sa11_reg[2]/P0001 ,
		_w8316_,
		_w8317_
	);
	LUT4 #(
		.INIT('h0002)
	) name7785 (
		\sa11_reg[2]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8318_
	);
	LUT4 #(
		.INIT('h002a)
	) name7786 (
		\sa11_reg[1]/P0001 ,
		_w6712_,
		_w7645_,
		_w8318_,
		_w8319_
	);
	LUT2 #(
		.INIT('h4)
	) name7787 (
		_w8317_,
		_w8319_,
		_w8320_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name7788 (
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8321_
	);
	LUT2 #(
		.INIT('h2)
	) name7789 (
		_w6730_,
		_w8321_,
		_w8322_
	);
	LUT3 #(
		.INIT('ha8)
	) name7790 (
		\sa11_reg[5]/P0001 ,
		_w6731_,
		_w6719_,
		_w8323_
	);
	LUT3 #(
		.INIT('h8a)
	) name7791 (
		\sa11_reg[0]/P0001 ,
		\sa11_reg[3]/P0001 ,
		_w6638_,
		_w8324_
	);
	LUT3 #(
		.INIT('h10)
	) name7792 (
		_w8322_,
		_w8323_,
		_w8324_,
		_w8325_
	);
	LUT3 #(
		.INIT('he0)
	) name7793 (
		_w8315_,
		_w8320_,
		_w8325_,
		_w8326_
	);
	LUT4 #(
		.INIT('hffda)
	) name7794 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8327_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7795 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[2]/P0001 ,
		_w7684_,
		_w8327_,
		_w8328_
	);
	LUT3 #(
		.INIT('h54)
	) name7796 (
		\sa11_reg[1]/P0001 ,
		_w7645_,
		_w7637_,
		_w8329_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name7797 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8330_
	);
	LUT4 #(
		.INIT('h3f1d)
	) name7798 (
		\sa11_reg[1]/P0001 ,
		_w6666_,
		_w6694_,
		_w8330_,
		_w8331_
	);
	LUT4 #(
		.INIT('h0105)
	) name7799 (
		\sa11_reg[0]/P0001 ,
		_w6730_,
		_w6704_,
		_w6910_,
		_w8332_
	);
	LUT4 #(
		.INIT('h0e00)
	) name7800 (
		\sa11_reg[2]/P0001 ,
		_w8331_,
		_w8329_,
		_w8332_,
		_w8333_
	);
	LUT2 #(
		.INIT('h4)
	) name7801 (
		_w8328_,
		_w8333_,
		_w8334_
	);
	LUT3 #(
		.INIT('h01)
	) name7802 (
		_w6667_,
		_w6677_,
		_w7477_,
		_w8335_
	);
	LUT3 #(
		.INIT('h02)
	) name7803 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w8336_
	);
	LUT3 #(
		.INIT('h07)
	) name7804 (
		_w6634_,
		_w6681_,
		_w8336_,
		_w8337_
	);
	LUT4 #(
		.INIT('h135f)
	) name7805 (
		_w7690_,
		_w7697_,
		_w8335_,
		_w8337_,
		_w8338_
	);
	LUT4 #(
		.INIT('h000b)
	) name7806 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		_w8339_
	);
	LUT2 #(
		.INIT('h4)
	) name7807 (
		_w7447_,
		_w8339_,
		_w8340_
	);
	LUT3 #(
		.INIT('h54)
	) name7808 (
		\sa11_reg[1]/P0001 ,
		_w8338_,
		_w8340_,
		_w8341_
	);
	LUT4 #(
		.INIT('h0400)
	) name7809 (
		\sa11_reg[3]/P0001 ,
		\sa11_reg[4]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8342_
	);
	LUT4 #(
		.INIT('h0007)
	) name7810 (
		_w6879_,
		_w6847_,
		_w6896_,
		_w8342_,
		_w8343_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name7811 (
		\sa11_reg[1]/P0001 ,
		\sa11_reg[2]/P0001 ,
		_w6680_,
		_w8343_,
		_w8344_
	);
	LUT4 #(
		.INIT('h0013)
	) name7812 (
		_w6634_,
		_w6725_,
		_w6861_,
		_w6910_,
		_w8345_
	);
	LUT3 #(
		.INIT('had)
	) name7813 (
		\sa11_reg[5]/P0001 ,
		\sa11_reg[6]/NET0131 ,
		\sa11_reg[7]/NET0131 ,
		_w8346_
	);
	LUT4 #(
		.INIT('h7707)
	) name7814 (
		_w6707_,
		_w6714_,
		_w7650_,
		_w8346_,
		_w8347_
	);
	LUT3 #(
		.INIT('hd0)
	) name7815 (
		_w7480_,
		_w8345_,
		_w8347_,
		_w8348_
	);
	LUT2 #(
		.INIT('h4)
	) name7816 (
		_w8344_,
		_w8348_,
		_w8349_
	);
	LUT4 #(
		.INIT('h5400)
	) name7817 (
		_w8341_,
		_w8326_,
		_w8334_,
		_w8349_,
		_w8350_
	);
	LUT3 #(
		.INIT('h54)
	) name7818 (
		\sa00_reg[2]/P0001 ,
		_w7214_,
		_w7208_,
		_w8351_
	);
	LUT4 #(
		.INIT('h0020)
	) name7819 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8352_
	);
	LUT4 #(
		.INIT('h0001)
	) name7820 (
		_w6799_,
		_w6751_,
		_w8096_,
		_w8352_,
		_w8353_
	);
	LUT3 #(
		.INIT('h01)
	) name7821 (
		\sa00_reg[1]/P0001 ,
		_w6808_,
		_w6785_,
		_w8354_
	);
	LUT3 #(
		.INIT('h40)
	) name7822 (
		_w8351_,
		_w8353_,
		_w8354_,
		_w8355_
	);
	LUT4 #(
		.INIT('hbbf3)
	) name7823 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w8356_
	);
	LUT2 #(
		.INIT('h1)
	) name7824 (
		\sa00_reg[2]/P0001 ,
		_w8356_,
		_w8357_
	);
	LUT4 #(
		.INIT('h0002)
	) name7825 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8358_
	);
	LUT4 #(
		.INIT('h002a)
	) name7826 (
		\sa00_reg[1]/P0001 ,
		_w7385_,
		_w7402_,
		_w8358_,
		_w8359_
	);
	LUT2 #(
		.INIT('h4)
	) name7827 (
		_w8357_,
		_w8359_,
		_w8360_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name7828 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8361_
	);
	LUT2 #(
		.INIT('h2)
	) name7829 (
		_w6831_,
		_w8361_,
		_w8362_
	);
	LUT2 #(
		.INIT('h8)
	) name7830 (
		_w6832_,
		_w7186_,
		_w8363_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name7831 (
		\sa00_reg[6]/NET0131 ,
		_w6769_,
		_w6770_,
		_w6783_,
		_w8364_
	);
	LUT3 #(
		.INIT('h10)
	) name7832 (
		_w8363_,
		_w8362_,
		_w8364_,
		_w8365_
	);
	LUT4 #(
		.INIT('h02aa)
	) name7833 (
		\sa00_reg[0]/P0001 ,
		_w8355_,
		_w8360_,
		_w8365_,
		_w8366_
	);
	LUT3 #(
		.INIT('h07)
	) name7834 (
		_w6738_,
		_w6788_,
		_w6781_,
		_w8367_
	);
	LUT4 #(
		.INIT('h0015)
	) name7835 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w6749_,
		_w8152_,
		_w8368_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name7836 (
		_w7421_,
		_w8161_,
		_w8367_,
		_w8368_,
		_w8369_
	);
	LUT4 #(
		.INIT('h000b)
	) name7837 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w8370_
	);
	LUT2 #(
		.INIT('h4)
	) name7838 (
		_w6818_,
		_w8370_,
		_w8371_
	);
	LUT3 #(
		.INIT('h15)
	) name7839 (
		\sa00_reg[1]/P0001 ,
		_w6805_,
		_w6770_,
		_w8372_
	);
	LUT2 #(
		.INIT('h4)
	) name7840 (
		_w8371_,
		_w8372_,
		_w8373_
	);
	LUT4 #(
		.INIT('h0007)
	) name7841 (
		_w6748_,
		_w6788_,
		_w7166_,
		_w7175_,
		_w8374_
	);
	LUT2 #(
		.INIT('h2)
	) name7842 (
		\sa00_reg[1]/P0001 ,
		_w6771_,
		_w8375_
	);
	LUT3 #(
		.INIT('he0)
	) name7843 (
		\sa00_reg[2]/P0001 ,
		_w8374_,
		_w8375_,
		_w8376_
	);
	LUT3 #(
		.INIT('h0b)
	) name7844 (
		_w8369_,
		_w8373_,
		_w8376_,
		_w8377_
	);
	LUT4 #(
		.INIT('hffda)
	) name7845 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8378_
	);
	LUT2 #(
		.INIT('h2)
	) name7846 (
		\sa00_reg[2]/P0001 ,
		_w8378_,
		_w8379_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name7847 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8380_
	);
	LUT3 #(
		.INIT('h51)
	) name7848 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w8381_
	);
	LUT3 #(
		.INIT('h45)
	) name7849 (
		_w7414_,
		_w8380_,
		_w8381_,
		_w8382_
	);
	LUT3 #(
		.INIT('h8a)
	) name7850 (
		\sa00_reg[1]/P0001 ,
		_w8379_,
		_w8382_,
		_w8383_
	);
	LUT4 #(
		.INIT('h0040)
	) name7851 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w8384_
	);
	LUT3 #(
		.INIT('h54)
	) name7852 (
		\sa00_reg[1]/P0001 ,
		_w8158_,
		_w8384_,
		_w8385_
	);
	LUT3 #(
		.INIT('h15)
	) name7853 (
		_w6802_,
		_w7387_,
		_w8081_,
		_w8386_
	);
	LUT3 #(
		.INIT('h10)
	) name7854 (
		_w7424_,
		_w8385_,
		_w8386_,
		_w8387_
	);
	LUT3 #(
		.INIT('h80)
	) name7855 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		_w8388_
	);
	LUT3 #(
		.INIT('had)
	) name7856 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8389_
	);
	LUT4 #(
		.INIT('h5f13)
	) name7857 (
		_w6839_,
		_w8111_,
		_w8388_,
		_w8389_,
		_w8390_
	);
	LUT4 #(
		.INIT('he2ee)
	) name7858 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w8391_
	);
	LUT3 #(
		.INIT('h80)
	) name7859 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[2]/P0001 ,
		\sa00_reg[7]/NET0131 ,
		_w8392_
	);
	LUT4 #(
		.INIT('h7077)
	) name7860 (
		_w6742_,
		_w7402_,
		_w8391_,
		_w8392_,
		_w8393_
	);
	LUT2 #(
		.INIT('h8)
	) name7861 (
		_w8390_,
		_w8393_,
		_w8394_
	);
	LUT4 #(
		.INIT('hba00)
	) name7862 (
		\sa00_reg[0]/P0001 ,
		_w8383_,
		_w8387_,
		_w8394_,
		_w8395_
	);
	LUT3 #(
		.INIT('h10)
	) name7863 (
		_w8377_,
		_w8366_,
		_w8395_,
		_w8396_
	);
	LUT4 #(
		.INIT('h9669)
	) name7864 (
		_w7706_,
		_w8169_,
		_w8350_,
		_w8396_,
		_w8397_
	);
	LUT3 #(
		.INIT('h82)
	) name7865 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[123]/P0001 ,
		\u0_w_reg[0][27]/P0001 ,
		_w8398_
	);
	LUT4 #(
		.INIT('h00be)
	) name7866 (
		\ld_r_reg/P0001 ,
		_w8310_,
		_w8397_,
		_w8398_,
		_w8399_
	);
	LUT4 #(
		.INIT('h6996)
	) name7867 (
		\u0_w_reg[0][19]/P0001 ,
		_w7908_,
		_w8262_,
		_w8309_,
		_w8400_
	);
	LUT4 #(
		.INIT('h0103)
	) name7868 (
		_w7000_,
		_w7230_,
		_w7256_,
		_w7497_,
		_w8401_
	);
	LUT4 #(
		.INIT('h0020)
	) name7869 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w8402_
	);
	LUT4 #(
		.INIT('h0001)
	) name7870 (
		_w7265_,
		_w7271_,
		_w7561_,
		_w8402_,
		_w8403_
	);
	LUT4 #(
		.INIT('h4555)
	) name7871 (
		\sa22_reg[1]/P0001 ,
		_w6960_,
		_w8403_,
		_w8401_,
		_w8404_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name7872 (
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w8405_
	);
	LUT2 #(
		.INIT('h2)
	) name7873 (
		_w7292_,
		_w8405_,
		_w8406_
	);
	LUT4 #(
		.INIT('hbbf3)
	) name7874 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		_w8407_
	);
	LUT4 #(
		.INIT('h1500)
	) name7875 (
		\sa22_reg[2]/P0001 ,
		_w6921_,
		_w6946_,
		_w8407_,
		_w8408_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7876 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w8409_
	);
	LUT2 #(
		.INIT('h2)
	) name7877 (
		\sa22_reg[1]/P0001 ,
		_w8409_,
		_w8410_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name7878 (
		\sa22_reg[3]/P0001 ,
		_w6953_,
		_w7023_,
		_w7240_,
		_w8411_
	);
	LUT4 #(
		.INIT('h4500)
	) name7879 (
		_w7819_,
		_w8408_,
		_w8410_,
		_w8411_,
		_w8412_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7880 (
		\sa22_reg[0]/P0001 ,
		_w8404_,
		_w8406_,
		_w8412_,
		_w8413_
	);
	LUT3 #(
		.INIT('h10)
	) name7881 (
		_w7019_,
		_w7249_,
		_w7566_,
		_w8414_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7882 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w8415_
	);
	LUT2 #(
		.INIT('h4)
	) name7883 (
		_w6930_,
		_w8415_,
		_w8416_
	);
	LUT4 #(
		.INIT('h888a)
	) name7884 (
		\sa22_reg[1]/P0001 ,
		_w7532_,
		_w8414_,
		_w8416_,
		_w8417_
	);
	LUT4 #(
		.INIT('h0040)
	) name7885 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		\sa22_reg[5]/P0001 ,
		\sa22_reg[7]/NET0131 ,
		_w8418_
	);
	LUT3 #(
		.INIT('h54)
	) name7886 (
		\sa22_reg[1]/P0001 ,
		_w7592_,
		_w8418_,
		_w8419_
	);
	LUT3 #(
		.INIT('h80)
	) name7887 (
		\sa22_reg[2]/P0001 ,
		_w6923_,
		_w7287_,
		_w8420_
	);
	LUT3 #(
		.INIT('h15)
	) name7888 (
		_w7008_,
		_w7240_,
		_w7520_,
		_w8421_
	);
	LUT3 #(
		.INIT('h10)
	) name7889 (
		_w8420_,
		_w8419_,
		_w8421_,
		_w8422_
	);
	LUT3 #(
		.INIT('h45)
	) name7890 (
		\sa22_reg[0]/P0001 ,
		_w8417_,
		_w8422_,
		_w8423_
	);
	LUT4 #(
		.INIT('h0400)
	) name7891 (
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w8424_
	);
	LUT4 #(
		.INIT('h0007)
	) name7892 (
		\sa22_reg[6]/NET0131 ,
		_w6986_,
		_w7003_,
		_w8424_,
		_w8425_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name7893 (
		\sa22_reg[1]/P0001 ,
		\sa22_reg[2]/P0001 ,
		_w6981_,
		_w8425_,
		_w8426_
	);
	LUT4 #(
		.INIT('h0007)
	) name7894 (
		_w6929_,
		_w6985_,
		_w7240_,
		_w7537_,
		_w8427_
	);
	LUT4 #(
		.INIT('h0015)
	) name7895 (
		_w6977_,
		_w6982_,
		_w7249_,
		_w7592_,
		_w8428_
	);
	LUT4 #(
		.INIT('h0013)
	) name7896 (
		_w6951_,
		_w7227_,
		_w7497_,
		_w7901_,
		_w8429_
	);
	LUT4 #(
		.INIT('hd800)
	) name7897 (
		\sa22_reg[2]/P0001 ,
		_w8428_,
		_w8427_,
		_w8429_,
		_w8430_
	);
	LUT4 #(
		.INIT('h0103)
	) name7898 (
		_w6921_,
		_w6959_,
		_w7023_,
		_w7500_,
		_w8431_
	);
	LUT3 #(
		.INIT('had)
	) name7899 (
		\sa22_reg[5]/P0001 ,
		\sa22_reg[6]/NET0131 ,
		\sa22_reg[7]/NET0131 ,
		_w8432_
	);
	LUT3 #(
		.INIT('h02)
	) name7900 (
		\sa22_reg[2]/P0001 ,
		\sa22_reg[3]/P0001 ,
		\sa22_reg[4]/P0001 ,
		_w8433_
	);
	LUT4 #(
		.INIT('h7077)
	) name7901 (
		_w7227_,
		_w7520_,
		_w8432_,
		_w8433_,
		_w8434_
	);
	LUT3 #(
		.INIT('hd0)
	) name7902 (
		_w7540_,
		_w8431_,
		_w8434_,
		_w8435_
	);
	LUT4 #(
		.INIT('h3200)
	) name7903 (
		\sa22_reg[1]/P0001 ,
		_w8426_,
		_w8430_,
		_w8435_,
		_w8436_
	);
	LUT3 #(
		.INIT('h10)
	) name7904 (
		_w8423_,
		_w8413_,
		_w8436_,
		_w8437_
	);
	LUT4 #(
		.INIT('h2e00)
	) name7905 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8438_
	);
	LUT3 #(
		.INIT('ha8)
	) name7906 (
		\sa00_reg[2]/P0001 ,
		_w7757_,
		_w8438_,
		_w8439_
	);
	LUT3 #(
		.INIT('h01)
	) name7907 (
		_w6802_,
		_w6817_,
		_w8158_,
		_w8440_
	);
	LUT4 #(
		.INIT('h0010)
	) name7908 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8441_
	);
	LUT2 #(
		.INIT('h1)
	) name7909 (
		_w8101_,
		_w8441_,
		_w8442_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name7910 (
		\sa00_reg[1]/P0001 ,
		_w8439_,
		_w8440_,
		_w8442_,
		_w8443_
	);
	LUT4 #(
		.INIT('hfd3f)
	) name7911 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8444_
	);
	LUT3 #(
		.INIT('h8a)
	) name7912 (
		\sa00_reg[2]/P0001 ,
		_w8116_,
		_w8444_,
		_w8445_
	);
	LUT4 #(
		.INIT('hefdf)
	) name7913 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8446_
	);
	LUT2 #(
		.INIT('h1)
	) name7914 (
		\sa00_reg[2]/P0001 ,
		_w8446_,
		_w8447_
	);
	LUT4 #(
		.INIT('h0007)
	) name7915 (
		_w6780_,
		_w6781_,
		_w7214_,
		_w7418_,
		_w8448_
	);
	LUT4 #(
		.INIT('h5455)
	) name7916 (
		\sa00_reg[1]/P0001 ,
		_w8447_,
		_w8445_,
		_w8448_,
		_w8449_
	);
	LUT4 #(
		.INIT('h0013)
	) name7917 (
		_w6780_,
		_w6783_,
		_w7757_,
		_w8084_,
		_w8450_
	);
	LUT4 #(
		.INIT('hf4cf)
	) name7918 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8451_
	);
	LUT2 #(
		.INIT('h8)
	) name7919 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[4]/P0001 ,
		_w8452_
	);
	LUT4 #(
		.INIT('h7077)
	) name7920 (
		_w6738_,
		_w7186_,
		_w8451_,
		_w8452_,
		_w8453_
	);
	LUT3 #(
		.INIT('he0)
	) name7921 (
		\sa00_reg[2]/P0001 ,
		_w8450_,
		_w8453_,
		_w8454_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7922 (
		\sa00_reg[0]/P0001 ,
		_w8449_,
		_w8443_,
		_w8454_,
		_w8455_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name7923 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w7170_,
		_w7396_,
		_w8456_
	);
	LUT3 #(
		.INIT('h13)
	) name7924 (
		\sa00_reg[5]/P0001 ,
		_w6813_,
		_w6823_,
		_w8457_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name7925 (
		\sa00_reg[2]/P0001 ,
		_w6748_,
		_w6788_,
		_w7159_,
		_w8458_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name7926 (
		\sa00_reg[1]/P0001 ,
		_w8456_,
		_w8457_,
		_w8458_,
		_w8459_
	);
	LUT3 #(
		.INIT('h13)
	) name7927 (
		_w6802_,
		_w6783_,
		_w7402_,
		_w8460_
	);
	LUT3 #(
		.INIT('he0)
	) name7928 (
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8461_
	);
	LUT4 #(
		.INIT('h23af)
	) name7929 (
		_w6805_,
		_w6832_,
		_w6764_,
		_w8461_,
		_w8462_
	);
	LUT3 #(
		.INIT('h15)
	) name7930 (
		\sa00_reg[1]/P0001 ,
		_w8460_,
		_w8462_,
		_w8463_
	);
	LUT4 #(
		.INIT('h5540)
	) name7931 (
		\sa00_reg[2]/P0001 ,
		_w6745_,
		_w6788_,
		_w6749_,
		_w8464_
	);
	LUT2 #(
		.INIT('h8)
	) name7932 (
		_w6831_,
		_w7170_,
		_w8465_
	);
	LUT4 #(
		.INIT('h47cf)
	) name7933 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w7152_,
		_w7419_,
		_w8466_
	);
	LUT3 #(
		.INIT('h10)
	) name7934 (
		_w8465_,
		_w8464_,
		_w8466_,
		_w8467_
	);
	LUT4 #(
		.INIT('h5455)
	) name7935 (
		\sa00_reg[0]/P0001 ,
		_w8459_,
		_w8463_,
		_w8467_,
		_w8468_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name7936 (
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		\sa00_reg[7]/NET0131 ,
		_w8469_
	);
	LUT2 #(
		.INIT('h2)
	) name7937 (
		_w8079_,
		_w8469_,
		_w8470_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name7938 (
		\sa00_reg[2]/P0001 ,
		\sa00_reg[3]/P0001 ,
		_w6802_,
		_w6742_,
		_w8471_
	);
	LUT3 #(
		.INIT('h8a)
	) name7939 (
		\sa00_reg[1]/P0001 ,
		_w8470_,
		_w8471_,
		_w8472_
	);
	LUT4 #(
		.INIT('h2000)
	) name7940 (
		\sa00_reg[3]/P0001 ,
		\sa00_reg[4]/P0001 ,
		\sa00_reg[5]/P0001 ,
		\sa00_reg[6]/NET0131 ,
		_w8473_
	);
	LUT3 #(
		.INIT('hc8)
	) name7941 (
		_w6817_,
		_w7738_,
		_w8473_,
		_w8474_
	);
	LUT4 #(
		.INIT('haabf)
	) name7942 (
		\sa00_reg[5]/P0001 ,
		_w6745_,
		_w6758_,
		_w7152_,
		_w8475_
	);
	LUT3 #(
		.INIT('h1d)
	) name7943 (
		\sa00_reg[1]/P0001 ,
		\sa00_reg[2]/P0001 ,
		\sa00_reg[5]/P0001 ,
		_w8476_
	);
	LUT4 #(
		.INIT('h135f)
	) name7944 (
		\sa00_reg[4]/P0001 ,
		_w6808_,
		_w7727_,
		_w8476_,
		_w8477_
	);
	LUT4 #(
		.INIT('h3100)
	) name7945 (
		_w7389_,
		_w7755_,
		_w8475_,
		_w8477_,
		_w8478_
	);
	LUT3 #(
		.INIT('h10)
	) name7946 (
		_w8472_,
		_w8474_,
		_w8478_,
		_w8479_
	);
	LUT3 #(
		.INIT('h10)
	) name7947 (
		_w8468_,
		_w8455_,
		_w8479_,
		_w8480_
	);
	LUT4 #(
		.INIT('h6996)
	) name7948 (
		_w7706_,
		_w8350_,
		_w8437_,
		_w8480_,
		_w8481_
	);
	LUT3 #(
		.INIT('h82)
	) name7949 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[115]/P0001 ,
		\u0_w_reg[0][19]/P0001 ,
		_w8482_
	);
	LUT4 #(
		.INIT('h00eb)
	) name7950 (
		\ld_r_reg/P0001 ,
		_w8400_,
		_w8481_,
		_w8482_,
		_w8483_
	);
	LUT4 #(
		.INIT('h6996)
	) name7951 (
		_w7908_,
		_w8218_,
		_w8437_,
		_w8480_,
		_w8484_
	);
	LUT3 #(
		.INIT('h2a)
	) name7952 (
		\sa33_reg[1]/P0001 ,
		_w7088_,
		_w7113_,
		_w8485_
	);
	LUT4 #(
		.INIT('h0002)
	) name7953 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8486_
	);
	LUT3 #(
		.INIT('h07)
	) name7954 (
		_w7764_,
		_w7984_,
		_w8486_,
		_w8487_
	);
	LUT2 #(
		.INIT('h8)
	) name7955 (
		_w8485_,
		_w8487_,
		_w8488_
	);
	LUT4 #(
		.INIT('h000b)
	) name7956 (
		\sa33_reg[2]/P0001 ,
		_w7070_,
		_w7336_,
		_w7976_,
		_w8489_
	);
	LUT3 #(
		.INIT('h01)
	) name7957 (
		\sa33_reg[1]/P0001 ,
		_w7340_,
		_w7321_,
		_w8490_
	);
	LUT3 #(
		.INIT('h08)
	) name7958 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8491_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name7959 (
		_w7053_,
		_w7344_,
		_w7916_,
		_w8491_,
		_w8492_
	);
	LUT3 #(
		.INIT('h80)
	) name7960 (
		_w8489_,
		_w8490_,
		_w8492_,
		_w8493_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name7961 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8494_
	);
	LUT2 #(
		.INIT('h2)
	) name7962 (
		_w7138_,
		_w8494_,
		_w8495_
	);
	LUT3 #(
		.INIT('h2a)
	) name7963 (
		\sa33_reg[0]/P0001 ,
		_w7066_,
		_w7139_,
		_w8496_
	);
	LUT4 #(
		.INIT('h135f)
	) name7964 (
		_w7055_,
		_w7107_,
		_w7056_,
		_w7123_,
		_w8497_
	);
	LUT3 #(
		.INIT('h40)
	) name7965 (
		_w8495_,
		_w8496_,
		_w8497_,
		_w8498_
	);
	LUT3 #(
		.INIT('he0)
	) name7966 (
		_w8488_,
		_w8493_,
		_w8498_,
		_w8499_
	);
	LUT4 #(
		.INIT('hffda)
	) name7967 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8500_
	);
	LUT2 #(
		.INIT('h2)
	) name7968 (
		\sa33_reg[2]/P0001 ,
		_w8500_,
		_w8501_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name7969 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8502_
	);
	LUT3 #(
		.INIT('h51)
	) name7970 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8503_
	);
	LUT4 #(
		.INIT('h2022)
	) name7971 (
		\sa33_reg[1]/P0001 ,
		_w7793_,
		_w8502_,
		_w8503_,
		_w8504_
	);
	LUT4 #(
		.INIT('h0040)
	) name7972 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8505_
	);
	LUT3 #(
		.INIT('h01)
	) name7973 (
		\sa33_reg[1]/P0001 ,
		_w7059_,
		_w8505_,
		_w8506_
	);
	LUT3 #(
		.INIT('h0b)
	) name7974 (
		_w8501_,
		_w8504_,
		_w8506_,
		_w8507_
	);
	LUT2 #(
		.INIT('h8)
	) name7975 (
		_w7353_,
		_w8277_,
		_w8508_
	);
	LUT4 #(
		.INIT('h0111)
	) name7976 (
		\sa33_reg[0]/P0001 ,
		_w7119_,
		_w7142_,
		_w7342_,
		_w8509_
	);
	LUT2 #(
		.INIT('h4)
	) name7977 (
		_w8508_,
		_w8509_,
		_w8510_
	);
	LUT2 #(
		.INIT('h4)
	) name7978 (
		_w8507_,
		_w8510_,
		_w8511_
	);
	LUT4 #(
		.INIT('h0800)
	) name7979 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8512_
	);
	LUT3 #(
		.INIT('h01)
	) name7980 (
		\sa33_reg[2]/P0001 ,
		_w7953_,
		_w8512_,
		_w8513_
	);
	LUT3 #(
		.INIT('h07)
	) name7981 (
		\sa33_reg[6]/P0001 ,
		_w7063_,
		_w7321_,
		_w8514_
	);
	LUT4 #(
		.INIT('haaa2)
	) name7982 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w8515_
	);
	LUT4 #(
		.INIT('h0700)
	) name7983 (
		_w7033_,
		_w7110_,
		_w7059_,
		_w8515_,
		_w8516_
	);
	LUT3 #(
		.INIT('h01)
	) name7984 (
		\sa33_reg[1]/P0001 ,
		_w7963_,
		_w7980_,
		_w8517_
	);
	LUT4 #(
		.INIT('hf800)
	) name7985 (
		_w8513_,
		_w8514_,
		_w8516_,
		_w8517_,
		_w8518_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name7986 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[5]/P0001 ,
		_w7938_,
		_w8293_,
		_w8519_
	);
	LUT2 #(
		.INIT('h2)
	) name7987 (
		\sa33_reg[6]/P0001 ,
		_w8519_,
		_w8520_
	);
	LUT3 #(
		.INIT('ha8)
	) name7988 (
		\sa33_reg[2]/P0001 ,
		_w7070_,
		_w7123_,
		_w8521_
	);
	LUT3 #(
		.INIT('h8a)
	) name7989 (
		\sa33_reg[1]/P0001 ,
		\sa33_reg[2]/P0001 ,
		_w7116_,
		_w8522_
	);
	LUT3 #(
		.INIT('h13)
	) name7990 (
		_w7049_,
		_w7141_,
		_w7302_,
		_w8523_
	);
	LUT3 #(
		.INIT('h40)
	) name7991 (
		_w8521_,
		_w8522_,
		_w8523_,
		_w8524_
	);
	LUT3 #(
		.INIT('had)
	) name7992 (
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8525_
	);
	LUT3 #(
		.INIT('h02)
	) name7993 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[3]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w8526_
	);
	LUT4 #(
		.INIT('h7077)
	) name7994 (
		_w7113_,
		_w7980_,
		_w8525_,
		_w8526_,
		_w8527_
	);
	LUT4 #(
		.INIT('hba00)
	) name7995 (
		_w8518_,
		_w8520_,
		_w8524_,
		_w8527_,
		_w8528_
	);
	LUT4 #(
		.INIT('ha955)
	) name7996 (
		\u0_w_reg[0][11]/P0001 ,
		_w8499_,
		_w8511_,
		_w8528_,
		_w8529_
	);
	LUT3 #(
		.INIT('h69)
	) name7997 (
		_w7971_,
		_w8309_,
		_w8529_,
		_w8530_
	);
	LUT3 #(
		.INIT('h82)
	) name7998 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[107]/P0001 ,
		\u0_w_reg[0][11]/P0001 ,
		_w8531_
	);
	LUT4 #(
		.INIT('h00eb)
	) name7999 (
		\ld_r_reg/P0001 ,
		_w8484_,
		_w8530_,
		_w8531_,
		_w8532_
	);
	LUT4 #(
		.INIT('h6996)
	) name8000 (
		\u0_w_reg[0][12]/P0001 ,
		_w7367_,
		_w7971_,
		_w8309_,
		_w8533_
	);
	LUT4 #(
		.INIT('h6996)
	) name8001 (
		_w6737_,
		_w6842_,
		_w7908_,
		_w8262_,
		_w8534_
	);
	LUT3 #(
		.INIT('h82)
	) name8002 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[108]/P0001 ,
		\u0_w_reg[0][12]/P0001 ,
		_w8535_
	);
	LUT4 #(
		.INIT('h00eb)
	) name8003 (
		\ld_r_reg/P0001 ,
		_w8533_,
		_w8534_,
		_w8535_,
		_w8536_
	);
	LUT4 #(
		.INIT('h6996)
	) name8004 (
		\u0_w_reg[0][4]/P0001 ,
		_w7295_,
		_w7971_,
		_w8309_,
		_w8537_
	);
	LUT4 #(
		.INIT('h6996)
	) name8005 (
		_w6737_,
		_w6842_,
		_w8169_,
		_w8480_,
		_w8538_
	);
	LUT3 #(
		.INIT('h82)
	) name8006 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[100]/P0001 ,
		\u0_w_reg[0][4]/P0001 ,
		_w8539_
	);
	LUT4 #(
		.INIT('h00eb)
	) name8007 (
		\ld_r_reg/P0001 ,
		_w8537_,
		_w8538_,
		_w8539_,
		_w8540_
	);
	LUT4 #(
		.INIT('h6996)
	) name8008 (
		\u0_w_reg[0][25]/P0001 ,
		_w7817_,
		_w7865_,
		_w8068_,
		_w8541_
	);
	LUT4 #(
		.INIT('h9669)
	) name8009 (
		_w7655_,
		_w7706_,
		_w8123_,
		_w8169_,
		_w8542_
	);
	LUT3 #(
		.INIT('h28)
	) name8010 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[121]/P0001 ,
		\u0_w_reg[0][25]/P0001 ,
		_w8543_
	);
	LUT4 #(
		.INIT('hff14)
	) name8011 (
		\ld_r_reg/P0001 ,
		_w8541_,
		_w8542_,
		_w8543_,
		_w8544_
	);
	LUT4 #(
		.INIT('h6996)
	) name8012 (
		\u0_w_reg[0][28]/P0001 ,
		_w6737_,
		_w7295_,
		_w7367_,
		_w8545_
	);
	LUT4 #(
		.INIT('h9669)
	) name8013 (
		_w7706_,
		_w8169_,
		_w8218_,
		_w8480_,
		_w8546_
	);
	LUT3 #(
		.INIT('h82)
	) name8014 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[124]/P0001 ,
		\u0_w_reg[0][28]/P0001 ,
		_w8547_
	);
	LUT4 #(
		.INIT('h00be)
	) name8015 (
		\ld_r_reg/P0001 ,
		_w8545_,
		_w8546_,
		_w8547_,
		_w8548_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name8016 (
		\u0_w_reg[0][24]/P0001 ,
		_w7991_,
		_w8004_,
		_w8017_,
		_w8549_
	);
	LUT4 #(
		.INIT('h9669)
	) name8017 (
		_w7603_,
		_w7655_,
		_w7706_,
		_w8169_,
		_w8550_
	);
	LUT3 #(
		.INIT('h28)
	) name8018 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[120]/P0001 ,
		\u0_w_reg[0][24]/P0001 ,
		_w8551_
	);
	LUT4 #(
		.INIT('hff14)
	) name8019 (
		\ld_r_reg/P0001 ,
		_w8549_,
		_w8550_,
		_w8551_,
		_w8552_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name8020 (
		\u0_w_reg[0][16]/P0001 ,
		_w7991_,
		_w8004_,
		_w8017_,
		_w8553_
	);
	LUT4 #(
		.INIT('h6996)
	) name8021 (
		_w7603_,
		_w7706_,
		_w7908_,
		_w8123_,
		_w8554_
	);
	LUT3 #(
		.INIT('h28)
	) name8022 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[112]/P0001 ,
		\u0_w_reg[0][16]/P0001 ,
		_w8555_
	);
	LUT4 #(
		.INIT('hff41)
	) name8023 (
		\ld_r_reg/P0001 ,
		_w8553_,
		_w8554_,
		_w8555_,
		_w8556_
	);
	LUT4 #(
		.INIT('h6996)
	) name8024 (
		_w6842_,
		_w7706_,
		_w8218_,
		_w8262_,
		_w8557_
	);
	LUT4 #(
		.INIT('h5655)
	) name8025 (
		\u0_w_reg[0][20]/P0001 ,
		_w7893_,
		_w7880_,
		_w7907_,
		_w8558_
	);
	LUT3 #(
		.INIT('h96)
	) name8026 (
		_w7295_,
		_w7367_,
		_w8558_,
		_w8559_
	);
	LUT3 #(
		.INIT('h82)
	) name8027 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[116]/P0001 ,
		\u0_w_reg[0][20]/P0001 ,
		_w8560_
	);
	LUT4 #(
		.INIT('h00be)
	) name8028 (
		\ld_r_reg/P0001 ,
		_w8557_,
		_w8559_,
		_w8560_,
		_w8561_
	);
	LUT4 #(
		.INIT('hb44b)
	) name8029 (
		_w6867_,
		_w6920_,
		_w7031_,
		_w7433_,
		_w8562_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name8030 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8563_
	);
	LUT4 #(
		.INIT('h80aa)
	) name8031 (
		\sa33_reg[2]/P0001 ,
		_w7069_,
		_w7123_,
		_w8563_,
		_w8564_
	);
	LUT2 #(
		.INIT('h8)
	) name8032 (
		_w7763_,
		_w7928_,
		_w8565_
	);
	LUT4 #(
		.INIT('haaa2)
	) name8033 (
		\sa33_reg[1]/P0001 ,
		_w7979_,
		_w8565_,
		_w8564_,
		_w8566_
	);
	LUT3 #(
		.INIT('ha8)
	) name8034 (
		\sa33_reg[2]/P0001 ,
		_w7067_,
		_w7938_,
		_w8567_
	);
	LUT3 #(
		.INIT('h13)
	) name8035 (
		_w7078_,
		_w7119_,
		_w7342_,
		_w8568_
	);
	LUT4 #(
		.INIT('h5155)
	) name8036 (
		\sa33_reg[1]/P0001 ,
		_w7117_,
		_w8567_,
		_w8568_,
		_w8569_
	);
	LUT3 #(
		.INIT('h54)
	) name8037 (
		\sa33_reg[2]/P0001 ,
		_w7088_,
		_w7079_,
		_w8570_
	);
	LUT2 #(
		.INIT('h1)
	) name8038 (
		_w7118_,
		_w7054_,
		_w8571_
	);
	LUT4 #(
		.INIT('h0d05)
	) name8039 (
		\sa33_reg[2]/P0001 ,
		_w8291_,
		_w8570_,
		_w8571_,
		_w8572_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8040 (
		\sa33_reg[0]/P0001 ,
		_w8569_,
		_w8566_,
		_w8572_,
		_w8573_
	);
	LUT4 #(
		.INIT('h0111)
	) name8041 (
		\sa33_reg[1]/P0001 ,
		_w7088_,
		_w7138_,
		_w7139_,
		_w8574_
	);
	LUT4 #(
		.INIT('hd8ff)
	) name8042 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8575_
	);
	LUT3 #(
		.INIT('h72)
	) name8043 (
		\sa33_reg[4]/P0001 ,
		_w7141_,
		_w8575_,
		_w8576_
	);
	LUT3 #(
		.INIT('h40)
	) name8044 (
		_w8005_,
		_w8574_,
		_w8576_,
		_w8577_
	);
	LUT3 #(
		.INIT('h7e)
	) name8045 (
		\sa33_reg[4]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8578_
	);
	LUT2 #(
		.INIT('h2)
	) name8046 (
		_w7055_,
		_w8578_,
		_w8579_
	);
	LUT2 #(
		.INIT('h8)
	) name8047 (
		_w7062_,
		_w7344_,
		_w8580_
	);
	LUT3 #(
		.INIT('h2a)
	) name8048 (
		\sa33_reg[1]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7063_,
		_w8581_
	);
	LUT3 #(
		.INIT('h10)
	) name8049 (
		_w8580_,
		_w8579_,
		_w8581_,
		_w8582_
	);
	LUT4 #(
		.INIT('h002a)
	) name8050 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[4]/P0001 ,
		_w7141_,
		_w8001_,
		_w8583_
	);
	LUT3 #(
		.INIT('h54)
	) name8051 (
		_w7043_,
		_w7358_,
		_w7914_,
		_w8584_
	);
	LUT4 #(
		.INIT('h0015)
	) name8052 (
		\sa33_reg[2]/P0001 ,
		\sa33_reg[6]/P0001 ,
		_w7134_,
		_w7353_,
		_w8585_
	);
	LUT3 #(
		.INIT('h45)
	) name8053 (
		_w8583_,
		_w8584_,
		_w8585_,
		_w8586_
	);
	LUT4 #(
		.INIT('h5501)
	) name8054 (
		\sa33_reg[0]/P0001 ,
		_w8577_,
		_w8582_,
		_w8586_,
		_w8587_
	);
	LUT3 #(
		.INIT('h02)
	) name8055 (
		\sa33_reg[2]/P0001 ,
		_w7311_,
		_w7965_,
		_w8588_
	);
	LUT4 #(
		.INIT('h0001)
	) name8056 (
		\sa33_reg[2]/P0001 ,
		_w7119_,
		_w7793_,
		_w7772_,
		_w8589_
	);
	LUT2 #(
		.INIT('h1)
	) name8057 (
		_w7962_,
		_w8512_,
		_w8590_
	);
	LUT4 #(
		.INIT('h0155)
	) name8058 (
		\sa33_reg[1]/P0001 ,
		_w8588_,
		_w8589_,
		_w8590_,
		_w8591_
	);
	LUT4 #(
		.INIT('hf7fa)
	) name8059 (
		\sa33_reg[3]/P0001 ,
		\sa33_reg[5]/P0001 ,
		\sa33_reg[6]/P0001 ,
		\sa33_reg[7]/NET0131 ,
		_w8592_
	);
	LUT4 #(
		.INIT('hc0d0)
	) name8060 (
		\sa33_reg[4]/P0001 ,
		_w7948_,
		_w7952_,
		_w8592_,
		_w8593_
	);
	LUT3 #(
		.INIT('h80)
	) name8061 (
		\sa33_reg[1]/P0001 ,
		_w7142_,
		_w7342_,
		_w8594_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name8062 (
		\sa33_reg[5]/P0001 ,
		_w7044_,
		_w7055_,
		_w7066_,
		_w8595_
	);
	LUT4 #(
		.INIT('h0777)
	) name8063 (
		_w7113_,
		_w7119_,
		_w7799_,
		_w8277_,
		_w8596_
	);
	LUT4 #(
		.INIT('h1000)
	) name8064 (
		_w8593_,
		_w8594_,
		_w8595_,
		_w8596_,
		_w8597_
	);
	LUT2 #(
		.INIT('h4)
	) name8065 (
		_w8591_,
		_w8597_,
		_w8598_
	);
	LUT3 #(
		.INIT('h10)
	) name8066 (
		_w8573_,
		_w8587_,
		_w8598_,
		_w8599_
	);
	LUT4 #(
		.INIT('h5655)
	) name8067 (
		\u0_w_reg[0][22]/P0001 ,
		_w8573_,
		_w8587_,
		_w8598_,
		_w8600_
	);
	LUT2 #(
		.INIT('h6)
	) name8068 (
		_w7551_,
		_w8600_,
		_w8601_
	);
	LUT3 #(
		.INIT('h82)
	) name8069 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[118]/P0001 ,
		\u0_w_reg[0][22]/P0001 ,
		_w8602_
	);
	LUT4 #(
		.INIT('h00eb)
	) name8070 (
		\ld_r_reg/P0001 ,
		_w8562_,
		_w8601_,
		_w8602_,
		_w8603_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name8071 (
		\u0_w_reg[0][8]/P0001 ,
		_w7991_,
		_w8004_,
		_w8017_,
		_w8604_
	);
	LUT4 #(
		.INIT('h9669)
	) name8072 (
		_w7655_,
		_w7908_,
		_w7971_,
		_w8123_,
		_w8605_
	);
	LUT3 #(
		.INIT('h82)
	) name8073 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[104]/P0001 ,
		\u0_w_reg[0][8]/P0001 ,
		_w8606_
	);
	LUT4 #(
		.INIT('h00be)
	) name8074 (
		\ld_r_reg/P0001 ,
		_w8604_,
		_w8605_,
		_w8606_,
		_w8607_
	);
	LUT4 #(
		.INIT('h6996)
	) name8075 (
		_w8169_,
		_w8218_,
		_w8396_,
		_w8480_,
		_w8608_
	);
	LUT4 #(
		.INIT('ha955)
	) name8076 (
		\u0_w_reg[0][3]/P0001 ,
		_w8499_,
		_w8511_,
		_w8528_,
		_w8609_
	);
	LUT3 #(
		.INIT('h96)
	) name8077 (
		_w7971_,
		_w8262_,
		_w8609_,
		_w8610_
	);
	LUT3 #(
		.INIT('h82)
	) name8078 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[99]/P0001 ,
		\u0_w_reg[0][3]/P0001 ,
		_w8611_
	);
	LUT4 #(
		.INIT('h00be)
	) name8079 (
		\ld_r_reg/P0001 ,
		_w8608_,
		_w8610_,
		_w8611_,
		_w8612_
	);
	LUT4 #(
		.INIT('ha955)
	) name8080 (
		\u0_w_reg[0][26]/P0001 ,
		_w8499_,
		_w8511_,
		_w8528_,
		_w8613_
	);
	LUT3 #(
		.INIT('h69)
	) name8081 (
		_w8350_,
		_w8437_,
		_w8613_,
		_w8614_
	);
	LUT3 #(
		.INIT('h28)
	) name8082 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[122]/P0001 ,
		\u0_w_reg[0][26]/P0001 ,
		_w8615_
	);
	LUT4 #(
		.INIT('hff14)
	) name8083 (
		\ld_r_reg/P0001 ,
		_w8069_,
		_w8614_,
		_w8615_,
		_w8616_
	);
	LUT4 #(
		.INIT('hb44b)
	) name8084 (
		_w7725_,
		_w7761_,
		_w8350_,
		_w8396_,
		_w8617_
	);
	LUT4 #(
		.INIT('h5655)
	) name8085 (
		\u0_w_reg[0][2]/P0001 ,
		_w8423_,
		_w8413_,
		_w8436_,
		_w8618_
	);
	LUT2 #(
		.INIT('h6)
	) name8086 (
		_w7817_,
		_w8618_,
		_w8619_
	);
	LUT3 #(
		.INIT('h82)
	) name8087 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[98]/P0001 ,
		\u0_w_reg[0][2]/P0001 ,
		_w8620_
	);
	LUT4 #(
		.INIT('h00eb)
	) name8088 (
		\ld_r_reg/P0001 ,
		_w8617_,
		_w8619_,
		_w8620_,
		_w8621_
	);
	LUT4 #(
		.INIT('h5655)
	) name8089 (
		\u0_w_reg[0][30]/P0001 ,
		_w8573_,
		_w8587_,
		_w8598_,
		_w8622_
	);
	LUT3 #(
		.INIT('h69)
	) name8090 (
		_w7491_,
		_w7551_,
		_w8622_,
		_w8623_
	);
	LUT3 #(
		.INIT('h28)
	) name8091 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[126]/P0001 ,
		\u0_w_reg[0][30]/P0001 ,
		_w8624_
	);
	LUT4 #(
		.INIT('hff14)
	) name8092 (
		\ld_r_reg/P0001 ,
		_w7300_,
		_w8623_,
		_w8624_,
		_w8625_
	);
	LUT2 #(
		.INIT('h9)
	) name8093 (
		\u0_w_reg[0][31]/P0001 ,
		_w7706_,
		_w8626_
	);
	LUT4 #(
		.INIT('h6996)
	) name8094 (
		_w7433_,
		_w7491_,
		_w7908_,
		_w7971_,
		_w8627_
	);
	LUT3 #(
		.INIT('h82)
	) name8095 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[127]/P0001 ,
		\u0_w_reg[0][31]/P0001 ,
		_w8628_
	);
	LUT4 #(
		.INIT('h00be)
	) name8096 (
		\ld_r_reg/P0001 ,
		_w8626_,
		_w8627_,
		_w8628_,
		_w8629_
	);
	LUT3 #(
		.INIT('h96)
	) name8097 (
		_w7865_,
		_w8068_,
		_w8396_,
		_w8630_
	);
	LUT4 #(
		.INIT('ha955)
	) name8098 (
		\u0_w_reg[0][18]/P0001 ,
		_w8499_,
		_w8511_,
		_w8528_,
		_w8631_
	);
	LUT2 #(
		.INIT('h6)
	) name8099 (
		_w8437_,
		_w8631_,
		_w8632_
	);
	LUT3 #(
		.INIT('h82)
	) name8100 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[114]/P0001 ,
		\u0_w_reg[0][18]/P0001 ,
		_w8633_
	);
	LUT4 #(
		.INIT('h00be)
	) name8101 (
		\ld_r_reg/P0001 ,
		_w8630_,
		_w8632_,
		_w8633_,
		_w8634_
	);
	LUT3 #(
		.INIT('h69)
	) name8102 (
		_w7491_,
		_w7551_,
		_w8169_,
		_w8635_
	);
	LUT3 #(
		.INIT('h69)
	) name8103 (
		\u0_w_reg[0][23]/P0001 ,
		_w7908_,
		_w7971_,
		_w8636_
	);
	LUT3 #(
		.INIT('h82)
	) name8104 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[119]/P0001 ,
		\u0_w_reg[0][23]/P0001 ,
		_w8637_
	);
	LUT4 #(
		.INIT('h00eb)
	) name8105 (
		\ld_r_reg/P0001 ,
		_w8635_,
		_w8636_,
		_w8637_,
		_w8638_
	);
	LUT3 #(
		.INIT('h69)
	) name8106 (
		_w7031_,
		_w7433_,
		_w7491_,
		_w8639_
	);
	LUT4 #(
		.INIT('h5655)
	) name8107 (
		\u0_w_reg[0][14]/P0001 ,
		_w8573_,
		_w8587_,
		_w8598_,
		_w8640_
	);
	LUT3 #(
		.INIT('hb4)
	) name8108 (
		_w7074_,
		_w7146_,
		_w8640_,
		_w8641_
	);
	LUT3 #(
		.INIT('h82)
	) name8109 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[110]/P0001 ,
		\u0_w_reg[0][14]/P0001 ,
		_w8642_
	);
	LUT4 #(
		.INIT('h00eb)
	) name8110 (
		\ld_r_reg/P0001 ,
		_w8639_,
		_w8641_,
		_w8642_,
		_w8643_
	);
	LUT3 #(
		.INIT('h69)
	) name8111 (
		_w7551_,
		_w7706_,
		_w8169_,
		_w8644_
	);
	LUT4 #(
		.INIT('h5655)
	) name8112 (
		\u0_w_reg[0][15]/P0001 ,
		_w7951_,
		_w7934_,
		_w7970_,
		_w8645_
	);
	LUT2 #(
		.INIT('h6)
	) name8113 (
		_w8599_,
		_w8645_,
		_w8646_
	);
	LUT3 #(
		.INIT('h82)
	) name8114 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[111]/P0001 ,
		\u0_w_reg[0][15]/P0001 ,
		_w8647_
	);
	LUT4 #(
		.INIT('h00eb)
	) name8115 (
		\ld_r_reg/P0001 ,
		_w8644_,
		_w8646_,
		_w8647_,
		_w8648_
	);
	LUT3 #(
		.INIT('h69)
	) name8116 (
		_w7433_,
		_w7706_,
		_w8169_,
		_w8649_
	);
	LUT4 #(
		.INIT('h5655)
	) name8117 (
		\u0_w_reg[0][7]/P0001 ,
		_w8573_,
		_w8587_,
		_w8598_,
		_w8650_
	);
	LUT2 #(
		.INIT('h6)
	) name8118 (
		_w7908_,
		_w8650_,
		_w8651_
	);
	LUT3 #(
		.INIT('h82)
	) name8119 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[103]/P0001 ,
		\u0_w_reg[0][7]/P0001 ,
		_w8652_
	);
	LUT4 #(
		.INIT('h00eb)
	) name8120 (
		\ld_r_reg/P0001 ,
		_w8649_,
		_w8651_,
		_w8652_,
		_w8653_
	);
	LUT2 #(
		.INIT('h4)
	) name8121 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w8654_
	);
	LUT4 #(
		.INIT('h0040)
	) name8122 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8655_
	);
	LUT2 #(
		.INIT('h2)
	) name8123 (
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8656_
	);
	LUT2 #(
		.INIT('h1)
	) name8124 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w8657_
	);
	LUT4 #(
		.INIT('h0010)
	) name8125 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8658_
	);
	LUT2 #(
		.INIT('h4)
	) name8126 (
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8659_
	);
	LUT4 #(
		.INIT('hf5ef)
	) name8127 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8660_
	);
	LUT3 #(
		.INIT('h45)
	) name8128 (
		\u0_w_reg[3][18]/P0001 ,
		_w8655_,
		_w8660_,
		_w8661_
	);
	LUT2 #(
		.INIT('h8)
	) name8129 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8662_
	);
	LUT4 #(
		.INIT('h1000)
	) name8130 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8663_
	);
	LUT2 #(
		.INIT('h2)
	) name8131 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8664_
	);
	LUT2 #(
		.INIT('h1)
	) name8132 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8665_
	);
	LUT4 #(
		.INIT('h0002)
	) name8133 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8666_
	);
	LUT3 #(
		.INIT('h0b)
	) name8134 (
		\u0_w_reg[3][23]/P0001 ,
		_w8663_,
		_w8666_,
		_w8667_
	);
	LUT3 #(
		.INIT('h40)
	) name8135 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8668_
	);
	LUT4 #(
		.INIT('h0400)
	) name8136 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8669_
	);
	LUT2 #(
		.INIT('h2)
	) name8137 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8670_
	);
	LUT4 #(
		.INIT('h0080)
	) name8138 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8671_
	);
	LUT3 #(
		.INIT('h13)
	) name8139 (
		\u0_w_reg[3][18]/P0001 ,
		_w8669_,
		_w8671_,
		_w8672_
	);
	LUT3 #(
		.INIT('h80)
	) name8140 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8673_
	);
	LUT2 #(
		.INIT('h1)
	) name8141 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w8674_
	);
	LUT2 #(
		.INIT('h8)
	) name8142 (
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8675_
	);
	LUT3 #(
		.INIT('h40)
	) name8143 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8676_
	);
	LUT4 #(
		.INIT('h1000)
	) name8144 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8677_
	);
	LUT3 #(
		.INIT('h0d)
	) name8145 (
		_w8673_,
		_w8674_,
		_w8677_,
		_w8678_
	);
	LUT4 #(
		.INIT('h4000)
	) name8146 (
		_w8661_,
		_w8667_,
		_w8672_,
		_w8678_,
		_w8679_
	);
	LUT2 #(
		.INIT('h1)
	) name8147 (
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8680_
	);
	LUT3 #(
		.INIT('h01)
	) name8148 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8681_
	);
	LUT4 #(
		.INIT('h0002)
	) name8149 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8682_
	);
	LUT2 #(
		.INIT('h4)
	) name8150 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8683_
	);
	LUT3 #(
		.INIT('h20)
	) name8151 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8684_
	);
	LUT4 #(
		.INIT('h0200)
	) name8152 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8685_
	);
	LUT3 #(
		.INIT('h54)
	) name8153 (
		\u0_w_reg[3][19]/P0001 ,
		_w8682_,
		_w8685_,
		_w8686_
	);
	LUT3 #(
		.INIT('h80)
	) name8154 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8687_
	);
	LUT3 #(
		.INIT('h01)
	) name8155 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8688_
	);
	LUT2 #(
		.INIT('h8)
	) name8156 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w8689_
	);
	LUT4 #(
		.INIT('h135f)
	) name8157 (
		_w8657_,
		_w8688_,
		_w8687_,
		_w8689_,
		_w8690_
	);
	LUT2 #(
		.INIT('h4)
	) name8158 (
		_w8686_,
		_w8690_,
		_w8691_
	);
	LUT2 #(
		.INIT('h1)
	) name8159 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8692_
	);
	LUT3 #(
		.INIT('h01)
	) name8160 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8693_
	);
	LUT3 #(
		.INIT('h80)
	) name8161 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8694_
	);
	LUT3 #(
		.INIT('h7e)
	) name8162 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8695_
	);
	LUT4 #(
		.INIT('h8002)
	) name8163 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8696_
	);
	LUT2 #(
		.INIT('h4)
	) name8164 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8697_
	);
	LUT4 #(
		.INIT('h0020)
	) name8165 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8698_
	);
	LUT3 #(
		.INIT('h01)
	) name8166 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8699_
	);
	LUT4 #(
		.INIT('h0023)
	) name8167 (
		\u0_w_reg[3][19]/P0001 ,
		_w8696_,
		_w8698_,
		_w8699_,
		_w8700_
	);
	LUT3 #(
		.INIT('h02)
	) name8168 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8701_
	);
	LUT4 #(
		.INIT('h0008)
	) name8169 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8702_
	);
	LUT2 #(
		.INIT('h4)
	) name8170 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8703_
	);
	LUT4 #(
		.INIT('h1000)
	) name8171 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8704_
	);
	LUT2 #(
		.INIT('h1)
	) name8172 (
		_w8702_,
		_w8704_,
		_w8705_
	);
	LUT3 #(
		.INIT('h54)
	) name8173 (
		\u0_w_reg[3][18]/P0001 ,
		_w8702_,
		_w8704_,
		_w8706_
	);
	LUT2 #(
		.INIT('h8)
	) name8174 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8707_
	);
	LUT4 #(
		.INIT('h0800)
	) name8175 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8708_
	);
	LUT4 #(
		.INIT('h0001)
	) name8176 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8709_
	);
	LUT3 #(
		.INIT('h0b)
	) name8177 (
		\u0_w_reg[3][18]/P0001 ,
		_w8708_,
		_w8709_,
		_w8710_
	);
	LUT4 #(
		.INIT('hd800)
	) name8178 (
		\u0_w_reg[3][18]/P0001 ,
		_w8700_,
		_w8705_,
		_w8710_,
		_w8711_
	);
	LUT4 #(
		.INIT('hd800)
	) name8179 (
		\u0_w_reg[3][17]/P0001 ,
		_w8679_,
		_w8691_,
		_w8711_,
		_w8712_
	);
	LUT2 #(
		.INIT('h1)
	) name8180 (
		\u0_w_reg[3][16]/P0001 ,
		_w8712_,
		_w8713_
	);
	LUT2 #(
		.INIT('h2)
	) name8181 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w8714_
	);
	LUT3 #(
		.INIT('h20)
	) name8182 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		_w8715_
	);
	LUT4 #(
		.INIT('hdfdc)
	) name8183 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8716_
	);
	LUT3 #(
		.INIT('h45)
	) name8184 (
		\u0_w_reg[3][18]/P0001 ,
		_w8701_,
		_w8716_,
		_w8717_
	);
	LUT4 #(
		.INIT('h0200)
	) name8185 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8718_
	);
	LUT3 #(
		.INIT('h13)
	) name8186 (
		_w8654_,
		_w8718_,
		_w8681_,
		_w8719_
	);
	LUT3 #(
		.INIT('h04)
	) name8187 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8720_
	);
	LUT2 #(
		.INIT('h2)
	) name8188 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8721_
	);
	LUT2 #(
		.INIT('h8)
	) name8189 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w8722_
	);
	LUT3 #(
		.INIT('h08)
	) name8190 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8723_
	);
	LUT4 #(
		.INIT('h153f)
	) name8191 (
		_w8721_,
		_w8707_,
		_w8720_,
		_w8723_,
		_w8724_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name8192 (
		\u0_w_reg[3][17]/P0001 ,
		_w8717_,
		_w8719_,
		_w8724_,
		_w8725_
	);
	LUT3 #(
		.INIT('h10)
	) name8193 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8726_
	);
	LUT4 #(
		.INIT('h0008)
	) name8194 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8727_
	);
	LUT3 #(
		.INIT('ha8)
	) name8195 (
		\u0_w_reg[3][18]/P0001 ,
		_w8726_,
		_w8727_,
		_w8728_
	);
	LUT2 #(
		.INIT('h4)
	) name8196 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w8729_
	);
	LUT3 #(
		.INIT('h10)
	) name8197 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8730_
	);
	LUT2 #(
		.INIT('h8)
	) name8198 (
		_w8729_,
		_w8730_,
		_w8731_
	);
	LUT2 #(
		.INIT('h2)
	) name8199 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w8732_
	);
	LUT3 #(
		.INIT('h08)
	) name8200 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8733_
	);
	LUT4 #(
		.INIT('h4000)
	) name8201 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8734_
	);
	LUT4 #(
		.INIT('h45cf)
	) name8202 (
		\u0_w_reg[3][22]/P0001 ,
		_w8732_,
		_w8733_,
		_w8734_,
		_w8735_
	);
	LUT4 #(
		.INIT('h5455)
	) name8203 (
		\u0_w_reg[3][17]/P0001 ,
		_w8728_,
		_w8731_,
		_w8735_,
		_w8736_
	);
	LUT4 #(
		.INIT('h0080)
	) name8204 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8737_
	);
	LUT4 #(
		.INIT('h0020)
	) name8205 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8738_
	);
	LUT3 #(
		.INIT('h04)
	) name8206 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8739_
	);
	LUT4 #(
		.INIT('h2000)
	) name8207 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8740_
	);
	LUT4 #(
		.INIT('hdfbb)
	) name8208 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8741_
	);
	LUT4 #(
		.INIT('h5455)
	) name8209 (
		\u0_w_reg[3][18]/P0001 ,
		_w8737_,
		_w8738_,
		_w8741_,
		_w8742_
	);
	LUT3 #(
		.INIT('h02)
	) name8210 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w8743_
	);
	LUT4 #(
		.INIT('h0002)
	) name8211 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		_w8744_
	);
	LUT4 #(
		.INIT('hf3fd)
	) name8212 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		_w8745_
	);
	LUT3 #(
		.INIT('h80)
	) name8213 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8746_
	);
	LUT4 #(
		.INIT('h8000)
	) name8214 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8747_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name8215 (
		_w8656_,
		_w8745_,
		_w8732_,
		_w8747_,
		_w8748_
	);
	LUT2 #(
		.INIT('h4)
	) name8216 (
		_w8742_,
		_w8748_,
		_w8749_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8217 (
		\u0_w_reg[3][16]/P0001 ,
		_w8736_,
		_w8725_,
		_w8749_,
		_w8750_
	);
	LUT4 #(
		.INIT('h0001)
	) name8218 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8751_
	);
	LUT3 #(
		.INIT('h04)
	) name8219 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8752_
	);
	LUT3 #(
		.INIT('heb)
	) name8220 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8753_
	);
	LUT2 #(
		.INIT('h2)
	) name8221 (
		_w8654_,
		_w8753_,
		_w8754_
	);
	LUT4 #(
		.INIT('h0080)
	) name8222 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8755_
	);
	LUT3 #(
		.INIT('h07)
	) name8223 (
		\u0_w_reg[3][22]/P0001 ,
		_w8734_,
		_w8755_,
		_w8756_
	);
	LUT4 #(
		.INIT('h1311)
	) name8224 (
		\u0_w_reg[3][18]/P0001 ,
		_w8751_,
		_w8754_,
		_w8756_,
		_w8757_
	);
	LUT2 #(
		.INIT('h1)
	) name8225 (
		\u0_w_reg[3][17]/P0001 ,
		_w8757_,
		_w8758_
	);
	LUT2 #(
		.INIT('h8)
	) name8226 (
		_w8732_,
		_w8671_,
		_w8759_
	);
	LUT3 #(
		.INIT('h02)
	) name8227 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		_w8760_
	);
	LUT4 #(
		.INIT('h23af)
	) name8228 (
		\u0_w_reg[3][18]/P0001 ,
		_w8680_,
		_w8708_,
		_w8760_,
		_w8761_
	);
	LUT3 #(
		.INIT('h8a)
	) name8229 (
		\u0_w_reg[3][17]/P0001 ,
		_w8759_,
		_w8761_,
		_w8762_
	);
	LUT3 #(
		.INIT('h40)
	) name8230 (
		\u0_w_reg[3][18]/P0001 ,
		_w8746_,
		_w8664_,
		_w8763_
	);
	LUT2 #(
		.INIT('h1)
	) name8231 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w8764_
	);
	LUT4 #(
		.INIT('haeaf)
	) name8232 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w8740_,
		_w8668_,
		_w8765_
	);
	LUT3 #(
		.INIT('h45)
	) name8233 (
		\u0_w_reg[3][17]/P0001 ,
		_w8763_,
		_w8765_,
		_w8766_
	);
	LUT4 #(
		.INIT('h0020)
	) name8234 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8767_
	);
	LUT2 #(
		.INIT('h4)
	) name8235 (
		\u0_w_reg[3][23]/P0001 ,
		_w8767_,
		_w8768_
	);
	LUT3 #(
		.INIT('h10)
	) name8236 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8767_,
		_w8769_
	);
	LUT4 #(
		.INIT('h0008)
	) name8237 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8770_
	);
	LUT2 #(
		.INIT('h8)
	) name8238 (
		_w8689_,
		_w8770_,
		_w8771_
	);
	LUT3 #(
		.INIT('h01)
	) name8239 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		_w8772_
	);
	LUT4 #(
		.INIT('h153f)
	) name8240 (
		_w8675_,
		_w8689_,
		_w8770_,
		_w8772_,
		_w8773_
	);
	LUT2 #(
		.INIT('h4)
	) name8241 (
		_w8769_,
		_w8773_,
		_w8774_
	);
	LUT3 #(
		.INIT('h10)
	) name8242 (
		_w8766_,
		_w8762_,
		_w8774_,
		_w8775_
	);
	LUT3 #(
		.INIT('h10)
	) name8243 (
		_w8750_,
		_w8758_,
		_w8775_,
		_w8776_
	);
	LUT3 #(
		.INIT('h65)
	) name8244 (
		\u0_r0_out_reg[29]/P0001 ,
		_w8713_,
		_w8776_,
		_w8777_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name8245 (
		\key[125]_pad ,
		ld_pad,
		\u0_w_reg[0][29]/P0001 ,
		_w8777_,
		_w8778_
	);
	LUT2 #(
		.INIT('h9)
	) name8246 (
		\u0_w_reg[0][29]/P0001 ,
		\u0_w_reg[1][29]/P0002 ,
		_w8779_
	);
	LUT3 #(
		.INIT('h69)
	) name8247 (
		\u0_w_reg[0][29]/P0001 ,
		\u0_w_reg[1][29]/P0002 ,
		\u0_w_reg[2][29]/P0001 ,
		_w8780_
	);
	LUT4 #(
		.INIT('h9a65)
	) name8248 (
		\u0_r0_out_reg[29]/P0001 ,
		_w8713_,
		_w8776_,
		_w8780_,
		_w8781_
	);
	LUT3 #(
		.INIT('h8b)
	) name8249 (
		\key[61]_pad ,
		ld_pad,
		_w8781_,
		_w8782_
	);
	LUT4 #(
		.INIT('hb88b)
	) name8250 (
		\key[29]_pad ,
		ld_pad,
		\u0_w_reg[3][29]/P0001 ,
		_w8781_,
		_w8783_
	);
	LUT3 #(
		.INIT('h08)
	) name8251 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8784_
	);
	LUT2 #(
		.INIT('h4)
	) name8252 (
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8785_
	);
	LUT3 #(
		.INIT('h20)
	) name8253 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8786_
	);
	LUT4 #(
		.INIT('h0200)
	) name8254 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8787_
	);
	LUT4 #(
		.INIT('hfd3f)
	) name8255 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8788_
	);
	LUT2 #(
		.INIT('h1)
	) name8256 (
		\u0_w_reg[3][10]/P0001 ,
		_w8788_,
		_w8789_
	);
	LUT2 #(
		.INIT('h8)
	) name8257 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		_w8790_
	);
	LUT2 #(
		.INIT('h1)
	) name8258 (
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8791_
	);
	LUT4 #(
		.INIT('h0008)
	) name8259 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8792_
	);
	LUT2 #(
		.INIT('h4)
	) name8260 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8793_
	);
	LUT3 #(
		.INIT('h10)
	) name8261 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8794_
	);
	LUT3 #(
		.INIT('ha8)
	) name8262 (
		\u0_w_reg[3][10]/P0001 ,
		_w8792_,
		_w8794_,
		_w8795_
	);
	LUT2 #(
		.INIT('h8)
	) name8263 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8796_
	);
	LUT3 #(
		.INIT('h80)
	) name8264 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8797_
	);
	LUT4 #(
		.INIT('h8000)
	) name8265 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8798_
	);
	LUT2 #(
		.INIT('h8)
	) name8266 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8799_
	);
	LUT4 #(
		.INIT('h0080)
	) name8267 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8800_
	);
	LUT4 #(
		.INIT('h0023)
	) name8268 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w8798_,
		_w8800_,
		_w8801_
	);
	LUT3 #(
		.INIT('h10)
	) name8269 (
		_w8795_,
		_w8789_,
		_w8801_,
		_w8802_
	);
	LUT2 #(
		.INIT('h1)
	) name8270 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8803_
	);
	LUT2 #(
		.INIT('h2)
	) name8271 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8804_
	);
	LUT4 #(
		.INIT('h0002)
	) name8272 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8805_
	);
	LUT3 #(
		.INIT('h8c)
	) name8273 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w8805_,
		_w8806_
	);
	LUT4 #(
		.INIT('h0200)
	) name8274 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8807_
	);
	LUT2 #(
		.INIT('h4)
	) name8275 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		_w8808_
	);
	LUT4 #(
		.INIT('h0400)
	) name8276 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8809_
	);
	LUT2 #(
		.INIT('h2)
	) name8277 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8810_
	);
	LUT3 #(
		.INIT('h08)
	) name8278 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8811_
	);
	LUT4 #(
		.INIT('h5d5f)
	) name8279 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8809_,
		_w8811_,
		_w8812_
	);
	LUT3 #(
		.INIT('h20)
	) name8280 (
		_w8806_,
		_w8807_,
		_w8812_,
		_w8813_
	);
	LUT3 #(
		.INIT('h8a)
	) name8281 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w8798_,
		_w8814_
	);
	LUT2 #(
		.INIT('h1)
	) name8282 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		_w8815_
	);
	LUT4 #(
		.INIT('h0100)
	) name8283 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8816_
	);
	LUT2 #(
		.INIT('h4)
	) name8284 (
		\u0_w_reg[3][15]/P0001 ,
		_w8816_,
		_w8817_
	);
	LUT4 #(
		.INIT('h0020)
	) name8285 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8818_
	);
	LUT3 #(
		.INIT('h04)
	) name8286 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8819_
	);
	LUT4 #(
		.INIT('h5545)
	) name8287 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8820_
	);
	LUT3 #(
		.INIT('h10)
	) name8288 (
		_w8800_,
		_w8818_,
		_w8820_,
		_w8821_
	);
	LUT3 #(
		.INIT('h0d)
	) name8289 (
		_w8814_,
		_w8817_,
		_w8821_,
		_w8822_
	);
	LUT2 #(
		.INIT('h4)
	) name8290 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w8823_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name8291 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w8824_
	);
	LUT2 #(
		.INIT('h2)
	) name8292 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		_w8825_
	);
	LUT3 #(
		.INIT('h20)
	) name8293 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		_w8826_
	);
	LUT3 #(
		.INIT('h8a)
	) name8294 (
		\u0_w_reg[3][8]/P0001 ,
		_w8824_,
		_w8826_,
		_w8827_
	);
	LUT3 #(
		.INIT('h10)
	) name8295 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8828_
	);
	LUT3 #(
		.INIT('h23)
	) name8296 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8829_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name8297 (
		_w8796_,
		_w8823_,
		_w8828_,
		_w8829_,
		_w8830_
	);
	LUT2 #(
		.INIT('h8)
	) name8298 (
		_w8827_,
		_w8830_,
		_w8831_
	);
	LUT4 #(
		.INIT('h5400)
	) name8299 (
		_w8822_,
		_w8802_,
		_w8813_,
		_w8831_,
		_w8832_
	);
	LUT4 #(
		.INIT('h0010)
	) name8300 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8833_
	);
	LUT4 #(
		.INIT('h0040)
	) name8301 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8834_
	);
	LUT4 #(
		.INIT('h5554)
	) name8302 (
		\u0_w_reg[3][10]/P0001 ,
		_w8786_,
		_w8833_,
		_w8834_,
		_w8835_
	);
	LUT3 #(
		.INIT('h80)
	) name8303 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8836_
	);
	LUT2 #(
		.INIT('h8)
	) name8304 (
		_w8804_,
		_w8836_,
		_w8837_
	);
	LUT3 #(
		.INIT('h40)
	) name8305 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8838_
	);
	LUT4 #(
		.INIT('h1000)
	) name8306 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8839_
	);
	LUT4 #(
		.INIT('h0002)
	) name8307 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8840_
	);
	LUT3 #(
		.INIT('h02)
	) name8308 (
		\u0_w_reg[3][9]/P0001 ,
		_w8839_,
		_w8840_,
		_w8841_
	);
	LUT4 #(
		.INIT('h0040)
	) name8309 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8842_
	);
	LUT2 #(
		.INIT('h4)
	) name8310 (
		\u0_w_reg[3][12]/P0001 ,
		_w8842_,
		_w8843_
	);
	LUT4 #(
		.INIT('h0400)
	) name8311 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8844_
	);
	LUT3 #(
		.INIT('h80)
	) name8312 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8845_
	);
	LUT2 #(
		.INIT('h1)
	) name8313 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		_w8846_
	);
	LUT3 #(
		.INIT('h51)
	) name8314 (
		_w8844_,
		_w8845_,
		_w8846_,
		_w8847_
	);
	LUT4 #(
		.INIT('h1000)
	) name8315 (
		_w8843_,
		_w8837_,
		_w8847_,
		_w8841_,
		_w8848_
	);
	LUT4 #(
		.INIT('h4000)
	) name8316 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8849_
	);
	LUT4 #(
		.INIT('h0200)
	) name8317 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8850_
	);
	LUT2 #(
		.INIT('h2)
	) name8318 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		_w8851_
	);
	LUT4 #(
		.INIT('h0002)
	) name8319 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8852_
	);
	LUT4 #(
		.INIT('h5554)
	) name8320 (
		\u0_w_reg[3][11]/P0001 ,
		_w8850_,
		_w8852_,
		_w8849_,
		_w8853_
	);
	LUT2 #(
		.INIT('h8)
	) name8321 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w8854_
	);
	LUT3 #(
		.INIT('h08)
	) name8322 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		_w8855_
	);
	LUT3 #(
		.INIT('h15)
	) name8323 (
		\u0_w_reg[3][9]/P0001 ,
		_w8803_,
		_w8855_,
		_w8856_
	);
	LUT2 #(
		.INIT('h4)
	) name8324 (
		_w8853_,
		_w8856_,
		_w8857_
	);
	LUT3 #(
		.INIT('h02)
	) name8325 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8858_
	);
	LUT4 #(
		.INIT('h0008)
	) name8326 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8859_
	);
	LUT4 #(
		.INIT('h1000)
	) name8327 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8860_
	);
	LUT4 #(
		.INIT('h0800)
	) name8328 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8861_
	);
	LUT4 #(
		.INIT('h0001)
	) name8329 (
		\u0_w_reg[3][10]/P0001 ,
		_w8859_,
		_w8860_,
		_w8861_,
		_w8862_
	);
	LUT2 #(
		.INIT('h1)
	) name8330 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8863_
	);
	LUT3 #(
		.INIT('h01)
	) name8331 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8864_
	);
	LUT3 #(
		.INIT('h7e)
	) name8332 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8865_
	);
	LUT4 #(
		.INIT('h8002)
	) name8333 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8866_
	);
	LUT4 #(
		.INIT('h0020)
	) name8334 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8867_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8335 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8868_
	);
	LUT4 #(
		.INIT('h2300)
	) name8336 (
		\u0_w_reg[3][11]/P0001 ,
		_w8866_,
		_w8867_,
		_w8868_,
		_w8869_
	);
	LUT4 #(
		.INIT('h0001)
	) name8337 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8870_
	);
	LUT2 #(
		.INIT('h1)
	) name8338 (
		\u0_w_reg[3][8]/P0001 ,
		_w8870_,
		_w8871_
	);
	LUT3 #(
		.INIT('he0)
	) name8339 (
		_w8862_,
		_w8869_,
		_w8871_,
		_w8872_
	);
	LUT4 #(
		.INIT('hf400)
	) name8340 (
		_w8835_,
		_w8848_,
		_w8857_,
		_w8872_,
		_w8873_
	);
	LUT4 #(
		.INIT('h0080)
	) name8341 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8874_
	);
	LUT3 #(
		.INIT('h04)
	) name8342 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8875_
	);
	LUT3 #(
		.INIT('h6b)
	) name8343 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8876_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name8344 (
		\u0_w_reg[3][10]/P0001 ,
		_w8808_,
		_w8874_,
		_w8876_,
		_w8877_
	);
	LUT2 #(
		.INIT('h4)
	) name8345 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w8878_
	);
	LUT3 #(
		.INIT('h08)
	) name8346 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8879_
	);
	LUT4 #(
		.INIT('h0080)
	) name8347 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8880_
	);
	LUT2 #(
		.INIT('h8)
	) name8348 (
		_w8878_,
		_w8880_,
		_w8881_
	);
	LUT3 #(
		.INIT('h40)
	) name8349 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8882_
	);
	LUT2 #(
		.INIT('h1)
	) name8350 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w8883_
	);
	LUT2 #(
		.INIT('h8)
	) name8351 (
		_w8882_,
		_w8883_,
		_w8884_
	);
	LUT4 #(
		.INIT('h0001)
	) name8352 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8885_
	);
	LUT3 #(
		.INIT('h07)
	) name8353 (
		_w8796_,
		_w8828_,
		_w8885_,
		_w8886_
	);
	LUT4 #(
		.INIT('h0100)
	) name8354 (
		_w8877_,
		_w8884_,
		_w8881_,
		_w8886_,
		_w8887_
	);
	LUT3 #(
		.INIT('h40)
	) name8355 (
		\u0_w_reg[3][11]/P0001 ,
		_w8804_,
		_w8836_,
		_w8888_
	);
	LUT4 #(
		.INIT('h0002)
	) name8356 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8889_
	);
	LUT4 #(
		.INIT('h8caf)
	) name8357 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		_w8861_,
		_w8889_,
		_w8890_
	);
	LUT2 #(
		.INIT('h4)
	) name8358 (
		_w8888_,
		_w8890_,
		_w8891_
	);
	LUT2 #(
		.INIT('h4)
	) name8359 (
		\u0_w_reg[3][10]/P0001 ,
		_w8839_,
		_w8892_
	);
	LUT4 #(
		.INIT('h0080)
	) name8360 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8893_
	);
	LUT2 #(
		.INIT('h2)
	) name8361 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8894_
	);
	LUT2 #(
		.INIT('h8)
	) name8362 (
		_w8893_,
		_w8894_,
		_w8895_
	);
	LUT3 #(
		.INIT('h02)
	) name8363 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8896_
	);
	LUT3 #(
		.INIT('h40)
	) name8364 (
		\u0_w_reg[3][10]/P0001 ,
		_w8810_,
		_w8896_,
		_w8897_
	);
	LUT3 #(
		.INIT('h01)
	) name8365 (
		_w8895_,
		_w8897_,
		_w8892_,
		_w8898_
	);
	LUT4 #(
		.INIT('he400)
	) name8366 (
		\u0_w_reg[3][9]/P0001 ,
		_w8887_,
		_w8891_,
		_w8898_,
		_w8899_
	);
	LUT4 #(
		.INIT('ha955)
	) name8367 (
		\u0_w_reg[0][21]/P0001 ,
		_w8832_,
		_w8873_,
		_w8899_,
		_w8900_
	);
	LUT2 #(
		.INIT('h9)
	) name8368 (
		\u0_w_reg[1][21]/P0001 ,
		\u0_w_reg[2][21]/P0001 ,
		_w8901_
	);
	LUT4 #(
		.INIT('hb88b)
	) name8369 (
		\key[53]_pad ,
		ld_pad,
		_w8900_,
		_w8901_,
		_w8902_
	);
	LUT2 #(
		.INIT('h4)
	) name8370 (
		\key[51]_pad ,
		ld_pad,
		_w8903_
	);
	LUT3 #(
		.INIT('h8a)
	) name8371 (
		\u0_w_reg[3][10]/P0001 ,
		_w8819_,
		_w8788_,
		_w8904_
	);
	LUT3 #(
		.INIT('h10)
	) name8372 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		_w8905_
	);
	LUT4 #(
		.INIT('h1000)
	) name8373 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8906_
	);
	LUT2 #(
		.INIT('h1)
	) name8374 (
		_w8885_,
		_w8906_,
		_w8907_
	);
	LUT4 #(
		.INIT('h3b3f)
	) name8375 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w8850_,
		_w8875_,
		_w8908_
	);
	LUT4 #(
		.INIT('h1000)
	) name8376 (
		_w8892_,
		_w8904_,
		_w8907_,
		_w8908_,
		_w8909_
	);
	LUT3 #(
		.INIT('h01)
	) name8377 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8910_
	);
	LUT3 #(
		.INIT('h04)
	) name8378 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8911_
	);
	LUT4 #(
		.INIT('h5545)
	) name8379 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8912_
	);
	LUT4 #(
		.INIT('h0c04)
	) name8380 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8913_
	);
	LUT3 #(
		.INIT('h20)
	) name8381 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8914_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name8382 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8915_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name8383 (
		_w8910_,
		_w8912_,
		_w8913_,
		_w8915_,
		_w8916_
	);
	LUT2 #(
		.INIT('h8)
	) name8384 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8917_
	);
	LUT4 #(
		.INIT('h2000)
	) name8385 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8918_
	);
	LUT4 #(
		.INIT('h4000)
	) name8386 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8919_
	);
	LUT3 #(
		.INIT('h01)
	) name8387 (
		_w8861_,
		_w8918_,
		_w8919_,
		_w8920_
	);
	LUT2 #(
		.INIT('h4)
	) name8388 (
		_w8916_,
		_w8920_,
		_w8921_
	);
	LUT4 #(
		.INIT('h0800)
	) name8389 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8922_
	);
	LUT4 #(
		.INIT('hfddf)
	) name8390 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8923_
	);
	LUT3 #(
		.INIT('h8a)
	) name8391 (
		\u0_w_reg[3][10]/P0001 ,
		_w8922_,
		_w8923_,
		_w8924_
	);
	LUT3 #(
		.INIT('h10)
	) name8392 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8925_
	);
	LUT4 #(
		.INIT('h0100)
	) name8393 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8926_
	);
	LUT4 #(
		.INIT('h8000)
	) name8394 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8927_
	);
	LUT3 #(
		.INIT('h54)
	) name8395 (
		\u0_w_reg[3][10]/P0001 ,
		_w8926_,
		_w8927_,
		_w8928_
	);
	LUT4 #(
		.INIT('h2000)
	) name8396 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8929_
	);
	LUT2 #(
		.INIT('h4)
	) name8397 (
		\u0_w_reg[3][15]/P0001 ,
		_w8929_,
		_w8930_
	);
	LUT3 #(
		.INIT('h10)
	) name8398 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w8861_,
		_w8931_
	);
	LUT4 #(
		.INIT('h0001)
	) name8399 (
		_w8928_,
		_w8930_,
		_w8931_,
		_w8924_,
		_w8932_
	);
	LUT4 #(
		.INIT('he400)
	) name8400 (
		\u0_w_reg[3][9]/P0001 ,
		_w8909_,
		_w8921_,
		_w8932_,
		_w8933_
	);
	LUT3 #(
		.INIT('h40)
	) name8401 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w8861_,
		_w8934_
	);
	LUT3 #(
		.INIT('hf4)
	) name8402 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8935_
	);
	LUT3 #(
		.INIT('h51)
	) name8403 (
		\u0_w_reg[3][9]/P0001 ,
		_w8804_,
		_w8935_,
		_w8936_
	);
	LUT2 #(
		.INIT('h2)
	) name8404 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w8937_
	);
	LUT3 #(
		.INIT('he0)
	) name8405 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8938_
	);
	LUT3 #(
		.INIT('h07)
	) name8406 (
		_w8937_,
		_w8938_,
		_w8926_,
		_w8939_
	);
	LUT3 #(
		.INIT('h40)
	) name8407 (
		_w8934_,
		_w8936_,
		_w8939_,
		_w8940_
	);
	LUT4 #(
		.INIT('h4000)
	) name8408 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w8941_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name8409 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8864_,
		_w8941_,
		_w8942_
	);
	LUT3 #(
		.INIT('h80)
	) name8410 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8943_
	);
	LUT3 #(
		.INIT('h6f)
	) name8411 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8944_
	);
	LUT2 #(
		.INIT('h2)
	) name8412 (
		_w8799_,
		_w8944_,
		_w8945_
	);
	LUT4 #(
		.INIT('h080c)
	) name8413 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w8787_,
		_w8844_,
		_w8946_
	);
	LUT3 #(
		.INIT('h10)
	) name8414 (
		_w8942_,
		_w8945_,
		_w8946_,
		_w8947_
	);
	LUT4 #(
		.INIT('h0080)
	) name8415 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8948_
	);
	LUT4 #(
		.INIT('h5510)
	) name8416 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w8798_,
		_w8948_,
		_w8949_
	);
	LUT4 #(
		.INIT('h0002)
	) name8417 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8950_
	);
	LUT3 #(
		.INIT('ha8)
	) name8418 (
		\u0_w_reg[3][10]/P0001 ,
		_w8849_,
		_w8950_,
		_w8951_
	);
	LUT3 #(
		.INIT('h01)
	) name8419 (
		_w8817_,
		_w8951_,
		_w8949_,
		_w8952_
	);
	LUT3 #(
		.INIT('he0)
	) name8420 (
		_w8940_,
		_w8947_,
		_w8952_,
		_w8953_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8421 (
		\u0_w_reg[3][10]/P0001 ,
		_w8861_,
		_w8918_,
		_w8929_,
		_w8954_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name8422 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8955_
	);
	LUT4 #(
		.INIT('h0100)
	) name8423 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8956_
	);
	LUT2 #(
		.INIT('h8)
	) name8424 (
		_w8878_,
		_w8956_,
		_w8957_
	);
	LUT4 #(
		.INIT('hbafe)
	) name8425 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w8955_,
		_w8956_,
		_w8958_
	);
	LUT3 #(
		.INIT('h8a)
	) name8426 (
		\u0_w_reg[3][9]/P0001 ,
		_w8954_,
		_w8958_,
		_w8959_
	);
	LUT4 #(
		.INIT('h2000)
	) name8427 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8960_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name8428 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		_w8850_,
		_w8960_,
		_w8961_
	);
	LUT2 #(
		.INIT('h2)
	) name8429 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w8962_
	);
	LUT3 #(
		.INIT('h02)
	) name8430 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w8963_
	);
	LUT4 #(
		.INIT('h0010)
	) name8431 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8964_
	);
	LUT4 #(
		.INIT('hffed)
	) name8432 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8965_
	);
	LUT2 #(
		.INIT('h2)
	) name8433 (
		_w8963_,
		_w8965_,
		_w8966_
	);
	LUT4 #(
		.INIT('h0010)
	) name8434 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w8967_
	);
	LUT3 #(
		.INIT('hc8)
	) name8435 (
		_w8858_,
		_w8917_,
		_w8967_,
		_w8968_
	);
	LUT4 #(
		.INIT('h000d)
	) name8436 (
		\u0_w_reg[3][10]/P0001 ,
		_w8961_,
		_w8966_,
		_w8968_,
		_w8969_
	);
	LUT2 #(
		.INIT('h4)
	) name8437 (
		_w8959_,
		_w8969_,
		_w8970_
	);
	LUT4 #(
		.INIT('he400)
	) name8438 (
		\u0_w_reg[3][8]/P0001 ,
		_w8953_,
		_w8933_,
		_w8970_,
		_w8971_
	);
	LUT2 #(
		.INIT('h9)
	) name8439 (
		\u0_w_reg[1][19]/P0001 ,
		\u0_w_reg[2][19]/P0001 ,
		_w8972_
	);
	LUT3 #(
		.INIT('h69)
	) name8440 (
		\u0_w_reg[0][19]/P0001 ,
		_w8971_,
		_w8972_,
		_w8973_
	);
	LUT4 #(
		.INIT('h1441)
	) name8441 (
		ld_pad,
		\u0_w_reg[0][19]/P0001 ,
		_w8971_,
		_w8972_,
		_w8974_
	);
	LUT2 #(
		.INIT('h1)
	) name8442 (
		_w8903_,
		_w8974_,
		_w8975_
	);
	LUT2 #(
		.INIT('h4)
	) name8443 (
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w8976_
	);
	LUT2 #(
		.INIT('h4)
	) name8444 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w8977_
	);
	LUT4 #(
		.INIT('h0400)
	) name8445 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w8978_
	);
	LUT2 #(
		.INIT('h1)
	) name8446 (
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w8979_
	);
	LUT3 #(
		.INIT('h01)
	) name8447 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w8980_
	);
	LUT4 #(
		.INIT('h0002)
	) name8448 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w8981_
	);
	LUT3 #(
		.INIT('h54)
	) name8449 (
		\u0_w_reg[3][29]/P0001 ,
		_w8978_,
		_w8981_,
		_w8982_
	);
	LUT2 #(
		.INIT('h8)
	) name8450 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w8983_
	);
	LUT3 #(
		.INIT('h80)
	) name8451 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w8984_
	);
	LUT4 #(
		.INIT('h4000)
	) name8452 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w8985_
	);
	LUT2 #(
		.INIT('h4)
	) name8453 (
		\u0_w_reg[3][28]/P0001 ,
		_w8985_,
		_w8986_
	);
	LUT2 #(
		.INIT('h1)
	) name8454 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w8987_
	);
	LUT3 #(
		.INIT('h01)
	) name8455 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w8988_
	);
	LUT2 #(
		.INIT('h8)
	) name8456 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w8989_
	);
	LUT3 #(
		.INIT('h15)
	) name8457 (
		\u0_w_reg[3][25]/P0001 ,
		_w8988_,
		_w8989_,
		_w8990_
	);
	LUT3 #(
		.INIT('h10)
	) name8458 (
		_w8982_,
		_w8986_,
		_w8990_,
		_w8991_
	);
	LUT4 #(
		.INIT('h0040)
	) name8459 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w8992_
	);
	LUT2 #(
		.INIT('h2)
	) name8460 (
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w8993_
	);
	LUT4 #(
		.INIT('h0a10)
	) name8461 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w8994_
	);
	LUT3 #(
		.INIT('h54)
	) name8462 (
		\u0_w_reg[3][26]/P0001 ,
		_w8992_,
		_w8994_,
		_w8995_
	);
	LUT2 #(
		.INIT('h8)
	) name8463 (
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w8996_
	);
	LUT3 #(
		.INIT('h40)
	) name8464 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w8997_
	);
	LUT4 #(
		.INIT('h1000)
	) name8465 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w8998_
	);
	LUT2 #(
		.INIT('h2)
	) name8466 (
		\u0_w_reg[3][25]/P0001 ,
		_w8998_,
		_w8999_
	);
	LUT2 #(
		.INIT('h4)
	) name8467 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		_w9000_
	);
	LUT3 #(
		.INIT('h04)
	) name8468 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9001_
	);
	LUT2 #(
		.INIT('h2)
	) name8469 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9002_
	);
	LUT4 #(
		.INIT('h0002)
	) name8470 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9003_
	);
	LUT4 #(
		.INIT('h0400)
	) name8471 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9004_
	);
	LUT4 #(
		.INIT('h0057)
	) name8472 (
		_w9000_,
		_w8976_,
		_w9001_,
		_w9003_,
		_w9005_
	);
	LUT2 #(
		.INIT('h2)
	) name8473 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9006_
	);
	LUT3 #(
		.INIT('h80)
	) name8474 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9007_
	);
	LUT3 #(
		.INIT('h80)
	) name8475 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9008_
	);
	LUT2 #(
		.INIT('h1)
	) name8476 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w9009_
	);
	LUT4 #(
		.INIT('h7707)
	) name8477 (
		_w9006_,
		_w9007_,
		_w9008_,
		_w9009_,
		_w9010_
	);
	LUT4 #(
		.INIT('h4000)
	) name8478 (
		_w8995_,
		_w8999_,
		_w9005_,
		_w9010_,
		_w9011_
	);
	LUT2 #(
		.INIT('h1)
	) name8479 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9012_
	);
	LUT4 #(
		.INIT('h0001)
	) name8480 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9013_
	);
	LUT2 #(
		.INIT('h4)
	) name8481 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9014_
	);
	LUT3 #(
		.INIT('h20)
	) name8482 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9015_
	);
	LUT4 #(
		.INIT('h0020)
	) name8483 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9016_
	);
	LUT2 #(
		.INIT('h4)
	) name8484 (
		\u0_w_reg[3][27]/P0001 ,
		_w9016_,
		_w9017_
	);
	LUT3 #(
		.INIT('h02)
	) name8485 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9018_
	);
	LUT4 #(
		.INIT('h0002)
	) name8486 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9019_
	);
	LUT2 #(
		.INIT('h8)
	) name8487 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w9020_
	);
	LUT3 #(
		.INIT('h80)
	) name8488 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9021_
	);
	LUT4 #(
		.INIT('h8000)
	) name8489 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9022_
	);
	LUT3 #(
		.INIT('h01)
	) name8490 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9023_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8491 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9024_
	);
	LUT3 #(
		.INIT('h04)
	) name8492 (
		_w9022_,
		_w9024_,
		_w9019_,
		_w9025_
	);
	LUT3 #(
		.INIT('h02)
	) name8493 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9026_
	);
	LUT4 #(
		.INIT('h0008)
	) name8494 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9027_
	);
	LUT4 #(
		.INIT('h1000)
	) name8495 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9028_
	);
	LUT2 #(
		.INIT('h1)
	) name8496 (
		_w9027_,
		_w9028_,
		_w9029_
	);
	LUT2 #(
		.INIT('h8)
	) name8497 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9030_
	);
	LUT4 #(
		.INIT('h0800)
	) name8498 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9031_
	);
	LUT4 #(
		.INIT('h0001)
	) name8499 (
		\u0_w_reg[3][26]/P0001 ,
		_w9031_,
		_w9027_,
		_w9028_,
		_w9032_
	);
	LUT4 #(
		.INIT('h5510)
	) name8500 (
		_w9013_,
		_w9017_,
		_w9025_,
		_w9032_,
		_w9033_
	);
	LUT4 #(
		.INIT('h0155)
	) name8501 (
		\u0_w_reg[3][24]/P0001 ,
		_w8991_,
		_w9011_,
		_w9033_,
		_w9034_
	);
	LUT3 #(
		.INIT('h08)
	) name8502 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9035_
	);
	LUT3 #(
		.INIT('h10)
	) name8503 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9036_
	);
	LUT4 #(
		.INIT('h0200)
	) name8504 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9037_
	);
	LUT4 #(
		.INIT('hfd3f)
	) name8505 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9038_
	);
	LUT2 #(
		.INIT('h1)
	) name8506 (
		\u0_w_reg[3][26]/P0001 ,
		_w9038_,
		_w9039_
	);
	LUT3 #(
		.INIT('h10)
	) name8507 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9040_
	);
	LUT4 #(
		.INIT('h0008)
	) name8508 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9041_
	);
	LUT3 #(
		.INIT('ha8)
	) name8509 (
		\u0_w_reg[3][26]/P0001 ,
		_w9040_,
		_w9041_,
		_w9042_
	);
	LUT4 #(
		.INIT('h0080)
	) name8510 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9043_
	);
	LUT4 #(
		.INIT('h4000)
	) name8511 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9044_
	);
	LUT3 #(
		.INIT('h13)
	) name8512 (
		\u0_w_reg[3][31]/P0001 ,
		_w9043_,
		_w9044_,
		_w9045_
	);
	LUT4 #(
		.INIT('h5455)
	) name8513 (
		\u0_w_reg[3][25]/P0001 ,
		_w9039_,
		_w9042_,
		_w9045_,
		_w9046_
	);
	LUT2 #(
		.INIT('h2)
	) name8514 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w9047_
	);
	LUT4 #(
		.INIT('h0200)
	) name8515 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9048_
	);
	LUT2 #(
		.INIT('h2)
	) name8516 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9049_
	);
	LUT3 #(
		.INIT('h08)
	) name8517 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9050_
	);
	LUT3 #(
		.INIT('h13)
	) name8518 (
		_w9049_,
		_w9048_,
		_w9050_,
		_w9051_
	);
	LUT3 #(
		.INIT('h20)
	) name8519 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9052_
	);
	LUT3 #(
		.INIT('h01)
	) name8520 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9053_
	);
	LUT3 #(
		.INIT('h57)
	) name8521 (
		_w8977_,
		_w9052_,
		_w9053_,
		_w9054_
	);
	LUT3 #(
		.INIT('h2a)
	) name8522 (
		\u0_w_reg[3][25]/P0001 ,
		_w9051_,
		_w9054_,
		_w9055_
	);
	LUT4 #(
		.INIT('h0020)
	) name8523 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9056_
	);
	LUT3 #(
		.INIT('h04)
	) name8524 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9057_
	);
	LUT4 #(
		.INIT('h2000)
	) name8525 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9058_
	);
	LUT4 #(
		.INIT('hdfbb)
	) name8526 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9059_
	);
	LUT4 #(
		.INIT('h5455)
	) name8527 (
		\u0_w_reg[3][26]/P0001 ,
		_w9043_,
		_w9056_,
		_w9059_,
		_w9060_
	);
	LUT4 #(
		.INIT('h0040)
	) name8528 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9061_
	);
	LUT2 #(
		.INIT('h8)
	) name8529 (
		\u0_w_reg[3][27]/P0001 ,
		_w9061_,
		_w9062_
	);
	LUT2 #(
		.INIT('h2)
	) name8530 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		_w9063_
	);
	LUT3 #(
		.INIT('h23)
	) name8531 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9064_
	);
	LUT4 #(
		.INIT('h0123)
	) name8532 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9065_
	);
	LUT3 #(
		.INIT('h20)
	) name8533 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		_w9066_
	);
	LUT3 #(
		.INIT('ha8)
	) name8534 (
		_w9063_,
		_w9065_,
		_w9066_,
		_w9067_
	);
	LUT2 #(
		.INIT('h2)
	) name8535 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w9068_
	);
	LUT4 #(
		.INIT('h8000)
	) name8536 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9069_
	);
	LUT4 #(
		.INIT('h0010)
	) name8537 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9070_
	);
	LUT4 #(
		.INIT('h7fef)
	) name8538 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9071_
	);
	LUT2 #(
		.INIT('h2)
	) name8539 (
		_w9068_,
		_w9071_,
		_w9072_
	);
	LUT4 #(
		.INIT('h0001)
	) name8540 (
		_w9060_,
		_w9062_,
		_w9067_,
		_w9072_,
		_w9073_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8541 (
		\u0_w_reg[3][24]/P0001 ,
		_w9055_,
		_w9046_,
		_w9073_,
		_w9074_
	);
	LUT4 #(
		.INIT('h0080)
	) name8542 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9075_
	);
	LUT3 #(
		.INIT('h04)
	) name8543 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9076_
	);
	LUT3 #(
		.INIT('h6b)
	) name8544 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9077_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name8545 (
		\u0_w_reg[3][26]/P0001 ,
		_w8977_,
		_w9075_,
		_w9077_,
		_w9078_
	);
	LUT4 #(
		.INIT('h0001)
	) name8546 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9079_
	);
	LUT3 #(
		.INIT('h54)
	) name8547 (
		\u0_w_reg[3][25]/P0001 ,
		_w9078_,
		_w9079_,
		_w9080_
	);
	LUT2 #(
		.INIT('h1)
	) name8548 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		_w9081_
	);
	LUT3 #(
		.INIT('h10)
	) name8549 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		_w9082_
	);
	LUT4 #(
		.INIT('h1000)
	) name8550 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9083_
	);
	LUT4 #(
		.INIT('h8000)
	) name8551 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9084_
	);
	LUT4 #(
		.INIT('h0023)
	) name8552 (
		\u0_w_reg[3][31]/P0001 ,
		_w9058_,
		_w9084_,
		_w9083_,
		_w9085_
	);
	LUT2 #(
		.INIT('h2)
	) name8553 (
		_w9081_,
		_w9085_,
		_w9086_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name8554 (
		\u0_w_reg[3][26]/P0001 ,
		_w9031_,
		_w9018_,
		_w8987_,
		_w9087_
	);
	LUT2 #(
		.INIT('h2)
	) name8555 (
		\u0_w_reg[3][25]/P0001 ,
		_w9087_,
		_w9088_
	);
	LUT2 #(
		.INIT('h4)
	) name8556 (
		\u0_w_reg[3][26]/P0001 ,
		_w8998_,
		_w9089_
	);
	LUT2 #(
		.INIT('h4)
	) name8557 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w9090_
	);
	LUT4 #(
		.INIT('h0004)
	) name8558 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9091_
	);
	LUT2 #(
		.INIT('h8)
	) name8559 (
		_w9090_,
		_w9091_,
		_w9092_
	);
	LUT4 #(
		.INIT('h0080)
	) name8560 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9093_
	);
	LUT2 #(
		.INIT('h2)
	) name8561 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9094_
	);
	LUT4 #(
		.INIT('h0020)
	) name8562 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9095_
	);
	LUT3 #(
		.INIT('h80)
	) name8563 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9096_
	);
	LUT4 #(
		.INIT('h0777)
	) name8564 (
		_w9093_,
		_w9094_,
		_w9095_,
		_w9096_,
		_w9097_
	);
	LUT3 #(
		.INIT('h10)
	) name8565 (
		_w9089_,
		_w9092_,
		_w9097_,
		_w9098_
	);
	LUT4 #(
		.INIT('h0100)
	) name8566 (
		_w9080_,
		_w9088_,
		_w9086_,
		_w9098_,
		_w9099_
	);
	LUT4 #(
		.INIT('h5655)
	) name8567 (
		\u0_w_reg[0][5]/P0001 ,
		_w9074_,
		_w9034_,
		_w9099_,
		_w9100_
	);
	LUT2 #(
		.INIT('h9)
	) name8568 (
		\u0_w_reg[1][5]/P0001 ,
		\u0_w_reg[2][5]/P0001 ,
		_w9101_
	);
	LUT4 #(
		.INIT('hb88b)
	) name8569 (
		\key[37]_pad ,
		ld_pad,
		_w9100_,
		_w9101_,
		_w9102_
	);
	LUT4 #(
		.INIT('ha955)
	) name8570 (
		\u0_w_reg[0][10]/P0001 ,
		_w8499_,
		_w8511_,
		_w8528_,
		_w9103_
	);
	LUT2 #(
		.INIT('h6)
	) name8571 (
		_w7817_,
		_w9103_,
		_w9104_
	);
	LUT3 #(
		.INIT('h69)
	) name8572 (
		_w7865_,
		_w8350_,
		_w8396_,
		_w9105_
	);
	LUT3 #(
		.INIT('h82)
	) name8573 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[106]/P0001 ,
		\u0_w_reg[0][10]/P0001 ,
		_w9106_
	);
	LUT4 #(
		.INIT('h00eb)
	) name8574 (
		\ld_r_reg/P0001 ,
		_w9104_,
		_w9105_,
		_w9106_,
		_w9107_
	);
	LUT4 #(
		.INIT('h0080)
	) name8575 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9108_
	);
	LUT3 #(
		.INIT('h07)
	) name8576 (
		\u0_w_reg[3][22]/P0001 ,
		_w8734_,
		_w9108_,
		_w9109_
	);
	LUT4 #(
		.INIT('h0015)
	) name8577 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8734_,
		_w9108_,
		_w9110_
	);
	LUT3 #(
		.INIT('h40)
	) name8578 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w9111_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name8579 (
		\u0_w_reg[3][17]/P0001 ,
		_w8721_,
		_w8693_,
		_w9111_,
		_w9112_
	);
	LUT4 #(
		.INIT('h0002)
	) name8580 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9113_
	);
	LUT4 #(
		.INIT('h4000)
	) name8581 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9114_
	);
	LUT3 #(
		.INIT('h02)
	) name8582 (
		\u0_w_reg[3][18]/P0001 ,
		_w9113_,
		_w9114_,
		_w9115_
	);
	LUT3 #(
		.INIT('h45)
	) name8583 (
		_w9110_,
		_w9112_,
		_w9115_,
		_w9116_
	);
	LUT2 #(
		.INIT('h4)
	) name8584 (
		\u0_w_reg[3][18]/P0001 ,
		_w8669_,
		_w9117_
	);
	LUT3 #(
		.INIT('h2a)
	) name8585 (
		\u0_w_reg[3][17]/P0001 ,
		_w8657_,
		_w8687_,
		_w9118_
	);
	LUT4 #(
		.INIT('h0200)
	) name8586 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9119_
	);
	LUT4 #(
		.INIT('h8000)
	) name8587 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9120_
	);
	LUT3 #(
		.INIT('h13)
	) name8588 (
		\u0_w_reg[3][20]/P0001 ,
		_w9119_,
		_w9120_,
		_w9121_
	);
	LUT3 #(
		.INIT('h40)
	) name8589 (
		_w9117_,
		_w9118_,
		_w9121_,
		_w9122_
	);
	LUT3 #(
		.INIT('h40)
	) name8590 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w8708_,
		_w9123_
	);
	LUT3 #(
		.INIT('hf4)
	) name8591 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w9124_
	);
	LUT2 #(
		.INIT('h2)
	) name8592 (
		_w8670_,
		_w9124_,
		_w9125_
	);
	LUT3 #(
		.INIT('h20)
	) name8593 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9126_
	);
	LUT4 #(
		.INIT('h0100)
	) name8594 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9127_
	);
	LUT4 #(
		.INIT('h0405)
	) name8595 (
		\u0_w_reg[3][17]/P0001 ,
		_w8665_,
		_w9127_,
		_w9126_,
		_w9128_
	);
	LUT3 #(
		.INIT('h10)
	) name8596 (
		_w9125_,
		_w9123_,
		_w9128_,
		_w9129_
	);
	LUT2 #(
		.INIT('h4)
	) name8597 (
		\u0_w_reg[3][21]/P0001 ,
		_w8658_,
		_w9130_
	);
	LUT4 #(
		.INIT('h000e)
	) name8598 (
		_w9122_,
		_w9129_,
		_w9116_,
		_w9130_,
		_w9131_
	);
	LUT4 #(
		.INIT('h0c04)
	) name8599 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9132_
	);
	LUT3 #(
		.INIT('ha8)
	) name8600 (
		\u0_w_reg[3][17]/P0001 ,
		_w8684_,
		_w9132_,
		_w9133_
	);
	LUT3 #(
		.INIT('h80)
	) name8601 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9134_
	);
	LUT4 #(
		.INIT('h0800)
	) name8602 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9135_
	);
	LUT4 #(
		.INIT('hfddf)
	) name8603 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9136_
	);
	LUT2 #(
		.INIT('h4)
	) name8604 (
		_w9135_,
		_w9136_,
		_w9137_
	);
	LUT3 #(
		.INIT('h8a)
	) name8605 (
		\u0_w_reg[3][18]/P0001 ,
		_w9133_,
		_w9137_,
		_w9138_
	);
	LUT4 #(
		.INIT('hff3b)
	) name8606 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9139_
	);
	LUT3 #(
		.INIT('h8a)
	) name8607 (
		\u0_w_reg[3][18]/P0001 ,
		_w9119_,
		_w9139_,
		_w9140_
	);
	LUT4 #(
		.INIT('h0105)
	) name8608 (
		_w8663_,
		_w8675_,
		_w8751_,
		_w8772_,
		_w9141_
	);
	LUT4 #(
		.INIT('h153f)
	) name8609 (
		_w8729_,
		_w8723_,
		_w8683_,
		_w8752_,
		_w9142_
	);
	LUT4 #(
		.INIT('h4555)
	) name8610 (
		\u0_w_reg[3][17]/P0001 ,
		_w9140_,
		_w9141_,
		_w9142_,
		_w9143_
	);
	LUT4 #(
		.INIT('h0001)
	) name8611 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9144_
	);
	LUT4 #(
		.INIT('h2000)
	) name8612 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9145_
	);
	LUT4 #(
		.INIT('h0010)
	) name8613 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9146_
	);
	LUT4 #(
		.INIT('h0001)
	) name8614 (
		_w8734_,
		_w8708_,
		_w9145_,
		_w9146_,
		_w9147_
	);
	LUT3 #(
		.INIT('h8a)
	) name8615 (
		\u0_w_reg[3][17]/P0001 ,
		_w9144_,
		_w9147_,
		_w9148_
	);
	LUT3 #(
		.INIT('h54)
	) name8616 (
		\u0_w_reg[3][18]/P0001 ,
		_w9127_,
		_w9120_,
		_w9149_
	);
	LUT2 #(
		.INIT('h8)
	) name8617 (
		_w8656_,
		_w8715_,
		_w9150_
	);
	LUT3 #(
		.INIT('h10)
	) name8618 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w8734_,
		_w9151_
	);
	LUT3 #(
		.INIT('h01)
	) name8619 (
		_w9150_,
		_w9151_,
		_w9149_,
		_w9152_
	);
	LUT4 #(
		.INIT('h0100)
	) name8620 (
		_w9143_,
		_w9148_,
		_w9138_,
		_w9152_,
		_w9153_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name8621 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9154_
	);
	LUT2 #(
		.INIT('h2)
	) name8622 (
		_w8764_,
		_w9154_,
		_w9155_
	);
	LUT3 #(
		.INIT('ha8)
	) name8623 (
		\u0_w_reg[3][18]/P0001 ,
		_w8708_,
		_w9145_,
		_w9156_
	);
	LUT3 #(
		.INIT('h08)
	) name8624 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w9157_
	);
	LUT2 #(
		.INIT('h4)
	) name8625 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9158_
	);
	LUT4 #(
		.INIT('h0100)
	) name8626 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9159_
	);
	LUT2 #(
		.INIT('h8)
	) name8627 (
		_w8729_,
		_w9159_,
		_w9160_
	);
	LUT4 #(
		.INIT('h135f)
	) name8628 (
		_w8662_,
		_w8729_,
		_w9157_,
		_w9159_,
		_w9161_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8629 (
		\u0_w_reg[3][17]/P0001 ,
		_w9156_,
		_w9155_,
		_w9161_,
		_w9162_
	);
	LUT3 #(
		.INIT('h04)
	) name8630 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w9163_
	);
	LUT4 #(
		.INIT('h0010)
	) name8631 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9164_
	);
	LUT4 #(
		.INIT('h0002)
	) name8632 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9165_
	);
	LUT4 #(
		.INIT('hffed)
	) name8633 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9166_
	);
	LUT2 #(
		.INIT('h2)
	) name8634 (
		_w9163_,
		_w9166_,
		_w9167_
	);
	LUT3 #(
		.INIT('h10)
	) name8635 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w9168_
	);
	LUT4 #(
		.INIT('h135f)
	) name8636 (
		\u0_w_reg[3][18]/P0001 ,
		_w8675_,
		_w9145_,
		_w9168_,
		_w9169_
	);
	LUT2 #(
		.INIT('h4)
	) name8637 (
		\u0_w_reg[3][21]/P0001 ,
		_w9108_,
		_w9170_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name8638 (
		\u0_w_reg[3][21]/P0001 ,
		_w8685_,
		_w8689_,
		_w9108_,
		_w9171_
	);
	LUT4 #(
		.INIT('h0e00)
	) name8639 (
		\u0_w_reg[3][20]/P0001 ,
		_w9169_,
		_w9167_,
		_w9171_,
		_w9172_
	);
	LUT2 #(
		.INIT('h4)
	) name8640 (
		_w9162_,
		_w9172_,
		_w9173_
	);
	LUT4 #(
		.INIT('hd800)
	) name8641 (
		\u0_w_reg[3][16]/P0001 ,
		_w9153_,
		_w9131_,
		_w9173_,
		_w9174_
	);
	LUT2 #(
		.INIT('h9)
	) name8642 (
		\u0_r0_out_reg[27]/P0001 ,
		\u0_w_reg[0][27]/P0001 ,
		_w9175_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name8643 (
		\key[123]_pad ,
		ld_pad,
		_w9174_,
		_w9175_,
		_w9176_
	);
	LUT3 #(
		.INIT('h96)
	) name8644 (
		\u0_r0_out_reg[27]/P0001 ,
		\u0_w_reg[0][27]/P0001 ,
		\u0_w_reg[1][27]/P0001 ,
		_w9177_
	);
	LUT4 #(
		.INIT('hb88b)
	) name8645 (
		\key[91]_pad ,
		ld_pad,
		_w9174_,
		_w9177_,
		_w9178_
	);
	LUT2 #(
		.INIT('h4)
	) name8646 (
		\key[59]_pad ,
		ld_pad,
		_w9179_
	);
	LUT3 #(
		.INIT('h96)
	) name8647 (
		\u0_w_reg[2][27]/P0001 ,
		_w9174_,
		_w9177_,
		_w9180_
	);
	LUT4 #(
		.INIT('h4114)
	) name8648 (
		ld_pad,
		\u0_w_reg[2][27]/P0001 ,
		_w9174_,
		_w9177_,
		_w9181_
	);
	LUT2 #(
		.INIT('h1)
	) name8649 (
		_w9179_,
		_w9181_,
		_w9182_
	);
	LUT4 #(
		.INIT('hb88b)
	) name8650 (
		\key[27]_pad ,
		ld_pad,
		\u0_w_reg[3][27]/P0001 ,
		_w9180_,
		_w9183_
	);
	LUT3 #(
		.INIT('h8a)
	) name8651 (
		\u0_w_reg[3][26]/P0001 ,
		_w9057_,
		_w9038_,
		_w9184_
	);
	LUT4 #(
		.INIT('h0105)
	) name8652 (
		\u0_w_reg[3][25]/P0001 ,
		_w9076_,
		_w9079_,
		_w9090_,
		_w9185_
	);
	LUT4 #(
		.INIT('h1000)
	) name8653 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9186_
	);
	LUT3 #(
		.INIT('h07)
	) name8654 (
		_w8987_,
		_w9021_,
		_w9186_,
		_w9187_
	);
	LUT4 #(
		.INIT('h1000)
	) name8655 (
		_w9089_,
		_w9184_,
		_w9185_,
		_w9187_,
		_w9188_
	);
	LUT3 #(
		.INIT('h20)
	) name8656 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9189_
	);
	LUT4 #(
		.INIT('h0c04)
	) name8657 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9190_
	);
	LUT3 #(
		.INIT('ha8)
	) name8658 (
		\u0_w_reg[3][26]/P0001 ,
		_w9189_,
		_w9190_,
		_w9191_
	);
	LUT4 #(
		.INIT('h0001)
	) name8659 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9192_
	);
	LUT2 #(
		.INIT('h2)
	) name8660 (
		\u0_w_reg[3][25]/P0001 ,
		_w9192_,
		_w9193_
	);
	LUT2 #(
		.INIT('h8)
	) name8661 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9194_
	);
	LUT4 #(
		.INIT('h2000)
	) name8662 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9195_
	);
	LUT4 #(
		.INIT('h4000)
	) name8663 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9196_
	);
	LUT2 #(
		.INIT('h1)
	) name8664 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w9197_
	);
	LUT4 #(
		.INIT('h0010)
	) name8665 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9198_
	);
	LUT4 #(
		.INIT('h0001)
	) name8666 (
		_w9031_,
		_w9196_,
		_w9198_,
		_w9195_,
		_w9199_
	);
	LUT3 #(
		.INIT('h20)
	) name8667 (
		_w9193_,
		_w9191_,
		_w9199_,
		_w9200_
	);
	LUT4 #(
		.INIT('h8000)
	) name8668 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9201_
	);
	LUT3 #(
		.INIT('h07)
	) name8669 (
		_w8977_,
		_w9052_,
		_w9201_,
		_w9202_
	);
	LUT3 #(
		.INIT('h10)
	) name8670 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9203_
	);
	LUT4 #(
		.INIT('h0100)
	) name8671 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9204_
	);
	LUT2 #(
		.INIT('h1)
	) name8672 (
		\u0_w_reg[3][26]/P0001 ,
		_w9204_,
		_w9205_
	);
	LUT4 #(
		.INIT('h0800)
	) name8673 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9206_
	);
	LUT4 #(
		.INIT('h0200)
	) name8674 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9207_
	);
	LUT4 #(
		.INIT('h0002)
	) name8675 (
		\u0_w_reg[3][26]/P0001 ,
		_w9016_,
		_w9207_,
		_w9206_,
		_w9208_
	);
	LUT4 #(
		.INIT('h5540)
	) name8676 (
		_w9062_,
		_w9202_,
		_w9205_,
		_w9208_,
		_w9209_
	);
	LUT4 #(
		.INIT('h02aa)
	) name8677 (
		\u0_w_reg[3][24]/P0001 ,
		_w9188_,
		_w9200_,
		_w9209_,
		_w9210_
	);
	LUT3 #(
		.INIT('h01)
	) name8678 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9211_
	);
	LUT4 #(
		.INIT('h0040)
	) name8679 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9212_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name8680 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9211_,
		_w9212_,
		_w9213_
	);
	LUT2 #(
		.INIT('h2)
	) name8681 (
		\u0_w_reg[3][25]/P0001 ,
		_w9037_,
		_w9214_
	);
	LUT2 #(
		.INIT('h6)
	) name8682 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w9215_
	);
	LUT4 #(
		.INIT('haf23)
	) name8683 (
		\u0_w_reg[3][26]/P0001 ,
		_w8984_,
		_w9004_,
		_w9215_,
		_w9216_
	);
	LUT3 #(
		.INIT('h40)
	) name8684 (
		_w9213_,
		_w9214_,
		_w9216_,
		_w9217_
	);
	LUT3 #(
		.INIT('h40)
	) name8685 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w9031_,
		_w9218_
	);
	LUT2 #(
		.INIT('h1)
	) name8686 (
		\u0_w_reg[3][25]/P0001 ,
		_w9204_,
		_w9219_
	);
	LUT3 #(
		.INIT('h20)
	) name8687 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9220_
	);
	LUT4 #(
		.INIT('h0a1f)
	) name8688 (
		_w8987_,
		_w9094_,
		_w9006_,
		_w9220_,
		_w9221_
	);
	LUT3 #(
		.INIT('h40)
	) name8689 (
		_w9218_,
		_w9219_,
		_w9221_,
		_w9222_
	);
	LUT4 #(
		.INIT('h4000)
	) name8690 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9223_
	);
	LUT3 #(
		.INIT('ha8)
	) name8691 (
		\u0_w_reg[3][26]/P0001 ,
		_w9019_,
		_w9223_,
		_w9224_
	);
	LUT4 #(
		.INIT('h0080)
	) name8692 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9225_
	);
	LUT4 #(
		.INIT('h5540)
	) name8693 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9044_,
		_w9225_,
		_w9226_
	);
	LUT2 #(
		.INIT('h4)
	) name8694 (
		\u0_w_reg[3][27]/P0001 ,
		_w9070_,
		_w9227_
	);
	LUT3 #(
		.INIT('h01)
	) name8695 (
		_w9226_,
		_w9224_,
		_w9227_,
		_w9228_
	);
	LUT4 #(
		.INIT('h0155)
	) name8696 (
		\u0_w_reg[3][24]/P0001 ,
		_w9217_,
		_w9222_,
		_w9228_,
		_w9229_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name8697 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9230_
	);
	LUT2 #(
		.INIT('h2)
	) name8698 (
		_w9197_,
		_w9230_,
		_w9231_
	);
	LUT3 #(
		.INIT('ha8)
	) name8699 (
		\u0_w_reg[3][26]/P0001 ,
		_w9031_,
		_w9195_,
		_w9232_
	);
	LUT4 #(
		.INIT('h0100)
	) name8700 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9233_
	);
	LUT4 #(
		.INIT('h135f)
	) name8701 (
		_w9047_,
		_w9090_,
		_w9007_,
		_w9233_,
		_w9234_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8702 (
		\u0_w_reg[3][25]/P0001 ,
		_w9232_,
		_w9231_,
		_w9234_,
		_w9235_
	);
	LUT4 #(
		.INIT('habaf)
	) name8703 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w9070_,
		_w9053_,
		_w9236_
	);
	LUT2 #(
		.INIT('h4)
	) name8704 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		_w9237_
	);
	LUT2 #(
		.INIT('h4)
	) name8705 (
		_w9236_,
		_w9237_,
		_w9238_
	);
	LUT4 #(
		.INIT('h2000)
	) name8706 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9239_
	);
	LUT4 #(
		.INIT('h1000)
	) name8707 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9240_
	);
	LUT3 #(
		.INIT('ha8)
	) name8708 (
		_w9047_,
		_w9239_,
		_w9240_,
		_w9241_
	);
	LUT2 #(
		.INIT('h8)
	) name8709 (
		_w9026_,
		_w9194_,
		_w9242_
	);
	LUT3 #(
		.INIT('h80)
	) name8710 (
		\u0_w_reg[3][26]/P0001 ,
		_w8987_,
		_w9021_,
		_w9243_
	);
	LUT3 #(
		.INIT('h01)
	) name8711 (
		_w9242_,
		_w9241_,
		_w9243_,
		_w9244_
	);
	LUT3 #(
		.INIT('h10)
	) name8712 (
		_w9235_,
		_w9238_,
		_w9244_,
		_w9245_
	);
	LUT4 #(
		.INIT('h5655)
	) name8713 (
		\u0_w_reg[0][3]/P0001 ,
		_w9210_,
		_w9229_,
		_w9245_,
		_w9246_
	);
	LUT2 #(
		.INIT('h9)
	) name8714 (
		\u0_w_reg[1][3]/P0001 ,
		\u0_w_reg[2][3]/P0001 ,
		_w9247_
	);
	LUT4 #(
		.INIT('hb88b)
	) name8715 (
		\key[35]_pad ,
		ld_pad,
		_w9246_,
		_w9247_,
		_w9248_
	);
	LUT2 #(
		.INIT('h1)
	) name8716 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9249_
	);
	LUT3 #(
		.INIT('h01)
	) name8717 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9250_
	);
	LUT4 #(
		.INIT('h0040)
	) name8718 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9251_
	);
	LUT4 #(
		.INIT('ha820)
	) name8719 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w9249_,
		_w9251_,
		_w9252_
	);
	LUT2 #(
		.INIT('h8)
	) name8720 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9253_
	);
	LUT2 #(
		.INIT('h4)
	) name8721 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9254_
	);
	LUT4 #(
		.INIT('h4000)
	) name8722 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9255_
	);
	LUT2 #(
		.INIT('h8)
	) name8723 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9256_
	);
	LUT4 #(
		.INIT('h0200)
	) name8724 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9257_
	);
	LUT4 #(
		.INIT('h008a)
	) name8725 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w9255_,
		_w9257_,
		_w9258_
	);
	LUT2 #(
		.INIT('h2)
	) name8726 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9259_
	);
	LUT4 #(
		.INIT('h0400)
	) name8727 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9260_
	);
	LUT2 #(
		.INIT('h8)
	) name8728 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9261_
	);
	LUT3 #(
		.INIT('h80)
	) name8729 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9262_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name8730 (
		\u0_w_reg[3][2]/P0001 ,
		_w9260_,
		_w9261_,
		_w9262_,
		_w9263_
	);
	LUT3 #(
		.INIT('h40)
	) name8731 (
		_w9252_,
		_w9258_,
		_w9263_,
		_w9264_
	);
	LUT3 #(
		.INIT('h10)
	) name8732 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9265_
	);
	LUT4 #(
		.INIT('h0100)
	) name8733 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9266_
	);
	LUT2 #(
		.INIT('h1)
	) name8734 (
		\u0_w_reg[3][1]/P0001 ,
		_w9266_,
		_w9267_
	);
	LUT2 #(
		.INIT('h2)
	) name8735 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w9268_
	);
	LUT3 #(
		.INIT('he0)
	) name8736 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9269_
	);
	LUT2 #(
		.INIT('h8)
	) name8737 (
		_w9268_,
		_w9269_,
		_w9270_
	);
	LUT2 #(
		.INIT('h2)
	) name8738 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9271_
	);
	LUT2 #(
		.INIT('h2)
	) name8739 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9272_
	);
	LUT3 #(
		.INIT('hf4)
	) name8740 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9273_
	);
	LUT2 #(
		.INIT('h4)
	) name8741 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w9274_
	);
	LUT4 #(
		.INIT('h4000)
	) name8742 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9275_
	);
	LUT2 #(
		.INIT('h8)
	) name8743 (
		_w9259_,
		_w9275_,
		_w9276_
	);
	LUT4 #(
		.INIT('h51f3)
	) name8744 (
		_w9259_,
		_w9271_,
		_w9273_,
		_w9275_,
		_w9277_
	);
	LUT3 #(
		.INIT('h40)
	) name8745 (
		_w9270_,
		_w9267_,
		_w9277_,
		_w9278_
	);
	LUT4 #(
		.INIT('h4000)
	) name8746 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9279_
	);
	LUT2 #(
		.INIT('h8)
	) name8747 (
		\u0_w_reg[3][6]/P0001 ,
		_w9279_,
		_w9280_
	);
	LUT3 #(
		.INIT('h08)
	) name8748 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9281_
	);
	LUT4 #(
		.INIT('h0080)
	) name8749 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9282_
	);
	LUT3 #(
		.INIT('h07)
	) name8750 (
		\u0_w_reg[3][6]/P0001 ,
		_w9279_,
		_w9282_,
		_w9283_
	);
	LUT4 #(
		.INIT('h4440)
	) name8751 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9279_,
		_w9281_,
		_w9284_
	);
	LUT2 #(
		.INIT('h1)
	) name8752 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w9285_
	);
	LUT2 #(
		.INIT('h4)
	) name8753 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9286_
	);
	LUT3 #(
		.INIT('h04)
	) name8754 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9287_
	);
	LUT3 #(
		.INIT('h15)
	) name8755 (
		\u0_w_reg[3][0]/P0001 ,
		_w9285_,
		_w9287_,
		_w9288_
	);
	LUT2 #(
		.INIT('h8)
	) name8756 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w9289_
	);
	LUT3 #(
		.INIT('h80)
	) name8757 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9290_
	);
	LUT4 #(
		.INIT('h153f)
	) name8758 (
		_w9254_,
		_w9250_,
		_w9289_,
		_w9290_,
		_w9291_
	);
	LUT3 #(
		.INIT('h40)
	) name8759 (
		_w9284_,
		_w9288_,
		_w9291_,
		_w9292_
	);
	LUT3 #(
		.INIT('he0)
	) name8760 (
		_w9264_,
		_w9278_,
		_w9292_,
		_w9293_
	);
	LUT3 #(
		.INIT('h20)
	) name8761 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9294_
	);
	LUT4 #(
		.INIT('h0c04)
	) name8762 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9295_
	);
	LUT3 #(
		.INIT('ha8)
	) name8763 (
		\u0_w_reg[3][2]/P0001 ,
		_w9294_,
		_w9295_,
		_w9296_
	);
	LUT2 #(
		.INIT('h8)
	) name8764 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9297_
	);
	LUT3 #(
		.INIT('h4c)
	) name8765 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9298_
	);
	LUT2 #(
		.INIT('h8)
	) name8766 (
		_w9253_,
		_w9298_,
		_w9299_
	);
	LUT4 #(
		.INIT('h2000)
	) name8767 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9300_
	);
	LUT2 #(
		.INIT('h1)
	) name8768 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9301_
	);
	LUT4 #(
		.INIT('h0001)
	) name8769 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9302_
	);
	LUT2 #(
		.INIT('h1)
	) name8770 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w9303_
	);
	LUT4 #(
		.INIT('h0010)
	) name8771 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9304_
	);
	LUT3 #(
		.INIT('h01)
	) name8772 (
		_w9302_,
		_w9304_,
		_w9300_,
		_w9305_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8773 (
		\u0_w_reg[3][1]/P0001 ,
		_w9299_,
		_w9296_,
		_w9305_,
		_w9306_
	);
	LUT3 #(
		.INIT('h40)
	) name8774 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9307_
	);
	LUT4 #(
		.INIT('h1000)
	) name8775 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9308_
	);
	LUT4 #(
		.INIT('h0020)
	) name8776 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9309_
	);
	LUT4 #(
		.INIT('hefdf)
	) name8777 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9310_
	);
	LUT2 #(
		.INIT('h1)
	) name8778 (
		\u0_w_reg[3][2]/P0001 ,
		_w9310_,
		_w9311_
	);
	LUT2 #(
		.INIT('h1)
	) name8779 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w9312_
	);
	LUT2 #(
		.INIT('h2)
	) name8780 (
		_w9257_,
		_w9312_,
		_w9313_
	);
	LUT2 #(
		.INIT('h1)
	) name8781 (
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9314_
	);
	LUT4 #(
		.INIT('h0001)
	) name8782 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9315_
	);
	LUT4 #(
		.INIT('h0080)
	) name8783 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9316_
	);
	LUT2 #(
		.INIT('h2)
	) name8784 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w9317_
	);
	LUT4 #(
		.INIT('h0020)
	) name8785 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9318_
	);
	LUT4 #(
		.INIT('h1000)
	) name8786 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9319_
	);
	LUT4 #(
		.INIT('h0001)
	) name8787 (
		_w9315_,
		_w9316_,
		_w9318_,
		_w9319_,
		_w9320_
	);
	LUT4 #(
		.INIT('h5455)
	) name8788 (
		\u0_w_reg[3][1]/P0001 ,
		_w9311_,
		_w9313_,
		_w9320_,
		_w9321_
	);
	LUT4 #(
		.INIT('h0800)
	) name8789 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9322_
	);
	LUT3 #(
		.INIT('h80)
	) name8790 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9323_
	);
	LUT4 #(
		.INIT('h8000)
	) name8791 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9324_
	);
	LUT3 #(
		.INIT('h0b)
	) name8792 (
		\u0_w_reg[3][3]/P0001 ,
		_w9322_,
		_w9324_,
		_w9325_
	);
	LUT2 #(
		.INIT('h1)
	) name8793 (
		\u0_w_reg[3][2]/P0001 ,
		_w9266_,
		_w9326_
	);
	LUT4 #(
		.INIT('h0020)
	) name8794 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9327_
	);
	LUT4 #(
		.INIT('h0200)
	) name8795 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9328_
	);
	LUT2 #(
		.INIT('h4)
	) name8796 (
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9329_
	);
	LUT4 #(
		.INIT('h0800)
	) name8797 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9330_
	);
	LUT4 #(
		.INIT('h0002)
	) name8798 (
		\u0_w_reg[3][2]/P0001 ,
		_w9330_,
		_w9327_,
		_w9328_,
		_w9331_
	);
	LUT3 #(
		.INIT('h04)
	) name8799 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9332_
	);
	LUT3 #(
		.INIT('h2a)
	) name8800 (
		\u0_w_reg[3][0]/P0001 ,
		_w9297_,
		_w9332_,
		_w9333_
	);
	LUT4 #(
		.INIT('hf800)
	) name8801 (
		_w9325_,
		_w9326_,
		_w9331_,
		_w9333_,
		_w9334_
	);
	LUT3 #(
		.INIT('h10)
	) name8802 (
		_w9321_,
		_w9306_,
		_w9334_,
		_w9335_
	);
	LUT3 #(
		.INIT('h02)
	) name8803 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9336_
	);
	LUT4 #(
		.INIT('hf9ad)
	) name8804 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9337_
	);
	LUT2 #(
		.INIT('h2)
	) name8805 (
		_w9303_,
		_w9337_,
		_w9338_
	);
	LUT2 #(
		.INIT('h2)
	) name8806 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w9339_
	);
	LUT4 #(
		.INIT('h2000)
	) name8807 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9340_
	);
	LUT3 #(
		.INIT('ha8)
	) name8808 (
		\u0_w_reg[3][2]/P0001 ,
		_w9322_,
		_w9340_,
		_w9341_
	);
	LUT4 #(
		.INIT('h153f)
	) name8809 (
		_w9257_,
		_w9289_,
		_w9307_,
		_w9312_,
		_w9342_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8810 (
		\u0_w_reg[3][1]/P0001 ,
		_w9338_,
		_w9341_,
		_w9342_,
		_w9343_
	);
	LUT2 #(
		.INIT('h4)
	) name8811 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		_w9344_
	);
	LUT3 #(
		.INIT('h01)
	) name8812 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9345_
	);
	LUT4 #(
		.INIT('h0001)
	) name8813 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9346_
	);
	LUT2 #(
		.INIT('h8)
	) name8814 (
		\u0_w_reg[3][4]/P0001 ,
		_w9346_,
		_w9347_
	);
	LUT4 #(
		.INIT('h23ef)
	) name8815 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w9287_,
		_w9346_,
		_w9348_
	);
	LUT4 #(
		.INIT('h0008)
	) name8816 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9349_
	);
	LUT2 #(
		.INIT('h8)
	) name8817 (
		\u0_w_reg[3][6]/P0001 ,
		_w9349_,
		_w9350_
	);
	LUT2 #(
		.INIT('h1)
	) name8818 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		_w9351_
	);
	LUT4 #(
		.INIT('h2000)
	) name8819 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9352_
	);
	LUT4 #(
		.INIT('h1000)
	) name8820 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9353_
	);
	LUT4 #(
		.INIT('hedff)
	) name8821 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9354_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8822 (
		_w9289_,
		_w9351_,
		_w9352_,
		_w9354_,
		_w9355_
	);
	LUT4 #(
		.INIT('h0d00)
	) name8823 (
		_w9344_,
		_w9348_,
		_w9350_,
		_w9355_,
		_w9356_
	);
	LUT2 #(
		.INIT('h4)
	) name8824 (
		_w9343_,
		_w9356_,
		_w9357_
	);
	LUT4 #(
		.INIT('ha955)
	) name8825 (
		\u0_w_reg[0][11]/P0001 ,
		_w9293_,
		_w9335_,
		_w9357_,
		_w9358_
	);
	LUT2 #(
		.INIT('h9)
	) name8826 (
		\u0_w_reg[1][11]/P0001 ,
		\u0_w_reg[2][11]/P0001 ,
		_w9359_
	);
	LUT4 #(
		.INIT('hb88b)
	) name8827 (
		\key[43]_pad ,
		ld_pad,
		_w9358_,
		_w9359_,
		_w9360_
	);
	LUT2 #(
		.INIT('h4)
	) name8828 (
		\key[44]_pad ,
		ld_pad,
		_w9361_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name8829 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9362_
	);
	LUT2 #(
		.INIT('h1)
	) name8830 (
		\u0_w_reg[3][2]/P0001 ,
		_w9362_,
		_w9363_
	);
	LUT4 #(
		.INIT('h0200)
	) name8831 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9364_
	);
	LUT2 #(
		.INIT('h1)
	) name8832 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9365_
	);
	LUT3 #(
		.INIT('h02)
	) name8833 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9366_
	);
	LUT3 #(
		.INIT('h13)
	) name8834 (
		_w9259_,
		_w9364_,
		_w9366_,
		_w9367_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8835 (
		\u0_w_reg[3][1]/P0001 ,
		_w9347_,
		_w9363_,
		_w9367_,
		_w9368_
	);
	LUT3 #(
		.INIT('h40)
	) name8836 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9369_
	);
	LUT4 #(
		.INIT('h0008)
	) name8837 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9370_
	);
	LUT3 #(
		.INIT('h54)
	) name8838 (
		\u0_w_reg[3][2]/P0001 ,
		_w9369_,
		_w9370_,
		_w9371_
	);
	LUT3 #(
		.INIT('h23)
	) name8839 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9372_
	);
	LUT2 #(
		.INIT('h2)
	) name8840 (
		_w9256_,
		_w9372_,
		_w9373_
	);
	LUT3 #(
		.INIT('h54)
	) name8841 (
		\u0_w_reg[3][1]/P0001 ,
		_w9371_,
		_w9373_,
		_w9374_
	);
	LUT2 #(
		.INIT('h4)
	) name8842 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w9375_
	);
	LUT3 #(
		.INIT('h04)
	) name8843 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9376_
	);
	LUT4 #(
		.INIT('h0023)
	) name8844 (
		\u0_w_reg[3][1]/P0001 ,
		_w9257_,
		_w9322_,
		_w9376_,
		_w9377_
	);
	LUT4 #(
		.INIT('h0001)
	) name8845 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9378_
	);
	LUT4 #(
		.INIT('h0020)
	) name8846 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9379_
	);
	LUT4 #(
		.INIT('h0203)
	) name8847 (
		\u0_w_reg[3][3]/P0001 ,
		_w9300_,
		_w9379_,
		_w9378_,
		_w9380_
	);
	LUT3 #(
		.INIT('h08)
	) name8848 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w9381_
	);
	LUT4 #(
		.INIT('h0008)
	) name8849 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9382_
	);
	LUT4 #(
		.INIT('h002a)
	) name8850 (
		\u0_w_reg[3][0]/P0001 ,
		_w9254_,
		_w9290_,
		_w9382_,
		_w9383_
	);
	LUT4 #(
		.INIT('he400)
	) name8851 (
		\u0_w_reg[3][2]/P0001 ,
		_w9380_,
		_w9377_,
		_w9383_,
		_w9384_
	);
	LUT3 #(
		.INIT('h10)
	) name8852 (
		_w9374_,
		_w9368_,
		_w9384_,
		_w9385_
	);
	LUT4 #(
		.INIT('h0100)
	) name8853 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9386_
	);
	LUT3 #(
		.INIT('h20)
	) name8854 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9387_
	);
	LUT4 #(
		.INIT('h5150)
	) name8855 (
		\u0_w_reg[3][2]/P0001 ,
		_w9339_,
		_w9386_,
		_w9387_,
		_w9388_
	);
	LUT4 #(
		.INIT('h0103)
	) name8856 (
		_w9268_,
		_w9282_,
		_w9316_,
		_w9294_,
		_w9389_
	);
	LUT3 #(
		.INIT('h8a)
	) name8857 (
		\u0_w_reg[3][1]/P0001 ,
		_w9388_,
		_w9389_,
		_w9390_
	);
	LUT2 #(
		.INIT('h8)
	) name8858 (
		\u0_w_reg[3][5]/P0001 ,
		_w9304_,
		_w9391_
	);
	LUT3 #(
		.INIT('h80)
	) name8859 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9392_
	);
	LUT4 #(
		.INIT('h8000)
	) name8860 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9393_
	);
	LUT2 #(
		.INIT('h2)
	) name8861 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		_w9394_
	);
	LUT4 #(
		.INIT('hf351)
	) name8862 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		_w9395_
	);
	LUT3 #(
		.INIT('h31)
	) name8863 (
		_w9314_,
		_w9393_,
		_w9395_,
		_w9396_
	);
	LUT3 #(
		.INIT('h45)
	) name8864 (
		\u0_w_reg[3][1]/P0001 ,
		_w9391_,
		_w9396_,
		_w9397_
	);
	LUT4 #(
		.INIT('h0004)
	) name8865 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9398_
	);
	LUT4 #(
		.INIT('h5540)
	) name8866 (
		\u0_w_reg[3][3]/P0001 ,
		_w9274_,
		_w9307_,
		_w9398_,
		_w9399_
	);
	LUT3 #(
		.INIT('h10)
	) name8867 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9400_
	);
	LUT4 #(
		.INIT('h0002)
	) name8868 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9401_
	);
	LUT3 #(
		.INIT('ha2)
	) name8869 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w9402_
	);
	LUT4 #(
		.INIT('h0155)
	) name8870 (
		\u0_w_reg[3][0]/P0001 ,
		_w9400_,
		_w9401_,
		_w9402_,
		_w9403_
	);
	LUT2 #(
		.INIT('h4)
	) name8871 (
		_w9399_,
		_w9403_,
		_w9404_
	);
	LUT3 #(
		.INIT('h10)
	) name8872 (
		_w9397_,
		_w9390_,
		_w9404_,
		_w9405_
	);
	LUT4 #(
		.INIT('haa80)
	) name8873 (
		\u0_w_reg[3][3]/P0001 ,
		_w9287_,
		_w9312_,
		_w9393_,
		_w9406_
	);
	LUT3 #(
		.INIT('h15)
	) name8874 (
		\u0_w_reg[3][2]/P0001 ,
		_w9297_,
		_w9369_,
		_w9407_
	);
	LUT3 #(
		.INIT('h10)
	) name8875 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9408_
	);
	LUT2 #(
		.INIT('h4)
	) name8876 (
		_w9365_,
		_w9408_,
		_w9409_
	);
	LUT3 #(
		.INIT('h8a)
	) name8877 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w9386_,
		_w9410_
	);
	LUT4 #(
		.INIT('h0080)
	) name8878 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9411_
	);
	LUT4 #(
		.INIT('h0020)
	) name8879 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9412_
	);
	LUT4 #(
		.INIT('h0007)
	) name8880 (
		_w9256_,
		_w9336_,
		_w9411_,
		_w9412_,
		_w9413_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name8881 (
		_w9407_,
		_w9409_,
		_w9410_,
		_w9413_,
		_w9414_
	);
	LUT4 #(
		.INIT('h2300)
	) name8882 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		_w9415_
	);
	LUT2 #(
		.INIT('h8)
	) name8883 (
		_w9314_,
		_w9415_,
		_w9416_
	);
	LUT3 #(
		.INIT('h15)
	) name8884 (
		\u0_w_reg[3][1]/P0001 ,
		_w9261_,
		_w9281_,
		_w9417_
	);
	LUT2 #(
		.INIT('h4)
	) name8885 (
		_w9416_,
		_w9417_,
		_w9418_
	);
	LUT4 #(
		.INIT('h555e)
	) name8886 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9419_
	);
	LUT4 #(
		.INIT('haf8c)
	) name8887 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		_w9255_,
		_w9419_,
		_w9420_
	);
	LUT2 #(
		.INIT('h1)
	) name8888 (
		\u0_w_reg[3][2]/P0001 ,
		_w9420_,
		_w9421_
	);
	LUT4 #(
		.INIT('h0020)
	) name8889 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9422_
	);
	LUT3 #(
		.INIT('ha8)
	) name8890 (
		\u0_w_reg[3][4]/P0001 ,
		_w9300_,
		_w9422_,
		_w9423_
	);
	LUT3 #(
		.INIT('h02)
	) name8891 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9424_
	);
	LUT2 #(
		.INIT('h8)
	) name8892 (
		_w9289_,
		_w9424_,
		_w9425_
	);
	LUT3 #(
		.INIT('h02)
	) name8893 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		_w9426_
	);
	LUT3 #(
		.INIT('h2a)
	) name8894 (
		\u0_w_reg[3][1]/P0001 ,
		_w9329_,
		_w9426_,
		_w9427_
	);
	LUT3 #(
		.INIT('h10)
	) name8895 (
		_w9423_,
		_w9425_,
		_w9427_,
		_w9428_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name8896 (
		_w9414_,
		_w9418_,
		_w9421_,
		_w9428_,
		_w9429_
	);
	LUT4 #(
		.INIT('h000e)
	) name8897 (
		_w9385_,
		_w9405_,
		_w9406_,
		_w9429_,
		_w9430_
	);
	LUT2 #(
		.INIT('h9)
	) name8898 (
		\u0_w_reg[1][12]/P0001 ,
		\u0_w_reg[2][12]/P0001 ,
		_w9431_
	);
	LUT3 #(
		.INIT('h69)
	) name8899 (
		\u0_w_reg[0][12]/P0001 ,
		_w9430_,
		_w9431_,
		_w9432_
	);
	LUT4 #(
		.INIT('h1441)
	) name8900 (
		ld_pad,
		\u0_w_reg[0][12]/P0001 ,
		_w9430_,
		_w9431_,
		_w9433_
	);
	LUT2 #(
		.INIT('h1)
	) name8901 (
		_w9361_,
		_w9433_,
		_w9434_
	);
	LUT3 #(
		.INIT('h54)
	) name8902 (
		\u0_w_reg[3][19]/P0001 ,
		_w8739_,
		_w8682_,
		_w9435_
	);
	LUT3 #(
		.INIT('h80)
	) name8903 (
		\u0_w_reg[3][20]/P0001 ,
		_w8659_,
		_w8772_,
		_w9436_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name8904 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9437_
	);
	LUT2 #(
		.INIT('h2)
	) name8905 (
		\u0_w_reg[3][18]/P0001 ,
		_w9437_,
		_w9438_
	);
	LUT3 #(
		.INIT('h01)
	) name8906 (
		\u0_w_reg[3][17]/P0001 ,
		_w8718_,
		_w8760_,
		_w9439_
	);
	LUT4 #(
		.INIT('h0100)
	) name8907 (
		_w9438_,
		_w9435_,
		_w9436_,
		_w9439_,
		_w9440_
	);
	LUT3 #(
		.INIT('h40)
	) name8908 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w9441_
	);
	LUT4 #(
		.INIT('h0002)
	) name8909 (
		\u0_w_reg[3][17]/P0001 ,
		_w8698_,
		_w9144_,
		_w9441_,
		_w9442_
	);
	LUT4 #(
		.INIT('h2000)
	) name8910 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9443_
	);
	LUT3 #(
		.INIT('h07)
	) name8911 (
		_w8721_,
		_w8723_,
		_w9443_,
		_w9444_
	);
	LUT4 #(
		.INIT('h002a)
	) name8912 (
		\u0_w_reg[3][18]/P0001 ,
		_w8707_,
		_w8720_,
		_w9159_,
		_w9445_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name8913 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9446_
	);
	LUT2 #(
		.INIT('h2)
	) name8914 (
		\u0_w_reg[3][19]/P0001 ,
		_w9446_,
		_w9447_
	);
	LUT4 #(
		.INIT('h0040)
	) name8915 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9448_
	);
	LUT3 #(
		.INIT('h01)
	) name8916 (
		\u0_w_reg[3][18]/P0001 ,
		_w8747_,
		_w9448_,
		_w9449_
	);
	LUT4 #(
		.INIT('h7077)
	) name8917 (
		_w9444_,
		_w9445_,
		_w9447_,
		_w9449_,
		_w9450_
	);
	LUT4 #(
		.INIT('h0040)
	) name8918 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9451_
	);
	LUT3 #(
		.INIT('h07)
	) name8919 (
		_w8659_,
		_w8760_,
		_w9451_,
		_w9452_
	);
	LUT4 #(
		.INIT('h5400)
	) name8920 (
		_w9450_,
		_w9440_,
		_w9442_,
		_w9452_,
		_w9453_
	);
	LUT3 #(
		.INIT('h80)
	) name8921 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w9454_
	);
	LUT3 #(
		.INIT('ha8)
	) name8922 (
		\u0_w_reg[3][23]/P0001 ,
		_w8772_,
		_w9454_,
		_w9455_
	);
	LUT4 #(
		.INIT('h0080)
	) name8923 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9456_
	);
	LUT4 #(
		.INIT('h0007)
	) name8924 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9457_
	);
	LUT4 #(
		.INIT('h002a)
	) name8925 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w9456_,
		_w9457_,
		_w9458_
	);
	LUT4 #(
		.INIT('hbfef)
	) name8926 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9459_
	);
	LUT2 #(
		.INIT('h1)
	) name8927 (
		\u0_w_reg[3][19]/P0001 ,
		_w9459_,
		_w9460_
	);
	LUT4 #(
		.INIT('h4c00)
	) name8928 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9461_
	);
	LUT4 #(
		.INIT('h0145)
	) name8929 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		_w8727_,
		_w9461_,
		_w9462_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name8930 (
		_w9455_,
		_w9458_,
		_w9460_,
		_w9462_,
		_w9463_
	);
	LUT3 #(
		.INIT('h02)
	) name8931 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9464_
	);
	LUT3 #(
		.INIT('hb9)
	) name8932 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9465_
	);
	LUT2 #(
		.INIT('h2)
	) name8933 (
		_w9157_,
		_w9465_,
		_w9466_
	);
	LUT4 #(
		.INIT('h0001)
	) name8934 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w9467_
	);
	LUT4 #(
		.INIT('h0007)
	) name8935 (
		_w8707_,
		_w8720_,
		_w9120_,
		_w9467_,
		_w9468_
	);
	LUT3 #(
		.INIT('h32)
	) name8936 (
		\u0_w_reg[3][18]/P0001 ,
		_w9466_,
		_w9468_,
		_w9469_
	);
	LUT2 #(
		.INIT('h4)
	) name8937 (
		_w9463_,
		_w9469_,
		_w9470_
	);
	LUT4 #(
		.INIT('h4000)
	) name8938 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9471_
	);
	LUT4 #(
		.INIT('haa80)
	) name8939 (
		\u0_w_reg[3][22]/P0001 ,
		_w8743_,
		_w8721_,
		_w9471_,
		_w9472_
	);
	LUT3 #(
		.INIT('h20)
	) name8940 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w9473_
	);
	LUT4 #(
		.INIT('hffde)
	) name8941 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w9474_
	);
	LUT4 #(
		.INIT('h4055)
	) name8942 (
		\u0_w_reg[3][23]/P0001 ,
		_w8732_,
		_w9473_,
		_w9474_,
		_w9475_
	);
	LUT2 #(
		.INIT('h8)
	) name8943 (
		_w8730_,
		_w8689_,
		_w9476_
	);
	LUT3 #(
		.INIT('h8a)
	) name8944 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		_w8734_,
		_w9477_
	);
	LUT3 #(
		.INIT('h10)
	) name8945 (
		_w9475_,
		_w9476_,
		_w9477_,
		_w9478_
	);
	LUT4 #(
		.INIT('h0004)
	) name8946 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9479_
	);
	LUT4 #(
		.INIT('hff4b)
	) name8947 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9480_
	);
	LUT2 #(
		.INIT('h2)
	) name8948 (
		_w8764_,
		_w9480_,
		_w9481_
	);
	LUT3 #(
		.INIT('h67)
	) name8949 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9482_
	);
	LUT2 #(
		.INIT('h2)
	) name8950 (
		_w8743_,
		_w9482_,
		_w9483_
	);
	LUT4 #(
		.INIT('h0040)
	) name8951 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9484_
	);
	LUT2 #(
		.INIT('h8)
	) name8952 (
		_w8729_,
		_w9484_,
		_w9485_
	);
	LUT3 #(
		.INIT('h15)
	) name8953 (
		\u0_w_reg[3][17]/P0001 ,
		_w8689_,
		_w8770_,
		_w9486_
	);
	LUT4 #(
		.INIT('h0100)
	) name8954 (
		_w9483_,
		_w9485_,
		_w9481_,
		_w9486_,
		_w9487_
	);
	LUT3 #(
		.INIT('h54)
	) name8955 (
		_w9472_,
		_w9478_,
		_w9487_,
		_w9488_
	);
	LUT4 #(
		.INIT('he400)
	) name8956 (
		\u0_w_reg[3][16]/P0001 ,
		_w9470_,
		_w9453_,
		_w9488_,
		_w9489_
	);
	LUT2 #(
		.INIT('h9)
	) name8957 (
		\u0_r0_out_reg[24]/P0001 ,
		\u0_w_reg[0][24]/P0001 ,
		_w9490_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name8958 (
		\key[120]_pad ,
		ld_pad,
		_w9489_,
		_w9490_,
		_w9491_
	);
	LUT3 #(
		.INIT('h0e)
	) name8959 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		_w9492_
	);
	LUT4 #(
		.INIT('h5054)
	) name8960 (
		\u0_w_reg[3][19]/P0001 ,
		_w8680_,
		_w8739_,
		_w9492_,
		_w9493_
	);
	LUT4 #(
		.INIT('h0020)
	) name8961 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9494_
	);
	LUT4 #(
		.INIT('h0200)
	) name8962 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9495_
	);
	LUT4 #(
		.INIT('h2000)
	) name8963 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9496_
	);
	LUT4 #(
		.INIT('h0001)
	) name8964 (
		\u0_w_reg[3][17]/P0001 ,
		_w9494_,
		_w9495_,
		_w9496_,
		_w9497_
	);
	LUT3 #(
		.INIT('h0b)
	) name8965 (
		\u0_w_reg[3][18]/P0001 ,
		_w8740_,
		_w9456_,
		_w9498_
	);
	LUT4 #(
		.INIT('h0002)
	) name8966 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9499_
	);
	LUT4 #(
		.INIT('h002a)
	) name8967 (
		\u0_w_reg[3][17]/P0001 ,
		_w8729_,
		_w9484_,
		_w9499_,
		_w9500_
	);
	LUT4 #(
		.INIT('h00bf)
	) name8968 (
		_w9493_,
		_w9497_,
		_w9498_,
		_w9500_,
		_w9501_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name8969 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9502_
	);
	LUT2 #(
		.INIT('h2)
	) name8970 (
		_w8689_,
		_w9502_,
		_w9503_
	);
	LUT2 #(
		.INIT('h2)
	) name8971 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		_w9504_
	);
	LUT4 #(
		.INIT('hbbf3)
	) name8972 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w9505_
	);
	LUT2 #(
		.INIT('h2)
	) name8973 (
		_w9504_,
		_w9505_,
		_w9506_
	);
	LUT3 #(
		.INIT('hed)
	) name8974 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9507_
	);
	LUT2 #(
		.INIT('h2)
	) name8975 (
		_w8657_,
		_w9507_,
		_w9508_
	);
	LUT3 #(
		.INIT('h2a)
	) name8976 (
		\u0_w_reg[3][16]/P0001 ,
		_w8732_,
		_w8733_,
		_w9509_
	);
	LUT4 #(
		.INIT('h0100)
	) name8977 (
		_w9503_,
		_w9508_,
		_w9506_,
		_w9509_,
		_w9510_
	);
	LUT4 #(
		.INIT('h0040)
	) name8978 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9511_
	);
	LUT3 #(
		.INIT('h01)
	) name8979 (
		\u0_w_reg[3][17]/P0001 ,
		_w8734_,
		_w9511_,
		_w9512_
	);
	LUT4 #(
		.INIT('h0800)
	) name8980 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9513_
	);
	LUT2 #(
		.INIT('h2)
	) name8981 (
		\u0_w_reg[3][17]/P0001 ,
		_w9513_,
		_w9514_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name8982 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9515_
	);
	LUT4 #(
		.INIT('hffda)
	) name8983 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9516_
	);
	LUT4 #(
		.INIT('hfe54)
	) name8984 (
		\u0_w_reg[3][18]/P0001 ,
		_w8721_,
		_w9515_,
		_w9516_,
		_w9517_
	);
	LUT3 #(
		.INIT('h15)
	) name8985 (
		_w9512_,
		_w9514_,
		_w9517_,
		_w9518_
	);
	LUT3 #(
		.INIT('h80)
	) name8986 (
		\u0_w_reg[3][22]/P0001 ,
		_w8684_,
		_w8689_,
		_w9519_
	);
	LUT2 #(
		.INIT('h1)
	) name8987 (
		\u0_w_reg[3][16]/P0001 ,
		_w8708_,
		_w9520_
	);
	LUT3 #(
		.INIT('h10)
	) name8988 (
		_w8769_,
		_w9519_,
		_w9520_,
		_w9521_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name8989 (
		_w9501_,
		_w9510_,
		_w9518_,
		_w9521_,
		_w9522_
	);
	LUT4 #(
		.INIT('h0007)
	) name8990 (
		_w8746_,
		_w8664_,
		_w9135_,
		_w9479_,
		_w9523_
	);
	LUT2 #(
		.INIT('h1)
	) name8991 (
		\u0_w_reg[3][18]/P0001 ,
		_w9523_,
		_w9524_
	);
	LUT4 #(
		.INIT('hbcfc)
	) name8992 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9525_
	);
	LUT2 #(
		.INIT('h2)
	) name8993 (
		_w8689_,
		_w9525_,
		_w9526_
	);
	LUT2 #(
		.INIT('h8)
	) name8994 (
		\u0_w_reg[3][18]/P0001 ,
		_w8734_,
		_w9527_
	);
	LUT4 #(
		.INIT('h000b)
	) name8995 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w9528_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name8996 (
		_w8692_,
		_w8764_,
		_w9464_,
		_w9528_,
		_w9529_
	);
	LUT3 #(
		.INIT('h10)
	) name8997 (
		_w9526_,
		_w9527_,
		_w9529_,
		_w9530_
	);
	LUT3 #(
		.INIT('h45)
	) name8998 (
		\u0_w_reg[3][17]/P0001 ,
		_w9524_,
		_w9530_,
		_w9531_
	);
	LUT3 #(
		.INIT('h13)
	) name8999 (
		\u0_w_reg[3][20]/P0001 ,
		_w8704_,
		_w9120_,
		_w9532_
	);
	LUT3 #(
		.INIT('h10)
	) name9000 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9533_
	);
	LUT4 #(
		.INIT('h0400)
	) name9001 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9534_
	);
	LUT4 #(
		.INIT('h0013)
	) name9002 (
		\u0_w_reg[3][20]/P0001 ,
		_w8704_,
		_w9120_,
		_w9534_,
		_w9535_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name9003 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		_w8677_,
		_w9535_,
		_w9536_
	);
	LUT2 #(
		.INIT('h2)
	) name9004 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9537_
	);
	LUT3 #(
		.INIT('h80)
	) name9005 (
		_w8697_,
		_w9157_,
		_w9537_,
		_w9538_
	);
	LUT3 #(
		.INIT('had)
	) name9006 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9539_
	);
	LUT4 #(
		.INIT('he2ee)
	) name9007 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w9540_
	);
	LUT2 #(
		.INIT('h8)
	) name9008 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		_w9541_
	);
	LUT3 #(
		.INIT('h80)
	) name9009 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9542_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name9010 (
		_w8743_,
		_w9539_,
		_w9540_,
		_w9542_,
		_w9543_
	);
	LUT3 #(
		.INIT('h10)
	) name9011 (
		_w9160_,
		_w9538_,
		_w9543_,
		_w9544_
	);
	LUT2 #(
		.INIT('h4)
	) name9012 (
		_w9536_,
		_w9544_,
		_w9545_
	);
	LUT4 #(
		.INIT('h5655)
	) name9013 (
		\u0_w_reg[0][26]/P0001 ,
		_w9531_,
		_w9522_,
		_w9545_,
		_w9546_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name9014 (
		\key[122]_pad ,
		ld_pad,
		\u0_r0_out_reg[26]/P0001 ,
		_w9546_,
		_w9547_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name9015 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9548_
	);
	LUT4 #(
		.INIT('h20aa)
	) name9016 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w8677_,
		_w9548_,
		_w9549_
	);
	LUT2 #(
		.INIT('h4)
	) name9017 (
		_w8703_,
		_w8772_,
		_w9550_
	);
	LUT4 #(
		.INIT('haaa2)
	) name9018 (
		\u0_w_reg[3][17]/P0001 ,
		_w9444_,
		_w9550_,
		_w9549_,
		_w9551_
	);
	LUT3 #(
		.INIT('ha8)
	) name9019 (
		\u0_w_reg[3][18]/P0001 ,
		_w8752_,
		_w9134_,
		_w9552_
	);
	LUT3 #(
		.INIT('h15)
	) name9020 (
		_w8708_,
		_w8764_,
		_w9464_,
		_w9553_
	);
	LUT4 #(
		.INIT('h5455)
	) name9021 (
		\u0_w_reg[3][17]/P0001 ,
		_w8706_,
		_w9552_,
		_w9553_,
		_w9554_
	);
	LUT3 #(
		.INIT('h54)
	) name9022 (
		\u0_w_reg[3][18]/P0001 ,
		_w8655_,
		_w9484_,
		_w9555_
	);
	LUT2 #(
		.INIT('h1)
	) name9023 (
		_w8709_,
		_w9119_,
		_w9556_
	);
	LUT4 #(
		.INIT('h0d05)
	) name9024 (
		\u0_w_reg[3][18]/P0001 ,
		_w9109_,
		_w9555_,
		_w9556_,
		_w9557_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9025 (
		\u0_w_reg[3][16]/P0001 ,
		_w9551_,
		_w9554_,
		_w9557_,
		_w9558_
	);
	LUT3 #(
		.INIT('h13)
	) name9026 (
		_w8721_,
		_w9145_,
		_w9111_,
		_w9559_
	);
	LUT4 #(
		.INIT('h0004)
	) name9027 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w9560_
	);
	LUT3 #(
		.INIT('h0b)
	) name9028 (
		_w8680_,
		_w8760_,
		_w9560_,
		_w9561_
	);
	LUT3 #(
		.INIT('h15)
	) name9029 (
		\u0_w_reg[3][18]/P0001 ,
		_w9559_,
		_w9561_,
		_w9562_
	);
	LUT3 #(
		.INIT('h9d)
	) name9030 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w9563_
	);
	LUT2 #(
		.INIT('h2)
	) name9031 (
		_w8683_,
		_w9563_,
		_w9564_
	);
	LUT3 #(
		.INIT('h01)
	) name9032 (
		\u0_w_reg[3][17]/P0001 ,
		_w9471_,
		_w9484_,
		_w9565_
	);
	LUT4 #(
		.INIT('h0100)
	) name9033 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9566_
	);
	LUT3 #(
		.INIT('h07)
	) name9034 (
		_w8689_,
		_w9464_,
		_w9566_,
		_w9567_
	);
	LUT3 #(
		.INIT('h40)
	) name9035 (
		_w9564_,
		_w9565_,
		_w9567_,
		_w9568_
	);
	LUT2 #(
		.INIT('h2)
	) name9036 (
		_w8732_,
		_w8695_,
		_w9569_
	);
	LUT2 #(
		.INIT('h4)
	) name9037 (
		\u0_w_reg[3][18]/P0001 ,
		_w8709_,
		_w9570_
	);
	LUT3 #(
		.INIT('h2a)
	) name9038 (
		\u0_w_reg[3][17]/P0001 ,
		_w8746_,
		_w8664_,
		_w9571_
	);
	LUT3 #(
		.INIT('h10)
	) name9039 (
		_w9569_,
		_w9570_,
		_w9571_,
		_w9572_
	);
	LUT4 #(
		.INIT('h4445)
	) name9040 (
		\u0_w_reg[3][16]/P0001 ,
		_w9562_,
		_w9568_,
		_w9572_,
		_w9573_
	);
	LUT3 #(
		.INIT('h20)
	) name9041 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9574_
	);
	LUT4 #(
		.INIT('h0103)
	) name9042 (
		_w8714_,
		_w8751_,
		_w9165_,
		_w9574_,
		_w9575_
	);
	LUT4 #(
		.INIT('h5540)
	) name9043 (
		\u0_w_reg[3][16]/P0001 ,
		_w8654_,
		_w8676_,
		_w9467_,
		_w9576_
	);
	LUT4 #(
		.INIT('h0301)
	) name9044 (
		\u0_w_reg[3][17]/P0001 ,
		_w9170_,
		_w9576_,
		_w9575_,
		_w9577_
	);
	LUT2 #(
		.INIT('h2)
	) name9045 (
		\u0_w_reg[3][18]/P0001 ,
		_w9577_,
		_w9578_
	);
	LUT2 #(
		.INIT('h8)
	) name9046 (
		_w8729_,
		_w9574_,
		_w9579_
	);
	LUT3 #(
		.INIT('h1b)
	) name9047 (
		\u0_w_reg[3][18]/P0001 ,
		_w8698_,
		_w9114_,
		_w9580_
	);
	LUT3 #(
		.INIT('h23)
	) name9048 (
		\u0_w_reg[3][18]/P0001 ,
		_w8663_,
		_w8708_,
		_w9581_
	);
	LUT3 #(
		.INIT('h13)
	) name9049 (
		_w8680_,
		_w9135_,
		_w9157_,
		_w9582_
	);
	LUT4 #(
		.INIT('h4000)
	) name9050 (
		_w9579_,
		_w9581_,
		_w9582_,
		_w9580_,
		_w9583_
	);
	LUT3 #(
		.INIT('h54)
	) name9051 (
		\u0_w_reg[3][19]/P0001 ,
		_w8682_,
		_w8709_,
		_w9584_
	);
	LUT4 #(
		.INIT('h0200)
	) name9052 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8767_,
		_w9585_
	);
	LUT3 #(
		.INIT('h01)
	) name9053 (
		_w9123_,
		_w9585_,
		_w9584_,
		_w9586_
	);
	LUT3 #(
		.INIT('he0)
	) name9054 (
		\u0_w_reg[3][17]/P0001 ,
		_w9583_,
		_w9586_,
		_w9587_
	);
	LUT4 #(
		.INIT('h0100)
	) name9055 (
		_w9558_,
		_w9573_,
		_w9578_,
		_w9587_,
		_w9588_
	);
	LUT4 #(
		.INIT('h1441)
	) name9056 (
		ld_pad,
		\u0_r0_out_reg[30]/P0001 ,
		\u0_w_reg[0][30]/P0001 ,
		_w9588_,
		_w9589_
	);
	LUT2 #(
		.INIT('h8)
	) name9057 (
		\key[126]_pad ,
		ld_pad,
		_w9590_
	);
	LUT2 #(
		.INIT('he)
	) name9058 (
		_w9589_,
		_w9590_,
		_w9591_
	);
	LUT3 #(
		.INIT('h40)
	) name9059 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9592_
	);
	LUT4 #(
		.INIT('ha7f7)
	) name9060 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9593_
	);
	LUT2 #(
		.INIT('h2)
	) name9061 (
		_w8732_,
		_w9593_,
		_w9594_
	);
	LUT3 #(
		.INIT('h07)
	) name9062 (
		\u0_w_reg[3][18]/P0001 ,
		_w8671_,
		_w9448_,
		_w9595_
	);
	LUT4 #(
		.INIT('h15bf)
	) name9063 (
		\u0_w_reg[3][20]/P0001 ,
		_w8697_,
		_w8689_,
		_w9146_,
		_w9596_
	);
	LUT3 #(
		.INIT('h40)
	) name9064 (
		_w9594_,
		_w9595_,
		_w9596_,
		_w9597_
	);
	LUT4 #(
		.INIT('h7d5d)
	) name9065 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9598_
	);
	LUT2 #(
		.INIT('h1)
	) name9066 (
		\u0_w_reg[3][18]/P0001 ,
		_w9598_,
		_w9599_
	);
	LUT4 #(
		.INIT('h3100)
	) name9067 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w9600_
	);
	LUT3 #(
		.INIT('h54)
	) name9068 (
		\u0_w_reg[3][23]/P0001 ,
		_w9441_,
		_w9600_,
		_w9601_
	);
	LUT3 #(
		.INIT('h07)
	) name9069 (
		\u0_w_reg[3][23]/P0001 ,
		_w8744_,
		_w8767_,
		_w9602_
	);
	LUT3 #(
		.INIT('h10)
	) name9070 (
		_w9601_,
		_w9599_,
		_w9602_,
		_w9603_
	);
	LUT4 #(
		.INIT('h3fbb)
	) name9071 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9604_
	);
	LUT2 #(
		.INIT('h2)
	) name9072 (
		_w8764_,
		_w9604_,
		_w9605_
	);
	LUT3 #(
		.INIT('h10)
	) name9073 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9606_
	);
	LUT4 #(
		.INIT('h0111)
	) name9074 (
		\u0_w_reg[3][17]/P0001 ,
		_w8734_,
		_w8729_,
		_w9606_,
		_w9607_
	);
	LUT2 #(
		.INIT('h4)
	) name9075 (
		_w9605_,
		_w9607_,
		_w9608_
	);
	LUT4 #(
		.INIT('hd500)
	) name9076 (
		\u0_w_reg[3][16]/P0001 ,
		_w9597_,
		_w9603_,
		_w9608_,
		_w9609_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name9077 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9610_
	);
	LUT3 #(
		.INIT('h51)
	) name9078 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w9610_,
		_w9611_
	);
	LUT3 #(
		.INIT('had)
	) name9079 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w9612_
	);
	LUT4 #(
		.INIT('hadfb)
	) name9080 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9613_
	);
	LUT2 #(
		.INIT('h1)
	) name9081 (
		\u0_w_reg[3][19]/P0001 ,
		_w9613_,
		_w9614_
	);
	LUT3 #(
		.INIT('h02)
	) name9082 (
		\u0_w_reg[3][18]/P0001 ,
		_w8737_,
		_w8704_,
		_w9615_
	);
	LUT3 #(
		.INIT('h45)
	) name9083 (
		_w9611_,
		_w9614_,
		_w9615_,
		_w9616_
	);
	LUT3 #(
		.INIT('hf6)
	) name9084 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9617_
	);
	LUT3 #(
		.INIT('h2a)
	) name9085 (
		\u0_w_reg[3][18]/P0001 ,
		_w9612_,
		_w9617_,
		_w9618_
	);
	LUT4 #(
		.INIT('h153f)
	) name9086 (
		_w8697_,
		_w8659_,
		_w8772_,
		_w9134_,
		_w9619_
	);
	LUT2 #(
		.INIT('h4)
	) name9087 (
		_w9618_,
		_w9619_,
		_w9620_
	);
	LUT4 #(
		.INIT('hc444)
	) name9088 (
		\u0_w_reg[3][16]/P0001 ,
		\u0_w_reg[3][17]/P0001 ,
		_w9597_,
		_w9620_,
		_w9621_
	);
	LUT3 #(
		.INIT('h45)
	) name9089 (
		_w9609_,
		_w9616_,
		_w9621_,
		_w9622_
	);
	LUT4 #(
		.INIT('h0020)
	) name9090 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9623_
	);
	LUT3 #(
		.INIT('h54)
	) name9091 (
		\u0_w_reg[3][18]/P0001 ,
		_w8723_,
		_w9623_,
		_w9624_
	);
	LUT4 #(
		.INIT('h153f)
	) name9092 (
		_w8732_,
		_w8654_,
		_w8676_,
		_w9473_,
		_w9625_
	);
	LUT3 #(
		.INIT('h20)
	) name9093 (
		_w9514_,
		_w9624_,
		_w9625_,
		_w9626_
	);
	LUT2 #(
		.INIT('h1)
	) name9094 (
		\u0_w_reg[3][17]/P0001 ,
		_w8682_,
		_w9627_
	);
	LUT3 #(
		.INIT('h07)
	) name9095 (
		_w8684_,
		_w8689_,
		_w9443_,
		_w9628_
	);
	LUT2 #(
		.INIT('h8)
	) name9096 (
		_w9627_,
		_w9628_,
		_w9629_
	);
	LUT4 #(
		.INIT('h153f)
	) name9097 (
		\u0_w_reg[3][20]/P0001 ,
		_w8680_,
		_w8760_,
		_w9120_,
		_w9630_
	);
	LUT2 #(
		.INIT('h2)
	) name9098 (
		\u0_w_reg[3][18]/P0001 ,
		_w9630_,
		_w9631_
	);
	LUT3 #(
		.INIT('h10)
	) name9099 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w9632_
	);
	LUT3 #(
		.INIT('h54)
	) name9100 (
		\u0_w_reg[3][18]/P0001 ,
		_w9165_,
		_w9632_,
		_w9633_
	);
	LUT4 #(
		.INIT('h0001)
	) name9101 (
		_w8763_,
		_w8771_,
		_w9605_,
		_w9633_,
		_w9634_
	);
	LUT4 #(
		.INIT('h0e00)
	) name9102 (
		_w9626_,
		_w9629_,
		_w9631_,
		_w9634_,
		_w9635_
	);
	LUT4 #(
		.INIT('h8caf)
	) name9103 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8727_,
		_w8663_,
		_w9636_
	);
	LUT4 #(
		.INIT('h4000)
	) name9104 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w9637_
	);
	LUT4 #(
		.INIT('h0013)
	) name9105 (
		_w8697_,
		_w8666_,
		_w9134_,
		_w9637_,
		_w9638_
	);
	LUT4 #(
		.INIT('hfcb8)
	) name9106 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		_w9636_,
		_w9638_,
		_w9639_
	);
	LUT3 #(
		.INIT('he0)
	) name9107 (
		\u0_w_reg[3][16]/P0001 ,
		_w9635_,
		_w9639_,
		_w9640_
	);
	LUT3 #(
		.INIT('h65)
	) name9108 (
		\u0_w_reg[0][31]/P0001 ,
		_w9622_,
		_w9640_,
		_w9641_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name9109 (
		\key[127]_pad ,
		ld_pad,
		\u0_r0_out_reg[31]/P0001 ,
		_w9641_,
		_w9642_
	);
	LUT2 #(
		.INIT('h9)
	) name9110 (
		\u0_r0_out_reg[26]/P0001 ,
		\u0_w_reg[1][26]/P0001 ,
		_w9643_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9111 (
		\key[90]_pad ,
		ld_pad,
		_w9546_,
		_w9643_,
		_w9644_
	);
	LUT2 #(
		.INIT('h9)
	) name9112 (
		\u0_w_reg[0][30]/P0001 ,
		\u0_w_reg[1][30]/P0001 ,
		_w9645_
	);
	LUT4 #(
		.INIT('h4114)
	) name9113 (
		ld_pad,
		\u0_r0_out_reg[30]/P0001 ,
		_w9588_,
		_w9645_,
		_w9646_
	);
	LUT2 #(
		.INIT('h8)
	) name9114 (
		\key[94]_pad ,
		ld_pad,
		_w9647_
	);
	LUT2 #(
		.INIT('he)
	) name9115 (
		_w9646_,
		_w9647_,
		_w9648_
	);
	LUT2 #(
		.INIT('h9)
	) name9116 (
		\u0_r0_out_reg[31]/P0001 ,
		\u0_w_reg[1][31]/P0001 ,
		_w9649_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9117 (
		\key[95]_pad ,
		ld_pad,
		_w9641_,
		_w9649_,
		_w9650_
	);
	LUT2 #(
		.INIT('h9)
	) name9118 (
		\u0_w_reg[1][24]/P0002 ,
		\u0_w_reg[2][24]/P0001 ,
		_w9651_
	);
	LUT4 #(
		.INIT('h9669)
	) name9119 (
		\u0_r0_out_reg[24]/P0001 ,
		\u0_w_reg[0][24]/P0001 ,
		\u0_w_reg[1][24]/P0002 ,
		\u0_w_reg[2][24]/P0001 ,
		_w9652_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name9120 (
		\key[56]_pad ,
		ld_pad,
		_w9489_,
		_w9652_,
		_w9653_
	);
	LUT3 #(
		.INIT('h69)
	) name9121 (
		\u0_r0_out_reg[26]/P0001 ,
		\u0_w_reg[1][26]/P0001 ,
		\u0_w_reg[2][26]/P0001 ,
		_w9654_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9122 (
		\key[58]_pad ,
		ld_pad,
		_w9546_,
		_w9654_,
		_w9655_
	);
	LUT2 #(
		.INIT('h4)
	) name9123 (
		\key[62]_pad ,
		ld_pad,
		_w9656_
	);
	LUT3 #(
		.INIT('h69)
	) name9124 (
		\u0_w_reg[0][30]/P0001 ,
		\u0_w_reg[1][30]/P0001 ,
		\u0_w_reg[2][30]/P0001 ,
		_w9657_
	);
	LUT3 #(
		.INIT('h69)
	) name9125 (
		\u0_r0_out_reg[30]/P0001 ,
		_w9588_,
		_w9657_,
		_w9658_
	);
	LUT4 #(
		.INIT('h1441)
	) name9126 (
		ld_pad,
		\u0_r0_out_reg[30]/P0001 ,
		_w9588_,
		_w9657_,
		_w9659_
	);
	LUT2 #(
		.INIT('h1)
	) name9127 (
		_w9656_,
		_w9659_,
		_w9660_
	);
	LUT3 #(
		.INIT('h69)
	) name9128 (
		\u0_r0_out_reg[31]/P0001 ,
		\u0_w_reg[1][31]/P0001 ,
		\u0_w_reg[2][31]/P0001 ,
		_w9661_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9129 (
		\u0_w_reg[0][31]/P0001 ,
		_w9622_,
		_w9640_,
		_w9661_,
		_w9662_
	);
	LUT3 #(
		.INIT('h8b)
	) name9130 (
		\key[63]_pad ,
		ld_pad,
		_w9662_,
		_w9663_
	);
	LUT3 #(
		.INIT('h96)
	) name9131 (
		\u0_w_reg[3][24]/P0001 ,
		_w9489_,
		_w9490_,
		_w9664_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9132 (
		\key[24]_pad ,
		ld_pad,
		_w9651_,
		_w9664_,
		_w9665_
	);
	LUT4 #(
		.INIT('h1441)
	) name9133 (
		ld_pad,
		\u0_w_reg[3][26]/P0001 ,
		_w9546_,
		_w9654_,
		_w9666_
	);
	LUT2 #(
		.INIT('h8)
	) name9134 (
		\key[26]_pad ,
		ld_pad,
		_w9667_
	);
	LUT2 #(
		.INIT('he)
	) name9135 (
		_w9666_,
		_w9667_,
		_w9668_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9136 (
		\key[30]_pad ,
		ld_pad,
		\u0_w_reg[3][30]/P0001 ,
		_w9658_,
		_w9669_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9137 (
		\key[31]_pad ,
		ld_pad,
		\u0_w_reg[3][31]/P0001 ,
		_w9662_,
		_w9670_
	);
	LUT3 #(
		.INIT('hb8)
	) name9138 (
		\key[117]_pad ,
		ld_pad,
		_w8900_,
		_w9671_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name9139 (
		\key[85]_pad ,
		ld_pad,
		\u0_w_reg[1][21]/P0001 ,
		_w8900_,
		_w9672_
	);
	LUT4 #(
		.INIT('h1441)
	) name9140 (
		ld_pad,
		\u0_w_reg[3][21]/P0001 ,
		_w8900_,
		_w8901_,
		_w9673_
	);
	LUT2 #(
		.INIT('h8)
	) name9141 (
		\key[21]_pad ,
		ld_pad,
		_w9674_
	);
	LUT2 #(
		.INIT('he)
	) name9142 (
		_w9673_,
		_w9674_,
		_w9675_
	);
	LUT3 #(
		.INIT('h15)
	) name9143 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9676_
	);
	LUT3 #(
		.INIT('ha2)
	) name9144 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9677_
	);
	LUT3 #(
		.INIT('h02)
	) name9145 (
		_w9068_,
		_w9677_,
		_w9676_,
		_w9678_
	);
	LUT3 #(
		.INIT('h07)
	) name9146 (
		_w9006_,
		_w9007_,
		_w9212_,
		_w9679_
	);
	LUT3 #(
		.INIT('h08)
	) name9147 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9680_
	);
	LUT3 #(
		.INIT('h08)
	) name9148 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w9681_
	);
	LUT4 #(
		.INIT('h153f)
	) name9149 (
		_w9014_,
		_w9197_,
		_w9680_,
		_w9681_,
		_w9682_
	);
	LUT3 #(
		.INIT('h40)
	) name9150 (
		_w9678_,
		_w9679_,
		_w9682_,
		_w9683_
	);
	LUT4 #(
		.INIT('h82a2)
	) name9151 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9684_
	);
	LUT4 #(
		.INIT('hff2f)
	) name9152 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9685_
	);
	LUT3 #(
		.INIT('h45)
	) name9153 (
		\u0_w_reg[3][26]/P0001 ,
		_w9684_,
		_w9685_,
		_w9686_
	);
	LUT3 #(
		.INIT('h10)
	) name9154 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9687_
	);
	LUT4 #(
		.INIT('h0040)
	) name9155 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9688_
	);
	LUT4 #(
		.INIT('h0020)
	) name9156 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9689_
	);
	LUT4 #(
		.INIT('h0103)
	) name9157 (
		_w9068_,
		_w9688_,
		_w9689_,
		_w9687_,
		_w9690_
	);
	LUT2 #(
		.INIT('h4)
	) name9158 (
		_w9686_,
		_w9690_,
		_w9691_
	);
	LUT3 #(
		.INIT('h2a)
	) name9159 (
		\u0_w_reg[3][24]/P0001 ,
		_w9683_,
		_w9691_,
		_w9692_
	);
	LUT4 #(
		.INIT('h0010)
	) name9160 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9693_
	);
	LUT2 #(
		.INIT('h1)
	) name9161 (
		_w8985_,
		_w9693_,
		_w9694_
	);
	LUT2 #(
		.INIT('h4)
	) name9162 (
		\u0_w_reg[3][29]/P0001 ,
		_w9041_,
		_w9695_
	);
	LUT3 #(
		.INIT('h15)
	) name9163 (
		\u0_w_reg[3][26]/P0001 ,
		_w9000_,
		_w9001_,
		_w9696_
	);
	LUT3 #(
		.INIT('h20)
	) name9164 (
		_w9694_,
		_w9695_,
		_w9696_,
		_w9697_
	);
	LUT2 #(
		.INIT('h8)
	) name9165 (
		_w9189_,
		_w9194_,
		_w9698_
	);
	LUT3 #(
		.INIT('h02)
	) name9166 (
		\u0_w_reg[3][26]/P0001 ,
		_w9044_,
		_w9003_,
		_w9699_
	);
	LUT2 #(
		.INIT('h4)
	) name9167 (
		_w9698_,
		_w9699_,
		_w9700_
	);
	LUT4 #(
		.INIT('h0105)
	) name9168 (
		\u0_w_reg[3][25]/P0001 ,
		_w9090_,
		_w9196_,
		_w9687_,
		_w9701_
	);
	LUT3 #(
		.INIT('he0)
	) name9169 (
		_w9697_,
		_w9700_,
		_w9701_,
		_w9702_
	);
	LUT3 #(
		.INIT('had)
	) name9170 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9703_
	);
	LUT4 #(
		.INIT('hadfb)
	) name9171 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9704_
	);
	LUT2 #(
		.INIT('h1)
	) name9172 (
		\u0_w_reg[3][27]/P0001 ,
		_w9704_,
		_w9705_
	);
	LUT3 #(
		.INIT('h02)
	) name9173 (
		\u0_w_reg[3][26]/P0001 ,
		_w9043_,
		_w9028_,
		_w9706_
	);
	LUT2 #(
		.INIT('h4)
	) name9174 (
		_w9705_,
		_w9706_,
		_w9707_
	);
	LUT4 #(
		.INIT('hbfef)
	) name9175 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9708_
	);
	LUT3 #(
		.INIT('h02)
	) name9176 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9709_
	);
	LUT4 #(
		.INIT('hbfe3)
	) name9177 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9710_
	);
	LUT2 #(
		.INIT('h2)
	) name9178 (
		\u0_w_reg[3][27]/P0001 ,
		_w9710_,
		_w9711_
	);
	LUT4 #(
		.INIT('h0010)
	) name9179 (
		_w9075_,
		_w9695_,
		_w9696_,
		_w9711_,
		_w9712_
	);
	LUT2 #(
		.INIT('h1)
	) name9180 (
		_w9707_,
		_w9712_,
		_w9713_
	);
	LUT3 #(
		.INIT('hf6)
	) name9181 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9714_
	);
	LUT3 #(
		.INIT('h2a)
	) name9182 (
		\u0_w_reg[3][26]/P0001 ,
		_w9703_,
		_w9714_,
		_w9715_
	);
	LUT4 #(
		.INIT('h0100)
	) name9183 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9716_
	);
	LUT4 #(
		.INIT('h4c7f)
	) name9184 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9189_,
		_w9716_,
		_w9717_
	);
	LUT2 #(
		.INIT('h4)
	) name9185 (
		_w9715_,
		_w9717_,
		_w9718_
	);
	LUT4 #(
		.INIT('hc444)
	) name9186 (
		\u0_w_reg[3][24]/P0001 ,
		\u0_w_reg[3][25]/P0001 ,
		_w9683_,
		_w9718_,
		_w9719_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name9187 (
		_w9692_,
		_w9702_,
		_w9713_,
		_w9719_,
		_w9720_
	);
	LUT3 #(
		.INIT('h45)
	) name9188 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9084_,
		_w9721_
	);
	LUT4 #(
		.INIT('h0002)
	) name9189 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9722_
	);
	LUT3 #(
		.INIT('h10)
	) name9190 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9723_
	);
	LUT4 #(
		.INIT('h0001)
	) name9191 (
		_w8985_,
		_w9693_,
		_w9722_,
		_w9723_,
		_w9724_
	);
	LUT2 #(
		.INIT('h8)
	) name9192 (
		_w8983_,
		_w9021_,
		_w9725_
	);
	LUT3 #(
		.INIT('h2a)
	) name9193 (
		\u0_w_reg[3][26]/P0001 ,
		_w9049_,
		_w9050_,
		_w9726_
	);
	LUT4 #(
		.INIT('h7077)
	) name9194 (
		_w9721_,
		_w9724_,
		_w9725_,
		_w9726_,
		_w9727_
	);
	LUT4 #(
		.INIT('h0800)
	) name9195 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9728_
	);
	LUT4 #(
		.INIT('h002a)
	) name9196 (
		\u0_w_reg[3][25]/P0001 ,
		_w9068_,
		_w9015_,
		_w9728_,
		_w9729_
	);
	LUT2 #(
		.INIT('h8)
	) name9197 (
		\u0_w_reg[3][28]/P0001 ,
		_w8998_,
		_w9730_
	);
	LUT4 #(
		.INIT('h0020)
	) name9198 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9731_
	);
	LUT3 #(
		.INIT('h54)
	) name9199 (
		\u0_w_reg[3][26]/P0001 ,
		_w9050_,
		_w9731_,
		_w9732_
	);
	LUT3 #(
		.INIT('h10)
	) name9200 (
		_w9730_,
		_w9732_,
		_w9729_,
		_w9733_
	);
	LUT4 #(
		.INIT('h2000)
	) name9201 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9734_
	);
	LUT2 #(
		.INIT('h1)
	) name9202 (
		\u0_w_reg[3][25]/P0001 ,
		_w9734_,
		_w9735_
	);
	LUT4 #(
		.INIT('h0002)
	) name9203 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9736_
	);
	LUT3 #(
		.INIT('h07)
	) name9204 (
		_w8989_,
		_w9189_,
		_w9736_,
		_w9737_
	);
	LUT2 #(
		.INIT('h8)
	) name9205 (
		_w9735_,
		_w9737_,
		_w9738_
	);
	LUT3 #(
		.INIT('h40)
	) name9206 (
		\u0_w_reg[3][31]/P0001 ,
		_w8988_,
		_w8989_,
		_w9739_
	);
	LUT4 #(
		.INIT('h000e)
	) name9207 (
		_w9733_,
		_w9738_,
		_w9739_,
		_w9727_,
		_w9740_
	);
	LUT2 #(
		.INIT('h1)
	) name9208 (
		\u0_w_reg[3][24]/P0001 ,
		_w9740_,
		_w9741_
	);
	LUT3 #(
		.INIT('h56)
	) name9209 (
		\u0_w_reg[0][7]/P0001 ,
		_w9720_,
		_w9741_,
		_w9742_
	);
	LUT2 #(
		.INIT('h9)
	) name9210 (
		\u0_w_reg[1][7]/P0001 ,
		\u0_w_reg[2][7]/P0001 ,
		_w9743_
	);
	LUT4 #(
		.INIT('ha956)
	) name9211 (
		\u0_w_reg[0][7]/P0001 ,
		_w9720_,
		_w9741_,
		_w9743_,
		_w9744_
	);
	LUT3 #(
		.INIT('h8b)
	) name9212 (
		\key[39]_pad ,
		ld_pad,
		_w9744_,
		_w9745_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9213 (
		\key[115]_pad ,
		ld_pad,
		\u0_w_reg[0][19]/P0001 ,
		_w8971_,
		_w9746_
	);
	LUT4 #(
		.INIT('h1441)
	) name9214 (
		ld_pad,
		\u0_w_reg[0][19]/P0001 ,
		\u0_w_reg[1][19]/P0001 ,
		_w8971_,
		_w9747_
	);
	LUT2 #(
		.INIT('h8)
	) name9215 (
		\key[83]_pad ,
		ld_pad,
		_w9748_
	);
	LUT2 #(
		.INIT('he)
	) name9216 (
		_w9747_,
		_w9748_,
		_w9749_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9217 (
		\key[19]_pad ,
		ld_pad,
		\u0_w_reg[3][19]/P0001 ,
		_w8973_,
		_w9750_
	);
	LUT3 #(
		.INIT('hb8)
	) name9218 (
		\key[101]_pad ,
		ld_pad,
		_w9100_,
		_w9751_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name9219 (
		\key[69]_pad ,
		ld_pad,
		\u0_w_reg[1][5]/P0001 ,
		_w9100_,
		_w9752_
	);
	LUT4 #(
		.INIT('h1441)
	) name9220 (
		ld_pad,
		\u0_w_reg[3][5]/P0001 ,
		_w9100_,
		_w9101_,
		_w9753_
	);
	LUT2 #(
		.INIT('h8)
	) name9221 (
		\key[5]_pad ,
		ld_pad,
		_w9754_
	);
	LUT2 #(
		.INIT('he)
	) name9222 (
		_w9753_,
		_w9754_,
		_w9755_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name9223 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9239_,
		_w9716_,
		_w9756_
	);
	LUT4 #(
		.INIT('h0001)
	) name9224 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9757_
	);
	LUT4 #(
		.INIT('h0080)
	) name9225 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9758_
	);
	LUT3 #(
		.INIT('ha8)
	) name9226 (
		\u0_w_reg[3][26]/P0001 ,
		_w9757_,
		_w9758_,
		_w9759_
	);
	LUT3 #(
		.INIT('h02)
	) name9227 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		_w9760_
	);
	LUT4 #(
		.INIT('h0001)
	) name9228 (
		\u0_w_reg[3][25]/P0001 ,
		_w9048_,
		_w9693_,
		_w9760_,
		_w9761_
	);
	LUT3 #(
		.INIT('h40)
	) name9229 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9762_
	);
	LUT4 #(
		.INIT('h0002)
	) name9230 (
		\u0_w_reg[3][25]/P0001 ,
		_w9016_,
		_w9192_,
		_w9762_,
		_w9763_
	);
	LUT4 #(
		.INIT('h00ef)
	) name9231 (
		_w9759_,
		_w9756_,
		_w9761_,
		_w9763_,
		_w9764_
	);
	LUT3 #(
		.INIT('h07)
	) name9232 (
		_w9049_,
		_w9050_,
		_w9734_,
		_w9765_
	);
	LUT4 #(
		.INIT('h002a)
	) name9233 (
		\u0_w_reg[3][26]/P0001 ,
		_w8977_,
		_w9052_,
		_w9233_,
		_w9766_
	);
	LUT4 #(
		.INIT('h5155)
	) name9234 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9767_
	);
	LUT4 #(
		.INIT('hff9d)
	) name9235 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9768_
	);
	LUT3 #(
		.INIT('h40)
	) name9236 (
		_w9069_,
		_w9767_,
		_w9768_,
		_w9769_
	);
	LUT4 #(
		.INIT('h0040)
	) name9237 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9770_
	);
	LUT4 #(
		.INIT('h008a)
	) name9238 (
		\u0_w_reg[3][24]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w9037_,
		_w9770_,
		_w9771_
	);
	LUT4 #(
		.INIT('hf800)
	) name9239 (
		_w9765_,
		_w9766_,
		_w9769_,
		_w9771_,
		_w9772_
	);
	LUT2 #(
		.INIT('h4)
	) name9240 (
		_w9764_,
		_w9772_,
		_w9773_
	);
	LUT2 #(
		.INIT('h1)
	) name9241 (
		\u0_w_reg[3][27]/P0001 ,
		_w9708_,
		_w9774_
	);
	LUT2 #(
		.INIT('h4)
	) name9242 (
		\u0_w_reg[3][26]/P0001 ,
		_w9041_,
		_w9775_
	);
	LUT3 #(
		.INIT('h80)
	) name9243 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9776_
	);
	LUT3 #(
		.INIT('h45)
	) name9244 (
		\u0_w_reg[3][25]/P0001 ,
		_w9194_,
		_w9776_,
		_w9777_
	);
	LUT3 #(
		.INIT('h10)
	) name9245 (
		_w9774_,
		_w9775_,
		_w9777_,
		_w9778_
	);
	LUT2 #(
		.INIT('h8)
	) name9246 (
		_w9002_,
		_w9007_,
		_w9779_
	);
	LUT4 #(
		.INIT('h7ff8)
	) name9247 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9780_
	);
	LUT3 #(
		.INIT('h20)
	) name9248 (
		\u0_w_reg[3][25]/P0001 ,
		_w9716_,
		_w9780_,
		_w9781_
	);
	LUT2 #(
		.INIT('h4)
	) name9249 (
		_w9779_,
		_w9781_,
		_w9782_
	);
	LUT4 #(
		.INIT('h0001)
	) name9250 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9783_
	);
	LUT4 #(
		.INIT('h0007)
	) name9251 (
		_w8977_,
		_w9052_,
		_w9201_,
		_w9783_,
		_w9784_
	);
	LUT3 #(
		.INIT('hb9)
	) name9252 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9785_
	);
	LUT3 #(
		.INIT('h51)
	) name9253 (
		\u0_w_reg[3][24]/P0001 ,
		_w9681_,
		_w9785_,
		_w9786_
	);
	LUT3 #(
		.INIT('he0)
	) name9254 (
		\u0_w_reg[3][26]/P0001 ,
		_w9784_,
		_w9786_,
		_w9787_
	);
	LUT3 #(
		.INIT('he0)
	) name9255 (
		_w9778_,
		_w9782_,
		_w9787_,
		_w9788_
	);
	LUT2 #(
		.INIT('h8)
	) name9256 (
		_w8979_,
		_w9082_,
		_w9789_
	);
	LUT3 #(
		.INIT('h7b)
	) name9257 (
		\u0_w_reg[3][27]/P0001 ,
		_w8993_,
		_w9000_,
		_w9790_
	);
	LUT3 #(
		.INIT('h02)
	) name9258 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w9791_
	);
	LUT3 #(
		.INIT('h67)
	) name9259 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9792_
	);
	LUT4 #(
		.INIT('h7707)
	) name9260 (
		_w9093_,
		_w9094_,
		_w9791_,
		_w9792_,
		_w9793_
	);
	LUT4 #(
		.INIT('hba00)
	) name9261 (
		\u0_w_reg[3][26]/P0001 ,
		_w9789_,
		_w9790_,
		_w9793_,
		_w9794_
	);
	LUT4 #(
		.INIT('h4000)
	) name9262 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9795_
	);
	LUT4 #(
		.INIT('haa80)
	) name9263 (
		\u0_w_reg[3][30]/P0001 ,
		_w9057_,
		_w9068_,
		_w9795_,
		_w9796_
	);
	LUT4 #(
		.INIT('ha280)
	) name9264 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w9036_,
		_w9016_,
		_w9797_
	);
	LUT2 #(
		.INIT('h4)
	) name9265 (
		\u0_w_reg[3][26]/P0001 ,
		_w9196_,
		_w9798_
	);
	LUT2 #(
		.INIT('h4)
	) name9266 (
		\u0_w_reg[3][31]/P0001 ,
		_w9783_,
		_w9799_
	);
	LUT2 #(
		.INIT('h8)
	) name9267 (
		\u0_w_reg[3][27]/P0001 ,
		_w9091_,
		_w9800_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name9268 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9091_,
		_w9783_,
		_w9801_
	);
	LUT3 #(
		.INIT('h10)
	) name9269 (
		_w9797_,
		_w9798_,
		_w9801_,
		_w9802_
	);
	LUT4 #(
		.INIT('h3120)
	) name9270 (
		\u0_w_reg[3][25]/P0001 ,
		_w9796_,
		_w9802_,
		_w9794_,
		_w9803_
	);
	LUT4 #(
		.INIT('ha955)
	) name9271 (
		\u0_w_reg[0][0]/P0001 ,
		_w9773_,
		_w9788_,
		_w9803_,
		_w9804_
	);
	LUT2 #(
		.INIT('h9)
	) name9272 (
		\u0_w_reg[1][0]/P0001 ,
		\u0_w_reg[2][0]/P0001 ,
		_w9805_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9273 (
		\key[32]_pad ,
		ld_pad,
		_w9804_,
		_w9805_,
		_w9806_
	);
	LUT4 #(
		.INIT('h0007)
	) name9274 (
		_w9261_,
		_w9281_,
		_w9330_,
		_w9398_,
		_w9807_
	);
	LUT2 #(
		.INIT('h1)
	) name9275 (
		\u0_w_reg[3][2]/P0001 ,
		_w9807_,
		_w9808_
	);
	LUT4 #(
		.INIT('hbcfc)
	) name9276 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9809_
	);
	LUT2 #(
		.INIT('h2)
	) name9277 (
		_w9289_,
		_w9809_,
		_w9810_
	);
	LUT4 #(
		.INIT('h0302)
	) name9278 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9811_
	);
	LUT3 #(
		.INIT('h45)
	) name9279 (
		\u0_w_reg[3][1]/P0001 ,
		_w9375_,
		_w9811_,
		_w9812_
	);
	LUT4 #(
		.INIT('h135f)
	) name9280 (
		_w9290_,
		_w9303_,
		_w9375_,
		_w9424_,
		_w9813_
	);
	LUT3 #(
		.INIT('h40)
	) name9281 (
		_w9810_,
		_w9812_,
		_w9813_,
		_w9814_
	);
	LUT3 #(
		.INIT('h07)
	) name9282 (
		_w9261_,
		_w9262_,
		_w9353_,
		_w9815_
	);
	LUT4 #(
		.INIT('h0400)
	) name9283 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9816_
	);
	LUT4 #(
		.INIT('h0007)
	) name9284 (
		_w9261_,
		_w9262_,
		_w9353_,
		_w9816_,
		_w9817_
	);
	LUT3 #(
		.INIT('h20)
	) name9285 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9818_
	);
	LUT4 #(
		.INIT('h2def)
	) name9286 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9286_,
		_w9819_
	);
	LUT2 #(
		.INIT('h2)
	) name9287 (
		\u0_w_reg[3][1]/P0001 ,
		_w9308_,
		_w9820_
	);
	LUT4 #(
		.INIT('hd800)
	) name9288 (
		\u0_w_reg[3][2]/P0001 ,
		_w9819_,
		_w9817_,
		_w9820_,
		_w9821_
	);
	LUT3 #(
		.INIT('h0b)
	) name9289 (
		_w9808_,
		_w9814_,
		_w9821_,
		_w9822_
	);
	LUT4 #(
		.INIT('h0010)
	) name9290 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9823_
	);
	LUT4 #(
		.INIT('h0001)
	) name9291 (
		_w9352_,
		_w9364_,
		_w9422_,
		_w9823_,
		_w9824_
	);
	LUT3 #(
		.INIT('h0e)
	) name9292 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		_w9825_
	);
	LUT2 #(
		.INIT('h2)
	) name9293 (
		_w9345_,
		_w9825_,
		_w9826_
	);
	LUT4 #(
		.INIT('h0015)
	) name9294 (
		\u0_w_reg[3][1]/P0001 ,
		_w9274_,
		_w9307_,
		_w9316_,
		_w9827_
	);
	LUT3 #(
		.INIT('h01)
	) name9295 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9828_
	);
	LUT4 #(
		.INIT('h0002)
	) name9296 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9829_
	);
	LUT2 #(
		.INIT('h4)
	) name9297 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w9830_
	);
	LUT4 #(
		.INIT('h0040)
	) name9298 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9831_
	);
	LUT4 #(
		.INIT('h002a)
	) name9299 (
		\u0_w_reg[3][1]/P0001 ,
		_w9830_,
		_w9831_,
		_w9829_,
		_w9832_
	);
	LUT4 #(
		.INIT('h00bf)
	) name9300 (
		_w9826_,
		_w9824_,
		_w9827_,
		_w9832_,
		_w9833_
	);
	LUT4 #(
		.INIT('h0008)
	) name9301 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9834_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name9302 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9835_
	);
	LUT2 #(
		.INIT('h2)
	) name9303 (
		_w9289_,
		_w9835_,
		_w9836_
	);
	LUT3 #(
		.INIT('h8a)
	) name9304 (
		\u0_w_reg[3][0]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w9386_,
		_w9837_
	);
	LUT2 #(
		.INIT('h4)
	) name9305 (
		\u0_w_reg[3][6]/P0001 ,
		_w9823_,
		_w9838_
	);
	LUT4 #(
		.INIT('h2202)
	) name9306 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9839_
	);
	LUT4 #(
		.INIT('h135f)
	) name9307 (
		\u0_w_reg[3][5]/P0001 ,
		_w9298_,
		_w9422_,
		_w9839_,
		_w9840_
	);
	LUT4 #(
		.INIT('h1000)
	) name9308 (
		_w9836_,
		_w9838_,
		_w9837_,
		_w9840_,
		_w9841_
	);
	LUT4 #(
		.INIT('h0800)
	) name9309 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9842_
	);
	LUT2 #(
		.INIT('h2)
	) name9310 (
		\u0_w_reg[3][1]/P0001 ,
		_w9842_,
		_w9843_
	);
	LUT4 #(
		.INIT('h5155)
	) name9311 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9844_
	);
	LUT3 #(
		.INIT('h80)
	) name9312 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9845_
	);
	LUT3 #(
		.INIT('h10)
	) name9313 (
		_w9250_,
		_w9845_,
		_w9844_,
		_w9846_
	);
	LUT4 #(
		.INIT('haaa8)
	) name9314 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9847_
	);
	LUT2 #(
		.INIT('h4)
	) name9315 (
		_w9379_,
		_w9847_,
		_w9848_
	);
	LUT4 #(
		.INIT('h0040)
	) name9316 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9849_
	);
	LUT3 #(
		.INIT('h01)
	) name9317 (
		\u0_w_reg[3][1]/P0001 ,
		_w9279_,
		_w9849_,
		_w9850_
	);
	LUT4 #(
		.INIT('h0057)
	) name9318 (
		_w9843_,
		_w9846_,
		_w9848_,
		_w9850_,
		_w9851_
	);
	LUT3 #(
		.INIT('h80)
	) name9319 (
		\u0_w_reg[3][4]/P0001 ,
		_w9289_,
		_w9307_,
		_w9852_
	);
	LUT2 #(
		.INIT('h8)
	) name9320 (
		_w9301_,
		_w9412_,
		_w9853_
	);
	LUT4 #(
		.INIT('h0111)
	) name9321 (
		\u0_w_reg[3][0]/P0001 ,
		_w9322_,
		_w9301_,
		_w9412_,
		_w9854_
	);
	LUT2 #(
		.INIT('h4)
	) name9322 (
		_w9852_,
		_w9854_,
		_w9855_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name9323 (
		_w9833_,
		_w9841_,
		_w9851_,
		_w9855_,
		_w9856_
	);
	LUT3 #(
		.INIT('had)
	) name9324 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9857_
	);
	LUT3 #(
		.INIT('h02)
	) name9325 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w9858_
	);
	LUT4 #(
		.INIT('h7077)
	) name9326 (
		_w9257_,
		_w9312_,
		_w9857_,
		_w9858_,
		_w9859_
	);
	LUT4 #(
		.INIT('h5655)
	) name9327 (
		\u0_w_reg[0][10]/P0001 ,
		_w9856_,
		_w9822_,
		_w9859_,
		_w9860_
	);
	LUT2 #(
		.INIT('h9)
	) name9328 (
		\u0_w_reg[1][10]/P0001 ,
		\u0_w_reg[2][10]/P0001 ,
		_w9861_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9329 (
		\key[42]_pad ,
		ld_pad,
		_w9860_,
		_w9861_,
		_w9862_
	);
	LUT4 #(
		.INIT('hbfef)
	) name9330 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9863_
	);
	LUT2 #(
		.INIT('h1)
	) name9331 (
		\u0_w_reg[3][11]/P0001 ,
		_w9863_,
		_w9864_
	);
	LUT3 #(
		.INIT('h80)
	) name9332 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9865_
	);
	LUT2 #(
		.INIT('h4)
	) name9333 (
		_w8917_,
		_w9865_,
		_w9866_
	);
	LUT3 #(
		.INIT('h23)
	) name9334 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w8792_,
		_w9867_
	);
	LUT3 #(
		.INIT('h10)
	) name9335 (
		_w9864_,
		_w9866_,
		_w9867_,
		_w9868_
	);
	LUT4 #(
		.INIT('h0080)
	) name9336 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9869_
	);
	LUT3 #(
		.INIT('ha8)
	) name9337 (
		\u0_w_reg[3][11]/P0001 ,
		_w8797_,
		_w9869_,
		_w9870_
	);
	LUT4 #(
		.INIT('hfe00)
	) name9338 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w9871_
	);
	LUT3 #(
		.INIT('h01)
	) name9339 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9872_
	);
	LUT4 #(
		.INIT('h0100)
	) name9340 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9873_
	);
	LUT3 #(
		.INIT('h10)
	) name9341 (
		_w9872_,
		_w9873_,
		_w9871_,
		_w9874_
	);
	LUT2 #(
		.INIT('h4)
	) name9342 (
		_w9870_,
		_w9874_,
		_w9875_
	);
	LUT4 #(
		.INIT('h0001)
	) name9343 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w9876_
	);
	LUT4 #(
		.INIT('h0007)
	) name9344 (
		\u0_w_reg[3][13]/P0001 ,
		_w8809_,
		_w8927_,
		_w9876_,
		_w9877_
	);
	LUT3 #(
		.INIT('h02)
	) name9345 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9878_
	);
	LUT3 #(
		.INIT('hb9)
	) name9346 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9879_
	);
	LUT3 #(
		.INIT('h51)
	) name9347 (
		\u0_w_reg[3][8]/P0001 ,
		_w8855_,
		_w9879_,
		_w9880_
	);
	LUT3 #(
		.INIT('he0)
	) name9348 (
		\u0_w_reg[3][10]/P0001 ,
		_w9877_,
		_w9880_,
		_w9881_
	);
	LUT3 #(
		.INIT('he0)
	) name9349 (
		_w9868_,
		_w9875_,
		_w9881_,
		_w9882_
	);
	LUT4 #(
		.INIT('h3ffa)
	) name9350 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9883_
	);
	LUT4 #(
		.INIT('h80a2)
	) name9351 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		_w8879_,
		_w9883_,
		_w9884_
	);
	LUT2 #(
		.INIT('h8)
	) name9352 (
		_w8850_,
		_w8883_,
		_w9885_
	);
	LUT4 #(
		.INIT('h0010)
	) name9353 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9886_
	);
	LUT3 #(
		.INIT('h8a)
	) name9354 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9887_
	);
	LUT3 #(
		.INIT('h31)
	) name9355 (
		_w8825_,
		_w9886_,
		_w9887_,
		_w9888_
	);
	LUT4 #(
		.INIT('h5455)
	) name9356 (
		\u0_w_reg[3][9]/P0001 ,
		_w9884_,
		_w9885_,
		_w9888_,
		_w9889_
	);
	LUT4 #(
		.INIT('h2000)
	) name9357 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9890_
	);
	LUT3 #(
		.INIT('h07)
	) name9358 (
		_w8810_,
		_w8811_,
		_w9890_,
		_w9891_
	);
	LUT4 #(
		.INIT('h002a)
	) name9359 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		_w8809_,
		_w8956_,
		_w9892_
	);
	LUT4 #(
		.INIT('h5155)
	) name9360 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w9893_
	);
	LUT4 #(
		.INIT('h0040)
	) name9361 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9894_
	);
	LUT4 #(
		.INIT('hff9d)
	) name9362 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9895_
	);
	LUT3 #(
		.INIT('h40)
	) name9363 (
		_w8798_,
		_w9893_,
		_w9895_,
		_w9896_
	);
	LUT3 #(
		.INIT('h07)
	) name9364 (
		_w9891_,
		_w9892_,
		_w9896_,
		_w9897_
	);
	LUT3 #(
		.INIT('h54)
	) name9365 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9898_
	);
	LUT4 #(
		.INIT('h4041)
	) name9366 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9899_
	);
	LUT3 #(
		.INIT('ha8)
	) name9367 (
		\u0_w_reg[3][9]/P0001 ,
		_w8867_,
		_w9899_,
		_w9900_
	);
	LUT4 #(
		.INIT('h0200)
	) name9368 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9901_
	);
	LUT4 #(
		.INIT('h080c)
	) name9369 (
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][8]/P0001 ,
		_w8842_,
		_w9901_,
		_w9902_
	);
	LUT2 #(
		.INIT('h4)
	) name9370 (
		_w9900_,
		_w9902_,
		_w9903_
	);
	LUT3 #(
		.INIT('h10)
	) name9371 (
		_w9889_,
		_w9897_,
		_w9903_,
		_w9904_
	);
	LUT4 #(
		.INIT('h4000)
	) name9372 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9905_
	);
	LUT4 #(
		.INIT('haa80)
	) name9373 (
		\u0_w_reg[3][14]/P0001 ,
		_w8819_,
		_w8937_,
		_w9905_,
		_w9906_
	);
	LUT4 #(
		.INIT('h0004)
	) name9374 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9907_
	);
	LUT4 #(
		.INIT('hff4b)
	) name9375 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9908_
	);
	LUT2 #(
		.INIT('h2)
	) name9376 (
		_w8883_,
		_w9908_,
		_w9909_
	);
	LUT4 #(
		.INIT('haa80)
	) name9377 (
		\u0_w_reg[3][10]/P0001 ,
		_w8803_,
		_w8925_,
		_w8906_,
		_w9910_
	);
	LUT4 #(
		.INIT('h0040)
	) name9378 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9911_
	);
	LUT2 #(
		.INIT('h8)
	) name9379 (
		_w8878_,
		_w9911_,
		_w9912_
	);
	LUT3 #(
		.INIT('h15)
	) name9380 (
		\u0_w_reg[3][9]/P0001 ,
		_w8893_,
		_w8894_,
		_w9913_
	);
	LUT4 #(
		.INIT('h0100)
	) name9381 (
		_w9912_,
		_w9910_,
		_w9909_,
		_w9913_,
		_w9914_
	);
	LUT3 #(
		.INIT('h20)
	) name9382 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w9915_
	);
	LUT4 #(
		.INIT('h0020)
	) name9383 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w9916_
	);
	LUT4 #(
		.INIT('hffde)
	) name9384 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w9917_
	);
	LUT4 #(
		.INIT('h4055)
	) name9385 (
		\u0_w_reg[3][15]/P0001 ,
		_w8937_,
		_w9915_,
		_w9917_,
		_w9918_
	);
	LUT2 #(
		.INIT('h8)
	) name9386 (
		_w8786_,
		_w8851_,
		_w9919_
	);
	LUT3 #(
		.INIT('h8c)
	) name9387 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w8919_,
		_w9920_
	);
	LUT3 #(
		.INIT('h10)
	) name9388 (
		_w9919_,
		_w9918_,
		_w9920_,
		_w9921_
	);
	LUT3 #(
		.INIT('h54)
	) name9389 (
		_w9906_,
		_w9914_,
		_w9921_,
		_w9922_
	);
	LUT4 #(
		.INIT('ha955)
	) name9390 (
		\u0_w_reg[0][16]/P0001 ,
		_w9882_,
		_w9904_,
		_w9922_,
		_w9923_
	);
	LUT2 #(
		.INIT('h9)
	) name9391 (
		\u0_w_reg[1][16]/P0001 ,
		\u0_w_reg[2][16]/P0001 ,
		_w9924_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9392 (
		\key[48]_pad ,
		ld_pad,
		_w9923_,
		_w9924_,
		_w9925_
	);
	LUT4 #(
		.INIT('h0020)
	) name9393 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9926_
	);
	LUT4 #(
		.INIT('h0200)
	) name9394 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9927_
	);
	LUT3 #(
		.INIT('h01)
	) name9395 (
		_w9886_,
		_w9927_,
		_w9926_,
		_w9928_
	);
	LUT3 #(
		.INIT('h07)
	) name9396 (
		_w8796_,
		_w8828_,
		_w9869_,
		_w9929_
	);
	LUT3 #(
		.INIT('h0e)
	) name9397 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		_w9930_
	);
	LUT4 #(
		.INIT('h1101)
	) name9398 (
		\u0_w_reg[3][9]/P0001 ,
		_w8960_,
		_w9872_,
		_w9930_,
		_w9931_
	);
	LUT4 #(
		.INIT('h0002)
	) name9399 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9932_
	);
	LUT4 #(
		.INIT('h002a)
	) name9400 (
		\u0_w_reg[3][9]/P0001 ,
		_w8878_,
		_w9911_,
		_w9932_,
		_w9933_
	);
	LUT4 #(
		.INIT('h007f)
	) name9401 (
		_w9928_,
		_w9929_,
		_w9931_,
		_w9933_,
		_w9934_
	);
	LUT4 #(
		.INIT('h0008)
	) name9402 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9935_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name9403 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9936_
	);
	LUT2 #(
		.INIT('h2)
	) name9404 (
		_w8854_,
		_w9936_,
		_w9937_
	);
	LUT2 #(
		.INIT('h8)
	) name9405 (
		\u0_w_reg[3][10]/P0001 ,
		_w8842_,
		_w9938_
	);
	LUT3 #(
		.INIT('h2a)
	) name9406 (
		\u0_w_reg[3][8]/P0001 ,
		_w8803_,
		_w8925_,
		_w9939_
	);
	LUT3 #(
		.INIT('h4c)
	) name9407 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w9940_
	);
	LUT4 #(
		.INIT('h5100)
	) name9408 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w9941_
	);
	LUT4 #(
		.INIT('h0777)
	) name9409 (
		_w8791_,
		_w8905_,
		_w9940_,
		_w9941_,
		_w9942_
	);
	LUT4 #(
		.INIT('h1000)
	) name9410 (
		_w9937_,
		_w9938_,
		_w9939_,
		_w9942_,
		_w9943_
	);
	LUT4 #(
		.INIT('h0040)
	) name9411 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9944_
	);
	LUT3 #(
		.INIT('h01)
	) name9412 (
		\u0_w_reg[3][9]/P0001 ,
		_w8919_,
		_w9944_,
		_w9945_
	);
	LUT3 #(
		.INIT('h80)
	) name9413 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9946_
	);
	LUT3 #(
		.INIT('h04)
	) name9414 (
		_w8864_,
		_w9893_,
		_w9946_,
		_w9947_
	);
	LUT3 #(
		.INIT('h02)
	) name9415 (
		\u0_w_reg[3][10]/P0001 ,
		_w8818_,
		_w9872_,
		_w9948_
	);
	LUT4 #(
		.INIT('h0800)
	) name9416 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9949_
	);
	LUT2 #(
		.INIT('h2)
	) name9417 (
		\u0_w_reg[3][9]/P0001 ,
		_w9949_,
		_w9950_
	);
	LUT4 #(
		.INIT('h0155)
	) name9418 (
		_w9945_,
		_w9947_,
		_w9948_,
		_w9950_,
		_w9951_
	);
	LUT3 #(
		.INIT('h80)
	) name9419 (
		\u0_w_reg[3][10]/P0001 ,
		_w8793_,
		_w8943_,
		_w9952_
	);
	LUT2 #(
		.INIT('h1)
	) name9420 (
		\u0_w_reg[3][8]/P0001 ,
		_w8861_,
		_w9953_
	);
	LUT3 #(
		.INIT('h10)
	) name9421 (
		_w8897_,
		_w9952_,
		_w9953_,
		_w9954_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name9422 (
		_w9934_,
		_w9943_,
		_w9951_,
		_w9954_,
		_w9955_
	);
	LUT3 #(
		.INIT('h3d)
	) name9423 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9956_
	);
	LUT2 #(
		.INIT('h2)
	) name9424 (
		_w8793_,
		_w9956_,
		_w9957_
	);
	LUT3 #(
		.INIT('had)
	) name9425 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9958_
	);
	LUT3 #(
		.INIT('h31)
	) name9426 (
		_w8815_,
		_w8925_,
		_w9958_,
		_w9959_
	);
	LUT4 #(
		.INIT('h4c44)
	) name9427 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w9957_,
		_w9959_,
		_w9960_
	);
	LUT4 #(
		.INIT('hbcfc)
	) name9428 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9961_
	);
	LUT2 #(
		.INIT('h2)
	) name9429 (
		\u0_w_reg[3][11]/P0001 ,
		_w9961_,
		_w9962_
	);
	LUT4 #(
		.INIT('h3010)
	) name9430 (
		_w8815_,
		_w8919_,
		_w8962_,
		_w9958_,
		_w9963_
	);
	LUT4 #(
		.INIT('h0004)
	) name9431 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9964_
	);
	LUT2 #(
		.INIT('h1)
	) name9432 (
		\u0_w_reg[3][10]/P0001 ,
		_w9964_,
		_w9965_
	);
	LUT4 #(
		.INIT('h8000)
	) name9433 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w9966_
	);
	LUT4 #(
		.INIT('h0203)
	) name9434 (
		\u0_w_reg[3][15]/P0001 ,
		_w8922_,
		_w9907_,
		_w9966_,
		_w9967_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name9435 (
		_w9962_,
		_w9963_,
		_w9965_,
		_w9967_,
		_w9968_
	);
	LUT4 #(
		.INIT('h000b)
	) name9436 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w9969_
	);
	LUT2 #(
		.INIT('h4)
	) name9437 (
		_w8863_,
		_w9969_,
		_w9970_
	);
	LUT3 #(
		.INIT('h54)
	) name9438 (
		_w9960_,
		_w9968_,
		_w9970_,
		_w9971_
	);
	LUT3 #(
		.INIT('h13)
	) name9439 (
		\u0_w_reg[3][15]/P0001 ,
		_w8860_,
		_w9966_,
		_w9972_
	);
	LUT4 #(
		.INIT('h0103)
	) name9440 (
		\u0_w_reg[3][15]/P0001 ,
		_w8809_,
		_w8860_,
		_w9966_,
		_w9973_
	);
	LUT4 #(
		.INIT('hc0c4)
	) name9441 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w8839_,
		_w9973_,
		_w9974_
	);
	LUT2 #(
		.INIT('h1)
	) name9442 (
		_w8957_,
		_w9974_,
		_w9975_
	);
	LUT4 #(
		.INIT('h5655)
	) name9443 (
		\u0_w_reg[0][18]/P0001 ,
		_w9971_,
		_w9955_,
		_w9975_,
		_w9976_
	);
	LUT2 #(
		.INIT('h9)
	) name9444 (
		\u0_w_reg[1][18]/P0001 ,
		\u0_w_reg[2][18]/P0001 ,
		_w9977_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9445 (
		\key[50]_pad ,
		ld_pad,
		_w9976_,
		_w9977_,
		_w9978_
	);
	LUT2 #(
		.INIT('h8)
	) name9446 (
		_w8980_,
		_w9009_,
		_w9979_
	);
	LUT3 #(
		.INIT('h04)
	) name9447 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9980_
	);
	LUT4 #(
		.INIT('h0004)
	) name9448 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9981_
	);
	LUT3 #(
		.INIT('h0b)
	) name9449 (
		\u0_w_reg[3][26]/P0001 ,
		_w9058_,
		_w9981_,
		_w9982_
	);
	LUT2 #(
		.INIT('h2)
	) name9450 (
		\u0_w_reg[3][26]/P0001 ,
		_w9685_,
		_w9983_
	);
	LUT4 #(
		.INIT('h0200)
	) name9451 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9984_
	);
	LUT4 #(
		.INIT('h2000)
	) name9452 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9985_
	);
	LUT4 #(
		.INIT('h0001)
	) name9453 (
		\u0_w_reg[3][25]/P0001 ,
		_w9693_,
		_w9984_,
		_w9985_,
		_w9986_
	);
	LUT4 #(
		.INIT('h1000)
	) name9454 (
		_w9983_,
		_w9979_,
		_w9986_,
		_w9982_,
		_w9987_
	);
	LUT4 #(
		.INIT('hea40)
	) name9455 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w9061_,
		_w9023_,
		_w9988_
	);
	LUT2 #(
		.INIT('h2)
	) name9456 (
		\u0_w_reg[3][25]/P0001 ,
		_w9988_,
		_w9989_
	);
	LUT4 #(
		.INIT('h0008)
	) name9457 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9990_
	);
	LUT4 #(
		.INIT('h3fd7)
	) name9458 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9991_
	);
	LUT2 #(
		.INIT('h2)
	) name9459 (
		_w8989_,
		_w9991_,
		_w9992_
	);
	LUT4 #(
		.INIT('h0100)
	) name9460 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9993_
	);
	LUT2 #(
		.INIT('h4)
	) name9461 (
		\u0_w_reg[3][29]/P0001 ,
		_w9993_,
		_w9994_
	);
	LUT3 #(
		.INIT('h2a)
	) name9462 (
		\u0_w_reg[3][24]/P0001 ,
		_w8979_,
		_w9082_,
		_w9995_
	);
	LUT4 #(
		.INIT('h0222)
	) name9463 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w9996_
	);
	LUT4 #(
		.INIT('h0777)
	) name9464 (
		_w9068_,
		_w9035_,
		_w9677_,
		_w9996_,
		_w9997_
	);
	LUT4 #(
		.INIT('h1000)
	) name9465 (
		_w9992_,
		_w9994_,
		_w9995_,
		_w9997_,
		_w9998_
	);
	LUT3 #(
		.INIT('he0)
	) name9466 (
		_w9987_,
		_w9989_,
		_w9998_,
		_w9999_
	);
	LUT3 #(
		.INIT('h80)
	) name9467 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10000_
	);
	LUT3 #(
		.INIT('h04)
	) name9468 (
		_w9211_,
		_w9767_,
		_w10000_,
		_w10001_
	);
	LUT3 #(
		.INIT('h02)
	) name9469 (
		\u0_w_reg[3][26]/P0001 ,
		_w9056_,
		_w8980_,
		_w10002_
	);
	LUT4 #(
		.INIT('h888a)
	) name9470 (
		\u0_w_reg[3][25]/P0001 ,
		_w9728_,
		_w10001_,
		_w10002_,
		_w10003_
	);
	LUT4 #(
		.INIT('h0040)
	) name9471 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10004_
	);
	LUT3 #(
		.INIT('h54)
	) name9472 (
		\u0_w_reg[3][25]/P0001 ,
		_w9196_,
		_w10004_,
		_w10005_
	);
	LUT2 #(
		.INIT('h8)
	) name9473 (
		_w9020_,
		_w9239_,
		_w10006_
	);
	LUT4 #(
		.INIT('h0111)
	) name9474 (
		\u0_w_reg[3][24]/P0001 ,
		_w9031_,
		_w9090_,
		_w9091_,
		_w10007_
	);
	LUT3 #(
		.INIT('h10)
	) name9475 (
		_w10006_,
		_w10005_,
		_w10007_,
		_w10008_
	);
	LUT2 #(
		.INIT('h4)
	) name9476 (
		_w10003_,
		_w10008_,
		_w10009_
	);
	LUT3 #(
		.INIT('h07)
	) name9477 (
		_w8983_,
		_w9021_,
		_w9028_,
		_w10010_
	);
	LUT4 #(
		.INIT('h0013)
	) name9478 (
		_w8983_,
		_w8978_,
		_w9021_,
		_w9028_,
		_w10011_
	);
	LUT3 #(
		.INIT('hc8)
	) name9479 (
		\u0_w_reg[3][26]/P0001 ,
		_w8999_,
		_w10011_,
		_w10012_
	);
	LUT2 #(
		.INIT('h1)
	) name9480 (
		_w9091_,
		_w9206_,
		_w10013_
	);
	LUT4 #(
		.INIT('hbcfc)
	) name9481 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10014_
	);
	LUT4 #(
		.INIT('h0a02)
	) name9482 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w9196_,
		_w10014_,
		_w10015_
	);
	LUT3 #(
		.INIT('h07)
	) name9483 (
		_w9721_,
		_w10013_,
		_w10015_,
		_w10016_
	);
	LUT3 #(
		.INIT('h15)
	) name9484 (
		\u0_w_reg[3][25]/P0001 ,
		_w9197_,
		_w9709_,
		_w10017_
	);
	LUT4 #(
		.INIT('h000b)
	) name9485 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w10018_
	);
	LUT2 #(
		.INIT('h4)
	) name9486 (
		_w9012_,
		_w10018_,
		_w10019_
	);
	LUT2 #(
		.INIT('h2)
	) name9487 (
		_w10017_,
		_w10019_,
		_w10020_
	);
	LUT3 #(
		.INIT('had)
	) name9488 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10021_
	);
	LUT2 #(
		.INIT('h2)
	) name9489 (
		_w9791_,
		_w10021_,
		_w10022_
	);
	LUT2 #(
		.INIT('h8)
	) name9490 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		_w10023_
	);
	LUT3 #(
		.INIT('he0)
	) name9491 (
		_w9058_,
		_w9203_,
		_w10023_,
		_w10024_
	);
	LUT3 #(
		.INIT('h80)
	) name9492 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w10025_
	);
	LUT4 #(
		.INIT('h153f)
	) name9493 (
		_w9070_,
		_w9090_,
		_w9233_,
		_w10025_,
		_w10026_
	);
	LUT3 #(
		.INIT('h10)
	) name9494 (
		_w10024_,
		_w10022_,
		_w10026_,
		_w10027_
	);
	LUT4 #(
		.INIT('hba00)
	) name9495 (
		_w10012_,
		_w10016_,
		_w10020_,
		_w10027_,
		_w10028_
	);
	LUT4 #(
		.INIT('ha955)
	) name9496 (
		\u0_w_reg[0][2]/P0001 ,
		_w9999_,
		_w10009_,
		_w10028_,
		_w10029_
	);
	LUT3 #(
		.INIT('h96)
	) name9497 (
		\u0_w_reg[1][2]/P0001 ,
		\u0_w_reg[2][2]/P0001 ,
		_w10029_,
		_w10030_
	);
	LUT4 #(
		.INIT('h4114)
	) name9498 (
		ld_pad,
		\u0_w_reg[1][2]/P0001 ,
		\u0_w_reg[2][2]/P0001 ,
		_w10029_,
		_w10031_
	);
	LUT2 #(
		.INIT('h8)
	) name9499 (
		\key[34]_pad ,
		ld_pad,
		_w10032_
	);
	LUT2 #(
		.INIT('he)
	) name9500 (
		_w10031_,
		_w10032_,
		_w10033_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name9501 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10034_
	);
	LUT4 #(
		.INIT('h20aa)
	) name9502 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w9353_,
		_w10034_,
		_w10035_
	);
	LUT2 #(
		.INIT('h8)
	) name9503 (
		_w9259_,
		_w9281_,
		_w10036_
	);
	LUT4 #(
		.INIT('h2000)
	) name9504 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10037_
	);
	LUT3 #(
		.INIT('h07)
	) name9505 (
		_w9303_,
		_w9372_,
		_w10037_,
		_w10038_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9506 (
		\u0_w_reg[3][1]/P0001 ,
		_w10036_,
		_w10035_,
		_w10038_,
		_w10039_
	);
	LUT2 #(
		.INIT('h1)
	) name9507 (
		_w9353_,
		_w9349_,
		_w10040_
	);
	LUT3 #(
		.INIT('h54)
	) name9508 (
		\u0_w_reg[3][2]/P0001 ,
		_w9353_,
		_w9349_,
		_w10041_
	);
	LUT3 #(
		.INIT('ha8)
	) name9509 (
		\u0_w_reg[3][2]/P0001 ,
		_w9262_,
		_w9287_,
		_w10042_
	);
	LUT3 #(
		.INIT('h15)
	) name9510 (
		_w9322_,
		_w9303_,
		_w9424_,
		_w10043_
	);
	LUT4 #(
		.INIT('h5455)
	) name9511 (
		\u0_w_reg[3][1]/P0001 ,
		_w10041_,
		_w10042_,
		_w10043_,
		_w10044_
	);
	LUT2 #(
		.INIT('h1)
	) name9512 (
		_w9257_,
		_w9378_,
		_w10045_
	);
	LUT3 #(
		.INIT('h08)
	) name9513 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w10046_
	);
	LUT3 #(
		.INIT('h40)
	) name9514 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w10047_
	);
	LUT4 #(
		.INIT('h135f)
	) name9515 (
		_w9303_,
		_w9365_,
		_w10046_,
		_w10047_,
		_w10048_
	);
	LUT4 #(
		.INIT('hd500)
	) name9516 (
		\u0_w_reg[3][2]/P0001 ,
		_w9283_,
		_w10045_,
		_w10048_,
		_w10049_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9517 (
		\u0_w_reg[3][0]/P0001 ,
		_w10044_,
		_w10039_,
		_w10049_,
		_w10050_
	);
	LUT4 #(
		.INIT('h0001)
	) name9518 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w10051_
	);
	LUT3 #(
		.INIT('h2a)
	) name9519 (
		\u0_w_reg[3][2]/P0001 ,
		_w9307_,
		_w9375_,
		_w10052_
	);
	LUT4 #(
		.INIT('h002a)
	) name9520 (
		\u0_w_reg[3][2]/P0001 ,
		_w9307_,
		_w9375_,
		_w10051_,
		_w10053_
	);
	LUT4 #(
		.INIT('h0015)
	) name9521 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w9251_,
		_w9300_,
		_w10054_
	);
	LUT4 #(
		.INIT('h0004)
	) name9522 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w10055_
	);
	LUT3 #(
		.INIT('h0b)
	) name9523 (
		_w9314_,
		_w9426_,
		_w10055_,
		_w10056_
	);
	LUT3 #(
		.INIT('h15)
	) name9524 (
		_w10053_,
		_w10054_,
		_w10056_,
		_w10057_
	);
	LUT4 #(
		.INIT('h0100)
	) name9525 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10058_
	);
	LUT4 #(
		.INIT('h0001)
	) name9526 (
		\u0_w_reg[3][1]/P0001 ,
		_w9275_,
		_w9831_,
		_w10058_,
		_w10059_
	);
	LUT4 #(
		.INIT('h0200)
	) name9527 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10060_
	);
	LUT4 #(
		.INIT('h153f)
	) name9528 (
		_w9289_,
		_w9307_,
		_w9375_,
		_w9424_,
		_w10061_
	);
	LUT3 #(
		.INIT('h40)
	) name9529 (
		_w10060_,
		_w10059_,
		_w10061_,
		_w10062_
	);
	LUT3 #(
		.INIT('h80)
	) name9530 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10063_
	);
	LUT3 #(
		.INIT('h7e)
	) name9531 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10064_
	);
	LUT4 #(
		.INIT('h0072)
	) name9532 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w9378_,
		_w10064_,
		_w10065_
	);
	LUT3 #(
		.INIT('h2a)
	) name9533 (
		\u0_w_reg[3][1]/P0001 ,
		_w9261_,
		_w9281_,
		_w10066_
	);
	LUT2 #(
		.INIT('h4)
	) name9534 (
		_w10065_,
		_w10066_,
		_w10067_
	);
	LUT4 #(
		.INIT('h4445)
	) name9535 (
		\u0_w_reg[3][0]/P0001 ,
		_w10057_,
		_w10062_,
		_w10067_,
		_w10068_
	);
	LUT4 #(
		.INIT('hf7fa)
	) name9536 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10069_
	);
	LUT4 #(
		.INIT('h0002)
	) name9537 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10070_
	);
	LUT4 #(
		.INIT('haa02)
	) name9538 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w10069_,
		_w10070_,
		_w10071_
	);
	LUT3 #(
		.INIT('ha8)
	) name9539 (
		\u0_w_reg[3][1]/P0001 ,
		_w9853_,
		_w10071_,
		_w10072_
	);
	LUT3 #(
		.INIT('h54)
	) name9540 (
		\u0_w_reg[3][2]/P0001 ,
		_w9327_,
		_w9842_,
		_w10073_
	);
	LUT4 #(
		.INIT('h0007)
	) name9541 (
		_w9254_,
		_w9290_,
		_w9319_,
		_w9330_,
		_w10074_
	);
	LUT4 #(
		.INIT('h23af)
	) name9542 (
		\u0_w_reg[3][2]/P0001 ,
		_w9314_,
		_w9322_,
		_w9381_,
		_w10075_
	);
	LUT4 #(
		.INIT('h4555)
	) name9543 (
		\u0_w_reg[3][1]/P0001 ,
		_w10073_,
		_w10074_,
		_w10075_,
		_w10076_
	);
	LUT4 #(
		.INIT('h3230)
	) name9544 (
		\u0_w_reg[3][6]/P0001 ,
		_w9274_,
		_w9346_,
		_w9349_,
		_w10077_
	);
	LUT2 #(
		.INIT('h1)
	) name9545 (
		_w9276_,
		_w10077_,
		_w10078_
	);
	LUT3 #(
		.INIT('h10)
	) name9546 (
		_w10072_,
		_w10076_,
		_w10078_,
		_w10079_
	);
	LUT4 #(
		.INIT('h5655)
	) name9547 (
		\u0_w_reg[0][14]/P0001 ,
		_w10068_,
		_w10050_,
		_w10079_,
		_w10080_
	);
	LUT2 #(
		.INIT('h9)
	) name9548 (
		\u0_w_reg[1][14]/P0001 ,
		\u0_w_reg[2][14]/P0001 ,
		_w10081_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9549 (
		\key[46]_pad ,
		ld_pad,
		_w10080_,
		_w10081_,
		_w10082_
	);
	LUT3 #(
		.INIT('h54)
	) name9550 (
		\u0_w_reg[3][10]/P0001 ,
		_w8859_,
		_w8860_,
		_w10083_
	);
	LUT4 #(
		.INIT('hfda8)
	) name9551 (
		\u0_w_reg[3][10]/P0001 ,
		_w8875_,
		_w8943_,
		_w9964_,
		_w10084_
	);
	LUT2 #(
		.INIT('h1)
	) name9552 (
		\u0_w_reg[3][9]/P0001 ,
		_w8861_,
		_w10085_
	);
	LUT3 #(
		.INIT('h10)
	) name9553 (
		_w10084_,
		_w10083_,
		_w10085_,
		_w10086_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name9554 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10087_
	);
	LUT4 #(
		.INIT('h80aa)
	) name9555 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8816_,
		_w10087_,
		_w10088_
	);
	LUT3 #(
		.INIT('h2a)
	) name9556 (
		\u0_w_reg[3][9]/P0001 ,
		_w8829_,
		_w8883_,
		_w10089_
	);
	LUT3 #(
		.INIT('h20)
	) name9557 (
		_w9891_,
		_w10088_,
		_w10089_,
		_w10090_
	);
	LUT3 #(
		.INIT('h01)
	) name9558 (
		_w8787_,
		_w8870_,
		_w8948_,
		_w10091_
	);
	LUT3 #(
		.INIT('h01)
	) name9559 (
		\u0_w_reg[3][10]/P0001 ,
		_w8834_,
		_w9911_,
		_w10092_
	);
	LUT3 #(
		.INIT('h07)
	) name9560 (
		_w8814_,
		_w10091_,
		_w10092_,
		_w10093_
	);
	LUT4 #(
		.INIT('haa02)
	) name9561 (
		\u0_w_reg[3][8]/P0001 ,
		_w10086_,
		_w10090_,
		_w10093_,
		_w10094_
	);
	LUT4 #(
		.INIT('h0100)
	) name9562 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10095_
	);
	LUT3 #(
		.INIT('h01)
	) name9563 (
		_w9905_,
		_w9911_,
		_w10095_,
		_w10096_
	);
	LUT2 #(
		.INIT('h8)
	) name9564 (
		_w8854_,
		_w9878_,
		_w10097_
	);
	LUT2 #(
		.INIT('h8)
	) name9565 (
		_w8808_,
		_w8838_,
		_w10098_
	);
	LUT4 #(
		.INIT('h0015)
	) name9566 (
		\u0_w_reg[3][9]/P0001 ,
		_w8808_,
		_w8838_,
		_w9901_,
		_w10099_
	);
	LUT3 #(
		.INIT('h40)
	) name9567 (
		_w10097_,
		_w10096_,
		_w10099_,
		_w10100_
	);
	LUT2 #(
		.INIT('h4)
	) name9568 (
		_w8865_,
		_w8937_,
		_w10101_
	);
	LUT2 #(
		.INIT('h4)
	) name9569 (
		\u0_w_reg[3][10]/P0001 ,
		_w8870_,
		_w10102_
	);
	LUT3 #(
		.INIT('h8c)
	) name9570 (
		\u0_w_reg[3][15]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w9966_,
		_w10103_
	);
	LUT3 #(
		.INIT('h10)
	) name9571 (
		_w10101_,
		_w10102_,
		_w10103_,
		_w10104_
	);
	LUT4 #(
		.INIT('haa80)
	) name9572 (
		\u0_w_reg[3][10]/P0001 ,
		_w8808_,
		_w8838_,
		_w9876_,
		_w10105_
	);
	LUT3 #(
		.INIT('he6)
	) name9573 (
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10106_
	);
	LUT2 #(
		.INIT('h2)
	) name9574 (
		_w8808_,
		_w10106_,
		_w10107_
	);
	LUT3 #(
		.INIT('h13)
	) name9575 (
		_w8825_,
		_w8918_,
		_w9898_,
		_w10108_
	);
	LUT4 #(
		.INIT('h2322)
	) name9576 (
		\u0_w_reg[3][10]/P0001 ,
		_w10105_,
		_w10107_,
		_w10108_,
		_w10109_
	);
	LUT4 #(
		.INIT('h0155)
	) name9577 (
		\u0_w_reg[3][8]/P0001 ,
		_w10100_,
		_w10104_,
		_w10109_,
		_w10110_
	);
	LUT3 #(
		.INIT('h02)
	) name9578 (
		\u0_w_reg[3][10]/P0001 ,
		_w8849_,
		_w8889_,
		_w10111_
	);
	LUT4 #(
		.INIT('h0001)
	) name9579 (
		\u0_w_reg[3][10]/P0001 ,
		_w8861_,
		_w8867_,
		_w9949_,
		_w10112_
	);
	LUT2 #(
		.INIT('h1)
	) name9580 (
		_w8906_,
		_w8922_,
		_w10113_
	);
	LUT4 #(
		.INIT('h0155)
	) name9581 (
		\u0_w_reg[3][9]/P0001 ,
		_w10111_,
		_w10112_,
		_w10113_,
		_w10114_
	);
	LUT2 #(
		.INIT('h8)
	) name9582 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w10115_
	);
	LUT4 #(
		.INIT('hf7fa)
	) name9583 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10116_
	);
	LUT4 #(
		.INIT('hc0d0)
	) name9584 (
		\u0_w_reg[3][12]/P0001 ,
		_w8805_,
		_w10115_,
		_w10116_,
		_w10117_
	);
	LUT2 #(
		.INIT('h4)
	) name9585 (
		\u0_w_reg[3][15]/P0001 ,
		_w9876_,
		_w10118_
	);
	LUT4 #(
		.INIT('hff7a)
	) name9586 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10119_
	);
	LUT2 #(
		.INIT('h2)
	) name9587 (
		_w8851_,
		_w10119_,
		_w10120_
	);
	LUT3 #(
		.INIT('h80)
	) name9588 (
		_w8810_,
		_w8823_,
		_w8896_,
		_w10121_
	);
	LUT4 #(
		.INIT('h0001)
	) name9589 (
		_w8934_,
		_w10118_,
		_w10120_,
		_w10121_,
		_w10122_
	);
	LUT3 #(
		.INIT('h10)
	) name9590 (
		_w10114_,
		_w10117_,
		_w10122_,
		_w10123_
	);
	LUT4 #(
		.INIT('h5655)
	) name9591 (
		\u0_w_reg[0][22]/P0001 ,
		_w10094_,
		_w10110_,
		_w10123_,
		_w10124_
	);
	LUT2 #(
		.INIT('h9)
	) name9592 (
		\u0_w_reg[1][22]/P0001 ,
		\u0_w_reg[2][22]/P0001 ,
		_w10125_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9593 (
		\key[54]_pad ,
		ld_pad,
		_w10124_,
		_w10125_,
		_w10126_
	);
	LUT2 #(
		.INIT('h4)
	) name9594 (
		\key[38]_pad ,
		ld_pad,
		_w10127_
	);
	LUT3 #(
		.INIT('h2a)
	) name9595 (
		\u0_w_reg[3][25]/P0001 ,
		_w9064_,
		_w9197_,
		_w10128_
	);
	LUT4 #(
		.INIT('h0111)
	) name9596 (
		\u0_w_reg[3][25]/P0001 ,
		_w9031_,
		_w9197_,
		_w9709_,
		_w10129_
	);
	LUT4 #(
		.INIT('h153f)
	) name9597 (
		_w9029_,
		_w9765_,
		_w10128_,
		_w10129_,
		_w10130_
	);
	LUT3 #(
		.INIT('h01)
	) name9598 (
		\u0_w_reg[3][26]/P0001 ,
		_w9061_,
		_w8992_,
		_w10131_
	);
	LUT2 #(
		.INIT('h4)
	) name9599 (
		_w10130_,
		_w10131_,
		_w10132_
	);
	LUT4 #(
		.INIT('hfb5f)
	) name9600 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10133_
	);
	LUT3 #(
		.INIT('h70)
	) name9601 (
		_w9014_,
		_w9203_,
		_w10133_,
		_w10134_
	);
	LUT3 #(
		.INIT('h80)
	) name9602 (
		_w9765_,
		_w10128_,
		_w10134_,
		_w10135_
	);
	LUT2 #(
		.INIT('h1)
	) name9603 (
		_w9076_,
		_w9021_,
		_w10136_
	);
	LUT2 #(
		.INIT('h8)
	) name9604 (
		_w10129_,
		_w10136_,
		_w10137_
	);
	LUT2 #(
		.INIT('h2)
	) name9605 (
		\u0_w_reg[3][26]/P0001 ,
		_w9037_,
		_w10138_
	);
	LUT4 #(
		.INIT('h0007)
	) name9606 (
		\u0_w_reg[3][31]/P0001 ,
		_w9044_,
		_w9013_,
		_w9225_,
		_w10139_
	);
	LUT2 #(
		.INIT('h8)
	) name9607 (
		_w10138_,
		_w10139_,
		_w10140_
	);
	LUT4 #(
		.INIT('h02aa)
	) name9608 (
		\u0_w_reg[3][24]/P0001 ,
		_w10135_,
		_w10137_,
		_w10140_,
		_w10141_
	);
	LUT4 #(
		.INIT('h115f)
	) name9609 (
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9212_,
		_w9760_,
		_w10142_
	);
	LUT2 #(
		.INIT('h1)
	) name9610 (
		\u0_w_reg[3][26]/P0001 ,
		_w9195_,
		_w10143_
	);
	LUT4 #(
		.INIT('h0004)
	) name9611 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w10144_
	);
	LUT3 #(
		.INIT('h01)
	) name9612 (
		\u0_w_reg[3][26]/P0001 ,
		_w9195_,
		_w10144_,
		_w10145_
	);
	LUT4 #(
		.INIT('h002a)
	) name9613 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w8998_,
		_w9783_,
		_w10146_
	);
	LUT3 #(
		.INIT('h07)
	) name9614 (
		_w10142_,
		_w10145_,
		_w10146_,
		_w10147_
	);
	LUT4 #(
		.INIT('h0200)
	) name9615 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10148_
	);
	LUT4 #(
		.INIT('h0007)
	) name9616 (
		_w8989_,
		_w9709_,
		_w9993_,
		_w10148_,
		_w10149_
	);
	LUT3 #(
		.INIT('h01)
	) name9617 (
		\u0_w_reg[3][25]/P0001 ,
		_w9061_,
		_w9795_,
		_w10150_
	);
	LUT3 #(
		.INIT('h40)
	) name9618 (
		_w9730_,
		_w10150_,
		_w10149_,
		_w10151_
	);
	LUT3 #(
		.INIT('h80)
	) name9619 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10152_
	);
	LUT3 #(
		.INIT('h7e)
	) name9620 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10153_
	);
	LUT2 #(
		.INIT('h2)
	) name9621 (
		_w9068_,
		_w10153_,
		_w10154_
	);
	LUT2 #(
		.INIT('h4)
	) name9622 (
		\u0_w_reg[3][26]/P0001 ,
		_w9013_,
		_w10155_
	);
	LUT3 #(
		.INIT('h8a)
	) name9623 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9084_,
		_w10156_
	);
	LUT3 #(
		.INIT('h10)
	) name9624 (
		_w10155_,
		_w10154_,
		_w10156_,
		_w10157_
	);
	LUT4 #(
		.INIT('h4445)
	) name9625 (
		\u0_w_reg[3][24]/P0001 ,
		_w10147_,
		_w10151_,
		_w10157_,
		_w10158_
	);
	LUT4 #(
		.INIT('h0001)
	) name9626 (
		\u0_w_reg[3][26]/P0001 ,
		_w9031_,
		_w9016_,
		_w9728_,
		_w10159_
	);
	LUT4 #(
		.INIT('h0002)
	) name9627 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10160_
	);
	LUT3 #(
		.INIT('h02)
	) name9628 (
		\u0_w_reg[3][26]/P0001 ,
		_w9223_,
		_w10160_,
		_w10161_
	);
	LUT2 #(
		.INIT('h1)
	) name9629 (
		_w9206_,
		_w9186_,
		_w10162_
	);
	LUT4 #(
		.INIT('h0155)
	) name9630 (
		\u0_w_reg[3][25]/P0001 ,
		_w10159_,
		_w10161_,
		_w10162_,
		_w10163_
	);
	LUT4 #(
		.INIT('hdff3)
	) name9631 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10164_
	);
	LUT4 #(
		.INIT('hc0d0)
	) name9632 (
		\u0_w_reg[3][30]/P0001 ,
		_w9079_,
		_w10023_,
		_w10164_,
		_w10165_
	);
	LUT4 #(
		.INIT('haa80)
	) name9633 (
		\u0_w_reg[3][26]/P0001 ,
		_w9026_,
		_w9194_,
		_w9757_,
		_w10166_
	);
	LUT3 #(
		.INIT('h80)
	) name9634 (
		\u0_w_reg[3][25]/P0001 ,
		_w9090_,
		_w9091_,
		_w10167_
	);
	LUT4 #(
		.INIT('h0001)
	) name9635 (
		_w9218_,
		_w9799_,
		_w10166_,
		_w10167_,
		_w10168_
	);
	LUT3 #(
		.INIT('h10)
	) name9636 (
		_w10163_,
		_w10165_,
		_w10168_,
		_w10169_
	);
	LUT4 #(
		.INIT('h0b00)
	) name9637 (
		_w10132_,
		_w10141_,
		_w10158_,
		_w10169_,
		_w10170_
	);
	LUT2 #(
		.INIT('h9)
	) name9638 (
		\u0_w_reg[1][6]/P0001 ,
		\u0_w_reg[2][6]/P0001 ,
		_w10171_
	);
	LUT3 #(
		.INIT('h69)
	) name9639 (
		\u0_w_reg[0][6]/P0001 ,
		_w10170_,
		_w10171_,
		_w10172_
	);
	LUT4 #(
		.INIT('h1441)
	) name9640 (
		ld_pad,
		\u0_w_reg[0][6]/P0001 ,
		_w10170_,
		_w10171_,
		_w10173_
	);
	LUT2 #(
		.INIT('h1)
	) name9641 (
		_w10127_,
		_w10173_,
		_w10174_
	);
	LUT2 #(
		.INIT('h4)
	) name9642 (
		\key[45]_pad ,
		ld_pad,
		_w10175_
	);
	LUT3 #(
		.INIT('h20)
	) name9643 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10176_
	);
	LUT4 #(
		.INIT('hf7a7)
	) name9644 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10177_
	);
	LUT4 #(
		.INIT('h4051)
	) name9645 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w9329_,
		_w10177_,
		_w10178_
	);
	LUT3 #(
		.INIT('h54)
	) name9646 (
		\u0_w_reg[3][7]/P0001 ,
		_w9319_,
		_w9393_,
		_w10179_
	);
	LUT2 #(
		.INIT('h4)
	) name9647 (
		_w9312_,
		_w9323_,
		_w10180_
	);
	LUT3 #(
		.INIT('h01)
	) name9648 (
		_w9260_,
		_w9308_,
		_w9401_,
		_w10181_
	);
	LUT4 #(
		.INIT('h0100)
	) name9649 (
		_w10178_,
		_w10179_,
		_w10180_,
		_w10181_,
		_w10182_
	);
	LUT3 #(
		.INIT('h54)
	) name9650 (
		\u0_w_reg[3][5]/P0001 ,
		_w9382_,
		_w9816_,
		_w10183_
	);
	LUT4 #(
		.INIT('h45cf)
	) name9651 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w9255_,
		_w9346_,
		_w10184_
	);
	LUT2 #(
		.INIT('h4)
	) name9652 (
		_w10183_,
		_w10184_,
		_w10185_
	);
	LUT4 #(
		.INIT('h8002)
	) name9653 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10186_
	);
	LUT4 #(
		.INIT('h0007)
	) name9654 (
		_w9286_,
		_w9376_,
		_w9828_,
		_w10186_,
		_w10187_
	);
	LUT3 #(
		.INIT('h0b)
	) name9655 (
		\u0_w_reg[3][2]/P0001 ,
		_w9322_,
		_w9378_,
		_w10188_
	);
	LUT4 #(
		.INIT('he400)
	) name9656 (
		\u0_w_reg[3][2]/P0001 ,
		_w10040_,
		_w10187_,
		_w10188_,
		_w10189_
	);
	LUT4 #(
		.INIT('hd800)
	) name9657 (
		\u0_w_reg[3][1]/P0001 ,
		_w10182_,
		_w10185_,
		_w10189_,
		_w10190_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name9658 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w9259_,
		_w10191_
	);
	LUT4 #(
		.INIT('h0200)
	) name9659 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10192_
	);
	LUT4 #(
		.INIT('h002a)
	) name9660 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		_w9346_,
		_w10192_,
		_w10193_
	);
	LUT2 #(
		.INIT('h8)
	) name9661 (
		_w10191_,
		_w10193_,
		_w10194_
	);
	LUT3 #(
		.INIT('ha8)
	) name9662 (
		\u0_w_reg[3][2]/P0001 ,
		_w9370_,
		_w9400_,
		_w10195_
	);
	LUT3 #(
		.INIT('h07)
	) name9663 (
		\u0_w_reg[3][6]/P0001 ,
		_w9279_,
		_w9411_,
		_w10196_
	);
	LUT4 #(
		.INIT('h0040)
	) name9664 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10197_
	);
	LUT4 #(
		.INIT('h0045)
	) name9665 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		_w9257_,
		_w10197_,
		_w10198_
	);
	LUT3 #(
		.INIT('h40)
	) name9666 (
		_w10195_,
		_w10196_,
		_w10198_,
		_w10199_
	);
	LUT3 #(
		.INIT('h02)
	) name9667 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10200_
	);
	LUT4 #(
		.INIT('h2023)
	) name9668 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w10201_
	);
	LUT3 #(
		.INIT('ha8)
	) name9669 (
		\u0_w_reg[3][1]/P0001 ,
		_w10200_,
		_w10201_,
		_w10202_
	);
	LUT4 #(
		.INIT('h5545)
	) name9670 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10203_
	);
	LUT3 #(
		.INIT('h10)
	) name9671 (
		_w9379_,
		_w9411_,
		_w10203_,
		_w10204_
	);
	LUT3 #(
		.INIT('h2a)
	) name9672 (
		\u0_w_reg[3][2]/P0001 ,
		_w9285_,
		_w9287_,
		_w10205_
	);
	LUT4 #(
		.INIT('h8acf)
	) name9673 (
		_w9280_,
		_w10202_,
		_w10204_,
		_w10205_,
		_w10206_
	);
	LUT4 #(
		.INIT('h0777)
	) name9674 (
		_w9274_,
		_w9307_,
		_w9297_,
		_w9332_,
		_w10207_
	);
	LUT4 #(
		.INIT('h5400)
	) name9675 (
		_w10206_,
		_w10194_,
		_w10199_,
		_w10207_,
		_w10208_
	);
	LUT4 #(
		.INIT('h0080)
	) name9676 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w10209_
	);
	LUT3 #(
		.INIT('h10)
	) name9677 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10210_
	);
	LUT3 #(
		.INIT('h6b)
	) name9678 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10211_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name9679 (
		\u0_w_reg[3][2]/P0001 ,
		_w9375_,
		_w10209_,
		_w10211_,
		_w10212_
	);
	LUT3 #(
		.INIT('h07)
	) name9680 (
		_w9274_,
		_w9307_,
		_w9315_,
		_w10213_
	);
	LUT4 #(
		.INIT('h153f)
	) name9681 (
		_w9274_,
		_w9303_,
		_w9369_,
		_w9411_,
		_w10214_
	);
	LUT4 #(
		.INIT('h4555)
	) name9682 (
		\u0_w_reg[3][1]/P0001 ,
		_w10212_,
		_w10213_,
		_w10214_,
		_w10215_
	);
	LUT4 #(
		.INIT('h23af)
	) name9683 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w9322_,
		_w9378_,
		_w10216_
	);
	LUT2 #(
		.INIT('h2)
	) name9684 (
		\u0_w_reg[3][1]/P0001 ,
		_w10216_,
		_w10217_
	);
	LUT4 #(
		.INIT('h5450)
	) name9685 (
		\u0_w_reg[3][2]/P0001 ,
		_w9259_,
		_w9308_,
		_w9366_,
		_w10218_
	);
	LUT2 #(
		.INIT('h8)
	) name9686 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		_w10219_
	);
	LUT3 #(
		.INIT('h80)
	) name9687 (
		\u0_w_reg[3][4]/P0001 ,
		_w9251_,
		_w10219_,
		_w10220_
	);
	LUT2 #(
		.INIT('h8)
	) name9688 (
		_w9272_,
		_w10209_,
		_w10221_
	);
	LUT3 #(
		.INIT('h01)
	) name9689 (
		_w10218_,
		_w10220_,
		_w10221_,
		_w10222_
	);
	LUT3 #(
		.INIT('h10)
	) name9690 (
		_w10215_,
		_w10217_,
		_w10222_,
		_w10223_
	);
	LUT4 #(
		.INIT('hd800)
	) name9691 (
		\u0_w_reg[3][0]/P0001 ,
		_w10208_,
		_w10190_,
		_w10223_,
		_w10224_
	);
	LUT2 #(
		.INIT('h9)
	) name9692 (
		\u0_w_reg[1][13]/P0001 ,
		\u0_w_reg[2][13]/P0001 ,
		_w10225_
	);
	LUT3 #(
		.INIT('h69)
	) name9693 (
		\u0_w_reg[0][13]/P0001 ,
		_w10224_,
		_w10225_,
		_w10226_
	);
	LUT4 #(
		.INIT('h1441)
	) name9694 (
		ld_pad,
		\u0_w_reg[0][13]/P0001 ,
		_w10224_,
		_w10225_,
		_w10227_
	);
	LUT2 #(
		.INIT('h1)
	) name9695 (
		_w10175_,
		_w10227_,
		_w10228_
	);
	LUT4 #(
		.INIT('hf5c5)
	) name9696 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10229_
	);
	LUT2 #(
		.INIT('h2)
	) name9697 (
		_w9830_,
		_w10229_,
		_w10230_
	);
	LUT2 #(
		.INIT('h8)
	) name9698 (
		_w9268_,
		_w9818_,
		_w10231_
	);
	LUT4 #(
		.INIT('h002a)
	) name9699 (
		\u0_w_reg[3][1]/P0001 ,
		_w9307_,
		_w9375_,
		_w9842_,
		_w10232_
	);
	LUT3 #(
		.INIT('h10)
	) name9700 (
		_w10231_,
		_w10230_,
		_w10232_,
		_w10233_
	);
	LUT2 #(
		.INIT('h8)
	) name9701 (
		_w9289_,
		_w9294_,
		_w10234_
	);
	LUT4 #(
		.INIT('h0002)
	) name9702 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10235_
	);
	LUT3 #(
		.INIT('h01)
	) name9703 (
		\u0_w_reg[3][1]/P0001 ,
		_w10037_,
		_w10235_,
		_w10236_
	);
	LUT2 #(
		.INIT('h4)
	) name9704 (
		_w10234_,
		_w10236_,
		_w10237_
	);
	LUT2 #(
		.INIT('h8)
	) name9705 (
		\u0_w_reg[3][4]/P0001 ,
		_w9302_,
		_w10238_
	);
	LUT4 #(
		.INIT('h0100)
	) name9706 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10239_
	);
	LUT4 #(
		.INIT('h0015)
	) name9707 (
		\u0_w_reg[3][0]/P0001 ,
		_w9274_,
		_w9411_,
		_w10239_,
		_w10240_
	);
	LUT4 #(
		.INIT('h8000)
	) name9708 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10241_
	);
	LUT4 #(
		.INIT('h7ffe)
	) name9709 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10242_
	);
	LUT2 #(
		.INIT('h2)
	) name9710 (
		_w9289_,
		_w10242_,
		_w10243_
	);
	LUT4 #(
		.INIT('h3fbb)
	) name9711 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10244_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9712 (
		_w9272_,
		_w9303_,
		_w10209_,
		_w10244_,
		_w10245_
	);
	LUT4 #(
		.INIT('h1000)
	) name9713 (
		_w10243_,
		_w10238_,
		_w10240_,
		_w10245_,
		_w10246_
	);
	LUT3 #(
		.INIT('he0)
	) name9714 (
		_w10233_,
		_w10237_,
		_w10246_,
		_w10247_
	);
	LUT4 #(
		.INIT('h7f5f)
	) name9715 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10248_
	);
	LUT4 #(
		.INIT('hd8dd)
	) name9716 (
		\u0_w_reg[3][2]/P0001 ,
		_w9266_,
		_w9336_,
		_w10248_,
		_w10249_
	);
	LUT3 #(
		.INIT('h04)
	) name9717 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10250_
	);
	LUT2 #(
		.INIT('h4)
	) name9718 (
		_w9317_,
		_w10250_,
		_w10251_
	);
	LUT3 #(
		.INIT('h01)
	) name9719 (
		\u0_w_reg[3][1]/P0001 ,
		_w9412_,
		_w10197_,
		_w10252_
	);
	LUT3 #(
		.INIT('h10)
	) name9720 (
		_w10249_,
		_w10251_,
		_w10252_,
		_w10253_
	);
	LUT3 #(
		.INIT('had)
	) name9721 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w10254_
	);
	LUT3 #(
		.INIT('hf6)
	) name9722 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10255_
	);
	LUT3 #(
		.INIT('h2a)
	) name9723 (
		\u0_w_reg[3][2]/P0001 ,
		_w10254_,
		_w10255_,
		_w10256_
	);
	LUT2 #(
		.INIT('h8)
	) name9724 (
		_w9262_,
		_w9286_,
		_w10257_
	);
	LUT3 #(
		.INIT('h2a)
	) name9725 (
		\u0_w_reg[3][1]/P0001 ,
		_w9303_,
		_w10210_,
		_w10258_
	);
	LUT3 #(
		.INIT('h10)
	) name9726 (
		_w10256_,
		_w10257_,
		_w10258_,
		_w10259_
	);
	LUT4 #(
		.INIT('h0040)
	) name9727 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10260_
	);
	LUT4 #(
		.INIT('h002a)
	) name9728 (
		\u0_w_reg[3][0]/P0001 ,
		_w9289_,
		_w9400_,
		_w10260_,
		_w10261_
	);
	LUT3 #(
		.INIT('ha8)
	) name9729 (
		\u0_w_reg[3][4]/P0001 ,
		_w9316_,
		_w9304_,
		_w10262_
	);
	LUT4 #(
		.INIT('ha7f7)
	) name9730 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10263_
	);
	LUT2 #(
		.INIT('h2)
	) name9731 (
		_w9268_,
		_w10263_,
		_w10264_
	);
	LUT3 #(
		.INIT('h10)
	) name9732 (
		_w10262_,
		_w10264_,
		_w10261_,
		_w10265_
	);
	LUT3 #(
		.INIT('he0)
	) name9733 (
		_w10253_,
		_w10259_,
		_w10265_,
		_w10266_
	);
	LUT4 #(
		.INIT('hadfb)
	) name9734 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10267_
	);
	LUT2 #(
		.INIT('h1)
	) name9735 (
		\u0_w_reg[3][3]/P0001 ,
		_w10267_,
		_w10268_
	);
	LUT3 #(
		.INIT('h02)
	) name9736 (
		\u0_w_reg[3][2]/P0001 ,
		_w9353_,
		_w9411_,
		_w10269_
	);
	LUT4 #(
		.INIT('h0010)
	) name9737 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10270_
	);
	LUT4 #(
		.INIT('hbfef)
	) name9738 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10271_
	);
	LUT4 #(
		.INIT('hb7e3)
	) name9739 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10272_
	);
	LUT4 #(
		.INIT('h88a8)
	) name9740 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w10272_,
		_w10273_
	);
	LUT3 #(
		.INIT('hb0)
	) name9741 (
		_w10268_,
		_w10269_,
		_w10273_,
		_w10274_
	);
	LUT2 #(
		.INIT('h4)
	) name9742 (
		\u0_w_reg[3][2]/P0001 ,
		_w10060_,
		_w10275_
	);
	LUT3 #(
		.INIT('h51)
	) name9743 (
		_w9279_,
		_w9303_,
		_w10244_,
		_w10276_
	);
	LUT3 #(
		.INIT('h45)
	) name9744 (
		\u0_w_reg[3][1]/P0001 ,
		_w10275_,
		_w10276_,
		_w10277_
	);
	LUT4 #(
		.INIT('hf080)
	) name9745 (
		_w9262_,
		_w9286_,
		_w9344_,
		_w9401_,
		_w10278_
	);
	LUT2 #(
		.INIT('h8)
	) name9746 (
		_w9830_,
		_w10070_,
		_w10279_
	);
	LUT4 #(
		.INIT('h135f)
	) name9747 (
		_w9344_,
		_w9365_,
		_w9392_,
		_w10047_,
		_w10280_
	);
	LUT4 #(
		.INIT('h0032)
	) name9748 (
		\u0_w_reg[3][3]/P0001 ,
		_w10279_,
		_w10280_,
		_w10278_,
		_w10281_
	);
	LUT3 #(
		.INIT('h10)
	) name9749 (
		_w10274_,
		_w10277_,
		_w10281_,
		_w10282_
	);
	LUT4 #(
		.INIT('ha955)
	) name9750 (
		\u0_w_reg[0][15]/P0001 ,
		_w10247_,
		_w10266_,
		_w10282_,
		_w10283_
	);
	LUT3 #(
		.INIT('h96)
	) name9751 (
		\u0_w_reg[1][15]/P0001 ,
		\u0_w_reg[2][15]/P0001 ,
		_w10283_,
		_w10284_
	);
	LUT4 #(
		.INIT('h4114)
	) name9752 (
		ld_pad,
		\u0_w_reg[1][15]/P0001 ,
		\u0_w_reg[2][15]/P0001 ,
		_w10283_,
		_w10285_
	);
	LUT2 #(
		.INIT('h8)
	) name9753 (
		\key[47]_pad ,
		ld_pad,
		_w10286_
	);
	LUT2 #(
		.INIT('he)
	) name9754 (
		_w10285_,
		_w10286_,
		_w10287_
	);
	LUT2 #(
		.INIT('h4)
	) name9755 (
		\key[40]_pad ,
		ld_pad,
		_w10288_
	);
	LUT2 #(
		.INIT('h1)
	) name9756 (
		\u0_w_reg[3][3]/P0001 ,
		_w10271_,
		_w10289_
	);
	LUT2 #(
		.INIT('h2)
	) name9757 (
		_w9290_,
		_w9297_,
		_w10290_
	);
	LUT3 #(
		.INIT('h45)
	) name9758 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		_w9370_,
		_w10291_
	);
	LUT3 #(
		.INIT('h10)
	) name9759 (
		_w10289_,
		_w10290_,
		_w10291_,
		_w10292_
	);
	LUT3 #(
		.INIT('h80)
	) name9760 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10293_
	);
	LUT3 #(
		.INIT('ha8)
	) name9761 (
		\u0_w_reg[3][3]/P0001 ,
		_w9316_,
		_w10293_,
		_w10294_
	);
	LUT4 #(
		.INIT('haaa8)
	) name9762 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10295_
	);
	LUT4 #(
		.INIT('h0100)
	) name9763 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10296_
	);
	LUT3 #(
		.INIT('h10)
	) name9764 (
		_w9828_,
		_w10296_,
		_w10295_,
		_w10297_
	);
	LUT2 #(
		.INIT('h4)
	) name9765 (
		_w10294_,
		_w10297_,
		_w10298_
	);
	LUT4 #(
		.INIT('h000b)
	) name9766 (
		\u0_w_reg[3][3]/P0001 ,
		_w9322_,
		_w9324_,
		_w10051_,
		_w10299_
	);
	LUT3 #(
		.INIT('hb9)
	) name9767 (
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10300_
	);
	LUT3 #(
		.INIT('h51)
	) name9768 (
		\u0_w_reg[3][0]/P0001 ,
		_w9381_,
		_w10300_,
		_w10301_
	);
	LUT3 #(
		.INIT('he0)
	) name9769 (
		\u0_w_reg[3][2]/P0001 ,
		_w10299_,
		_w10301_,
		_w10302_
	);
	LUT3 #(
		.INIT('he0)
	) name9770 (
		_w10292_,
		_w10298_,
		_w10302_,
		_w10303_
	);
	LUT4 #(
		.INIT('ha888)
	) name9771 (
		\u0_w_reg[3][4]/P0001 ,
		_w9316_,
		_w9303_,
		_w10210_,
		_w10304_
	);
	LUT4 #(
		.INIT('h3ffa)
	) name9772 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10305_
	);
	LUT2 #(
		.INIT('h2)
	) name9773 (
		_w9394_,
		_w10305_,
		_w10306_
	);
	LUT4 #(
		.INIT('h5551)
	) name9774 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		_w10307_
	);
	LUT3 #(
		.INIT('h10)
	) name9775 (
		_w9823_,
		_w10192_,
		_w10307_,
		_w10308_
	);
	LUT4 #(
		.INIT('h0002)
	) name9776 (
		\u0_w_reg[3][1]/P0001 ,
		_w9327_,
		_w9302_,
		_w10047_,
		_w10309_
	);
	LUT4 #(
		.INIT('h00ef)
	) name9777 (
		_w10306_,
		_w10304_,
		_w10308_,
		_w10309_,
		_w10310_
	);
	LUT4 #(
		.INIT('h0004)
	) name9778 (
		_w9366_,
		_w9844_,
		_w10241_,
		_w10260_,
		_w10311_
	);
	LUT3 #(
		.INIT('h02)
	) name9779 (
		\u0_w_reg[3][2]/P0001 ,
		_w9386_,
		_w10037_,
		_w10312_
	);
	LUT4 #(
		.INIT('h0222)
	) name9780 (
		\u0_w_reg[3][0]/P0001 ,
		_w9251_,
		_w9329_,
		_w9426_,
		_w10313_
	);
	LUT4 #(
		.INIT('hec00)
	) name9781 (
		_w10191_,
		_w10311_,
		_w10312_,
		_w10313_,
		_w10314_
	);
	LUT2 #(
		.INIT('h4)
	) name9782 (
		_w10310_,
		_w10314_,
		_w10315_
	);
	LUT2 #(
		.INIT('h4)
	) name9783 (
		\u0_w_reg[3][3]/P0001 ,
		_w9831_,
		_w10316_
	);
	LUT3 #(
		.INIT('h15)
	) name9784 (
		_w9257_,
		_w9286_,
		_w9376_,
		_w10317_
	);
	LUT3 #(
		.INIT('h8a)
	) name9785 (
		\u0_w_reg[3][2]/P0001 ,
		_w10316_,
		_w10317_,
		_w10318_
	);
	LUT3 #(
		.INIT('h8a)
	) name9786 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w9378_,
		_w10319_
	);
	LUT4 #(
		.INIT('h23af)
	) name9787 (
		\u0_w_reg[3][2]/P0001 ,
		_w9259_,
		_w9279_,
		_w9366_,
		_w10320_
	);
	LUT2 #(
		.INIT('h8)
	) name9788 (
		_w10319_,
		_w10320_,
		_w10321_
	);
	LUT3 #(
		.INIT('h07)
	) name9789 (
		_w9259_,
		_w9281_,
		_w9319_,
		_w10322_
	);
	LUT4 #(
		.INIT('hff4f)
	) name9790 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10323_
	);
	LUT2 #(
		.INIT('h1)
	) name9791 (
		\u0_w_reg[3][3]/P0001 ,
		_w10323_,
		_w10324_
	);
	LUT3 #(
		.INIT('h45)
	) name9792 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w9823_,
		_w10325_
	);
	LUT4 #(
		.INIT('h7077)
	) name9793 (
		_w9410_,
		_w10322_,
		_w10324_,
		_w10325_,
		_w10326_
	);
	LUT3 #(
		.INIT('h15)
	) name9794 (
		\u0_w_reg[3][1]/P0001 ,
		_w9830_,
		_w9831_,
		_w10327_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name9795 (
		_w10318_,
		_w10321_,
		_w10326_,
		_w10327_,
		_w10328_
	);
	LUT2 #(
		.INIT('h8)
	) name9796 (
		_w9274_,
		_w9845_,
		_w10329_
	);
	LUT4 #(
		.INIT('h1110)
	) name9797 (
		_w10328_,
		_w10329_,
		_w10303_,
		_w10315_,
		_w10330_
	);
	LUT2 #(
		.INIT('h9)
	) name9798 (
		\u0_w_reg[1][8]/P0001 ,
		\u0_w_reg[2][8]/P0001 ,
		_w10331_
	);
	LUT3 #(
		.INIT('h69)
	) name9799 (
		\u0_w_reg[0][8]/P0001 ,
		_w10330_,
		_w10331_,
		_w10332_
	);
	LUT4 #(
		.INIT('h1441)
	) name9800 (
		ld_pad,
		\u0_w_reg[0][8]/P0001 ,
		_w10330_,
		_w10331_,
		_w10333_
	);
	LUT2 #(
		.INIT('h1)
	) name9801 (
		_w10288_,
		_w10333_,
		_w10334_
	);
	LUT4 #(
		.INIT('h4000)
	) name9802 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10335_
	);
	LUT3 #(
		.INIT('ha8)
	) name9803 (
		\u0_w_reg[3][18]/P0001 ,
		_w8694_,
		_w10335_,
		_w10336_
	);
	LUT4 #(
		.INIT('h0800)
	) name9804 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w10337_
	);
	LUT4 #(
		.INIT('h5554)
	) name9805 (
		\u0_w_reg[3][18]/P0001 ,
		_w8688_,
		_w9533_,
		_w10337_,
		_w10338_
	);
	LUT4 #(
		.INIT('h0002)
	) name9806 (
		\u0_w_reg[3][17]/P0001 ,
		_w8737_,
		_w8738_,
		_w8666_,
		_w10339_
	);
	LUT3 #(
		.INIT('h10)
	) name9807 (
		_w10338_,
		_w10336_,
		_w10339_,
		_w10340_
	);
	LUT2 #(
		.INIT('h8)
	) name9808 (
		_w8772_,
		_w9592_,
		_w10341_
	);
	LUT4 #(
		.INIT('h8caf)
	) name9809 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w8698_,
		_w9120_,
		_w10342_
	);
	LUT3 #(
		.INIT('h15)
	) name9810 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		_w9145_,
		_w10343_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name9811 (
		\u0_w_reg[3][21]/P0001 ,
		_w8656_,
		_w8732_,
		_w8722_,
		_w10344_
	);
	LUT4 #(
		.INIT('h4000)
	) name9812 (
		_w10341_,
		_w10343_,
		_w10344_,
		_w10342_,
		_w10345_
	);
	LUT2 #(
		.INIT('h8)
	) name9813 (
		_w8729_,
		_w9114_,
		_w10346_
	);
	LUT3 #(
		.INIT('h13)
	) name9814 (
		_w8689_,
		_w8751_,
		_w8770_,
		_w10347_
	);
	LUT4 #(
		.INIT('hffa8)
	) name9815 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10348_
	);
	LUT2 #(
		.INIT('h2)
	) name9816 (
		_w8732_,
		_w10348_,
		_w10349_
	);
	LUT4 #(
		.INIT('h0100)
	) name9817 (
		_w9151_,
		_w10346_,
		_w10349_,
		_w10347_,
		_w10350_
	);
	LUT4 #(
		.INIT('h0155)
	) name9818 (
		\u0_w_reg[3][16]/P0001 ,
		_w10340_,
		_w10345_,
		_w10350_,
		_w10351_
	);
	LUT3 #(
		.INIT('h80)
	) name9819 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10352_
	);
	LUT4 #(
		.INIT('hcedf)
	) name9820 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10353_
	);
	LUT3 #(
		.INIT('h8a)
	) name9821 (
		\u0_w_reg[3][18]/P0001 ,
		_w10352_,
		_w10353_,
		_w10354_
	);
	LUT3 #(
		.INIT('ha2)
	) name9822 (
		\u0_w_reg[3][17]/P0001 ,
		_w9532_,
		_w10354_,
		_w10355_
	);
	LUT3 #(
		.INIT('hc5)
	) name9823 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10356_
	);
	LUT2 #(
		.INIT('h2)
	) name9824 (
		_w8722_,
		_w10356_,
		_w10357_
	);
	LUT4 #(
		.INIT('h0400)
	) name9825 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10358_
	);
	LUT3 #(
		.INIT('h07)
	) name9826 (
		_w8720_,
		_w9158_,
		_w10358_,
		_w10359_
	);
	LUT3 #(
		.INIT('h45)
	) name9827 (
		\u0_w_reg[3][17]/P0001 ,
		_w10357_,
		_w10359_,
		_w10360_
	);
	LUT4 #(
		.INIT('hf7bf)
	) name9828 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10361_
	);
	LUT2 #(
		.INIT('h1)
	) name9829 (
		\u0_w_reg[3][18]/P0001 ,
		_w10361_,
		_w10362_
	);
	LUT2 #(
		.INIT('h2)
	) name9830 (
		_w9164_,
		_w9541_,
		_w10363_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name9831 (
		_w8674_,
		_w8677_,
		_w8689_,
		_w8770_,
		_w10364_
	);
	LUT3 #(
		.INIT('h10)
	) name9832 (
		_w10362_,
		_w10363_,
		_w10364_,
		_w10365_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9833 (
		\u0_w_reg[3][16]/P0001 ,
		_w10355_,
		_w10360_,
		_w10365_,
		_w10366_
	);
	LUT4 #(
		.INIT('h0007)
	) name9834 (
		_w8654_,
		_w8681_,
		_w9443_,
		_w9623_,
		_w10367_
	);
	LUT3 #(
		.INIT('h9f)
	) name9835 (
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w8723_,
		_w10368_
	);
	LUT4 #(
		.INIT('h0155)
	) name9836 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		_w10367_,
		_w10368_,
		_w10369_
	);
	LUT3 #(
		.INIT('h54)
	) name9837 (
		_w8707_,
		_w8720_,
		_w8709_,
		_w10370_
	);
	LUT2 #(
		.INIT('h1)
	) name9838 (
		_w8666_,
		_w9484_,
		_w10371_
	);
	LUT3 #(
		.INIT('h8a)
	) name9839 (
		_w9504_,
		_w10370_,
		_w10371_,
		_w10372_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name9840 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10373_
	);
	LUT4 #(
		.INIT('hbf15)
	) name9841 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		_w8676_,
		_w10373_,
		_w10374_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name9842 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10375_
	);
	LUT4 #(
		.INIT('h7cfa)
	) name9843 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10376_
	);
	LUT4 #(
		.INIT('hf531)
	) name9844 (
		_w8689_,
		_w9163_,
		_w10375_,
		_w10376_,
		_w10377_
	);
	LUT3 #(
		.INIT('hd0)
	) name9845 (
		_w9541_,
		_w10374_,
		_w10377_,
		_w10378_
	);
	LUT3 #(
		.INIT('h10)
	) name9846 (
		_w10372_,
		_w10369_,
		_w10378_,
		_w10379_
	);
	LUT4 #(
		.INIT('h5655)
	) name9847 (
		\u0_w_reg[0][25]/P0001 ,
		_w10366_,
		_w10351_,
		_w10379_,
		_w10380_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name9848 (
		\key[121]_pad ,
		ld_pad,
		\u0_r0_out_reg[25]/P0001 ,
		_w10380_,
		_w10381_
	);
	LUT2 #(
		.INIT('h9)
	) name9849 (
		\u0_r0_out_reg[25]/P0001 ,
		\u0_w_reg[1][25]/P0001 ,
		_w10382_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9850 (
		\key[89]_pad ,
		ld_pad,
		_w10380_,
		_w10382_,
		_w10383_
	);
	LUT3 #(
		.INIT('h69)
	) name9851 (
		\u0_r0_out_reg[25]/P0001 ,
		\u0_w_reg[1][25]/P0001 ,
		\u0_w_reg[2][25]/P0001 ,
		_w10384_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9852 (
		\key[57]_pad ,
		ld_pad,
		_w10380_,
		_w10384_,
		_w10385_
	);
	LUT4 #(
		.INIT('h1441)
	) name9853 (
		ld_pad,
		\u0_w_reg[3][25]/P0001 ,
		_w10380_,
		_w10384_,
		_w10386_
	);
	LUT2 #(
		.INIT('h8)
	) name9854 (
		\key[25]_pad ,
		ld_pad,
		_w10387_
	);
	LUT2 #(
		.INIT('he)
	) name9855 (
		_w10386_,
		_w10387_,
		_w10388_
	);
	LUT4 #(
		.INIT('h0020)
	) name9856 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10389_
	);
	LUT3 #(
		.INIT('h54)
	) name9857 (
		\u0_w_reg[3][10]/P0001 ,
		_w8811_,
		_w10389_,
		_w10390_
	);
	LUT3 #(
		.INIT('h07)
	) name9858 (
		_w8937_,
		_w9915_,
		_w9949_,
		_w10391_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9859 (
		\u0_w_reg[3][9]/P0001 ,
		_w10098_,
		_w10390_,
		_w10391_,
		_w10392_
	);
	LUT3 #(
		.INIT('h80)
	) name9860 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w9966_,
		_w10393_
	);
	LUT4 #(
		.INIT('h0015)
	) name9861 (
		\u0_w_reg[3][8]/P0001 ,
		_w8893_,
		_w8894_,
		_w8967_,
		_w10394_
	);
	LUT4 #(
		.INIT('h1101)
	) name9862 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10395_
	);
	LUT4 #(
		.INIT('h0777)
	) name9863 (
		_w8851_,
		_w8889_,
		_w9887_,
		_w10395_,
		_w10396_
	);
	LUT3 #(
		.INIT('h40)
	) name9864 (
		_w10393_,
		_w10394_,
		_w10396_,
		_w10397_
	);
	LUT4 #(
		.INIT('h0013)
	) name9865 (
		_w8854_,
		_w8852_,
		_w8914_,
		_w9890_,
		_w10398_
	);
	LUT4 #(
		.INIT('h5150)
	) name9866 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w8805_,
		_w9966_,
		_w10399_
	);
	LUT3 #(
		.INIT('h0e)
	) name9867 (
		\u0_w_reg[3][9]/P0001 ,
		_w10398_,
		_w10399_,
		_w10400_
	);
	LUT3 #(
		.INIT('h40)
	) name9868 (
		_w10392_,
		_w10397_,
		_w10400_,
		_w10401_
	);
	LUT4 #(
		.INIT('h4151)
	) name9869 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10402_
	);
	LUT3 #(
		.INIT('ha8)
	) name9870 (
		\u0_w_reg[3][12]/P0001 ,
		_w8911_,
		_w10402_,
		_w10403_
	);
	LUT4 #(
		.INIT('h0010)
	) name9871 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10404_
	);
	LUT3 #(
		.INIT('h01)
	) name9872 (
		\u0_w_reg[3][9]/P0001 ,
		_w9916_,
		_w10404_,
		_w10405_
	);
	LUT4 #(
		.INIT('h0040)
	) name9873 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10406_
	);
	LUT3 #(
		.INIT('h07)
	) name9874 (
		_w8851_,
		_w8925_,
		_w10406_,
		_w10407_
	);
	LUT3 #(
		.INIT('h40)
	) name9875 (
		_w10403_,
		_w10405_,
		_w10407_,
		_w10408_
	);
	LUT3 #(
		.INIT('had)
	) name9876 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w10409_
	);
	LUT3 #(
		.INIT('hf6)
	) name9877 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10410_
	);
	LUT3 #(
		.INIT('h2a)
	) name9878 (
		\u0_w_reg[3][10]/P0001 ,
		_w10409_,
		_w10410_,
		_w10411_
	);
	LUT3 #(
		.INIT('h2a)
	) name9879 (
		\u0_w_reg[3][9]/P0001 ,
		_w8793_,
		_w8943_,
		_w10412_
	);
	LUT2 #(
		.INIT('h4)
	) name9880 (
		\u0_w_reg[3][14]/P0001 ,
		_w9873_,
		_w10413_
	);
	LUT3 #(
		.INIT('h04)
	) name9881 (
		_w10411_,
		_w10412_,
		_w10413_,
		_w10414_
	);
	LUT4 #(
		.INIT('ha7f7)
	) name9882 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10415_
	);
	LUT2 #(
		.INIT('h2)
	) name9883 (
		_w8937_,
		_w10415_,
		_w10416_
	);
	LUT4 #(
		.INIT('h002a)
	) name9884 (
		\u0_w_reg[3][8]/P0001 ,
		_w8804_,
		_w8836_,
		_w9894_,
		_w10417_
	);
	LUT4 #(
		.INIT('h15bf)
	) name9885 (
		\u0_w_reg[3][12]/P0001 ,
		_w8793_,
		_w8854_,
		_w10404_,
		_w10418_
	);
	LUT3 #(
		.INIT('h40)
	) name9886 (
		_w10416_,
		_w10417_,
		_w10418_,
		_w10419_
	);
	LUT3 #(
		.INIT('he0)
	) name9887 (
		_w10408_,
		_w10414_,
		_w10419_,
		_w10420_
	);
	LUT4 #(
		.INIT('hadfb)
	) name9888 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10421_
	);
	LUT2 #(
		.INIT('h1)
	) name9889 (
		\u0_w_reg[3][11]/P0001 ,
		_w10421_,
		_w10422_
	);
	LUT3 #(
		.INIT('h02)
	) name9890 (
		\u0_w_reg[3][10]/P0001 ,
		_w8800_,
		_w8860_,
		_w10423_
	);
	LUT4 #(
		.INIT('hbfe3)
	) name9891 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10424_
	);
	LUT4 #(
		.INIT('h0501)
	) name9892 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w8874_,
		_w10424_,
		_w10425_
	);
	LUT4 #(
		.INIT('h2022)
	) name9893 (
		\u0_w_reg[3][9]/P0001 ,
		_w10425_,
		_w10422_,
		_w10423_,
		_w10426_
	);
	LUT3 #(
		.INIT('h10)
	) name9894 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10427_
	);
	LUT2 #(
		.INIT('h8)
	) name9895 (
		_w8878_,
		_w10427_,
		_w10428_
	);
	LUT3 #(
		.INIT('h15)
	) name9896 (
		_w8919_,
		_w9887_,
		_w10395_,
		_w10429_
	);
	LUT3 #(
		.INIT('h45)
	) name9897 (
		\u0_w_reg[3][9]/P0001 ,
		_w10428_,
		_w10429_,
		_w10430_
	);
	LUT4 #(
		.INIT('h67ef)
	) name9898 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		_w8784_,
		_w8910_,
		_w10431_
	);
	LUT4 #(
		.INIT('h0103)
	) name9899 (
		_w8793_,
		_w8840_,
		_w8941_,
		_w8943_,
		_w10432_
	);
	LUT4 #(
		.INIT('hfad8)
	) name9900 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w10431_,
		_w10432_,
		_w10433_
	);
	LUT3 #(
		.INIT('h10)
	) name9901 (
		_w10426_,
		_w10430_,
		_w10433_,
		_w10434_
	);
	LUT4 #(
		.INIT('ha955)
	) name9902 (
		\u0_w_reg[0][23]/P0001 ,
		_w10401_,
		_w10420_,
		_w10434_,
		_w10435_
	);
	LUT3 #(
		.INIT('h96)
	) name9903 (
		\u0_w_reg[1][23]/P0001 ,
		\u0_w_reg[2][23]/P0001 ,
		_w10435_,
		_w10436_
	);
	LUT4 #(
		.INIT('h4114)
	) name9904 (
		ld_pad,
		\u0_w_reg[1][23]/P0001 ,
		\u0_w_reg[2][23]/P0001 ,
		_w10435_,
		_w10437_
	);
	LUT2 #(
		.INIT('h8)
	) name9905 (
		\key[55]_pad ,
		ld_pad,
		_w10438_
	);
	LUT2 #(
		.INIT('he)
	) name9906 (
		_w10437_,
		_w10438_,
		_w10439_
	);
	LUT3 #(
		.INIT('hb8)
	) name9907 (
		\key[99]_pad ,
		ld_pad,
		_w9246_,
		_w10440_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name9908 (
		\key[67]_pad ,
		ld_pad,
		\u0_w_reg[1][3]/P0001 ,
		_w9246_,
		_w10441_
	);
	LUT4 #(
		.INIT('h1441)
	) name9909 (
		ld_pad,
		\u0_w_reg[3][3]/P0001 ,
		_w9246_,
		_w9247_,
		_w10442_
	);
	LUT2 #(
		.INIT('h8)
	) name9910 (
		\key[3]_pad ,
		ld_pad,
		_w10443_
	);
	LUT2 #(
		.INIT('he)
	) name9911 (
		_w10442_,
		_w10443_,
		_w10444_
	);
	LUT3 #(
		.INIT('hb8)
	) name9912 (
		\key[107]_pad ,
		ld_pad,
		_w9358_,
		_w10445_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name9913 (
		\key[75]_pad ,
		ld_pad,
		\u0_w_reg[1][11]/P0001 ,
		_w9358_,
		_w10446_
	);
	LUT4 #(
		.INIT('h1441)
	) name9914 (
		ld_pad,
		\u0_w_reg[3][11]/P0001 ,
		_w9358_,
		_w9359_,
		_w10447_
	);
	LUT2 #(
		.INIT('h8)
	) name9915 (
		\key[11]_pad ,
		ld_pad,
		_w10448_
	);
	LUT2 #(
		.INIT('he)
	) name9916 (
		_w10447_,
		_w10448_,
		_w10449_
	);
	LUT4 #(
		.INIT('haaa8)
	) name9917 (
		\u0_w_reg[3][10]/P0001 ,
		_w9915_,
		_w9946_,
		_w10427_,
		_w10450_
	);
	LUT3 #(
		.INIT('ha2)
	) name9918 (
		\u0_w_reg[3][9]/P0001 ,
		_w9972_,
		_w10450_,
		_w10451_
	);
	LUT4 #(
		.INIT('h0001)
	) name9919 (
		_w8842_,
		_w8964_,
		_w9935_,
		_w9949_,
		_w10452_
	);
	LUT2 #(
		.INIT('h1)
	) name9920 (
		\u0_w_reg[3][10]/P0001 ,
		_w10452_,
		_w10453_
	);
	LUT4 #(
		.INIT('h383b)
	) name9921 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		_w10454_
	);
	LUT4 #(
		.INIT('h0f01)
	) name9922 (
		_w8785_,
		_w8893_,
		_w8964_,
		_w10454_,
		_w10455_
	);
	LUT4 #(
		.INIT('h5510)
	) name9923 (
		\u0_w_reg[3][11]/P0001 ,
		_w8846_,
		_w8838_,
		_w9935_,
		_w10456_
	);
	LUT3 #(
		.INIT('h0e)
	) name9924 (
		\u0_w_reg[3][9]/P0001 ,
		_w10455_,
		_w10456_,
		_w10457_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9925 (
		\u0_w_reg[3][8]/P0001 ,
		_w10451_,
		_w10453_,
		_w10457_,
		_w10458_
	);
	LUT4 #(
		.INIT('h0803)
	) name9926 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w10459_
	);
	LUT4 #(
		.INIT('h5455)
	) name9927 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10460_
	);
	LUT4 #(
		.INIT('h4000)
	) name9928 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10461_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name9929 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10462_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name9930 (
		_w10459_,
		_w10460_,
		_w10461_,
		_w10462_,
		_w10463_
	);
	LUT4 #(
		.INIT('h0002)
	) name9931 (
		\u0_w_reg[3][9]/P0001 ,
		_w8800_,
		_w8818_,
		_w8840_,
		_w10464_
	);
	LUT2 #(
		.INIT('h4)
	) name9932 (
		_w10463_,
		_w10464_,
		_w10465_
	);
	LUT3 #(
		.INIT('h15)
	) name9933 (
		\u0_w_reg[3][9]/P0001 ,
		_w8838_,
		_w8854_,
		_w10466_
	);
	LUT3 #(
		.INIT('hbd)
	) name9934 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10467_
	);
	LUT3 #(
		.INIT('he3)
	) name9935 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10468_
	);
	LUT4 #(
		.INIT('hf351)
	) name9936 (
		_w8828_,
		_w8917_,
		_w10467_,
		_w10468_,
		_w10469_
	);
	LUT3 #(
		.INIT('h40)
	) name9937 (
		_w9938_,
		_w10466_,
		_w10469_,
		_w10470_
	);
	LUT2 #(
		.INIT('h8)
	) name9938 (
		_w8849_,
		_w8878_,
		_w10471_
	);
	LUT3 #(
		.INIT('h15)
	) name9939 (
		_w8885_,
		_w8893_,
		_w8894_,
		_w10472_
	);
	LUT4 #(
		.INIT('hffa8)
	) name9940 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10473_
	);
	LUT4 #(
		.INIT('hefcd)
	) name9941 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w8861_,
		_w10473_,
		_w10474_
	);
	LUT3 #(
		.INIT('h40)
	) name9942 (
		_w10471_,
		_w10472_,
		_w10474_,
		_w10475_
	);
	LUT4 #(
		.INIT('h0155)
	) name9943 (
		\u0_w_reg[3][8]/P0001 ,
		_w10465_,
		_w10470_,
		_w10475_,
		_w10476_
	);
	LUT4 #(
		.INIT('h000b)
	) name9944 (
		\u0_w_reg[3][11]/P0001 ,
		_w8805_,
		_w9890_,
		_w10389_,
		_w10477_
	);
	LUT4 #(
		.INIT('h153f)
	) name9945 (
		\u0_w_reg[3][11]/P0001 ,
		_w8810_,
		_w8811_,
		_w8850_,
		_w10478_
	);
	LUT4 #(
		.INIT('h0133)
	) name9946 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w10477_,
		_w10478_,
		_w10479_
	);
	LUT3 #(
		.INIT('h0b)
	) name9947 (
		\u0_w_reg[3][13]/P0001 ,
		_w8960_,
		_w9966_,
		_w10480_
	);
	LUT3 #(
		.INIT('h8c)
	) name9948 (
		_w10098_,
		_w10115_,
		_w10480_,
		_w10481_
	);
	LUT4 #(
		.INIT('hefec)
	) name9949 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10482_
	);
	LUT2 #(
		.INIT('h1)
	) name9950 (
		\u0_w_reg[3][14]/P0001 ,
		_w10482_,
		_w10483_
	);
	LUT3 #(
		.INIT('h01)
	) name9951 (
		_w8840_,
		_w9911_,
		_w9964_,
		_w10484_
	);
	LUT4 #(
		.INIT('hf7fd)
	) name9952 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10485_
	);
	LUT4 #(
		.INIT('h7cfa)
	) name9953 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10486_
	);
	LUT4 #(
		.INIT('hf531)
	) name9954 (
		_w8851_,
		_w8963_,
		_w10485_,
		_w10486_,
		_w10487_
	);
	LUT4 #(
		.INIT('h7500)
	) name9955 (
		_w8823_,
		_w10483_,
		_w10484_,
		_w10487_,
		_w10488_
	);
	LUT3 #(
		.INIT('h10)
	) name9956 (
		_w10481_,
		_w10479_,
		_w10488_,
		_w10489_
	);
	LUT4 #(
		.INIT('h5655)
	) name9957 (
		\u0_w_reg[0][17]/P0001 ,
		_w10476_,
		_w10458_,
		_w10489_,
		_w10490_
	);
	LUT2 #(
		.INIT('h9)
	) name9958 (
		\u0_w_reg[1][17]/P0001 ,
		\u0_w_reg[2][17]/P0001 ,
		_w10491_
	);
	LUT4 #(
		.INIT('hb88b)
	) name9959 (
		\key[49]_pad ,
		ld_pad,
		_w10490_,
		_w10491_,
		_w10492_
	);
	LUT2 #(
		.INIT('h2)
	) name9960 (
		\u0_w_reg[3][26]/P0001 ,
		_w9195_,
		_w10493_
	);
	LUT4 #(
		.INIT('h0105)
	) name9961 (
		\u0_w_reg[3][26]/P0001 ,
		_w9014_,
		_w9016_,
		_w9203_,
		_w10494_
	);
	LUT3 #(
		.INIT('h15)
	) name9962 (
		\u0_w_reg[3][25]/P0001 ,
		_w9026_,
		_w9194_,
		_w10495_
	);
	LUT4 #(
		.INIT('h153f)
	) name9963 (
		_w9066_,
		_w9068_,
		_w9035_,
		_w8996_,
		_w10496_
	);
	LUT4 #(
		.INIT('he000)
	) name9964 (
		_w10493_,
		_w10494_,
		_w10495_,
		_w10496_,
		_w10497_
	);
	LUT4 #(
		.INIT('h0800)
	) name9965 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w10498_
	);
	LUT3 #(
		.INIT('h10)
	) name9966 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10499_
	);
	LUT4 #(
		.INIT('h5554)
	) name9967 (
		\u0_w_reg[3][26]/P0001 ,
		_w8988_,
		_w10499_,
		_w10498_,
		_w10500_
	);
	LUT3 #(
		.INIT('ha8)
	) name9968 (
		\u0_w_reg[3][26]/P0001 ,
		_w8985_,
		_w10152_,
		_w10501_
	);
	LUT4 #(
		.INIT('h0002)
	) name9969 (
		\u0_w_reg[3][25]/P0001 ,
		_w9043_,
		_w9056_,
		_w9003_,
		_w10502_
	);
	LUT3 #(
		.INIT('h10)
	) name9970 (
		_w10501_,
		_w10500_,
		_w10502_,
		_w10503_
	);
	LUT4 #(
		.INIT('hffa8)
	) name9971 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10504_
	);
	LUT2 #(
		.INIT('h2)
	) name9972 (
		_w9068_,
		_w10504_,
		_w10505_
	);
	LUT3 #(
		.INIT('h15)
	) name9973 (
		_w9079_,
		_w9093_,
		_w9094_,
		_w10506_
	);
	LUT4 #(
		.INIT('habef)
	) name9974 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w9031_,
		_w9223_,
		_w10507_
	);
	LUT3 #(
		.INIT('h40)
	) name9975 (
		_w10505_,
		_w10506_,
		_w10507_,
		_w10508_
	);
	LUT4 #(
		.INIT('h0155)
	) name9976 (
		\u0_w_reg[3][24]/P0001 ,
		_w10497_,
		_w10503_,
		_w10508_,
		_w10509_
	);
	LUT4 #(
		.INIT('hcedf)
	) name9977 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10510_
	);
	LUT3 #(
		.INIT('h8a)
	) name9978 (
		\u0_w_reg[3][26]/P0001 ,
		_w10000_,
		_w10510_,
		_w10511_
	);
	LUT3 #(
		.INIT('ha2)
	) name9979 (
		\u0_w_reg[3][25]/P0001 ,
		_w10010_,
		_w10511_,
		_w10512_
	);
	LUT4 #(
		.INIT('h0001)
	) name9980 (
		_w9070_,
		_w9728_,
		_w9770_,
		_w9990_,
		_w10513_
	);
	LUT2 #(
		.INIT('h1)
	) name9981 (
		\u0_w_reg[3][26]/P0001 ,
		_w10513_,
		_w10514_
	);
	LUT4 #(
		.INIT('h383b)
	) name9982 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		_w10515_
	);
	LUT4 #(
		.INIT('h5501)
	) name9983 (
		_w9070_,
		_w8976_,
		_w9093_,
		_w10515_,
		_w10516_
	);
	LUT4 #(
		.INIT('h5504)
	) name9984 (
		\u0_w_reg[3][27]/P0001 ,
		_w8997_,
		_w9009_,
		_w9990_,
		_w10517_
	);
	LUT3 #(
		.INIT('h0e)
	) name9985 (
		\u0_w_reg[3][25]/P0001 ,
		_w10516_,
		_w10517_,
		_w10518_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9986 (
		\u0_w_reg[3][24]/P0001 ,
		_w10512_,
		_w10514_,
		_w10518_,
		_w10519_
	);
	LUT4 #(
		.INIT('h0007)
	) name9987 (
		_w8977_,
		_w9053_,
		_w9731_,
		_w9734_,
		_w10520_
	);
	LUT4 #(
		.INIT('hedff)
	) name9988 (
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9020_,
		_w10521_
	);
	LUT4 #(
		.INIT('h0155)
	) name9989 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		_w10520_,
		_w10521_,
		_w10522_
	);
	LUT2 #(
		.INIT('h4)
	) name9990 (
		\u0_w_reg[3][31]/P0001 ,
		_w10018_,
		_w10523_
	);
	LUT3 #(
		.INIT('h23)
	) name9991 (
		_w9030_,
		_w9061_,
		_w9980_,
		_w10524_
	);
	LUT3 #(
		.INIT('h8a)
	) name9992 (
		_w9063_,
		_w10523_,
		_w10524_,
		_w10525_
	);
	LUT4 #(
		.INIT('h7cfa)
	) name9993 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10526_
	);
	LUT3 #(
		.INIT('h04)
	) name9994 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w10527_
	);
	LUT2 #(
		.INIT('h4)
	) name9995 (
		_w10526_,
		_w10527_,
		_w10528_
	);
	LUT4 #(
		.INIT('hec00)
	) name9996 (
		_w8997_,
		_w9084_,
		_w9215_,
		_w10023_,
		_w10529_
	);
	LUT4 #(
		.INIT('h0001)
	) name9997 (
		_w9243_,
		_w9739_,
		_w10529_,
		_w10528_,
		_w10530_
	);
	LUT3 #(
		.INIT('h10)
	) name9998 (
		_w10525_,
		_w10522_,
		_w10530_,
		_w10531_
	);
	LUT4 #(
		.INIT('h5655)
	) name9999 (
		\u0_w_reg[0][1]/P0001 ,
		_w10519_,
		_w10509_,
		_w10531_,
		_w10532_
	);
	LUT2 #(
		.INIT('h9)
	) name10000 (
		\u0_w_reg[1][1]/P0001 ,
		\u0_w_reg[2][1]/P0001 ,
		_w10533_
	);
	LUT4 #(
		.INIT('hb88b)
	) name10001 (
		\key[33]_pad ,
		ld_pad,
		_w10532_,
		_w10533_,
		_w10534_
	);
	LUT2 #(
		.INIT('h8)
	) name10002 (
		_w9303_,
		_w9353_,
		_w10535_
	);
	LUT4 #(
		.INIT('h153f)
	) name10003 (
		\u0_w_reg[3][5]/P0001 ,
		_w9297_,
		_w9369_,
		_w9422_,
		_w10536_
	);
	LUT2 #(
		.INIT('h4)
	) name10004 (
		_w9268_,
		_w9327_,
		_w10537_
	);
	LUT3 #(
		.INIT('h15)
	) name10005 (
		\u0_w_reg[3][1]/P0001 ,
		_w9289_,
		_w9307_,
		_w10538_
	);
	LUT4 #(
		.INIT('h1000)
	) name10006 (
		_w10537_,
		_w10535_,
		_w10538_,
		_w10536_,
		_w10539_
	);
	LUT3 #(
		.INIT('h10)
	) name10007 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10540_
	);
	LUT4 #(
		.INIT('h0803)
	) name10008 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		_w10541_
	);
	LUT3 #(
		.INIT('h54)
	) name10009 (
		\u0_w_reg[3][2]/P0001 ,
		_w10540_,
		_w10541_,
		_w10542_
	);
	LUT4 #(
		.INIT('h4000)
	) name10010 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10543_
	);
	LUT3 #(
		.INIT('ha8)
	) name10011 (
		\u0_w_reg[3][2]/P0001 ,
		_w10063_,
		_w10543_,
		_w10544_
	);
	LUT4 #(
		.INIT('h0002)
	) name10012 (
		\u0_w_reg[3][1]/P0001 ,
		_w9379_,
		_w9401_,
		_w9411_,
		_w10545_
	);
	LUT3 #(
		.INIT('h10)
	) name10013 (
		_w10542_,
		_w10544_,
		_w10545_,
		_w10546_
	);
	LUT3 #(
		.INIT('h2a)
	) name10014 (
		\u0_w_reg[3][2]/P0001 ,
		_w9259_,
		_w9281_,
		_w10547_
	);
	LUT3 #(
		.INIT('h10)
	) name10015 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w9322_,
		_w10548_
	);
	LUT3 #(
		.INIT('hf4)
	) name10016 (
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10549_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10017 (
		\u0_w_reg[3][2]/P0001 ,
		_w9285_,
		_w9346_,
		_w10549_,
		_w10550_
	);
	LUT4 #(
		.INIT('h3200)
	) name10018 (
		_w9407_,
		_w10548_,
		_w10547_,
		_w10550_,
		_w10551_
	);
	LUT4 #(
		.INIT('h0155)
	) name10019 (
		\u0_w_reg[3][0]/P0001 ,
		_w10539_,
		_w10546_,
		_w10551_,
		_w10552_
	);
	LUT4 #(
		.INIT('haaa8)
	) name10020 (
		\u0_w_reg[3][2]/P0001 ,
		_w9265_,
		_w9845_,
		_w9818_,
		_w10553_
	);
	LUT3 #(
		.INIT('ha2)
	) name10021 (
		\u0_w_reg[3][1]/P0001 ,
		_w9815_,
		_w10553_,
		_w10554_
	);
	LUT4 #(
		.INIT('hfe77)
	) name10022 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10555_
	);
	LUT2 #(
		.INIT('h2)
	) name10023 (
		\u0_w_reg[3][5]/P0001 ,
		_w10555_,
		_w10556_
	);
	LUT3 #(
		.INIT('h0b)
	) name10024 (
		_w9317_,
		_w10176_,
		_w10270_,
		_w10557_
	);
	LUT3 #(
		.INIT('h45)
	) name10025 (
		\u0_w_reg[3][1]/P0001 ,
		_w10556_,
		_w10557_,
		_w10558_
	);
	LUT4 #(
		.INIT('h5504)
	) name10026 (
		\u0_w_reg[3][3]/P0001 ,
		_w9307_,
		_w9312_,
		_w9834_,
		_w10559_
	);
	LUT4 #(
		.INIT('h0001)
	) name10027 (
		_w9251_,
		_w9834_,
		_w9842_,
		_w10270_,
		_w10560_
	);
	LUT3 #(
		.INIT('h32)
	) name10028 (
		\u0_w_reg[3][2]/P0001 ,
		_w10559_,
		_w10560_,
		_w10561_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10029 (
		\u0_w_reg[3][0]/P0001 ,
		_w10554_,
		_w10558_,
		_w10561_,
		_w10562_
	);
	LUT4 #(
		.INIT('h0013)
	) name10030 (
		\u0_w_reg[3][4]/P0001 ,
		_w9309_,
		_w9346_,
		_w10037_,
		_w10563_
	);
	LUT4 #(
		.INIT('h135f)
	) name10031 (
		_w9259_,
		_w9256_,
		_w9281_,
		_w9336_,
		_w10564_
	);
	LUT4 #(
		.INIT('h0155)
	) name10032 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		_w10563_,
		_w10564_,
		_w10565_
	);
	LUT4 #(
		.INIT('hafac)
	) name10033 (
		\u0_w_reg[3][3]/P0001 ,
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10566_
	);
	LUT3 #(
		.INIT('h13)
	) name10034 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10567_
	);
	LUT2 #(
		.INIT('h4)
	) name10035 (
		_w10566_,
		_w10567_,
		_w10568_
	);
	LUT3 #(
		.INIT('h01)
	) name10036 (
		\u0_w_reg[3][2]/P0001 ,
		_w9401_,
		_w9831_,
		_w10569_
	);
	LUT2 #(
		.INIT('h4)
	) name10037 (
		_w10568_,
		_w10569_,
		_w10570_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name10038 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10571_
	);
	LUT2 #(
		.INIT('h2)
	) name10039 (
		\u0_w_reg[3][3]/P0001 ,
		_w10571_,
		_w10572_
	);
	LUT3 #(
		.INIT('ha2)
	) name10040 (
		\u0_w_reg[3][1]/P0001 ,
		_w10052_,
		_w10572_,
		_w10573_
	);
	LUT4 #(
		.INIT('h5040)
	) name10041 (
		\u0_w_reg[3][6]/P0001 ,
		_w9250_,
		_w9289_,
		_w9294_,
		_w10574_
	);
	LUT4 #(
		.INIT('h7cfa)
	) name10042 (
		\u0_w_reg[3][4]/P0001 ,
		\u0_w_reg[3][5]/P0001 ,
		\u0_w_reg[3][6]/P0001 ,
		\u0_w_reg[3][7]/P0001 ,
		_w10575_
	);
	LUT3 #(
		.INIT('h04)
	) name10043 (
		\u0_w_reg[3][1]/P0001 ,
		\u0_w_reg[3][2]/P0001 ,
		\u0_w_reg[3][3]/P0001 ,
		_w10576_
	);
	LUT2 #(
		.INIT('h4)
	) name10044 (
		_w10575_,
		_w10576_,
		_w10577_
	);
	LUT2 #(
		.INIT('h1)
	) name10045 (
		_w10574_,
		_w10577_,
		_w10578_
	);
	LUT4 #(
		.INIT('h4500)
	) name10046 (
		_w10565_,
		_w10570_,
		_w10573_,
		_w10578_,
		_w10579_
	);
	LUT4 #(
		.INIT('h5655)
	) name10047 (
		\u0_w_reg[0][9]/P0001 ,
		_w10562_,
		_w10552_,
		_w10579_,
		_w10580_
	);
	LUT2 #(
		.INIT('h9)
	) name10048 (
		\u0_w_reg[1][9]/P0001 ,
		\u0_w_reg[2][9]/P0001 ,
		_w10581_
	);
	LUT4 #(
		.INIT('hb88b)
	) name10049 (
		\key[41]_pad ,
		ld_pad,
		_w10580_,
		_w10581_,
		_w10582_
	);
	LUT4 #(
		.INIT('hb88b)
	) name10050 (
		\key[108]_pad ,
		ld_pad,
		\u0_w_reg[0][12]/P0001 ,
		_w9430_,
		_w10583_
	);
	LUT4 #(
		.INIT('h1441)
	) name10051 (
		ld_pad,
		\u0_w_reg[0][12]/P0001 ,
		\u0_w_reg[1][12]/P0001 ,
		_w9430_,
		_w10584_
	);
	LUT2 #(
		.INIT('h8)
	) name10052 (
		\key[76]_pad ,
		ld_pad,
		_w10585_
	);
	LUT2 #(
		.INIT('he)
	) name10053 (
		_w10584_,
		_w10585_,
		_w10586_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name10054 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10587_
	);
	LUT2 #(
		.INIT('h1)
	) name10055 (
		\u0_w_reg[3][10]/P0001 ,
		_w10587_,
		_w10588_
	);
	LUT3 #(
		.INIT('h07)
	) name10056 (
		_w8810_,
		_w8896_,
		_w9927_,
		_w10589_
	);
	LUT3 #(
		.INIT('h20)
	) name10057 (
		_w8806_,
		_w10588_,
		_w10589_,
		_w10590_
	);
	LUT3 #(
		.INIT('h54)
	) name10058 (
		\u0_w_reg[3][10]/P0001 ,
		_w8792_,
		_w8882_,
		_w10591_
	);
	LUT3 #(
		.INIT('h01)
	) name10059 (
		\u0_w_reg[3][9]/P0001 ,
		_w8845_,
		_w8960_,
		_w10592_
	);
	LUT2 #(
		.INIT('h4)
	) name10060 (
		_w10591_,
		_w10592_,
		_w10593_
	);
	LUT3 #(
		.INIT('h04)
	) name10061 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10594_
	);
	LUT4 #(
		.INIT('haaa8)
	) name10062 (
		\u0_w_reg[3][10]/P0001 ,
		_w8849_,
		_w8896_,
		_w10594_,
		_w10595_
	);
	LUT4 #(
		.INIT('h0203)
	) name10063 (
		\u0_w_reg[3][15]/P0001 ,
		_w8818_,
		_w8918_,
		_w9876_,
		_w10596_
	);
	LUT2 #(
		.INIT('h8)
	) name10064 (
		_w8861_,
		_w8962_,
		_w10597_
	);
	LUT3 #(
		.INIT('h2a)
	) name10065 (
		\u0_w_reg[3][8]/P0001 ,
		_w8786_,
		_w8851_,
		_w10598_
	);
	LUT4 #(
		.INIT('h0e00)
	) name10066 (
		\u0_w_reg[3][10]/P0001 ,
		_w10596_,
		_w10597_,
		_w10598_,
		_w10599_
	);
	LUT4 #(
		.INIT('h5400)
	) name10067 (
		_w10595_,
		_w10590_,
		_w10593_,
		_w10599_,
		_w10600_
	);
	LUT3 #(
		.INIT('hd0)
	) name10068 (
		\u0_w_reg[3][11]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		_w10601_
	);
	LUT4 #(
		.INIT('h5450)
	) name10069 (
		\u0_w_reg[3][10]/P0001 ,
		_w8785_,
		_w8956_,
		_w10601_,
		_w10602_
	);
	LUT2 #(
		.INIT('h8)
	) name10070 (
		_w8937_,
		_w8914_,
		_w10603_
	);
	LUT3 #(
		.INIT('h02)
	) name10071 (
		\u0_w_reg[3][9]/P0001 ,
		_w8948_,
		_w9869_,
		_w10604_
	);
	LUT3 #(
		.INIT('h10)
	) name10072 (
		_w10602_,
		_w10603_,
		_w10604_,
		_w10605_
	);
	LUT3 #(
		.INIT('h01)
	) name10073 (
		\u0_w_reg[3][9]/P0001 ,
		_w8852_,
		_w8889_,
		_w10606_
	);
	LUT4 #(
		.INIT('h8000)
	) name10074 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		_w10607_
	);
	LUT3 #(
		.INIT('h07)
	) name10075 (
		_w8784_,
		_w8883_,
		_w10607_,
		_w10608_
	);
	LUT2 #(
		.INIT('h8)
	) name10076 (
		_w10606_,
		_w10608_,
		_w10609_
	);
	LUT4 #(
		.INIT('ha888)
	) name10077 (
		\u0_w_reg[3][10]/P0001 ,
		_w8816_,
		_w8790_,
		_w8910_,
		_w10610_
	);
	LUT4 #(
		.INIT('h5540)
	) name10078 (
		\u0_w_reg[3][11]/P0001 ,
		_w8796_,
		_w8828_,
		_w9907_,
		_w10611_
	);
	LUT3 #(
		.INIT('h01)
	) name10079 (
		\u0_w_reg[3][8]/P0001 ,
		_w10611_,
		_w10610_,
		_w10612_
	);
	LUT3 #(
		.INIT('he0)
	) name10080 (
		_w10605_,
		_w10609_,
		_w10612_,
		_w10613_
	);
	LUT4 #(
		.INIT('hcc40)
	) name10081 (
		\u0_w_reg[3][10]/P0001 ,
		\u0_w_reg[3][11]/P0001 ,
		_w8964_,
		_w10607_,
		_w10614_
	);
	LUT2 #(
		.INIT('h2)
	) name10082 (
		_w8803_,
		_w8944_,
		_w10615_
	);
	LUT3 #(
		.INIT('h01)
	) name10083 (
		_w8800_,
		_w9916_,
		_w9964_,
		_w10616_
	);
	LUT3 #(
		.INIT('h8a)
	) name10084 (
		\u0_w_reg[3][10]/P0001 ,
		_w10615_,
		_w10616_,
		_w10617_
	);
	LUT3 #(
		.INIT('h23)
	) name10085 (
		\u0_w_reg[3][15]/P0001 ,
		\u0_w_reg[3][9]/P0001 ,
		_w9966_,
		_w10618_
	);
	LUT4 #(
		.INIT('h3020)
	) name10086 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10619_
	);
	LUT2 #(
		.INIT('h8)
	) name10087 (
		_w8883_,
		_w10619_,
		_w10620_
	);
	LUT4 #(
		.INIT('h153f)
	) name10088 (
		_w8791_,
		_w8849_,
		_w8878_,
		_w8905_,
		_w10621_
	);
	LUT3 #(
		.INIT('h40)
	) name10089 (
		_w10620_,
		_w10618_,
		_w10621_,
		_w10622_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name10090 (
		\u0_w_reg[3][14]/P0001 ,
		_w8854_,
		_w9878_,
		_w9901_,
		_w10623_
	);
	LUT4 #(
		.INIT('h153f)
	) name10091 (
		\u0_w_reg[3][12]/P0001 ,
		_w8878_,
		_w9898_,
		_w9926_,
		_w10624_
	);
	LUT4 #(
		.INIT('hbffe)
	) name10092 (
		\u0_w_reg[3][12]/P0001 ,
		\u0_w_reg[3][13]/P0001 ,
		\u0_w_reg[3][14]/P0001 ,
		\u0_w_reg[3][15]/P0001 ,
		_w10625_
	);
	LUT2 #(
		.INIT('h2)
	) name10093 (
		_w8883_,
		_w10625_,
		_w10626_
	);
	LUT4 #(
		.INIT('h2000)
	) name10094 (
		_w10412_,
		_w10626_,
		_w10623_,
		_w10624_,
		_w10627_
	);
	LUT4 #(
		.INIT('h5510)
	) name10095 (
		_w10614_,
		_w10617_,
		_w10622_,
		_w10627_,
		_w10628_
	);
	LUT4 #(
		.INIT('ha955)
	) name10096 (
		\u0_w_reg[0][20]/P0001 ,
		_w10600_,
		_w10613_,
		_w10628_,
		_w10629_
	);
	LUT3 #(
		.INIT('h96)
	) name10097 (
		\u0_w_reg[1][20]/P0001 ,
		\u0_w_reg[2][20]/P0001 ,
		_w10629_,
		_w10630_
	);
	LUT4 #(
		.INIT('h4114)
	) name10098 (
		ld_pad,
		\u0_w_reg[1][20]/P0001 ,
		\u0_w_reg[2][20]/P0001 ,
		_w10629_,
		_w10631_
	);
	LUT2 #(
		.INIT('h8)
	) name10099 (
		\key[52]_pad ,
		ld_pad,
		_w10632_
	);
	LUT2 #(
		.INIT('he)
	) name10100 (
		_w10631_,
		_w10632_,
		_w10633_
	);
	LUT4 #(
		.INIT('h5510)
	) name10101 (
		\u0_w_reg[3][26]/P0001 ,
		_w9047_,
		_w9052_,
		_w9233_,
		_w10634_
	);
	LUT4 #(
		.INIT('h0080)
	) name10102 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10635_
	);
	LUT4 #(
		.INIT('h0007)
	) name10103 (
		_w9068_,
		_w9189_,
		_w9225_,
		_w10635_,
		_w10636_
	);
	LUT3 #(
		.INIT('h8a)
	) name10104 (
		\u0_w_reg[3][25]/P0001 ,
		_w10634_,
		_w10636_,
		_w10637_
	);
	LUT2 #(
		.INIT('h4)
	) name10105 (
		\u0_w_reg[3][26]/P0001 ,
		_w9770_,
		_w10638_
	);
	LUT4 #(
		.INIT('h8000)
	) name10106 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w10639_
	);
	LUT3 #(
		.INIT('h01)
	) name10107 (
		_w9736_,
		_w10160_,
		_w10639_,
		_w10640_
	);
	LUT3 #(
		.INIT('h45)
	) name10108 (
		\u0_w_reg[3][25]/P0001 ,
		_w10638_,
		_w10640_,
		_w10641_
	);
	LUT4 #(
		.INIT('h3310)
	) name10109 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w9058_,
		_w9091_,
		_w10642_
	);
	LUT4 #(
		.INIT('h0100)
	) name10110 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w10643_
	);
	LUT4 #(
		.INIT('haa20)
	) name10111 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		_w9041_,
		_w10643_,
		_w10644_
	);
	LUT2 #(
		.INIT('h1)
	) name10112 (
		_w10642_,
		_w10644_,
		_w10645_
	);
	LUT4 #(
		.INIT('h5455)
	) name10113 (
		\u0_w_reg[3][24]/P0001 ,
		_w10641_,
		_w10637_,
		_w10645_,
		_w10646_
	);
	LUT3 #(
		.INIT('h40)
	) name10114 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10647_
	);
	LUT3 #(
		.INIT('h54)
	) name10115 (
		\u0_w_reg[3][26]/P0001 ,
		_w9041_,
		_w10647_,
		_w10648_
	);
	LUT4 #(
		.INIT('h1555)
	) name10116 (
		\u0_w_reg[3][25]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10649_
	);
	LUT2 #(
		.INIT('h4)
	) name10117 (
		_w9985_,
		_w10649_,
		_w10650_
	);
	LUT2 #(
		.INIT('h4)
	) name10118 (
		_w10648_,
		_w10650_,
		_w10651_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name10119 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10652_
	);
	LUT2 #(
		.INIT('h1)
	) name10120 (
		\u0_w_reg[3][26]/P0001 ,
		_w10652_,
		_w10653_
	);
	LUT4 #(
		.INIT('h002a)
	) name10121 (
		\u0_w_reg[3][25]/P0001 ,
		_w8977_,
		_w9053_,
		_w9984_,
		_w10654_
	);
	LUT3 #(
		.INIT('h10)
	) name10122 (
		_w9800_,
		_w10653_,
		_w10654_,
		_w10655_
	);
	LUT3 #(
		.INIT('h0b)
	) name10123 (
		\u0_w_reg[3][25]/P0001 ,
		_w9031_,
		_w9223_,
		_w10656_
	);
	LUT3 #(
		.INIT('h23)
	) name10124 (
		\u0_w_reg[3][31]/P0001 ,
		_w9056_,
		_w9783_,
		_w10657_
	);
	LUT4 #(
		.INIT('h135f)
	) name10125 (
		_w10138_,
		_w10143_,
		_w10656_,
		_w10657_,
		_w10658_
	);
	LUT4 #(
		.INIT('h0008)
	) name10126 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		_w10659_
	);
	LUT2 #(
		.INIT('h1)
	) name10127 (
		_w9095_,
		_w10659_,
		_w10660_
	);
	LUT4 #(
		.INIT('h5400)
	) name10128 (
		_w10658_,
		_w10651_,
		_w10655_,
		_w10660_,
		_w10661_
	);
	LUT4 #(
		.INIT('h0015)
	) name10129 (
		_w9043_,
		_w8987_,
		_w9021_,
		_w9689_,
		_w10662_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10130 (
		\u0_w_reg[3][26]/P0001 ,
		_w9981_,
		_w9994_,
		_w10662_,
		_w10663_
	);
	LUT4 #(
		.INIT('hcecf)
	) name10131 (
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w9084_,
		_w9082_,
		_w10664_
	);
	LUT4 #(
		.INIT('h3020)
	) name10132 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10665_
	);
	LUT4 #(
		.INIT('haebf)
	) name10133 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w9223_,
		_w10665_,
		_w10666_
	);
	LUT2 #(
		.INIT('h8)
	) name10134 (
		_w10664_,
		_w10666_,
		_w10667_
	);
	LUT3 #(
		.INIT('h45)
	) name10135 (
		\u0_w_reg[3][25]/P0001 ,
		_w10663_,
		_w10667_,
		_w10668_
	);
	LUT4 #(
		.INIT('h4440)
	) name10136 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10669_
	);
	LUT4 #(
		.INIT('h7dff)
	) name10137 (
		\u0_w_reg[3][27]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10670_
	);
	LUT3 #(
		.INIT('h45)
	) name10138 (
		\u0_w_reg[3][29]/P0001 ,
		_w10669_,
		_w10670_,
		_w10671_
	);
	LUT4 #(
		.INIT('hbffe)
	) name10139 (
		\u0_w_reg[3][28]/P0001 ,
		\u0_w_reg[3][29]/P0001 ,
		\u0_w_reg[3][30]/P0001 ,
		\u0_w_reg[3][31]/P0001 ,
		_w10672_
	);
	LUT2 #(
		.INIT('h2)
	) name10140 (
		_w9197_,
		_w10672_,
		_w10673_
	);
	LUT4 #(
		.INIT('h57df)
	) name10141 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w9680_,
		_w9709_,
		_w10674_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10142 (
		\u0_w_reg[3][25]/P0001 ,
		_w10673_,
		_w10671_,
		_w10674_,
		_w10675_
	);
	LUT4 #(
		.INIT('hcc40)
	) name10143 (
		\u0_w_reg[3][26]/P0001 ,
		\u0_w_reg[3][27]/P0001 ,
		_w9070_,
		_w10639_,
		_w10676_
	);
	LUT2 #(
		.INIT('h1)
	) name10144 (
		_w10675_,
		_w10676_,
		_w10677_
	);
	LUT4 #(
		.INIT('h3100)
	) name10145 (
		\u0_w_reg[3][24]/P0001 ,
		_w10668_,
		_w10661_,
		_w10677_,
		_w10678_
	);
	LUT3 #(
		.INIT('h65)
	) name10146 (
		\u0_w_reg[0][4]/P0001 ,
		_w10646_,
		_w10678_,
		_w10679_
	);
	LUT2 #(
		.INIT('h9)
	) name10147 (
		\u0_w_reg[1][4]/P0001 ,
		\u0_w_reg[2][4]/P0001 ,
		_w10680_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10148 (
		\u0_w_reg[0][4]/P0001 ,
		_w10646_,
		_w10678_,
		_w10680_,
		_w10681_
	);
	LUT3 #(
		.INIT('h8b)
	) name10149 (
		\key[36]_pad ,
		ld_pad,
		_w10681_,
		_w10682_
	);
	LUT4 #(
		.INIT('hb88b)
	) name10150 (
		\key[12]_pad ,
		ld_pad,
		\u0_w_reg[3][12]/P0001 ,
		_w9432_,
		_w10683_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name10151 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10684_
	);
	LUT2 #(
		.INIT('h1)
	) name10152 (
		\u0_w_reg[3][18]/P0001 ,
		_w10684_,
		_w10685_
	);
	LUT3 #(
		.INIT('h07)
	) name10153 (
		_w8654_,
		_w8681_,
		_w9495_,
		_w10686_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10154 (
		\u0_w_reg[3][17]/P0001 ,
		_w8768_,
		_w10685_,
		_w10686_,
		_w10687_
	);
	LUT3 #(
		.INIT('h54)
	) name10155 (
		\u0_w_reg[3][18]/P0001 ,
		_w8727_,
		_w8668_,
		_w10688_
	);
	LUT2 #(
		.INIT('h1)
	) name10156 (
		_w8673_,
		_w9496_,
		_w10689_
	);
	LUT3 #(
		.INIT('h45)
	) name10157 (
		\u0_w_reg[3][17]/P0001 ,
		_w10688_,
		_w10689_,
		_w10690_
	);
	LUT4 #(
		.INIT('h5ffe)
	) name10158 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10691_
	);
	LUT4 #(
		.INIT('h5051)
	) name10159 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		_w8738_,
		_w10691_,
		_w10692_
	);
	LUT4 #(
		.INIT('h0008)
	) name10160 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w10693_
	);
	LUT4 #(
		.INIT('h0020)
	) name10161 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10694_
	);
	LUT4 #(
		.INIT('h0007)
	) name10162 (
		_w8730_,
		_w8689_,
		_w10693_,
		_w10694_,
		_w10695_
	);
	LUT4 #(
		.INIT('h33bf)
	) name10163 (
		\u0_w_reg[3][17]/P0001 ,
		\u0_w_reg[3][18]/P0001 ,
		_w8708_,
		_w9114_,
		_w10696_
	);
	LUT3 #(
		.INIT('h40)
	) name10164 (
		_w10692_,
		_w10695_,
		_w10696_,
		_w10697_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10165 (
		\u0_w_reg[3][16]/P0001 ,
		_w10690_,
		_w10687_,
		_w10697_,
		_w10698_
	);
	LUT4 #(
		.INIT('h5150)
	) name10166 (
		\u0_w_reg[3][18]/P0001 ,
		_w8714_,
		_w9159_,
		_w9574_,
		_w10699_
	);
	LUT2 #(
		.INIT('h8)
	) name10167 (
		_w8732_,
		_w8684_,
		_w10700_
	);
	LUT3 #(
		.INIT('h02)
	) name10168 (
		\u0_w_reg[3][17]/P0001 ,
		_w9108_,
		_w9456_,
		_w10701_
	);
	LUT3 #(
		.INIT('h10)
	) name10169 (
		_w10699_,
		_w10700_,
		_w10701_,
		_w10702_
	);
	LUT2 #(
		.INIT('h4)
	) name10170 (
		\u0_w_reg[3][18]/P0001 ,
		_w9451_,
		_w10703_
	);
	LUT4 #(
		.INIT('h8000)
	) name10171 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w10704_
	);
	LUT4 #(
		.INIT('h0002)
	) name10172 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10705_
	);
	LUT4 #(
		.INIT('h0001)
	) name10173 (
		\u0_w_reg[3][17]/P0001 ,
		_w8682_,
		_w10704_,
		_w10705_,
		_w10706_
	);
	LUT2 #(
		.INIT('h4)
	) name10174 (
		_w10703_,
		_w10706_,
		_w10707_
	);
	LUT4 #(
		.INIT('h0100)
	) name10175 (
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		_w10708_
	);
	LUT4 #(
		.INIT('haa20)
	) name10176 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		_w8727_,
		_w10708_,
		_w10709_
	);
	LUT4 #(
		.INIT('h3310)
	) name10177 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w8740_,
		_w9479_,
		_w10710_
	);
	LUT2 #(
		.INIT('h1)
	) name10178 (
		_w10709_,
		_w10710_,
		_w10711_
	);
	LUT4 #(
		.INIT('h0155)
	) name10179 (
		\u0_w_reg[3][16]/P0001 ,
		_w10702_,
		_w10707_,
		_w10711_,
		_w10712_
	);
	LUT4 #(
		.INIT('hfef3)
	) name10180 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10713_
	);
	LUT2 #(
		.INIT('h1)
	) name10181 (
		\u0_w_reg[3][19]/P0001 ,
		_w10713_,
		_w10714_
	);
	LUT4 #(
		.INIT('h0015)
	) name10182 (
		_w8737_,
		_w8723_,
		_w8683_,
		_w8767_,
		_w10715_
	);
	LUT3 #(
		.INIT('h8a)
	) name10183 (
		\u0_w_reg[3][18]/P0001 ,
		_w10714_,
		_w10715_,
		_w10716_
	);
	LUT4 #(
		.INIT('h135f)
	) name10184 (
		_w8746_,
		_w8729_,
		_w8664_,
		_w9114_,
		_w10717_
	);
	LUT3 #(
		.INIT('hc8)
	) name10185 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10718_
	);
	LUT4 #(
		.INIT('h2777)
	) name10186 (
		\u0_w_reg[3][21]/P0001 ,
		_w8751_,
		_w8764_,
		_w10718_,
		_w10719_
	);
	LUT2 #(
		.INIT('h8)
	) name10187 (
		_w10717_,
		_w10719_,
		_w10720_
	);
	LUT3 #(
		.INIT('h45)
	) name10188 (
		\u0_w_reg[3][17]/P0001 ,
		_w10716_,
		_w10720_,
		_w10721_
	);
	LUT4 #(
		.INIT('hc480)
	) name10189 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		_w8746_,
		_w9164_,
		_w10722_
	);
	LUT2 #(
		.INIT('h8)
	) name10190 (
		\u0_w_reg[3][20]/P0001 ,
		_w9494_,
		_w10723_
	);
	LUT4 #(
		.INIT('h135f)
	) name10191 (
		_w8697_,
		_w8689_,
		_w9134_,
		_w9464_,
		_w10724_
	);
	LUT4 #(
		.INIT('h4440)
	) name10192 (
		\u0_w_reg[3][18]/P0001 ,
		\u0_w_reg[3][19]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10725_
	);
	LUT3 #(
		.INIT('h54)
	) name10193 (
		\u0_w_reg[3][21]/P0001 ,
		_w8718_,
		_w10725_,
		_w10726_
	);
	LUT4 #(
		.INIT('hbffe)
	) name10194 (
		\u0_w_reg[3][20]/P0001 ,
		\u0_w_reg[3][21]/P0001 ,
		\u0_w_reg[3][22]/P0001 ,
		\u0_w_reg[3][23]/P0001 ,
		_w10727_
	);
	LUT2 #(
		.INIT('h2)
	) name10195 (
		_w8764_,
		_w10727_,
		_w10728_
	);
	LUT4 #(
		.INIT('h0100)
	) name10196 (
		_w10723_,
		_w10726_,
		_w10728_,
		_w10724_,
		_w10729_
	);
	LUT3 #(
		.INIT('h31)
	) name10197 (
		\u0_w_reg[3][17]/P0001 ,
		_w10722_,
		_w10729_,
		_w10730_
	);
	LUT4 #(
		.INIT('h0100)
	) name10198 (
		_w10698_,
		_w10721_,
		_w10712_,
		_w10730_,
		_w10731_
	);
	LUT3 #(
		.INIT('h69)
	) name10199 (
		\u0_r0_out_reg[28]/P0001 ,
		\u0_w_reg[0][28]/P0001 ,
		_w10731_,
		_w10732_
	);
	LUT4 #(
		.INIT('h1441)
	) name10200 (
		ld_pad,
		\u0_r0_out_reg[28]/P0001 ,
		\u0_w_reg[0][28]/P0001 ,
		_w10731_,
		_w10733_
	);
	LUT2 #(
		.INIT('h8)
	) name10201 (
		\key[124]_pad ,
		ld_pad,
		_w10734_
	);
	LUT2 #(
		.INIT('he)
	) name10202 (
		_w10733_,
		_w10734_,
		_w10735_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10203 (
		\key[92]_pad ,
		ld_pad,
		\u0_w_reg[1][28]/P0001 ,
		_w10732_,
		_w10736_
	);
	LUT2 #(
		.INIT('h9)
	) name10204 (
		\u0_w_reg[0][28]/P0001 ,
		\u0_w_reg[2][28]/P0001 ,
		_w10737_
	);
	LUT3 #(
		.INIT('h69)
	) name10205 (
		\u0_r0_out_reg[28]/P0001 ,
		_w10731_,
		_w10737_,
		_w10738_
	);
	LUT4 #(
		.INIT('hb88b)
	) name10206 (
		\key[60]_pad ,
		ld_pad,
		\u0_w_reg[1][28]/P0001 ,
		_w10738_,
		_w10739_
	);
	LUT2 #(
		.INIT('h9)
	) name10207 (
		\u0_w_reg[1][28]/P0001 ,
		\u0_w_reg[3][28]/P0001 ,
		_w10740_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10208 (
		\key[28]_pad ,
		ld_pad,
		_w10738_,
		_w10740_,
		_w10741_
	);
	LUT4 #(
		.INIT('h1114)
	) name10209 (
		ld_pad,
		\u0_w_reg[0][7]/P0001 ,
		_w9720_,
		_w9741_,
		_w10742_
	);
	LUT2 #(
		.INIT('h8)
	) name10210 (
		\key[103]_pad ,
		ld_pad,
		_w10743_
	);
	LUT2 #(
		.INIT('he)
	) name10211 (
		_w10742_,
		_w10743_,
		_w10744_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10212 (
		\key[71]_pad ,
		ld_pad,
		\u0_w_reg[1][7]/P0001 ,
		_w9742_,
		_w10745_
	);
	LUT4 #(
		.INIT('hb88b)
	) name10213 (
		\key[7]_pad ,
		ld_pad,
		\u0_w_reg[3][7]/P0001 ,
		_w9744_,
		_w10746_
	);
	LUT3 #(
		.INIT('hb8)
	) name10214 (
		\key[96]_pad ,
		ld_pad,
		_w9804_,
		_w10747_
	);
	LUT3 #(
		.INIT('hb8)
	) name10215 (
		\key[106]_pad ,
		ld_pad,
		_w9860_,
		_w10748_
	);
	LUT3 #(
		.INIT('hb8)
	) name10216 (
		\key[112]_pad ,
		ld_pad,
		_w9923_,
		_w10749_
	);
	LUT3 #(
		.INIT('hb8)
	) name10217 (
		\key[114]_pad ,
		ld_pad,
		_w9976_,
		_w10750_
	);
	LUT3 #(
		.INIT('hb8)
	) name10218 (
		\key[98]_pad ,
		ld_pad,
		_w10029_,
		_w10751_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10219 (
		\key[64]_pad ,
		ld_pad,
		\u0_w_reg[1][0]/P0001 ,
		_w9804_,
		_w10752_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10220 (
		\key[74]_pad ,
		ld_pad,
		\u0_w_reg[1][10]/P0001 ,
		_w9860_,
		_w10753_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10221 (
		\key[80]_pad ,
		ld_pad,
		\u0_w_reg[1][16]/P0001 ,
		_w9923_,
		_w10754_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10222 (
		\key[82]_pad ,
		ld_pad,
		\u0_w_reg[1][18]/P0001 ,
		_w9976_,
		_w10755_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10223 (
		\key[66]_pad ,
		ld_pad,
		\u0_w_reg[1][2]/P0001 ,
		_w10029_,
		_w10756_
	);
	LUT4 #(
		.INIT('h1441)
	) name10224 (
		ld_pad,
		\u0_w_reg[3][0]/P0001 ,
		_w9804_,
		_w9805_,
		_w10757_
	);
	LUT2 #(
		.INIT('h8)
	) name10225 (
		\key[0]_pad ,
		ld_pad,
		_w10758_
	);
	LUT2 #(
		.INIT('he)
	) name10226 (
		_w10757_,
		_w10758_,
		_w10759_
	);
	LUT4 #(
		.INIT('h1441)
	) name10227 (
		ld_pad,
		\u0_w_reg[3][10]/P0001 ,
		_w9860_,
		_w9861_,
		_w10760_
	);
	LUT2 #(
		.INIT('h8)
	) name10228 (
		\key[10]_pad ,
		ld_pad,
		_w10761_
	);
	LUT2 #(
		.INIT('he)
	) name10229 (
		_w10760_,
		_w10761_,
		_w10762_
	);
	LUT4 #(
		.INIT('h1441)
	) name10230 (
		ld_pad,
		\u0_w_reg[3][16]/P0001 ,
		_w9923_,
		_w9924_,
		_w10763_
	);
	LUT2 #(
		.INIT('h8)
	) name10231 (
		\key[16]_pad ,
		ld_pad,
		_w10764_
	);
	LUT2 #(
		.INIT('he)
	) name10232 (
		_w10763_,
		_w10764_,
		_w10765_
	);
	LUT4 #(
		.INIT('h1441)
	) name10233 (
		ld_pad,
		\u0_w_reg[3][18]/P0001 ,
		_w9976_,
		_w9977_,
		_w10766_
	);
	LUT2 #(
		.INIT('h8)
	) name10234 (
		\key[18]_pad ,
		ld_pad,
		_w10767_
	);
	LUT2 #(
		.INIT('he)
	) name10235 (
		_w10766_,
		_w10767_,
		_w10768_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10236 (
		\key[2]_pad ,
		ld_pad,
		\u0_w_reg[3][2]/P0001 ,
		_w10030_,
		_w10769_
	);
	LUT3 #(
		.INIT('h65)
	) name10237 (
		\u0_w_reg[0][5]/P0001 ,
		_w7074_,
		_w7146_,
		_w10770_
	);
	LUT3 #(
		.INIT('hb8)
	) name10238 (
		\key[110]_pad ,
		ld_pad,
		_w10080_,
		_w10771_
	);
	LUT3 #(
		.INIT('hb8)
	) name10239 (
		\key[118]_pad ,
		ld_pad,
		_w10124_,
		_w10772_
	);
	LUT4 #(
		.INIT('hb88b)
	) name10240 (
		\key[102]_pad ,
		ld_pad,
		\u0_w_reg[0][6]/P0001 ,
		_w10170_,
		_w10773_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10241 (
		\key[78]_pad ,
		ld_pad,
		\u0_w_reg[1][14]/P0001 ,
		_w10080_,
		_w10774_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10242 (
		\key[86]_pad ,
		ld_pad,
		\u0_w_reg[1][22]/P0001 ,
		_w10124_,
		_w10775_
	);
	LUT4 #(
		.INIT('h1441)
	) name10243 (
		ld_pad,
		\u0_w_reg[0][6]/P0001 ,
		\u0_w_reg[1][6]/P0001 ,
		_w10170_,
		_w10776_
	);
	LUT2 #(
		.INIT('h8)
	) name10244 (
		\key[70]_pad ,
		ld_pad,
		_w10777_
	);
	LUT2 #(
		.INIT('he)
	) name10245 (
		_w10776_,
		_w10777_,
		_w10778_
	);
	LUT4 #(
		.INIT('h1441)
	) name10246 (
		ld_pad,
		\u0_w_reg[3][14]/P0001 ,
		_w10080_,
		_w10081_,
		_w10779_
	);
	LUT2 #(
		.INIT('h8)
	) name10247 (
		\key[14]_pad ,
		ld_pad,
		_w10780_
	);
	LUT2 #(
		.INIT('he)
	) name10248 (
		_w10779_,
		_w10780_,
		_w10781_
	);
	LUT4 #(
		.INIT('h1441)
	) name10249 (
		ld_pad,
		\u0_w_reg[3][22]/P0001 ,
		_w10124_,
		_w10125_,
		_w10782_
	);
	LUT2 #(
		.INIT('h8)
	) name10250 (
		\key[22]_pad ,
		ld_pad,
		_w10783_
	);
	LUT2 #(
		.INIT('he)
	) name10251 (
		_w10782_,
		_w10783_,
		_w10784_
	);
	LUT4 #(
		.INIT('hb88b)
	) name10252 (
		\key[6]_pad ,
		ld_pad,
		\u0_w_reg[3][6]/P0001 ,
		_w10172_,
		_w10785_
	);
	LUT4 #(
		.INIT('hb88b)
	) name10253 (
		\key[109]_pad ,
		ld_pad,
		\u0_w_reg[0][13]/P0001 ,
		_w10224_,
		_w10786_
	);
	LUT3 #(
		.INIT('hb8)
	) name10254 (
		\key[111]_pad ,
		ld_pad,
		_w10283_,
		_w10787_
	);
	LUT4 #(
		.INIT('hb88b)
	) name10255 (
		\key[104]_pad ,
		ld_pad,
		\u0_w_reg[0][8]/P0001 ,
		_w10330_,
		_w10788_
	);
	LUT4 #(
		.INIT('h1441)
	) name10256 (
		ld_pad,
		\u0_w_reg[0][13]/P0001 ,
		\u0_w_reg[1][13]/P0001 ,
		_w10224_,
		_w10789_
	);
	LUT2 #(
		.INIT('h8)
	) name10257 (
		\key[77]_pad ,
		ld_pad,
		_w10790_
	);
	LUT2 #(
		.INIT('he)
	) name10258 (
		_w10789_,
		_w10790_,
		_w10791_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10259 (
		\key[79]_pad ,
		ld_pad,
		\u0_w_reg[1][15]/P0001 ,
		_w10283_,
		_w10792_
	);
	LUT4 #(
		.INIT('h1441)
	) name10260 (
		ld_pad,
		\u0_w_reg[0][8]/P0001 ,
		\u0_w_reg[1][8]/P0001 ,
		_w10330_,
		_w10793_
	);
	LUT2 #(
		.INIT('h8)
	) name10261 (
		\key[72]_pad ,
		ld_pad,
		_w10794_
	);
	LUT2 #(
		.INIT('he)
	) name10262 (
		_w10793_,
		_w10794_,
		_w10795_
	);
	LUT4 #(
		.INIT('hb88b)
	) name10263 (
		\key[13]_pad ,
		ld_pad,
		\u0_w_reg[3][13]/P0001 ,
		_w10226_,
		_w10796_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10264 (
		\key[15]_pad ,
		ld_pad,
		\u0_w_reg[3][15]/P0001 ,
		_w10284_,
		_w10797_
	);
	LUT4 #(
		.INIT('hb88b)
	) name10265 (
		\key[8]_pad ,
		ld_pad,
		\u0_w_reg[3][8]/P0001 ,
		_w10332_,
		_w10798_
	);
	LUT2 #(
		.INIT('h9)
	) name10266 (
		\u0_w_reg[0][29]/P0001 ,
		_w7224_,
		_w10799_
	);
	LUT4 #(
		.INIT('h5655)
	) name10267 (
		\u0_w_reg[3][29]/P0001 ,
		_w1129_,
		_w1086_,
		_w1148_,
		_w10800_
	);
	LUT2 #(
		.INIT('h9)
	) name10268 (
		\u0_w_reg[2][29]/P0001 ,
		_w933_,
		_w10801_
	);
	LUT2 #(
		.INIT('h9)
	) name10269 (
		\u0_w_reg[1][29]/P0002 ,
		_w5389_,
		_w10802_
	);
	LUT3 #(
		.INIT('hb8)
	) name10270 (
		\key[119]_pad ,
		ld_pad,
		_w10435_,
		_w10803_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10271 (
		\key[87]_pad ,
		ld_pad,
		\u0_w_reg[1][23]/P0001 ,
		_w10435_,
		_w10804_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10272 (
		\key[23]_pad ,
		ld_pad,
		\u0_w_reg[3][23]/P0001 ,
		_w10436_,
		_w10805_
	);
	LUT4 #(
		.INIT('h5655)
	) name10273 (
		\u0_w_reg[3][8]/P0001 ,
		_w2376_,
		_w2360_,
		_w2387_,
		_w10806_
	);
	LUT2 #(
		.INIT('h9)
	) name10274 (
		\u0_w_reg[0][11]/P0001 ,
		_w8262_,
		_w10807_
	);
	LUT4 #(
		.INIT('h5655)
	) name10275 (
		\u0_w_reg[3][11]/P0001 ,
		_w2625_,
		_w2612_,
		_w2640_,
		_w10808_
	);
	LUT2 #(
		.INIT('h9)
	) name10276 (
		\u0_w_reg[2][11]/P0001 ,
		_w4236_,
		_w10809_
	);
	LUT4 #(
		.INIT('h5655)
	) name10277 (
		\u0_w_reg[1][11]/P0001 ,
		_w6181_,
		_w6164_,
		_w6194_,
		_w10810_
	);
	LUT2 #(
		.INIT('h9)
	) name10278 (
		\u0_w_reg[0][12]/P0001 ,
		_w7295_,
		_w10811_
	);
	LUT2 #(
		.INIT('h9)
	) name10279 (
		\u0_w_reg[2][12]/P0001 ,
		_w3616_,
		_w10812_
	);
	LUT2 #(
		.INIT('h9)
	) name10280 (
		\u0_w_reg[1][12]/P0001 ,
		_w5517_,
		_w10813_
	);
	LUT4 #(
		.INIT('h5655)
	) name10281 (
		\u0_w_reg[0][8]/P0001 ,
		_w7574_,
		_w7590_,
		_w7602_,
		_w10814_
	);
	LUT4 #(
		.INIT('h5655)
	) name10282 (
		\u0_w_reg[0][24]/P0001 ,
		_w8108_,
		_w8090_,
		_w8122_,
		_w10815_
	);
	LUT4 #(
		.INIT('h5655)
	) name10283 (
		\u0_w_reg[0][27]/P0001 ,
		_w8468_,
		_w8455_,
		_w8479_,
		_w10816_
	);
	LUT2 #(
		.INIT('h9)
	) name10284 (
		\u0_w_reg[3][24]/P0001 ,
		_w2685_,
		_w10817_
	);
	LUT4 #(
		.INIT('h5655)
	) name10285 (
		\u0_w_reg[3][27]/P0001 ,
		_w2521_,
		_w2534_,
		_w2546_,
		_w10818_
	);
	LUT4 #(
		.INIT('h5655)
	) name10286 (
		\u0_w_reg[2][8]/P0001 ,
		_w4066_,
		_w4080_,
		_w4092_,
		_w10819_
	);
	LUT2 #(
		.INIT('h9)
	) name10287 (
		\u0_w_reg[2][24]/P0001 ,
		_w3841_,
		_w10820_
	);
	LUT4 #(
		.INIT('h5655)
	) name10288 (
		\u0_w_reg[2][27]/P0001 ,
		_w4131_,
		_w4118_,
		_w4144_,
		_w10821_
	);
	LUT3 #(
		.INIT('h65)
	) name10289 (
		\u0_w_reg[1][8]/P0001 ,
		_w6316_,
		_w6342_,
		_w10822_
	);
	LUT2 #(
		.INIT('h9)
	) name10290 (
		\u0_w_reg[1][24]/P0002 ,
		_w5909_,
		_w10823_
	);
	LUT2 #(
		.INIT('h9)
	) name10291 (
		\u0_w_reg[1][27]/P0001 ,
		_w6102_,
		_w10824_
	);
	LUT3 #(
		.INIT('hb8)
	) name10292 (
		\key[113]_pad ,
		ld_pad,
		_w10490_,
		_w10825_
	);
	LUT3 #(
		.INIT('hb8)
	) name10293 (
		\key[97]_pad ,
		ld_pad,
		_w10532_,
		_w10826_
	);
	LUT3 #(
		.INIT('hb8)
	) name10294 (
		\key[105]_pad ,
		ld_pad,
		_w10580_,
		_w10827_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10295 (
		\key[81]_pad ,
		ld_pad,
		\u0_w_reg[1][17]/P0001 ,
		_w10490_,
		_w10828_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10296 (
		\key[65]_pad ,
		ld_pad,
		\u0_w_reg[1][1]/P0001 ,
		_w10532_,
		_w10829_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10297 (
		\key[73]_pad ,
		ld_pad,
		\u0_w_reg[1][9]/P0001 ,
		_w10580_,
		_w10830_
	);
	LUT4 #(
		.INIT('h1441)
	) name10298 (
		ld_pad,
		\u0_w_reg[3][17]/P0001 ,
		_w10490_,
		_w10491_,
		_w10831_
	);
	LUT2 #(
		.INIT('h8)
	) name10299 (
		\key[17]_pad ,
		ld_pad,
		_w10832_
	);
	LUT2 #(
		.INIT('he)
	) name10300 (
		_w10831_,
		_w10832_,
		_w10833_
	);
	LUT4 #(
		.INIT('h1441)
	) name10301 (
		ld_pad,
		\u0_w_reg[3][1]/P0001 ,
		_w10532_,
		_w10533_,
		_w10834_
	);
	LUT2 #(
		.INIT('h8)
	) name10302 (
		\key[1]_pad ,
		ld_pad,
		_w10835_
	);
	LUT2 #(
		.INIT('he)
	) name10303 (
		_w10834_,
		_w10835_,
		_w10836_
	);
	LUT4 #(
		.INIT('h1441)
	) name10304 (
		ld_pad,
		\u0_w_reg[3][9]/P0001 ,
		_w10580_,
		_w10581_,
		_w10837_
	);
	LUT2 #(
		.INIT('h8)
	) name10305 (
		\key[9]_pad ,
		ld_pad,
		_w10838_
	);
	LUT2 #(
		.INIT('he)
	) name10306 (
		_w10837_,
		_w10838_,
		_w10839_
	);
	LUT2 #(
		.INIT('h9)
	) name10307 (
		\u0_w_reg[0][19]/P0001 ,
		_w8218_,
		_w10840_
	);
	LUT4 #(
		.INIT('h5655)
	) name10308 (
		\u0_w_reg[3][19]/P0001 ,
		_w2578_,
		_w2565_,
		_w2591_,
		_w10841_
	);
	LUT4 #(
		.INIT('h5655)
	) name10309 (
		\u0_w_reg[2][19]/P0001 ,
		_w4175_,
		_w4161_,
		_w4188_,
		_w10842_
	);
	LUT4 #(
		.INIT('h5655)
	) name10310 (
		\u0_w_reg[1][19]/P0001 ,
		_w6134_,
		_w6120_,
		_w6146_,
		_w10843_
	);
	LUT2 #(
		.INIT('h9)
	) name10311 (
		\u0_w_reg[0][9]/P0001 ,
		_w7865_,
		_w10844_
	);
	LUT4 #(
		.INIT('h5655)
	) name10312 (
		\u0_w_reg[2][9]/P0001 ,
		_w3979_,
		_w3962_,
		_w3995_,
		_w10845_
	);
	LUT4 #(
		.INIT('ha955)
	) name10313 (
		\u0_w_reg[1][9]/P0001 ,
		_w6023_,
		_w6040_,
		_w6052_,
		_w10846_
	);
	LUT2 #(
		.INIT('h9)
	) name10314 (
		\u0_w_reg[0][13]/P0001 ,
		_w7031_,
		_w10847_
	);
	LUT3 #(
		.INIT('h65)
	) name10315 (
		\u0_w_reg[0][21]/P0001 ,
		_w6867_,
		_w6920_,
		_w10848_
	);
	LUT2 #(
		.INIT('h9)
	) name10316 (
		\u0_w_reg[3][13]/P0001 ,
		_w2059_,
		_w10849_
	);
	LUT2 #(
		.INIT('h9)
	) name10317 (
		\u0_w_reg[3][21]/P0001 ,
		_w2002_,
		_w10850_
	);
	LUT4 #(
		.INIT('ha955)
	) name10318 (
		\u0_w_reg[2][13]/P0001 ,
		_w3520_,
		_w3543_,
		_w3556_,
		_w10851_
	);
	LUT3 #(
		.INIT('h65)
	) name10319 (
		\u0_w_reg[2][21]/P0001 ,
		_w775_,
		_w821_,
		_w10852_
	);
	LUT3 #(
		.INIT('h65)
	) name10320 (
		\u0_w_reg[1][13]/P0001 ,
		_w4942_,
		_w5003_,
		_w10853_
	);
	LUT3 #(
		.INIT('h65)
	) name10321 (
		\u0_w_reg[1][21]/P0001 ,
		_w4841_,
		_w4886_,
		_w10854_
	);
	LUT3 #(
		.INIT('hb8)
	) name10322 (
		\key[116]_pad ,
		ld_pad,
		_w10629_,
		_w10855_
	);
	LUT4 #(
		.INIT('h1411)
	) name10323 (
		ld_pad,
		\u0_w_reg[0][4]/P0001 ,
		_w10646_,
		_w10678_,
		_w10856_
	);
	LUT2 #(
		.INIT('h8)
	) name10324 (
		\key[100]_pad ,
		ld_pad,
		_w10857_
	);
	LUT2 #(
		.INIT('he)
	) name10325 (
		_w10856_,
		_w10857_,
		_w10858_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10326 (
		\key[84]_pad ,
		ld_pad,
		\u0_w_reg[1][20]/P0001 ,
		_w10629_,
		_w10859_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10327 (
		\key[68]_pad ,
		ld_pad,
		\u0_w_reg[1][4]/P0001 ,
		_w10679_,
		_w10860_
	);
	LUT4 #(
		.INIT('h8bb8)
	) name10328 (
		\key[20]_pad ,
		ld_pad,
		\u0_w_reg[3][20]/P0001 ,
		_w10630_,
		_w10861_
	);
	LUT4 #(
		.INIT('hb88b)
	) name10329 (
		\key[4]_pad ,
		ld_pad,
		\u0_w_reg[3][4]/P0001 ,
		_w10681_,
		_w10862_
	);
	LUT2 #(
		.INIT('h9)
	) name10330 (
		\u0_w_reg[0][3]/P0001 ,
		_w8309_,
		_w10863_
	);
	LUT4 #(
		.INIT('h5655)
	) name10331 (
		\u0_w_reg[3][9]/P0001 ,
		_w2715_,
		_w2699_,
		_w2731_,
		_w10864_
	);
	LUT2 #(
		.INIT('h9)
	) name10332 (
		\u0_w_reg[0][17]/P0001 ,
		_w8068_,
		_w10865_
	);
	LUT2 #(
		.INIT('h9)
	) name10333 (
		\u0_w_reg[3][17]/P0001 ,
		_w2437_,
		_w10866_
	);
	LUT2 #(
		.INIT('h9)
	) name10334 (
		\u0_w_reg[2][17]/P0001 ,
		_w3745_,
		_w10867_
	);
	LUT4 #(
		.INIT('h5655)
	) name10335 (
		\u0_w_reg[1][17]/P0001 ,
		_w5792_,
		_w5780_,
		_w5810_,
		_w10868_
	);
	LUT2 #(
		.INIT('h9)
	) name10336 (
		\u0_w_reg[0][4]/P0001 ,
		_w7367_,
		_w10869_
	);
	LUT2 #(
		.INIT('h9)
	) name10337 (
		\u0_w_reg[3][12]/P0001 ,
		_w2121_,
		_w10870_
	);
	LUT2 #(
		.INIT('h9)
	) name10338 (
		\u0_w_reg[0][16]/P0001 ,
		_w7655_,
		_w10871_
	);
	LUT2 #(
		.INIT('h9)
	) name10339 (
		\u0_w_reg[3][16]/P0001 ,
		_w2952_,
		_w10872_
	);
	LUT2 #(
		.INIT('h9)
	) name10340 (
		\u0_w_reg[2][16]/P0001 ,
		_w4331_,
		_w10873_
	);
	LUT4 #(
		.INIT('h5655)
	) name10341 (
		\u0_w_reg[1][16]/P0001 ,
		_w6269_,
		_w6283_,
		_w6297_,
		_w10874_
	);
	LUT4 #(
		.INIT('h5655)
	) name10342 (
		\u0_w_reg[0][1]/P0001 ,
		_w7797_,
		_w7782_,
		_w7816_,
		_w10875_
	);
	LUT4 #(
		.INIT('h5655)
	) name10343 (
		\u0_w_reg[0][6]/P0001 ,
		_w8573_,
		_w8587_,
		_w8598_,
		_w10876_
	);
	LUT4 #(
		.INIT('h5655)
	) name10344 (
		\u0_w_reg[0][0]/P0001 ,
		_w7991_,
		_w8004_,
		_w8017_,
		_w10877_
	);
	LUT4 #(
		.INIT('h5655)
	) name10345 (
		\u0_w_reg[0][10]/P0001 ,
		_w8423_,
		_w8413_,
		_w8436_,
		_w10878_
	);
	LUT4 #(
		.INIT('h5655)
	) name10346 (
		\u0_w_reg[0][15]/P0001 ,
		_w7893_,
		_w7880_,
		_w7907_,
		_w10879_
	);
	LUT4 #(
		.INIT('h5655)
	) name10347 (
		\u0_w_reg[0][31]/P0001 ,
		_w8151_,
		_w8138_,
		_w8168_,
		_w10880_
	);
	LUT4 #(
		.INIT('ha955)
	) name10348 (
		\u0_w_reg[3][31]/P0001 ,
		_w1643_,
		_w1667_,
		_w1684_,
		_w10881_
	);
	LUT2 #(
		.INIT('h9)
	) name10349 (
		\u0_w_reg[2][10]/P0001 ,
		_w4466_,
		_w10882_
	);
	LUT2 #(
		.INIT('h9)
	) name10350 (
		\u0_w_reg[2][15]/P0001 ,
		_w3389_,
		_w10883_
	);
	LUT2 #(
		.INIT('h9)
	) name10351 (
		\u0_w_reg[2][31]/P0001 ,
		_w3265_,
		_w10884_
	);
	LUT2 #(
		.INIT('h9)
	) name10352 (
		\u0_w_reg[1][10]/P0001 ,
		_w6507_,
		_w10885_
	);
	LUT4 #(
		.INIT('h5655)
	) name10353 (
		\u0_w_reg[1][15]/P0001 ,
		_w5717_,
		_w5738_,
		_w5757_,
		_w10886_
	);
	LUT3 #(
		.INIT('h65)
	) name10354 (
		\u0_w_reg[1][31]/P0001 ,
		_w5599_,
		_w5642_,
		_w10887_
	);
	LUT2 #(
		.INIT('h9)
	) name10355 (
		\u0_w_reg[0][18]/P0001 ,
		_w8350_,
		_w10888_
	);
	LUT2 #(
		.INIT('h9)
	) name10356 (
		\u0_w_reg[3][18]/P0001 ,
		_w2824_,
		_w10889_
	);
	LUT4 #(
		.INIT('h5655)
	) name10357 (
		\u0_w_reg[2][18]/P0001 ,
		_w4350_,
		_w4361_,
		_w4377_,
		_w10890_
	);
	LUT4 #(
		.INIT('h5655)
	) name10358 (
		\u0_w_reg[1][18]/P0001 ,
		_w6410_,
		_w6396_,
		_w6425_,
		_w10891_
	);
	LUT2 #(
		.INIT('h9)
	) name10359 (
		\u0_w_reg[0][23]/P0001 ,
		_w7706_,
		_w10892_
	);
	LUT2 #(
		.INIT('h9)
	) name10360 (
		\u0_w_reg[3][15]/P0001 ,
		_w1830_,
		_w10893_
	);
	LUT2 #(
		.INIT('h9)
	) name10361 (
		\u0_w_reg[3][23]/P0001 ,
		_w1619_,
		_w10894_
	);
	LUT2 #(
		.INIT('h9)
	) name10362 (
		\u0_w_reg[2][23]/P0001 ,
		_w3324_,
		_w10895_
	);
	LUT2 #(
		.INIT('h9)
	) name10363 (
		\u0_w_reg[1][23]/P0001 ,
		_w5695_,
		_w10896_
	);
	LUT4 #(
		.INIT('h5655)
	) name10364 (
		\u0_w_reg[0][26]/P0001 ,
		_w8377_,
		_w8366_,
		_w8395_,
		_w10897_
	);
	LUT2 #(
		.INIT('h9)
	) name10365 (
		\u0_w_reg[3][26]/P0001 ,
		_w2867_,
		_w10898_
	);
	LUT4 #(
		.INIT('h5655)
	) name10366 (
		\u0_w_reg[2][26]/P0001 ,
		_w4391_,
		_w4403_,
		_w4421_,
		_w10899_
	);
	LUT2 #(
		.INIT('h9)
	) name10367 (
		\u0_w_reg[1][26]/P0001 ,
		_w6469_,
		_w10900_
	);
	LUT4 #(
		.INIT('h5655)
	) name10368 (
		\u0_w_reg[0][7]/P0001 ,
		_w7951_,
		_w7934_,
		_w7970_,
		_w10901_
	);
	LUT2 #(
		.INIT('h9)
	) name10369 (
		\u0_w_reg[0][30]/P0001 ,
		_w7433_,
		_w10902_
	);
	LUT2 #(
		.INIT('h9)
	) name10370 (
		\u0_w_reg[3][30]/P0001 ,
		_w1214_,
		_w10903_
	);
	LUT4 #(
		.INIT('h5655)
	) name10371 (
		\u0_w_reg[2][30]/P0001 ,
		_w3095_,
		_w3117_,
		_w3141_,
		_w10904_
	);
	LUT2 #(
		.INIT('h9)
	) name10372 (
		\u0_w_reg[1][30]/P0001 ,
		_w5454_,
		_w10905_
	);
	LUT4 #(
		.INIT('ha955)
	) name10373 (
		\u0_w_reg[3][10]/P0001 ,
		_w2884_,
		_w2894_,
		_w2908_,
		_w10906_
	);
	LUT4 #(
		.INIT('h5655)
	) name10374 (
		\u0_w_reg[0][14]/P0001 ,
		_w7509_,
		_w7531_,
		_w7550_,
		_w10907_
	);
	LUT4 #(
		.INIT('h5655)
	) name10375 (
		\u0_w_reg[0][22]/P0001 ,
		_w7453_,
		_w7473_,
		_w7490_,
		_w10908_
	);
	LUT2 #(
		.INIT('h9)
	) name10376 (
		\u0_w_reg[3][14]/P0001 ,
		_w1438_,
		_w10909_
	);
	LUT4 #(
		.INIT('h5655)
	) name10377 (
		\u0_w_reg[3][22]/P0001 ,
		_w1261_,
		_w1293_,
		_w1322_,
		_w10910_
	);
	LUT4 #(
		.INIT('h5655)
	) name10378 (
		\u0_w_reg[2][14]/P0001 ,
		_w685_,
		_w714_,
		_w744_,
		_w10911_
	);
	LUT4 #(
		.INIT('h5655)
	) name10379 (
		\u0_w_reg[2][22]/P0001 ,
		_w582_,
		_w612_,
		_w636_,
		_w10912_
	);
	LUT2 #(
		.INIT('h9)
	) name10380 (
		\u0_w_reg[1][14]/P0001 ,
		_w5316_,
		_w10913_
	);
	LUT4 #(
		.INIT('h5655)
	) name10381 (
		\u0_w_reg[1][22]/P0001 ,
		_w5213_,
		_w5229_,
		_w5247_,
		_w10914_
	);
	LUT4 #(
		.INIT('ha955)
	) name10382 (
		\u0_w_reg[0][2]/P0001 ,
		_w8499_,
		_w8511_,
		_w8528_,
		_w10915_
	);
	LUT3 #(
		.INIT('h65)
	) name10383 (
		\u0_w_reg[0][25]/P0001 ,
		_w7725_,
		_w7761_,
		_w10916_
	);
	LUT2 #(
		.INIT('h9)
	) name10384 (
		\u0_w_reg[3][25]/P0001 ,
		_w2489_,
		_w10917_
	);
	LUT2 #(
		.INIT('h9)
	) name10385 (
		\u0_w_reg[2][25]/P0001 ,
		_w3795_,
		_w10918_
	);
	LUT2 #(
		.INIT('h9)
	) name10386 (
		\u0_w_reg[1][25]/P0001 ,
		_w5861_,
		_w10919_
	);
	LUT2 #(
		.INIT('h9)
	) name10387 (
		\u0_w_reg[0][20]/P0001 ,
		_w6737_,
		_w10920_
	);
	LUT2 #(
		.INIT('h9)
	) name10388 (
		\u0_w_reg[3][20]/P0001 ,
		_w1895_,
		_w10921_
	);
	LUT2 #(
		.INIT('h9)
	) name10389 (
		\u0_w_reg[2][20]/P0001 ,
		_w3445_,
		_w10922_
	);
	LUT2 #(
		.INIT('h9)
	) name10390 (
		\u0_w_reg[1][20]/P0001 ,
		_w4691_,
		_w10923_
	);
	LUT2 #(
		.INIT('h9)
	) name10391 (
		\u0_w_reg[0][28]/P0001 ,
		_w6842_,
		_w10924_
	);
	LUT2 #(
		.INIT('h9)
	) name10392 (
		\u0_w_reg[3][28]/P0001 ,
		_w1948_,
		_w10925_
	);
	LUT2 #(
		.INIT('h9)
	) name10393 (
		\u0_w_reg[2][28]/P0001 ,
		_w3496_,
		_w10926_
	);
	LUT2 #(
		.INIT('h9)
	) name10394 (
		\u0_w_reg[1][28]/P0001 ,
		_w4804_,
		_w10927_
	);
	LUT4 #(
		.INIT('h0078)
	) name10395 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		\u0_r0_rcnt_reg[1]/P0001 ,
		\u0_r0_rcnt_reg[2]/P0001 ,
		\u0_r0_rcnt_reg[3]/P0001 ,
		_w10928_
	);
	LUT4 #(
		.INIT('h807f)
	) name10396 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		\u0_r0_rcnt_reg[1]/P0001 ,
		\u0_r0_rcnt_reg[2]/P0001 ,
		\u0_r0_rcnt_reg[3]/P0001 ,
		_w10929_
	);
	LUT4 #(
		.INIT('hfe67)
	) name10397 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		\u0_r0_rcnt_reg[1]/P0001 ,
		\u0_r0_rcnt_reg[2]/P0001 ,
		\u0_r0_rcnt_reg[3]/P0001 ,
		_w10930_
	);
	LUT4 #(
		.INIT('h5455)
	) name10398 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		\u0_r0_rcnt_reg[1]/P0001 ,
		\u0_r0_rcnt_reg[2]/P0001 ,
		\u0_r0_rcnt_reg[3]/P0001 ,
		_w10931_
	);
	LUT3 #(
		.INIT('h01)
	) name10399 (
		ld_pad,
		_w10930_,
		_w10931_,
		_w10932_
	);
	LUT4 #(
		.INIT('haaa8)
	) name10400 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		\u0_r0_rcnt_reg[1]/P0001 ,
		\u0_r0_rcnt_reg[2]/P0001 ,
		\u0_r0_rcnt_reg[3]/P0001 ,
		_w10933_
	);
	LUT3 #(
		.INIT('h01)
	) name10401 (
		ld_pad,
		_w10931_,
		_w10933_,
		_w10934_
	);
	LUT4 #(
		.INIT('haa2a)
	) name10402 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		\u0_r0_rcnt_reg[1]/P0001 ,
		\u0_r0_rcnt_reg[2]/P0001 ,
		\u0_r0_rcnt_reg[3]/P0001 ,
		_w10935_
	);
	LUT4 #(
		.INIT('h5551)
	) name10403 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		\u0_r0_rcnt_reg[1]/P0001 ,
		\u0_r0_rcnt_reg[2]/P0001 ,
		\u0_r0_rcnt_reg[3]/P0001 ,
		_w10936_
	);
	LUT3 #(
		.INIT('h01)
	) name10404 (
		ld_pad,
		_w10936_,
		_w10935_,
		_w10937_
	);
	LUT2 #(
		.INIT('h1)
	) name10405 (
		ld_pad,
		\u0_r0_rcnt_reg[0]/P0001 ,
		_w10938_
	);
	LUT2 #(
		.INIT('h4)
	) name10406 (
		_w10930_,
		_w10938_,
		_w10939_
	);
	LUT4 #(
		.INIT('hfe7e)
	) name10407 (
		\u0_r0_rcnt_reg[0]/P0001 ,
		\u0_r0_rcnt_reg[1]/P0001 ,
		\u0_r0_rcnt_reg[2]/P0001 ,
		\u0_r0_rcnt_reg[3]/P0001 ,
		_w10940_
	);
	LUT2 #(
		.INIT('h1)
	) name10408 (
		ld_pad,
		_w10940_,
		_w10941_
	);
	LUT3 #(
		.INIT('h14)
	) name10409 (
		ld_pad,
		\u0_r0_rcnt_reg[0]/P0001 ,
		\u0_r0_rcnt_reg[1]/P0001 ,
		_w10942_
	);
	LUT3 #(
		.INIT('h10)
	) name10410 (
		ld_pad,
		\u0_r0_rcnt_reg[0]/P0001 ,
		\u0_r0_rcnt_reg[1]/P0001 ,
		_w10943_
	);
	LUT2 #(
		.INIT('h8)
	) name10411 (
		_w10928_,
		_w10943_,
		_w10944_
	);
	LUT3 #(
		.INIT('h04)
	) name10412 (
		ld_pad,
		\u0_r0_rcnt_reg[0]/P0001 ,
		\u0_r0_rcnt_reg[1]/P0001 ,
		_w10945_
	);
	LUT2 #(
		.INIT('h8)
	) name10413 (
		_w10928_,
		_w10945_,
		_w10946_
	);
	LUT4 #(
		.INIT('hfe00)
	) name10414 (
		\dcnt_reg[0]/P0001 ,
		\dcnt_reg[1]/P0001 ,
		\dcnt_reg[2]/P0001 ,
		\dcnt_reg[3]/P0001 ,
		_w10947_
	);
	LUT3 #(
		.INIT('hc8)
	) name10415 (
		ld_pad,
		rst_pad,
		_w10947_,
		_w10948_
	);
	LUT2 #(
		.INIT('h1)
	) name10416 (
		ld_pad,
		_w10929_,
		_w10949_
	);
	LUT4 #(
		.INIT('heaaa)
	) name10417 (
		ld_pad,
		\u0_r0_rcnt_reg[0]/P0001 ,
		\u0_r0_rcnt_reg[1]/P0001 ,
		\u0_r0_rcnt_reg[2]/P0001 ,
		_w10950_
	);
	LUT4 #(
		.INIT('h1e1f)
	) name10418 (
		\dcnt_reg[0]/P0001 ,
		\dcnt_reg[1]/P0001 ,
		\dcnt_reg[2]/P0001 ,
		\dcnt_reg[3]/P0001 ,
		_w10951_
	);
	LUT2 #(
		.INIT('h4)
	) name10419 (
		ld_pad,
		rst_pad,
		_w10952_
	);
	LUT2 #(
		.INIT('h4)
	) name10420 (
		_w10951_,
		_w10952_,
		_w10953_
	);
	LUT2 #(
		.INIT('h1)
	) name10421 (
		\dcnt_reg[2]/P0001 ,
		\dcnt_reg[3]/P0001 ,
		_w10954_
	);
	LUT4 #(
		.INIT('h0001)
	) name10422 (
		\dcnt_reg[0]/P0001 ,
		\dcnt_reg[1]/P0001 ,
		\dcnt_reg[2]/P0001 ,
		\dcnt_reg[3]/P0001 ,
		_w10955_
	);
	LUT4 #(
		.INIT('hc0d0)
	) name10423 (
		\dcnt_reg[0]/P0001 ,
		ld_pad,
		rst_pad,
		_w10955_,
		_w10956_
	);
	LUT2 #(
		.INIT('h6)
	) name10424 (
		\dcnt_reg[0]/P0001 ,
		\dcnt_reg[1]/P0001 ,
		_w10957_
	);
	LUT4 #(
		.INIT('h888c)
	) name10425 (
		ld_pad,
		rst_pad,
		_w10955_,
		_w10957_,
		_w10958_
	);
	LUT4 #(
		.INIT('h1540)
	) name10426 (
		ld_pad,
		\u0_r0_rcnt_reg[0]/P0001 ,
		\u0_r0_rcnt_reg[1]/P0001 ,
		\u0_r0_rcnt_reg[2]/P0001 ,
		_w10959_
	);
	LUT3 #(
		.INIT('h02)
	) name10427 (
		\dcnt_reg[0]/P0001 ,
		\dcnt_reg[1]/P0001 ,
		ld_pad,
		_w10960_
	);
	LUT2 #(
		.INIT('h8)
	) name10428 (
		_w10954_,
		_w10960_,
		_w10961_
	);
	LUT4 #(
		.INIT('h5655)
	) name10429 (
		\u0_w_reg[1][9]/P0001 ,
		_w6370_,
		_w6359_,
		_w6382_,
		_w10962_
	);
	LUT3 #(
		.INIT('h69)
	) name10430 (
		_w5961_,
		_w6012_,
		_w10962_,
		_w10963_
	);
	LUT4 #(
		.INIT('h4114)
	) name10431 (
		\ld_r_reg/P0001 ,
		_w5862_,
		_w6593_,
		_w10963_,
		_w10964_
	);
	LUT3 #(
		.INIT('h28)
	) name10432 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[73]/P0001 ,
		\u0_w_reg[1][9]/P0001 ,
		_w10965_
	);
	LUT2 #(
		.INIT('he)
	) name10433 (
		_w10964_,
		_w10965_,
		_w10966_
	);
	LUT4 #(
		.INIT('h5655)
	) name10434 (
		\u0_w_reg[0][0]/P0001 ,
		_w7951_,
		_w7934_,
		_w7970_,
		_w10967_
	);
	LUT4 #(
		.INIT('h9669)
	) name10435 (
		_w7603_,
		_w7655_,
		_w8123_,
		_w8169_,
		_w10968_
	);
	LUT3 #(
		.INIT('h82)
	) name10436 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[96]/P0001 ,
		\u0_w_reg[0][0]/P0001 ,
		_w10969_
	);
	LUT4 #(
		.INIT('h00eb)
	) name10437 (
		\ld_r_reg/P0001 ,
		_w10967_,
		_w10968_,
		_w10969_,
		_w10970_
	);
	LUT2 #(
		.INIT('h9)
	) name10438 (
		\u0_w_reg[1][0]/P0001 ,
		_w6012_,
		_w10971_
	);
	LUT4 #(
		.INIT('h4114)
	) name10439 (
		\ld_r_reg/P0001 ,
		_w5910_,
		_w6608_,
		_w10971_,
		_w10972_
	);
	LUT3 #(
		.INIT('h82)
	) name10440 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[64]/P0001 ,
		\u0_w_reg[1][0]/P0001 ,
		_w10973_
	);
	LUT2 #(
		.INIT('h1)
	) name10441 (
		_w10972_,
		_w10973_,
		_w10974_
	);
	LUT2 #(
		.INIT('h9)
	) name10442 (
		\u0_w_reg[2][0]/P0001 ,
		_w3949_,
		_w10975_
	);
	LUT4 #(
		.INIT('h9669)
	) name10443 (
		_w3265_,
		_w3841_,
		_w4093_,
		_w4331_,
		_w10976_
	);
	LUT3 #(
		.INIT('h82)
	) name10444 (
		\ld_r_reg/P0001 ,
		\text_in_r_reg[32]/P0001 ,
		\u0_w_reg[2][0]/P0001 ,
		_w10977_
	);
	LUT4 #(
		.INIT('h00eb)
	) name10445 (
		\ld_r_reg/P0001 ,
		_w10975_,
		_w10976_,
		_w10977_,
		_w10978_
	);
	LUT4 #(
		.INIT('h4114)
	) name10446 (
		ld_pad,
		\u0_w_reg[1][24]/P0002 ,
		_w9489_,
		_w9490_,
		_w10979_
	);
	LUT2 #(
		.INIT('h8)
	) name10447 (
		\key[88]_pad ,
		ld_pad,
		_w10980_
	);
	LUT2 #(
		.INIT('he)
	) name10448 (
		_w10979_,
		_w10980_,
		_w10981_
	);
	LUT4 #(
		.INIT('hb88b)
	) name10449 (
		\key[93]_pad ,
		ld_pad,
		_w8777_,
		_w8779_,
		_w10982_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g21/_0_  = _w1043_ ;
	assign \g56610/_0_  = _w1555_ ;
	assign \g56611/_0_  = _w1833_ ;
	assign \g56612/_0_  = _w2064_ ;
	assign \g56613/_0_  = _w2069_ ;
	assign \g56614/_0_  = _w2125_ ;
	assign \g56615/_0_  = _w2130_ ;
	assign \g56616/_0_  = _w2188_ ;
	assign \g56617/_0_  = _w2193_ ;
	assign \g56630/_0_  = _w2493_ ;
	assign \g56631/_0_  = _w2497_ ;
	assign \g56632/_0_  = _w2595_ ;
	assign \g56633/_0_  = _w2645_ ;
	assign \g56634/_0_  = _w2736_ ;
	assign \g56635/_0_  = _w2783_ ;
	assign \g56645/_0_  = _w2913_ ;
	assign \g56646/_0_  = _w2955_ ;
	assign \g56647/_0_  = _w2960_ ;
	assign \g56648/_0_  = _w2964_ ;
	assign \g56649/_0_  = _w2969_ ;
	assign \g56650/_0_  = _w2974_ ;
	assign \g56651/_0_  = _w2979_ ;
	assign \g56652/_0_  = _w3022_ ;
	assign \g56666/_0_  = _w3026_ ;
	assign \g56667/_0_  = _w3031_ ;
	assign \g56668/_0_  = _w3035_ ;
	assign \g56669/_0_  = _w3038_ ;
	assign \g56670/_0_  = _w3042_ ;
	assign \g56671/_0_  = _w3047_ ;
	assign \g56672/_0_  = _w3051_ ;
	assign \g56674/_0_  = _w3056_ ;
	assign \g56675/_0_  = _w3060_ ;
	assign \g56704/_0_  = _w3064_ ;
	assign \g56739/_0_  = _w3065_ ;
	assign \g56743/_0_  = _w3066_ ;
	assign \g56763/_0_  = _w3067_ ;
	assign \g56776/_0_  = _w3068_ ;
	assign \g56812/_0_  = _w3069_ ;
	assign \g56818/_0_  = _w3070_ ;
	assign \g56861/_0_  = _w3071_ ;
	assign \g56874/_0_  = _w3072_ ;
	assign \g56919/_0_  = _w3208_ ;
	assign \g56920/_0_  = _w3392_ ;
	assign \g56921/_0_  = _w3562_ ;
	assign \g56923/_0_  = _w3567_ ;
	assign \g56924/_0_  = _w3620_ ;
	assign \g56925/_0_  = _w3689_ ;
	assign \g56926/_0_  = _w3694_ ;
	assign \g56956/_0_  = _w4000_ ;
	assign \g56957/_0_  = _w4096_ ;
	assign \g56958/_0_  = _w4100_ ;
	assign \g56959/_0_  = _w4192_ ;
	assign \g56960/_0_  = _w4240_ ;
	assign \g56961/_0_  = _w4289_ ;
	assign \g56972/_0_  = _w4336_ ;
	assign \g56973/_0_  = _w4469_ ;
	assign \g56974/_0_  = _w4474_ ;
	assign \g56976/_0_  = _w4478_ ;
	assign \g56977/_0_  = _w4482_ ;
	assign \g56978/_0_  = _w4486_ ;
	assign \g56979/_0_  = _w4490_ ;
	assign \g56980/_0_  = _w4539_ ;
	assign \g57008/_0_  = _w4543_ ;
	assign \g57010/_0_  = _w4547_ ;
	assign \g57011/_0_  = _w4551_ ;
	assign \g57012/_0_  = _w4555_ ;
	assign \g57013/_0_  = _w4559_ ;
	assign \g57014/_0_  = _w4564_ ;
	assign \g57015/_0_  = _w4568_ ;
	assign \g57016/_0_  = _w4572_ ;
	assign \g57017/_0_  = _w4577_ ;
	assign \g57086/_0_  = _w4578_ ;
	assign \g57091/_0_  = _w4579_ ;
	assign \g57114/_0_  = _w4580_ ;
	assign \g57129/_0_  = _w4581_ ;
	assign \g57163/_0_  = _w4582_ ;
	assign \g57171/_0_  = _w4583_ ;
	assign \g57204/_0_  = _w4584_ ;
	assign \g57218/_0_  = _w4585_ ;
	assign \g57262/_0_  = _w5125_ ;
	assign \g57263/_0_  = _w5393_ ;
	assign \g57264/_0_  = _w5459_ ;
	assign \g57265/_0_  = _w5521_ ;
	assign \g57266/_0_  = _w5583_ ;
	assign \g57267/_0_  = _w5588_ ;
	assign \g57268/_0_  = _w5592_ ;
	assign \g57269/_0_  = _w5762_ ;
	assign \g57300/_0_  = _w6058_ ;
	assign \g57301/_0_  = _w6151_ ;
	assign \g57302/_0_  = _w6200_ ;
	assign \g57303/_0_  = _w6204_ ;
	assign \g57304/_0_  = _w6251_ ;
	assign \g57316/_0_  = _w6388_ ;
	assign \g57317/_0_  = _w6510_ ;
	assign \g57319/_0_  = _w6515_ ;
	assign \g57320/_0_  = _w6519_ ;
	assign \g57321/_0_  = _w6526_ ;
	assign \g57322/_0_  = _w6531_ ;
	assign \g57323/_0_  = _w6578_ ;
	assign \g57324/_0_  = _w6583_ ;
	assign \g57350/_0_  = _w6587_ ;
	assign \g57353/_0_  = _w6591_ ;
	assign \g57354/_0_  = _w6597_ ;
	assign \g57355/_0_  = _w6602_ ;
	assign \g57356/_0_  = _w6606_ ;
	assign \g57357/_0_  = _w6611_ ;
	assign \g57358/_0_  = _w6615_ ;
	assign \g57359/_0_  = _w6620_ ;
	assign \g57360/_0_  = _w6625_ ;
	assign \g57427/_0_  = _w6626_ ;
	assign \g57432/_0_  = _w6627_ ;
	assign \g57456/_0_  = _w6628_ ;
	assign \g57471/_0_  = _w6629_ ;
	assign \g57506/_0_  = _w6630_ ;
	assign \g57512/_0_  = _w6631_ ;
	assign \g57540/_0_  = _w6632_ ;
	assign \g57547/_0_  = _w6633_ ;
	assign \g57654/_0_  = _w7150_ ;
	assign \g57655/_0_  = _w7299_ ;
	assign \g57656/_0_  = _w7370_ ;
	assign \g57657/_0_  = _w7374_ ;
	assign \g57658/_0_  = _w7555_ ;
	assign \g57676/_0_  = _w7913_ ;
	assign \g57677/_0_  = _w8072_ ;
	assign \g57678/_0_  = _w8173_ ;
	assign \g57679/_0_  = _w8399_ ;
	assign \g57680/_0_  = _w8483_ ;
	assign \g57681/_0_  = _w8532_ ;
	assign \g57682/_0_  = _w8536_ ;
	assign \g57683/_0_  = _w8540_ ;
	assign \g57684/_0_  = _w8544_ ;
	assign \g57685/_0_  = _w8548_ ;
	assign \g57686/_0_  = _w8552_ ;
	assign \g57687/_0_  = _w8556_ ;
	assign \g57688/_0_  = _w8561_ ;
	assign \g57689/_0_  = _w8603_ ;
	assign \g57690/_0_  = _w8607_ ;
	assign \g57691/_0_  = _w8612_ ;
	assign \g57700/_0_  = _w8616_ ;
	assign \g57701/_0_  = _w8621_ ;
	assign \g57702/_0_  = _w8625_ ;
	assign \g57703/_0_  = _w8629_ ;
	assign \g57704/_0_  = _w8634_ ;
	assign \g57705/_0_  = _w8638_ ;
	assign \g57706/_0_  = _w8643_ ;
	assign \g57707/_0_  = _w8648_ ;
	assign \g57708/_0_  = _w8653_ ;
	assign \g57709/_3_  = _w8778_ ;
	assign \g57710/_3_  = _w8782_ ;
	assign \g57711/_0_  = _w8783_ ;
	assign \g57712/_3_  = _w8902_ ;
	assign \g57715/_3_  = _w8975_ ;
	assign \g57716/_3_  = _w9102_ ;
	assign \g57767/_0_  = _w9107_ ;
	assign \g57768/_3_  = _w9176_ ;
	assign \g57769/_3_  = _w9178_ ;
	assign \g57770/_3_  = _w9182_ ;
	assign \g57771/_3_  = _w9183_ ;
	assign \g57777/_3_  = _w9248_ ;
	assign \g57779/_3_  = _w9360_ ;
	assign \g57804/_3_  = _w9434_ ;
	assign \g57805/_3_  = _w9491_ ;
	assign \g57806/_3_  = _w9547_ ;
	assign \g57807/_3_  = _w9591_ ;
	assign \g57808/_3_  = _w9642_ ;
	assign \g57809/_3_  = _w9644_ ;
	assign \g57810/_3_  = _w9648_ ;
	assign \g57811/_3_  = _w9650_ ;
	assign \g57812/_3_  = _w9653_ ;
	assign \g57813/_3_  = _w9655_ ;
	assign \g57814/_3_  = _w9660_ ;
	assign \g57815/_3_  = _w9663_ ;
	assign \g57816/_0_  = _w9665_ ;
	assign \g57817/_3_  = _w9668_ ;
	assign \g57818/_3_  = _w9669_ ;
	assign \g57819/_3_  = _w9670_ ;
	assign \g57822/_3_  = _w9671_ ;
	assign \g57823/_3_  = _w9672_ ;
	assign \g57824/_3_  = _w9675_ ;
	assign \g57830/_3_  = _w9745_ ;
	assign \g57835/_3_  = _w9746_ ;
	assign \g57836/_3_  = _w9749_ ;
	assign \g57837/_3_  = _w9750_ ;
	assign \g57841/_3_  = _w9751_ ;
	assign \g57842/_3_  = _w9752_ ;
	assign \g57843/_3_  = _w9755_ ;
	assign \g57854/_3_  = _w9806_ ;
	assign \g57855/_3_  = _w9862_ ;
	assign \g57856/_3_  = _w9925_ ;
	assign \g57857/_3_  = _w9978_ ;
	assign \g57858/_3_  = _w10033_ ;
	assign \g57859/_3_  = _w10082_ ;
	assign \g57860/_3_  = _w10126_ ;
	assign \g57861/_3_  = _w10174_ ;
	assign \g57871/_3_  = _w10228_ ;
	assign \g57872/_3_  = _w10287_ ;
	assign \g57874/_3_  = _w10334_ ;
	assign \g57968/_3_  = _w10381_ ;
	assign \g57969/_3_  = _w10383_ ;
	assign \g57970/_3_  = _w10385_ ;
	assign \g57971/_3_  = _w10388_ ;
	assign \g57980/_3_  = _w10439_ ;
	assign \g57983/_3_  = _w10440_ ;
	assign \g57984/_3_  = _w10441_ ;
	assign \g57985/_3_  = _w10444_ ;
	assign \g58012/_3_  = _w10445_ ;
	assign \g58013/_3_  = _w10446_ ;
	assign \g58015/_3_  = _w10449_ ;
	assign \g58057/_3_  = _w10492_ ;
	assign \g58058/_3_  = _w10534_ ;
	assign \g58059/_3_  = _w10582_ ;
	assign \g58189/_3_  = _w10583_ ;
	assign \g58190/_3_  = _w10586_ ;
	assign \g58191/_3_  = _w10633_ ;
	assign \g58192/_3_  = _w10682_ ;
	assign \g58193/_3_  = _w10683_ ;
	assign \g58194/_3_  = _w10735_ ;
	assign \g58195/_3_  = _w10736_ ;
	assign \g58196/_3_  = _w10739_ ;
	assign \g58197/_3_  = _w10741_ ;
	assign \g58224/_3_  = _w10744_ ;
	assign \g58226/_3_  = _w10745_ ;
	assign \g58229/_3_  = _w10746_ ;
	assign \g58255/_3_  = _w10747_ ;
	assign \g58256/_3_  = _w10748_ ;
	assign \g58257/_3_  = _w10749_ ;
	assign \g58258/_3_  = _w10750_ ;
	assign \g58259/_3_  = _w10751_ ;
	assign \g58260/_3_  = _w10752_ ;
	assign \g58261/_3_  = _w10753_ ;
	assign \g58262/_3_  = _w10754_ ;
	assign \g58263/_3_  = _w10755_ ;
	assign \g58264/_3_  = _w10756_ ;
	assign \g58265/_3_  = _w10759_ ;
	assign \g58266/_3_  = _w10762_ ;
	assign \g58267/_3_  = _w10765_ ;
	assign \g58268/_3_  = _w10768_ ;
	assign \g58269/_3_  = _w10769_ ;
	assign \g58270/_0_  = _w10770_ ;
	assign \g58271/_3_  = _w10771_ ;
	assign \g58272/_3_  = _w10772_ ;
	assign \g58273/_3_  = _w10773_ ;
	assign \g58274/_3_  = _w10774_ ;
	assign \g58275/_3_  = _w10775_ ;
	assign \g58276/_3_  = _w10778_ ;
	assign \g58277/_3_  = _w10781_ ;
	assign \g58278/_3_  = _w10784_ ;
	assign \g58279/_3_  = _w10785_ ;
	assign \g58285/_3_  = _w10786_ ;
	assign \g58286/_3_  = _w10787_ ;
	assign \g58288/_3_  = _w10788_ ;
	assign \g58289/_3_  = _w10791_ ;
	assign \g58290/_3_  = _w10792_ ;
	assign \g58292/_3_  = _w10795_ ;
	assign \g58294/_3_  = _w10796_ ;
	assign \g58295/_3_  = _w10797_ ;
	assign \g58297/_3_  = _w10798_ ;
	assign \g58330/_0_  = _w10799_ ;
	assign \g58331/_0_  = _w10800_ ;
	assign \g58332/_0_  = _w10801_ ;
	assign \g58333/_0_  = _w10802_ ;
	assign \g58444/_3_  = _w10803_ ;
	assign \g58445/_3_  = _w10804_ ;
	assign \g58446/_3_  = _w10805_ ;
	assign \g58462/_0_  = _w10806_ ;
	assign \g58506/_0_  = _w10807_ ;
	assign \g58507/_0_  = _w10808_ ;
	assign \g58508/_0_  = _w10809_ ;
	assign \g58509/_0_  = _w10810_ ;
	assign \g58531/_0_  = _w10811_ ;
	assign \g58532/_0_  = _w10812_ ;
	assign \g58533/_0_  = _w10813_ ;
	assign \g58550/_0_  = _w10814_ ;
	assign \g58551/_0_  = _w10815_ ;
	assign \g58552/_0_  = _w10816_ ;
	assign \g58553/_0_  = _w10817_ ;
	assign \g58554/_0_  = _w10818_ ;
	assign \g58555/_0_  = _w10819_ ;
	assign \g58556/_0_  = _w10820_ ;
	assign \g58557/_0_  = _w10821_ ;
	assign \g58558/_0_  = _w10822_ ;
	assign \g58559/_0_  = _w10823_ ;
	assign \g58560/_0_  = _w10824_ ;
	assign \g58600/_3_  = _w10825_ ;
	assign \g58601/_3_  = _w10826_ ;
	assign \g58602/_3_  = _w10827_ ;
	assign \g58603/_3_  = _w10828_ ;
	assign \g58604/_3_  = _w10829_ ;
	assign \g58605/_3_  = _w10830_ ;
	assign \g58606/_3_  = _w10833_ ;
	assign \g58607/_3_  = _w10836_ ;
	assign \g58608/_3_  = _w10839_ ;
	assign \g58611/_0_  = _w10840_ ;
	assign \g58612/_0_  = _w10841_ ;
	assign \g58613/_0_  = _w10842_ ;
	assign \g58614/_0_  = _w10843_ ;
	assign \g58617/_0_  = _w10844_ ;
	assign \g58618/_0_  = _w10845_ ;
	assign \g58619/_0_  = _w10846_ ;
	assign \g58634/_0_  = _w10847_ ;
	assign \g58635/_0_  = _w10848_ ;
	assign \g58636/_0_  = _w10849_ ;
	assign \g58637/_0_  = _w10850_ ;
	assign \g58638/_0_  = _w10851_ ;
	assign \g58639/_0_  = _w10852_ ;
	assign \g58640/_0_  = _w10853_ ;
	assign \g58641/_0_  = _w10854_ ;
	assign \g58829/_3_  = _w10855_ ;
	assign \g58830/_3_  = _w10858_ ;
	assign \g58831/_3_  = _w10859_ ;
	assign \g58832/_3_  = _w10860_ ;
	assign \g58833/_3_  = _w10861_ ;
	assign \g58834/_3_  = _w10862_ ;
	assign \g58835/_0_  = _w10863_ ;
	assign \g58844/_0_  = _w10864_ ;
	assign \g58902/_0_  = _w10865_ ;
	assign \g58903/_0_  = _w10866_ ;
	assign \g58904/_0_  = _w10867_ ;
	assign \g58905/_0_  = _w10868_ ;
	assign \g58910/_0_  = _w10869_ ;
	assign \g58913/_0_  = _w10870_ ;
	assign \g58934/_0_  = _w10871_ ;
	assign \g58935/_0_  = _w10872_ ;
	assign \g58936/_0_  = _w10873_ ;
	assign \g58937/_0_  = _w10874_ ;
	assign \g58938/_0_  = _w10875_ ;
	assign \g58970/_0_  = _w10876_ ;
	assign \g58972/_0_  = _w10877_ ;
	assign \g58994/_0_  = _w10878_ ;
	assign \g58995/_0_  = _w10879_ ;
	assign \g58996/_0_  = _w10880_ ;
	assign \g58997/_0_  = _w10881_ ;
	assign \g58998/_0_  = _w10882_ ;
	assign \g58999/_0_  = _w10883_ ;
	assign \g59000/_0_  = _w10884_ ;
	assign \g59002/_0_  = _w10885_ ;
	assign \g59003/_0_  = _w10886_ ;
	assign \g59004/_0_  = _w10887_ ;
	assign \g59254/_0_  = _w10888_ ;
	assign \g59257/_0_  = _w10889_ ;
	assign \g59258/_0_  = _w10890_ ;
	assign \g59259/_0_  = _w10891_ ;
	assign \g59276/_0_  = _w10892_ ;
	assign \g59277/_0_  = _w10893_ ;
	assign \g59278/_0_  = _w10894_ ;
	assign \g59279/_0_  = _w10895_ ;
	assign \g59280/_0_  = _w10896_ ;
	assign \g59291/_0_  = _w10897_ ;
	assign \g59292/_0_  = _w10898_ ;
	assign \g59293/_0_  = _w10899_ ;
	assign \g59294/_0_  = _w10900_ ;
	assign \g59295/_0_  = _w10901_ ;
	assign \g59308/_0_  = _w10902_ ;
	assign \g59309/_0_  = _w10903_ ;
	assign \g59310/_0_  = _w10904_ ;
	assign \g59311/_0_  = _w10905_ ;
	assign \g59330/_0_  = _w10906_ ;
	assign \g59331/_0_  = _w10907_ ;
	assign \g59332/_0_  = _w10908_ ;
	assign \g59333/_0_  = _w10909_ ;
	assign \g59334/_0_  = _w10910_ ;
	assign \g59335/_0_  = _w10911_ ;
	assign \g59336/_0_  = _w10912_ ;
	assign \g59337/_0_  = _w10913_ ;
	assign \g59338/_0_  = _w10914_ ;
	assign \g59339/_0_  = _w10915_ ;
	assign \g59596/_0_  = _w10916_ ;
	assign \g59597/_0_  = _w10917_ ;
	assign \g59598/_0_  = _w10918_ ;
	assign \g59599/_0_  = _w10919_ ;
	assign \g59625/_0_  = _w10920_ ;
	assign \g59626/_0_  = _w10921_ ;
	assign \g59627/_0_  = _w10922_ ;
	assign \g59628/_0_  = _w10923_ ;
	assign \g59837/_0_  = _w10924_ ;
	assign \g59838/_0_  = _w10925_ ;
	assign \g59839/_0_  = _w10926_ ;
	assign \g59840/_0_  = _w10927_ ;
	assign \g60090/_0_  = _w10932_ ;
	assign \g60320/_0_  = _w10934_ ;
	assign \g60321/_0_  = _w10937_ ;
	assign \g60409/_0_  = _w10939_ ;
	assign \g60539/_0_  = _w10941_ ;
	assign \g60860/_0_  = _w10944_ ;
	assign \g60977/_0_  = _w10946_ ;
	assign \g61012/_0_  = _w10948_ ;
	assign \g61185/_0_  = _w10949_ ;
	assign \g61524/_2_  = _w10950_ ;
	assign \g61776/_0_  = _w10953_ ;
	assign \g61895/_0_  = _w10956_ ;
	assign \g61897/_0_  = _w10958_ ;
	assign \g62220/_0_  = _w10959_ ;
	assign \g65958/_0_  = _w10942_ ;
	assign \g72347/_3_  = _w10961_ ;
	assign \g77848/_0_  = _w10938_ ;
	assign \g85056/_0_  = _w10966_ ;
	assign \sa30_reg[0]/_05_  = _w10970_ ;
	assign \sa31_reg[0]/_05_  = _w10974_ ;
	assign \sa32_reg[0]/_05_  = _w10978_ ;
	assign \u0_w_reg[1][24]/_05_  = _w10981_ ;
	assign \u0_w_reg[1][29]/_05_  = _w10982_ ;
endmodule;