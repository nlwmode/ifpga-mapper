module top( \DataOut_i[0]_pad  , \DataOut_i[1]_pad  , \DataOut_i[2]_pad  , \DataOut_i[3]_pad  , \DataOut_i[4]_pad  , \DataOut_i[5]_pad  , \DataOut_i[6]_pad  , \DataOut_i[7]_pad  , \LineState_o[0]_pad  , \LineState_o[1]_pad  , RxActive_o_pad , RxValid_o_pad , TxValid_i_pad , \i_rx_phy_bit_cnt_reg[0]/NET0131  , \i_rx_phy_bit_cnt_reg[1]/NET0131  , \i_rx_phy_bit_cnt_reg[2]/NET0131  , \i_rx_phy_bit_stuff_err_reg/P0001  , \i_rx_phy_byte_err_reg/P0001  , \i_rx_phy_dpll_state_reg[0]/P0001  , \i_rx_phy_dpll_state_reg[1]/NET0131  , \i_rx_phy_fs_ce_reg/P0001  , \i_rx_phy_fs_state_reg[0]/NET0131  , \i_rx_phy_fs_state_reg[1]/P0001  , \i_rx_phy_fs_state_reg[2]/NET0131  , \i_rx_phy_one_cnt_reg[0]/NET0131  , \i_rx_phy_one_cnt_reg[1]/NET0131  , \i_rx_phy_one_cnt_reg[2]/NET0131  , \i_rx_phy_rx_en_reg/NET0131  , \i_rx_phy_rx_valid1_reg/P0001  , \i_rx_phy_rx_valid_r_reg/P0001  , \i_rx_phy_rxd_r_reg/NET0131  , \i_rx_phy_rxd_s0_reg/P0001  , \i_rx_phy_rxd_s1_reg/P0001  , \i_rx_phy_rxd_s_reg/P0001  , \i_rx_phy_rxdn_s0_reg/P0001  , \i_rx_phy_rxdn_s_r_reg/P0001  , \i_rx_phy_rxdn_s_reg/NET0131  , \i_rx_phy_rxdp_s0_reg/P0001  , \i_rx_phy_rxdp_s_r_reg/P0001  , \i_rx_phy_rxdp_s_reg/NET0131  , \i_rx_phy_sd_nrzi_reg/NET0131  , \i_rx_phy_sd_r_reg/NET0131  , \i_rx_phy_se0_r_reg/P0001  , \i_rx_phy_se0_s_reg/NET0131  , \i_rx_phy_shift_en_reg/NET0131  , \i_rx_phy_sync_err_reg/P0001  , \i_tx_phy_append_eop_reg/P0001  , \i_tx_phy_append_eop_sync1_reg/P0001  , \i_tx_phy_append_eop_sync2_reg/P0001  , \i_tx_phy_append_eop_sync3_reg/NET0131  , \i_tx_phy_append_eop_sync4_reg/P0001  , \i_tx_phy_bit_cnt_reg[0]/NET0131  , \i_tx_phy_bit_cnt_reg[1]/NET0131  , \i_tx_phy_bit_cnt_reg[2]/P0001  , \i_tx_phy_data_done_reg/NET0131  , \i_tx_phy_hold_reg_d_reg[0]/P0001  , \i_tx_phy_hold_reg_d_reg[1]/P0001  , \i_tx_phy_hold_reg_d_reg[2]/P0001  , \i_tx_phy_hold_reg_d_reg[3]/P0001  , \i_tx_phy_hold_reg_d_reg[4]/P0001  , \i_tx_phy_hold_reg_d_reg[5]/P0001  , \i_tx_phy_hold_reg_d_reg[6]/P0001  , \i_tx_phy_hold_reg_d_reg[7]/P0001  , \i_tx_phy_hold_reg_reg[0]/P0001  , \i_tx_phy_hold_reg_reg[1]/P0001  , \i_tx_phy_hold_reg_reg[2]/P0001  , \i_tx_phy_hold_reg_reg[3]/P0001  , \i_tx_phy_hold_reg_reg[4]/P0001  , \i_tx_phy_hold_reg_reg[5]/P0001  , \i_tx_phy_hold_reg_reg[6]/P0001  , \i_tx_phy_hold_reg_reg[7]/P0001  , \i_tx_phy_ld_data_reg/NET0131  , \i_tx_phy_one_cnt_reg[0]/NET0131  , \i_tx_phy_one_cnt_reg[1]/NET0131  , \i_tx_phy_one_cnt_reg[2]/NET0131  , \i_tx_phy_sd_bs_o_reg/NET0131  , \i_tx_phy_sd_nrzi_o_reg/NET0131  , \i_tx_phy_sd_raw_o_reg/NET0131  , \i_tx_phy_sft_done_r_reg/NET0131  , \i_tx_phy_sft_done_reg/NET0131  , \i_tx_phy_state_reg[0]/P0001  , \i_tx_phy_state_reg[1]/P0001  , \i_tx_phy_state_reg[2]/NET0131  , \i_tx_phy_tx_ip_reg/P0001  , \i_tx_phy_tx_ip_sync_reg/P0001  , \i_tx_phy_txoe_r1_reg/P0001  , \i_tx_phy_txoe_r2_reg/P0001  , phy_tx_mode_pad , \rst_cnt_reg[0]/NET0131  , \rst_cnt_reg[1]/NET0131  , \rst_cnt_reg[2]/NET0131  , \rst_cnt_reg[3]/NET0131  , \rst_cnt_reg[4]/NET0131  , rst_pad , txdn_pad , txdp_pad , txoe_pad , usb_rst_pad , RxError_o_pad , \_al_n0  , \_al_n1  , \g1661/_0_  , \g1680/_0_  , \g1695/_0_  , \g1703/_1_  , \g1707/_0_  , \g1725/_0_  , \g1728/_0_  , \g1729/_0_  , \g1736/_0_  , \g1737/_0_  , \g1738/_0_  , \g1739/_0_  , \g1740/_0_  , \g1741/_0_  , \g1742/_0_  , \g1743/_0_  , \g1747/_3_  , \g1748/_0_  , \g1757/_0_  , \g1758/_0_  , \g1763/_0_  , \g1764/_0_  , \g1811/_0_  , \g1812/_0_  , \g1815/_0_  , \g1816/_0_  , \g1820/_1_  , \g1821/_0_  , \g1837/_0_  , \g1838/_0_  , \g1841/_0_  , \g1842/_0_  , \g1843/_0_  , \g1844/_0_  , \g1845/_0_  , \g1846/_0_  , \g1848/_0_  , \g1851/_0_  , \g1852/_0_  , \g1853/_0_  , \g1857/_0_  , \g1858/_0_  , \g1865/_0_  , \g1869/_0_  , \g1871/_0_  , \g1872/_0_  , \g1873/_0_  , \g1876/_0_  , \g1878/_0_  , \g1897/_1_  , \g1901/_0_  , \g1904/_0_  , \g1928/_0_  , \g1936/_3_  , \g1961/_0_  , \g1962/_0_  , \g1963/_0_  , \g1966/_0_  , \g1967/_0_  , \g1968/_0_  , \g1975/_0_  , \g1980/_0_  , \g2055/_0_  , \g2112/_0_  , \g2411/_2_  , \g2463/_0_  , \g2501/_0_  , \g2620/_0_  , \g2650/_0_  , \g2657/_0_  , \g2671/_0_  , \i_rx_phy_sd_r_reg/NET0131_reg_syn_3  );
  input \DataOut_i[0]_pad  ;
  input \DataOut_i[1]_pad  ;
  input \DataOut_i[2]_pad  ;
  input \DataOut_i[3]_pad  ;
  input \DataOut_i[4]_pad  ;
  input \DataOut_i[5]_pad  ;
  input \DataOut_i[6]_pad  ;
  input \DataOut_i[7]_pad  ;
  input \LineState_o[0]_pad  ;
  input \LineState_o[1]_pad  ;
  input RxActive_o_pad ;
  input RxValid_o_pad ;
  input TxValid_i_pad ;
  input \i_rx_phy_bit_cnt_reg[0]/NET0131  ;
  input \i_rx_phy_bit_cnt_reg[1]/NET0131  ;
  input \i_rx_phy_bit_cnt_reg[2]/NET0131  ;
  input \i_rx_phy_bit_stuff_err_reg/P0001  ;
  input \i_rx_phy_byte_err_reg/P0001  ;
  input \i_rx_phy_dpll_state_reg[0]/P0001  ;
  input \i_rx_phy_dpll_state_reg[1]/NET0131  ;
  input \i_rx_phy_fs_ce_reg/P0001  ;
  input \i_rx_phy_fs_state_reg[0]/NET0131  ;
  input \i_rx_phy_fs_state_reg[1]/P0001  ;
  input \i_rx_phy_fs_state_reg[2]/NET0131  ;
  input \i_rx_phy_one_cnt_reg[0]/NET0131  ;
  input \i_rx_phy_one_cnt_reg[1]/NET0131  ;
  input \i_rx_phy_one_cnt_reg[2]/NET0131  ;
  input \i_rx_phy_rx_en_reg/NET0131  ;
  input \i_rx_phy_rx_valid1_reg/P0001  ;
  input \i_rx_phy_rx_valid_r_reg/P0001  ;
  input \i_rx_phy_rxd_r_reg/NET0131  ;
  input \i_rx_phy_rxd_s0_reg/P0001  ;
  input \i_rx_phy_rxd_s1_reg/P0001  ;
  input \i_rx_phy_rxd_s_reg/P0001  ;
  input \i_rx_phy_rxdn_s0_reg/P0001  ;
  input \i_rx_phy_rxdn_s_r_reg/P0001  ;
  input \i_rx_phy_rxdn_s_reg/NET0131  ;
  input \i_rx_phy_rxdp_s0_reg/P0001  ;
  input \i_rx_phy_rxdp_s_r_reg/P0001  ;
  input \i_rx_phy_rxdp_s_reg/NET0131  ;
  input \i_rx_phy_sd_nrzi_reg/NET0131  ;
  input \i_rx_phy_sd_r_reg/NET0131  ;
  input \i_rx_phy_se0_r_reg/P0001  ;
  input \i_rx_phy_se0_s_reg/NET0131  ;
  input \i_rx_phy_shift_en_reg/NET0131  ;
  input \i_rx_phy_sync_err_reg/P0001  ;
  input \i_tx_phy_append_eop_reg/P0001  ;
  input \i_tx_phy_append_eop_sync1_reg/P0001  ;
  input \i_tx_phy_append_eop_sync2_reg/P0001  ;
  input \i_tx_phy_append_eop_sync3_reg/NET0131  ;
  input \i_tx_phy_append_eop_sync4_reg/P0001  ;
  input \i_tx_phy_bit_cnt_reg[0]/NET0131  ;
  input \i_tx_phy_bit_cnt_reg[1]/NET0131  ;
  input \i_tx_phy_bit_cnt_reg[2]/P0001  ;
  input \i_tx_phy_data_done_reg/NET0131  ;
  input \i_tx_phy_hold_reg_d_reg[0]/P0001  ;
  input \i_tx_phy_hold_reg_d_reg[1]/P0001  ;
  input \i_tx_phy_hold_reg_d_reg[2]/P0001  ;
  input \i_tx_phy_hold_reg_d_reg[3]/P0001  ;
  input \i_tx_phy_hold_reg_d_reg[4]/P0001  ;
  input \i_tx_phy_hold_reg_d_reg[5]/P0001  ;
  input \i_tx_phy_hold_reg_d_reg[6]/P0001  ;
  input \i_tx_phy_hold_reg_d_reg[7]/P0001  ;
  input \i_tx_phy_hold_reg_reg[0]/P0001  ;
  input \i_tx_phy_hold_reg_reg[1]/P0001  ;
  input \i_tx_phy_hold_reg_reg[2]/P0001  ;
  input \i_tx_phy_hold_reg_reg[3]/P0001  ;
  input \i_tx_phy_hold_reg_reg[4]/P0001  ;
  input \i_tx_phy_hold_reg_reg[5]/P0001  ;
  input \i_tx_phy_hold_reg_reg[6]/P0001  ;
  input \i_tx_phy_hold_reg_reg[7]/P0001  ;
  input \i_tx_phy_ld_data_reg/NET0131  ;
  input \i_tx_phy_one_cnt_reg[0]/NET0131  ;
  input \i_tx_phy_one_cnt_reg[1]/NET0131  ;
  input \i_tx_phy_one_cnt_reg[2]/NET0131  ;
  input \i_tx_phy_sd_bs_o_reg/NET0131  ;
  input \i_tx_phy_sd_nrzi_o_reg/NET0131  ;
  input \i_tx_phy_sd_raw_o_reg/NET0131  ;
  input \i_tx_phy_sft_done_r_reg/NET0131  ;
  input \i_tx_phy_sft_done_reg/NET0131  ;
  input \i_tx_phy_state_reg[0]/P0001  ;
  input \i_tx_phy_state_reg[1]/P0001  ;
  input \i_tx_phy_state_reg[2]/NET0131  ;
  input \i_tx_phy_tx_ip_reg/P0001  ;
  input \i_tx_phy_tx_ip_sync_reg/P0001  ;
  input \i_tx_phy_txoe_r1_reg/P0001  ;
  input \i_tx_phy_txoe_r2_reg/P0001  ;
  input phy_tx_mode_pad ;
  input \rst_cnt_reg[0]/NET0131  ;
  input \rst_cnt_reg[1]/NET0131  ;
  input \rst_cnt_reg[2]/NET0131  ;
  input \rst_cnt_reg[3]/NET0131  ;
  input \rst_cnt_reg[4]/NET0131  ;
  input rst_pad ;
  input txdn_pad ;
  input txdp_pad ;
  input txoe_pad ;
  input usb_rst_pad ;
  output RxError_o_pad ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1661/_0_  ;
  output \g1680/_0_  ;
  output \g1695/_0_  ;
  output \g1703/_1_  ;
  output \g1707/_0_  ;
  output \g1725/_0_  ;
  output \g1728/_0_  ;
  output \g1729/_0_  ;
  output \g1736/_0_  ;
  output \g1737/_0_  ;
  output \g1738/_0_  ;
  output \g1739/_0_  ;
  output \g1740/_0_  ;
  output \g1741/_0_  ;
  output \g1742/_0_  ;
  output \g1743/_0_  ;
  output \g1747/_3_  ;
  output \g1748/_0_  ;
  output \g1757/_0_  ;
  output \g1758/_0_  ;
  output \g1763/_0_  ;
  output \g1764/_0_  ;
  output \g1811/_0_  ;
  output \g1812/_0_  ;
  output \g1815/_0_  ;
  output \g1816/_0_  ;
  output \g1820/_1_  ;
  output \g1821/_0_  ;
  output \g1837/_0_  ;
  output \g1838/_0_  ;
  output \g1841/_0_  ;
  output \g1842/_0_  ;
  output \g1843/_0_  ;
  output \g1844/_0_  ;
  output \g1845/_0_  ;
  output \g1846/_0_  ;
  output \g1848/_0_  ;
  output \g1851/_0_  ;
  output \g1852/_0_  ;
  output \g1853/_0_  ;
  output \g1857/_0_  ;
  output \g1858/_0_  ;
  output \g1865/_0_  ;
  output \g1869/_0_  ;
  output \g1871/_0_  ;
  output \g1872/_0_  ;
  output \g1873/_0_  ;
  output \g1876/_0_  ;
  output \g1878/_0_  ;
  output \g1897/_1_  ;
  output \g1901/_0_  ;
  output \g1904/_0_  ;
  output \g1928/_0_  ;
  output \g1936/_3_  ;
  output \g1961/_0_  ;
  output \g1962/_0_  ;
  output \g1963/_0_  ;
  output \g1966/_0_  ;
  output \g1967/_0_  ;
  output \g1968/_0_  ;
  output \g1975/_0_  ;
  output \g1980/_0_  ;
  output \g2055/_0_  ;
  output \g2112/_0_  ;
  output \g2411/_2_  ;
  output \g2463/_0_  ;
  output \g2501/_0_  ;
  output \g2620/_0_  ;
  output \g2650/_0_  ;
  output \g2657/_0_  ;
  output \g2671/_0_  ;
  output \i_rx_phy_sd_r_reg/NET0131_reg_syn_3  ;
  wire n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 ;
  assign n99 = ~\i_rx_phy_bit_stuff_err_reg/P0001  & ~\i_rx_phy_byte_err_reg/P0001  ;
  assign n100 = ~\i_rx_phy_sync_err_reg/P0001  & n99 ;
  assign n101 = \i_rx_phy_rxdn_s_reg/NET0131  & ~\i_rx_phy_rxdp_s_reg/NET0131  ;
  assign n102 = \i_rx_phy_rx_en_reg/NET0131  & n101 ;
  assign n103 = ~\i_rx_phy_fs_state_reg[0]/NET0131  & n102 ;
  assign n104 = ~\i_rx_phy_rxdn_s_reg/NET0131  & ~\i_rx_phy_rxdp_s_reg/NET0131  ;
  assign n105 = \i_rx_phy_fs_ce_reg/P0001  & ~n104 ;
  assign n106 = ~RxActive_o_pad & ~\i_rx_phy_se0_s_reg/NET0131  ;
  assign n107 = n105 & n106 ;
  assign n108 = ~n103 & n107 ;
  assign n109 = \i_rx_phy_fs_state_reg[1]/P0001  & ~n108 ;
  assign n110 = \i_rx_phy_rx_en_reg/NET0131  & ~\i_rx_phy_rxdn_s_reg/NET0131  ;
  assign n111 = \i_rx_phy_rxdp_s_reg/NET0131  & n110 ;
  assign n112 = \i_rx_phy_fs_state_reg[0]/NET0131  & ~\i_rx_phy_fs_state_reg[1]/P0001  ;
  assign n113 = n111 & n112 ;
  assign n114 = n107 & n113 ;
  assign n115 = ~n109 & ~n114 ;
  assign n116 = rst_pad & ~n115 ;
  assign n117 = \i_rx_phy_fs_ce_reg/P0001  & ~usb_rst_pad ;
  assign n118 = \rst_cnt_reg[0]/NET0131  & n117 ;
  assign n119 = \rst_cnt_reg[1]/NET0131  & n118 ;
  assign n120 = \rst_cnt_reg[2]/NET0131  & n119 ;
  assign n121 = ~\rst_cnt_reg[3]/NET0131  & ~n120 ;
  assign n122 = ~\LineState_o[0]_pad  & ~\LineState_o[1]_pad  ;
  assign n123 = rst_pad & n122 ;
  assign n124 = \rst_cnt_reg[2]/NET0131  & \rst_cnt_reg[3]/NET0131  ;
  assign n125 = n119 & n124 ;
  assign n126 = n123 & ~n125 ;
  assign n127 = ~n121 & n126 ;
  assign n128 = ~\i_tx_phy_state_reg[0]/P0001  & ~\i_tx_phy_state_reg[1]/P0001  ;
  assign n129 = \i_tx_phy_state_reg[2]/NET0131  & n128 ;
  assign n130 = \i_rx_phy_fs_ce_reg/P0001  & ~\i_tx_phy_append_eop_sync3_reg/NET0131  ;
  assign n131 = n129 & n130 ;
  assign n137 = TxValid_i_pad & ~\i_tx_phy_state_reg[2]/NET0131  ;
  assign n138 = n128 & n137 ;
  assign n147 = ~n131 & ~n138 ;
  assign n132 = ~\i_tx_phy_sft_done_r_reg/NET0131  & \i_tx_phy_sft_done_reg/NET0131  ;
  assign n143 = ~\i_tx_phy_state_reg[2]/NET0131  & n132 ;
  assign n142 = \i_tx_phy_state_reg[0]/P0001  & ~\i_tx_phy_state_reg[1]/P0001  ;
  assign n144 = \i_rx_phy_fs_ce_reg/P0001  & \i_tx_phy_state_reg[2]/NET0131  ;
  assign n145 = n142 & ~n144 ;
  assign n146 = ~n143 & n145 ;
  assign n133 = ~\i_tx_phy_state_reg[0]/P0001  & \i_tx_phy_state_reg[1]/P0001  ;
  assign n134 = ~\i_tx_phy_state_reg[2]/NET0131  & n133 ;
  assign n135 = ~\i_tx_phy_data_done_reg/NET0131  & n132 ;
  assign n136 = n134 & n135 ;
  assign n139 = \i_tx_phy_state_reg[0]/P0001  & \i_tx_phy_state_reg[1]/P0001  ;
  assign n140 = ~\i_tx_phy_state_reg[2]/NET0131  & n139 ;
  assign n141 = ~\i_tx_phy_append_eop_sync3_reg/NET0131  & n140 ;
  assign n148 = ~n136 & ~n141 ;
  assign n149 = ~n146 & n148 ;
  assign n150 = n147 & n149 ;
  assign n151 = rst_pad & ~n150 ;
  assign n153 = \rst_cnt_reg[4]/NET0131  & n125 ;
  assign n152 = ~\rst_cnt_reg[4]/NET0131  & ~n125 ;
  assign n154 = n123 & ~n152 ;
  assign n155 = ~n153 & n154 ;
  assign n156 = ~\i_rx_phy_bit_cnt_reg[1]/NET0131  & ~\i_rx_phy_bit_cnt_reg[2]/NET0131  ;
  assign n157 = RxActive_o_pad & ~\i_rx_phy_se0_r_reg/P0001  ;
  assign n158 = n104 & n157 ;
  assign n159 = ~n156 & n158 ;
  assign n160 = ~\rst_cnt_reg[2]/NET0131  & ~n119 ;
  assign n161 = ~n120 & n123 ;
  assign n162 = ~n160 & n161 ;
  assign n163 = \i_tx_phy_hold_reg_reg[7]/P0001  & ~\i_tx_phy_ld_data_reg/NET0131  ;
  assign n164 = \DataOut_i[7]_pad  & \i_tx_phy_ld_data_reg/NET0131  ;
  assign n165 = ~n163 & ~n164 ;
  assign n166 = ~n138 & n165 ;
  assign n168 = ~\i_rx_phy_one_cnt_reg[0]/NET0131  & \i_rx_phy_one_cnt_reg[1]/NET0131  ;
  assign n169 = \i_rx_phy_one_cnt_reg[2]/NET0131  & n168 ;
  assign n170 = \i_rx_phy_fs_ce_reg/P0001  & ~n169 ;
  assign n171 = \i_rx_phy_bit_cnt_reg[0]/NET0131  & n170 ;
  assign n172 = \i_rx_phy_bit_cnt_reg[1]/NET0131  & n171 ;
  assign n174 = ~\i_rx_phy_bit_cnt_reg[2]/NET0131  & ~n172 ;
  assign n167 = \i_rx_phy_shift_en_reg/NET0131  & rst_pad ;
  assign n173 = \i_rx_phy_bit_cnt_reg[2]/NET0131  & n172 ;
  assign n175 = n167 & ~n173 ;
  assign n176 = ~n174 & n175 ;
  assign n192 = \i_tx_phy_bit_cnt_reg[1]/NET0131  & ~\i_tx_phy_hold_reg_d_reg[7]/P0001  ;
  assign n191 = ~\i_tx_phy_bit_cnt_reg[1]/NET0131  & ~\i_tx_phy_hold_reg_d_reg[5]/P0001  ;
  assign n193 = \i_tx_phy_bit_cnt_reg[0]/NET0131  & ~n191 ;
  assign n194 = ~n192 & n193 ;
  assign n188 = \i_tx_phy_bit_cnt_reg[1]/NET0131  & ~\i_tx_phy_hold_reg_d_reg[6]/P0001  ;
  assign n187 = ~\i_tx_phy_bit_cnt_reg[1]/NET0131  & ~\i_tx_phy_hold_reg_d_reg[4]/P0001  ;
  assign n189 = ~\i_tx_phy_bit_cnt_reg[0]/NET0131  & ~n187 ;
  assign n190 = ~n188 & n189 ;
  assign n195 = \i_tx_phy_bit_cnt_reg[2]/P0001  & ~n190 ;
  assign n196 = ~n194 & n195 ;
  assign n182 = \i_tx_phy_bit_cnt_reg[0]/NET0131  & ~\i_tx_phy_hold_reg_d_reg[1]/P0001  ;
  assign n181 = ~\i_tx_phy_bit_cnt_reg[0]/NET0131  & ~\i_tx_phy_hold_reg_d_reg[0]/P0001  ;
  assign n183 = ~\i_tx_phy_bit_cnt_reg[1]/NET0131  & ~n181 ;
  assign n184 = ~n182 & n183 ;
  assign n178 = \i_tx_phy_bit_cnt_reg[0]/NET0131  & ~\i_tx_phy_hold_reg_d_reg[3]/P0001  ;
  assign n177 = ~\i_tx_phy_bit_cnt_reg[0]/NET0131  & ~\i_tx_phy_hold_reg_d_reg[2]/P0001  ;
  assign n179 = \i_tx_phy_bit_cnt_reg[1]/NET0131  & ~n177 ;
  assign n180 = ~n178 & n179 ;
  assign n185 = ~\i_tx_phy_bit_cnt_reg[2]/P0001  & ~n180 ;
  assign n186 = ~n184 & n185 ;
  assign n197 = \i_tx_phy_tx_ip_sync_reg/P0001  & ~n186 ;
  assign n198 = ~n196 & n197 ;
  assign n199 = ~\i_tx_phy_hold_reg_reg[0]/P0001  & ~\i_tx_phy_ld_data_reg/NET0131  ;
  assign n200 = ~\DataOut_i[0]_pad  & \i_tx_phy_ld_data_reg/NET0131  ;
  assign n201 = ~n199 & ~n200 ;
  assign n202 = ~n138 & n201 ;
  assign n203 = ~\i_tx_phy_hold_reg_reg[1]/P0001  & ~\i_tx_phy_ld_data_reg/NET0131  ;
  assign n204 = ~\DataOut_i[1]_pad  & \i_tx_phy_ld_data_reg/NET0131  ;
  assign n205 = ~n203 & ~n204 ;
  assign n206 = ~n138 & n205 ;
  assign n207 = ~\i_tx_phy_hold_reg_reg[2]/P0001  & ~\i_tx_phy_ld_data_reg/NET0131  ;
  assign n208 = ~\DataOut_i[2]_pad  & \i_tx_phy_ld_data_reg/NET0131  ;
  assign n209 = ~n207 & ~n208 ;
  assign n210 = ~n138 & n209 ;
  assign n211 = ~\i_tx_phy_hold_reg_reg[3]/P0001  & ~\i_tx_phy_ld_data_reg/NET0131  ;
  assign n212 = ~\DataOut_i[3]_pad  & \i_tx_phy_ld_data_reg/NET0131  ;
  assign n213 = ~n211 & ~n212 ;
  assign n214 = ~n138 & n213 ;
  assign n215 = ~\i_tx_phy_hold_reg_reg[4]/P0001  & ~\i_tx_phy_ld_data_reg/NET0131  ;
  assign n216 = ~\DataOut_i[4]_pad  & \i_tx_phy_ld_data_reg/NET0131  ;
  assign n217 = ~n215 & ~n216 ;
  assign n218 = ~n138 & n217 ;
  assign n219 = ~\i_tx_phy_hold_reg_reg[5]/P0001  & ~\i_tx_phy_ld_data_reg/NET0131  ;
  assign n220 = ~\DataOut_i[5]_pad  & \i_tx_phy_ld_data_reg/NET0131  ;
  assign n221 = ~n219 & ~n220 ;
  assign n222 = ~n138 & n221 ;
  assign n223 = ~\i_tx_phy_hold_reg_reg[6]/P0001  & ~\i_tx_phy_ld_data_reg/NET0131  ;
  assign n224 = ~\DataOut_i[6]_pad  & \i_tx_phy_ld_data_reg/NET0131  ;
  assign n225 = ~n223 & ~n224 ;
  assign n226 = ~n138 & n225 ;
  assign n227 = RxActive_o_pad & \i_rx_phy_fs_ce_reg/P0001  ;
  assign n228 = \i_rx_phy_sd_nrzi_reg/NET0131  & ~n104 ;
  assign n229 = n227 & n228 ;
  assign n230 = n169 & n229 ;
  assign n231 = ~\i_rx_phy_fs_ce_reg/P0001  & ~\i_rx_phy_se0_s_reg/NET0131  ;
  assign n232 = ~n105 & ~n231 ;
  assign n233 = n142 & n143 ;
  assign n234 = ~n134 & ~n233 ;
  assign n235 = ~n141 & n234 ;
  assign n236 = rst_pad & ~n235 ;
  assign n237 = \i_tx_phy_append_eop_sync3_reg/NET0131  & n140 ;
  assign n238 = ~\i_rx_phy_fs_ce_reg/P0001  & \i_tx_phy_state_reg[2]/NET0131  ;
  assign n239 = n142 & n238 ;
  assign n240 = ~n129 & ~n239 ;
  assign n241 = ~n237 & n240 ;
  assign n242 = rst_pad & ~n241 ;
  assign n243 = \i_tx_phy_one_cnt_reg[0]/NET0131  & \i_tx_phy_one_cnt_reg[1]/NET0131  ;
  assign n244 = ~\i_tx_phy_one_cnt_reg[0]/NET0131  & \i_tx_phy_one_cnt_reg[1]/NET0131  ;
  assign n245 = \i_tx_phy_one_cnt_reg[2]/NET0131  & n244 ;
  assign n246 = \i_rx_phy_fs_ce_reg/P0001  & ~n245 ;
  assign n247 = \i_tx_phy_sd_raw_o_reg/NET0131  & n246 ;
  assign n251 = ~n243 & n247 ;
  assign n252 = \i_rx_phy_fs_ce_reg/P0001  & \i_tx_phy_one_cnt_reg[2]/NET0131  ;
  assign n253 = ~n251 & n252 ;
  assign n248 = n243 & n247 ;
  assign n249 = ~\i_tx_phy_one_cnt_reg[2]/NET0131  & ~n248 ;
  assign n250 = \i_tx_phy_tx_ip_sync_reg/P0001  & rst_pad ;
  assign n254 = ~n249 & n250 ;
  assign n255 = ~n253 & n254 ;
  assign n256 = \i_rx_phy_rx_valid1_reg/P0001  & ~n170 ;
  assign n257 = ~n173 & ~n256 ;
  assign n258 = rst_pad & ~n257 ;
  assign n259 = \i_tx_phy_bit_cnt_reg[0]/NET0131  & n246 ;
  assign n260 = \i_tx_phy_bit_cnt_reg[1]/NET0131  & n259 ;
  assign n262 = \i_tx_phy_bit_cnt_reg[2]/P0001  & n260 ;
  assign n261 = ~\i_tx_phy_bit_cnt_reg[2]/P0001  & ~n260 ;
  assign n263 = n250 & ~n261 ;
  assign n264 = ~n262 & n263 ;
  assign n265 = ~\i_rx_phy_fs_ce_reg/P0001  & \i_rx_phy_one_cnt_reg[1]/NET0131  ;
  assign n266 = ~\i_rx_phy_one_cnt_reg[0]/NET0131  & ~\i_rx_phy_one_cnt_reg[1]/NET0131  ;
  assign n267 = \i_rx_phy_sd_nrzi_reg/NET0131  & n170 ;
  assign n268 = \i_rx_phy_one_cnt_reg[0]/NET0131  & \i_rx_phy_one_cnt_reg[1]/NET0131  ;
  assign n269 = n267 & ~n268 ;
  assign n270 = ~n266 & n269 ;
  assign n271 = ~n265 & ~n270 ;
  assign n272 = n167 & ~n271 ;
  assign n273 = ~\i_rx_phy_fs_ce_reg/P0001  & \i_tx_phy_one_cnt_reg[1]/NET0131  ;
  assign n274 = ~\i_tx_phy_one_cnt_reg[0]/NET0131  & ~\i_tx_phy_one_cnt_reg[1]/NET0131  ;
  assign n275 = n251 & ~n274 ;
  assign n276 = ~n273 & ~n275 ;
  assign n277 = n250 & ~n276 ;
  assign n278 = \i_rx_phy_rxd_r_reg/NET0131  & ~\i_rx_phy_rxd_s_reg/P0001  ;
  assign n279 = ~\i_rx_phy_rxd_r_reg/NET0131  & \i_rx_phy_rxd_s_reg/P0001  ;
  assign n280 = ~n278 & ~n279 ;
  assign n281 = \i_rx_phy_rx_en_reg/NET0131  & ~n280 ;
  assign n284 = ~\i_rx_phy_dpll_state_reg[0]/P0001  & ~n281 ;
  assign n282 = \i_rx_phy_dpll_state_reg[0]/P0001  & ~\i_rx_phy_dpll_state_reg[1]/NET0131  ;
  assign n283 = n281 & n282 ;
  assign n285 = rst_pad & ~n283 ;
  assign n286 = ~n284 & n285 ;
  assign n287 = \i_rx_phy_dpll_state_reg[1]/NET0131  & n284 ;
  assign n288 = ~n282 & ~n287 ;
  assign n289 = rst_pad & ~n288 ;
  assign n290 = \i_tx_phy_append_eop_reg/P0001  & ~\i_tx_phy_append_eop_sync2_reg/P0001  ;
  assign n291 = ~n136 & ~n290 ;
  assign n292 = rst_pad & ~n291 ;
  assign n293 = ~\rst_cnt_reg[1]/NET0131  & ~n118 ;
  assign n294 = ~n119 & n123 ;
  assign n295 = ~n293 & n294 ;
  assign n296 = ~\i_rx_phy_bit_cnt_reg[0]/NET0131  & ~n170 ;
  assign n297 = n167 & ~n171 ;
  assign n298 = ~n296 & n297 ;
  assign n300 = \i_tx_phy_append_eop_sync3_reg/NET0131  & phy_tx_mode_pad ;
  assign n301 = \i_rx_phy_fs_ce_reg/P0001  & ~n300 ;
  assign n302 = \i_tx_phy_sd_nrzi_o_reg/NET0131  & n301 ;
  assign n299 = ~\i_rx_phy_fs_ce_reg/P0001  & txdp_pad ;
  assign n303 = rst_pad & ~n299 ;
  assign n304 = ~n302 & n303 ;
  assign n305 = ~\i_tx_phy_bit_cnt_reg[0]/NET0131  & ~n246 ;
  assign n306 = n250 & ~n259 ;
  assign n307 = ~n305 & n306 ;
  assign n308 = ~\i_tx_phy_bit_cnt_reg[1]/NET0131  & ~n259 ;
  assign n309 = n250 & ~n260 ;
  assign n310 = ~n308 & n309 ;
  assign n312 = ~\i_rx_phy_one_cnt_reg[0]/NET0131  & ~n267 ;
  assign n311 = \i_rx_phy_fs_ce_reg/P0001  & \i_rx_phy_one_cnt_reg[0]/NET0131  ;
  assign n313 = n167 & ~n311 ;
  assign n314 = ~n312 & n313 ;
  assign n315 = ~\i_rx_phy_bit_cnt_reg[1]/NET0131  & ~n171 ;
  assign n316 = n167 & ~n172 ;
  assign n317 = ~n315 & n316 ;
  assign n319 = ~\i_tx_phy_one_cnt_reg[0]/NET0131  & ~n247 ;
  assign n318 = \i_rx_phy_fs_ce_reg/P0001  & \i_tx_phy_one_cnt_reg[0]/NET0131  ;
  assign n320 = n250 & ~n318 ;
  assign n321 = ~n319 & n320 ;
  assign n322 = ~\i_rx_phy_rxd_s_reg/P0001  & ~\i_rx_phy_sd_r_reg/NET0131  ;
  assign n323 = \i_rx_phy_rxd_s_reg/P0001  & \i_rx_phy_sd_r_reg/NET0131  ;
  assign n324 = ~n322 & ~n323 ;
  assign n325 = \i_rx_phy_fs_ce_reg/P0001  & ~n324 ;
  assign n326 = ~\i_rx_phy_fs_ce_reg/P0001  & \i_rx_phy_sd_nrzi_reg/NET0131  ;
  assign n327 = RxActive_o_pad & ~n326 ;
  assign n328 = ~n325 & n327 ;
  assign n329 = rst_pad & ~n328 ;
  assign n332 = ~n133 & ~n233 ;
  assign n330 = \i_tx_phy_data_done_reg/NET0131  & n132 ;
  assign n331 = n133 & ~n330 ;
  assign n333 = TxValid_i_pad & rst_pad ;
  assign n334 = ~n331 & n333 ;
  assign n335 = ~n332 & n334 ;
  assign n336 = ~\i_rx_phy_fs_ce_reg/P0001  & txdn_pad ;
  assign n337 = ~\i_tx_phy_sd_nrzi_o_reg/NET0131  & phy_tx_mode_pad ;
  assign n338 = ~\i_tx_phy_append_eop_sync3_reg/NET0131  & ~n337 ;
  assign n339 = n301 & ~n338 ;
  assign n340 = ~n336 & ~n339 ;
  assign n341 = rst_pad & ~n340 ;
  assign n342 = ~\i_rx_phy_fs_ce_reg/P0001  & \i_rx_phy_rx_valid_r_reg/P0001  ;
  assign n343 = ~RxValid_o_pad & ~n342 ;
  assign n344 = \i_rx_phy_fs_ce_reg/P0001  & ~\i_tx_phy_sd_bs_o_reg/NET0131  ;
  assign n346 = ~\i_tx_phy_sd_nrzi_o_reg/NET0131  & n344 ;
  assign n345 = \i_tx_phy_sd_nrzi_o_reg/NET0131  & ~n344 ;
  assign n347 = \i_tx_phy_txoe_r1_reg/P0001  & n250 ;
  assign n348 = ~n345 & n347 ;
  assign n349 = ~n346 & n348 ;
  assign n350 = \rst_cnt_reg[0]/NET0131  & \rst_cnt_reg[1]/NET0131  ;
  assign n351 = \rst_cnt_reg[4]/NET0131  & n350 ;
  assign n352 = n124 & n351 ;
  assign n353 = ~\rst_cnt_reg[0]/NET0131  & ~n117 ;
  assign n354 = ~n118 & n123 ;
  assign n355 = ~n353 & n354 ;
  assign n356 = \LineState_o[1]_pad  & \i_rx_phy_rxdn_s0_reg/P0001  ;
  assign n357 = ~\i_rx_phy_rxdn_s_r_reg/P0001  & ~n356 ;
  assign n358 = \LineState_o[0]_pad  & \i_rx_phy_rxdp_s0_reg/P0001  ;
  assign n359 = ~\i_rx_phy_rxdp_s_r_reg/P0001  & ~n358 ;
  assign n360 = \i_rx_phy_fs_ce_reg/P0001  & \i_tx_phy_append_eop_sync4_reg/P0001  ;
  assign n361 = \i_tx_phy_append_eop_sync3_reg/NET0131  & ~n360 ;
  assign n362 = \i_rx_phy_fs_ce_reg/P0001  & \i_tx_phy_append_eop_sync2_reg/P0001  ;
  assign n363 = ~n361 & ~n362 ;
  assign n364 = rst_pad & ~n363 ;
  assign n365 = ~\i_rx_phy_fs_ce_reg/P0001  & \i_tx_phy_sd_bs_o_reg/NET0131  ;
  assign n366 = \i_tx_phy_tx_ip_sync_reg/P0001  & n247 ;
  assign n367 = ~n365 & ~n366 ;
  assign n368 = rst_pad & ~n367 ;
  assign n369 = ~n233 & ~n330 ;
  assign n370 = ~n234 & ~n369 ;
  assign n371 = \i_rx_phy_shift_en_reg/NET0131  & n170 ;
  assign n372 = \i_rx_phy_rx_valid1_reg/P0001  & n170 ;
  assign n373 = \i_rx_phy_fs_ce_reg/P0001  & ~\i_tx_phy_txoe_r1_reg/P0001  ;
  assign n374 = ~\i_tx_phy_txoe_r2_reg/P0001  & n373 ;
  assign n375 = ~\i_rx_phy_fs_ce_reg/P0001  & txoe_pad ;
  assign n376 = rst_pad & ~n375 ;
  assign n377 = ~n374 & n376 ;
  assign n378 = \i_rx_phy_rxd_s0_reg/P0001  & \i_rx_phy_rxd_s_reg/P0001  ;
  assign n379 = ~\i_rx_phy_rxd_s0_reg/P0001  & ~\i_rx_phy_rxd_s_reg/P0001  ;
  assign n380 = \i_rx_phy_rxd_s1_reg/P0001  & ~n379 ;
  assign n381 = ~n378 & ~n380 ;
  assign n382 = \i_tx_phy_bit_cnt_reg[0]/NET0131  & \i_tx_phy_bit_cnt_reg[1]/NET0131  ;
  assign n383 = \i_tx_phy_bit_cnt_reg[2]/P0001  & n382 ;
  assign n384 = ~n245 & n383 ;
  assign n386 = \i_rx_phy_fs_ce_reg/P0001  & ~\i_tx_phy_tx_ip_sync_reg/P0001  ;
  assign n385 = ~\i_rx_phy_fs_ce_reg/P0001  & ~\i_tx_phy_txoe_r1_reg/P0001  ;
  assign n387 = rst_pad & ~n385 ;
  assign n388 = ~n386 & n387 ;
  assign n390 = \i_rx_phy_fs_ce_reg/P0001  & ~\i_tx_phy_tx_ip_reg/P0001  ;
  assign n389 = ~\i_rx_phy_fs_ce_reg/P0001  & ~\i_tx_phy_tx_ip_sync_reg/P0001  ;
  assign n391 = rst_pad & ~n389 ;
  assign n392 = ~n390 & n391 ;
  assign n393 = ~\i_rx_phy_fs_ce_reg/P0001  & ~\i_tx_phy_txoe_r2_reg/P0001  ;
  assign n394 = rst_pad & ~n373 ;
  assign n395 = ~n393 & n394 ;
  assign n397 = \i_rx_phy_fs_ce_reg/P0001  & ~\i_tx_phy_append_eop_reg/P0001  ;
  assign n396 = ~\i_rx_phy_fs_ce_reg/P0001  & ~\i_tx_phy_append_eop_sync1_reg/P0001  ;
  assign n398 = rst_pad & ~n396 ;
  assign n399 = ~n397 & n398 ;
  assign n401 = \i_rx_phy_fs_ce_reg/P0001  & ~\i_tx_phy_append_eop_sync1_reg/P0001  ;
  assign n400 = ~\i_rx_phy_fs_ce_reg/P0001  & ~\i_tx_phy_append_eop_sync2_reg/P0001  ;
  assign n402 = rst_pad & ~n400 ;
  assign n403 = ~n401 & n402 ;
  assign n404 = ~\i_rx_phy_fs_ce_reg/P0001  & ~\i_tx_phy_append_eop_sync4_reg/P0001  ;
  assign n405 = rst_pad & ~n130 ;
  assign n406 = ~n404 & n405 ;
  assign n407 = ~\i_tx_phy_data_done_reg/NET0131  & \i_tx_phy_tx_ip_reg/P0001  ;
  assign n408 = n333 & ~n407 ;
  assign n409 = ~\i_rx_phy_fs_state_reg[0]/NET0131  & ~n107 ;
  assign n410 = rst_pad & ~n108 ;
  assign n411 = ~n409 & n410 ;
  assign n412 = \i_rx_phy_rx_valid_r_reg/P0001  & n104 ;
  assign n413 = RxActive_o_pad & ~n412 ;
  assign n415 = ~\i_rx_phy_fs_state_reg[1]/P0001  & ~\i_rx_phy_rx_en_reg/NET0131  ;
  assign n414 = \i_rx_phy_fs_state_reg[0]/NET0131  & \i_rx_phy_fs_state_reg[2]/NET0131  ;
  assign n416 = n101 & n414 ;
  assign n417 = ~n415 & n416 ;
  assign n418 = n107 & n417 ;
  assign n419 = \i_rx_phy_rx_en_reg/NET0131  & n418 ;
  assign n420 = ~n413 & ~n419 ;
  assign n421 = rst_pad & ~n420 ;
  assign n428 = \i_rx_phy_fs_state_reg[2]/NET0131  & n103 ;
  assign n424 = \i_rx_phy_fs_state_reg[0]/NET0131  & ~\i_rx_phy_fs_state_reg[2]/NET0131  ;
  assign n425 = \i_rx_phy_fs_state_reg[1]/P0001  & ~n424 ;
  assign n423 = ~\i_rx_phy_fs_state_reg[1]/P0001  & ~n414 ;
  assign n426 = n111 & ~n423 ;
  assign n427 = ~n425 & n426 ;
  assign n429 = n107 & ~n427 ;
  assign n430 = ~n428 & n429 ;
  assign n422 = ~\i_rx_phy_fs_state_reg[2]/NET0131  & ~n107 ;
  assign n431 = rst_pad & ~n422 ;
  assign n432 = ~n430 & n431 ;
  assign n433 = ~n111 & n424 ;
  assign n435 = ~\i_rx_phy_fs_state_reg[1]/P0001  & ~n111 ;
  assign n436 = \i_rx_phy_fs_state_reg[0]/NET0131  & ~n435 ;
  assign n434 = ~\i_rx_phy_fs_state_reg[1]/P0001  & ~\i_rx_phy_fs_state_reg[2]/NET0131  ;
  assign n437 = ~n102 & ~n434 ;
  assign n438 = ~n436 & n437 ;
  assign n439 = ~n433 & ~n438 ;
  assign n440 = n107 & ~n439 ;
  assign n443 = n267 & n268 ;
  assign n444 = ~\i_rx_phy_one_cnt_reg[2]/NET0131  & ~n443 ;
  assign n441 = \i_rx_phy_fs_ce_reg/P0001  & \i_rx_phy_one_cnt_reg[2]/NET0131  ;
  assign n442 = ~n269 & n441 ;
  assign n445 = n167 & ~n442 ;
  assign n446 = ~n444 & n445 ;
  assign n447 = ~\i_tx_phy_append_eop_sync3_reg/NET0131  & \i_tx_phy_tx_ip_reg/P0001  ;
  assign n448 = ~n138 & ~n447 ;
  assign n449 = rst_pad & ~n448 ;
  assign n450 = ~\i_rx_phy_fs_ce_reg/P0001  & \i_rx_phy_shift_en_reg/NET0131  ;
  assign n451 = ~n227 & ~n450 ;
  assign n452 = ~n418 & n451 ;
  assign n453 = \i_rx_phy_fs_ce_reg/P0001  & \i_rx_phy_rxd_s_reg/P0001  ;
  assign n454 = ~\i_rx_phy_fs_ce_reg/P0001  & \i_rx_phy_sd_r_reg/NET0131  ;
  assign n455 = ~n453 & ~n454 ;
  assign RxError_o_pad = ~n100 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1661/_0_  = n116 ;
  assign \g1680/_0_  = n127 ;
  assign \g1695/_0_  = n151 ;
  assign \g1703/_1_  = n155 ;
  assign \g1707/_0_  = n159 ;
  assign \g1725/_0_  = n162 ;
  assign \g1728/_0_  = ~n166 ;
  assign \g1729/_0_  = n176 ;
  assign \g1736/_0_  = n198 ;
  assign \g1737/_0_  = n202 ;
  assign \g1738/_0_  = n206 ;
  assign \g1739/_0_  = n210 ;
  assign \g1740/_0_  = n214 ;
  assign \g1741/_0_  = n218 ;
  assign \g1742/_0_  = n222 ;
  assign \g1743/_0_  = n226 ;
  assign \g1747/_3_  = n230 ;
  assign \g1748/_0_  = n232 ;
  assign \g1757/_0_  = n236 ;
  assign \g1758/_0_  = n242 ;
  assign \g1763/_0_  = n255 ;
  assign \g1764/_0_  = n258 ;
  assign \g1811/_0_  = n264 ;
  assign \g1812/_0_  = n272 ;
  assign \g1815/_0_  = n277 ;
  assign \g1816/_0_  = ~n286 ;
  assign \g1820/_1_  = n104 ;
  assign \g1821/_0_  = n289 ;
  assign \g1837/_0_  = n292 ;
  assign \g1838/_0_  = n295 ;
  assign \g1841/_0_  = n298 ;
  assign \g1842/_0_  = ~n304 ;
  assign \g1843/_0_  = n307 ;
  assign \g1844/_0_  = n310 ;
  assign \g1845/_0_  = n314 ;
  assign \g1846/_0_  = n317 ;
  assign \g1848/_0_  = n321 ;
  assign \g1851/_0_  = n329 ;
  assign \g1852/_0_  = n335 ;
  assign \g1853/_0_  = n341 ;
  assign \g1857/_0_  = ~n343 ;
  assign \g1858/_0_  = ~n349 ;
  assign \g1865/_0_  = n352 ;
  assign \g1869/_0_  = n355 ;
  assign \g1871/_0_  = ~n357 ;
  assign \g1872/_0_  = ~n359 ;
  assign \g1873/_0_  = n364 ;
  assign \g1876/_0_  = n368 ;
  assign \g1878/_0_  = n370 ;
  assign \g1897/_1_  = n371 ;
  assign \g1901/_0_  = n372 ;
  assign \g1904/_0_  = ~n377 ;
  assign \g1928/_0_  = ~n381 ;
  assign \g1936/_3_  = n384 ;
  assign \g1961/_0_  = n388 ;
  assign \g1962/_0_  = n392 ;
  assign \g1963/_0_  = n395 ;
  assign \g1966/_0_  = n399 ;
  assign \g1967/_0_  = n403 ;
  assign \g1968/_0_  = n406 ;
  assign \g1975/_0_  = n358 ;
  assign \g1980/_0_  = n356 ;
  assign \g2055/_0_  = n408 ;
  assign \g2112/_0_  = n282 ;
  assign \g2411/_2_  = n411 ;
  assign \g2463/_0_  = n421 ;
  assign \g2501/_0_  = n432 ;
  assign \g2620/_0_  = n440 ;
  assign \g2650/_0_  = n446 ;
  assign \g2657/_0_  = n449 ;
  assign \g2671/_0_  = ~n452 ;
  assign \i_rx_phy_sd_r_reg/NET0131_reg_syn_3  = ~n455 ;
endmodule
