module top (\P1_B_reg/NET0131 , \P1_IR_reg[0]/NET0131 , \P1_IR_reg[10]/NET0131 , \P1_IR_reg[11]/NET0131 , \P1_IR_reg[12]/NET0131 , \P1_IR_reg[13]/NET0131 , \P1_IR_reg[14]/NET0131 , \P1_IR_reg[15]/NET0131 , \P1_IR_reg[16]/NET0131 , \P1_IR_reg[17]/NET0131 , \P1_IR_reg[18]/NET0131 , \P1_IR_reg[19]/NET0131 , \P1_IR_reg[1]/NET0131 , \P1_IR_reg[20]/NET0131 , \P1_IR_reg[21]/NET0131 , \P1_IR_reg[22]/NET0131 , \P1_IR_reg[23]/NET0131 , \P1_IR_reg[24]/NET0131 , \P1_IR_reg[25]/NET0131 , \P1_IR_reg[26]/NET0131 , \P1_IR_reg[27]/NET0131 , \P1_IR_reg[28]/NET0131 , \P1_IR_reg[29]/NET0131 , \P1_IR_reg[2]/NET0131 , \P1_IR_reg[30]/NET0131 , \P1_IR_reg[31]/NET0131 , \P1_IR_reg[3]/NET0131 , \P1_IR_reg[4]/NET0131 , \P1_IR_reg[5]/NET0131 , \P1_IR_reg[6]/NET0131 , \P1_IR_reg[7]/NET0131 , \P1_IR_reg[8]/NET0131 , \P1_IR_reg[9]/NET0131 , \P1_addr_reg[0]/NET0131 , \P1_addr_reg[10]/NET0131 , \P1_addr_reg[11]/NET0131 , \P1_addr_reg[12]/NET0131 , \P1_addr_reg[13]/NET0131 , \P1_addr_reg[14]/NET0131 , \P1_addr_reg[15]/NET0131 , \P1_addr_reg[16]/NET0131 , \P1_addr_reg[17]/NET0131 , \P1_addr_reg[18]/NET0131 , \P1_addr_reg[19]/NET0131 , \P1_addr_reg[1]/NET0131 , \P1_addr_reg[2]/NET0131 , \P1_addr_reg[3]/NET0131 , \P1_addr_reg[4]/NET0131 , \P1_addr_reg[5]/NET0131 , \P1_addr_reg[6]/NET0131 , \P1_addr_reg[7]/NET0131 , \P1_addr_reg[8]/NET0131 , \P1_addr_reg[9]/NET0131 , \P1_d_reg[0]/NET0131 , \P1_d_reg[1]/NET0131 , \P1_datao_reg[0]/NET0131 , \P1_datao_reg[10]/NET0131 , \P1_datao_reg[11]/NET0131 , \P1_datao_reg[12]/NET0131 , \P1_datao_reg[13]/NET0131 , \P1_datao_reg[14]/NET0131 , \P1_datao_reg[15]/NET0131 , \P1_datao_reg[16]/NET0131 , \P1_datao_reg[17]/NET0131 , \P1_datao_reg[18]/NET0131 , \P1_datao_reg[19]/NET0131 , \P1_datao_reg[1]/NET0131 , \P1_datao_reg[20]/NET0131 , \P1_datao_reg[21]/NET0131 , \P1_datao_reg[22]/NET0131 , \P1_datao_reg[23]/NET0131 , \P1_datao_reg[24]/NET0131 , \P1_datao_reg[25]/NET0131 , \P1_datao_reg[26]/NET0131 , \P1_datao_reg[27]/NET0131 , \P1_datao_reg[28]/NET0131 , \P1_datao_reg[29]/NET0131 , \P1_datao_reg[2]/NET0131 , \P1_datao_reg[30]/NET0131 , \P1_datao_reg[31]/NET0131 , \P1_datao_reg[3]/NET0131 , \P1_datao_reg[4]/NET0131 , \P1_datao_reg[5]/NET0131 , \P1_datao_reg[6]/NET0131 , \P1_datao_reg[7]/NET0131 , \P1_datao_reg[8]/NET0131 , \P1_datao_reg[9]/NET0131 , \P1_rd_reg/NET0131 , \P1_reg0_reg[0]/NET0131 , \P1_reg0_reg[10]/NET0131 , \P1_reg0_reg[11]/NET0131 , \P1_reg0_reg[12]/NET0131 , \P1_reg0_reg[13]/NET0131 , \P1_reg0_reg[14]/NET0131 , \P1_reg0_reg[15]/NET0131 , \P1_reg0_reg[16]/NET0131 , \P1_reg0_reg[17]/NET0131 , \P1_reg0_reg[18]/NET0131 , \P1_reg0_reg[19]/NET0131 , \P1_reg0_reg[1]/NET0131 , \P1_reg0_reg[20]/NET0131 , \P1_reg0_reg[21]/NET0131 , \P1_reg0_reg[22]/NET0131 , \P1_reg0_reg[23]/NET0131 , \P1_reg0_reg[24]/NET0131 , \P1_reg0_reg[25]/NET0131 , \P1_reg0_reg[26]/NET0131 , \P1_reg0_reg[27]/NET0131 , \P1_reg0_reg[28]/NET0131 , \P1_reg0_reg[29]/NET0131 , \P1_reg0_reg[2]/NET0131 , \P1_reg0_reg[30]/NET0131 , \P1_reg0_reg[31]/NET0131 , \P1_reg0_reg[3]/NET0131 , \P1_reg0_reg[4]/NET0131 , \P1_reg0_reg[5]/NET0131 , \P1_reg0_reg[6]/NET0131 , \P1_reg0_reg[7]/NET0131 , \P1_reg0_reg[8]/NET0131 , \P1_reg0_reg[9]/NET0131 , \P1_reg1_reg[0]/NET0131 , \P1_reg1_reg[10]/NET0131 , \P1_reg1_reg[11]/NET0131 , \P1_reg1_reg[12]/NET0131 , \P1_reg1_reg[13]/NET0131 , \P1_reg1_reg[14]/NET0131 , \P1_reg1_reg[15]/NET0131 , \P1_reg1_reg[16]/NET0131 , \P1_reg1_reg[17]/NET0131 , \P1_reg1_reg[18]/NET0131 , \P1_reg1_reg[19]/NET0131 , \P1_reg1_reg[1]/NET0131 , \P1_reg1_reg[20]/NET0131 , \P1_reg1_reg[21]/NET0131 , \P1_reg1_reg[22]/NET0131 , \P1_reg1_reg[23]/NET0131 , \P1_reg1_reg[24]/NET0131 , \P1_reg1_reg[25]/NET0131 , \P1_reg1_reg[26]/NET0131 , \P1_reg1_reg[27]/NET0131 , \P1_reg1_reg[28]/NET0131 , \P1_reg1_reg[29]/NET0131 , \P1_reg1_reg[2]/NET0131 , \P1_reg1_reg[30]/NET0131 , \P1_reg1_reg[31]/NET0131 , \P1_reg1_reg[3]/NET0131 , \P1_reg1_reg[4]/NET0131 , \P1_reg1_reg[5]/NET0131 , \P1_reg1_reg[6]/NET0131 , \P1_reg1_reg[7]/NET0131 , \P1_reg1_reg[8]/NET0131 , \P1_reg1_reg[9]/NET0131 , \P1_reg2_reg[0]/NET0131 , \P1_reg2_reg[10]/NET0131 , \P1_reg2_reg[11]/NET0131 , \P1_reg2_reg[12]/NET0131 , \P1_reg2_reg[13]/NET0131 , \P1_reg2_reg[14]/NET0131 , \P1_reg2_reg[15]/NET0131 , \P1_reg2_reg[16]/NET0131 , \P1_reg2_reg[17]/NET0131 , \P1_reg2_reg[18]/NET0131 , \P1_reg2_reg[19]/NET0131 , \P1_reg2_reg[1]/NET0131 , \P1_reg2_reg[20]/NET0131 , \P1_reg2_reg[21]/NET0131 , \P1_reg2_reg[22]/NET0131 , \P1_reg2_reg[23]/NET0131 , \P1_reg2_reg[24]/NET0131 , \P1_reg2_reg[25]/NET0131 , \P1_reg2_reg[26]/NET0131 , \P1_reg2_reg[27]/NET0131 , \P1_reg2_reg[28]/NET0131 , \P1_reg2_reg[29]/NET0131 , \P1_reg2_reg[2]/NET0131 , \P1_reg2_reg[30]/NET0131 , \P1_reg2_reg[31]/NET0131 , \P1_reg2_reg[3]/NET0131 , \P1_reg2_reg[4]/NET0131 , \P1_reg2_reg[5]/NET0131 , \P1_reg2_reg[6]/NET0131 , \P1_reg2_reg[7]/NET0131 , \P1_reg2_reg[8]/NET0131 , \P1_reg2_reg[9]/NET0131 , \P1_reg3_reg[0]/NET0131 , \P1_reg3_reg[10]/NET0131 , \P1_reg3_reg[11]/NET0131 , \P1_reg3_reg[12]/NET0131 , \P1_reg3_reg[13]/NET0131 , \P1_reg3_reg[14]/NET0131 , \P1_reg3_reg[15]/NET0131 , \P1_reg3_reg[16]/NET0131 , \P1_reg3_reg[17]/NET0131 , \P1_reg3_reg[18]/NET0131 , \P1_reg3_reg[19]/NET0131 , \P1_reg3_reg[1]/NET0131 , \P1_reg3_reg[20]/NET0131 , \P1_reg3_reg[21]/NET0131 , \P1_reg3_reg[22]/NET0131 , \P1_reg3_reg[23]/NET0131 , \P1_reg3_reg[24]/NET0131 , \P1_reg3_reg[25]/NET0131 , \P1_reg3_reg[26]/NET0131 , \P1_reg3_reg[27]/NET0131 , \P1_reg3_reg[28]/NET0131 , \P1_reg3_reg[2]/NET0131 , \P1_reg3_reg[3]/NET0131 , \P1_reg3_reg[4]/NET0131 , \P1_reg3_reg[5]/NET0131 , \P1_reg3_reg[6]/NET0131 , \P1_reg3_reg[7]/NET0131 , \P1_reg3_reg[8]/NET0131 , \P1_reg3_reg[9]/NET0131 , \P1_state_reg[0]/NET0131 , \P1_wr_reg/NET0131 , \P2_B_reg/NET0131 , \P2_IR_reg[0]/NET0131 , \P2_IR_reg[10]/NET0131 , \P2_IR_reg[11]/NET0131 , \P2_IR_reg[12]/NET0131 , \P2_IR_reg[13]/NET0131 , \P2_IR_reg[14]/NET0131 , \P2_IR_reg[15]/NET0131 , \P2_IR_reg[16]/NET0131 , \P2_IR_reg[17]/NET0131 , \P2_IR_reg[18]/NET0131 , \P2_IR_reg[19]/NET0131 , \P2_IR_reg[1]/NET0131 , \P2_IR_reg[20]/NET0131 , \P2_IR_reg[21]/NET0131 , \P2_IR_reg[22]/NET0131 , \P2_IR_reg[23]/NET0131 , \P2_IR_reg[24]/NET0131 , \P2_IR_reg[25]/NET0131 , \P2_IR_reg[26]/NET0131 , \P2_IR_reg[27]/NET0131 , \P2_IR_reg[28]/NET0131 , \P2_IR_reg[29]/NET0131 , \P2_IR_reg[2]/NET0131 , \P2_IR_reg[30]/NET0131 , \P2_IR_reg[31]/NET0131 , \P2_IR_reg[3]/NET0131 , \P2_IR_reg[4]/NET0131 , \P2_IR_reg[5]/NET0131 , \P2_IR_reg[6]/NET0131 , \P2_IR_reg[7]/NET0131 , \P2_IR_reg[8]/NET0131 , \P2_IR_reg[9]/NET0131 , \P2_addr_reg[0]/NET0131 , \P2_addr_reg[10]/NET0131 , \P2_addr_reg[11]/NET0131 , \P2_addr_reg[12]/NET0131 , \P2_addr_reg[13]/NET0131 , \P2_addr_reg[14]/NET0131 , \P2_addr_reg[15]/NET0131 , \P2_addr_reg[16]/NET0131 , \P2_addr_reg[17]/NET0131 , \P2_addr_reg[18]/NET0131 , \P2_addr_reg[19]/NET0131 , \P2_addr_reg[1]/NET0131 , \P2_addr_reg[2]/NET0131 , \P2_addr_reg[3]/NET0131 , \P2_addr_reg[4]/NET0131 , \P2_addr_reg[5]/NET0131 , \P2_addr_reg[6]/NET0131 , \P2_addr_reg[7]/NET0131 , \P2_addr_reg[8]/NET0131 , \P2_addr_reg[9]/NET0131 , \P2_d_reg[0]/NET0131 , \P2_d_reg[1]/NET0131 , \P2_datao_reg[0]/NET0131 , \P2_datao_reg[10]/NET0131 , \P2_datao_reg[11]/NET0131 , \P2_datao_reg[12]/NET0131 , \P2_datao_reg[13]/NET0131 , \P2_datao_reg[14]/NET0131 , \P2_datao_reg[15]/NET0131 , \P2_datao_reg[16]/NET0131 , \P2_datao_reg[17]/NET0131 , \P2_datao_reg[18]/NET0131 , \P2_datao_reg[19]/NET0131 , \P2_datao_reg[1]/NET0131 , \P2_datao_reg[20]/NET0131 , \P2_datao_reg[21]/NET0131 , \P2_datao_reg[22]/NET0131 , \P2_datao_reg[23]/NET0131 , \P2_datao_reg[24]/NET0131 , \P2_datao_reg[25]/NET0131 , \P2_datao_reg[26]/NET0131 , \P2_datao_reg[27]/NET0131 , \P2_datao_reg[28]/NET0131 , \P2_datao_reg[29]/NET0131 , \P2_datao_reg[2]/NET0131 , \P2_datao_reg[30]/NET0131 , \P2_datao_reg[31]/NET0131 , \P2_datao_reg[3]/NET0131 , \P2_datao_reg[4]/NET0131 , \P2_datao_reg[5]/NET0131 , \P2_datao_reg[6]/NET0131 , \P2_datao_reg[7]/NET0131 , \P2_datao_reg[8]/NET0131 , \P2_datao_reg[9]/NET0131 , \P2_rd_reg/NET0131 , \P2_reg0_reg[0]/NET0131 , \P2_reg0_reg[10]/NET0131 , \P2_reg0_reg[11]/NET0131 , \P2_reg0_reg[12]/NET0131 , \P2_reg0_reg[13]/NET0131 , \P2_reg0_reg[14]/NET0131 , \P2_reg0_reg[15]/NET0131 , \P2_reg0_reg[16]/NET0131 , \P2_reg0_reg[17]/NET0131 , \P2_reg0_reg[18]/NET0131 , \P2_reg0_reg[19]/NET0131 , \P2_reg0_reg[1]/NET0131 , \P2_reg0_reg[20]/NET0131 , \P2_reg0_reg[21]/NET0131 , \P2_reg0_reg[22]/NET0131 , \P2_reg0_reg[23]/NET0131 , \P2_reg0_reg[24]/NET0131 , \P2_reg0_reg[25]/NET0131 , \P2_reg0_reg[26]/NET0131 , \P2_reg0_reg[27]/NET0131 , \P2_reg0_reg[28]/NET0131 , \P2_reg0_reg[29]/NET0131 , \P2_reg0_reg[2]/NET0131 , \P2_reg0_reg[30]/NET0131 , \P2_reg0_reg[31]/NET0131 , \P2_reg0_reg[3]/NET0131 , \P2_reg0_reg[4]/NET0131 , \P2_reg0_reg[5]/NET0131 , \P2_reg0_reg[6]/NET0131 , \P2_reg0_reg[7]/NET0131 , \P2_reg0_reg[8]/NET0131 , \P2_reg0_reg[9]/NET0131 , \P2_reg1_reg[0]/NET0131 , \P2_reg1_reg[10]/NET0131 , \P2_reg1_reg[11]/NET0131 , \P2_reg1_reg[12]/NET0131 , \P2_reg1_reg[13]/NET0131 , \P2_reg1_reg[14]/NET0131 , \P2_reg1_reg[15]/NET0131 , \P2_reg1_reg[16]/NET0131 , \P2_reg1_reg[17]/NET0131 , \P2_reg1_reg[18]/NET0131 , \P2_reg1_reg[19]/NET0131 , \P2_reg1_reg[1]/NET0131 , \P2_reg1_reg[20]/NET0131 , \P2_reg1_reg[21]/NET0131 , \P2_reg1_reg[22]/NET0131 , \P2_reg1_reg[23]/NET0131 , \P2_reg1_reg[24]/NET0131 , \P2_reg1_reg[25]/NET0131 , \P2_reg1_reg[26]/NET0131 , \P2_reg1_reg[27]/NET0131 , \P2_reg1_reg[28]/NET0131 , \P2_reg1_reg[29]/NET0131 , \P2_reg1_reg[2]/NET0131 , \P2_reg1_reg[30]/NET0131 , \P2_reg1_reg[31]/NET0131 , \P2_reg1_reg[3]/NET0131 , \P2_reg1_reg[4]/NET0131 , \P2_reg1_reg[5]/NET0131 , \P2_reg1_reg[6]/NET0131 , \P2_reg1_reg[7]/NET0131 , \P2_reg1_reg[8]/NET0131 , \P2_reg1_reg[9]/NET0131 , \P2_reg2_reg[0]/NET0131 , \P2_reg2_reg[10]/NET0131 , \P2_reg2_reg[11]/NET0131 , \P2_reg2_reg[12]/NET0131 , \P2_reg2_reg[13]/NET0131 , \P2_reg2_reg[14]/NET0131 , \P2_reg2_reg[15]/NET0131 , \P2_reg2_reg[16]/NET0131 , \P2_reg2_reg[17]/NET0131 , \P2_reg2_reg[18]/NET0131 , \P2_reg2_reg[19]/NET0131 , \P2_reg2_reg[1]/NET0131 , \P2_reg2_reg[20]/NET0131 , \P2_reg2_reg[21]/NET0131 , \P2_reg2_reg[22]/NET0131 , \P2_reg2_reg[23]/NET0131 , \P2_reg2_reg[24]/NET0131 , \P2_reg2_reg[25]/NET0131 , \P2_reg2_reg[26]/NET0131 , \P2_reg2_reg[27]/NET0131 , \P2_reg2_reg[28]/NET0131 , \P2_reg2_reg[29]/NET0131 , \P2_reg2_reg[2]/NET0131 , \P2_reg2_reg[30]/NET0131 , \P2_reg2_reg[31]/NET0131 , \P2_reg2_reg[3]/NET0131 , \P2_reg2_reg[4]/NET0131 , \P2_reg2_reg[5]/NET0131 , \P2_reg2_reg[6]/NET0131 , \P2_reg2_reg[7]/NET0131 , \P2_reg2_reg[8]/NET0131 , \P2_reg2_reg[9]/NET0131 , \P2_reg3_reg[0]/NET0131 , \P2_reg3_reg[10]/NET0131 , \P2_reg3_reg[11]/NET0131 , \P2_reg3_reg[12]/NET0131 , \P2_reg3_reg[13]/NET0131 , \P2_reg3_reg[14]/NET0131 , \P2_reg3_reg[15]/NET0131 , \P2_reg3_reg[16]/NET0131 , \P2_reg3_reg[17]/NET0131 , \P2_reg3_reg[18]/NET0131 , \P2_reg3_reg[19]/NET0131 , \P2_reg3_reg[1]/NET0131 , \P2_reg3_reg[20]/NET0131 , \P2_reg3_reg[21]/NET0131 , \P2_reg3_reg[22]/NET0131 , \P2_reg3_reg[23]/NET0131 , \P2_reg3_reg[24]/NET0131 , \P2_reg3_reg[25]/NET0131 , \P2_reg3_reg[26]/NET0131 , \P2_reg3_reg[27]/NET0131 , \P2_reg3_reg[28]/NET0131 , \P2_reg3_reg[2]/NET0131 , \P2_reg3_reg[3]/NET0131 , \P2_reg3_reg[4]/NET0131 , \P2_reg3_reg[5]/NET0131 , \P2_reg3_reg[6]/NET0131 , \P2_reg3_reg[7]/NET0131 , \P2_reg3_reg[8]/NET0131 , \P2_reg3_reg[9]/NET0131 , \P2_wr_reg/NET0131 , \si[0]_pad , \si[10]_pad , \si[11]_pad , \si[12]_pad , \si[13]_pad , \si[14]_pad , \si[15]_pad , \si[16]_pad , \si[17]_pad , \si[18]_pad , \si[19]_pad , \si[1]_pad , \si[20]_pad , \si[21]_pad , \si[22]_pad , \si[23]_pad , \si[24]_pad , \si[25]_pad , \si[26]_pad , \si[27]_pad , \si[28]_pad , \si[29]_pad , \si[2]_pad , \si[30]_pad , \si[31]_pad , \si[3]_pad , \si[4]_pad , \si[5]_pad , \si[6]_pad , \si[7]_pad , \si[8]_pad , \si[9]_pad , \P1_state_reg[0]/NET0131_syn_2 , \_al_n0 , \_al_n1 , \g70791/_0_ , \g70792/_0_ , \g70793/_0_ , \g70794/_0_ , \g70795/_0_ , \g70796/_0_ , \g70813/_0_ , \g70814/_0_ , \g70848/_0_ , \g70849/_0_ , \g70850/_0_ , \g70851/_0_ , \g70852/_0_ , \g70856/_0_ , \g70857/_0_ , \g70858/_0_ , \g70859/_0_ , \g70860/_0_ , \g70861/_0_ , \g70862/_0_ , \g70896/_0_ , \g70902/_0_ , \g70903/_0_ , \g70904/_0_ , \g70906/_0_ , \g70907/_0_ , \g70908/_0_ , \g70909/_0_ , \g70910/_0_ , \g70911/_0_ , \g70912/_0_ , \g70913/_0_ , \g70914/_0_ , \g70915/_0_ , \g70916/_0_ , \g70917/_0_ , \g70918/_0_ , \g70919/_0_ , \g70920/_0_ , \g70921/_0_ , \g70922/_0_ , \g70923/_0_ , \g70924/_0_ , \g70925/_0_ , \g70926/_0_ , \g70927/_0_ , \g70987/_0_ , \g70988/_0_ , \g70989/_0_ , \g70990/_0_ , \g70991/_0_ , \g71006/_0_ , \g71007/_0_ , \g71009/_0_ , \g71010/_0_ , \g71011/_0_ , \g71012/_0_ , \g71013/_0_ , \g71014/_0_ , \g71015/_0_ , \g71016/_0_ , \g71017/_0_ , \g71018/_0_ , \g71019/_0_ , \g71020/_0_ , \g71021/_0_ , \g71022/_0_ , \g71023/_0_ , \g71090/_0_ , \g71091/_0_ , \g71092/_0_ , \g71093/_0_ , \g71094/_0_ , \g71125/_0_ , \g71130/_0_ , \g71131/_0_ , \g71132/_0_ , \g71133/_0_ , \g71134/_0_ , \g71135/_0_ , \g71136/_0_ , \g71137/_0_ , \g71138/_0_ , \g71139/_0_ , \g71140/_0_ , \g71141/_0_ , \g71142/_0_ , \g71143/_0_ , \g71144/_0_ , \g71145/_0_ , \g71150/_0_ , \g71151/_0_ , \g71152/_0_ , \g71153/_0_ , \g71154/_0_ , \g71155/_0_ , \g71156/_0_ , \g71157/_0_ , \g71158/_0_ , \g71230/_0_ , \g71231/_0_ , \g71232/_0_ , \g71233/_0_ , \g71234/_0_ , \g71235/_0_ , \g71236/_0_ , \g71238/_0_ , \g71239/_0_ , \g71270/_0_ , \g71275/_0_ , \g71276/_0_ , \g71277/_0_ , \g71278/_0_ , \g71279/_0_ , \g71280/_0_ , \g71281/_0_ , \g71282/_0_ , \g71283/_0_ , \g71284/_0_ , \g71285/_0_ , \g71286/_0_ , \g71287/_0_ , \g71288/_0_ , \g71289/_0_ , \g71290/_0_ , \g71291/_0_ , \g71292/_0_ , \g71293/_0_ , \g71294/_0_ , \g71295/_0_ , \g71296/_0_ , \g71297/_0_ , \g71298/_0_ , \g71299/_0_ , \g71300/_0_ , \g71301/_0_ , \g71302/_0_ , \g71303/_0_ , \g71304/_0_ , \g71305/_0_ , \g71306/_0_ , \g71307/_0_ , \g71382/_0_ , \g71384/_0_ , \g71385/_0_ , \g71387/_0_ , \g71388/_0_ , \g71389/_0_ , \g71439/_0_ , \g71440/_0_ , \g71441/_0_ , \g71442/_0_ , \g71443/_0_ , \g71444/_0_ , \g71445/_0_ , \g71446/_0_ , \g71447/_0_ , \g71448/_0_ , \g71449/_0_ , \g71450/_0_ , \g71451/_0_ , \g71452/_0_ , \g71453/_0_ , \g71454/_0_ , \g71455/_0_ , \g71456/_0_ , \g71457/_0_ , \g71458/_0_ , \g71459/_0_ , \g71460/_0_ , \g71461/_0_ , \g71536/_0_ , \g71537/_0_ , \g71538/_0_ , \g71540/_0_ , \g71541/_0_ , \g71542/_0_ , \g71602/_0_ , \g71604/_0_ , \g71610/_0_ , \g71611/_0_ , \g71618/_0_ , \g71619/_0_ , \g71620/_0_ , \g71621/_0_ , \g71622/_0_ , \g71623/_0_ , \g71624/_0_ , \g71625/_0_ , \g71626/_0_ , \g71627/_0_ , \g71629/_0_ , \g71630/_0_ , \g71631/_0_ , \g71632/_0_ , \g71633/_0_ , \g71634/_0_ , \g71635/_0_ , \g71636/_0_ , \g71710/_0_ , \g71711/_0_ , \g71782/_0_ , \g71785/_0_ , \g71786/_0_ , \g71787/_0_ , \g71788/_0_ , \g71789/_0_ , \g71790/_0_ , \g71791/_0_ , \g71792/_0_ , \g71793/_0_ , \g71794/_0_ , \g71795/_0_ , \g71796/_0_ , \g71797/_0_ , \g71798/_0_ , \g71799/_0_ , \g71883/_0_ , \g72000/_0_ , \g72001/_0_ , \g72002/_0_ , \g72003/_0_ , \g72004/_0_ , \g72005/_0_ , \g72236/_0_ , \g72237/_0_ , \g72238/_0_ , \g72239/_0_ , \g72240/_0_ , \g72372/_0_ , \g72376/_0_ , \g72383/_0_ , \g72561/_0_ , \g72562/_0_ , \g72563/_0_ , \g72564/_0_ , \g72970/_0_ , \g72980/_0_ , \g72981/_0_ , \g72982/_0_ , \g72983/_0_ , \g74234/_0_ , \g74260/_0_ , \g75086/_0_ , \g75087/_0_ , \g75088/_0_ , \g75089/_0_ , \g75091/_0_ , \g75092/_0_ , \g80304/_3_ , \g80305/_3_ , \g80306/_3_ , \g80307/_3_ , \g80308/_0_ , \g80309/_0_ , \g80815/_0_ , \g80816/_0_ , \g80817/_0_ , \g80818/_0_ , \g80819/_0_ , \g80820/_0_ , \g80821/_0_ , \g80822/_0_ , \g80823/_0_ , \g80824/_0_ , \g80825/_0_ , \g80826/_3_ , \g80827/_0_ , \g80828/_0_ , \g80829/_0_ , \g80830/_0_ , \g80831/_0_ , \g80832/_0_ , \g80833/_0_ , \g80834/_0_ , \g80835/_0_ , \g80836/_0_ , \g80837/_0_ , \g80838/_3_ , \g80839/_0_ , \g80840/_3_ , \g80841/_0_ , \g80859/_3_ , \g80860/_3_ , \g80861/_3_ , \g80862/_3_ , \g80863/_3_ , \g80864/_3_ , \g80865/_3_ , \g80866/_3_ , \g80867/_3_ , \g80868/_3_ , \g80869/_3_ , \g80870/_3_ , \g80871/_3_ , \g80872/_3_ , \g80873/_3_ , \g80874/_3_ , \g80875/_3_ , \g80876/_3_ , \g80877/_3_ , \g80878/_3_ , \g80879/_0_ , \g80880/_3_ , \g80881/_3_ , \g80882/_3_ , \g80883/_3_ , \g80884/_3_ , \g80885/_3_ , \g80886/_3_ , \g80888/_0_ , \g81262/_0_ , \g81278/_0_ , \g81884/_0_ , \g81893/_0_ , \g81896/_0_ , \g81897/_0_ , \g81898/_0_ , \g81899/_0_ , \g81900/_0_ , \g81901/_0_ , \g81902/_0_ , \g81903/_0_ , \g81904/_0_ , \g81905/_0_ , \g81906/_0_ , \g81907/_0_ , \g81908/_0_ , \g81909/_0_ , \g81910/_0_ , \g81911/_0_ , \g81923/_0_ , \g81924/_0_ , \g81925/_0_ , \g81926/_0_ , \g82414/_0_ , \g82532/_0_ , \g83134/_0_ , \g83135/_0_ , \g83141/_0_ , \g83142/_0_ , \g83145/_0_ , \g83146/_0_ , \g83147/_0_ , \g83148/_0_ , \g83152/_0_ , \g83153/_0_ , \g83154/_0_ , \g83155/_0_ , \g83156/_0_ , \g83157/_0_ , \g83158/_0_ , \g83159/_0_ , \g83164/_0_ , \g83165/_0_ , \g83177/_0_ , \g83178/_0_ , \g83409/_0_ , \g83411/_0_ , \g83807/u3_syn_4 , \g84138/u3_syn_4 , \g85062/_0_ , \g85079/_2_ , \g85113/_0_ , \g85121/_0_ , \g85594/_0_ , \g85663/_0_ , \g85669/_0_ , \g85749/_0_ , \g85784/_0_ , \g85809/_0_ , \g85817/_0_ , \g85828/_0_ , \g85845/_0_ , \g85851/_0_ , \g85858/_0_ , \g85871/_0_ , \g85882_dup/_0_ , \g85891/_0_ , \g85900/_0_ , \g85905/_0_ , \g85917/_0_ , \g85934/_0_ , \g85949/_0_ , \g85971/_0_ , \g85997/_0_ , \g86044/_0_ , \g86053/_0_ , \g86063/_0_ , \g86082/_0_ , \g86088/_0_ , \g86098/_0_ , \g86105/_0_ , \g86179/_0_ , \g86256_dup/_0_ , \g86264/_0_ , \g86273/_0_ , \g86281/_0_ , \g86288/_0_ , \g86297/_0_ , \g86304/_0_ , \g86310/_0_ , \g86320/_0_ , \g86328/_0_ , \g86339/_0_ , \g86353/_0_ , \g86360/_0_ , \g86368/_0_ , \g86373/_0_ , \g86385/_0_ , \g86392/_0_ , \g86399/_0_ , \g86421/_0_ , \g86432/_0_ , \g87592/_1__syn_2 , \g87632/_1_ , \g92847/_0_ , \g92957/_0_ , \g93056/_0_ , \g93289/_0_ , \g93538_dup95061/_0_ , \g93856/_0_ , \g93870/_0_ , \g94004/_0_ , \g94128/_0_ , \g94173/_0_ , \g94187/_0_ , \g94191/_0_ , \g94318/_0_ , \g94505/_0_ , rd_pad, \so[0]_pad , \so[10]_pad , \so[11]_pad , \so[12]_pad , \so[13]_pad , \so[14]_pad , \so[15]_pad , \so[16]_pad , \so[17]_pad , \so[18]_pad , \so[19]_pad , \so[1]_pad , \so[2]_pad , \so[3]_pad , \so[4]_pad , \so[5]_pad , \so[6]_pad , \so[7]_pad , \so[8]_pad , \so[9]_pad , wr_pad);
	input \P1_B_reg/NET0131  ;
	input \P1_IR_reg[0]/NET0131  ;
	input \P1_IR_reg[10]/NET0131  ;
	input \P1_IR_reg[11]/NET0131  ;
	input \P1_IR_reg[12]/NET0131  ;
	input \P1_IR_reg[13]/NET0131  ;
	input \P1_IR_reg[14]/NET0131  ;
	input \P1_IR_reg[15]/NET0131  ;
	input \P1_IR_reg[16]/NET0131  ;
	input \P1_IR_reg[17]/NET0131  ;
	input \P1_IR_reg[18]/NET0131  ;
	input \P1_IR_reg[19]/NET0131  ;
	input \P1_IR_reg[1]/NET0131  ;
	input \P1_IR_reg[20]/NET0131  ;
	input \P1_IR_reg[21]/NET0131  ;
	input \P1_IR_reg[22]/NET0131  ;
	input \P1_IR_reg[23]/NET0131  ;
	input \P1_IR_reg[24]/NET0131  ;
	input \P1_IR_reg[25]/NET0131  ;
	input \P1_IR_reg[26]/NET0131  ;
	input \P1_IR_reg[27]/NET0131  ;
	input \P1_IR_reg[28]/NET0131  ;
	input \P1_IR_reg[29]/NET0131  ;
	input \P1_IR_reg[2]/NET0131  ;
	input \P1_IR_reg[30]/NET0131  ;
	input \P1_IR_reg[31]/NET0131  ;
	input \P1_IR_reg[3]/NET0131  ;
	input \P1_IR_reg[4]/NET0131  ;
	input \P1_IR_reg[5]/NET0131  ;
	input \P1_IR_reg[6]/NET0131  ;
	input \P1_IR_reg[7]/NET0131  ;
	input \P1_IR_reg[8]/NET0131  ;
	input \P1_IR_reg[9]/NET0131  ;
	input \P1_addr_reg[0]/NET0131  ;
	input \P1_addr_reg[10]/NET0131  ;
	input \P1_addr_reg[11]/NET0131  ;
	input \P1_addr_reg[12]/NET0131  ;
	input \P1_addr_reg[13]/NET0131  ;
	input \P1_addr_reg[14]/NET0131  ;
	input \P1_addr_reg[15]/NET0131  ;
	input \P1_addr_reg[16]/NET0131  ;
	input \P1_addr_reg[17]/NET0131  ;
	input \P1_addr_reg[18]/NET0131  ;
	input \P1_addr_reg[19]/NET0131  ;
	input \P1_addr_reg[1]/NET0131  ;
	input \P1_addr_reg[2]/NET0131  ;
	input \P1_addr_reg[3]/NET0131  ;
	input \P1_addr_reg[4]/NET0131  ;
	input \P1_addr_reg[5]/NET0131  ;
	input \P1_addr_reg[6]/NET0131  ;
	input \P1_addr_reg[7]/NET0131  ;
	input \P1_addr_reg[8]/NET0131  ;
	input \P1_addr_reg[9]/NET0131  ;
	input \P1_d_reg[0]/NET0131  ;
	input \P1_d_reg[1]/NET0131  ;
	input \P1_datao_reg[0]/NET0131  ;
	input \P1_datao_reg[10]/NET0131  ;
	input \P1_datao_reg[11]/NET0131  ;
	input \P1_datao_reg[12]/NET0131  ;
	input \P1_datao_reg[13]/NET0131  ;
	input \P1_datao_reg[14]/NET0131  ;
	input \P1_datao_reg[15]/NET0131  ;
	input \P1_datao_reg[16]/NET0131  ;
	input \P1_datao_reg[17]/NET0131  ;
	input \P1_datao_reg[18]/NET0131  ;
	input \P1_datao_reg[19]/NET0131  ;
	input \P1_datao_reg[1]/NET0131  ;
	input \P1_datao_reg[20]/NET0131  ;
	input \P1_datao_reg[21]/NET0131  ;
	input \P1_datao_reg[22]/NET0131  ;
	input \P1_datao_reg[23]/NET0131  ;
	input \P1_datao_reg[24]/NET0131  ;
	input \P1_datao_reg[25]/NET0131  ;
	input \P1_datao_reg[26]/NET0131  ;
	input \P1_datao_reg[27]/NET0131  ;
	input \P1_datao_reg[28]/NET0131  ;
	input \P1_datao_reg[29]/NET0131  ;
	input \P1_datao_reg[2]/NET0131  ;
	input \P1_datao_reg[30]/NET0131  ;
	input \P1_datao_reg[31]/NET0131  ;
	input \P1_datao_reg[3]/NET0131  ;
	input \P1_datao_reg[4]/NET0131  ;
	input \P1_datao_reg[5]/NET0131  ;
	input \P1_datao_reg[6]/NET0131  ;
	input \P1_datao_reg[7]/NET0131  ;
	input \P1_datao_reg[8]/NET0131  ;
	input \P1_datao_reg[9]/NET0131  ;
	input \P1_rd_reg/NET0131  ;
	input \P1_reg0_reg[0]/NET0131  ;
	input \P1_reg0_reg[10]/NET0131  ;
	input \P1_reg0_reg[11]/NET0131  ;
	input \P1_reg0_reg[12]/NET0131  ;
	input \P1_reg0_reg[13]/NET0131  ;
	input \P1_reg0_reg[14]/NET0131  ;
	input \P1_reg0_reg[15]/NET0131  ;
	input \P1_reg0_reg[16]/NET0131  ;
	input \P1_reg0_reg[17]/NET0131  ;
	input \P1_reg0_reg[18]/NET0131  ;
	input \P1_reg0_reg[19]/NET0131  ;
	input \P1_reg0_reg[1]/NET0131  ;
	input \P1_reg0_reg[20]/NET0131  ;
	input \P1_reg0_reg[21]/NET0131  ;
	input \P1_reg0_reg[22]/NET0131  ;
	input \P1_reg0_reg[23]/NET0131  ;
	input \P1_reg0_reg[24]/NET0131  ;
	input \P1_reg0_reg[25]/NET0131  ;
	input \P1_reg0_reg[26]/NET0131  ;
	input \P1_reg0_reg[27]/NET0131  ;
	input \P1_reg0_reg[28]/NET0131  ;
	input \P1_reg0_reg[29]/NET0131  ;
	input \P1_reg0_reg[2]/NET0131  ;
	input \P1_reg0_reg[30]/NET0131  ;
	input \P1_reg0_reg[31]/NET0131  ;
	input \P1_reg0_reg[3]/NET0131  ;
	input \P1_reg0_reg[4]/NET0131  ;
	input \P1_reg0_reg[5]/NET0131  ;
	input \P1_reg0_reg[6]/NET0131  ;
	input \P1_reg0_reg[7]/NET0131  ;
	input \P1_reg0_reg[8]/NET0131  ;
	input \P1_reg0_reg[9]/NET0131  ;
	input \P1_reg1_reg[0]/NET0131  ;
	input \P1_reg1_reg[10]/NET0131  ;
	input \P1_reg1_reg[11]/NET0131  ;
	input \P1_reg1_reg[12]/NET0131  ;
	input \P1_reg1_reg[13]/NET0131  ;
	input \P1_reg1_reg[14]/NET0131  ;
	input \P1_reg1_reg[15]/NET0131  ;
	input \P1_reg1_reg[16]/NET0131  ;
	input \P1_reg1_reg[17]/NET0131  ;
	input \P1_reg1_reg[18]/NET0131  ;
	input \P1_reg1_reg[19]/NET0131  ;
	input \P1_reg1_reg[1]/NET0131  ;
	input \P1_reg1_reg[20]/NET0131  ;
	input \P1_reg1_reg[21]/NET0131  ;
	input \P1_reg1_reg[22]/NET0131  ;
	input \P1_reg1_reg[23]/NET0131  ;
	input \P1_reg1_reg[24]/NET0131  ;
	input \P1_reg1_reg[25]/NET0131  ;
	input \P1_reg1_reg[26]/NET0131  ;
	input \P1_reg1_reg[27]/NET0131  ;
	input \P1_reg1_reg[28]/NET0131  ;
	input \P1_reg1_reg[29]/NET0131  ;
	input \P1_reg1_reg[2]/NET0131  ;
	input \P1_reg1_reg[30]/NET0131  ;
	input \P1_reg1_reg[31]/NET0131  ;
	input \P1_reg1_reg[3]/NET0131  ;
	input \P1_reg1_reg[4]/NET0131  ;
	input \P1_reg1_reg[5]/NET0131  ;
	input \P1_reg1_reg[6]/NET0131  ;
	input \P1_reg1_reg[7]/NET0131  ;
	input \P1_reg1_reg[8]/NET0131  ;
	input \P1_reg1_reg[9]/NET0131  ;
	input \P1_reg2_reg[0]/NET0131  ;
	input \P1_reg2_reg[10]/NET0131  ;
	input \P1_reg2_reg[11]/NET0131  ;
	input \P1_reg2_reg[12]/NET0131  ;
	input \P1_reg2_reg[13]/NET0131  ;
	input \P1_reg2_reg[14]/NET0131  ;
	input \P1_reg2_reg[15]/NET0131  ;
	input \P1_reg2_reg[16]/NET0131  ;
	input \P1_reg2_reg[17]/NET0131  ;
	input \P1_reg2_reg[18]/NET0131  ;
	input \P1_reg2_reg[19]/NET0131  ;
	input \P1_reg2_reg[1]/NET0131  ;
	input \P1_reg2_reg[20]/NET0131  ;
	input \P1_reg2_reg[21]/NET0131  ;
	input \P1_reg2_reg[22]/NET0131  ;
	input \P1_reg2_reg[23]/NET0131  ;
	input \P1_reg2_reg[24]/NET0131  ;
	input \P1_reg2_reg[25]/NET0131  ;
	input \P1_reg2_reg[26]/NET0131  ;
	input \P1_reg2_reg[27]/NET0131  ;
	input \P1_reg2_reg[28]/NET0131  ;
	input \P1_reg2_reg[29]/NET0131  ;
	input \P1_reg2_reg[2]/NET0131  ;
	input \P1_reg2_reg[30]/NET0131  ;
	input \P1_reg2_reg[31]/NET0131  ;
	input \P1_reg2_reg[3]/NET0131  ;
	input \P1_reg2_reg[4]/NET0131  ;
	input \P1_reg2_reg[5]/NET0131  ;
	input \P1_reg2_reg[6]/NET0131  ;
	input \P1_reg2_reg[7]/NET0131  ;
	input \P1_reg2_reg[8]/NET0131  ;
	input \P1_reg2_reg[9]/NET0131  ;
	input \P1_reg3_reg[0]/NET0131  ;
	input \P1_reg3_reg[10]/NET0131  ;
	input \P1_reg3_reg[11]/NET0131  ;
	input \P1_reg3_reg[12]/NET0131  ;
	input \P1_reg3_reg[13]/NET0131  ;
	input \P1_reg3_reg[14]/NET0131  ;
	input \P1_reg3_reg[15]/NET0131  ;
	input \P1_reg3_reg[16]/NET0131  ;
	input \P1_reg3_reg[17]/NET0131  ;
	input \P1_reg3_reg[18]/NET0131  ;
	input \P1_reg3_reg[19]/NET0131  ;
	input \P1_reg3_reg[1]/NET0131  ;
	input \P1_reg3_reg[20]/NET0131  ;
	input \P1_reg3_reg[21]/NET0131  ;
	input \P1_reg3_reg[22]/NET0131  ;
	input \P1_reg3_reg[23]/NET0131  ;
	input \P1_reg3_reg[24]/NET0131  ;
	input \P1_reg3_reg[25]/NET0131  ;
	input \P1_reg3_reg[26]/NET0131  ;
	input \P1_reg3_reg[27]/NET0131  ;
	input \P1_reg3_reg[28]/NET0131  ;
	input \P1_reg3_reg[2]/NET0131  ;
	input \P1_reg3_reg[3]/NET0131  ;
	input \P1_reg3_reg[4]/NET0131  ;
	input \P1_reg3_reg[5]/NET0131  ;
	input \P1_reg3_reg[6]/NET0131  ;
	input \P1_reg3_reg[7]/NET0131  ;
	input \P1_reg3_reg[8]/NET0131  ;
	input \P1_reg3_reg[9]/NET0131  ;
	input \P1_state_reg[0]/NET0131  ;
	input \P1_wr_reg/NET0131  ;
	input \P2_B_reg/NET0131  ;
	input \P2_IR_reg[0]/NET0131  ;
	input \P2_IR_reg[10]/NET0131  ;
	input \P2_IR_reg[11]/NET0131  ;
	input \P2_IR_reg[12]/NET0131  ;
	input \P2_IR_reg[13]/NET0131  ;
	input \P2_IR_reg[14]/NET0131  ;
	input \P2_IR_reg[15]/NET0131  ;
	input \P2_IR_reg[16]/NET0131  ;
	input \P2_IR_reg[17]/NET0131  ;
	input \P2_IR_reg[18]/NET0131  ;
	input \P2_IR_reg[19]/NET0131  ;
	input \P2_IR_reg[1]/NET0131  ;
	input \P2_IR_reg[20]/NET0131  ;
	input \P2_IR_reg[21]/NET0131  ;
	input \P2_IR_reg[22]/NET0131  ;
	input \P2_IR_reg[23]/NET0131  ;
	input \P2_IR_reg[24]/NET0131  ;
	input \P2_IR_reg[25]/NET0131  ;
	input \P2_IR_reg[26]/NET0131  ;
	input \P2_IR_reg[27]/NET0131  ;
	input \P2_IR_reg[28]/NET0131  ;
	input \P2_IR_reg[29]/NET0131  ;
	input \P2_IR_reg[2]/NET0131  ;
	input \P2_IR_reg[30]/NET0131  ;
	input \P2_IR_reg[31]/NET0131  ;
	input \P2_IR_reg[3]/NET0131  ;
	input \P2_IR_reg[4]/NET0131  ;
	input \P2_IR_reg[5]/NET0131  ;
	input \P2_IR_reg[6]/NET0131  ;
	input \P2_IR_reg[7]/NET0131  ;
	input \P2_IR_reg[8]/NET0131  ;
	input \P2_IR_reg[9]/NET0131  ;
	input \P2_addr_reg[0]/NET0131  ;
	input \P2_addr_reg[10]/NET0131  ;
	input \P2_addr_reg[11]/NET0131  ;
	input \P2_addr_reg[12]/NET0131  ;
	input \P2_addr_reg[13]/NET0131  ;
	input \P2_addr_reg[14]/NET0131  ;
	input \P2_addr_reg[15]/NET0131  ;
	input \P2_addr_reg[16]/NET0131  ;
	input \P2_addr_reg[17]/NET0131  ;
	input \P2_addr_reg[18]/NET0131  ;
	input \P2_addr_reg[19]/NET0131  ;
	input \P2_addr_reg[1]/NET0131  ;
	input \P2_addr_reg[2]/NET0131  ;
	input \P2_addr_reg[3]/NET0131  ;
	input \P2_addr_reg[4]/NET0131  ;
	input \P2_addr_reg[5]/NET0131  ;
	input \P2_addr_reg[6]/NET0131  ;
	input \P2_addr_reg[7]/NET0131  ;
	input \P2_addr_reg[8]/NET0131  ;
	input \P2_addr_reg[9]/NET0131  ;
	input \P2_d_reg[0]/NET0131  ;
	input \P2_d_reg[1]/NET0131  ;
	input \P2_datao_reg[0]/NET0131  ;
	input \P2_datao_reg[10]/NET0131  ;
	input \P2_datao_reg[11]/NET0131  ;
	input \P2_datao_reg[12]/NET0131  ;
	input \P2_datao_reg[13]/NET0131  ;
	input \P2_datao_reg[14]/NET0131  ;
	input \P2_datao_reg[15]/NET0131  ;
	input \P2_datao_reg[16]/NET0131  ;
	input \P2_datao_reg[17]/NET0131  ;
	input \P2_datao_reg[18]/NET0131  ;
	input \P2_datao_reg[19]/NET0131  ;
	input \P2_datao_reg[1]/NET0131  ;
	input \P2_datao_reg[20]/NET0131  ;
	input \P2_datao_reg[21]/NET0131  ;
	input \P2_datao_reg[22]/NET0131  ;
	input \P2_datao_reg[23]/NET0131  ;
	input \P2_datao_reg[24]/NET0131  ;
	input \P2_datao_reg[25]/NET0131  ;
	input \P2_datao_reg[26]/NET0131  ;
	input \P2_datao_reg[27]/NET0131  ;
	input \P2_datao_reg[28]/NET0131  ;
	input \P2_datao_reg[29]/NET0131  ;
	input \P2_datao_reg[2]/NET0131  ;
	input \P2_datao_reg[30]/NET0131  ;
	input \P2_datao_reg[31]/NET0131  ;
	input \P2_datao_reg[3]/NET0131  ;
	input \P2_datao_reg[4]/NET0131  ;
	input \P2_datao_reg[5]/NET0131  ;
	input \P2_datao_reg[6]/NET0131  ;
	input \P2_datao_reg[7]/NET0131  ;
	input \P2_datao_reg[8]/NET0131  ;
	input \P2_datao_reg[9]/NET0131  ;
	input \P2_rd_reg/NET0131  ;
	input \P2_reg0_reg[0]/NET0131  ;
	input \P2_reg0_reg[10]/NET0131  ;
	input \P2_reg0_reg[11]/NET0131  ;
	input \P2_reg0_reg[12]/NET0131  ;
	input \P2_reg0_reg[13]/NET0131  ;
	input \P2_reg0_reg[14]/NET0131  ;
	input \P2_reg0_reg[15]/NET0131  ;
	input \P2_reg0_reg[16]/NET0131  ;
	input \P2_reg0_reg[17]/NET0131  ;
	input \P2_reg0_reg[18]/NET0131  ;
	input \P2_reg0_reg[19]/NET0131  ;
	input \P2_reg0_reg[1]/NET0131  ;
	input \P2_reg0_reg[20]/NET0131  ;
	input \P2_reg0_reg[21]/NET0131  ;
	input \P2_reg0_reg[22]/NET0131  ;
	input \P2_reg0_reg[23]/NET0131  ;
	input \P2_reg0_reg[24]/NET0131  ;
	input \P2_reg0_reg[25]/NET0131  ;
	input \P2_reg0_reg[26]/NET0131  ;
	input \P2_reg0_reg[27]/NET0131  ;
	input \P2_reg0_reg[28]/NET0131  ;
	input \P2_reg0_reg[29]/NET0131  ;
	input \P2_reg0_reg[2]/NET0131  ;
	input \P2_reg0_reg[30]/NET0131  ;
	input \P2_reg0_reg[31]/NET0131  ;
	input \P2_reg0_reg[3]/NET0131  ;
	input \P2_reg0_reg[4]/NET0131  ;
	input \P2_reg0_reg[5]/NET0131  ;
	input \P2_reg0_reg[6]/NET0131  ;
	input \P2_reg0_reg[7]/NET0131  ;
	input \P2_reg0_reg[8]/NET0131  ;
	input \P2_reg0_reg[9]/NET0131  ;
	input \P2_reg1_reg[0]/NET0131  ;
	input \P2_reg1_reg[10]/NET0131  ;
	input \P2_reg1_reg[11]/NET0131  ;
	input \P2_reg1_reg[12]/NET0131  ;
	input \P2_reg1_reg[13]/NET0131  ;
	input \P2_reg1_reg[14]/NET0131  ;
	input \P2_reg1_reg[15]/NET0131  ;
	input \P2_reg1_reg[16]/NET0131  ;
	input \P2_reg1_reg[17]/NET0131  ;
	input \P2_reg1_reg[18]/NET0131  ;
	input \P2_reg1_reg[19]/NET0131  ;
	input \P2_reg1_reg[1]/NET0131  ;
	input \P2_reg1_reg[20]/NET0131  ;
	input \P2_reg1_reg[21]/NET0131  ;
	input \P2_reg1_reg[22]/NET0131  ;
	input \P2_reg1_reg[23]/NET0131  ;
	input \P2_reg1_reg[24]/NET0131  ;
	input \P2_reg1_reg[25]/NET0131  ;
	input \P2_reg1_reg[26]/NET0131  ;
	input \P2_reg1_reg[27]/NET0131  ;
	input \P2_reg1_reg[28]/NET0131  ;
	input \P2_reg1_reg[29]/NET0131  ;
	input \P2_reg1_reg[2]/NET0131  ;
	input \P2_reg1_reg[30]/NET0131  ;
	input \P2_reg1_reg[31]/NET0131  ;
	input \P2_reg1_reg[3]/NET0131  ;
	input \P2_reg1_reg[4]/NET0131  ;
	input \P2_reg1_reg[5]/NET0131  ;
	input \P2_reg1_reg[6]/NET0131  ;
	input \P2_reg1_reg[7]/NET0131  ;
	input \P2_reg1_reg[8]/NET0131  ;
	input \P2_reg1_reg[9]/NET0131  ;
	input \P2_reg2_reg[0]/NET0131  ;
	input \P2_reg2_reg[10]/NET0131  ;
	input \P2_reg2_reg[11]/NET0131  ;
	input \P2_reg2_reg[12]/NET0131  ;
	input \P2_reg2_reg[13]/NET0131  ;
	input \P2_reg2_reg[14]/NET0131  ;
	input \P2_reg2_reg[15]/NET0131  ;
	input \P2_reg2_reg[16]/NET0131  ;
	input \P2_reg2_reg[17]/NET0131  ;
	input \P2_reg2_reg[18]/NET0131  ;
	input \P2_reg2_reg[19]/NET0131  ;
	input \P2_reg2_reg[1]/NET0131  ;
	input \P2_reg2_reg[20]/NET0131  ;
	input \P2_reg2_reg[21]/NET0131  ;
	input \P2_reg2_reg[22]/NET0131  ;
	input \P2_reg2_reg[23]/NET0131  ;
	input \P2_reg2_reg[24]/NET0131  ;
	input \P2_reg2_reg[25]/NET0131  ;
	input \P2_reg2_reg[26]/NET0131  ;
	input \P2_reg2_reg[27]/NET0131  ;
	input \P2_reg2_reg[28]/NET0131  ;
	input \P2_reg2_reg[29]/NET0131  ;
	input \P2_reg2_reg[2]/NET0131  ;
	input \P2_reg2_reg[30]/NET0131  ;
	input \P2_reg2_reg[31]/NET0131  ;
	input \P2_reg2_reg[3]/NET0131  ;
	input \P2_reg2_reg[4]/NET0131  ;
	input \P2_reg2_reg[5]/NET0131  ;
	input \P2_reg2_reg[6]/NET0131  ;
	input \P2_reg2_reg[7]/NET0131  ;
	input \P2_reg2_reg[8]/NET0131  ;
	input \P2_reg2_reg[9]/NET0131  ;
	input \P2_reg3_reg[0]/NET0131  ;
	input \P2_reg3_reg[10]/NET0131  ;
	input \P2_reg3_reg[11]/NET0131  ;
	input \P2_reg3_reg[12]/NET0131  ;
	input \P2_reg3_reg[13]/NET0131  ;
	input \P2_reg3_reg[14]/NET0131  ;
	input \P2_reg3_reg[15]/NET0131  ;
	input \P2_reg3_reg[16]/NET0131  ;
	input \P2_reg3_reg[17]/NET0131  ;
	input \P2_reg3_reg[18]/NET0131  ;
	input \P2_reg3_reg[19]/NET0131  ;
	input \P2_reg3_reg[1]/NET0131  ;
	input \P2_reg3_reg[20]/NET0131  ;
	input \P2_reg3_reg[21]/NET0131  ;
	input \P2_reg3_reg[22]/NET0131  ;
	input \P2_reg3_reg[23]/NET0131  ;
	input \P2_reg3_reg[24]/NET0131  ;
	input \P2_reg3_reg[25]/NET0131  ;
	input \P2_reg3_reg[26]/NET0131  ;
	input \P2_reg3_reg[27]/NET0131  ;
	input \P2_reg3_reg[28]/NET0131  ;
	input \P2_reg3_reg[2]/NET0131  ;
	input \P2_reg3_reg[3]/NET0131  ;
	input \P2_reg3_reg[4]/NET0131  ;
	input \P2_reg3_reg[5]/NET0131  ;
	input \P2_reg3_reg[6]/NET0131  ;
	input \P2_reg3_reg[7]/NET0131  ;
	input \P2_reg3_reg[8]/NET0131  ;
	input \P2_reg3_reg[9]/NET0131  ;
	input \P2_wr_reg/NET0131  ;
	input \si[0]_pad  ;
	input \si[10]_pad  ;
	input \si[11]_pad  ;
	input \si[12]_pad  ;
	input \si[13]_pad  ;
	input \si[14]_pad  ;
	input \si[15]_pad  ;
	input \si[16]_pad  ;
	input \si[17]_pad  ;
	input \si[18]_pad  ;
	input \si[19]_pad  ;
	input \si[1]_pad  ;
	input \si[20]_pad  ;
	input \si[21]_pad  ;
	input \si[22]_pad  ;
	input \si[23]_pad  ;
	input \si[24]_pad  ;
	input \si[25]_pad  ;
	input \si[26]_pad  ;
	input \si[27]_pad  ;
	input \si[28]_pad  ;
	input \si[29]_pad  ;
	input \si[2]_pad  ;
	input \si[30]_pad  ;
	input \si[31]_pad  ;
	input \si[3]_pad  ;
	input \si[4]_pad  ;
	input \si[5]_pad  ;
	input \si[6]_pad  ;
	input \si[7]_pad  ;
	input \si[8]_pad  ;
	input \si[9]_pad  ;
	output \P1_state_reg[0]/NET0131_syn_2  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g70791/_0_  ;
	output \g70792/_0_  ;
	output \g70793/_0_  ;
	output \g70794/_0_  ;
	output \g70795/_0_  ;
	output \g70796/_0_  ;
	output \g70813/_0_  ;
	output \g70814/_0_  ;
	output \g70848/_0_  ;
	output \g70849/_0_  ;
	output \g70850/_0_  ;
	output \g70851/_0_  ;
	output \g70852/_0_  ;
	output \g70856/_0_  ;
	output \g70857/_0_  ;
	output \g70858/_0_  ;
	output \g70859/_0_  ;
	output \g70860/_0_  ;
	output \g70861/_0_  ;
	output \g70862/_0_  ;
	output \g70896/_0_  ;
	output \g70902/_0_  ;
	output \g70903/_0_  ;
	output \g70904/_0_  ;
	output \g70906/_0_  ;
	output \g70907/_0_  ;
	output \g70908/_0_  ;
	output \g70909/_0_  ;
	output \g70910/_0_  ;
	output \g70911/_0_  ;
	output \g70912/_0_  ;
	output \g70913/_0_  ;
	output \g70914/_0_  ;
	output \g70915/_0_  ;
	output \g70916/_0_  ;
	output \g70917/_0_  ;
	output \g70918/_0_  ;
	output \g70919/_0_  ;
	output \g70920/_0_  ;
	output \g70921/_0_  ;
	output \g70922/_0_  ;
	output \g70923/_0_  ;
	output \g70924/_0_  ;
	output \g70925/_0_  ;
	output \g70926/_0_  ;
	output \g70927/_0_  ;
	output \g70987/_0_  ;
	output \g70988/_0_  ;
	output \g70989/_0_  ;
	output \g70990/_0_  ;
	output \g70991/_0_  ;
	output \g71006/_0_  ;
	output \g71007/_0_  ;
	output \g71009/_0_  ;
	output \g71010/_0_  ;
	output \g71011/_0_  ;
	output \g71012/_0_  ;
	output \g71013/_0_  ;
	output \g71014/_0_  ;
	output \g71015/_0_  ;
	output \g71016/_0_  ;
	output \g71017/_0_  ;
	output \g71018/_0_  ;
	output \g71019/_0_  ;
	output \g71020/_0_  ;
	output \g71021/_0_  ;
	output \g71022/_0_  ;
	output \g71023/_0_  ;
	output \g71090/_0_  ;
	output \g71091/_0_  ;
	output \g71092/_0_  ;
	output \g71093/_0_  ;
	output \g71094/_0_  ;
	output \g71125/_0_  ;
	output \g71130/_0_  ;
	output \g71131/_0_  ;
	output \g71132/_0_  ;
	output \g71133/_0_  ;
	output \g71134/_0_  ;
	output \g71135/_0_  ;
	output \g71136/_0_  ;
	output \g71137/_0_  ;
	output \g71138/_0_  ;
	output \g71139/_0_  ;
	output \g71140/_0_  ;
	output \g71141/_0_  ;
	output \g71142/_0_  ;
	output \g71143/_0_  ;
	output \g71144/_0_  ;
	output \g71145/_0_  ;
	output \g71150/_0_  ;
	output \g71151/_0_  ;
	output \g71152/_0_  ;
	output \g71153/_0_  ;
	output \g71154/_0_  ;
	output \g71155/_0_  ;
	output \g71156/_0_  ;
	output \g71157/_0_  ;
	output \g71158/_0_  ;
	output \g71230/_0_  ;
	output \g71231/_0_  ;
	output \g71232/_0_  ;
	output \g71233/_0_  ;
	output \g71234/_0_  ;
	output \g71235/_0_  ;
	output \g71236/_0_  ;
	output \g71238/_0_  ;
	output \g71239/_0_  ;
	output \g71270/_0_  ;
	output \g71275/_0_  ;
	output \g71276/_0_  ;
	output \g71277/_0_  ;
	output \g71278/_0_  ;
	output \g71279/_0_  ;
	output \g71280/_0_  ;
	output \g71281/_0_  ;
	output \g71282/_0_  ;
	output \g71283/_0_  ;
	output \g71284/_0_  ;
	output \g71285/_0_  ;
	output \g71286/_0_  ;
	output \g71287/_0_  ;
	output \g71288/_0_  ;
	output \g71289/_0_  ;
	output \g71290/_0_  ;
	output \g71291/_0_  ;
	output \g71292/_0_  ;
	output \g71293/_0_  ;
	output \g71294/_0_  ;
	output \g71295/_0_  ;
	output \g71296/_0_  ;
	output \g71297/_0_  ;
	output \g71298/_0_  ;
	output \g71299/_0_  ;
	output \g71300/_0_  ;
	output \g71301/_0_  ;
	output \g71302/_0_  ;
	output \g71303/_0_  ;
	output \g71304/_0_  ;
	output \g71305/_0_  ;
	output \g71306/_0_  ;
	output \g71307/_0_  ;
	output \g71382/_0_  ;
	output \g71384/_0_  ;
	output \g71385/_0_  ;
	output \g71387/_0_  ;
	output \g71388/_0_  ;
	output \g71389/_0_  ;
	output \g71439/_0_  ;
	output \g71440/_0_  ;
	output \g71441/_0_  ;
	output \g71442/_0_  ;
	output \g71443/_0_  ;
	output \g71444/_0_  ;
	output \g71445/_0_  ;
	output \g71446/_0_  ;
	output \g71447/_0_  ;
	output \g71448/_0_  ;
	output \g71449/_0_  ;
	output \g71450/_0_  ;
	output \g71451/_0_  ;
	output \g71452/_0_  ;
	output \g71453/_0_  ;
	output \g71454/_0_  ;
	output \g71455/_0_  ;
	output \g71456/_0_  ;
	output \g71457/_0_  ;
	output \g71458/_0_  ;
	output \g71459/_0_  ;
	output \g71460/_0_  ;
	output \g71461/_0_  ;
	output \g71536/_0_  ;
	output \g71537/_0_  ;
	output \g71538/_0_  ;
	output \g71540/_0_  ;
	output \g71541/_0_  ;
	output \g71542/_0_  ;
	output \g71602/_0_  ;
	output \g71604/_0_  ;
	output \g71610/_0_  ;
	output \g71611/_0_  ;
	output \g71618/_0_  ;
	output \g71619/_0_  ;
	output \g71620/_0_  ;
	output \g71621/_0_  ;
	output \g71622/_0_  ;
	output \g71623/_0_  ;
	output \g71624/_0_  ;
	output \g71625/_0_  ;
	output \g71626/_0_  ;
	output \g71627/_0_  ;
	output \g71629/_0_  ;
	output \g71630/_0_  ;
	output \g71631/_0_  ;
	output \g71632/_0_  ;
	output \g71633/_0_  ;
	output \g71634/_0_  ;
	output \g71635/_0_  ;
	output \g71636/_0_  ;
	output \g71710/_0_  ;
	output \g71711/_0_  ;
	output \g71782/_0_  ;
	output \g71785/_0_  ;
	output \g71786/_0_  ;
	output \g71787/_0_  ;
	output \g71788/_0_  ;
	output \g71789/_0_  ;
	output \g71790/_0_  ;
	output \g71791/_0_  ;
	output \g71792/_0_  ;
	output \g71793/_0_  ;
	output \g71794/_0_  ;
	output \g71795/_0_  ;
	output \g71796/_0_  ;
	output \g71797/_0_  ;
	output \g71798/_0_  ;
	output \g71799/_0_  ;
	output \g71883/_0_  ;
	output \g72000/_0_  ;
	output \g72001/_0_  ;
	output \g72002/_0_  ;
	output \g72003/_0_  ;
	output \g72004/_0_  ;
	output \g72005/_0_  ;
	output \g72236/_0_  ;
	output \g72237/_0_  ;
	output \g72238/_0_  ;
	output \g72239/_0_  ;
	output \g72240/_0_  ;
	output \g72372/_0_  ;
	output \g72376/_0_  ;
	output \g72383/_0_  ;
	output \g72561/_0_  ;
	output \g72562/_0_  ;
	output \g72563/_0_  ;
	output \g72564/_0_  ;
	output \g72970/_0_  ;
	output \g72980/_0_  ;
	output \g72981/_0_  ;
	output \g72982/_0_  ;
	output \g72983/_0_  ;
	output \g74234/_0_  ;
	output \g74260/_0_  ;
	output \g75086/_0_  ;
	output \g75087/_0_  ;
	output \g75088/_0_  ;
	output \g75089/_0_  ;
	output \g75091/_0_  ;
	output \g75092/_0_  ;
	output \g80304/_3_  ;
	output \g80305/_3_  ;
	output \g80306/_3_  ;
	output \g80307/_3_  ;
	output \g80308/_0_  ;
	output \g80309/_0_  ;
	output \g80815/_0_  ;
	output \g80816/_0_  ;
	output \g80817/_0_  ;
	output \g80818/_0_  ;
	output \g80819/_0_  ;
	output \g80820/_0_  ;
	output \g80821/_0_  ;
	output \g80822/_0_  ;
	output \g80823/_0_  ;
	output \g80824/_0_  ;
	output \g80825/_0_  ;
	output \g80826/_3_  ;
	output \g80827/_0_  ;
	output \g80828/_0_  ;
	output \g80829/_0_  ;
	output \g80830/_0_  ;
	output \g80831/_0_  ;
	output \g80832/_0_  ;
	output \g80833/_0_  ;
	output \g80834/_0_  ;
	output \g80835/_0_  ;
	output \g80836/_0_  ;
	output \g80837/_0_  ;
	output \g80838/_3_  ;
	output \g80839/_0_  ;
	output \g80840/_3_  ;
	output \g80841/_0_  ;
	output \g80859/_3_  ;
	output \g80860/_3_  ;
	output \g80861/_3_  ;
	output \g80862/_3_  ;
	output \g80863/_3_  ;
	output \g80864/_3_  ;
	output \g80865/_3_  ;
	output \g80866/_3_  ;
	output \g80867/_3_  ;
	output \g80868/_3_  ;
	output \g80869/_3_  ;
	output \g80870/_3_  ;
	output \g80871/_3_  ;
	output \g80872/_3_  ;
	output \g80873/_3_  ;
	output \g80874/_3_  ;
	output \g80875/_3_  ;
	output \g80876/_3_  ;
	output \g80877/_3_  ;
	output \g80878/_3_  ;
	output \g80879/_0_  ;
	output \g80880/_3_  ;
	output \g80881/_3_  ;
	output \g80882/_3_  ;
	output \g80883/_3_  ;
	output \g80884/_3_  ;
	output \g80885/_3_  ;
	output \g80886/_3_  ;
	output \g80888/_0_  ;
	output \g81262/_0_  ;
	output \g81278/_0_  ;
	output \g81884/_0_  ;
	output \g81893/_0_  ;
	output \g81896/_0_  ;
	output \g81897/_0_  ;
	output \g81898/_0_  ;
	output \g81899/_0_  ;
	output \g81900/_0_  ;
	output \g81901/_0_  ;
	output \g81902/_0_  ;
	output \g81903/_0_  ;
	output \g81904/_0_  ;
	output \g81905/_0_  ;
	output \g81906/_0_  ;
	output \g81907/_0_  ;
	output \g81908/_0_  ;
	output \g81909/_0_  ;
	output \g81910/_0_  ;
	output \g81911/_0_  ;
	output \g81923/_0_  ;
	output \g81924/_0_  ;
	output \g81925/_0_  ;
	output \g81926/_0_  ;
	output \g82414/_0_  ;
	output \g82532/_0_  ;
	output \g83134/_0_  ;
	output \g83135/_0_  ;
	output \g83141/_0_  ;
	output \g83142/_0_  ;
	output \g83145/_0_  ;
	output \g83146/_0_  ;
	output \g83147/_0_  ;
	output \g83148/_0_  ;
	output \g83152/_0_  ;
	output \g83153/_0_  ;
	output \g83154/_0_  ;
	output \g83155/_0_  ;
	output \g83156/_0_  ;
	output \g83157/_0_  ;
	output \g83158/_0_  ;
	output \g83159/_0_  ;
	output \g83164/_0_  ;
	output \g83165/_0_  ;
	output \g83177/_0_  ;
	output \g83178/_0_  ;
	output \g83409/_0_  ;
	output \g83411/_0_  ;
	output \g83807/u3_syn_4  ;
	output \g84138/u3_syn_4  ;
	output \g85062/_0_  ;
	output \g85079/_2_  ;
	output \g85113/_0_  ;
	output \g85121/_0_  ;
	output \g85594/_0_  ;
	output \g85663/_0_  ;
	output \g85669/_0_  ;
	output \g85749/_0_  ;
	output \g85784/_0_  ;
	output \g85809/_0_  ;
	output \g85817/_0_  ;
	output \g85828/_0_  ;
	output \g85845/_0_  ;
	output \g85851/_0_  ;
	output \g85858/_0_  ;
	output \g85871/_0_  ;
	output \g85882_dup/_0_  ;
	output \g85891/_0_  ;
	output \g85900/_0_  ;
	output \g85905/_0_  ;
	output \g85917/_0_  ;
	output \g85934/_0_  ;
	output \g85949/_0_  ;
	output \g85971/_0_  ;
	output \g85997/_0_  ;
	output \g86044/_0_  ;
	output \g86053/_0_  ;
	output \g86063/_0_  ;
	output \g86082/_0_  ;
	output \g86088/_0_  ;
	output \g86098/_0_  ;
	output \g86105/_0_  ;
	output \g86179/_0_  ;
	output \g86256_dup/_0_  ;
	output \g86264/_0_  ;
	output \g86273/_0_  ;
	output \g86281/_0_  ;
	output \g86288/_0_  ;
	output \g86297/_0_  ;
	output \g86304/_0_  ;
	output \g86310/_0_  ;
	output \g86320/_0_  ;
	output \g86328/_0_  ;
	output \g86339/_0_  ;
	output \g86353/_0_  ;
	output \g86360/_0_  ;
	output \g86368/_0_  ;
	output \g86373/_0_  ;
	output \g86385/_0_  ;
	output \g86392/_0_  ;
	output \g86399/_0_  ;
	output \g86421/_0_  ;
	output \g86432/_0_  ;
	output \g87592/_1__syn_2  ;
	output \g87632/_1_  ;
	output \g92847/_0_  ;
	output \g92957/_0_  ;
	output \g93056/_0_  ;
	output \g93289/_0_  ;
	output \g93538_dup95061/_0_  ;
	output \g93856/_0_  ;
	output \g93870/_0_  ;
	output \g94004/_0_  ;
	output \g94128/_0_  ;
	output \g94173/_0_  ;
	output \g94187/_0_  ;
	output \g94191/_0_  ;
	output \g94318/_0_  ;
	output \g94505/_0_  ;
	output rd_pad ;
	output \so[0]_pad  ;
	output \so[10]_pad  ;
	output \so[11]_pad  ;
	output \so[12]_pad  ;
	output \so[13]_pad  ;
	output \so[14]_pad  ;
	output \so[15]_pad  ;
	output \so[16]_pad  ;
	output \so[17]_pad  ;
	output \so[18]_pad  ;
	output \so[19]_pad  ;
	output \so[1]_pad  ;
	output \so[2]_pad  ;
	output \so[3]_pad  ;
	output \so[4]_pad  ;
	output \so[5]_pad  ;
	output \so[6]_pad  ;
	output \so[7]_pad  ;
	output \so[8]_pad  ;
	output \so[9]_pad  ;
	output wr_pad ;
	wire _w6603_ ;
	wire _w6602_ ;
	wire _w6601_ ;
	wire _w6600_ ;
	wire _w6599_ ;
	wire _w6598_ ;
	wire _w6597_ ;
	wire _w6596_ ;
	wire _w6595_ ;
	wire _w6594_ ;
	wire _w6593_ ;
	wire _w6592_ ;
	wire _w6591_ ;
	wire _w6590_ ;
	wire _w6589_ ;
	wire _w6588_ ;
	wire _w6587_ ;
	wire _w6586_ ;
	wire _w6585_ ;
	wire _w6584_ ;
	wire _w6583_ ;
	wire _w6582_ ;
	wire _w6581_ ;
	wire _w6580_ ;
	wire _w6579_ ;
	wire _w6578_ ;
	wire _w6577_ ;
	wire _w6576_ ;
	wire _w6575_ ;
	wire _w6574_ ;
	wire _w6573_ ;
	wire _w6572_ ;
	wire _w6571_ ;
	wire _w6570_ ;
	wire _w6569_ ;
	wire _w6568_ ;
	wire _w6567_ ;
	wire _w6566_ ;
	wire _w6565_ ;
	wire _w6564_ ;
	wire _w6563_ ;
	wire _w6562_ ;
	wire _w6561_ ;
	wire _w6560_ ;
	wire _w6559_ ;
	wire _w6558_ ;
	wire _w6557_ ;
	wire _w6556_ ;
	wire _w6555_ ;
	wire _w6554_ ;
	wire _w6553_ ;
	wire _w6552_ ;
	wire _w6551_ ;
	wire _w6550_ ;
	wire _w6549_ ;
	wire _w6548_ ;
	wire _w6547_ ;
	wire _w6546_ ;
	wire _w6545_ ;
	wire _w6544_ ;
	wire _w6543_ ;
	wire _w6542_ ;
	wire _w6541_ ;
	wire _w6540_ ;
	wire _w6539_ ;
	wire _w6538_ ;
	wire _w6537_ ;
	wire _w6536_ ;
	wire _w6535_ ;
	wire _w6534_ ;
	wire _w6533_ ;
	wire _w6532_ ;
	wire _w6531_ ;
	wire _w6530_ ;
	wire _w6529_ ;
	wire _w6528_ ;
	wire _w6527_ ;
	wire _w6526_ ;
	wire _w6525_ ;
	wire _w6524_ ;
	wire _w6523_ ;
	wire _w6522_ ;
	wire _w6521_ ;
	wire _w6520_ ;
	wire _w6519_ ;
	wire _w6518_ ;
	wire _w6517_ ;
	wire _w6516_ ;
	wire _w6515_ ;
	wire _w6514_ ;
	wire _w6513_ ;
	wire _w6512_ ;
	wire _w6511_ ;
	wire _w6510_ ;
	wire _w6509_ ;
	wire _w6508_ ;
	wire _w6507_ ;
	wire _w6506_ ;
	wire _w6505_ ;
	wire _w6504_ ;
	wire _w6503_ ;
	wire _w6502_ ;
	wire _w6501_ ;
	wire _w6500_ ;
	wire _w6499_ ;
	wire _w6498_ ;
	wire _w6497_ ;
	wire _w6496_ ;
	wire _w6495_ ;
	wire _w6494_ ;
	wire _w6493_ ;
	wire _w6492_ ;
	wire _w6491_ ;
	wire _w6490_ ;
	wire _w6489_ ;
	wire _w6488_ ;
	wire _w6487_ ;
	wire _w6486_ ;
	wire _w6485_ ;
	wire _w6484_ ;
	wire _w6483_ ;
	wire _w6482_ ;
	wire _w6481_ ;
	wire _w6480_ ;
	wire _w6479_ ;
	wire _w6478_ ;
	wire _w6477_ ;
	wire _w6476_ ;
	wire _w6475_ ;
	wire _w6474_ ;
	wire _w6473_ ;
	wire _w6472_ ;
	wire _w6471_ ;
	wire _w6470_ ;
	wire _w6469_ ;
	wire _w6468_ ;
	wire _w6467_ ;
	wire _w6466_ ;
	wire _w6465_ ;
	wire _w6464_ ;
	wire _w6463_ ;
	wire _w6462_ ;
	wire _w6461_ ;
	wire _w6460_ ;
	wire _w6459_ ;
	wire _w6458_ ;
	wire _w6457_ ;
	wire _w6456_ ;
	wire _w6455_ ;
	wire _w6454_ ;
	wire _w6453_ ;
	wire _w6452_ ;
	wire _w6451_ ;
	wire _w6450_ ;
	wire _w6449_ ;
	wire _w6448_ ;
	wire _w6447_ ;
	wire _w6446_ ;
	wire _w6445_ ;
	wire _w6444_ ;
	wire _w6443_ ;
	wire _w6442_ ;
	wire _w6441_ ;
	wire _w6440_ ;
	wire _w6439_ ;
	wire _w6438_ ;
	wire _w6437_ ;
	wire _w6436_ ;
	wire _w6435_ ;
	wire _w6434_ ;
	wire _w6433_ ;
	wire _w6432_ ;
	wire _w6431_ ;
	wire _w6430_ ;
	wire _w6429_ ;
	wire _w6428_ ;
	wire _w6427_ ;
	wire _w6426_ ;
	wire _w6425_ ;
	wire _w6424_ ;
	wire _w6423_ ;
	wire _w6422_ ;
	wire _w6421_ ;
	wire _w6420_ ;
	wire _w6419_ ;
	wire _w6418_ ;
	wire _w6417_ ;
	wire _w6416_ ;
	wire _w6415_ ;
	wire _w6414_ ;
	wire _w6413_ ;
	wire _w6412_ ;
	wire _w6411_ ;
	wire _w6410_ ;
	wire _w6409_ ;
	wire _w6408_ ;
	wire _w6407_ ;
	wire _w6406_ ;
	wire _w6405_ ;
	wire _w6404_ ;
	wire _w6403_ ;
	wire _w6402_ ;
	wire _w6401_ ;
	wire _w6400_ ;
	wire _w6399_ ;
	wire _w6398_ ;
	wire _w6397_ ;
	wire _w6396_ ;
	wire _w6395_ ;
	wire _w6394_ ;
	wire _w6393_ ;
	wire _w6392_ ;
	wire _w6391_ ;
	wire _w6390_ ;
	wire _w6389_ ;
	wire _w6388_ ;
	wire _w6387_ ;
	wire _w6386_ ;
	wire _w6385_ ;
	wire _w6384_ ;
	wire _w6383_ ;
	wire _w6382_ ;
	wire _w6381_ ;
	wire _w6380_ ;
	wire _w6379_ ;
	wire _w6378_ ;
	wire _w6377_ ;
	wire _w6376_ ;
	wire _w6375_ ;
	wire _w6374_ ;
	wire _w6373_ ;
	wire _w6372_ ;
	wire _w6371_ ;
	wire _w6370_ ;
	wire _w6369_ ;
	wire _w6368_ ;
	wire _w6367_ ;
	wire _w6366_ ;
	wire _w6365_ ;
	wire _w6364_ ;
	wire _w6363_ ;
	wire _w6362_ ;
	wire _w6361_ ;
	wire _w6360_ ;
	wire _w6359_ ;
	wire _w6358_ ;
	wire _w6357_ ;
	wire _w6356_ ;
	wire _w6355_ ;
	wire _w6354_ ;
	wire _w6353_ ;
	wire _w6352_ ;
	wire _w6351_ ;
	wire _w6350_ ;
	wire _w6349_ ;
	wire _w6348_ ;
	wire _w6347_ ;
	wire _w6346_ ;
	wire _w6345_ ;
	wire _w6344_ ;
	wire _w6343_ ;
	wire _w6342_ ;
	wire _w6341_ ;
	wire _w6340_ ;
	wire _w6339_ ;
	wire _w6338_ ;
	wire _w6337_ ;
	wire _w6336_ ;
	wire _w6335_ ;
	wire _w6334_ ;
	wire _w6333_ ;
	wire _w6332_ ;
	wire _w6331_ ;
	wire _w6330_ ;
	wire _w6329_ ;
	wire _w6328_ ;
	wire _w6327_ ;
	wire _w6326_ ;
	wire _w6325_ ;
	wire _w6324_ ;
	wire _w6323_ ;
	wire _w6322_ ;
	wire _w6321_ ;
	wire _w6320_ ;
	wire _w6319_ ;
	wire _w6318_ ;
	wire _w6317_ ;
	wire _w6316_ ;
	wire _w6315_ ;
	wire _w6314_ ;
	wire _w6313_ ;
	wire _w6312_ ;
	wire _w6311_ ;
	wire _w6310_ ;
	wire _w6309_ ;
	wire _w6308_ ;
	wire _w6307_ ;
	wire _w6306_ ;
	wire _w6305_ ;
	wire _w6304_ ;
	wire _w6303_ ;
	wire _w6302_ ;
	wire _w6301_ ;
	wire _w6300_ ;
	wire _w6299_ ;
	wire _w6298_ ;
	wire _w6297_ ;
	wire _w6296_ ;
	wire _w6295_ ;
	wire _w6294_ ;
	wire _w6293_ ;
	wire _w6292_ ;
	wire _w6291_ ;
	wire _w6290_ ;
	wire _w6289_ ;
	wire _w6288_ ;
	wire _w6287_ ;
	wire _w6286_ ;
	wire _w6285_ ;
	wire _w6284_ ;
	wire _w6283_ ;
	wire _w6282_ ;
	wire _w6281_ ;
	wire _w6280_ ;
	wire _w6279_ ;
	wire _w6278_ ;
	wire _w6277_ ;
	wire _w6276_ ;
	wire _w6275_ ;
	wire _w6274_ ;
	wire _w6273_ ;
	wire _w6272_ ;
	wire _w6271_ ;
	wire _w6270_ ;
	wire _w6269_ ;
	wire _w6268_ ;
	wire _w6267_ ;
	wire _w6266_ ;
	wire _w6265_ ;
	wire _w6264_ ;
	wire _w6263_ ;
	wire _w6262_ ;
	wire _w6261_ ;
	wire _w6260_ ;
	wire _w6259_ ;
	wire _w6258_ ;
	wire _w6257_ ;
	wire _w6256_ ;
	wire _w6255_ ;
	wire _w6254_ ;
	wire _w6253_ ;
	wire _w6252_ ;
	wire _w6251_ ;
	wire _w6250_ ;
	wire _w6249_ ;
	wire _w6248_ ;
	wire _w6247_ ;
	wire _w6246_ ;
	wire _w6245_ ;
	wire _w6244_ ;
	wire _w6243_ ;
	wire _w6242_ ;
	wire _w6241_ ;
	wire _w6240_ ;
	wire _w6239_ ;
	wire _w6238_ ;
	wire _w6237_ ;
	wire _w6236_ ;
	wire _w6235_ ;
	wire _w6234_ ;
	wire _w6233_ ;
	wire _w6232_ ;
	wire _w6231_ ;
	wire _w6230_ ;
	wire _w6229_ ;
	wire _w6228_ ;
	wire _w6227_ ;
	wire _w6226_ ;
	wire _w6225_ ;
	wire _w6224_ ;
	wire _w6223_ ;
	wire _w6222_ ;
	wire _w6221_ ;
	wire _w6220_ ;
	wire _w6219_ ;
	wire _w6218_ ;
	wire _w6217_ ;
	wire _w6216_ ;
	wire _w6215_ ;
	wire _w6214_ ;
	wire _w6213_ ;
	wire _w6212_ ;
	wire _w6211_ ;
	wire _w6210_ ;
	wire _w6209_ ;
	wire _w6208_ ;
	wire _w6207_ ;
	wire _w6206_ ;
	wire _w6205_ ;
	wire _w6204_ ;
	wire _w6203_ ;
	wire _w6202_ ;
	wire _w6201_ ;
	wire _w6200_ ;
	wire _w6199_ ;
	wire _w6198_ ;
	wire _w6197_ ;
	wire _w6196_ ;
	wire _w6195_ ;
	wire _w6194_ ;
	wire _w6193_ ;
	wire _w6192_ ;
	wire _w6191_ ;
	wire _w6190_ ;
	wire _w6189_ ;
	wire _w6188_ ;
	wire _w6187_ ;
	wire _w6186_ ;
	wire _w6185_ ;
	wire _w6184_ ;
	wire _w6183_ ;
	wire _w6182_ ;
	wire _w6181_ ;
	wire _w6180_ ;
	wire _w6179_ ;
	wire _w6178_ ;
	wire _w6177_ ;
	wire _w6176_ ;
	wire _w6175_ ;
	wire _w6174_ ;
	wire _w6173_ ;
	wire _w6172_ ;
	wire _w6171_ ;
	wire _w6170_ ;
	wire _w6169_ ;
	wire _w6168_ ;
	wire _w6167_ ;
	wire _w6166_ ;
	wire _w6165_ ;
	wire _w6164_ ;
	wire _w6163_ ;
	wire _w6162_ ;
	wire _w6161_ ;
	wire _w6160_ ;
	wire _w6159_ ;
	wire _w6158_ ;
	wire _w6157_ ;
	wire _w6156_ ;
	wire _w6155_ ;
	wire _w6154_ ;
	wire _w6153_ ;
	wire _w6152_ ;
	wire _w6151_ ;
	wire _w6150_ ;
	wire _w6149_ ;
	wire _w6148_ ;
	wire _w6147_ ;
	wire _w6146_ ;
	wire _w6145_ ;
	wire _w6144_ ;
	wire _w6143_ ;
	wire _w6142_ ;
	wire _w6141_ ;
	wire _w6140_ ;
	wire _w6139_ ;
	wire _w6138_ ;
	wire _w6137_ ;
	wire _w6136_ ;
	wire _w6135_ ;
	wire _w6134_ ;
	wire _w6133_ ;
	wire _w6132_ ;
	wire _w6131_ ;
	wire _w6130_ ;
	wire _w6129_ ;
	wire _w6128_ ;
	wire _w6127_ ;
	wire _w6126_ ;
	wire _w6125_ ;
	wire _w6124_ ;
	wire _w6123_ ;
	wire _w6122_ ;
	wire _w6121_ ;
	wire _w6120_ ;
	wire _w6119_ ;
	wire _w6118_ ;
	wire _w6117_ ;
	wire _w6116_ ;
	wire _w6115_ ;
	wire _w6114_ ;
	wire _w6113_ ;
	wire _w6112_ ;
	wire _w6111_ ;
	wire _w6110_ ;
	wire _w6109_ ;
	wire _w6108_ ;
	wire _w6107_ ;
	wire _w6106_ ;
	wire _w6105_ ;
	wire _w6104_ ;
	wire _w6103_ ;
	wire _w6102_ ;
	wire _w6101_ ;
	wire _w6100_ ;
	wire _w6099_ ;
	wire _w6098_ ;
	wire _w6097_ ;
	wire _w6096_ ;
	wire _w6095_ ;
	wire _w6094_ ;
	wire _w6093_ ;
	wire _w6092_ ;
	wire _w6091_ ;
	wire _w6090_ ;
	wire _w6089_ ;
	wire _w6088_ ;
	wire _w6087_ ;
	wire _w6086_ ;
	wire _w6085_ ;
	wire _w6084_ ;
	wire _w6083_ ;
	wire _w6082_ ;
	wire _w6081_ ;
	wire _w6080_ ;
	wire _w6079_ ;
	wire _w6078_ ;
	wire _w6077_ ;
	wire _w6076_ ;
	wire _w6075_ ;
	wire _w6074_ ;
	wire _w6073_ ;
	wire _w6072_ ;
	wire _w6071_ ;
	wire _w6070_ ;
	wire _w6069_ ;
	wire _w6068_ ;
	wire _w6067_ ;
	wire _w6066_ ;
	wire _w6065_ ;
	wire _w6064_ ;
	wire _w6063_ ;
	wire _w6062_ ;
	wire _w6061_ ;
	wire _w6060_ ;
	wire _w6059_ ;
	wire _w6058_ ;
	wire _w6057_ ;
	wire _w6056_ ;
	wire _w6055_ ;
	wire _w6054_ ;
	wire _w6053_ ;
	wire _w6052_ ;
	wire _w6051_ ;
	wire _w6050_ ;
	wire _w6049_ ;
	wire _w6048_ ;
	wire _w6047_ ;
	wire _w6046_ ;
	wire _w6045_ ;
	wire _w6044_ ;
	wire _w6043_ ;
	wire _w6042_ ;
	wire _w6041_ ;
	wire _w6040_ ;
	wire _w6039_ ;
	wire _w6038_ ;
	wire _w6037_ ;
	wire _w6036_ ;
	wire _w6035_ ;
	wire _w6034_ ;
	wire _w6033_ ;
	wire _w6032_ ;
	wire _w6031_ ;
	wire _w6030_ ;
	wire _w6029_ ;
	wire _w6028_ ;
	wire _w6027_ ;
	wire _w6026_ ;
	wire _w6025_ ;
	wire _w6024_ ;
	wire _w6023_ ;
	wire _w6022_ ;
	wire _w6021_ ;
	wire _w6020_ ;
	wire _w6019_ ;
	wire _w6018_ ;
	wire _w6017_ ;
	wire _w6016_ ;
	wire _w6015_ ;
	wire _w6014_ ;
	wire _w6013_ ;
	wire _w6012_ ;
	wire _w6011_ ;
	wire _w6010_ ;
	wire _w6009_ ;
	wire _w6008_ ;
	wire _w6007_ ;
	wire _w6006_ ;
	wire _w6005_ ;
	wire _w6004_ ;
	wire _w6003_ ;
	wire _w6002_ ;
	wire _w6001_ ;
	wire _w6000_ ;
	wire _w5999_ ;
	wire _w5998_ ;
	wire _w5997_ ;
	wire _w5996_ ;
	wire _w5995_ ;
	wire _w5994_ ;
	wire _w5993_ ;
	wire _w5992_ ;
	wire _w5991_ ;
	wire _w5990_ ;
	wire _w5989_ ;
	wire _w5988_ ;
	wire _w5987_ ;
	wire _w5986_ ;
	wire _w5985_ ;
	wire _w5984_ ;
	wire _w5983_ ;
	wire _w5982_ ;
	wire _w5981_ ;
	wire _w5980_ ;
	wire _w5979_ ;
	wire _w5978_ ;
	wire _w5977_ ;
	wire _w5976_ ;
	wire _w5975_ ;
	wire _w5974_ ;
	wire _w5973_ ;
	wire _w5972_ ;
	wire _w5971_ ;
	wire _w5970_ ;
	wire _w5969_ ;
	wire _w5968_ ;
	wire _w5967_ ;
	wire _w5966_ ;
	wire _w5965_ ;
	wire _w5964_ ;
	wire _w5963_ ;
	wire _w5962_ ;
	wire _w5961_ ;
	wire _w5960_ ;
	wire _w5959_ ;
	wire _w5958_ ;
	wire _w5957_ ;
	wire _w5956_ ;
	wire _w5955_ ;
	wire _w5954_ ;
	wire _w5953_ ;
	wire _w5952_ ;
	wire _w5951_ ;
	wire _w5950_ ;
	wire _w5949_ ;
	wire _w5948_ ;
	wire _w5947_ ;
	wire _w5946_ ;
	wire _w5945_ ;
	wire _w5944_ ;
	wire _w5943_ ;
	wire _w5942_ ;
	wire _w5941_ ;
	wire _w5940_ ;
	wire _w5939_ ;
	wire _w5938_ ;
	wire _w5937_ ;
	wire _w5936_ ;
	wire _w5935_ ;
	wire _w5934_ ;
	wire _w5933_ ;
	wire _w5932_ ;
	wire _w5931_ ;
	wire _w5930_ ;
	wire _w5929_ ;
	wire _w5928_ ;
	wire _w5927_ ;
	wire _w5926_ ;
	wire _w5925_ ;
	wire _w5924_ ;
	wire _w5923_ ;
	wire _w5922_ ;
	wire _w5921_ ;
	wire _w5920_ ;
	wire _w5919_ ;
	wire _w5918_ ;
	wire _w5917_ ;
	wire _w5916_ ;
	wire _w5915_ ;
	wire _w5914_ ;
	wire _w5913_ ;
	wire _w5912_ ;
	wire _w5911_ ;
	wire _w5910_ ;
	wire _w5909_ ;
	wire _w5908_ ;
	wire _w5907_ ;
	wire _w5906_ ;
	wire _w5905_ ;
	wire _w5904_ ;
	wire _w5903_ ;
	wire _w5902_ ;
	wire _w5901_ ;
	wire _w5900_ ;
	wire _w5899_ ;
	wire _w5898_ ;
	wire _w5897_ ;
	wire _w5896_ ;
	wire _w5895_ ;
	wire _w5894_ ;
	wire _w5893_ ;
	wire _w5892_ ;
	wire _w5891_ ;
	wire _w5890_ ;
	wire _w5889_ ;
	wire _w5888_ ;
	wire _w5887_ ;
	wire _w5886_ ;
	wire _w5885_ ;
	wire _w5884_ ;
	wire _w5883_ ;
	wire _w5882_ ;
	wire _w5881_ ;
	wire _w5880_ ;
	wire _w5879_ ;
	wire _w5878_ ;
	wire _w5877_ ;
	wire _w5876_ ;
	wire _w5875_ ;
	wire _w5874_ ;
	wire _w5873_ ;
	wire _w5872_ ;
	wire _w5871_ ;
	wire _w5870_ ;
	wire _w5869_ ;
	wire _w5868_ ;
	wire _w5867_ ;
	wire _w5866_ ;
	wire _w5865_ ;
	wire _w5864_ ;
	wire _w5863_ ;
	wire _w5862_ ;
	wire _w5861_ ;
	wire _w5860_ ;
	wire _w5859_ ;
	wire _w5858_ ;
	wire _w5857_ ;
	wire _w5856_ ;
	wire _w5855_ ;
	wire _w5854_ ;
	wire _w5853_ ;
	wire _w5852_ ;
	wire _w5851_ ;
	wire _w5850_ ;
	wire _w5849_ ;
	wire _w5848_ ;
	wire _w5847_ ;
	wire _w5846_ ;
	wire _w5845_ ;
	wire _w5844_ ;
	wire _w5843_ ;
	wire _w5842_ ;
	wire _w5841_ ;
	wire _w5840_ ;
	wire _w5839_ ;
	wire _w5838_ ;
	wire _w5837_ ;
	wire _w5836_ ;
	wire _w5835_ ;
	wire _w5834_ ;
	wire _w5833_ ;
	wire _w5832_ ;
	wire _w5831_ ;
	wire _w5830_ ;
	wire _w5829_ ;
	wire _w5828_ ;
	wire _w5827_ ;
	wire _w5826_ ;
	wire _w5825_ ;
	wire _w5824_ ;
	wire _w5823_ ;
	wire _w5822_ ;
	wire _w5821_ ;
	wire _w5820_ ;
	wire _w5819_ ;
	wire _w5818_ ;
	wire _w5817_ ;
	wire _w5816_ ;
	wire _w5815_ ;
	wire _w5814_ ;
	wire _w5813_ ;
	wire _w5812_ ;
	wire _w5811_ ;
	wire _w5810_ ;
	wire _w5809_ ;
	wire _w5808_ ;
	wire _w5807_ ;
	wire _w5806_ ;
	wire _w5805_ ;
	wire _w5804_ ;
	wire _w5803_ ;
	wire _w5802_ ;
	wire _w5801_ ;
	wire _w5800_ ;
	wire _w5799_ ;
	wire _w5798_ ;
	wire _w5797_ ;
	wire _w5796_ ;
	wire _w5795_ ;
	wire _w5794_ ;
	wire _w5793_ ;
	wire _w5792_ ;
	wire _w5791_ ;
	wire _w5790_ ;
	wire _w5789_ ;
	wire _w5788_ ;
	wire _w5787_ ;
	wire _w5786_ ;
	wire _w5785_ ;
	wire _w5784_ ;
	wire _w5783_ ;
	wire _w5782_ ;
	wire _w5781_ ;
	wire _w5780_ ;
	wire _w5779_ ;
	wire _w5778_ ;
	wire _w5777_ ;
	wire _w5776_ ;
	wire _w5775_ ;
	wire _w5774_ ;
	wire _w5773_ ;
	wire _w5772_ ;
	wire _w5771_ ;
	wire _w5770_ ;
	wire _w5769_ ;
	wire _w5768_ ;
	wire _w5767_ ;
	wire _w5766_ ;
	wire _w5765_ ;
	wire _w5764_ ;
	wire _w5763_ ;
	wire _w5762_ ;
	wire _w5761_ ;
	wire _w5760_ ;
	wire _w5759_ ;
	wire _w5758_ ;
	wire _w5757_ ;
	wire _w5756_ ;
	wire _w5755_ ;
	wire _w5754_ ;
	wire _w5753_ ;
	wire _w5752_ ;
	wire _w5751_ ;
	wire _w5750_ ;
	wire _w5749_ ;
	wire _w5748_ ;
	wire _w5747_ ;
	wire _w5746_ ;
	wire _w5745_ ;
	wire _w5744_ ;
	wire _w5743_ ;
	wire _w5742_ ;
	wire _w5741_ ;
	wire _w5740_ ;
	wire _w5739_ ;
	wire _w5738_ ;
	wire _w5737_ ;
	wire _w5736_ ;
	wire _w5735_ ;
	wire _w5734_ ;
	wire _w5733_ ;
	wire _w5732_ ;
	wire _w5731_ ;
	wire _w5730_ ;
	wire _w5729_ ;
	wire _w5728_ ;
	wire _w5727_ ;
	wire _w5726_ ;
	wire _w5725_ ;
	wire _w5724_ ;
	wire _w5723_ ;
	wire _w5722_ ;
	wire _w5721_ ;
	wire _w5720_ ;
	wire _w5719_ ;
	wire _w5718_ ;
	wire _w5717_ ;
	wire _w5716_ ;
	wire _w5715_ ;
	wire _w5714_ ;
	wire _w5713_ ;
	wire _w5712_ ;
	wire _w5711_ ;
	wire _w5710_ ;
	wire _w5709_ ;
	wire _w5708_ ;
	wire _w5707_ ;
	wire _w5706_ ;
	wire _w5705_ ;
	wire _w5704_ ;
	wire _w5703_ ;
	wire _w5702_ ;
	wire _w5701_ ;
	wire _w5700_ ;
	wire _w5699_ ;
	wire _w5698_ ;
	wire _w5697_ ;
	wire _w5696_ ;
	wire _w5695_ ;
	wire _w5694_ ;
	wire _w5693_ ;
	wire _w5692_ ;
	wire _w5691_ ;
	wire _w5690_ ;
	wire _w5689_ ;
	wire _w5688_ ;
	wire _w5687_ ;
	wire _w5686_ ;
	wire _w5685_ ;
	wire _w5684_ ;
	wire _w5683_ ;
	wire _w5682_ ;
	wire _w5681_ ;
	wire _w5680_ ;
	wire _w5679_ ;
	wire _w5678_ ;
	wire _w5677_ ;
	wire _w5676_ ;
	wire _w5675_ ;
	wire _w5674_ ;
	wire _w5673_ ;
	wire _w5672_ ;
	wire _w5671_ ;
	wire _w5670_ ;
	wire _w5669_ ;
	wire _w5668_ ;
	wire _w5667_ ;
	wire _w5666_ ;
	wire _w5665_ ;
	wire _w5664_ ;
	wire _w5663_ ;
	wire _w5662_ ;
	wire _w5661_ ;
	wire _w5660_ ;
	wire _w5659_ ;
	wire _w5658_ ;
	wire _w5657_ ;
	wire _w5656_ ;
	wire _w5655_ ;
	wire _w5654_ ;
	wire _w5653_ ;
	wire _w5652_ ;
	wire _w5651_ ;
	wire _w5650_ ;
	wire _w5649_ ;
	wire _w5648_ ;
	wire _w5647_ ;
	wire _w5646_ ;
	wire _w5645_ ;
	wire _w5644_ ;
	wire _w5643_ ;
	wire _w5642_ ;
	wire _w5641_ ;
	wire _w5640_ ;
	wire _w5639_ ;
	wire _w5638_ ;
	wire _w5637_ ;
	wire _w5636_ ;
	wire _w5635_ ;
	wire _w5634_ ;
	wire _w5633_ ;
	wire _w5632_ ;
	wire _w5631_ ;
	wire _w5630_ ;
	wire _w5629_ ;
	wire _w5628_ ;
	wire _w5627_ ;
	wire _w5626_ ;
	wire _w5625_ ;
	wire _w5624_ ;
	wire _w5623_ ;
	wire _w5622_ ;
	wire _w5621_ ;
	wire _w5620_ ;
	wire _w5619_ ;
	wire _w5618_ ;
	wire _w5617_ ;
	wire _w5616_ ;
	wire _w5615_ ;
	wire _w5614_ ;
	wire _w5613_ ;
	wire _w5612_ ;
	wire _w5611_ ;
	wire _w5610_ ;
	wire _w5609_ ;
	wire _w5608_ ;
	wire _w5607_ ;
	wire _w5606_ ;
	wire _w5605_ ;
	wire _w5604_ ;
	wire _w5603_ ;
	wire _w5602_ ;
	wire _w5601_ ;
	wire _w5600_ ;
	wire _w5599_ ;
	wire _w5598_ ;
	wire _w5597_ ;
	wire _w5596_ ;
	wire _w5595_ ;
	wire _w5594_ ;
	wire _w5593_ ;
	wire _w5592_ ;
	wire _w5591_ ;
	wire _w5590_ ;
	wire _w5589_ ;
	wire _w5588_ ;
	wire _w5587_ ;
	wire _w5586_ ;
	wire _w5585_ ;
	wire _w5584_ ;
	wire _w5583_ ;
	wire _w5582_ ;
	wire _w5581_ ;
	wire _w5580_ ;
	wire _w5579_ ;
	wire _w5578_ ;
	wire _w5577_ ;
	wire _w5576_ ;
	wire _w5575_ ;
	wire _w5574_ ;
	wire _w5573_ ;
	wire _w5572_ ;
	wire _w5571_ ;
	wire _w5570_ ;
	wire _w5569_ ;
	wire _w5568_ ;
	wire _w5567_ ;
	wire _w5566_ ;
	wire _w5565_ ;
	wire _w5564_ ;
	wire _w5563_ ;
	wire _w5562_ ;
	wire _w5561_ ;
	wire _w5560_ ;
	wire _w5559_ ;
	wire _w5558_ ;
	wire _w5557_ ;
	wire _w5556_ ;
	wire _w5555_ ;
	wire _w5554_ ;
	wire _w5553_ ;
	wire _w5552_ ;
	wire _w5551_ ;
	wire _w5550_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w2809_ ;
	wire _w2808_ ;
	wire _w2807_ ;
	wire _w2806_ ;
	wire _w2805_ ;
	wire _w2804_ ;
	wire _w2803_ ;
	wire _w2802_ ;
	wire _w2801_ ;
	wire _w2800_ ;
	wire _w2799_ ;
	wire _w2798_ ;
	wire _w2797_ ;
	wire _w2796_ ;
	wire _w2795_ ;
	wire _w2794_ ;
	wire _w2793_ ;
	wire _w2792_ ;
	wire _w2791_ ;
	wire _w2790_ ;
	wire _w2789_ ;
	wire _w2788_ ;
	wire _w2787_ ;
	wire _w2786_ ;
	wire _w2785_ ;
	wire _w2784_ ;
	wire _w2783_ ;
	wire _w2782_ ;
	wire _w2781_ ;
	wire _w2780_ ;
	wire _w2779_ ;
	wire _w2778_ ;
	wire _w2777_ ;
	wire _w2776_ ;
	wire _w2775_ ;
	wire _w2774_ ;
	wire _w2773_ ;
	wire _w2772_ ;
	wire _w2771_ ;
	wire _w2770_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2485_ ;
	wire _w2484_ ;
	wire _w2483_ ;
	wire _w2482_ ;
	wire _w2481_ ;
	wire _w2480_ ;
	wire _w2479_ ;
	wire _w2478_ ;
	wire _w2477_ ;
	wire _w2476_ ;
	wire _w2475_ ;
	wire _w2474_ ;
	wire _w2473_ ;
	wire _w2472_ ;
	wire _w2471_ ;
	wire _w2470_ ;
	wire _w2469_ ;
	wire _w2468_ ;
	wire _w2467_ ;
	wire _w2466_ ;
	wire _w2465_ ;
	wire _w2464_ ;
	wire _w2463_ ;
	wire _w2462_ ;
	wire _w2461_ ;
	wire _w2460_ ;
	wire _w2459_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w511_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w757_ ;
	wire _w2573_ ;
	wire _w216_ ;
	wire _w5303_ ;
	wire _w1325_ ;
	wire _w473_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w1501_ ;
	wire _w1502_ ;
	wire _w1503_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3177_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3195_ ;
	wire _w3196_ ;
	wire _w3197_ ;
	wire _w3198_ ;
	wire _w3199_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3202_ ;
	wire _w3203_ ;
	wire _w3204_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3210_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3217_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w3255_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w3338_ ;
	wire _w3339_ ;
	wire _w3340_ ;
	wire _w3341_ ;
	wire _w3342_ ;
	wire _w3343_ ;
	wire _w3344_ ;
	wire _w3345_ ;
	wire _w3346_ ;
	wire _w3347_ ;
	wire _w3348_ ;
	wire _w3349_ ;
	wire _w3350_ ;
	wire _w3351_ ;
	wire _w3352_ ;
	wire _w3353_ ;
	wire _w3354_ ;
	wire _w3355_ ;
	wire _w3356_ ;
	wire _w3357_ ;
	wire _w3358_ ;
	wire _w3359_ ;
	wire _w3360_ ;
	wire _w3361_ ;
	wire _w3362_ ;
	wire _w3363_ ;
	wire _w3364_ ;
	wire _w3365_ ;
	wire _w3366_ ;
	wire _w3367_ ;
	wire _w3368_ ;
	wire _w3369_ ;
	wire _w3370_ ;
	wire _w3371_ ;
	wire _w3372_ ;
	wire _w3373_ ;
	wire _w3374_ ;
	wire _w3375_ ;
	wire _w3376_ ;
	wire _w3377_ ;
	wire _w3378_ ;
	wire _w3379_ ;
	wire _w3380_ ;
	wire _w3381_ ;
	wire _w3382_ ;
	wire _w3383_ ;
	wire _w3384_ ;
	wire _w3385_ ;
	wire _w3386_ ;
	wire _w3387_ ;
	wire _w3388_ ;
	wire _w3389_ ;
	wire _w3390_ ;
	wire _w3391_ ;
	wire _w3392_ ;
	wire _w3393_ ;
	wire _w3394_ ;
	wire _w3395_ ;
	wire _w3396_ ;
	wire _w3397_ ;
	wire _w3398_ ;
	wire _w3399_ ;
	wire _w3400_ ;
	wire _w3401_ ;
	wire _w3402_ ;
	wire _w3403_ ;
	wire _w3404_ ;
	wire _w3405_ ;
	wire _w3406_ ;
	wire _w3407_ ;
	wire _w3408_ ;
	wire _w3409_ ;
	wire _w3410_ ;
	wire _w3411_ ;
	wire _w3412_ ;
	wire _w3413_ ;
	wire _w3414_ ;
	wire _w3415_ ;
	wire _w3416_ ;
	wire _w3417_ ;
	wire _w3418_ ;
	wire _w3419_ ;
	wire _w3420_ ;
	wire _w3421_ ;
	wire _w3422_ ;
	wire _w3423_ ;
	wire _w3424_ ;
	wire _w3425_ ;
	wire _w3426_ ;
	wire _w3427_ ;
	wire _w3428_ ;
	wire _w3429_ ;
	wire _w3430_ ;
	wire _w3431_ ;
	wire _w3432_ ;
	wire _w3433_ ;
	wire _w3434_ ;
	wire _w3435_ ;
	wire _w3436_ ;
	wire _w3437_ ;
	wire _w3438_ ;
	wire _w3439_ ;
	wire _w3440_ ;
	wire _w3441_ ;
	wire _w3442_ ;
	wire _w3443_ ;
	wire _w3444_ ;
	wire _w3445_ ;
	wire _w3446_ ;
	wire _w3447_ ;
	wire _w3448_ ;
	wire _w3449_ ;
	wire _w3450_ ;
	wire _w3451_ ;
	wire _w3452_ ;
	wire _w3453_ ;
	wire _w3454_ ;
	wire _w3455_ ;
	wire _w3456_ ;
	wire _w3457_ ;
	wire _w3458_ ;
	wire _w3459_ ;
	wire _w3460_ ;
	wire _w3461_ ;
	wire _w3462_ ;
	wire _w3463_ ;
	wire _w3464_ ;
	wire _w3465_ ;
	wire _w3466_ ;
	wire _w3467_ ;
	wire _w3468_ ;
	wire _w3469_ ;
	wire _w3470_ ;
	wire _w3471_ ;
	wire _w3472_ ;
	wire _w3473_ ;
	wire _w3474_ ;
	wire _w3475_ ;
	wire _w3476_ ;
	wire _w3477_ ;
	wire _w3478_ ;
	wire _w3479_ ;
	wire _w3480_ ;
	wire _w3481_ ;
	wire _w3482_ ;
	wire _w3483_ ;
	wire _w3484_ ;
	wire _w3485_ ;
	wire _w3486_ ;
	wire _w3487_ ;
	wire _w3488_ ;
	wire _w3489_ ;
	wire _w3490_ ;
	wire _w3491_ ;
	wire _w3492_ ;
	wire _w3493_ ;
	wire _w3494_ ;
	wire _w3495_ ;
	wire _w3496_ ;
	wire _w3497_ ;
	wire _w3498_ ;
	wire _w3499_ ;
	wire _w3500_ ;
	wire _w3501_ ;
	wire _w3502_ ;
	wire _w3503_ ;
	wire _w3504_ ;
	wire _w3505_ ;
	wire _w3506_ ;
	wire _w3507_ ;
	wire _w3508_ ;
	wire _w3509_ ;
	wire _w3510_ ;
	wire _w3511_ ;
	wire _w3512_ ;
	wire _w3513_ ;
	wire _w3514_ ;
	wire _w3515_ ;
	wire _w3516_ ;
	wire _w3517_ ;
	wire _w3518_ ;
	wire _w3519_ ;
	wire _w3520_ ;
	wire _w3521_ ;
	wire _w3522_ ;
	wire _w3523_ ;
	wire _w3524_ ;
	wire _w3525_ ;
	wire _w3526_ ;
	wire _w3527_ ;
	wire _w3528_ ;
	wire _w3529_ ;
	wire _w3530_ ;
	wire _w3531_ ;
	wire _w3532_ ;
	wire _w3533_ ;
	wire _w3534_ ;
	wire _w3535_ ;
	wire _w3536_ ;
	wire _w3537_ ;
	wire _w3538_ ;
	wire _w3539_ ;
	wire _w3540_ ;
	wire _w3541_ ;
	wire _w3542_ ;
	wire _w3543_ ;
	wire _w3544_ ;
	wire _w3545_ ;
	wire _w3546_ ;
	wire _w3547_ ;
	wire _w3548_ ;
	wire _w3549_ ;
	wire _w3550_ ;
	wire _w3551_ ;
	wire _w3552_ ;
	wire _w3553_ ;
	wire _w3554_ ;
	wire _w3555_ ;
	wire _w3556_ ;
	wire _w3557_ ;
	wire _w3558_ ;
	wire _w3559_ ;
	wire _w3560_ ;
	wire _w3561_ ;
	wire _w3562_ ;
	wire _w3563_ ;
	wire _w3564_ ;
	wire _w3565_ ;
	wire _w3566_ ;
	wire _w3567_ ;
	wire _w3568_ ;
	wire _w3569_ ;
	wire _w3570_ ;
	wire _w3571_ ;
	wire _w3572_ ;
	wire _w3573_ ;
	wire _w3574_ ;
	wire _w3575_ ;
	wire _w3576_ ;
	wire _w3577_ ;
	wire _w3578_ ;
	wire _w3579_ ;
	wire _w3580_ ;
	wire _w3581_ ;
	wire _w3582_ ;
	wire _w3583_ ;
	wire _w3584_ ;
	wire _w3585_ ;
	wire _w3586_ ;
	wire _w3587_ ;
	wire _w3588_ ;
	wire _w3589_ ;
	wire _w3590_ ;
	wire _w3591_ ;
	wire _w3592_ ;
	wire _w3593_ ;
	wire _w3594_ ;
	wire _w3595_ ;
	wire _w3596_ ;
	wire _w3597_ ;
	wire _w3598_ ;
	wire _w3599_ ;
	wire _w3600_ ;
	wire _w3601_ ;
	wire _w3602_ ;
	wire _w3603_ ;
	wire _w3604_ ;
	wire _w3605_ ;
	wire _w3606_ ;
	wire _w3607_ ;
	wire _w3608_ ;
	wire _w3609_ ;
	wire _w3610_ ;
	wire _w3611_ ;
	wire _w3612_ ;
	wire _w3613_ ;
	wire _w3614_ ;
	wire _w3615_ ;
	wire _w3616_ ;
	wire _w3617_ ;
	wire _w3618_ ;
	wire _w3619_ ;
	wire _w3620_ ;
	wire _w3621_ ;
	wire _w3622_ ;
	wire _w3623_ ;
	wire _w3624_ ;
	wire _w3625_ ;
	wire _w3626_ ;
	wire _w3627_ ;
	wire _w3628_ ;
	wire _w3629_ ;
	wire _w3630_ ;
	wire _w3631_ ;
	wire _w3632_ ;
	wire _w3633_ ;
	wire _w3634_ ;
	wire _w3635_ ;
	wire _w3636_ ;
	wire _w3637_ ;
	wire _w3638_ ;
	wire _w3639_ ;
	wire _w3640_ ;
	wire _w3641_ ;
	wire _w3642_ ;
	wire _w3643_ ;
	wire _w3644_ ;
	wire _w3645_ ;
	wire _w3646_ ;
	wire _w3647_ ;
	wire _w3648_ ;
	wire _w3649_ ;
	wire _w3650_ ;
	wire _w3651_ ;
	wire _w3652_ ;
	wire _w3653_ ;
	wire _w3654_ ;
	wire _w3655_ ;
	wire _w3656_ ;
	wire _w3657_ ;
	wire _w3658_ ;
	wire _w3659_ ;
	wire _w3660_ ;
	wire _w3661_ ;
	wire _w3662_ ;
	wire _w3663_ ;
	wire _w3664_ ;
	wire _w3665_ ;
	wire _w3666_ ;
	wire _w3667_ ;
	wire _w3668_ ;
	wire _w3669_ ;
	wire _w3670_ ;
	wire _w3671_ ;
	wire _w3672_ ;
	wire _w3673_ ;
	wire _w3674_ ;
	wire _w3675_ ;
	wire _w3676_ ;
	wire _w3677_ ;
	wire _w3678_ ;
	wire _w3679_ ;
	wire _w3680_ ;
	wire _w3681_ ;
	wire _w3682_ ;
	wire _w3683_ ;
	wire _w3684_ ;
	wire _w3685_ ;
	wire _w3686_ ;
	wire _w3687_ ;
	wire _w3688_ ;
	wire _w3689_ ;
	wire _w3690_ ;
	wire _w3691_ ;
	wire _w3692_ ;
	wire _w3693_ ;
	wire _w3694_ ;
	wire _w3695_ ;
	wire _w3696_ ;
	wire _w3697_ ;
	wire _w3698_ ;
	wire _w3699_ ;
	wire _w3700_ ;
	wire _w3701_ ;
	wire _w3702_ ;
	wire _w3703_ ;
	wire _w3704_ ;
	wire _w3705_ ;
	wire _w3706_ ;
	wire _w3707_ ;
	wire _w3708_ ;
	wire _w3709_ ;
	wire _w3710_ ;
	wire _w3711_ ;
	wire _w3712_ ;
	wire _w3713_ ;
	wire _w3714_ ;
	wire _w3715_ ;
	wire _w3716_ ;
	wire _w3717_ ;
	wire _w3718_ ;
	wire _w3719_ ;
	wire _w3720_ ;
	wire _w3721_ ;
	wire _w3722_ ;
	wire _w3723_ ;
	wire _w3724_ ;
	wire _w3725_ ;
	wire _w3726_ ;
	wire _w3727_ ;
	wire _w3728_ ;
	wire _w3729_ ;
	wire _w3730_ ;
	wire _w3731_ ;
	wire _w3732_ ;
	wire _w3733_ ;
	wire _w3734_ ;
	wire _w3735_ ;
	wire _w3736_ ;
	wire _w3737_ ;
	wire _w3738_ ;
	wire _w3739_ ;
	wire _w3740_ ;
	wire _w3741_ ;
	wire _w3742_ ;
	wire _w3743_ ;
	wire _w3744_ ;
	wire _w3745_ ;
	wire _w3746_ ;
	wire _w3747_ ;
	wire _w3748_ ;
	wire _w3749_ ;
	wire _w3750_ ;
	wire _w3751_ ;
	wire _w3752_ ;
	wire _w3753_ ;
	wire _w3754_ ;
	wire _w3755_ ;
	wire _w3756_ ;
	wire _w3757_ ;
	wire _w3758_ ;
	wire _w3759_ ;
	wire _w3760_ ;
	wire _w3761_ ;
	wire _w3762_ ;
	wire _w3763_ ;
	wire _w3764_ ;
	wire _w3765_ ;
	wire _w3766_ ;
	wire _w3767_ ;
	wire _w3768_ ;
	wire _w3769_ ;
	wire _w3770_ ;
	wire _w3771_ ;
	wire _w3772_ ;
	wire _w3773_ ;
	wire _w3774_ ;
	wire _w3775_ ;
	wire _w3776_ ;
	wire _w3777_ ;
	wire _w3778_ ;
	wire _w3779_ ;
	wire _w3780_ ;
	wire _w3781_ ;
	wire _w3782_ ;
	wire _w3783_ ;
	wire _w3784_ ;
	wire _w3785_ ;
	wire _w3786_ ;
	wire _w3787_ ;
	wire _w3788_ ;
	wire _w3789_ ;
	wire _w3790_ ;
	wire _w3791_ ;
	wire _w3792_ ;
	wire _w3793_ ;
	wire _w3794_ ;
	wire _w3795_ ;
	wire _w3796_ ;
	wire _w3797_ ;
	wire _w3798_ ;
	wire _w3799_ ;
	wire _w3800_ ;
	wire _w3801_ ;
	wire _w3802_ ;
	wire _w3803_ ;
	wire _w3804_ ;
	wire _w3805_ ;
	wire _w3806_ ;
	wire _w3807_ ;
	wire _w3808_ ;
	wire _w3809_ ;
	wire _w3810_ ;
	wire _w3811_ ;
	wire _w3812_ ;
	wire _w3813_ ;
	wire _w3814_ ;
	wire _w3815_ ;
	wire _w3816_ ;
	wire _w3817_ ;
	wire _w3818_ ;
	wire _w3819_ ;
	wire _w3820_ ;
	wire _w3821_ ;
	wire _w3822_ ;
	wire _w3823_ ;
	wire _w3824_ ;
	wire _w3825_ ;
	wire _w3826_ ;
	wire _w3827_ ;
	wire _w3828_ ;
	wire _w3829_ ;
	wire _w3830_ ;
	wire _w3831_ ;
	wire _w3832_ ;
	wire _w3833_ ;
	wire _w3834_ ;
	wire _w3835_ ;
	wire _w3836_ ;
	wire _w3837_ ;
	wire _w3838_ ;
	wire _w3839_ ;
	wire _w3840_ ;
	wire _w3841_ ;
	wire _w3842_ ;
	wire _w3843_ ;
	wire _w3844_ ;
	wire _w3845_ ;
	wire _w3846_ ;
	wire _w3847_ ;
	wire _w3848_ ;
	wire _w3849_ ;
	wire _w3850_ ;
	wire _w3851_ ;
	wire _w3852_ ;
	wire _w3853_ ;
	wire _w3854_ ;
	wire _w3855_ ;
	wire _w3856_ ;
	wire _w3857_ ;
	wire _w3858_ ;
	wire _w3859_ ;
	wire _w3860_ ;
	wire _w3861_ ;
	wire _w3862_ ;
	wire _w3863_ ;
	wire _w3864_ ;
	wire _w3865_ ;
	wire _w3866_ ;
	wire _w3867_ ;
	wire _w3868_ ;
	wire _w3869_ ;
	wire _w3870_ ;
	wire _w3871_ ;
	wire _w3872_ ;
	wire _w3873_ ;
	wire _w3874_ ;
	wire _w3875_ ;
	wire _w3876_ ;
	wire _w3877_ ;
	wire _w3878_ ;
	wire _w3879_ ;
	wire _w3880_ ;
	wire _w3881_ ;
	wire _w3882_ ;
	wire _w3883_ ;
	wire _w3884_ ;
	wire _w3885_ ;
	wire _w3886_ ;
	wire _w3887_ ;
	wire _w3888_ ;
	wire _w3889_ ;
	wire _w3890_ ;
	wire _w3891_ ;
	wire _w3892_ ;
	wire _w3893_ ;
	wire _w3894_ ;
	wire _w3895_ ;
	wire _w3896_ ;
	wire _w3897_ ;
	wire _w3898_ ;
	wire _w3899_ ;
	wire _w3900_ ;
	wire _w3901_ ;
	wire _w3902_ ;
	wire _w3903_ ;
	wire _w3904_ ;
	wire _w3905_ ;
	wire _w3906_ ;
	wire _w3907_ ;
	wire _w3908_ ;
	wire _w3909_ ;
	wire _w3910_ ;
	wire _w3911_ ;
	wire _w3912_ ;
	wire _w3913_ ;
	wire _w3914_ ;
	wire _w3915_ ;
	wire _w3916_ ;
	wire _w3917_ ;
	wire _w3918_ ;
	wire _w3919_ ;
	wire _w3920_ ;
	wire _w3921_ ;
	wire _w3922_ ;
	wire _w3923_ ;
	wire _w3924_ ;
	wire _w3925_ ;
	wire _w3926_ ;
	wire _w3927_ ;
	wire _w3928_ ;
	wire _w3929_ ;
	wire _w3930_ ;
	wire _w3931_ ;
	wire _w3932_ ;
	wire _w3933_ ;
	wire _w3934_ ;
	wire _w3935_ ;
	wire _w3936_ ;
	wire _w3937_ ;
	wire _w3938_ ;
	wire _w3939_ ;
	wire _w3940_ ;
	wire _w3941_ ;
	wire _w3942_ ;
	wire _w3943_ ;
	wire _w3944_ ;
	wire _w3945_ ;
	wire _w3946_ ;
	wire _w3947_ ;
	wire _w3948_ ;
	wire _w3949_ ;
	wire _w3950_ ;
	wire _w3951_ ;
	wire _w3952_ ;
	wire _w3953_ ;
	wire _w3954_ ;
	wire _w3955_ ;
	wire _w3956_ ;
	wire _w3957_ ;
	wire _w3958_ ;
	wire _w3959_ ;
	wire _w3960_ ;
	wire _w3961_ ;
	wire _w3962_ ;
	wire _w3963_ ;
	wire _w3964_ ;
	wire _w3965_ ;
	wire _w3966_ ;
	wire _w3967_ ;
	wire _w3968_ ;
	wire _w3969_ ;
	wire _w3970_ ;
	wire _w3971_ ;
	wire _w3972_ ;
	wire _w3973_ ;
	wire _w3974_ ;
	wire _w3975_ ;
	wire _w3976_ ;
	wire _w3977_ ;
	wire _w3978_ ;
	wire _w3979_ ;
	wire _w3980_ ;
	wire _w3981_ ;
	wire _w3982_ ;
	wire _w3983_ ;
	wire _w3984_ ;
	wire _w3985_ ;
	wire _w3986_ ;
	wire _w3987_ ;
	wire _w3988_ ;
	wire _w3989_ ;
	wire _w3990_ ;
	wire _w3991_ ;
	wire _w3992_ ;
	wire _w3993_ ;
	wire _w3994_ ;
	wire _w3995_ ;
	wire _w3996_ ;
	wire _w3997_ ;
	wire _w3998_ ;
	wire _w3999_ ;
	wire _w4000_ ;
	wire _w4001_ ;
	wire _w4002_ ;
	wire _w4003_ ;
	wire _w4004_ ;
	wire _w4005_ ;
	wire _w4006_ ;
	wire _w4007_ ;
	wire _w4008_ ;
	wire _w4009_ ;
	wire _w4010_ ;
	wire _w4011_ ;
	wire _w4012_ ;
	wire _w4013_ ;
	wire _w4014_ ;
	wire _w4015_ ;
	wire _w4016_ ;
	wire _w4017_ ;
	wire _w4018_ ;
	wire _w4019_ ;
	wire _w4020_ ;
	wire _w4021_ ;
	wire _w4022_ ;
	wire _w4023_ ;
	wire _w4024_ ;
	wire _w4025_ ;
	wire _w4026_ ;
	wire _w4027_ ;
	wire _w4028_ ;
	wire _w4029_ ;
	wire _w4030_ ;
	wire _w4031_ ;
	wire _w4032_ ;
	wire _w4033_ ;
	wire _w4034_ ;
	wire _w4035_ ;
	wire _w4036_ ;
	wire _w4037_ ;
	wire _w4038_ ;
	wire _w4039_ ;
	wire _w4040_ ;
	wire _w4041_ ;
	wire _w4042_ ;
	wire _w4043_ ;
	wire _w4044_ ;
	wire _w4045_ ;
	wire _w4046_ ;
	wire _w4047_ ;
	wire _w4048_ ;
	wire _w4049_ ;
	wire _w4050_ ;
	wire _w4051_ ;
	wire _w4052_ ;
	wire _w4053_ ;
	wire _w4054_ ;
	wire _w4055_ ;
	wire _w4056_ ;
	wire _w4057_ ;
	wire _w4058_ ;
	wire _w4059_ ;
	wire _w4060_ ;
	wire _w4061_ ;
	wire _w4062_ ;
	wire _w4063_ ;
	wire _w4064_ ;
	wire _w4065_ ;
	wire _w4066_ ;
	wire _w4067_ ;
	wire _w4068_ ;
	wire _w4069_ ;
	wire _w4070_ ;
	wire _w4071_ ;
	wire _w4072_ ;
	wire _w4073_ ;
	wire _w4074_ ;
	wire _w4075_ ;
	wire _w4076_ ;
	wire _w4077_ ;
	wire _w4078_ ;
	wire _w4079_ ;
	wire _w4080_ ;
	wire _w4081_ ;
	wire _w4082_ ;
	wire _w4083_ ;
	wire _w4084_ ;
	wire _w4085_ ;
	wire _w4086_ ;
	wire _w4087_ ;
	wire _w4088_ ;
	wire _w4089_ ;
	wire _w4090_ ;
	wire _w4091_ ;
	wire _w4092_ ;
	wire _w4093_ ;
	wire _w4094_ ;
	wire _w4095_ ;
	wire _w4096_ ;
	wire _w4097_ ;
	wire _w4098_ ;
	wire _w4099_ ;
	wire _w4100_ ;
	wire _w4101_ ;
	wire _w4102_ ;
	wire _w4103_ ;
	wire _w4104_ ;
	wire _w4105_ ;
	wire _w4106_ ;
	wire _w4107_ ;
	wire _w4108_ ;
	wire _w4109_ ;
	wire _w4110_ ;
	wire _w4111_ ;
	wire _w4112_ ;
	wire _w4113_ ;
	wire _w4114_ ;
	wire _w4115_ ;
	wire _w4116_ ;
	wire _w4117_ ;
	wire _w4118_ ;
	wire _w4119_ ;
	wire _w4120_ ;
	wire _w4121_ ;
	wire _w4122_ ;
	wire _w4123_ ;
	wire _w4124_ ;
	wire _w4125_ ;
	wire _w4126_ ;
	wire _w4127_ ;
	wire _w4128_ ;
	wire _w4129_ ;
	wire _w4130_ ;
	wire _w4131_ ;
	wire _w4132_ ;
	wire _w4133_ ;
	wire _w4134_ ;
	wire _w4135_ ;
	wire _w4136_ ;
	wire _w4137_ ;
	wire _w4138_ ;
	wire _w4139_ ;
	wire _w4140_ ;
	wire _w4141_ ;
	wire _w4142_ ;
	wire _w4143_ ;
	wire _w4144_ ;
	wire _w4145_ ;
	wire _w4146_ ;
	wire _w4147_ ;
	wire _w4148_ ;
	wire _w4149_ ;
	wire _w4150_ ;
	wire _w4151_ ;
	wire _w4152_ ;
	wire _w4153_ ;
	wire _w4154_ ;
	wire _w4155_ ;
	wire _w4156_ ;
	wire _w4157_ ;
	wire _w4158_ ;
	wire _w4159_ ;
	wire _w4160_ ;
	wire _w4161_ ;
	wire _w4162_ ;
	wire _w4163_ ;
	wire _w4164_ ;
	wire _w4165_ ;
	wire _w4166_ ;
	wire _w4167_ ;
	wire _w4168_ ;
	wire _w4169_ ;
	wire _w4170_ ;
	wire _w4171_ ;
	wire _w4172_ ;
	wire _w4173_ ;
	wire _w4174_ ;
	wire _w4175_ ;
	wire _w4176_ ;
	wire _w4177_ ;
	wire _w4178_ ;
	wire _w4179_ ;
	wire _w4180_ ;
	wire _w4181_ ;
	wire _w4182_ ;
	wire _w4183_ ;
	wire _w4184_ ;
	wire _w4185_ ;
	wire _w4186_ ;
	wire _w4187_ ;
	wire _w4188_ ;
	wire _w4189_ ;
	wire _w4190_ ;
	wire _w4191_ ;
	wire _w4192_ ;
	wire _w4193_ ;
	wire _w4194_ ;
	wire _w4195_ ;
	wire _w4196_ ;
	wire _w4197_ ;
	wire _w4198_ ;
	wire _w4199_ ;
	wire _w4200_ ;
	wire _w4201_ ;
	wire _w4202_ ;
	wire _w4203_ ;
	wire _w4204_ ;
	wire _w4205_ ;
	wire _w4206_ ;
	wire _w4207_ ;
	wire _w4208_ ;
	wire _w4209_ ;
	wire _w4210_ ;
	wire _w4211_ ;
	wire _w4212_ ;
	wire _w4213_ ;
	wire _w4214_ ;
	wire _w4215_ ;
	wire _w4216_ ;
	wire _w4217_ ;
	wire _w4218_ ;
	wire _w4219_ ;
	wire _w4220_ ;
	wire _w4221_ ;
	wire _w4222_ ;
	wire _w4223_ ;
	wire _w4224_ ;
	wire _w4225_ ;
	wire _w4226_ ;
	wire _w4227_ ;
	wire _w4228_ ;
	wire _w4229_ ;
	wire _w4230_ ;
	wire _w4231_ ;
	wire _w4232_ ;
	wire _w4233_ ;
	wire _w4234_ ;
	wire _w4235_ ;
	wire _w4236_ ;
	wire _w4237_ ;
	wire _w4238_ ;
	wire _w4239_ ;
	wire _w4240_ ;
	wire _w4241_ ;
	wire _w4242_ ;
	wire _w4243_ ;
	wire _w4244_ ;
	wire _w4245_ ;
	wire _w4246_ ;
	wire _w4247_ ;
	wire _w4248_ ;
	wire _w4249_ ;
	wire _w4250_ ;
	wire _w4251_ ;
	wire _w4252_ ;
	wire _w4253_ ;
	wire _w4254_ ;
	wire _w4255_ ;
	wire _w4256_ ;
	wire _w4257_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4304_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4335_ ;
	wire _w4336_ ;
	wire _w4337_ ;
	wire _w4338_ ;
	wire _w4339_ ;
	wire _w4340_ ;
	wire _w4341_ ;
	wire _w4342_ ;
	wire _w4343_ ;
	wire _w4344_ ;
	wire _w4345_ ;
	wire _w4346_ ;
	wire _w4347_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4363_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4383_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4433_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4574_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w5156_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5166_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5190_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5262_ ;
	wire _w5263_ ;
	wire _w5264_ ;
	wire _w5265_ ;
	wire _w5266_ ;
	wire _w5267_ ;
	wire _w5268_ ;
	wire _w5269_ ;
	wire _w5270_ ;
	wire _w5271_ ;
	wire _w5272_ ;
	wire _w5273_ ;
	wire _w5274_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5290_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	wire _w5301_ ;
	wire _w5302_ ;
	wire _w5304_ ;
	wire _w5305_ ;
	wire _w5306_ ;
	wire _w5307_ ;
	wire _w5308_ ;
	wire _w5309_ ;
	wire _w5310_ ;
	wire _w5311_ ;
	wire _w5312_ ;
	wire _w5313_ ;
	wire _w5314_ ;
	wire _w5315_ ;
	wire _w5316_ ;
	wire _w5317_ ;
	wire _w5318_ ;
	wire _w5319_ ;
	wire _w5320_ ;
	wire _w5321_ ;
	wire _w5322_ ;
	wire _w5323_ ;
	wire _w5324_ ;
	wire _w5325_ ;
	wire _w5326_ ;
	wire _w5327_ ;
	wire _w5328_ ;
	wire _w5329_ ;
	wire _w5330_ ;
	wire _w5331_ ;
	wire _w5332_ ;
	wire _w5333_ ;
	wire _w5334_ ;
	wire _w5335_ ;
	wire _w5336_ ;
	wire _w5337_ ;
	wire _w5338_ ;
	wire _w5339_ ;
	wire _w5340_ ;
	wire _w5341_ ;
	wire _w5342_ ;
	wire _w5343_ ;
	wire _w5344_ ;
	wire _w5345_ ;
	wire _w5346_ ;
	wire _w5347_ ;
	wire _w5348_ ;
	wire _w5349_ ;
	wire _w5350_ ;
	wire _w5351_ ;
	wire _w5352_ ;
	wire _w5353_ ;
	wire _w5354_ ;
	wire _w5355_ ;
	wire _w5356_ ;
	wire _w5357_ ;
	wire _w5358_ ;
	wire _w5359_ ;
	wire _w5360_ ;
	wire _w5361_ ;
	wire _w5362_ ;
	wire _w5363_ ;
	wire _w5364_ ;
	wire _w5365_ ;
	wire _w5366_ ;
	wire _w5367_ ;
	wire _w5368_ ;
	wire _w5369_ ;
	wire _w5370_ ;
	wire _w5371_ ;
	wire _w5372_ ;
	wire _w5373_ ;
	wire _w5374_ ;
	wire _w5375_ ;
	wire _w5376_ ;
	wire _w5377_ ;
	wire _w5378_ ;
	wire _w5379_ ;
	wire _w5380_ ;
	wire _w5381_ ;
	wire _w5382_ ;
	wire _w5383_ ;
	wire _w5384_ ;
	wire _w5385_ ;
	wire _w5386_ ;
	wire _w5387_ ;
	wire _w5388_ ;
	wire _w5389_ ;
	wire _w5390_ ;
	wire _w5391_ ;
	wire _w5392_ ;
	wire _w5393_ ;
	wire _w5394_ ;
	wire _w5395_ ;
	wire _w5396_ ;
	wire _w5397_ ;
	wire _w5398_ ;
	wire _w5399_ ;
	wire _w5400_ ;
	wire _w5401_ ;
	wire _w5402_ ;
	wire _w5403_ ;
	wire _w5404_ ;
	wire _w5405_ ;
	wire _w5406_ ;
	wire _w5407_ ;
	wire _w5408_ ;
	wire _w5409_ ;
	wire _w5410_ ;
	wire _w5411_ ;
	wire _w5412_ ;
	wire _w5413_ ;
	wire _w5414_ ;
	wire _w5415_ ;
	wire _w5416_ ;
	wire _w5417_ ;
	wire _w5418_ ;
	wire _w5419_ ;
	wire _w5420_ ;
	wire _w5421_ ;
	wire _w5422_ ;
	wire _w5423_ ;
	wire _w5424_ ;
	wire _w5425_ ;
	wire _w5426_ ;
	wire _w5427_ ;
	wire _w5428_ ;
	wire _w5429_ ;
	wire _w5430_ ;
	wire _w5431_ ;
	wire _w5432_ ;
	wire _w5433_ ;
	wire _w5434_ ;
	wire _w5435_ ;
	wire _w5436_ ;
	wire _w5437_ ;
	wire _w5438_ ;
	wire _w5439_ ;
	wire _w5440_ ;
	wire _w5441_ ;
	wire _w5442_ ;
	wire _w5443_ ;
	wire _w5444_ ;
	wire _w5445_ ;
	wire _w5446_ ;
	wire _w5447_ ;
	wire _w5448_ ;
	wire _w5449_ ;
	wire _w5450_ ;
	wire _w5451_ ;
	wire _w5452_ ;
	wire _w5453_ ;
	wire _w5454_ ;
	wire _w5455_ ;
	wire _w5456_ ;
	wire _w5457_ ;
	wire _w5458_ ;
	wire _w5459_ ;
	wire _w5460_ ;
	wire _w5461_ ;
	wire _w5462_ ;
	wire _w5463_ ;
	wire _w5464_ ;
	wire _w5465_ ;
	wire _w5466_ ;
	wire _w5467_ ;
	wire _w5468_ ;
	wire _w5469_ ;
	wire _w5470_ ;
	wire _w5471_ ;
	wire _w5472_ ;
	wire _w5473_ ;
	wire _w5474_ ;
	wire _w5475_ ;
	wire _w5476_ ;
	wire _w5477_ ;
	wire _w5478_ ;
	wire _w5479_ ;
	wire _w5480_ ;
	wire _w5481_ ;
	wire _w5482_ ;
	wire _w5483_ ;
	wire _w5484_ ;
	wire _w5485_ ;
	wire _w5486_ ;
	wire _w5487_ ;
	wire _w5488_ ;
	wire _w5489_ ;
	wire _w5490_ ;
	wire _w5491_ ;
	wire _w5492_ ;
	wire _w5493_ ;
	wire _w5494_ ;
	wire _w5495_ ;
	wire _w5496_ ;
	wire _w5497_ ;
	wire _w5498_ ;
	wire _w5499_ ;
	wire _w5500_ ;
	wire _w5501_ ;
	wire _w5502_ ;
	wire _w5503_ ;
	wire _w5504_ ;
	wire _w5505_ ;
	wire _w5506_ ;
	wire _w5507_ ;
	wire _w5508_ ;
	wire _w5509_ ;
	wire _w5510_ ;
	wire _w5511_ ;
	wire _w5512_ ;
	wire _w5513_ ;
	wire _w5514_ ;
	wire _w5515_ ;
	wire _w5516_ ;
	wire _w5517_ ;
	wire _w5518_ ;
	wire _w5519_ ;
	wire _w5520_ ;
	wire _w5521_ ;
	wire _w5522_ ;
	wire _w5523_ ;
	wire _w5524_ ;
	wire _w5525_ ;
	wire _w5526_ ;
	wire _w5527_ ;
	wire _w5528_ ;
	wire _w5529_ ;
	wire _w5530_ ;
	wire _w5531_ ;
	wire _w5532_ ;
	wire _w5533_ ;
	wire _w5534_ ;
	wire _w5535_ ;
	wire _w5536_ ;
	wire _w5537_ ;
	wire _w5538_ ;
	wire _w5539_ ;
	wire _w5540_ ;
	wire _w5541_ ;
	wire _w5542_ ;
	wire _w5543_ ;
	wire _w5544_ ;
	wire _w5545_ ;
	wire _w5546_ ;
	wire _w5547_ ;
	wire _w5548_ ;
	wire _w5549_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\P1_state_reg[0]/NET0131 ,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		_w464_
	);
	LUT3 #(
		.INIT('h01)
	) name2 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[8]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		_w465_
	);
	LUT4 #(
		.INIT('h0001)
	) name3 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[2]/NET0131 ,
		\P1_IR_reg[3]/NET0131 ,
		_w466_
	);
	LUT3 #(
		.INIT('h01)
	) name4 (
		\P1_IR_reg[5]/NET0131 ,
		\P1_IR_reg[6]/NET0131 ,
		\P1_IR_reg[7]/NET0131 ,
		_w467_
	);
	LUT3 #(
		.INIT('h40)
	) name5 (
		\P1_IR_reg[4]/NET0131 ,
		_w466_,
		_w467_,
		_w468_
	);
	LUT4 #(
		.INIT('h4000)
	) name6 (
		\P1_IR_reg[4]/NET0131 ,
		_w465_,
		_w466_,
		_w467_,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[12]/NET0131 ,
		_w470_
	);
	LUT3 #(
		.INIT('h01)
	) name8 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[12]/NET0131 ,
		\P1_IR_reg[13]/NET0131 ,
		_w471_
	);
	LUT4 #(
		.INIT('h0001)
	) name9 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[12]/NET0131 ,
		\P1_IR_reg[13]/NET0131 ,
		\P1_IR_reg[14]/NET0131 ,
		_w472_
	);
	LUT4 #(
		.INIT('h0001)
	) name10 (
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[17]/NET0131 ,
		\P1_IR_reg[18]/NET0131 ,
		_w473_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w472_,
		_w473_,
		_w474_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		_w475_
	);
	LUT4 #(
		.INIT('h0001)
	) name13 (
		\P1_IR_reg[19]/NET0131 ,
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		\P1_IR_reg[22]/NET0131 ,
		_w476_
	);
	LUT4 #(
		.INIT('h0001)
	) name14 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		\P1_IR_reg[25]/NET0131 ,
		\P1_IR_reg[26]/NET0131 ,
		_w477_
	);
	LUT4 #(
		.INIT('h8000)
	) name15 (
		_w469_,
		_w474_,
		_w476_,
		_w477_,
		_w478_
	);
	LUT3 #(
		.INIT('h59)
	) name16 (
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[15]/NET0131 ,
		_w480_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		_w465_,
		_w471_,
		_w481_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name19 (
		\P1_IR_reg[31]/NET0131 ,
		_w468_,
		_w480_,
		_w481_,
		_w482_
	);
	LUT4 #(
		.INIT('h0001)
	) name20 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[17]/NET0131 ,
		\P1_IR_reg[18]/NET0131 ,
		\P1_IR_reg[19]/NET0131 ,
		_w483_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\P1_IR_reg[22]/NET0131 ,
		\P1_IR_reg[23]/NET0131 ,
		_w484_
	);
	LUT4 #(
		.INIT('h0001)
	) name22 (
		\P1_IR_reg[24]/NET0131 ,
		\P1_IR_reg[25]/NET0131 ,
		\P1_IR_reg[26]/NET0131 ,
		\P1_IR_reg[27]/NET0131 ,
		_w485_
	);
	LUT4 #(
		.INIT('h8000)
	) name23 (
		_w483_,
		_w475_,
		_w484_,
		_w485_,
		_w486_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\P1_IR_reg[31]/NET0131 ,
		_w486_,
		_w487_
	);
	LUT3 #(
		.INIT('h56)
	) name25 (
		\P1_IR_reg[28]/NET0131 ,
		_w482_,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		_w479_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\P2_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w490_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		\P2_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w491_
	);
	LUT4 #(
		.INIT('hec80)
	) name29 (
		\P2_datao_reg[0]/NET0131 ,
		\P2_datao_reg[1]/NET0131 ,
		\si[0]_pad ,
		\si[1]_pad ,
		_w492_
	);
	LUT3 #(
		.INIT('h17)
	) name30 (
		\P2_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		\P2_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w494_
	);
	LUT4 #(
		.INIT('hfac8)
	) name32 (
		\P2_datao_reg[5]/NET0131 ,
		\P2_datao_reg[6]/NET0131 ,
		\si[5]_pad ,
		\si[6]_pad ,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\P2_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w496_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		\P2_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w497_
	);
	LUT4 #(
		.INIT('hfac8)
	) name35 (
		\P2_datao_reg[3]/NET0131 ,
		\P2_datao_reg[4]/NET0131 ,
		\si[3]_pad ,
		\si[4]_pad ,
		_w498_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w495_,
		_w498_,
		_w499_
	);
	LUT4 #(
		.INIT('hec80)
	) name37 (
		\P2_datao_reg[5]/NET0131 ,
		\P2_datao_reg[6]/NET0131 ,
		\si[5]_pad ,
		\si[6]_pad ,
		_w500_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\P2_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w501_
	);
	LUT4 #(
		.INIT('h135f)
	) name39 (
		\P2_datao_reg[3]/NET0131 ,
		\P2_datao_reg[4]/NET0131 ,
		\si[3]_pad ,
		\si[4]_pad ,
		_w502_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name40 (
		_w495_,
		_w496_,
		_w500_,
		_w502_,
		_w503_
	);
	LUT3 #(
		.INIT('hb0)
	) name41 (
		_w493_,
		_w499_,
		_w503_,
		_w504_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		\P2_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w505_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\P2_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w506_
	);
	LUT4 #(
		.INIT('hfac8)
	) name44 (
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		\si[10]_pad ,
		\si[9]_pad ,
		_w507_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		\P2_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w508_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		\P2_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w509_
	);
	LUT4 #(
		.INIT('hfac8)
	) name47 (
		\P2_datao_reg[7]/NET0131 ,
		\P2_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w510_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		_w507_,
		_w510_,
		_w511_
	);
	LUT4 #(
		.INIT('h4f00)
	) name49 (
		_w493_,
		_w499_,
		_w503_,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		\P2_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w513_
	);
	LUT4 #(
		.INIT('he8a0)
	) name51 (
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		\si[10]_pad ,
		\si[9]_pad ,
		_w514_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		\P2_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w515_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\P2_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w516_
	);
	LUT4 #(
		.INIT('h135f)
	) name54 (
		\P2_datao_reg[7]/NET0131 ,
		\P2_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w517_
	);
	LUT4 #(
		.INIT('h5551)
	) name55 (
		_w514_,
		_w507_,
		_w508_,
		_w517_,
		_w518_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\P2_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w519_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		\P2_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w520_
	);
	LUT4 #(
		.INIT('hfac8)
	) name58 (
		\P2_datao_reg[13]/NET0131 ,
		\P2_datao_reg[14]/NET0131 ,
		\si[13]_pad ,
		\si[14]_pad ,
		_w521_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		\P2_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w522_
	);
	LUT3 #(
		.INIT('h04)
	) name60 (
		_w519_,
		_w521_,
		_w522_,
		_w523_
	);
	LUT4 #(
		.INIT('hec80)
	) name61 (
		\P2_datao_reg[13]/NET0131 ,
		\P2_datao_reg[14]/NET0131 ,
		\si[13]_pad ,
		\si[14]_pad ,
		_w524_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		\P2_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w525_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		\P2_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w526_
	);
	LUT4 #(
		.INIT('h135f)
	) name64 (
		\P2_datao_reg[11]/NET0131 ,
		\P2_datao_reg[12]/NET0131 ,
		\si[11]_pad ,
		\si[12]_pad ,
		_w527_
	);
	LUT4 #(
		.INIT('h5545)
	) name65 (
		_w524_,
		_w519_,
		_w521_,
		_w527_,
		_w528_
	);
	LUT4 #(
		.INIT('h4f00)
	) name66 (
		_w512_,
		_w518_,
		_w523_,
		_w528_,
		_w529_
	);
	LUT4 #(
		.INIT('hfac8)
	) name67 (
		\P2_datao_reg[17]/NET0131 ,
		\P2_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w530_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		\P2_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w531_
	);
	LUT4 #(
		.INIT('hfac8)
	) name69 (
		\P2_datao_reg[15]/NET0131 ,
		\P2_datao_reg[16]/NET0131 ,
		\si[15]_pad ,
		\si[16]_pad ,
		_w532_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		_w530_,
		_w532_,
		_w533_
	);
	LUT4 #(
		.INIT('hfac8)
	) name71 (
		\P2_datao_reg[21]/NET0131 ,
		\P2_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w534_
	);
	LUT4 #(
		.INIT('hfac8)
	) name72 (
		\P2_datao_reg[19]/NET0131 ,
		\P2_datao_reg[20]/NET0131 ,
		\si[19]_pad ,
		\si[20]_pad ,
		_w535_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		_w534_,
		_w535_,
		_w536_
	);
	LUT4 #(
		.INIT('hec80)
	) name74 (
		\P2_datao_reg[21]/NET0131 ,
		\P2_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w537_
	);
	LUT4 #(
		.INIT('hec80)
	) name75 (
		\P2_datao_reg[19]/NET0131 ,
		\P2_datao_reg[20]/NET0131 ,
		\si[19]_pad ,
		\si[20]_pad ,
		_w538_
	);
	LUT3 #(
		.INIT('h13)
	) name76 (
		_w534_,
		_w537_,
		_w538_,
		_w539_
	);
	LUT4 #(
		.INIT('hec80)
	) name77 (
		\P2_datao_reg[17]/NET0131 ,
		\P2_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w540_
	);
	LUT4 #(
		.INIT('hec80)
	) name78 (
		\P2_datao_reg[15]/NET0131 ,
		\P2_datao_reg[16]/NET0131 ,
		\si[15]_pad ,
		\si[16]_pad ,
		_w541_
	);
	LUT3 #(
		.INIT('h13)
	) name79 (
		_w530_,
		_w540_,
		_w541_,
		_w542_
	);
	LUT3 #(
		.INIT('hb0)
	) name80 (
		_w542_,
		_w536_,
		_w539_,
		_w543_
	);
	LUT4 #(
		.INIT('hbf00)
	) name81 (
		_w529_,
		_w533_,
		_w536_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		\P2_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w545_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		\P2_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		\P2_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w547_
	);
	LUT4 #(
		.INIT('hfac8)
	) name85 (
		\P2_datao_reg[24]/NET0131 ,
		\P2_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w548_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		_w546_,
		_w548_,
		_w549_
	);
	LUT3 #(
		.INIT('h10)
	) name87 (
		_w545_,
		_w546_,
		_w548_,
		_w550_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		\P2_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		\P2_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w552_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		\P2_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w553_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		\P2_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w554_
	);
	LUT4 #(
		.INIT('hfac8)
	) name92 (
		\P2_datao_reg[27]/NET0131 ,
		\P2_datao_reg[28]/NET0131 ,
		\si[27]_pad ,
		\si[28]_pad ,
		_w555_
	);
	LUT3 #(
		.INIT('h04)
	) name93 (
		_w552_,
		_w555_,
		_w551_,
		_w556_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		_w550_,
		_w556_,
		_w557_
	);
	LUT4 #(
		.INIT('hec80)
	) name95 (
		\P2_datao_reg[25]/NET0131 ,
		\P2_datao_reg[26]/NET0131 ,
		\si[25]_pad ,
		\si[26]_pad ,
		_w558_
	);
	LUT4 #(
		.INIT('h135f)
	) name96 (
		\P2_datao_reg[23]/NET0131 ,
		\P2_datao_reg[24]/NET0131 ,
		\si[23]_pad ,
		\si[24]_pad ,
		_w559_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name97 (
		_w546_,
		_w548_,
		_w558_,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		\P2_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w561_
	);
	LUT4 #(
		.INIT('h135f)
	) name99 (
		\P2_datao_reg[27]/NET0131 ,
		\P2_datao_reg[28]/NET0131 ,
		\si[27]_pad ,
		\si[28]_pad ,
		_w562_
	);
	LUT4 #(
		.INIT('hfac8)
	) name100 (
		\P2_datao_reg[28]/NET0131 ,
		\P2_datao_reg[29]/NET0131 ,
		\si[28]_pad ,
		\si[29]_pad ,
		_w563_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name101 (
		_w561_,
		_w562_,
		_w551_,
		_w563_,
		_w564_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		\P2_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w565_
	);
	LUT4 #(
		.INIT('h000b)
	) name103 (
		_w560_,
		_w556_,
		_w564_,
		_w565_,
		_w566_
	);
	LUT3 #(
		.INIT('hb0)
	) name104 (
		_w544_,
		_w557_,
		_w566_,
		_w567_
	);
	LUT4 #(
		.INIT('hfe5e)
	) name105 (
		\P1_addr_reg[19]/NET0131 ,
		\P1_rd_reg/NET0131 ,
		\P2_addr_reg[19]/NET0131 ,
		\P2_rd_reg/NET0131 ,
		_w568_
	);
	LUT4 #(
		.INIT('ha6a9)
	) name106 (
		\P2_datao_reg[31]/NET0131 ,
		\si[31]_pad ,
		_w568_,
		_w567_,
		_w569_
	);
	LUT2 #(
		.INIT('h4)
	) name107 (
		_w489_,
		_w569_,
		_w570_
	);
	LUT4 #(
		.INIT('h0001)
	) name108 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		\P1_IR_reg[25]/NET0131 ,
		_w571_
	);
	LUT4 #(
		.INIT('h8000)
	) name109 (
		_w483_,
		_w475_,
		_w484_,
		_w571_,
		_w572_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name110 (
		\P1_IR_reg[31]/NET0131 ,
		_w468_,
		_w481_,
		_w572_,
		_w573_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[28]/NET0131 ,
		_w574_
	);
	LUT4 #(
		.INIT('h0001)
	) name112 (
		\P1_IR_reg[26]/NET0131 ,
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[28]/NET0131 ,
		\P1_IR_reg[29]/NET0131 ,
		_w575_
	);
	LUT2 #(
		.INIT('h2)
	) name113 (
		\P1_IR_reg[31]/NET0131 ,
		_w575_,
		_w576_
	);
	LUT3 #(
		.INIT('h56)
	) name114 (
		\P1_IR_reg[30]/NET0131 ,
		_w573_,
		_w576_,
		_w577_
	);
	LUT4 #(
		.INIT('h0001)
	) name115 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_IR_reg[18]/NET0131 ,
		\P1_IR_reg[19]/NET0131 ,
		\P1_IR_reg[20]/NET0131 ,
		_w578_
	);
	LUT4 #(
		.INIT('h0001)
	) name116 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[16]/NET0131 ,
		_w579_
	);
	LUT4 #(
		.INIT('h0001)
	) name117 (
		\P1_IR_reg[21]/NET0131 ,
		\P1_IR_reg[22]/NET0131 ,
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		_w580_
	);
	LUT4 #(
		.INIT('h0001)
	) name118 (
		\P1_IR_reg[25]/NET0131 ,
		\P1_IR_reg[26]/NET0131 ,
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[28]/NET0131 ,
		_w581_
	);
	LUT4 #(
		.INIT('h8000)
	) name119 (
		_w579_,
		_w578_,
		_w580_,
		_w581_,
		_w582_
	);
	LUT4 #(
		.INIT('hd555)
	) name120 (
		\P1_IR_reg[31]/NET0131 ,
		_w469_,
		_w470_,
		_w582_,
		_w583_
	);
	LUT2 #(
		.INIT('h9)
	) name121 (
		\P1_IR_reg[29]/NET0131 ,
		_w583_,
		_w584_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		_w577_,
		_w584_,
		_w585_
	);
	LUT4 #(
		.INIT('h8000)
	) name123 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		\P1_reg3_reg[5]/NET0131 ,
		\P1_reg3_reg[6]/NET0131 ,
		_w586_
	);
	LUT4 #(
		.INIT('h8000)
	) name124 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_reg3_reg[8]/NET0131 ,
		\P1_reg3_reg[9]/NET0131 ,
		_w586_,
		_w587_
	);
	LUT4 #(
		.INIT('h8000)
	) name125 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_reg3_reg[11]/NET0131 ,
		\P1_reg3_reg[12]/NET0131 ,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		\P1_reg3_reg[13]/NET0131 ,
		\P1_reg3_reg[14]/NET0131 ,
		_w589_
	);
	LUT3 #(
		.INIT('h80)
	) name127 (
		\P1_reg3_reg[15]/NET0131 ,
		\P1_reg3_reg[16]/NET0131 ,
		\P1_reg3_reg[17]/NET0131 ,
		_w590_
	);
	LUT3 #(
		.INIT('h80)
	) name128 (
		_w588_,
		_w589_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\P1_reg3_reg[18]/NET0131 ,
		\P1_reg3_reg[19]/NET0131 ,
		_w592_
	);
	LUT4 #(
		.INIT('h8000)
	) name130 (
		_w588_,
		_w589_,
		_w590_,
		_w592_,
		_w593_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		\P1_reg3_reg[20]/NET0131 ,
		\P1_reg3_reg[21]/NET0131 ,
		_w594_
	);
	LUT3 #(
		.INIT('h80)
	) name132 (
		\P1_reg3_reg[22]/NET0131 ,
		\P1_reg3_reg[23]/NET0131 ,
		\P1_reg3_reg[24]/NET0131 ,
		_w595_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		_w594_,
		_w595_,
		_w596_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		_w593_,
		_w596_,
		_w597_
	);
	LUT4 #(
		.INIT('h8000)
	) name135 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_reg3_reg[26]/NET0131 ,
		\P1_reg3_reg[27]/NET0131 ,
		\P1_reg3_reg[28]/NET0131 ,
		_w598_
	);
	LUT3 #(
		.INIT('h80)
	) name136 (
		_w593_,
		_w596_,
		_w598_,
		_w599_
	);
	LUT3 #(
		.INIT('h02)
	) name137 (
		\P1_reg0_reg[31]/NET0131 ,
		_w577_,
		_w584_,
		_w600_
	);
	LUT4 #(
		.INIT('hf53f)
	) name138 (
		\P1_reg1_reg[31]/NET0131 ,
		\P1_reg2_reg[31]/NET0131 ,
		_w577_,
		_w584_,
		_w601_
	);
	LUT4 #(
		.INIT('h0700)
	) name139 (
		_w585_,
		_w599_,
		_w600_,
		_w601_,
		_w602_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name140 (
		_w585_,
		_w599_,
		_w600_,
		_w601_,
		_w603_
	);
	LUT3 #(
		.INIT('h40)
	) name141 (
		_w489_,
		_w569_,
		_w602_,
		_w604_
	);
	LUT4 #(
		.INIT('h135f)
	) name142 (
		\P2_datao_reg[2]/NET0131 ,
		\P2_datao_reg[3]/NET0131 ,
		\si[2]_pad ,
		\si[3]_pad ,
		_w605_
	);
	LUT4 #(
		.INIT('h40f0)
	) name143 (
		_w490_,
		_w492_,
		_w498_,
		_w605_,
		_w606_
	);
	LUT4 #(
		.INIT('h135f)
	) name144 (
		\P2_datao_reg[4]/NET0131 ,
		\P2_datao_reg[5]/NET0131 ,
		\si[4]_pad ,
		\si[5]_pad ,
		_w607_
	);
	LUT3 #(
		.INIT('h40)
	) name145 (
		_w506_,
		_w495_,
		_w510_,
		_w608_
	);
	LUT4 #(
		.INIT('hec80)
	) name146 (
		\P2_datao_reg[8]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		\si[8]_pad ,
		\si[9]_pad ,
		_w609_
	);
	LUT4 #(
		.INIT('h135f)
	) name147 (
		\P2_datao_reg[6]/NET0131 ,
		\P2_datao_reg[7]/NET0131 ,
		\si[6]_pad ,
		\si[7]_pad ,
		_w610_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name148 (
		_w506_,
		_w510_,
		_w609_,
		_w610_,
		_w611_
	);
	LUT4 #(
		.INIT('h4f00)
	) name149 (
		_w606_,
		_w607_,
		_w608_,
		_w611_,
		_w612_
	);
	LUT4 #(
		.INIT('hfac8)
	) name150 (
		\P2_datao_reg[11]/NET0131 ,
		\P2_datao_reg[12]/NET0131 ,
		\si[11]_pad ,
		\si[12]_pad ,
		_w613_
	);
	LUT3 #(
		.INIT('h10)
	) name151 (
		_w520_,
		_w505_,
		_w613_,
		_w614_
	);
	LUT4 #(
		.INIT('hec80)
	) name152 (
		\P2_datao_reg[12]/NET0131 ,
		\P2_datao_reg[13]/NET0131 ,
		\si[12]_pad ,
		\si[13]_pad ,
		_w615_
	);
	LUT4 #(
		.INIT('h135f)
	) name153 (
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w616_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name154 (
		_w520_,
		_w613_,
		_w615_,
		_w616_,
		_w617_
	);
	LUT3 #(
		.INIT('hb0)
	) name155 (
		_w612_,
		_w614_,
		_w617_,
		_w618_
	);
	LUT4 #(
		.INIT('hfac8)
	) name156 (
		\P2_datao_reg[16]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w619_
	);
	LUT4 #(
		.INIT('hfac8)
	) name157 (
		\P2_datao_reg[14]/NET0131 ,
		\P2_datao_reg[15]/NET0131 ,
		\si[14]_pad ,
		\si[15]_pad ,
		_w620_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		_w619_,
		_w620_,
		_w621_
	);
	LUT4 #(
		.INIT('hfac8)
	) name159 (
		\P2_datao_reg[20]/NET0131 ,
		\P2_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w622_
	);
	LUT4 #(
		.INIT('hfac8)
	) name160 (
		\P2_datao_reg[18]/NET0131 ,
		\P2_datao_reg[19]/NET0131 ,
		\si[18]_pad ,
		\si[19]_pad ,
		_w623_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		_w622_,
		_w623_,
		_w624_
	);
	LUT4 #(
		.INIT('h8000)
	) name162 (
		_w619_,
		_w620_,
		_w622_,
		_w623_,
		_w625_
	);
	LUT4 #(
		.INIT('h4f00)
	) name163 (
		_w612_,
		_w614_,
		_w617_,
		_w625_,
		_w626_
	);
	LUT4 #(
		.INIT('hec80)
	) name164 (
		\P2_datao_reg[20]/NET0131 ,
		\P2_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w627_
	);
	LUT4 #(
		.INIT('hec80)
	) name165 (
		\P2_datao_reg[18]/NET0131 ,
		\P2_datao_reg[19]/NET0131 ,
		\si[18]_pad ,
		\si[19]_pad ,
		_w628_
	);
	LUT3 #(
		.INIT('h13)
	) name166 (
		_w622_,
		_w627_,
		_w628_,
		_w629_
	);
	LUT4 #(
		.INIT('hec80)
	) name167 (
		\P2_datao_reg[16]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w630_
	);
	LUT4 #(
		.INIT('hec80)
	) name168 (
		\P2_datao_reg[14]/NET0131 ,
		\P2_datao_reg[15]/NET0131 ,
		\si[14]_pad ,
		\si[15]_pad ,
		_w631_
	);
	LUT3 #(
		.INIT('h15)
	) name169 (
		_w630_,
		_w619_,
		_w631_,
		_w632_
	);
	LUT3 #(
		.INIT('hb0)
	) name170 (
		_w632_,
		_w624_,
		_w629_,
		_w633_
	);
	LUT4 #(
		.INIT('hfac8)
	) name171 (
		\P2_datao_reg[22]/NET0131 ,
		\P2_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w634_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		_w548_,
		_w634_,
		_w635_
	);
	LUT3 #(
		.INIT('h10)
	) name173 (
		_w546_,
		_w552_,
		_w555_,
		_w636_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		_w635_,
		_w636_,
		_w637_
	);
	LUT4 #(
		.INIT('hec80)
	) name175 (
		\P2_datao_reg[24]/NET0131 ,
		\P2_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w638_
	);
	LUT4 #(
		.INIT('hec80)
	) name176 (
		\P2_datao_reg[22]/NET0131 ,
		\P2_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w639_
	);
	LUT3 #(
		.INIT('h15)
	) name177 (
		_w638_,
		_w548_,
		_w639_,
		_w640_
	);
	LUT4 #(
		.INIT('h135f)
	) name178 (
		\P2_datao_reg[26]/NET0131 ,
		\P2_datao_reg[27]/NET0131 ,
		\si[26]_pad ,
		\si[27]_pad ,
		_w641_
	);
	LUT4 #(
		.INIT('h137f)
	) name179 (
		\P2_datao_reg[28]/NET0131 ,
		\P2_datao_reg[29]/NET0131 ,
		\si[28]_pad ,
		\si[29]_pad ,
		_w642_
	);
	LUT4 #(
		.INIT('hfb00)
	) name180 (
		_w552_,
		_w555_,
		_w641_,
		_w642_,
		_w643_
	);
	LUT3 #(
		.INIT('hb0)
	) name181 (
		_w640_,
		_w636_,
		_w643_,
		_w644_
	);
	LUT4 #(
		.INIT('h4f00)
	) name182 (
		_w626_,
		_w633_,
		_w637_,
		_w644_,
		_w645_
	);
	LUT4 #(
		.INIT('h5956)
	) name183 (
		\P2_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w568_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		_w489_,
		_w646_,
		_w647_
	);
	LUT3 #(
		.INIT('h08)
	) name185 (
		\P1_reg2_reg[30]/NET0131 ,
		_w577_,
		_w584_,
		_w648_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name186 (
		\P1_reg0_reg[30]/NET0131 ,
		\P1_reg1_reg[30]/NET0131 ,
		_w577_,
		_w584_,
		_w649_
	);
	LUT4 #(
		.INIT('h0700)
	) name187 (
		_w585_,
		_w599_,
		_w648_,
		_w649_,
		_w650_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name188 (
		_w585_,
		_w599_,
		_w648_,
		_w649_,
		_w651_
	);
	LUT3 #(
		.INIT('h10)
	) name189 (
		_w489_,
		_w646_,
		_w650_,
		_w652_
	);
	LUT4 #(
		.INIT('h00f4)
	) name190 (
		_w489_,
		_w569_,
		_w602_,
		_w652_,
		_w653_
	);
	LUT3 #(
		.INIT('hd0)
	) name191 (
		_w537_,
		_w545_,
		_w559_,
		_w654_
	);
	LUT4 #(
		.INIT('h4454)
	) name192 (
		_w553_,
		_w558_,
		_w549_,
		_w654_,
		_w655_
	);
	LUT3 #(
		.INIT('h51)
	) name193 (
		_w554_,
		_w562_,
		_w655_,
		_w656_
	);
	LUT4 #(
		.INIT('h0155)
	) name194 (
		_w525_,
		_w526_,
		_w514_,
		_w613_,
		_w657_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		_w495_,
		_w510_,
		_w658_
	);
	LUT4 #(
		.INIT('h0155)
	) name196 (
		_w515_,
		_w516_,
		_w500_,
		_w510_,
		_w659_
	);
	LUT4 #(
		.INIT('h1f00)
	) name197 (
		_w501_,
		_w606_,
		_w658_,
		_w659_,
		_w660_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		_w507_,
		_w613_,
		_w661_
	);
	LUT3 #(
		.INIT('h8a)
	) name199 (
		_w657_,
		_w660_,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		_w521_,
		_w532_,
		_w663_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		_w530_,
		_w535_,
		_w664_
	);
	LUT4 #(
		.INIT('h8000)
	) name202 (
		_w521_,
		_w530_,
		_w532_,
		_w535_,
		_w665_
	);
	LUT4 #(
		.INIT('h7500)
	) name203 (
		_w657_,
		_w660_,
		_w661_,
		_w665_,
		_w666_
	);
	LUT3 #(
		.INIT('h07)
	) name204 (
		_w540_,
		_w535_,
		_w538_,
		_w667_
	);
	LUT3 #(
		.INIT('h07)
	) name205 (
		_w524_,
		_w532_,
		_w541_,
		_w668_
	);
	LUT3 #(
		.INIT('hb0)
	) name206 (
		_w668_,
		_w664_,
		_w667_,
		_w669_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		_w534_,
		_w555_,
		_w670_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		_w550_,
		_w670_,
		_w671_
	);
	LUT4 #(
		.INIT('h040f)
	) name209 (
		_w666_,
		_w669_,
		_w656_,
		_w671_,
		_w672_
	);
	LUT4 #(
		.INIT('h5956)
	) name210 (
		\P2_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w568_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		_w489_,
		_w673_,
		_w674_
	);
	LUT3 #(
		.INIT('h08)
	) name212 (
		\P1_reg2_reg[29]/NET0131 ,
		_w577_,
		_w584_,
		_w675_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name213 (
		\P1_reg0_reg[29]/NET0131 ,
		\P1_reg1_reg[29]/NET0131 ,
		_w577_,
		_w584_,
		_w676_
	);
	LUT4 #(
		.INIT('h0700)
	) name214 (
		_w585_,
		_w599_,
		_w675_,
		_w676_,
		_w677_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name215 (
		_w585_,
		_w599_,
		_w675_,
		_w676_,
		_w678_
	);
	LUT3 #(
		.INIT('h10)
	) name216 (
		_w489_,
		_w673_,
		_w677_,
		_w679_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		\P2_datao_reg[28]/NET0131 ,
		_w568_,
		_w680_
	);
	LUT2 #(
		.INIT('h6)
	) name218 (
		\P2_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w681_
	);
	LUT3 #(
		.INIT('h07)
	) name219 (
		_w630_,
		_w623_,
		_w628_,
		_w682_
	);
	LUT3 #(
		.INIT('h04)
	) name220 (
		_w519_,
		_w521_,
		_w531_,
		_w683_
	);
	LUT3 #(
		.INIT('hc4)
	) name221 (
		_w495_,
		_w610_,
		_w607_,
		_w684_
	);
	LUT4 #(
		.INIT('h2033)
	) name222 (
		_w495_,
		_w509_,
		_w606_,
		_w684_,
		_w685_
	);
	LUT3 #(
		.INIT('h02)
	) name223 (
		_w507_,
		_w508_,
		_w522_,
		_w686_
	);
	LUT4 #(
		.INIT('hfac8)
	) name224 (
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w687_
	);
	LUT4 #(
		.INIT('h0155)
	) name225 (
		_w526_,
		_w513_,
		_w609_,
		_w687_,
		_w688_
	);
	LUT3 #(
		.INIT('h15)
	) name226 (
		_w631_,
		_w615_,
		_w620_,
		_w689_
	);
	LUT3 #(
		.INIT('hd0)
	) name227 (
		_w683_,
		_w688_,
		_w689_,
		_w690_
	);
	LUT4 #(
		.INIT('h7f00)
	) name228 (
		_w683_,
		_w685_,
		_w686_,
		_w690_,
		_w691_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		_w619_,
		_w623_,
		_w692_
	);
	LUT3 #(
		.INIT('h8c)
	) name230 (
		_w691_,
		_w682_,
		_w692_,
		_w693_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		_w622_,
		_w634_,
		_w694_
	);
	LUT3 #(
		.INIT('h04)
	) name232 (
		_w546_,
		_w548_,
		_w553_,
		_w695_
	);
	LUT2 #(
		.INIT('h8)
	) name233 (
		_w694_,
		_w695_,
		_w696_
	);
	LUT4 #(
		.INIT('h7300)
	) name234 (
		_w691_,
		_w682_,
		_w692_,
		_w696_,
		_w697_
	);
	LUT3 #(
		.INIT('h13)
	) name235 (
		_w627_,
		_w639_,
		_w634_,
		_w698_
	);
	LUT3 #(
		.INIT('hb0)
	) name236 (
		_w546_,
		_w638_,
		_w641_,
		_w699_
	);
	LUT4 #(
		.INIT('h0455)
	) name237 (
		_w553_,
		_w549_,
		_w698_,
		_w699_,
		_w700_
	);
	LUT4 #(
		.INIT('h1114)
	) name238 (
		_w568_,
		_w681_,
		_w697_,
		_w700_,
		_w701_
	);
	LUT3 #(
		.INIT('h54)
	) name239 (
		_w489_,
		_w680_,
		_w701_,
		_w702_
	);
	LUT4 #(
		.INIT('h8000)
	) name240 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_reg3_reg[26]/NET0131 ,
		_w593_,
		_w596_,
		_w703_
	);
	LUT4 #(
		.INIT('h00ec)
	) name241 (
		\P1_reg3_reg[27]/NET0131 ,
		\P1_reg3_reg[28]/NET0131 ,
		_w703_,
		_w599_,
		_w704_
	);
	LUT3 #(
		.INIT('h08)
	) name242 (
		\P1_reg2_reg[28]/NET0131 ,
		_w577_,
		_w584_,
		_w705_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name243 (
		\P1_reg0_reg[28]/NET0131 ,
		\P1_reg1_reg[28]/NET0131 ,
		_w577_,
		_w584_,
		_w706_
	);
	LUT2 #(
		.INIT('h4)
	) name244 (
		_w705_,
		_w706_,
		_w707_
	);
	LUT3 #(
		.INIT('h70)
	) name245 (
		_w585_,
		_w704_,
		_w707_,
		_w708_
	);
	LUT3 #(
		.INIT('h8f)
	) name246 (
		_w585_,
		_w704_,
		_w707_,
		_w709_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		_w702_,
		_w708_,
		_w710_
	);
	LUT3 #(
		.INIT('h01)
	) name248 (
		_w679_,
		_w702_,
		_w708_,
		_w711_
	);
	LUT3 #(
		.INIT('h0e)
	) name249 (
		_w489_,
		_w646_,
		_w650_,
		_w712_
	);
	LUT3 #(
		.INIT('h0e)
	) name250 (
		_w489_,
		_w673_,
		_w677_,
		_w713_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		_w712_,
		_w713_,
		_w714_
	);
	LUT4 #(
		.INIT('h1303)
	) name252 (
		_w711_,
		_w604_,
		_w653_,
		_w714_,
		_w715_
	);
	LUT3 #(
		.INIT('hb0)
	) name253 (
		_w529_,
		_w533_,
		_w542_,
		_w716_
	);
	LUT4 #(
		.INIT('h5956)
	) name254 (
		\P2_datao_reg[19]/NET0131 ,
		\si[19]_pad ,
		_w568_,
		_w716_,
		_w717_
	);
	LUT4 #(
		.INIT('h5999)
	) name255 (
		\P1_IR_reg[19]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w469_,
		_w474_,
		_w718_
	);
	LUT3 #(
		.INIT('h04)
	) name256 (
		_w718_,
		_w479_,
		_w488_,
		_w719_
	);
	LUT3 #(
		.INIT('h0e)
	) name257 (
		_w489_,
		_w717_,
		_w719_,
		_w720_
	);
	LUT3 #(
		.INIT('h6c)
	) name258 (
		\P1_reg3_reg[18]/NET0131 ,
		\P1_reg3_reg[19]/NET0131 ,
		_w591_,
		_w721_
	);
	LUT3 #(
		.INIT('h08)
	) name259 (
		\P1_reg2_reg[19]/NET0131 ,
		_w577_,
		_w584_,
		_w722_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name260 (
		\P1_reg0_reg[19]/NET0131 ,
		\P1_reg1_reg[19]/NET0131 ,
		_w577_,
		_w584_,
		_w723_
	);
	LUT4 #(
		.INIT('h1500)
	) name261 (
		_w722_,
		_w585_,
		_w721_,
		_w723_,
		_w724_
	);
	LUT4 #(
		.INIT('heaff)
	) name262 (
		_w722_,
		_w585_,
		_w721_,
		_w723_,
		_w725_
	);
	LUT4 #(
		.INIT('hf100)
	) name263 (
		_w489_,
		_w717_,
		_w719_,
		_w724_,
		_w726_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		\P2_datao_reg[18]/NET0131 ,
		_w568_,
		_w727_
	);
	LUT2 #(
		.INIT('h6)
	) name265 (
		\P2_datao_reg[18]/NET0131 ,
		\si[18]_pad ,
		_w728_
	);
	LUT4 #(
		.INIT('h4f00)
	) name266 (
		_w612_,
		_w614_,
		_w617_,
		_w621_,
		_w729_
	);
	LUT4 #(
		.INIT('h1141)
	) name267 (
		_w568_,
		_w728_,
		_w632_,
		_w729_,
		_w730_
	);
	LUT3 #(
		.INIT('he0)
	) name268 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[17]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w731_
	);
	LUT3 #(
		.INIT('h56)
	) name269 (
		\P1_IR_reg[18]/NET0131 ,
		_w482_,
		_w731_,
		_w732_
	);
	LUT3 #(
		.INIT('h20)
	) name270 (
		_w479_,
		_w488_,
		_w732_,
		_w733_
	);
	LUT4 #(
		.INIT('h00ab)
	) name271 (
		_w489_,
		_w727_,
		_w730_,
		_w733_,
		_w734_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name272 (
		\P1_reg3_reg[18]/NET0131 ,
		_w588_,
		_w589_,
		_w590_,
		_w735_
	);
	LUT3 #(
		.INIT('h80)
	) name273 (
		_w577_,
		_w584_,
		_w735_,
		_w736_
	);
	LUT3 #(
		.INIT('h20)
	) name274 (
		\P1_reg1_reg[18]/NET0131 ,
		_w577_,
		_w584_,
		_w737_
	);
	LUT4 #(
		.INIT('hff35)
	) name275 (
		\P1_reg0_reg[18]/NET0131 ,
		\P1_reg2_reg[18]/NET0131 ,
		_w577_,
		_w584_,
		_w738_
	);
	LUT3 #(
		.INIT('h10)
	) name276 (
		_w737_,
		_w736_,
		_w738_,
		_w739_
	);
	LUT3 #(
		.INIT('hef)
	) name277 (
		_w737_,
		_w736_,
		_w738_,
		_w740_
	);
	LUT2 #(
		.INIT('h4)
	) name278 (
		_w734_,
		_w739_,
		_w741_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		\P2_datao_reg[17]/NET0131 ,
		_w568_,
		_w742_
	);
	LUT2 #(
		.INIT('h6)
	) name280 (
		\P2_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w743_
	);
	LUT4 #(
		.INIT('h7500)
	) name281 (
		_w657_,
		_w660_,
		_w661_,
		_w663_,
		_w744_
	);
	LUT4 #(
		.INIT('h1141)
	) name282 (
		_w568_,
		_w743_,
		_w668_,
		_w744_,
		_w745_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name283 (
		\P1_IR_reg[31]/NET0131 ,
		_w469_,
		_w470_,
		_w579_,
		_w746_
	);
	LUT2 #(
		.INIT('h6)
	) name284 (
		\P1_IR_reg[17]/NET0131 ,
		_w746_,
		_w747_
	);
	LUT3 #(
		.INIT('h20)
	) name285 (
		_w479_,
		_w488_,
		_w747_,
		_w748_
	);
	LUT4 #(
		.INIT('h00ab)
	) name286 (
		_w489_,
		_w742_,
		_w745_,
		_w748_,
		_w749_
	);
	LUT4 #(
		.INIT('h8000)
	) name287 (
		\P1_reg3_reg[15]/NET0131 ,
		\P1_reg3_reg[16]/NET0131 ,
		_w588_,
		_w589_,
		_w750_
	);
	LUT3 #(
		.INIT('h32)
	) name288 (
		\P1_reg3_reg[17]/NET0131 ,
		_w591_,
		_w750_,
		_w751_
	);
	LUT3 #(
		.INIT('h20)
	) name289 (
		\P1_reg1_reg[17]/NET0131 ,
		_w577_,
		_w584_,
		_w752_
	);
	LUT4 #(
		.INIT('hff35)
	) name290 (
		\P1_reg0_reg[17]/NET0131 ,
		\P1_reg2_reg[17]/NET0131 ,
		_w577_,
		_w584_,
		_w753_
	);
	LUT4 #(
		.INIT('h1300)
	) name291 (
		_w585_,
		_w752_,
		_w751_,
		_w753_,
		_w754_
	);
	LUT4 #(
		.INIT('hecff)
	) name292 (
		_w585_,
		_w752_,
		_w751_,
		_w753_,
		_w755_
	);
	LUT4 #(
		.INIT('h5956)
	) name293 (
		\P2_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w568_,
		_w691_,
		_w756_
	);
	LUT2 #(
		.INIT('h6)
	) name294 (
		\P1_IR_reg[16]/NET0131 ,
		_w482_,
		_w757_
	);
	LUT3 #(
		.INIT('h20)
	) name295 (
		_w479_,
		_w488_,
		_w757_,
		_w758_
	);
	LUT3 #(
		.INIT('h0e)
	) name296 (
		_w489_,
		_w756_,
		_w758_,
		_w759_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name297 (
		\P1_reg3_reg[15]/NET0131 ,
		\P1_reg3_reg[16]/NET0131 ,
		_w588_,
		_w589_,
		_w760_
	);
	LUT3 #(
		.INIT('h80)
	) name298 (
		_w577_,
		_w584_,
		_w760_,
		_w761_
	);
	LUT3 #(
		.INIT('h08)
	) name299 (
		\P1_reg2_reg[16]/NET0131 ,
		_w577_,
		_w584_,
		_w762_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name300 (
		\P1_reg0_reg[16]/NET0131 ,
		\P1_reg1_reg[16]/NET0131 ,
		_w577_,
		_w584_,
		_w763_
	);
	LUT3 #(
		.INIT('h10)
	) name301 (
		_w762_,
		_w761_,
		_w763_,
		_w764_
	);
	LUT3 #(
		.INIT('hef)
	) name302 (
		_w762_,
		_w761_,
		_w763_,
		_w765_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name303 (
		_w749_,
		_w754_,
		_w759_,
		_w764_,
		_w766_
	);
	LUT4 #(
		.INIT('h22b2)
	) name304 (
		_w749_,
		_w754_,
		_w759_,
		_w764_,
		_w767_
	);
	LUT3 #(
		.INIT('h10)
	) name305 (
		_w726_,
		_w741_,
		_w767_,
		_w768_
	);
	LUT2 #(
		.INIT('h2)
	) name306 (
		_w734_,
		_w739_,
		_w769_
	);
	LUT4 #(
		.INIT('h000e)
	) name307 (
		_w489_,
		_w717_,
		_w719_,
		_w724_,
		_w770_
	);
	LUT3 #(
		.INIT('h54)
	) name308 (
		_w726_,
		_w769_,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		_w768_,
		_w771_,
		_w772_
	);
	LUT2 #(
		.INIT('h8)
	) name310 (
		\P2_datao_reg[22]/NET0131 ,
		_w568_,
		_w773_
	);
	LUT2 #(
		.INIT('h6)
	) name311 (
		\P2_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w774_
	);
	LUT4 #(
		.INIT('h1045)
	) name312 (
		_w568_,
		_w626_,
		_w633_,
		_w774_,
		_w775_
	);
	LUT3 #(
		.INIT('h54)
	) name313 (
		_w489_,
		_w773_,
		_w775_,
		_w776_
	);
	LUT3 #(
		.INIT('h6a)
	) name314 (
		\P1_reg3_reg[22]/NET0131 ,
		_w593_,
		_w594_,
		_w777_
	);
	LUT3 #(
		.INIT('h02)
	) name315 (
		\P1_reg0_reg[22]/NET0131 ,
		_w577_,
		_w584_,
		_w778_
	);
	LUT4 #(
		.INIT('hf53f)
	) name316 (
		\P1_reg1_reg[22]/NET0131 ,
		\P1_reg2_reg[22]/NET0131 ,
		_w577_,
		_w584_,
		_w779_
	);
	LUT4 #(
		.INIT('h1300)
	) name317 (
		_w585_,
		_w778_,
		_w777_,
		_w779_,
		_w780_
	);
	LUT4 #(
		.INIT('hecff)
	) name318 (
		_w585_,
		_w778_,
		_w777_,
		_w779_,
		_w781_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		_w776_,
		_w780_,
		_w782_
	);
	LUT4 #(
		.INIT('h5956)
	) name320 (
		\P2_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w568_,
		_w544_,
		_w783_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		_w489_,
		_w783_,
		_w784_
	);
	LUT4 #(
		.INIT('h8000)
	) name322 (
		\P1_reg3_reg[22]/NET0131 ,
		\P1_reg3_reg[23]/NET0131 ,
		_w593_,
		_w594_,
		_w785_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name323 (
		\P1_reg3_reg[22]/NET0131 ,
		\P1_reg3_reg[23]/NET0131 ,
		_w593_,
		_w594_,
		_w786_
	);
	LUT3 #(
		.INIT('h08)
	) name324 (
		\P1_reg2_reg[23]/NET0131 ,
		_w577_,
		_w584_,
		_w787_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name325 (
		\P1_reg0_reg[23]/NET0131 ,
		\P1_reg1_reg[23]/NET0131 ,
		_w577_,
		_w584_,
		_w788_
	);
	LUT4 #(
		.INIT('h1300)
	) name326 (
		_w585_,
		_w787_,
		_w786_,
		_w788_,
		_w789_
	);
	LUT4 #(
		.INIT('hecff)
	) name327 (
		_w585_,
		_w787_,
		_w786_,
		_w788_,
		_w790_
	);
	LUT3 #(
		.INIT('h10)
	) name328 (
		_w489_,
		_w783_,
		_w789_,
		_w791_
	);
	LUT2 #(
		.INIT('h1)
	) name329 (
		_w782_,
		_w791_,
		_w792_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		\P2_datao_reg[21]/NET0131 ,
		_w568_,
		_w793_
	);
	LUT2 #(
		.INIT('h6)
	) name331 (
		\P2_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w794_
	);
	LUT4 #(
		.INIT('h1045)
	) name332 (
		_w568_,
		_w666_,
		_w669_,
		_w794_,
		_w795_
	);
	LUT3 #(
		.INIT('h54)
	) name333 (
		_w489_,
		_w793_,
		_w795_,
		_w796_
	);
	LUT3 #(
		.INIT('h6c)
	) name334 (
		\P1_reg3_reg[20]/NET0131 ,
		\P1_reg3_reg[21]/NET0131 ,
		_w593_,
		_w797_
	);
	LUT3 #(
		.INIT('h08)
	) name335 (
		\P1_reg2_reg[21]/NET0131 ,
		_w577_,
		_w584_,
		_w798_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name336 (
		\P1_reg0_reg[21]/NET0131 ,
		\P1_reg1_reg[21]/NET0131 ,
		_w577_,
		_w584_,
		_w799_
	);
	LUT4 #(
		.INIT('h1300)
	) name337 (
		_w585_,
		_w798_,
		_w797_,
		_w799_,
		_w800_
	);
	LUT4 #(
		.INIT('hecff)
	) name338 (
		_w585_,
		_w798_,
		_w797_,
		_w799_,
		_w801_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		_w796_,
		_w800_,
		_w802_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		_w796_,
		_w800_,
		_w803_
	);
	LUT4 #(
		.INIT('h5956)
	) name341 (
		\P2_datao_reg[20]/NET0131 ,
		\si[20]_pad ,
		_w568_,
		_w693_,
		_w804_
	);
	LUT2 #(
		.INIT('h1)
	) name342 (
		_w489_,
		_w804_,
		_w805_
	);
	LUT2 #(
		.INIT('h6)
	) name343 (
		\P1_reg3_reg[20]/NET0131 ,
		_w593_,
		_w806_
	);
	LUT4 #(
		.INIT('h4080)
	) name344 (
		\P1_reg3_reg[20]/NET0131 ,
		_w577_,
		_w584_,
		_w593_,
		_w807_
	);
	LUT3 #(
		.INIT('h02)
	) name345 (
		\P1_reg0_reg[20]/NET0131 ,
		_w577_,
		_w584_,
		_w808_
	);
	LUT4 #(
		.INIT('hf53f)
	) name346 (
		\P1_reg1_reg[20]/NET0131 ,
		\P1_reg2_reg[20]/NET0131 ,
		_w577_,
		_w584_,
		_w809_
	);
	LUT3 #(
		.INIT('h10)
	) name347 (
		_w808_,
		_w807_,
		_w809_,
		_w810_
	);
	LUT3 #(
		.INIT('hef)
	) name348 (
		_w808_,
		_w807_,
		_w809_,
		_w811_
	);
	LUT3 #(
		.INIT('h0e)
	) name349 (
		_w489_,
		_w804_,
		_w810_,
		_w812_
	);
	LUT3 #(
		.INIT('h54)
	) name350 (
		_w802_,
		_w803_,
		_w812_,
		_w813_
	);
	LUT3 #(
		.INIT('h0e)
	) name351 (
		_w489_,
		_w783_,
		_w789_,
		_w814_
	);
	LUT2 #(
		.INIT('h1)
	) name352 (
		_w776_,
		_w780_,
		_w815_
	);
	LUT3 #(
		.INIT('h54)
	) name353 (
		_w791_,
		_w814_,
		_w815_,
		_w816_
	);
	LUT3 #(
		.INIT('h07)
	) name354 (
		_w792_,
		_w813_,
		_w816_,
		_w817_
	);
	LUT3 #(
		.INIT('h10)
	) name355 (
		_w489_,
		_w804_,
		_w810_,
		_w818_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w802_,
		_w818_,
		_w819_
	);
	LUT4 #(
		.INIT('heee0)
	) name357 (
		_w776_,
		_w780_,
		_w796_,
		_w800_,
		_w820_
	);
	LUT3 #(
		.INIT('he0)
	) name358 (
		_w802_,
		_w818_,
		_w820_,
		_w821_
	);
	LUT3 #(
		.INIT('h31)
	) name359 (
		_w792_,
		_w814_,
		_w821_,
		_w822_
	);
	LUT3 #(
		.INIT('h07)
	) name360 (
		_w772_,
		_w817_,
		_w822_,
		_w823_
	);
	LUT4 #(
		.INIT('hf53f)
	) name361 (
		\P1_reg1_reg[15]/NET0131 ,
		\P1_reg2_reg[15]/NET0131 ,
		_w577_,
		_w584_,
		_w824_
	);
	LUT3 #(
		.INIT('h6a)
	) name362 (
		\P1_reg3_reg[15]/NET0131 ,
		_w588_,
		_w589_,
		_w825_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name363 (
		\P1_reg0_reg[15]/NET0131 ,
		_w577_,
		_w584_,
		_w825_,
		_w826_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		_w824_,
		_w826_,
		_w827_
	);
	LUT2 #(
		.INIT('h7)
	) name365 (
		_w824_,
		_w826_,
		_w828_
	);
	LUT4 #(
		.INIT('h5956)
	) name366 (
		\P2_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w568_,
		_w529_,
		_w829_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		\P1_IR_reg[31]/NET0131 ,
		_w472_,
		_w830_
	);
	LUT4 #(
		.INIT('h55a6)
	) name368 (
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w469_,
		_w830_,
		_w831_
	);
	LUT3 #(
		.INIT('h20)
	) name369 (
		_w479_,
		_w488_,
		_w831_,
		_w832_
	);
	LUT3 #(
		.INIT('h0e)
	) name370 (
		_w489_,
		_w829_,
		_w832_,
		_w833_
	);
	LUT4 #(
		.INIT('hff35)
	) name371 (
		\P1_reg0_reg[14]/NET0131 ,
		\P1_reg2_reg[14]/NET0131 ,
		_w577_,
		_w584_,
		_w834_
	);
	LUT3 #(
		.INIT('h6c)
	) name372 (
		\P1_reg3_reg[13]/NET0131 ,
		\P1_reg3_reg[14]/NET0131 ,
		_w588_,
		_w835_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name373 (
		\P1_reg1_reg[14]/NET0131 ,
		_w577_,
		_w584_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h8)
	) name374 (
		_w834_,
		_w836_,
		_w837_
	);
	LUT2 #(
		.INIT('h7)
	) name375 (
		_w834_,
		_w836_,
		_w838_
	);
	LUT4 #(
		.INIT('h5956)
	) name376 (
		\P2_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w568_,
		_w618_,
		_w839_
	);
	LUT4 #(
		.INIT('h5999)
	) name377 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w468_,
		_w481_,
		_w840_
	);
	LUT3 #(
		.INIT('h02)
	) name378 (
		_w479_,
		_w488_,
		_w840_,
		_w841_
	);
	LUT3 #(
		.INIT('h0e)
	) name379 (
		_w489_,
		_w839_,
		_w841_,
		_w842_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name380 (
		_w827_,
		_w833_,
		_w837_,
		_w842_,
		_w843_
	);
	LUT2 #(
		.INIT('h6)
	) name381 (
		\P1_reg3_reg[13]/NET0131 ,
		_w588_,
		_w844_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name382 (
		\P1_reg0_reg[13]/NET0131 ,
		_w577_,
		_w584_,
		_w844_,
		_w845_
	);
	LUT4 #(
		.INIT('hf53f)
	) name383 (
		\P1_reg1_reg[13]/NET0131 ,
		\P1_reg2_reg[13]/NET0131 ,
		_w577_,
		_w584_,
		_w846_
	);
	LUT2 #(
		.INIT('h8)
	) name384 (
		_w845_,
		_w846_,
		_w847_
	);
	LUT2 #(
		.INIT('h7)
	) name385 (
		_w845_,
		_w846_,
		_w848_
	);
	LUT4 #(
		.INIT('h5956)
	) name386 (
		\P2_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w568_,
		_w662_,
		_w849_
	);
	LUT4 #(
		.INIT('ha666)
	) name387 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w469_,
		_w470_,
		_w850_
	);
	LUT3 #(
		.INIT('h20)
	) name388 (
		_w479_,
		_w488_,
		_w850_,
		_w851_
	);
	LUT3 #(
		.INIT('h0e)
	) name389 (
		_w489_,
		_w849_,
		_w851_,
		_w852_
	);
	LUT4 #(
		.INIT('h78f0)
	) name390 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_reg3_reg[11]/NET0131 ,
		\P1_reg3_reg[12]/NET0131 ,
		_w587_,
		_w853_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name391 (
		\P1_reg1_reg[12]/NET0131 ,
		_w577_,
		_w584_,
		_w853_,
		_w854_
	);
	LUT4 #(
		.INIT('hff35)
	) name392 (
		\P1_reg0_reg[12]/NET0131 ,
		\P1_reg2_reg[12]/NET0131 ,
		_w577_,
		_w584_,
		_w855_
	);
	LUT2 #(
		.INIT('h8)
	) name393 (
		_w854_,
		_w855_,
		_w856_
	);
	LUT2 #(
		.INIT('h7)
	) name394 (
		_w854_,
		_w855_,
		_w857_
	);
	LUT3 #(
		.INIT('h70)
	) name395 (
		_w685_,
		_w686_,
		_w688_,
		_w858_
	);
	LUT4 #(
		.INIT('h5956)
	) name396 (
		\P2_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w568_,
		_w858_,
		_w859_
	);
	LUT4 #(
		.INIT('h4000)
	) name397 (
		\P1_IR_reg[4]/NET0131 ,
		_w464_,
		_w466_,
		_w467_,
		_w860_
	);
	LUT3 #(
		.INIT('he0)
	) name398 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w861_
	);
	LUT4 #(
		.INIT('h55a6)
	) name399 (
		\P1_IR_reg[12]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w860_,
		_w861_,
		_w862_
	);
	LUT3 #(
		.INIT('h20)
	) name400 (
		_w479_,
		_w488_,
		_w862_,
		_w863_
	);
	LUT3 #(
		.INIT('h0e)
	) name401 (
		_w489_,
		_w859_,
		_w863_,
		_w864_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name402 (
		_w847_,
		_w852_,
		_w856_,
		_w864_,
		_w865_
	);
	LUT4 #(
		.INIT('h4d44)
	) name403 (
		_w847_,
		_w852_,
		_w856_,
		_w864_,
		_w866_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		_w827_,
		_w833_,
		_w867_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name405 (
		_w827_,
		_w833_,
		_w837_,
		_w842_,
		_w868_
	);
	LUT4 #(
		.INIT('h4d44)
	) name406 (
		_w827_,
		_w833_,
		_w837_,
		_w842_,
		_w869_
	);
	LUT3 #(
		.INIT('h07)
	) name407 (
		_w843_,
		_w866_,
		_w869_,
		_w870_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name408 (
		_w847_,
		_w852_,
		_w856_,
		_w864_,
		_w871_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		_w843_,
		_w871_,
		_w872_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name410 (
		\P1_reg0_reg[11]/NET0131 ,
		\P1_reg1_reg[11]/NET0131 ,
		_w577_,
		_w584_,
		_w873_
	);
	LUT3 #(
		.INIT('h6c)
	) name411 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_reg3_reg[11]/NET0131 ,
		_w587_,
		_w874_
	);
	LUT4 #(
		.INIT('h37f7)
	) name412 (
		\P1_reg2_reg[11]/NET0131 ,
		_w577_,
		_w584_,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		_w873_,
		_w875_,
		_w876_
	);
	LUT2 #(
		.INIT('h7)
	) name414 (
		_w873_,
		_w875_,
		_w877_
	);
	LUT2 #(
		.INIT('h8)
	) name415 (
		\P2_datao_reg[11]/NET0131 ,
		_w568_,
		_w878_
	);
	LUT2 #(
		.INIT('h6)
	) name416 (
		\P2_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w879_
	);
	LUT4 #(
		.INIT('h1045)
	) name417 (
		_w568_,
		_w512_,
		_w518_,
		_w879_,
		_w880_
	);
	LUT4 #(
		.INIT('hddd0)
	) name418 (
		_w479_,
		_w488_,
		_w878_,
		_w880_,
		_w881_
	);
	LUT3 #(
		.INIT('ha6)
	) name419 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w469_,
		_w882_
	);
	LUT3 #(
		.INIT('h20)
	) name420 (
		_w479_,
		_w488_,
		_w882_,
		_w883_
	);
	LUT2 #(
		.INIT('h1)
	) name421 (
		_w881_,
		_w883_,
		_w884_
	);
	LUT4 #(
		.INIT('h8880)
	) name422 (
		_w873_,
		_w875_,
		_w881_,
		_w883_,
		_w885_
	);
	LUT2 #(
		.INIT('h6)
	) name423 (
		\P1_reg3_reg[10]/NET0131 ,
		_w587_,
		_w886_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name424 (
		\P1_reg0_reg[10]/NET0131 ,
		_w577_,
		_w584_,
		_w886_,
		_w887_
	);
	LUT4 #(
		.INIT('hf53f)
	) name425 (
		\P1_reg1_reg[10]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w577_,
		_w584_,
		_w888_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		_w887_,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h7)
	) name427 (
		_w887_,
		_w888_,
		_w890_
	);
	LUT4 #(
		.INIT('h5956)
	) name428 (
		\P2_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w568_,
		_w612_,
		_w891_
	);
	LUT3 #(
		.INIT('h59)
	) name429 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w860_,
		_w892_
	);
	LUT4 #(
		.INIT('hf2d0)
	) name430 (
		_w479_,
		_w488_,
		_w891_,
		_w892_,
		_w893_
	);
	LUT3 #(
		.INIT('h08)
	) name431 (
		_w887_,
		_w888_,
		_w893_,
		_w894_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w885_,
		_w894_,
		_w895_
	);
	LUT4 #(
		.INIT('hf53f)
	) name433 (
		\P1_reg1_reg[9]/NET0131 ,
		\P1_reg2_reg[9]/NET0131 ,
		_w577_,
		_w584_,
		_w896_
	);
	LUT4 #(
		.INIT('h78f0)
	) name434 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_reg3_reg[8]/NET0131 ,
		\P1_reg3_reg[9]/NET0131 ,
		_w586_,
		_w897_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name435 (
		\P1_reg0_reg[9]/NET0131 ,
		_w577_,
		_w584_,
		_w897_,
		_w898_
	);
	LUT2 #(
		.INIT('h8)
	) name436 (
		_w896_,
		_w898_,
		_w899_
	);
	LUT2 #(
		.INIT('h7)
	) name437 (
		_w896_,
		_w898_,
		_w900_
	);
	LUT4 #(
		.INIT('h5956)
	) name438 (
		\P2_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w568_,
		_w660_,
		_w901_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name439 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		_w466_,
		_w467_,
		_w902_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[8]/NET0131 ,
		_w903_
	);
	LUT3 #(
		.INIT('h56)
	) name441 (
		\P1_IR_reg[9]/NET0131 ,
		_w902_,
		_w903_,
		_w904_
	);
	LUT4 #(
		.INIT('hd0f2)
	) name442 (
		_w479_,
		_w488_,
		_w901_,
		_w904_,
		_w905_
	);
	LUT3 #(
		.INIT('h08)
	) name443 (
		_w896_,
		_w898_,
		_w905_,
		_w906_
	);
	LUT3 #(
		.INIT('h70)
	) name444 (
		_w896_,
		_w898_,
		_w905_,
		_w907_
	);
	LUT3 #(
		.INIT('h6c)
	) name445 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_reg3_reg[8]/NET0131 ,
		_w586_,
		_w908_
	);
	LUT4 #(
		.INIT('h37f7)
	) name446 (
		\P1_reg2_reg[8]/NET0131 ,
		_w577_,
		_w584_,
		_w908_,
		_w909_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name447 (
		\P1_reg0_reg[8]/NET0131 ,
		\P1_reg1_reg[8]/NET0131 ,
		_w577_,
		_w584_,
		_w910_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		_w909_,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h7)
	) name449 (
		_w909_,
		_w910_,
		_w912_
	);
	LUT4 #(
		.INIT('h5659)
	) name450 (
		\P2_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w568_,
		_w685_,
		_w913_
	);
	LUT2 #(
		.INIT('h9)
	) name451 (
		\P1_IR_reg[8]/NET0131 ,
		_w902_,
		_w914_
	);
	LUT4 #(
		.INIT('hf2d0)
	) name452 (
		_w479_,
		_w488_,
		_w913_,
		_w914_,
		_w915_
	);
	LUT3 #(
		.INIT('h70)
	) name453 (
		_w909_,
		_w910_,
		_w915_,
		_w916_
	);
	LUT3 #(
		.INIT('h54)
	) name454 (
		_w906_,
		_w907_,
		_w916_,
		_w917_
	);
	LUT3 #(
		.INIT('h70)
	) name455 (
		_w887_,
		_w888_,
		_w893_,
		_w918_
	);
	LUT4 #(
		.INIT('h0007)
	) name456 (
		_w873_,
		_w875_,
		_w881_,
		_w883_,
		_w919_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		_w918_,
		_w919_,
		_w920_
	);
	LUT3 #(
		.INIT('h54)
	) name458 (
		_w885_,
		_w918_,
		_w919_,
		_w921_
	);
	LUT3 #(
		.INIT('h07)
	) name459 (
		_w895_,
		_w917_,
		_w921_,
		_w922_
	);
	LUT3 #(
		.INIT('ha2)
	) name460 (
		_w870_,
		_w872_,
		_w922_,
		_w923_
	);
	LUT4 #(
		.INIT('hff35)
	) name461 (
		\P1_reg0_reg[6]/NET0131 ,
		\P1_reg2_reg[6]/NET0131 ,
		_w577_,
		_w584_,
		_w924_
	);
	LUT4 #(
		.INIT('h7f80)
	) name462 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		\P1_reg3_reg[5]/NET0131 ,
		\P1_reg3_reg[6]/NET0131 ,
		_w925_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name463 (
		\P1_reg1_reg[6]/NET0131 ,
		_w577_,
		_w584_,
		_w925_,
		_w926_
	);
	LUT2 #(
		.INIT('h8)
	) name464 (
		_w924_,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h7)
	) name465 (
		_w924_,
		_w926_,
		_w928_
	);
	LUT3 #(
		.INIT('h45)
	) name466 (
		_w494_,
		_w606_,
		_w607_,
		_w929_
	);
	LUT4 #(
		.INIT('h5659)
	) name467 (
		\P2_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w568_,
		_w929_,
		_w930_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name468 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_IR_reg[5]/NET0131 ,
		_w466_,
		_w931_
	);
	LUT2 #(
		.INIT('h6)
	) name469 (
		\P1_IR_reg[6]/NET0131 ,
		_w931_,
		_w932_
	);
	LUT4 #(
		.INIT('hd0f2)
	) name470 (
		_w479_,
		_w488_,
		_w930_,
		_w932_,
		_w933_
	);
	LUT3 #(
		.INIT('h08)
	) name471 (
		_w924_,
		_w926_,
		_w933_,
		_w934_
	);
	LUT4 #(
		.INIT('hff35)
	) name472 (
		\P1_reg0_reg[7]/NET0131 ,
		\P1_reg2_reg[7]/NET0131 ,
		_w577_,
		_w584_,
		_w935_
	);
	LUT2 #(
		.INIT('h6)
	) name473 (
		\P1_reg3_reg[7]/NET0131 ,
		_w586_,
		_w936_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name474 (
		\P1_reg1_reg[7]/NET0131 ,
		_w577_,
		_w584_,
		_w936_,
		_w937_
	);
	LUT2 #(
		.INIT('h8)
	) name475 (
		_w935_,
		_w937_,
		_w938_
	);
	LUT2 #(
		.INIT('h7)
	) name476 (
		_w935_,
		_w937_,
		_w939_
	);
	LUT4 #(
		.INIT('h5956)
	) name477 (
		\P2_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w568_,
		_w504_,
		_w940_
	);
	LUT2 #(
		.INIT('h8)
	) name478 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[6]/NET0131 ,
		_w941_
	);
	LUT3 #(
		.INIT('h56)
	) name479 (
		\P1_IR_reg[7]/NET0131 ,
		_w931_,
		_w941_,
		_w942_
	);
	LUT4 #(
		.INIT('hd0f2)
	) name480 (
		_w479_,
		_w488_,
		_w940_,
		_w942_,
		_w943_
	);
	LUT3 #(
		.INIT('h08)
	) name481 (
		_w935_,
		_w937_,
		_w943_,
		_w944_
	);
	LUT2 #(
		.INIT('h1)
	) name482 (
		_w934_,
		_w944_,
		_w945_
	);
	LUT4 #(
		.INIT('hff35)
	) name483 (
		\P1_reg0_reg[5]/NET0131 ,
		\P1_reg2_reg[5]/NET0131 ,
		_w577_,
		_w584_,
		_w946_
	);
	LUT3 #(
		.INIT('h78)
	) name484 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		\P1_reg3_reg[5]/NET0131 ,
		_w947_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name485 (
		\P1_reg1_reg[5]/NET0131 ,
		_w577_,
		_w584_,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h8)
	) name486 (
		_w946_,
		_w948_,
		_w949_
	);
	LUT2 #(
		.INIT('h7)
	) name487 (
		_w946_,
		_w948_,
		_w950_
	);
	LUT2 #(
		.INIT('h8)
	) name488 (
		\P2_datao_reg[5]/NET0131 ,
		_w568_,
		_w951_
	);
	LUT2 #(
		.INIT('h6)
	) name489 (
		\P2_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w952_
	);
	LUT4 #(
		.INIT('h0154)
	) name490 (
		_w568_,
		_w501_,
		_w606_,
		_w952_,
		_w953_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		_w951_,
		_w953_,
		_w954_
	);
	LUT4 #(
		.INIT('h87a5)
	) name492 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_IR_reg[5]/NET0131 ,
		_w466_,
		_w955_
	);
	LUT4 #(
		.INIT('hf2d0)
	) name493 (
		_w479_,
		_w488_,
		_w954_,
		_w955_,
		_w956_
	);
	LUT3 #(
		.INIT('h08)
	) name494 (
		_w946_,
		_w948_,
		_w956_,
		_w957_
	);
	LUT2 #(
		.INIT('h6)
	) name495 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		_w958_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name496 (
		\P1_reg1_reg[4]/NET0131 ,
		_w577_,
		_w584_,
		_w958_,
		_w959_
	);
	LUT4 #(
		.INIT('hff35)
	) name497 (
		\P1_reg0_reg[4]/NET0131 ,
		\P1_reg2_reg[4]/NET0131 ,
		_w577_,
		_w584_,
		_w960_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		_w959_,
		_w960_,
		_w961_
	);
	LUT2 #(
		.INIT('h7)
	) name499 (
		_w959_,
		_w960_,
		_w962_
	);
	LUT3 #(
		.INIT('hc6)
	) name500 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		_w466_,
		_w963_
	);
	LUT4 #(
		.INIT('h040f)
	) name501 (
		_w490_,
		_w492_,
		_w497_,
		_w605_,
		_w964_
	);
	LUT4 #(
		.INIT('ha9a6)
	) name502 (
		\P2_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w568_,
		_w964_,
		_w965_
	);
	LUT4 #(
		.INIT('h02df)
	) name503 (
		_w479_,
		_w488_,
		_w963_,
		_w965_,
		_w966_
	);
	LUT3 #(
		.INIT('h08)
	) name504 (
		_w959_,
		_w960_,
		_w966_,
		_w967_
	);
	LUT2 #(
		.INIT('h1)
	) name505 (
		_w957_,
		_w967_,
		_w968_
	);
	LUT4 #(
		.INIT('hcff5)
	) name506 (
		\P1_reg0_reg[3]/NET0131 ,
		\P1_reg3_reg[3]/NET0131 ,
		_w577_,
		_w584_,
		_w969_
	);
	LUT4 #(
		.INIT('hf53f)
	) name507 (
		\P1_reg1_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w577_,
		_w584_,
		_w970_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		_w969_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h7)
	) name509 (
		_w969_,
		_w970_,
		_w972_
	);
	LUT4 #(
		.INIT('h5956)
	) name510 (
		\P2_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w568_,
		_w493_,
		_w973_
	);
	LUT4 #(
		.INIT('hfe00)
	) name511 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[2]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w974_
	);
	LUT2 #(
		.INIT('h6)
	) name512 (
		\P1_IR_reg[3]/NET0131 ,
		_w974_,
		_w975_
	);
	LUT4 #(
		.INIT('hd0f2)
	) name513 (
		_w479_,
		_w488_,
		_w973_,
		_w975_,
		_w976_
	);
	LUT3 #(
		.INIT('h08)
	) name514 (
		_w969_,
		_w970_,
		_w976_,
		_w977_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name515 (
		\P1_reg0_reg[2]/NET0131 ,
		\P1_reg1_reg[2]/NET0131 ,
		_w577_,
		_w584_,
		_w978_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name516 (
		\P1_reg2_reg[2]/NET0131 ,
		\P1_reg3_reg[2]/NET0131 ,
		_w577_,
		_w584_,
		_w979_
	);
	LUT2 #(
		.INIT('h8)
	) name517 (
		_w978_,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h7)
	) name518 (
		_w978_,
		_w979_,
		_w981_
	);
	LUT4 #(
		.INIT('h5659)
	) name519 (
		\P2_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w568_,
		_w492_,
		_w982_
	);
	LUT4 #(
		.INIT('h1ef0)
	) name520 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[2]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w983_
	);
	LUT4 #(
		.INIT('hd0f2)
	) name521 (
		_w479_,
		_w488_,
		_w982_,
		_w983_,
		_w984_
	);
	LUT3 #(
		.INIT('h08)
	) name522 (
		_w978_,
		_w979_,
		_w984_,
		_w985_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		_w977_,
		_w985_,
		_w986_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name524 (
		\P1_reg2_reg[1]/NET0131 ,
		\P1_reg3_reg[1]/NET0131 ,
		_w577_,
		_w584_,
		_w987_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name525 (
		\P1_reg0_reg[1]/NET0131 ,
		\P1_reg1_reg[1]/NET0131 ,
		_w577_,
		_w584_,
		_w988_
	);
	LUT2 #(
		.INIT('h8)
	) name526 (
		_w987_,
		_w988_,
		_w989_
	);
	LUT2 #(
		.INIT('h7)
	) name527 (
		_w987_,
		_w988_,
		_w990_
	);
	LUT3 #(
		.INIT('h93)
	) name528 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w991_
	);
	LUT4 #(
		.INIT('ha9a6)
	) name529 (
		\P2_datao_reg[1]/NET0131 ,
		\si[1]_pad ,
		_w568_,
		_w491_,
		_w992_
	);
	LUT4 #(
		.INIT('h20fd)
	) name530 (
		_w479_,
		_w488_,
		_w991_,
		_w992_,
		_w993_
	);
	LUT3 #(
		.INIT('h70)
	) name531 (
		_w987_,
		_w988_,
		_w993_,
		_w994_
	);
	LUT3 #(
		.INIT('h08)
	) name532 (
		_w987_,
		_w988_,
		_w993_,
		_w995_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name533 (
		\P1_reg0_reg[0]/NET0131 ,
		\P1_reg1_reg[0]/NET0131 ,
		_w577_,
		_w584_,
		_w996_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name534 (
		\P1_reg2_reg[0]/NET0131 ,
		\P1_reg3_reg[0]/NET0131 ,
		_w577_,
		_w584_,
		_w997_
	);
	LUT2 #(
		.INIT('h8)
	) name535 (
		_w996_,
		_w997_,
		_w998_
	);
	LUT2 #(
		.INIT('h7)
	) name536 (
		_w996_,
		_w997_,
		_w999_
	);
	LUT3 #(
		.INIT('ha6)
	) name537 (
		\P2_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w568_,
		_w1000_
	);
	LUT4 #(
		.INIT('h04f7)
	) name538 (
		\P1_IR_reg[0]/NET0131 ,
		_w479_,
		_w488_,
		_w1000_,
		_w1001_
	);
	LUT3 #(
		.INIT('h08)
	) name539 (
		_w996_,
		_w997_,
		_w1001_,
		_w1002_
	);
	LUT3 #(
		.INIT('h54)
	) name540 (
		_w994_,
		_w995_,
		_w1002_,
		_w1003_
	);
	LUT3 #(
		.INIT('h70)
	) name541 (
		_w969_,
		_w970_,
		_w976_,
		_w1004_
	);
	LUT3 #(
		.INIT('h70)
	) name542 (
		_w978_,
		_w979_,
		_w984_,
		_w1005_
	);
	LUT3 #(
		.INIT('h23)
	) name543 (
		_w977_,
		_w1004_,
		_w1005_,
		_w1006_
	);
	LUT4 #(
		.INIT('h08aa)
	) name544 (
		_w968_,
		_w986_,
		_w1003_,
		_w1006_,
		_w1007_
	);
	LUT3 #(
		.INIT('h70)
	) name545 (
		_w946_,
		_w948_,
		_w956_,
		_w1008_
	);
	LUT3 #(
		.INIT('h70)
	) name546 (
		_w959_,
		_w960_,
		_w966_,
		_w1009_
	);
	LUT3 #(
		.INIT('h23)
	) name547 (
		_w957_,
		_w1008_,
		_w1009_,
		_w1010_
	);
	LUT3 #(
		.INIT('h70)
	) name548 (
		_w935_,
		_w937_,
		_w943_,
		_w1011_
	);
	LUT3 #(
		.INIT('h70)
	) name549 (
		_w924_,
		_w926_,
		_w933_,
		_w1012_
	);
	LUT3 #(
		.INIT('h54)
	) name550 (
		_w944_,
		_w1011_,
		_w1012_,
		_w1013_
	);
	LUT3 #(
		.INIT('h0d)
	) name551 (
		_w945_,
		_w1010_,
		_w1013_,
		_w1014_
	);
	LUT3 #(
		.INIT('h70)
	) name552 (
		_w945_,
		_w1007_,
		_w1014_,
		_w1015_
	);
	LUT3 #(
		.INIT('h08)
	) name553 (
		_w909_,
		_w910_,
		_w915_,
		_w1016_
	);
	LUT2 #(
		.INIT('h1)
	) name554 (
		_w906_,
		_w1016_,
		_w1017_
	);
	LUT4 #(
		.INIT('h0001)
	) name555 (
		_w885_,
		_w894_,
		_w906_,
		_w1016_,
		_w1018_
	);
	LUT4 #(
		.INIT('h8f00)
	) name556 (
		_w945_,
		_w1007_,
		_w1014_,
		_w1018_,
		_w1019_
	);
	LUT3 #(
		.INIT('h4c)
	) name557 (
		_w872_,
		_w923_,
		_w1019_,
		_w1020_
	);
	LUT4 #(
		.INIT('h0001)
	) name558 (
		_w782_,
		_w791_,
		_w802_,
		_w818_,
		_w1021_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name559 (
		_w749_,
		_w754_,
		_w759_,
		_w764_,
		_w1022_
	);
	LUT3 #(
		.INIT('h10)
	) name560 (
		_w726_,
		_w741_,
		_w1022_,
		_w1023_
	);
	LUT2 #(
		.INIT('h8)
	) name561 (
		_w1021_,
		_w1023_,
		_w1024_
	);
	LUT4 #(
		.INIT('hb300)
	) name562 (
		_w872_,
		_w923_,
		_w1019_,
		_w1024_,
		_w1025_
	);
	LUT3 #(
		.INIT('h40)
	) name563 (
		_w612_,
		_w614_,
		_w625_,
		_w1026_
	);
	LUT4 #(
		.INIT('h7500)
	) name564 (
		_w632_,
		_w617_,
		_w621_,
		_w624_,
		_w1027_
	);
	LUT2 #(
		.INIT('h2)
	) name565 (
		_w629_,
		_w1027_,
		_w1028_
	);
	LUT4 #(
		.INIT('h2a22)
	) name566 (
		_w640_,
		_w635_,
		_w1026_,
		_w1028_,
		_w1029_
	);
	LUT4 #(
		.INIT('h5956)
	) name567 (
		\P2_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w568_,
		_w1029_,
		_w1030_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		_w489_,
		_w1030_,
		_w1031_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name569 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_reg3_reg[26]/NET0131 ,
		_w593_,
		_w596_,
		_w1032_
	);
	LUT3 #(
		.INIT('h20)
	) name570 (
		\P1_reg1_reg[26]/NET0131 ,
		_w577_,
		_w584_,
		_w1033_
	);
	LUT4 #(
		.INIT('hff35)
	) name571 (
		\P1_reg0_reg[26]/NET0131 ,
		\P1_reg2_reg[26]/NET0131 ,
		_w577_,
		_w584_,
		_w1034_
	);
	LUT4 #(
		.INIT('h1300)
	) name572 (
		_w585_,
		_w1033_,
		_w1032_,
		_w1034_,
		_w1035_
	);
	LUT4 #(
		.INIT('hecff)
	) name573 (
		_w585_,
		_w1033_,
		_w1032_,
		_w1034_,
		_w1036_
	);
	LUT3 #(
		.INIT('h10)
	) name574 (
		_w489_,
		_w1030_,
		_w1035_,
		_w1037_
	);
	LUT4 #(
		.INIT('h4f00)
	) name575 (
		_w529_,
		_w533_,
		_w542_,
		_w536_,
		_w1038_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name576 (
		_w539_,
		_w560_,
		_w550_,
		_w1038_,
		_w1039_
	);
	LUT4 #(
		.INIT('h5956)
	) name577 (
		\P2_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w568_,
		_w1039_,
		_w1040_
	);
	LUT2 #(
		.INIT('h1)
	) name578 (
		_w489_,
		_w1040_,
		_w1041_
	);
	LUT2 #(
		.INIT('h6)
	) name579 (
		\P1_reg3_reg[27]/NET0131 ,
		_w703_,
		_w1042_
	);
	LUT3 #(
		.INIT('h48)
	) name580 (
		\P1_reg3_reg[27]/NET0131 ,
		_w585_,
		_w703_,
		_w1043_
	);
	LUT3 #(
		.INIT('h08)
	) name581 (
		\P1_reg2_reg[27]/NET0131 ,
		_w577_,
		_w584_,
		_w1044_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name582 (
		\P1_reg0_reg[27]/NET0131 ,
		\P1_reg1_reg[27]/NET0131 ,
		_w577_,
		_w584_,
		_w1045_
	);
	LUT2 #(
		.INIT('h4)
	) name583 (
		_w1044_,
		_w1045_,
		_w1046_
	);
	LUT2 #(
		.INIT('h4)
	) name584 (
		_w1043_,
		_w1046_,
		_w1047_
	);
	LUT2 #(
		.INIT('hb)
	) name585 (
		_w1043_,
		_w1046_,
		_w1048_
	);
	LUT3 #(
		.INIT('h10)
	) name586 (
		_w489_,
		_w1040_,
		_w1047_,
		_w1049_
	);
	LUT4 #(
		.INIT('h3233)
	) name587 (
		_w489_,
		_w1037_,
		_w1040_,
		_w1047_,
		_w1050_
	);
	LUT4 #(
		.INIT('h020f)
	) name588 (
		_w537_,
		_w545_,
		_w547_,
		_w559_,
		_w1051_
	);
	LUT3 #(
		.INIT('h40)
	) name589 (
		_w660_,
		_w661_,
		_w665_,
		_w1052_
	);
	LUT4 #(
		.INIT('h7500)
	) name590 (
		_w668_,
		_w657_,
		_w663_,
		_w664_,
		_w1053_
	);
	LUT2 #(
		.INIT('h2)
	) name591 (
		_w667_,
		_w1053_,
		_w1054_
	);
	LUT4 #(
		.INIT('hfac8)
	) name592 (
		\P2_datao_reg[23]/NET0131 ,
		\P2_datao_reg[24]/NET0131 ,
		\si[23]_pad ,
		\si[24]_pad ,
		_w1055_
	);
	LUT2 #(
		.INIT('h8)
	) name593 (
		_w534_,
		_w1055_,
		_w1056_
	);
	LUT4 #(
		.INIT('h1055)
	) name594 (
		_w1051_,
		_w1052_,
		_w1054_,
		_w1056_,
		_w1057_
	);
	LUT4 #(
		.INIT('h5956)
	) name595 (
		\P2_datao_reg[25]/NET0131 ,
		\si[25]_pad ,
		_w568_,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		_w489_,
		_w1058_,
		_w1059_
	);
	LUT3 #(
		.INIT('h6a)
	) name597 (
		\P1_reg3_reg[25]/NET0131 ,
		_w593_,
		_w596_,
		_w1060_
	);
	LUT3 #(
		.INIT('h08)
	) name598 (
		\P1_reg2_reg[25]/NET0131 ,
		_w577_,
		_w584_,
		_w1061_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name599 (
		\P1_reg0_reg[25]/NET0131 ,
		\P1_reg1_reg[25]/NET0131 ,
		_w577_,
		_w584_,
		_w1062_
	);
	LUT4 #(
		.INIT('h1300)
	) name600 (
		_w585_,
		_w1061_,
		_w1060_,
		_w1062_,
		_w1063_
	);
	LUT4 #(
		.INIT('hecff)
	) name601 (
		_w585_,
		_w1061_,
		_w1060_,
		_w1062_,
		_w1064_
	);
	LUT3 #(
		.INIT('h10)
	) name602 (
		_w489_,
		_w1058_,
		_w1063_,
		_w1065_
	);
	LUT2 #(
		.INIT('h8)
	) name603 (
		\P2_datao_reg[24]/NET0131 ,
		_w568_,
		_w1066_
	);
	LUT2 #(
		.INIT('h6)
	) name604 (
		\P2_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w1067_
	);
	LUT4 #(
		.INIT('h8000)
	) name605 (
		_w619_,
		_w622_,
		_w623_,
		_w634_,
		_w1068_
	);
	LUT4 #(
		.INIT('h8000)
	) name606 (
		_w683_,
		_w685_,
		_w686_,
		_w1068_,
		_w1069_
	);
	LUT4 #(
		.INIT('h2f00)
	) name607 (
		_w683_,
		_w688_,
		_w689_,
		_w692_,
		_w1070_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name608 (
		_w682_,
		_w698_,
		_w694_,
		_w1070_,
		_w1071_
	);
	LUT4 #(
		.INIT('h1411)
	) name609 (
		_w568_,
		_w1067_,
		_w1069_,
		_w1071_,
		_w1072_
	);
	LUT3 #(
		.INIT('h54)
	) name610 (
		_w489_,
		_w1066_,
		_w1072_,
		_w1073_
	);
	LUT3 #(
		.INIT('h0e)
	) name611 (
		\P1_reg3_reg[24]/NET0131 ,
		_w785_,
		_w597_,
		_w1074_
	);
	LUT4 #(
		.INIT('h00c8)
	) name612 (
		\P1_reg3_reg[24]/NET0131 ,
		_w585_,
		_w785_,
		_w597_,
		_w1075_
	);
	LUT3 #(
		.INIT('h02)
	) name613 (
		\P1_reg0_reg[24]/NET0131 ,
		_w577_,
		_w584_,
		_w1076_
	);
	LUT4 #(
		.INIT('hf53f)
	) name614 (
		\P1_reg1_reg[24]/NET0131 ,
		\P1_reg2_reg[24]/NET0131 ,
		_w577_,
		_w584_,
		_w1077_
	);
	LUT2 #(
		.INIT('h4)
	) name615 (
		_w1076_,
		_w1077_,
		_w1078_
	);
	LUT2 #(
		.INIT('h4)
	) name616 (
		_w1075_,
		_w1078_,
		_w1079_
	);
	LUT2 #(
		.INIT('hb)
	) name617 (
		_w1075_,
		_w1078_,
		_w1080_
	);
	LUT3 #(
		.INIT('h20)
	) name618 (
		_w1073_,
		_w1075_,
		_w1078_,
		_w1081_
	);
	LUT2 #(
		.INIT('h1)
	) name619 (
		_w1065_,
		_w1081_,
		_w1082_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		_w1050_,
		_w1082_,
		_w1083_
	);
	LUT3 #(
		.INIT('h0e)
	) name621 (
		_w489_,
		_w1040_,
		_w1047_,
		_w1084_
	);
	LUT3 #(
		.INIT('h0e)
	) name622 (
		_w489_,
		_w1030_,
		_w1035_,
		_w1085_
	);
	LUT3 #(
		.INIT('h0e)
	) name623 (
		_w489_,
		_w1058_,
		_w1063_,
		_w1086_
	);
	LUT3 #(
		.INIT('h45)
	) name624 (
		_w1073_,
		_w1075_,
		_w1078_,
		_w1087_
	);
	LUT3 #(
		.INIT('h23)
	) name625 (
		_w1065_,
		_w1086_,
		_w1087_,
		_w1088_
	);
	LUT4 #(
		.INIT('h080e)
	) name626 (
		_w1059_,
		_w1063_,
		_w1085_,
		_w1087_,
		_w1089_
	);
	LUT3 #(
		.INIT('h31)
	) name627 (
		_w1050_,
		_w1084_,
		_w1089_,
		_w1090_
	);
	LUT4 #(
		.INIT('h1f00)
	) name628 (
		_w823_,
		_w1025_,
		_w1083_,
		_w1090_,
		_w1091_
	);
	LUT2 #(
		.INIT('h8)
	) name629 (
		_w702_,
		_w708_,
		_w1092_
	);
	LUT3 #(
		.INIT('h15)
	) name630 (
		_w679_,
		_w702_,
		_w708_,
		_w1093_
	);
	LUT4 #(
		.INIT('hbf00)
	) name631 (
		_w1091_,
		_w1093_,
		_w653_,
		_w715_,
		_w1094_
	);
	LUT2 #(
		.INIT('h2)
	) name632 (
		\P1_IR_reg[31]/NET0131 ,
		_w578_,
		_w1095_
	);
	LUT3 #(
		.INIT('h56)
	) name633 (
		\P1_IR_reg[21]/NET0131 ,
		_w746_,
		_w1095_,
		_w1096_
	);
	LUT3 #(
		.INIT('h2a)
	) name634 (
		\P1_IR_reg[31]/NET0131 ,
		_w483_,
		_w475_,
		_w1097_
	);
	LUT3 #(
		.INIT('h56)
	) name635 (
		\P1_IR_reg[22]/NET0131 ,
		_w482_,
		_w1097_,
		_w1098_
	);
	LUT2 #(
		.INIT('h2)
	) name636 (
		\P1_IR_reg[31]/NET0131 ,
		_w483_,
		_w1099_
	);
	LUT3 #(
		.INIT('h56)
	) name637 (
		\P1_IR_reg[20]/NET0131 ,
		_w482_,
		_w1099_,
		_w1100_
	);
	LUT4 #(
		.INIT('h00a9)
	) name638 (
		\P1_IR_reg[20]/NET0131 ,
		_w482_,
		_w1099_,
		_w718_,
		_w1101_
	);
	LUT3 #(
		.INIT('h40)
	) name639 (
		_w1096_,
		_w1098_,
		_w1101_,
		_w1102_
	);
	LUT3 #(
		.INIT('hb0)
	) name640 (
		\P1_B_reg/NET0131 ,
		_w1094_,
		_w1102_,
		_w1103_
	);
	LUT4 #(
		.INIT('h0504)
	) name641 (
		_w489_,
		_w602_,
		_w646_,
		_w650_,
		_w1104_
	);
	LUT4 #(
		.INIT('h00f4)
	) name642 (
		_w489_,
		_w569_,
		_w602_,
		_w1104_,
		_w1105_
	);
	LUT4 #(
		.INIT('h3301)
	) name643 (
		_w489_,
		_w602_,
		_w646_,
		_w650_,
		_w1106_
	);
	LUT3 #(
		.INIT('h04)
	) name644 (
		_w489_,
		_w569_,
		_w1106_,
		_w1107_
	);
	LUT4 #(
		.INIT('heee8)
	) name645 (
		_w674_,
		_w677_,
		_w702_,
		_w708_,
		_w1108_
	);
	LUT3 #(
		.INIT('h31)
	) name646 (
		_w1105_,
		_w1107_,
		_w1108_,
		_w1109_
	);
	LUT4 #(
		.INIT('hbf00)
	) name647 (
		_w1091_,
		_w1093_,
		_w1105_,
		_w1109_,
		_w1110_
	);
	LUT4 #(
		.INIT('h0056)
	) name648 (
		\P1_IR_reg[22]/NET0131 ,
		_w482_,
		_w1097_,
		_w718_,
		_w1111_
	);
	LUT3 #(
		.INIT('h80)
	) name649 (
		_w1096_,
		_w1100_,
		_w1111_,
		_w1112_
	);
	LUT4 #(
		.INIT('h5600)
	) name650 (
		\P1_IR_reg[22]/NET0131 ,
		_w482_,
		_w1097_,
		_w718_,
		_w1113_
	);
	LUT3 #(
		.INIT('h80)
	) name651 (
		_w1096_,
		_w1100_,
		_w1113_,
		_w1114_
	);
	LUT4 #(
		.INIT('h014f)
	) name652 (
		\P1_B_reg/NET0131 ,
		_w1110_,
		_w1112_,
		_w1114_,
		_w1115_
	);
	LUT2 #(
		.INIT('h4)
	) name653 (
		_w1103_,
		_w1115_,
		_w1116_
	);
	LUT3 #(
		.INIT('h08)
	) name654 (
		_w1096_,
		_w1100_,
		_w1098_,
		_w1117_
	);
	LUT3 #(
		.INIT('h90)
	) name655 (
		_w718_,
		_w1110_,
		_w1117_,
		_w1118_
	);
	LUT2 #(
		.INIT('h1)
	) name656 (
		_w1096_,
		_w1098_,
		_w1119_
	);
	LUT3 #(
		.INIT('h10)
	) name657 (
		_w1096_,
		_w1098_,
		_w1101_,
		_w1120_
	);
	LUT2 #(
		.INIT('h4)
	) name658 (
		_w1094_,
		_w1120_,
		_w1121_
	);
	LUT4 #(
		.INIT('ha900)
	) name659 (
		\P1_IR_reg[20]/NET0131 ,
		_w482_,
		_w1099_,
		_w718_,
		_w1122_
	);
	LUT2 #(
		.INIT('h4)
	) name660 (
		_w1096_,
		_w1122_,
		_w1123_
	);
	LUT2 #(
		.INIT('h8)
	) name661 (
		_w1094_,
		_w1123_,
		_w1124_
	);
	LUT4 #(
		.INIT('h1303)
	) name662 (
		_w1093_,
		_w604_,
		_w653_,
		_w714_,
		_w1125_
	);
	LUT4 #(
		.INIT('h00e8)
	) name663 (
		_w1059_,
		_w1063_,
		_w1081_,
		_w1085_,
		_w1126_
	);
	LUT3 #(
		.INIT('h31)
	) name664 (
		_w1050_,
		_w1084_,
		_w1126_,
		_w1127_
	);
	LUT3 #(
		.INIT('ha8)
	) name665 (
		_w715_,
		_w1125_,
		_w1127_,
		_w1128_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name666 (
		_w734_,
		_w739_,
		_w749_,
		_w754_,
		_w1129_
	);
	LUT4 #(
		.INIT('h1011)
	) name667 (
		_w726_,
		_w741_,
		_w1022_,
		_w1129_,
		_w1130_
	);
	LUT2 #(
		.INIT('h1)
	) name668 (
		_w770_,
		_w1130_,
		_w1131_
	);
	LUT3 #(
		.INIT('ha8)
	) name669 (
		_w817_,
		_w822_,
		_w1131_,
		_w1132_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name670 (
		_w837_,
		_w842_,
		_w847_,
		_w852_,
		_w1133_
	);
	LUT4 #(
		.INIT('h1311)
	) name671 (
		_w843_,
		_w867_,
		_w871_,
		_w1133_,
		_w1134_
	);
	LUT4 #(
		.INIT('h0b02)
	) name672 (
		_w899_,
		_w905_,
		_w918_,
		_w1016_,
		_w1135_
	);
	LUT3 #(
		.INIT('h31)
	) name673 (
		_w895_,
		_w919_,
		_w1135_,
		_w1136_
	);
	LUT3 #(
		.INIT('ha8)
	) name674 (
		_w870_,
		_w1134_,
		_w1136_,
		_w1137_
	);
	LUT3 #(
		.INIT('h70)
	) name675 (
		_w996_,
		_w997_,
		_w1001_,
		_w1138_
	);
	LUT4 #(
		.INIT('h020b)
	) name676 (
		_w989_,
		_w993_,
		_w1005_,
		_w1138_,
		_w1139_
	);
	LUT4 #(
		.INIT('h0001)
	) name677 (
		_w1004_,
		_w1008_,
		_w1009_,
		_w1012_,
		_w1140_
	);
	LUT3 #(
		.INIT('hd0)
	) name678 (
		_w986_,
		_w1139_,
		_w1140_,
		_w1141_
	);
	LUT4 #(
		.INIT('h00b2)
	) name679 (
		_w949_,
		_w956_,
		_w967_,
		_w1012_,
		_w1142_
	);
	LUT2 #(
		.INIT('h2)
	) name680 (
		_w945_,
		_w1142_,
		_w1143_
	);
	LUT3 #(
		.INIT('h01)
	) name681 (
		_w907_,
		_w916_,
		_w1011_,
		_w1144_
	);
	LUT4 #(
		.INIT('h8000)
	) name682 (
		_w865_,
		_w868_,
		_w920_,
		_w1144_,
		_w1145_
	);
	LUT3 #(
		.INIT('hb0)
	) name683 (
		_w1141_,
		_w1143_,
		_w1145_,
		_w1146_
	);
	LUT3 #(
		.INIT('h02)
	) name684 (
		_w766_,
		_w769_,
		_w770_,
		_w1147_
	);
	LUT4 #(
		.INIT('h0001)
	) name685 (
		_w803_,
		_w812_,
		_w814_,
		_w815_,
		_w1148_
	);
	LUT2 #(
		.INIT('h8)
	) name686 (
		_w1147_,
		_w1148_,
		_w1149_
	);
	LUT3 #(
		.INIT('he0)
	) name687 (
		_w1137_,
		_w1146_,
		_w1149_,
		_w1150_
	);
	LUT3 #(
		.INIT('h01)
	) name688 (
		_w1085_,
		_w1086_,
		_w1087_,
		_w1151_
	);
	LUT3 #(
		.INIT('h40)
	) name689 (
		_w710_,
		_w714_,
		_w1151_,
		_w1152_
	);
	LUT2 #(
		.INIT('h1)
	) name690 (
		_w1084_,
		_w604_,
		_w1153_
	);
	LUT2 #(
		.INIT('h8)
	) name691 (
		_w1152_,
		_w1153_,
		_w1154_
	);
	LUT4 #(
		.INIT('h0155)
	) name692 (
		_w1128_,
		_w1132_,
		_w1150_,
		_w1154_,
		_w1155_
	);
	LUT3 #(
		.INIT('h02)
	) name693 (
		_w1096_,
		_w1100_,
		_w1098_,
		_w1156_
	);
	LUT3 #(
		.INIT('h60)
	) name694 (
		_w718_,
		_w1155_,
		_w1156_,
		_w1157_
	);
	LUT2 #(
		.INIT('h4)
	) name695 (
		_w702_,
		_w708_,
		_w1158_
	);
	LUT2 #(
		.INIT('h2)
	) name696 (
		_w702_,
		_w708_,
		_w1159_
	);
	LUT2 #(
		.INIT('h9)
	) name697 (
		_w702_,
		_w708_,
		_w1160_
	);
	LUT3 #(
		.INIT('hb4)
	) name698 (
		_w489_,
		_w569_,
		_w602_,
		_w1161_
	);
	LUT2 #(
		.INIT('h4)
	) name699 (
		_w1160_,
		_w1161_,
		_w1162_
	);
	LUT3 #(
		.INIT('h01)
	) name700 (
		_w489_,
		_w1040_,
		_w1047_,
		_w1163_
	);
	LUT3 #(
		.INIT('he0)
	) name701 (
		_w489_,
		_w1040_,
		_w1047_,
		_w1164_
	);
	LUT3 #(
		.INIT('h1e)
	) name702 (
		_w489_,
		_w1040_,
		_w1047_,
		_w1165_
	);
	LUT2 #(
		.INIT('h9)
	) name703 (
		_w847_,
		_w852_,
		_w1166_
	);
	LUT2 #(
		.INIT('h6)
	) name704 (
		_w856_,
		_w864_,
		_w1167_
	);
	LUT2 #(
		.INIT('h6)
	) name705 (
		_w827_,
		_w833_,
		_w1168_
	);
	LUT4 #(
		.INIT('h9009)
	) name706 (
		_w827_,
		_w833_,
		_w856_,
		_w864_,
		_w1169_
	);
	LUT2 #(
		.INIT('h8)
	) name707 (
		_w1166_,
		_w1169_,
		_w1170_
	);
	LUT3 #(
		.INIT('h80)
	) name708 (
		_w896_,
		_w898_,
		_w905_,
		_w1171_
	);
	LUT3 #(
		.INIT('h07)
	) name709 (
		_w896_,
		_w898_,
		_w905_,
		_w1172_
	);
	LUT3 #(
		.INIT('h78)
	) name710 (
		_w896_,
		_w898_,
		_w905_,
		_w1173_
	);
	LUT4 #(
		.INIT('h7778)
	) name711 (
		_w873_,
		_w875_,
		_w881_,
		_w883_,
		_w1174_
	);
	LUT3 #(
		.INIT('h07)
	) name712 (
		_w959_,
		_w960_,
		_w966_,
		_w1175_
	);
	LUT3 #(
		.INIT('h80)
	) name713 (
		_w959_,
		_w960_,
		_w966_,
		_w1176_
	);
	LUT3 #(
		.INIT('h78)
	) name714 (
		_w959_,
		_w960_,
		_w966_,
		_w1177_
	);
	LUT3 #(
		.INIT('h87)
	) name715 (
		_w887_,
		_w888_,
		_w893_,
		_w1178_
	);
	LUT4 #(
		.INIT('h0400)
	) name716 (
		_w1173_,
		_w1174_,
		_w1177_,
		_w1178_,
		_w1179_
	);
	LUT3 #(
		.INIT('h87)
	) name717 (
		_w996_,
		_w997_,
		_w1001_,
		_w1180_
	);
	LUT3 #(
		.INIT('h87)
	) name718 (
		_w924_,
		_w926_,
		_w933_,
		_w1181_
	);
	LUT3 #(
		.INIT('h80)
	) name719 (
		_w935_,
		_w937_,
		_w943_,
		_w1182_
	);
	LUT3 #(
		.INIT('h07)
	) name720 (
		_w935_,
		_w937_,
		_w943_,
		_w1183_
	);
	LUT3 #(
		.INIT('h78)
	) name721 (
		_w935_,
		_w937_,
		_w943_,
		_w1184_
	);
	LUT3 #(
		.INIT('h80)
	) name722 (
		_w969_,
		_w970_,
		_w976_,
		_w1185_
	);
	LUT3 #(
		.INIT('h07)
	) name723 (
		_w969_,
		_w970_,
		_w976_,
		_w1186_
	);
	LUT3 #(
		.INIT('h78)
	) name724 (
		_w969_,
		_w970_,
		_w976_,
		_w1187_
	);
	LUT4 #(
		.INIT('h0008)
	) name725 (
		_w1180_,
		_w1181_,
		_w1184_,
		_w1187_,
		_w1188_
	);
	LUT2 #(
		.INIT('h9)
	) name726 (
		_w837_,
		_w842_,
		_w1189_
	);
	LUT3 #(
		.INIT('h87)
	) name727 (
		_w987_,
		_w988_,
		_w993_,
		_w1190_
	);
	LUT3 #(
		.INIT('h87)
	) name728 (
		_w909_,
		_w910_,
		_w915_,
		_w1191_
	);
	LUT3 #(
		.INIT('h87)
	) name729 (
		_w946_,
		_w948_,
		_w956_,
		_w1192_
	);
	LUT3 #(
		.INIT('h87)
	) name730 (
		_w978_,
		_w979_,
		_w984_,
		_w1193_
	);
	LUT4 #(
		.INIT('h8000)
	) name731 (
		_w1190_,
		_w1191_,
		_w1192_,
		_w1193_,
		_w1194_
	);
	LUT4 #(
		.INIT('h8000)
	) name732 (
		_w1189_,
		_w1194_,
		_w1179_,
		_w1188_,
		_w1195_
	);
	LUT3 #(
		.INIT('he1)
	) name733 (
		_w489_,
		_w646_,
		_w650_,
		_w1196_
	);
	LUT3 #(
		.INIT('he1)
	) name734 (
		_w489_,
		_w673_,
		_w677_,
		_w1197_
	);
	LUT2 #(
		.INIT('h9)
	) name735 (
		_w759_,
		_w764_,
		_w1198_
	);
	LUT2 #(
		.INIT('h4)
	) name736 (
		_w776_,
		_w780_,
		_w1199_
	);
	LUT2 #(
		.INIT('h2)
	) name737 (
		_w776_,
		_w780_,
		_w1200_
	);
	LUT2 #(
		.INIT('h9)
	) name738 (
		_w776_,
		_w780_,
		_w1201_
	);
	LUT2 #(
		.INIT('h4)
	) name739 (
		_w796_,
		_w800_,
		_w1202_
	);
	LUT2 #(
		.INIT('h2)
	) name740 (
		_w796_,
		_w800_,
		_w1203_
	);
	LUT2 #(
		.INIT('h9)
	) name741 (
		_w796_,
		_w800_,
		_w1204_
	);
	LUT4 #(
		.INIT('h0660)
	) name742 (
		_w776_,
		_w780_,
		_w796_,
		_w800_,
		_w1205_
	);
	LUT3 #(
		.INIT('h80)
	) name743 (
		_w1197_,
		_w1198_,
		_w1205_,
		_w1206_
	);
	LUT4 #(
		.INIT('h8000)
	) name744 (
		_w1170_,
		_w1195_,
		_w1196_,
		_w1206_,
		_w1207_
	);
	LUT3 #(
		.INIT('h10)
	) name745 (
		_w1073_,
		_w1075_,
		_w1078_,
		_w1208_
	);
	LUT3 #(
		.INIT('h8a)
	) name746 (
		_w1073_,
		_w1075_,
		_w1078_,
		_w1209_
	);
	LUT3 #(
		.INIT('h65)
	) name747 (
		_w1073_,
		_w1075_,
		_w1078_,
		_w1210_
	);
	LUT3 #(
		.INIT('he0)
	) name748 (
		_w489_,
		_w783_,
		_w789_,
		_w1211_
	);
	LUT3 #(
		.INIT('h01)
	) name749 (
		_w489_,
		_w783_,
		_w789_,
		_w1212_
	);
	LUT3 #(
		.INIT('h1e)
	) name750 (
		_w489_,
		_w783_,
		_w789_,
		_w1213_
	);
	LUT2 #(
		.INIT('h1)
	) name751 (
		_w734_,
		_w739_,
		_w1214_
	);
	LUT2 #(
		.INIT('h8)
	) name752 (
		_w734_,
		_w739_,
		_w1215_
	);
	LUT2 #(
		.INIT('h6)
	) name753 (
		_w734_,
		_w739_,
		_w1216_
	);
	LUT4 #(
		.INIT('h0ef1)
	) name754 (
		_w489_,
		_w717_,
		_w719_,
		_w724_,
		_w1217_
	);
	LUT4 #(
		.INIT('h0100)
	) name755 (
		_w1210_,
		_w1213_,
		_w1216_,
		_w1217_,
		_w1218_
	);
	LUT3 #(
		.INIT('he0)
	) name756 (
		_w489_,
		_w1058_,
		_w1063_,
		_w1219_
	);
	LUT3 #(
		.INIT('h01)
	) name757 (
		_w489_,
		_w1058_,
		_w1063_,
		_w1220_
	);
	LUT3 #(
		.INIT('h1e)
	) name758 (
		_w489_,
		_w1058_,
		_w1063_,
		_w1221_
	);
	LUT3 #(
		.INIT('he0)
	) name759 (
		_w489_,
		_w1030_,
		_w1035_,
		_w1222_
	);
	LUT3 #(
		.INIT('h01)
	) name760 (
		_w489_,
		_w1030_,
		_w1035_,
		_w1223_
	);
	LUT3 #(
		.INIT('h1e)
	) name761 (
		_w489_,
		_w1030_,
		_w1035_,
		_w1224_
	);
	LUT2 #(
		.INIT('h9)
	) name762 (
		_w749_,
		_w754_,
		_w1225_
	);
	LUT3 #(
		.INIT('h01)
	) name763 (
		_w489_,
		_w804_,
		_w810_,
		_w1226_
	);
	LUT3 #(
		.INIT('he0)
	) name764 (
		_w489_,
		_w804_,
		_w810_,
		_w1227_
	);
	LUT3 #(
		.INIT('h1e)
	) name765 (
		_w489_,
		_w804_,
		_w810_,
		_w1228_
	);
	LUT4 #(
		.INIT('h0010)
	) name766 (
		_w1221_,
		_w1224_,
		_w1225_,
		_w1228_,
		_w1229_
	);
	LUT2 #(
		.INIT('h8)
	) name767 (
		_w1218_,
		_w1229_,
		_w1230_
	);
	LUT4 #(
		.INIT('h4000)
	) name768 (
		_w1165_,
		_w1207_,
		_w1230_,
		_w1162_,
		_w1231_
	);
	LUT4 #(
		.INIT('h2228)
	) name769 (
		\P1_B_reg/NET0131 ,
		\P1_IR_reg[22]/NET0131 ,
		_w482_,
		_w1097_,
		_w1232_
	);
	LUT2 #(
		.INIT('h4)
	) name770 (
		_w1101_,
		_w1232_,
		_w1233_
	);
	LUT4 #(
		.INIT('h007d)
	) name771 (
		_w1100_,
		_w718_,
		_w1231_,
		_w1233_,
		_w1234_
	);
	LUT2 #(
		.INIT('h1)
	) name772 (
		_w1096_,
		_w1234_,
		_w1235_
	);
	LUT2 #(
		.INIT('h8)
	) name773 (
		_w1096_,
		_w1098_,
		_w1236_
	);
	LUT3 #(
		.INIT('h80)
	) name774 (
		_w1096_,
		_w1098_,
		_w1122_,
		_w1237_
	);
	LUT3 #(
		.INIT('h80)
	) name775 (
		_w1096_,
		_w1098_,
		_w1101_,
		_w1238_
	);
	LUT4 #(
		.INIT('h014f)
	) name776 (
		\P1_B_reg/NET0131 ,
		_w1155_,
		_w1237_,
		_w1238_,
		_w1239_
	);
	LUT3 #(
		.INIT('h10)
	) name777 (
		_w1235_,
		_w1157_,
		_w1239_,
		_w1240_
	);
	LUT4 #(
		.INIT('h0100)
	) name778 (
		_w1118_,
		_w1124_,
		_w1121_,
		_w1240_,
		_w1241_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name779 (
		\P1_IR_reg[31]/NET0131 ,
		_w469_,
		_w474_,
		_w476_,
		_w1242_
	);
	LUT2 #(
		.INIT('h6)
	) name780 (
		\P1_IR_reg[23]/NET0131 ,
		_w1242_,
		_w1243_
	);
	LUT3 #(
		.INIT('h48)
	) name781 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w1244_
	);
	LUT2 #(
		.INIT('h4)
	) name782 (
		_w479_,
		_w488_,
		_w1245_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name783 (
		\P1_IR_reg[31]/NET0131 ,
		_w579_,
		_w578_,
		_w580_,
		_w1246_
	);
	LUT4 #(
		.INIT('h00d5)
	) name784 (
		\P1_IR_reg[31]/NET0131 ,
		_w469_,
		_w470_,
		_w1246_,
		_w1247_
	);
	LUT2 #(
		.INIT('h9)
	) name785 (
		\P1_IR_reg[25]/NET0131 ,
		_w1247_,
		_w1248_
	);
	LUT2 #(
		.INIT('h9)
	) name786 (
		\P1_IR_reg[26]/NET0131 ,
		_w573_,
		_w1249_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name787 (
		\P1_IR_reg[31]/NET0131 ,
		_w483_,
		_w475_,
		_w484_,
		_w1250_
	);
	LUT3 #(
		.INIT('h56)
	) name788 (
		\P1_IR_reg[24]/NET0131 ,
		_w482_,
		_w1250_,
		_w1251_
	);
	LUT3 #(
		.INIT('h40)
	) name789 (
		_w1249_,
		_w1251_,
		_w1248_,
		_w1252_
	);
	LUT4 #(
		.INIT('h3313)
	) name790 (
		_w1237_,
		_w1243_,
		_w1245_,
		_w1252_,
		_w1253_
	);
	LUT3 #(
		.INIT('ha2)
	) name791 (
		\P1_B_reg/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1253_,
		_w1254_
	);
	LUT4 #(
		.INIT('hff70)
	) name792 (
		_w1116_,
		_w1241_,
		_w1244_,
		_w1254_,
		_w1255_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_IR_reg[18]/NET0131 ,
		_w1256_
	);
	LUT3 #(
		.INIT('h01)
	) name794 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w1257_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[12]/NET0131 ,
		_w1258_
	);
	LUT4 #(
		.INIT('h0001)
	) name796 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[2]/NET0131 ,
		\P2_IR_reg[3]/NET0131 ,
		_w1259_
	);
	LUT4 #(
		.INIT('h0001)
	) name797 (
		\P2_IR_reg[4]/NET0131 ,
		\P2_IR_reg[5]/NET0131 ,
		\P2_IR_reg[6]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		_w1260_
	);
	LUT2 #(
		.INIT('h8)
	) name798 (
		_w1259_,
		_w1260_,
		_w1261_
	);
	LUT4 #(
		.INIT('h8000)
	) name799 (
		_w1257_,
		_w1258_,
		_w1259_,
		_w1260_,
		_w1262_
	);
	LUT4 #(
		.INIT('h0001)
	) name800 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[16]/NET0131 ,
		_w1263_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name801 (
		\P2_IR_reg[31]/NET0131 ,
		_w1256_,
		_w1262_,
		_w1263_,
		_w1264_
	);
	LUT4 #(
		.INIT('h0001)
	) name802 (
		\P2_IR_reg[19]/NET0131 ,
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		_w1265_
	);
	LUT2 #(
		.INIT('h2)
	) name803 (
		\P2_IR_reg[31]/NET0131 ,
		_w1265_,
		_w1266_
	);
	LUT3 #(
		.INIT('h56)
	) name804 (
		\P2_IR_reg[23]/NET0131 ,
		_w1264_,
		_w1266_,
		_w1267_
	);
	LUT3 #(
		.INIT('h40)
	) name805 (
		\P2_IR_reg[13]/NET0131 ,
		_w1257_,
		_w1258_,
		_w1268_
	);
	LUT4 #(
		.INIT('h0001)
	) name806 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[16]/NET0131 ,
		\P2_IR_reg[17]/NET0131 ,
		_w1269_
	);
	LUT2 #(
		.INIT('h1)
	) name807 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_IR_reg[19]/NET0131 ,
		_w1270_
	);
	LUT2 #(
		.INIT('h8)
	) name808 (
		_w1269_,
		_w1270_,
		_w1271_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name809 (
		\P2_IR_reg[31]/NET0131 ,
		_w1261_,
		_w1268_,
		_w1271_,
		_w1272_
	);
	LUT4 #(
		.INIT('h0001)
	) name810 (
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1273_
	);
	LUT2 #(
		.INIT('h2)
	) name811 (
		\P2_IR_reg[31]/NET0131 ,
		_w1273_,
		_w1274_
	);
	LUT3 #(
		.INIT('h56)
	) name812 (
		\P2_IR_reg[24]/NET0131 ,
		_w1272_,
		_w1274_,
		_w1275_
	);
	LUT2 #(
		.INIT('h4)
	) name813 (
		\P2_IR_reg[24]/NET0131 ,
		_w1273_,
		_w1276_
	);
	LUT3 #(
		.INIT('h01)
	) name814 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_IR_reg[18]/NET0131 ,
		\P2_IR_reg[19]/NET0131 ,
		_w1277_
	);
	LUT4 #(
		.INIT('h4000)
	) name815 (
		\P2_IR_reg[24]/NET0131 ,
		_w1263_,
		_w1273_,
		_w1277_,
		_w1278_
	);
	LUT4 #(
		.INIT('h5999)
	) name816 (
		\P2_IR_reg[25]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1262_,
		_w1278_,
		_w1279_
	);
	LUT3 #(
		.INIT('h40)
	) name817 (
		\P2_IR_reg[25]/NET0131 ,
		_w1269_,
		_w1270_,
		_w1280_
	);
	LUT4 #(
		.INIT('h8000)
	) name818 (
		_w1261_,
		_w1276_,
		_w1268_,
		_w1280_,
		_w1281_
	);
	LUT3 #(
		.INIT('h59)
	) name819 (
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1281_,
		_w1282_
	);
	LUT4 #(
		.INIT('h0a06)
	) name820 (
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1279_,
		_w1281_,
		_w1283_
	);
	LUT2 #(
		.INIT('h8)
	) name821 (
		_w1275_,
		_w1283_,
		_w1284_
	);
	LUT3 #(
		.INIT('h15)
	) name822 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1285_
	);
	LUT4 #(
		.INIT('ha060)
	) name823 (
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1279_,
		_w1281_,
		_w1286_
	);
	LUT4 #(
		.INIT('h8882)
	) name824 (
		\P2_B_reg/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		_w1272_,
		_w1274_,
		_w1287_
	);
	LUT2 #(
		.INIT('h8)
	) name825 (
		_w1286_,
		_w1287_,
		_w1288_
	);
	LUT4 #(
		.INIT('h1114)
	) name826 (
		\P2_B_reg/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		_w1272_,
		_w1274_,
		_w1289_
	);
	LUT2 #(
		.INIT('h8)
	) name827 (
		_w1286_,
		_w1289_,
		_w1290_
	);
	LUT3 #(
		.INIT('h35)
	) name828 (
		\P2_d_reg[0]/NET0131 ,
		_w1275_,
		_w1282_,
		_w1291_
	);
	LUT3 #(
		.INIT('hef)
	) name829 (
		_w1290_,
		_w1288_,
		_w1291_,
		_w1292_
	);
	LUT4 #(
		.INIT('ha060)
	) name830 (
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_d_reg[1]/NET0131 ,
		_w1281_,
		_w1293_
	);
	LUT4 #(
		.INIT('h0509)
	) name831 (
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1279_,
		_w1281_,
		_w1294_
	);
	LUT2 #(
		.INIT('h1)
	) name832 (
		_w1293_,
		_w1294_,
		_w1295_
	);
	LUT4 #(
		.INIT('hc1c5)
	) name833 (
		\P2_d_reg[1]/NET0131 ,
		_w1279_,
		_w1282_,
		_w1289_,
		_w1296_
	);
	LUT2 #(
		.INIT('hb)
	) name834 (
		_w1288_,
		_w1296_,
		_w1297_
	);
	LUT4 #(
		.INIT('h0010)
	) name835 (
		_w1290_,
		_w1288_,
		_w1291_,
		_w1295_,
		_w1298_
	);
	LUT4 #(
		.INIT('h0001)
	) name836 (
		\P2_IR_reg[23]/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		\P2_IR_reg[25]/NET0131 ,
		\P2_IR_reg[26]/NET0131 ,
		_w1299_
	);
	LUT2 #(
		.INIT('h8)
	) name837 (
		_w1265_,
		_w1299_,
		_w1300_
	);
	LUT4 #(
		.INIT('h8000)
	) name838 (
		_w1256_,
		_w1262_,
		_w1263_,
		_w1300_,
		_w1301_
	);
	LUT3 #(
		.INIT('ha6)
	) name839 (
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1301_,
		_w1302_
	);
	LUT4 #(
		.INIT('h0001)
	) name840 (
		\P2_IR_reg[24]/NET0131 ,
		\P2_IR_reg[25]/NET0131 ,
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		_w1303_
	);
	LUT4 #(
		.INIT('h8000)
	) name841 (
		_w1261_,
		_w1268_,
		_w1271_,
		_w1303_,
		_w1304_
	);
	LUT4 #(
		.INIT('h5a56)
	) name842 (
		\P2_IR_reg[28]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1274_,
		_w1304_,
		_w1305_
	);
	LUT2 #(
		.INIT('h1)
	) name843 (
		_w1302_,
		_w1305_,
		_w1306_
	);
	LUT2 #(
		.INIT('h8)
	) name844 (
		\P1_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w1307_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		\P1_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w1308_
	);
	LUT2 #(
		.INIT('h8)
	) name846 (
		\P1_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w1309_
	);
	LUT2 #(
		.INIT('h1)
	) name847 (
		\P1_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w1310_
	);
	LUT4 #(
		.INIT('hfac8)
	) name848 (
		\P1_datao_reg[11]/NET0131 ,
		\P1_datao_reg[12]/NET0131 ,
		\si[11]_pad ,
		\si[12]_pad ,
		_w1311_
	);
	LUT2 #(
		.INIT('h8)
	) name849 (
		\P1_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w1312_
	);
	LUT2 #(
		.INIT('h1)
	) name850 (
		\P1_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w1313_
	);
	LUT2 #(
		.INIT('h8)
	) name851 (
		\P1_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w1314_
	);
	LUT4 #(
		.INIT('he8a0)
	) name852 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\si[10]_pad ,
		\si[9]_pad ,
		_w1315_
	);
	LUT4 #(
		.INIT('h1115)
	) name853 (
		_w1309_,
		_w1311_,
		_w1312_,
		_w1315_,
		_w1316_
	);
	LUT2 #(
		.INIT('h1)
	) name854 (
		\P1_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w1317_
	);
	LUT2 #(
		.INIT('h1)
	) name855 (
		\P1_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w1318_
	);
	LUT2 #(
		.INIT('h8)
	) name856 (
		\P1_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w1319_
	);
	LUT4 #(
		.INIT('hec80)
	) name857 (
		\P1_datao_reg[0]/NET0131 ,
		\P1_datao_reg[1]/NET0131 ,
		\si[0]_pad ,
		\si[1]_pad ,
		_w1320_
	);
	LUT4 #(
		.INIT('h135f)
	) name858 (
		\P1_datao_reg[2]/NET0131 ,
		\P1_datao_reg[3]/NET0131 ,
		\si[2]_pad ,
		\si[3]_pad ,
		_w1321_
	);
	LUT4 #(
		.INIT('h1055)
	) name859 (
		_w1317_,
		_w1318_,
		_w1320_,
		_w1321_,
		_w1322_
	);
	LUT3 #(
		.INIT('he8)
	) name860 (
		\P1_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w1322_,
		_w1323_
	);
	LUT4 #(
		.INIT('hfac8)
	) name861 (
		\P1_datao_reg[7]/NET0131 ,
		\P1_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w1324_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		\P1_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w1325_
	);
	LUT4 #(
		.INIT('hfac8)
	) name863 (
		\P1_datao_reg[5]/NET0131 ,
		\P1_datao_reg[6]/NET0131 ,
		\si[5]_pad ,
		\si[6]_pad ,
		_w1326_
	);
	LUT2 #(
		.INIT('h8)
	) name864 (
		_w1324_,
		_w1326_,
		_w1327_
	);
	LUT4 #(
		.INIT('he800)
	) name865 (
		\P1_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w1322_,
		_w1327_,
		_w1328_
	);
	LUT2 #(
		.INIT('h8)
	) name866 (
		\P1_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w1329_
	);
	LUT2 #(
		.INIT('h8)
	) name867 (
		\P1_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w1330_
	);
	LUT2 #(
		.INIT('h8)
	) name868 (
		\P1_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w1331_
	);
	LUT4 #(
		.INIT('hec80)
	) name869 (
		\P1_datao_reg[5]/NET0131 ,
		\P1_datao_reg[6]/NET0131 ,
		\si[5]_pad ,
		\si[6]_pad ,
		_w1332_
	);
	LUT4 #(
		.INIT('h1115)
	) name870 (
		_w1329_,
		_w1324_,
		_w1330_,
		_w1332_,
		_w1333_
	);
	LUT2 #(
		.INIT('h1)
	) name871 (
		\P1_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w1334_
	);
	LUT4 #(
		.INIT('hfac8)
	) name872 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\si[10]_pad ,
		\si[9]_pad ,
		_w1335_
	);
	LUT2 #(
		.INIT('h8)
	) name873 (
		_w1311_,
		_w1335_,
		_w1336_
	);
	LUT4 #(
		.INIT('h20aa)
	) name874 (
		_w1316_,
		_w1328_,
		_w1333_,
		_w1336_,
		_w1337_
	);
	LUT4 #(
		.INIT('hfac8)
	) name875 (
		\P1_datao_reg[19]/NET0131 ,
		\P1_datao_reg[20]/NET0131 ,
		\si[19]_pad ,
		\si[20]_pad ,
		_w1338_
	);
	LUT4 #(
		.INIT('hfac8)
	) name876 (
		\P1_datao_reg[17]/NET0131 ,
		\P1_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w1339_
	);
	LUT2 #(
		.INIT('h8)
	) name877 (
		_w1338_,
		_w1339_,
		_w1340_
	);
	LUT2 #(
		.INIT('h1)
	) name878 (
		\P1_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w1341_
	);
	LUT4 #(
		.INIT('hfac8)
	) name879 (
		\P1_datao_reg[15]/NET0131 ,
		\P1_datao_reg[16]/NET0131 ,
		\si[15]_pad ,
		\si[16]_pad ,
		_w1342_
	);
	LUT2 #(
		.INIT('h1)
	) name880 (
		\P1_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w1343_
	);
	LUT2 #(
		.INIT('h1)
	) name881 (
		\P1_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w1344_
	);
	LUT4 #(
		.INIT('hfac8)
	) name882 (
		\P1_datao_reg[13]/NET0131 ,
		\P1_datao_reg[14]/NET0131 ,
		\si[13]_pad ,
		\si[14]_pad ,
		_w1345_
	);
	LUT2 #(
		.INIT('h8)
	) name883 (
		_w1342_,
		_w1345_,
		_w1346_
	);
	LUT4 #(
		.INIT('h8000)
	) name884 (
		_w1338_,
		_w1339_,
		_w1342_,
		_w1345_,
		_w1347_
	);
	LUT4 #(
		.INIT('hec80)
	) name885 (
		\P1_datao_reg[19]/NET0131 ,
		\P1_datao_reg[20]/NET0131 ,
		\si[19]_pad ,
		\si[20]_pad ,
		_w1348_
	);
	LUT4 #(
		.INIT('hec80)
	) name886 (
		\P1_datao_reg[17]/NET0131 ,
		\P1_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w1349_
	);
	LUT3 #(
		.INIT('h15)
	) name887 (
		_w1348_,
		_w1338_,
		_w1349_,
		_w1350_
	);
	LUT4 #(
		.INIT('hec80)
	) name888 (
		\P1_datao_reg[15]/NET0131 ,
		\P1_datao_reg[16]/NET0131 ,
		\si[15]_pad ,
		\si[16]_pad ,
		_w1351_
	);
	LUT4 #(
		.INIT('hec80)
	) name889 (
		\P1_datao_reg[13]/NET0131 ,
		\P1_datao_reg[14]/NET0131 ,
		\si[13]_pad ,
		\si[14]_pad ,
		_w1352_
	);
	LUT3 #(
		.INIT('h15)
	) name890 (
		_w1351_,
		_w1342_,
		_w1352_,
		_w1353_
	);
	LUT3 #(
		.INIT('ha2)
	) name891 (
		_w1350_,
		_w1340_,
		_w1353_,
		_w1354_
	);
	LUT3 #(
		.INIT('hb0)
	) name892 (
		_w1337_,
		_w1347_,
		_w1354_,
		_w1355_
	);
	LUT2 #(
		.INIT('h1)
	) name893 (
		\P1_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w1356_
	);
	LUT2 #(
		.INIT('h1)
	) name894 (
		\P1_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w1357_
	);
	LUT4 #(
		.INIT('hfac8)
	) name895 (
		\P1_datao_reg[25]/NET0131 ,
		\P1_datao_reg[26]/NET0131 ,
		\si[25]_pad ,
		\si[26]_pad ,
		_w1358_
	);
	LUT2 #(
		.INIT('h1)
	) name896 (
		\P1_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w1359_
	);
	LUT4 #(
		.INIT('hfac8)
	) name897 (
		\P1_datao_reg[23]/NET0131 ,
		\P1_datao_reg[24]/NET0131 ,
		\si[23]_pad ,
		\si[24]_pad ,
		_w1360_
	);
	LUT4 #(
		.INIT('hfac8)
	) name898 (
		\P1_datao_reg[21]/NET0131 ,
		\P1_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w1361_
	);
	LUT2 #(
		.INIT('h8)
	) name899 (
		_w1360_,
		_w1361_,
		_w1362_
	);
	LUT4 #(
		.INIT('h4000)
	) name900 (
		_w1356_,
		_w1358_,
		_w1360_,
		_w1361_,
		_w1363_
	);
	LUT4 #(
		.INIT('h4f00)
	) name901 (
		_w1337_,
		_w1347_,
		_w1354_,
		_w1363_,
		_w1364_
	);
	LUT4 #(
		.INIT('h135f)
	) name902 (
		\P1_datao_reg[27]/NET0131 ,
		\P1_datao_reg[28]/NET0131 ,
		\si[27]_pad ,
		\si[28]_pad ,
		_w1365_
	);
	LUT4 #(
		.INIT('hec80)
	) name903 (
		\P1_datao_reg[25]/NET0131 ,
		\P1_datao_reg[26]/NET0131 ,
		\si[25]_pad ,
		\si[26]_pad ,
		_w1366_
	);
	LUT4 #(
		.INIT('hec80)
	) name904 (
		\P1_datao_reg[23]/NET0131 ,
		\P1_datao_reg[24]/NET0131 ,
		\si[23]_pad ,
		\si[24]_pad ,
		_w1367_
	);
	LUT4 #(
		.INIT('hec80)
	) name905 (
		\P1_datao_reg[21]/NET0131 ,
		\P1_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w1368_
	);
	LUT3 #(
		.INIT('h13)
	) name906 (
		_w1360_,
		_w1367_,
		_w1368_,
		_w1369_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name907 (
		_w1358_,
		_w1360_,
		_w1367_,
		_w1368_,
		_w1370_
	);
	LUT4 #(
		.INIT('h888c)
	) name908 (
		_w1356_,
		_w1365_,
		_w1366_,
		_w1370_,
		_w1371_
	);
	LUT3 #(
		.INIT('h45)
	) name909 (
		_w1308_,
		_w1364_,
		_w1371_,
		_w1372_
	);
	LUT4 #(
		.INIT('h6595)
	) name910 (
		\P1_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w568_,
		_w1372_,
		_w1373_
	);
	LUT2 #(
		.INIT('h1)
	) name911 (
		_w1306_,
		_w1373_,
		_w1374_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[28]/NET0131 ,
		_w1375_
	);
	LUT4 #(
		.INIT('h0001)
	) name913 (
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[28]/NET0131 ,
		\P2_IR_reg[29]/NET0131 ,
		_w1376_
	);
	LUT2 #(
		.INIT('h2)
	) name914 (
		\P2_IR_reg[31]/NET0131 ,
		_w1376_,
		_w1377_
	);
	LUT4 #(
		.INIT('h55a6)
	) name915 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1281_,
		_w1377_,
		_w1378_
	);
	LUT4 #(
		.INIT('h0001)
	) name916 (
		\P2_IR_reg[25]/NET0131 ,
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[28]/NET0131 ,
		_w1379_
	);
	LUT2 #(
		.INIT('h2)
	) name917 (
		\P2_IR_reg[31]/NET0131 ,
		_w1379_,
		_w1380_
	);
	LUT4 #(
		.INIT('h00d5)
	) name918 (
		\P2_IR_reg[31]/NET0131 ,
		_w1262_,
		_w1278_,
		_w1380_,
		_w1381_
	);
	LUT2 #(
		.INIT('h9)
	) name919 (
		\P2_IR_reg[29]/NET0131 ,
		_w1381_,
		_w1382_
	);
	LUT2 #(
		.INIT('h8)
	) name920 (
		_w1378_,
		_w1382_,
		_w1383_
	);
	LUT4 #(
		.INIT('h8000)
	) name921 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		\P2_reg3_reg[6]/NET0131 ,
		_w1384_
	);
	LUT4 #(
		.INIT('h8000)
	) name922 (
		\P2_reg3_reg[7]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		\P2_reg3_reg[9]/NET0131 ,
		_w1384_,
		_w1385_
	);
	LUT3 #(
		.INIT('h80)
	) name923 (
		\P2_reg3_reg[11]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		\P2_reg3_reg[13]/NET0131 ,
		_w1386_
	);
	LUT3 #(
		.INIT('h80)
	) name924 (
		\P2_reg3_reg[10]/NET0131 ,
		_w1385_,
		_w1386_,
		_w1387_
	);
	LUT4 #(
		.INIT('h8000)
	) name925 (
		\P2_reg3_reg[10]/NET0131 ,
		\P2_reg3_reg[14]/NET0131 ,
		_w1385_,
		_w1386_,
		_w1388_
	);
	LUT2 #(
		.INIT('h8)
	) name926 (
		\P2_reg3_reg[15]/NET0131 ,
		\P2_reg3_reg[16]/NET0131 ,
		_w1389_
	);
	LUT2 #(
		.INIT('h8)
	) name927 (
		\P2_reg3_reg[17]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		_w1390_
	);
	LUT2 #(
		.INIT('h8)
	) name928 (
		\P2_reg3_reg[20]/NET0131 ,
		\P2_reg3_reg[21]/NET0131 ,
		_w1391_
	);
	LUT4 #(
		.INIT('h8000)
	) name929 (
		\P2_reg3_reg[19]/NET0131 ,
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		\P2_reg3_reg[24]/NET0131 ,
		_w1392_
	);
	LUT2 #(
		.INIT('h8)
	) name930 (
		_w1391_,
		_w1392_,
		_w1393_
	);
	LUT4 #(
		.INIT('h8000)
	) name931 (
		_w1388_,
		_w1389_,
		_w1390_,
		_w1393_,
		_w1394_
	);
	LUT4 #(
		.INIT('h8000)
	) name932 (
		\P2_reg3_reg[25]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w1395_
	);
	LUT2 #(
		.INIT('h8)
	) name933 (
		_w1394_,
		_w1395_,
		_w1396_
	);
	LUT4 #(
		.INIT('h8000)
	) name934 (
		_w1378_,
		_w1382_,
		_w1394_,
		_w1395_,
		_w1397_
	);
	LUT3 #(
		.INIT('h02)
	) name935 (
		\P2_reg0_reg[29]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1398_
	);
	LUT4 #(
		.INIT('hf53f)
	) name936 (
		\P2_reg1_reg[29]/NET0131 ,
		\P2_reg2_reg[29]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1399_
	);
	LUT3 #(
		.INIT('h10)
	) name937 (
		_w1398_,
		_w1397_,
		_w1399_,
		_w1400_
	);
	LUT3 #(
		.INIT('hef)
	) name938 (
		_w1398_,
		_w1397_,
		_w1399_,
		_w1401_
	);
	LUT3 #(
		.INIT('h10)
	) name939 (
		_w1306_,
		_w1373_,
		_w1400_,
		_w1402_
	);
	LUT3 #(
		.INIT('h0e)
	) name940 (
		_w1306_,
		_w1373_,
		_w1400_,
		_w1403_
	);
	LUT3 #(
		.INIT('he1)
	) name941 (
		_w1306_,
		_w1373_,
		_w1400_,
		_w1404_
	);
	LUT4 #(
		.INIT('h135f)
	) name942 (
		\P1_datao_reg[26]/NET0131 ,
		\P1_datao_reg[27]/NET0131 ,
		\si[26]_pad ,
		\si[27]_pad ,
		_w1405_
	);
	LUT4 #(
		.INIT('hec80)
	) name943 (
		\P1_datao_reg[24]/NET0131 ,
		\P1_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w1406_
	);
	LUT4 #(
		.INIT('h1505)
	) name944 (
		_w1356_,
		_w1357_,
		_w1405_,
		_w1406_,
		_w1407_
	);
	LUT3 #(
		.INIT('h10)
	) name945 (
		_w1341_,
		_w1310_,
		_w1345_,
		_w1408_
	);
	LUT4 #(
		.INIT('hfac8)
	) name946 (
		\P1_datao_reg[4]/NET0131 ,
		\P1_datao_reg[5]/NET0131 ,
		\si[4]_pad ,
		\si[5]_pad ,
		_w1409_
	);
	LUT4 #(
		.INIT('hfac8)
	) name947 (
		\P1_datao_reg[6]/NET0131 ,
		\P1_datao_reg[7]/NET0131 ,
		\si[6]_pad ,
		\si[7]_pad ,
		_w1410_
	);
	LUT4 #(
		.INIT('hec80)
	) name948 (
		\P1_datao_reg[4]/NET0131 ,
		\P1_datao_reg[5]/NET0131 ,
		\si[4]_pad ,
		\si[5]_pad ,
		_w1411_
	);
	LUT4 #(
		.INIT('h0515)
	) name949 (
		_w1330_,
		_w1331_,
		_w1410_,
		_w1411_,
		_w1412_
	);
	LUT4 #(
		.INIT('h7f00)
	) name950 (
		_w1322_,
		_w1409_,
		_w1410_,
		_w1412_,
		_w1413_
	);
	LUT4 #(
		.INIT('hfac8)
	) name951 (
		\P1_datao_reg[8]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\si[8]_pad ,
		\si[9]_pad ,
		_w1414_
	);
	LUT4 #(
		.INIT('hfac8)
	) name952 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w1415_
	);
	LUT2 #(
		.INIT('h8)
	) name953 (
		_w1414_,
		_w1415_,
		_w1416_
	);
	LUT4 #(
		.INIT('hec80)
	) name954 (
		\P1_datao_reg[8]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\si[8]_pad ,
		\si[9]_pad ,
		_w1417_
	);
	LUT4 #(
		.INIT('h0515)
	) name955 (
		_w1312_,
		_w1314_,
		_w1415_,
		_w1417_,
		_w1418_
	);
	LUT4 #(
		.INIT('hfac8)
	) name956 (
		\P1_datao_reg[14]/NET0131 ,
		\P1_datao_reg[15]/NET0131 ,
		\si[14]_pad ,
		\si[15]_pad ,
		_w1419_
	);
	LUT4 #(
		.INIT('hec80)
	) name957 (
		\P1_datao_reg[12]/NET0131 ,
		\P1_datao_reg[13]/NET0131 ,
		\si[12]_pad ,
		\si[13]_pad ,
		_w1420_
	);
	LUT4 #(
		.INIT('hec80)
	) name958 (
		\P1_datao_reg[14]/NET0131 ,
		\P1_datao_reg[15]/NET0131 ,
		\si[14]_pad ,
		\si[15]_pad ,
		_w1421_
	);
	LUT3 #(
		.INIT('h07)
	) name959 (
		_w1419_,
		_w1420_,
		_w1421_,
		_w1422_
	);
	LUT3 #(
		.INIT('hd0)
	) name960 (
		_w1408_,
		_w1418_,
		_w1422_,
		_w1423_
	);
	LUT4 #(
		.INIT('hdf00)
	) name961 (
		_w1408_,
		_w1413_,
		_w1416_,
		_w1423_,
		_w1424_
	);
	LUT4 #(
		.INIT('hfac8)
	) name962 (
		\P1_datao_reg[18]/NET0131 ,
		\P1_datao_reg[19]/NET0131 ,
		\si[18]_pad ,
		\si[19]_pad ,
		_w1425_
	);
	LUT4 #(
		.INIT('hfac8)
	) name963 (
		\P1_datao_reg[16]/NET0131 ,
		\P1_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w1426_
	);
	LUT2 #(
		.INIT('h8)
	) name964 (
		_w1425_,
		_w1426_,
		_w1427_
	);
	LUT4 #(
		.INIT('hec80)
	) name965 (
		\P1_datao_reg[18]/NET0131 ,
		\P1_datao_reg[19]/NET0131 ,
		\si[18]_pad ,
		\si[19]_pad ,
		_w1428_
	);
	LUT4 #(
		.INIT('hec80)
	) name966 (
		\P1_datao_reg[16]/NET0131 ,
		\P1_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w1429_
	);
	LUT3 #(
		.INIT('h13)
	) name967 (
		_w1425_,
		_w1428_,
		_w1429_,
		_w1430_
	);
	LUT3 #(
		.INIT('hb0)
	) name968 (
		_w1424_,
		_w1427_,
		_w1430_,
		_w1431_
	);
	LUT4 #(
		.INIT('hfac8)
	) name969 (
		\P1_datao_reg[22]/NET0131 ,
		\P1_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w1432_
	);
	LUT4 #(
		.INIT('hfac8)
	) name970 (
		\P1_datao_reg[20]/NET0131 ,
		\P1_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w1433_
	);
	LUT2 #(
		.INIT('h8)
	) name971 (
		_w1432_,
		_w1433_,
		_w1434_
	);
	LUT4 #(
		.INIT('h4f00)
	) name972 (
		_w1424_,
		_w1427_,
		_w1430_,
		_w1434_,
		_w1435_
	);
	LUT4 #(
		.INIT('hec80)
	) name973 (
		\P1_datao_reg[22]/NET0131 ,
		\P1_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w1436_
	);
	LUT4 #(
		.INIT('hec80)
	) name974 (
		\P1_datao_reg[20]/NET0131 ,
		\P1_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w1437_
	);
	LUT3 #(
		.INIT('h13)
	) name975 (
		_w1432_,
		_w1436_,
		_w1437_,
		_w1438_
	);
	LUT3 #(
		.INIT('h04)
	) name976 (
		_w1356_,
		_w1358_,
		_w1359_,
		_w1439_
	);
	LUT4 #(
		.INIT('h1055)
	) name977 (
		_w1407_,
		_w1435_,
		_w1438_,
		_w1439_,
		_w1440_
	);
	LUT4 #(
		.INIT('h9565)
	) name978 (
		\P1_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w568_,
		_w1440_,
		_w1441_
	);
	LUT2 #(
		.INIT('h1)
	) name979 (
		_w1306_,
		_w1441_,
		_w1442_
	);
	LUT4 #(
		.INIT('h8000)
	) name980 (
		\P2_reg3_reg[25]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		\P2_reg3_reg[27]/NET0131 ,
		_w1394_,
		_w1443_
	);
	LUT2 #(
		.INIT('h6)
	) name981 (
		\P2_reg3_reg[28]/NET0131 ,
		_w1443_,
		_w1444_
	);
	LUT3 #(
		.INIT('h48)
	) name982 (
		\P2_reg3_reg[28]/NET0131 ,
		_w1383_,
		_w1443_,
		_w1445_
	);
	LUT3 #(
		.INIT('h02)
	) name983 (
		\P2_reg0_reg[28]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1446_
	);
	LUT4 #(
		.INIT('hf53f)
	) name984 (
		\P2_reg1_reg[28]/NET0131 ,
		\P2_reg2_reg[28]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1447_
	);
	LUT2 #(
		.INIT('h4)
	) name985 (
		_w1446_,
		_w1447_,
		_w1448_
	);
	LUT2 #(
		.INIT('h4)
	) name986 (
		_w1445_,
		_w1448_,
		_w1449_
	);
	LUT2 #(
		.INIT('hb)
	) name987 (
		_w1445_,
		_w1448_,
		_w1450_
	);
	LUT3 #(
		.INIT('he0)
	) name988 (
		_w1306_,
		_w1441_,
		_w1449_,
		_w1451_
	);
	LUT2 #(
		.INIT('h2)
	) name989 (
		\P1_datao_reg[27]/NET0131 ,
		_w568_,
		_w1452_
	);
	LUT2 #(
		.INIT('h6)
	) name990 (
		\P1_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w1453_
	);
	LUT3 #(
		.INIT('h13)
	) name991 (
		_w1358_,
		_w1366_,
		_w1367_,
		_w1454_
	);
	LUT2 #(
		.INIT('h8)
	) name992 (
		_w1358_,
		_w1360_,
		_w1455_
	);
	LUT2 #(
		.INIT('h8)
	) name993 (
		_w1361_,
		_w1338_,
		_w1456_
	);
	LUT2 #(
		.INIT('h8)
	) name994 (
		_w1339_,
		_w1342_,
		_w1457_
	);
	LUT4 #(
		.INIT('h8000)
	) name995 (
		_w1361_,
		_w1338_,
		_w1339_,
		_w1342_,
		_w1458_
	);
	LUT3 #(
		.INIT('h17)
	) name996 (
		\P1_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w1320_,
		_w1459_
	);
	LUT4 #(
		.INIT('h0e08)
	) name997 (
		\P1_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w1317_,
		_w1320_,
		_w1460_
	);
	LUT4 #(
		.INIT('h135f)
	) name998 (
		\P1_datao_reg[3]/NET0131 ,
		\P1_datao_reg[4]/NET0131 ,
		\si[3]_pad ,
		\si[4]_pad ,
		_w1461_
	);
	LUT2 #(
		.INIT('h4)
	) name999 (
		_w1325_,
		_w1409_,
		_w1462_
	);
	LUT4 #(
		.INIT('h1055)
	) name1000 (
		_w1332_,
		_w1460_,
		_w1461_,
		_w1462_,
		_w1463_
	);
	LUT3 #(
		.INIT('h04)
	) name1001 (
		_w1313_,
		_w1324_,
		_w1334_,
		_w1464_
	);
	LUT4 #(
		.INIT('h135f)
	) name1002 (
		\P1_datao_reg[7]/NET0131 ,
		\P1_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w1465_
	);
	LUT4 #(
		.INIT('h3323)
	) name1003 (
		_w1313_,
		_w1315_,
		_w1414_,
		_w1465_,
		_w1466_
	);
	LUT3 #(
		.INIT('hb0)
	) name1004 (
		_w1463_,
		_w1464_,
		_w1466_,
		_w1467_
	);
	LUT3 #(
		.INIT('h04)
	) name1005 (
		_w1343_,
		_w1311_,
		_w1344_,
		_w1468_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1006 (
		_w1463_,
		_w1464_,
		_w1466_,
		_w1468_,
		_w1469_
	);
	LUT3 #(
		.INIT('h07)
	) name1007 (
		_w1361_,
		_w1348_,
		_w1368_,
		_w1470_
	);
	LUT4 #(
		.INIT('h135f)
	) name1008 (
		\P1_datao_reg[11]/NET0131 ,
		\P1_datao_reg[12]/NET0131 ,
		\si[11]_pad ,
		\si[12]_pad ,
		_w1471_
	);
	LUT4 #(
		.INIT('h5545)
	) name1009 (
		_w1352_,
		_w1310_,
		_w1345_,
		_w1471_,
		_w1472_
	);
	LUT3 #(
		.INIT('h15)
	) name1010 (
		_w1349_,
		_w1339_,
		_w1351_,
		_w1473_
	);
	LUT3 #(
		.INIT('hd0)
	) name1011 (
		_w1457_,
		_w1472_,
		_w1473_,
		_w1474_
	);
	LUT4 #(
		.INIT('h08aa)
	) name1012 (
		_w1456_,
		_w1457_,
		_w1472_,
		_w1473_,
		_w1475_
	);
	LUT2 #(
		.INIT('h2)
	) name1013 (
		_w1470_,
		_w1475_,
		_w1476_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1014 (
		_w1455_,
		_w1458_,
		_w1469_,
		_w1476_,
		_w1477_
	);
	LUT4 #(
		.INIT('h2282)
	) name1015 (
		_w568_,
		_w1453_,
		_w1454_,
		_w1477_,
		_w1478_
	);
	LUT3 #(
		.INIT('h54)
	) name1016 (
		_w1306_,
		_w1452_,
		_w1478_,
		_w1479_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1017 (
		\P2_reg3_reg[25]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		\P2_reg3_reg[27]/NET0131 ,
		_w1394_,
		_w1480_
	);
	LUT3 #(
		.INIT('h20)
	) name1018 (
		\P2_reg1_reg[27]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1481_
	);
	LUT4 #(
		.INIT('hff35)
	) name1019 (
		\P2_reg0_reg[27]/NET0131 ,
		\P2_reg2_reg[27]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1482_
	);
	LUT4 #(
		.INIT('h1300)
	) name1020 (
		_w1383_,
		_w1481_,
		_w1480_,
		_w1482_,
		_w1483_
	);
	LUT4 #(
		.INIT('hecff)
	) name1021 (
		_w1383_,
		_w1481_,
		_w1480_,
		_w1482_,
		_w1484_
	);
	LUT4 #(
		.INIT('hab00)
	) name1022 (
		_w1306_,
		_w1452_,
		_w1478_,
		_w1483_,
		_w1485_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1023 (
		\P1_datao_reg[24]/NET0131 ,
		\P1_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w1486_
	);
	LUT3 #(
		.INIT('h15)
	) name1024 (
		_w1406_,
		_w1436_,
		_w1486_,
		_w1487_
	);
	LUT2 #(
		.INIT('h8)
	) name1025 (
		_w1432_,
		_w1486_,
		_w1488_
	);
	LUT3 #(
		.INIT('h07)
	) name1026 (
		_w1428_,
		_w1433_,
		_w1437_,
		_w1489_
	);
	LUT2 #(
		.INIT('h8)
	) name1027 (
		_w1419_,
		_w1426_,
		_w1490_
	);
	LUT3 #(
		.INIT('h07)
	) name1028 (
		_w1322_,
		_w1409_,
		_w1411_,
		_w1491_
	);
	LUT2 #(
		.INIT('h8)
	) name1029 (
		_w1410_,
		_w1414_,
		_w1492_
	);
	LUT4 #(
		.INIT('hf800)
	) name1030 (
		_w1322_,
		_w1409_,
		_w1411_,
		_w1492_,
		_w1493_
	);
	LUT4 #(
		.INIT('h135f)
	) name1031 (
		\P1_datao_reg[6]/NET0131 ,
		\P1_datao_reg[7]/NET0131 ,
		\si[6]_pad ,
		\si[7]_pad ,
		_w1494_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1032 (
		_w1324_,
		_w1334_,
		_w1417_,
		_w1494_,
		_w1495_
	);
	LUT3 #(
		.INIT('h02)
	) name1033 (
		_w1311_,
		_w1313_,
		_w1344_,
		_w1496_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1034 (
		_w1490_,
		_w1493_,
		_w1495_,
		_w1496_,
		_w1497_
	);
	LUT4 #(
		.INIT('h135f)
	) name1035 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w1498_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1036 (
		_w1311_,
		_w1344_,
		_w1420_,
		_w1498_,
		_w1499_
	);
	LUT3 #(
		.INIT('h07)
	) name1037 (
		_w1421_,
		_w1426_,
		_w1429_,
		_w1500_
	);
	LUT3 #(
		.INIT('hd0)
	) name1038 (
		_w1490_,
		_w1499_,
		_w1500_,
		_w1501_
	);
	LUT2 #(
		.INIT('h8)
	) name1039 (
		_w1425_,
		_w1433_,
		_w1502_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1040 (
		_w1489_,
		_w1497_,
		_w1501_,
		_w1502_,
		_w1503_
	);
	LUT3 #(
		.INIT('ha2)
	) name1041 (
		_w1487_,
		_w1488_,
		_w1503_,
		_w1504_
	);
	LUT4 #(
		.INIT('h9565)
	) name1042 (
		\P1_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w568_,
		_w1504_,
		_w1505_
	);
	LUT2 #(
		.INIT('h1)
	) name1043 (
		_w1306_,
		_w1505_,
		_w1506_
	);
	LUT3 #(
		.INIT('h6c)
	) name1044 (
		\P2_reg3_reg[25]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		_w1394_,
		_w1507_
	);
	LUT3 #(
		.INIT('h08)
	) name1045 (
		\P2_reg2_reg[26]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1508_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1046 (
		\P2_reg0_reg[26]/NET0131 ,
		\P2_reg1_reg[26]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1509_
	);
	LUT4 #(
		.INIT('h1300)
	) name1047 (
		_w1383_,
		_w1508_,
		_w1507_,
		_w1509_,
		_w1510_
	);
	LUT4 #(
		.INIT('hecff)
	) name1048 (
		_w1383_,
		_w1508_,
		_w1507_,
		_w1509_,
		_w1511_
	);
	LUT3 #(
		.INIT('he0)
	) name1049 (
		_w1306_,
		_w1505_,
		_w1510_,
		_w1512_
	);
	LUT4 #(
		.INIT('h0133)
	) name1050 (
		_w1306_,
		_w1485_,
		_w1505_,
		_w1510_,
		_w1513_
	);
	LUT2 #(
		.INIT('h2)
	) name1051 (
		\P1_datao_reg[25]/NET0131 ,
		_w568_,
		_w1514_
	);
	LUT2 #(
		.INIT('h6)
	) name1052 (
		\P1_datao_reg[25]/NET0131 ,
		\si[25]_pad ,
		_w1515_
	);
	LUT4 #(
		.INIT('hb000)
	) name1053 (
		_w1328_,
		_w1333_,
		_w1336_,
		_w1346_,
		_w1516_
	);
	LUT3 #(
		.INIT('h8a)
	) name1054 (
		_w1353_,
		_w1316_,
		_w1346_,
		_w1517_
	);
	LUT4 #(
		.INIT('h2a22)
	) name1055 (
		_w1340_,
		_w1353_,
		_w1316_,
		_w1346_,
		_w1518_
	);
	LUT2 #(
		.INIT('h2)
	) name1056 (
		_w1350_,
		_w1518_,
		_w1519_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1057 (
		_w1362_,
		_w1340_,
		_w1516_,
		_w1519_,
		_w1520_
	);
	LUT4 #(
		.INIT('h0a82)
	) name1058 (
		_w568_,
		_w1369_,
		_w1515_,
		_w1520_,
		_w1521_
	);
	LUT3 #(
		.INIT('h54)
	) name1059 (
		_w1306_,
		_w1514_,
		_w1521_,
		_w1522_
	);
	LUT2 #(
		.INIT('h6)
	) name1060 (
		\P2_reg3_reg[25]/NET0131 ,
		_w1394_,
		_w1523_
	);
	LUT4 #(
		.INIT('h4080)
	) name1061 (
		\P2_reg3_reg[25]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1394_,
		_w1524_
	);
	LUT3 #(
		.INIT('h02)
	) name1062 (
		\P2_reg0_reg[25]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1525_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1063 (
		\P2_reg1_reg[25]/NET0131 ,
		\P2_reg2_reg[25]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1526_
	);
	LUT3 #(
		.INIT('h10)
	) name1064 (
		_w1525_,
		_w1524_,
		_w1526_,
		_w1527_
	);
	LUT3 #(
		.INIT('hef)
	) name1065 (
		_w1525_,
		_w1524_,
		_w1526_,
		_w1528_
	);
	LUT4 #(
		.INIT('hab00)
	) name1066 (
		_w1306_,
		_w1514_,
		_w1521_,
		_w1527_,
		_w1529_
	);
	LUT2 #(
		.INIT('h2)
	) name1067 (
		_w1513_,
		_w1529_,
		_w1530_
	);
	LUT2 #(
		.INIT('h2)
	) name1068 (
		\P1_datao_reg[24]/NET0131 ,
		_w568_,
		_w1531_
	);
	LUT2 #(
		.INIT('h6)
	) name1069 (
		\P1_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w1532_
	);
	LUT4 #(
		.INIT('h208a)
	) name1070 (
		_w568_,
		_w1435_,
		_w1438_,
		_w1532_,
		_w1533_
	);
	LUT3 #(
		.INIT('h54)
	) name1071 (
		_w1306_,
		_w1531_,
		_w1533_,
		_w1534_
	);
	LUT4 #(
		.INIT('h8000)
	) name1072 (
		\P2_reg3_reg[19]/NET0131 ,
		_w1388_,
		_w1389_,
		_w1390_,
		_w1535_
	);
	LUT4 #(
		.INIT('h8000)
	) name1073 (
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		_w1391_,
		_w1535_,
		_w1536_
	);
	LUT3 #(
		.INIT('h32)
	) name1074 (
		\P2_reg3_reg[24]/NET0131 ,
		_w1394_,
		_w1536_,
		_w1537_
	);
	LUT4 #(
		.INIT('h0c08)
	) name1075 (
		\P2_reg3_reg[24]/NET0131 ,
		_w1383_,
		_w1394_,
		_w1536_,
		_w1538_
	);
	LUT3 #(
		.INIT('h20)
	) name1076 (
		\P2_reg1_reg[24]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1539_
	);
	LUT4 #(
		.INIT('hff35)
	) name1077 (
		\P2_reg0_reg[24]/NET0131 ,
		\P2_reg2_reg[24]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1540_
	);
	LUT2 #(
		.INIT('h4)
	) name1078 (
		_w1539_,
		_w1540_,
		_w1541_
	);
	LUT2 #(
		.INIT('h4)
	) name1079 (
		_w1538_,
		_w1541_,
		_w1542_
	);
	LUT2 #(
		.INIT('hb)
	) name1080 (
		_w1538_,
		_w1541_,
		_w1543_
	);
	LUT3 #(
		.INIT('ha2)
	) name1081 (
		_w1470_,
		_w1456_,
		_w1473_,
		_w1544_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1082 (
		_w1472_,
		_w1458_,
		_w1469_,
		_w1544_,
		_w1545_
	);
	LUT4 #(
		.INIT('h9565)
	) name1083 (
		\P1_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w568_,
		_w1545_,
		_w1546_
	);
	LUT2 #(
		.INIT('h1)
	) name1084 (
		_w1306_,
		_w1546_,
		_w1547_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1085 (
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		_w1391_,
		_w1535_,
		_w1548_
	);
	LUT3 #(
		.INIT('h08)
	) name1086 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1549_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1087 (
		\P2_reg0_reg[23]/NET0131 ,
		\P2_reg1_reg[23]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1550_
	);
	LUT4 #(
		.INIT('h1300)
	) name1088 (
		_w1383_,
		_w1549_,
		_w1548_,
		_w1550_,
		_w1551_
	);
	LUT4 #(
		.INIT('hecff)
	) name1089 (
		_w1383_,
		_w1549_,
		_w1548_,
		_w1550_,
		_w1552_
	);
	LUT3 #(
		.INIT('he0)
	) name1090 (
		_w1306_,
		_w1546_,
		_w1551_,
		_w1553_
	);
	LUT3 #(
		.INIT('h0b)
	) name1091 (
		_w1534_,
		_w1542_,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('h2)
	) name1092 (
		\P1_datao_reg[22]/NET0131 ,
		_w568_,
		_w1555_
	);
	LUT2 #(
		.INIT('h6)
	) name1093 (
		\P1_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w1556_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1094 (
		_w1493_,
		_w1495_,
		_w1496_,
		_w1499_,
		_w1557_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1095 (
		_w1490_,
		_w1500_,
		_w1502_,
		_w1557_,
		_w1558_
	);
	LUT4 #(
		.INIT('h0a82)
	) name1096 (
		_w568_,
		_w1489_,
		_w1556_,
		_w1558_,
		_w1559_
	);
	LUT3 #(
		.INIT('h54)
	) name1097 (
		_w1306_,
		_w1555_,
		_w1559_,
		_w1560_
	);
	LUT3 #(
		.INIT('h6a)
	) name1098 (
		\P2_reg3_reg[22]/NET0131 ,
		_w1391_,
		_w1535_,
		_w1561_
	);
	LUT3 #(
		.INIT('h20)
	) name1099 (
		\P2_reg1_reg[22]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1562_
	);
	LUT4 #(
		.INIT('hff35)
	) name1100 (
		\P2_reg0_reg[22]/NET0131 ,
		\P2_reg2_reg[22]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1563_
	);
	LUT4 #(
		.INIT('h1300)
	) name1101 (
		_w1383_,
		_w1562_,
		_w1561_,
		_w1563_,
		_w1564_
	);
	LUT4 #(
		.INIT('hecff)
	) name1102 (
		_w1383_,
		_w1562_,
		_w1561_,
		_w1563_,
		_w1565_
	);
	LUT4 #(
		.INIT('h0054)
	) name1103 (
		_w1306_,
		_w1555_,
		_w1559_,
		_w1564_,
		_w1566_
	);
	LUT4 #(
		.INIT('hab00)
	) name1104 (
		_w1306_,
		_w1555_,
		_w1559_,
		_w1564_,
		_w1567_
	);
	LUT4 #(
		.INIT('h9565)
	) name1105 (
		\P1_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w568_,
		_w1355_,
		_w1568_
	);
	LUT2 #(
		.INIT('h1)
	) name1106 (
		_w1306_,
		_w1568_,
		_w1569_
	);
	LUT3 #(
		.INIT('h6c)
	) name1107 (
		\P2_reg3_reg[20]/NET0131 ,
		\P2_reg3_reg[21]/NET0131 ,
		_w1535_,
		_w1570_
	);
	LUT3 #(
		.INIT('h02)
	) name1108 (
		\P2_reg0_reg[21]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1571_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1109 (
		\P2_reg1_reg[21]/NET0131 ,
		\P2_reg2_reg[21]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1572_
	);
	LUT4 #(
		.INIT('h1300)
	) name1110 (
		_w1383_,
		_w1571_,
		_w1570_,
		_w1572_,
		_w1573_
	);
	LUT4 #(
		.INIT('hecff)
	) name1111 (
		_w1383_,
		_w1571_,
		_w1570_,
		_w1572_,
		_w1574_
	);
	LUT3 #(
		.INIT('h01)
	) name1112 (
		_w1306_,
		_w1568_,
		_w1573_,
		_w1575_
	);
	LUT3 #(
		.INIT('h45)
	) name1113 (
		_w1566_,
		_w1567_,
		_w1575_,
		_w1576_
	);
	LUT3 #(
		.INIT('h01)
	) name1114 (
		_w1306_,
		_w1546_,
		_w1551_,
		_w1577_
	);
	LUT3 #(
		.INIT('h4d)
	) name1115 (
		_w1534_,
		_w1542_,
		_w1577_,
		_w1578_
	);
	LUT3 #(
		.INIT('hd0)
	) name1116 (
		_w1554_,
		_w1576_,
		_w1578_,
		_w1579_
	);
	LUT4 #(
		.INIT('h0054)
	) name1117 (
		_w1306_,
		_w1514_,
		_w1521_,
		_w1527_,
		_w1580_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1118 (
		_w1306_,
		_w1505_,
		_w1510_,
		_w1580_,
		_w1581_
	);
	LUT4 #(
		.INIT('h0054)
	) name1119 (
		_w1306_,
		_w1452_,
		_w1478_,
		_w1483_,
		_w1582_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1120 (
		_w1306_,
		_w1441_,
		_w1449_,
		_w1582_,
		_w1583_
	);
	LUT3 #(
		.INIT('hd0)
	) name1121 (
		_w1513_,
		_w1581_,
		_w1583_,
		_w1584_
	);
	LUT4 #(
		.INIT('h0455)
	) name1122 (
		_w1451_,
		_w1530_,
		_w1579_,
		_w1584_,
		_w1585_
	);
	LUT4 #(
		.INIT('h9565)
	) name1123 (
		\P1_datao_reg[20]/NET0131 ,
		\si[20]_pad ,
		_w568_,
		_w1431_,
		_w1586_
	);
	LUT2 #(
		.INIT('h1)
	) name1124 (
		_w1306_,
		_w1586_,
		_w1587_
	);
	LUT2 #(
		.INIT('h6)
	) name1125 (
		\P2_reg3_reg[20]/NET0131 ,
		_w1535_,
		_w1588_
	);
	LUT4 #(
		.INIT('h4080)
	) name1126 (
		\P2_reg3_reg[20]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1535_,
		_w1589_
	);
	LUT3 #(
		.INIT('h08)
	) name1127 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1590_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1128 (
		\P2_reg0_reg[20]/NET0131 ,
		\P2_reg1_reg[20]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1591_
	);
	LUT3 #(
		.INIT('h10)
	) name1129 (
		_w1590_,
		_w1589_,
		_w1591_,
		_w1592_
	);
	LUT3 #(
		.INIT('hef)
	) name1130 (
		_w1590_,
		_w1589_,
		_w1591_,
		_w1593_
	);
	LUT3 #(
		.INIT('he0)
	) name1131 (
		_w1306_,
		_w1586_,
		_w1592_,
		_w1594_
	);
	LUT2 #(
		.INIT('h6)
	) name1132 (
		\P2_IR_reg[19]/NET0131 ,
		_w1264_,
		_w1595_
	);
	LUT3 #(
		.INIT('h01)
	) name1133 (
		_w1302_,
		_w1305_,
		_w1595_,
		_w1596_
	);
	LUT3 #(
		.INIT('h4c)
	) name1134 (
		_w1457_,
		_w1474_,
		_w1469_,
		_w1597_
	);
	LUT4 #(
		.INIT('h9565)
	) name1135 (
		\P1_datao_reg[19]/NET0131 ,
		\si[19]_pad ,
		_w568_,
		_w1597_,
		_w1598_
	);
	LUT3 #(
		.INIT('h23)
	) name1136 (
		_w1306_,
		_w1596_,
		_w1598_,
		_w1599_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1137 (
		\P2_reg3_reg[19]/NET0131 ,
		_w1388_,
		_w1389_,
		_w1390_,
		_w1600_
	);
	LUT3 #(
		.INIT('h80)
	) name1138 (
		_w1378_,
		_w1382_,
		_w1600_,
		_w1601_
	);
	LUT3 #(
		.INIT('h08)
	) name1139 (
		\P2_reg2_reg[19]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1602_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1140 (
		\P2_reg0_reg[19]/NET0131 ,
		\P2_reg1_reg[19]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1603_
	);
	LUT3 #(
		.INIT('h10)
	) name1141 (
		_w1602_,
		_w1601_,
		_w1603_,
		_w1604_
	);
	LUT3 #(
		.INIT('hef)
	) name1142 (
		_w1602_,
		_w1601_,
		_w1603_,
		_w1605_
	);
	LUT4 #(
		.INIT('hdc00)
	) name1143 (
		_w1306_,
		_w1596_,
		_w1598_,
		_w1604_,
		_w1606_
	);
	LUT4 #(
		.INIT('ha666)
	) name1144 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1262_,
		_w1263_,
		_w1607_
	);
	LUT3 #(
		.INIT('h01)
	) name1145 (
		_w1302_,
		_w1305_,
		_w1607_,
		_w1608_
	);
	LUT2 #(
		.INIT('h2)
	) name1146 (
		\P1_datao_reg[17]/NET0131 ,
		_w568_,
		_w1609_
	);
	LUT2 #(
		.INIT('h6)
	) name1147 (
		\P1_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w1610_
	);
	LUT4 #(
		.INIT('h208a)
	) name1148 (
		_w568_,
		_w1516_,
		_w1517_,
		_w1610_,
		_w1611_
	);
	LUT4 #(
		.INIT('h3332)
	) name1149 (
		_w1306_,
		_w1608_,
		_w1609_,
		_w1611_,
		_w1612_
	);
	LUT3 #(
		.INIT('h6a)
	) name1150 (
		\P2_reg3_reg[17]/NET0131 ,
		_w1388_,
		_w1389_,
		_w1613_
	);
	LUT3 #(
		.INIT('h80)
	) name1151 (
		_w1378_,
		_w1382_,
		_w1613_,
		_w1614_
	);
	LUT3 #(
		.INIT('h02)
	) name1152 (
		\P2_reg0_reg[17]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1615_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1153 (
		\P2_reg1_reg[17]/NET0131 ,
		\P2_reg2_reg[17]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1616_
	);
	LUT3 #(
		.INIT('h10)
	) name1154 (
		_w1615_,
		_w1614_,
		_w1616_,
		_w1617_
	);
	LUT3 #(
		.INIT('hef)
	) name1155 (
		_w1615_,
		_w1614_,
		_w1616_,
		_w1618_
	);
	LUT2 #(
		.INIT('h2)
	) name1156 (
		\P2_IR_reg[31]/NET0131 ,
		_w1269_,
		_w1619_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1157 (
		\P2_IR_reg[31]/NET0131 ,
		_w1261_,
		_w1268_,
		_w1619_,
		_w1620_
	);
	LUT2 #(
		.INIT('h9)
	) name1158 (
		\P2_IR_reg[18]/NET0131 ,
		_w1620_,
		_w1621_
	);
	LUT3 #(
		.INIT('h01)
	) name1159 (
		_w1302_,
		_w1305_,
		_w1621_,
		_w1622_
	);
	LUT2 #(
		.INIT('h2)
	) name1160 (
		\P1_datao_reg[18]/NET0131 ,
		_w568_,
		_w1623_
	);
	LUT2 #(
		.INIT('h6)
	) name1161 (
		\P1_datao_reg[18]/NET0131 ,
		\si[18]_pad ,
		_w1624_
	);
	LUT4 #(
		.INIT('h208a)
	) name1162 (
		_w568_,
		_w1497_,
		_w1501_,
		_w1624_,
		_w1625_
	);
	LUT4 #(
		.INIT('h3332)
	) name1163 (
		_w1306_,
		_w1622_,
		_w1623_,
		_w1625_,
		_w1626_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1164 (
		\P2_reg3_reg[17]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		_w1388_,
		_w1389_,
		_w1627_
	);
	LUT3 #(
		.INIT('h80)
	) name1165 (
		_w1378_,
		_w1382_,
		_w1627_,
		_w1628_
	);
	LUT3 #(
		.INIT('h20)
	) name1166 (
		\P2_reg1_reg[18]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1629_
	);
	LUT4 #(
		.INIT('hff35)
	) name1167 (
		\P2_reg0_reg[18]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1630_
	);
	LUT3 #(
		.INIT('h10)
	) name1168 (
		_w1629_,
		_w1628_,
		_w1630_,
		_w1631_
	);
	LUT3 #(
		.INIT('hef)
	) name1169 (
		_w1629_,
		_w1628_,
		_w1630_,
		_w1632_
	);
	LUT2 #(
		.INIT('h4)
	) name1170 (
		_w1626_,
		_w1631_,
		_w1633_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1171 (
		_w1612_,
		_w1617_,
		_w1626_,
		_w1631_,
		_w1634_
	);
	LUT3 #(
		.INIT('h10)
	) name1172 (
		_w1594_,
		_w1606_,
		_w1634_,
		_w1635_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1173 (
		\P2_reg2_reg[2]/NET0131 ,
		\P2_reg3_reg[2]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1636_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1174 (
		\P2_reg0_reg[2]/NET0131 ,
		\P2_reg1_reg[2]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1637_
	);
	LUT2 #(
		.INIT('h8)
	) name1175 (
		_w1636_,
		_w1637_,
		_w1638_
	);
	LUT2 #(
		.INIT('h7)
	) name1176 (
		_w1636_,
		_w1637_,
		_w1639_
	);
	LUT4 #(
		.INIT('h6595)
	) name1177 (
		\P1_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w568_,
		_w1320_,
		_w1640_
	);
	LUT4 #(
		.INIT('h1ef0)
	) name1178 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[2]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1641_
	);
	LUT3 #(
		.INIT('h10)
	) name1179 (
		_w1302_,
		_w1305_,
		_w1641_,
		_w1642_
	);
	LUT4 #(
		.INIT('he0f1)
	) name1180 (
		_w1302_,
		_w1305_,
		_w1640_,
		_w1641_,
		_w1643_
	);
	LUT3 #(
		.INIT('h07)
	) name1181 (
		_w1636_,
		_w1637_,
		_w1643_,
		_w1644_
	);
	LUT3 #(
		.INIT('h80)
	) name1182 (
		_w1636_,
		_w1637_,
		_w1643_,
		_w1645_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1183 (
		\P2_reg0_reg[1]/NET0131 ,
		\P2_reg1_reg[1]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1646_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1184 (
		\P2_reg2_reg[1]/NET0131 ,
		\P2_reg3_reg[1]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1647_
	);
	LUT2 #(
		.INIT('h8)
	) name1185 (
		_w1646_,
		_w1647_,
		_w1648_
	);
	LUT2 #(
		.INIT('h7)
	) name1186 (
		_w1646_,
		_w1647_,
		_w1649_
	);
	LUT4 #(
		.INIT('h9a6a)
	) name1187 (
		\P1_datao_reg[1]/NET0131 ,
		\si[1]_pad ,
		_w568_,
		_w1319_,
		_w1650_
	);
	LUT3 #(
		.INIT('h93)
	) name1188 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1651_
	);
	LUT3 #(
		.INIT('h01)
	) name1189 (
		_w1302_,
		_w1305_,
		_w1651_,
		_w1652_
	);
	LUT4 #(
		.INIT('h1f0e)
	) name1190 (
		_w1302_,
		_w1305_,
		_w1650_,
		_w1651_,
		_w1653_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1191 (
		\P2_reg1_reg[0]/NET0131 ,
		\P2_reg3_reg[0]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1654_
	);
	LUT4 #(
		.INIT('hff35)
	) name1192 (
		\P2_reg0_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1655_
	);
	LUT2 #(
		.INIT('h8)
	) name1193 (
		_w1654_,
		_w1655_,
		_w1656_
	);
	LUT2 #(
		.INIT('h7)
	) name1194 (
		_w1654_,
		_w1655_,
		_w1657_
	);
	LUT3 #(
		.INIT('h6a)
	) name1195 (
		\P1_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w568_,
		_w1658_
	);
	LUT3 #(
		.INIT('h02)
	) name1196 (
		\P2_IR_reg[0]/NET0131 ,
		_w1302_,
		_w1305_,
		_w1659_
	);
	LUT4 #(
		.INIT('h01fd)
	) name1197 (
		\P2_IR_reg[0]/NET0131 ,
		_w1302_,
		_w1305_,
		_w1658_,
		_w1660_
	);
	LUT3 #(
		.INIT('h07)
	) name1198 (
		_w1654_,
		_w1655_,
		_w1660_,
		_w1661_
	);
	LUT4 #(
		.INIT('h1501)
	) name1199 (
		_w1645_,
		_w1648_,
		_w1653_,
		_w1661_,
		_w1662_
	);
	LUT4 #(
		.INIT('h9a6a)
	) name1200 (
		\P1_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w568_,
		_w1322_,
		_w1663_
	);
	LUT3 #(
		.INIT('h39)
	) name1201 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		_w1259_,
		_w1664_
	);
	LUT3 #(
		.INIT('h01)
	) name1202 (
		_w1302_,
		_w1305_,
		_w1664_,
		_w1665_
	);
	LUT4 #(
		.INIT('h1f0e)
	) name1203 (
		_w1302_,
		_w1305_,
		_w1663_,
		_w1664_,
		_w1666_
	);
	LUT4 #(
		.INIT('hff35)
	) name1204 (
		\P2_reg0_reg[4]/NET0131 ,
		\P2_reg2_reg[4]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1667_
	);
	LUT2 #(
		.INIT('h6)
	) name1205 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		_w1668_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1206 (
		\P2_reg1_reg[4]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1668_,
		_w1669_
	);
	LUT2 #(
		.INIT('h8)
	) name1207 (
		_w1667_,
		_w1669_,
		_w1670_
	);
	LUT2 #(
		.INIT('h7)
	) name1208 (
		_w1667_,
		_w1669_,
		_w1671_
	);
	LUT3 #(
		.INIT('h80)
	) name1209 (
		_w1666_,
		_w1667_,
		_w1669_,
		_w1672_
	);
	LUT4 #(
		.INIT('hff35)
	) name1210 (
		\P2_reg0_reg[3]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1673_
	);
	LUT4 #(
		.INIT('hc5ff)
	) name1211 (
		\P2_reg1_reg[3]/NET0131 ,
		\P2_reg3_reg[3]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1674_
	);
	LUT2 #(
		.INIT('h8)
	) name1212 (
		_w1673_,
		_w1674_,
		_w1675_
	);
	LUT2 #(
		.INIT('h7)
	) name1213 (
		_w1673_,
		_w1674_,
		_w1676_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1214 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[2]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1677_
	);
	LUT2 #(
		.INIT('h6)
	) name1215 (
		\P2_IR_reg[3]/NET0131 ,
		_w1677_,
		_w1678_
	);
	LUT3 #(
		.INIT('h10)
	) name1216 (
		_w1302_,
		_w1305_,
		_w1678_,
		_w1679_
	);
	LUT4 #(
		.INIT('h9565)
	) name1217 (
		\P1_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w568_,
		_w1459_,
		_w1680_
	);
	LUT4 #(
		.INIT('hef01)
	) name1218 (
		_w1302_,
		_w1305_,
		_w1678_,
		_w1680_,
		_w1681_
	);
	LUT3 #(
		.INIT('h80)
	) name1219 (
		_w1673_,
		_w1674_,
		_w1681_,
		_w1682_
	);
	LUT2 #(
		.INIT('h1)
	) name1220 (
		_w1672_,
		_w1682_,
		_w1683_
	);
	LUT3 #(
		.INIT('h15)
	) name1221 (
		_w1666_,
		_w1667_,
		_w1669_,
		_w1684_
	);
	LUT3 #(
		.INIT('h07)
	) name1222 (
		_w1673_,
		_w1674_,
		_w1681_,
		_w1685_
	);
	LUT3 #(
		.INIT('h23)
	) name1223 (
		_w1672_,
		_w1684_,
		_w1685_,
		_w1686_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1224 (
		_w1644_,
		_w1662_,
		_w1683_,
		_w1686_,
		_w1687_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1225 (
		\P2_reg0_reg[8]/NET0131 ,
		\P2_reg1_reg[8]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1688_
	);
	LUT3 #(
		.INIT('h6c)
	) name1226 (
		\P2_reg3_reg[7]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		_w1384_,
		_w1689_
	);
	LUT4 #(
		.INIT('h37f7)
	) name1227 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1689_,
		_w1690_
	);
	LUT2 #(
		.INIT('h8)
	) name1228 (
		_w1688_,
		_w1690_,
		_w1691_
	);
	LUT2 #(
		.INIT('h7)
	) name1229 (
		_w1688_,
		_w1690_,
		_w1692_
	);
	LUT4 #(
		.INIT('hc666)
	) name1230 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		_w1259_,
		_w1260_,
		_w1693_
	);
	LUT4 #(
		.INIT('h9565)
	) name1231 (
		\P1_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w568_,
		_w1413_,
		_w1694_
	);
	LUT4 #(
		.INIT('h10fe)
	) name1232 (
		_w1302_,
		_w1305_,
		_w1693_,
		_w1694_,
		_w1695_
	);
	LUT3 #(
		.INIT('h08)
	) name1233 (
		_w1688_,
		_w1690_,
		_w1695_,
		_w1696_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1234 (
		\P2_reg1_reg[7]/NET0131 ,
		\P2_reg2_reg[7]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1697_
	);
	LUT2 #(
		.INIT('h6)
	) name1235 (
		\P2_reg3_reg[7]/NET0131 ,
		_w1384_,
		_w1698_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1236 (
		\P2_reg0_reg[7]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1698_,
		_w1699_
	);
	LUT2 #(
		.INIT('h8)
	) name1237 (
		_w1697_,
		_w1699_,
		_w1700_
	);
	LUT2 #(
		.INIT('h7)
	) name1238 (
		_w1697_,
		_w1699_,
		_w1701_
	);
	LUT3 #(
		.INIT('ha8)
	) name1239 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[5]/NET0131 ,
		\P2_IR_reg[6]/NET0131 ,
		_w1702_
	);
	LUT4 #(
		.INIT('h0075)
	) name1240 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		_w1259_,
		_w1702_,
		_w1703_
	);
	LUT2 #(
		.INIT('h9)
	) name1241 (
		\P2_IR_reg[7]/NET0131 ,
		_w1703_,
		_w1704_
	);
	LUT4 #(
		.INIT('h9565)
	) name1242 (
		\P1_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w568_,
		_w1463_,
		_w1705_
	);
	LUT4 #(
		.INIT('h10fe)
	) name1243 (
		_w1302_,
		_w1305_,
		_w1704_,
		_w1705_,
		_w1706_
	);
	LUT3 #(
		.INIT('h08)
	) name1244 (
		_w1697_,
		_w1699_,
		_w1706_,
		_w1707_
	);
	LUT2 #(
		.INIT('h1)
	) name1245 (
		_w1696_,
		_w1707_,
		_w1708_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1246 (
		\P2_reg1_reg[6]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1709_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1247 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		\P2_reg3_reg[6]/NET0131 ,
		_w1710_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1248 (
		\P2_reg0_reg[6]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1710_,
		_w1711_
	);
	LUT2 #(
		.INIT('h8)
	) name1249 (
		_w1709_,
		_w1711_,
		_w1712_
	);
	LUT2 #(
		.INIT('h7)
	) name1250 (
		_w1709_,
		_w1711_,
		_w1713_
	);
	LUT4 #(
		.INIT('h5755)
	) name1251 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_IR_reg[5]/NET0131 ,
		_w1259_,
		_w1714_
	);
	LUT2 #(
		.INIT('h9)
	) name1252 (
		\P2_IR_reg[6]/NET0131 ,
		_w1714_,
		_w1715_
	);
	LUT4 #(
		.INIT('h9565)
	) name1253 (
		\P1_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w568_,
		_w1491_,
		_w1716_
	);
	LUT4 #(
		.INIT('h10fe)
	) name1254 (
		_w1302_,
		_w1305_,
		_w1715_,
		_w1716_,
		_w1717_
	);
	LUT3 #(
		.INIT('h08)
	) name1255 (
		_w1709_,
		_w1711_,
		_w1717_,
		_w1718_
	);
	LUT3 #(
		.INIT('h78)
	) name1256 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		_w1719_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1257 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1719_,
		_w1720_
	);
	LUT4 #(
		.INIT('hff35)
	) name1258 (
		\P2_reg0_reg[5]/NET0131 ,
		\P2_reg2_reg[5]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1721_
	);
	LUT2 #(
		.INIT('h8)
	) name1259 (
		_w1720_,
		_w1721_,
		_w1722_
	);
	LUT2 #(
		.INIT('h7)
	) name1260 (
		_w1720_,
		_w1721_,
		_w1723_
	);
	LUT4 #(
		.INIT('h87a5)
	) name1261 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_IR_reg[5]/NET0131 ,
		_w1259_,
		_w1724_
	);
	LUT4 #(
		.INIT('h6595)
	) name1262 (
		\P1_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w568_,
		_w1323_,
		_w1725_
	);
	LUT4 #(
		.INIT('h01ef)
	) name1263 (
		_w1302_,
		_w1305_,
		_w1724_,
		_w1725_,
		_w1726_
	);
	LUT3 #(
		.INIT('h08)
	) name1264 (
		_w1720_,
		_w1721_,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('h1)
	) name1265 (
		_w1718_,
		_w1727_,
		_w1728_
	);
	LUT4 #(
		.INIT('h0001)
	) name1266 (
		_w1696_,
		_w1707_,
		_w1718_,
		_w1727_,
		_w1729_
	);
	LUT3 #(
		.INIT('h70)
	) name1267 (
		_w1709_,
		_w1711_,
		_w1717_,
		_w1730_
	);
	LUT3 #(
		.INIT('h70)
	) name1268 (
		_w1720_,
		_w1721_,
		_w1726_,
		_w1731_
	);
	LUT3 #(
		.INIT('h23)
	) name1269 (
		_w1718_,
		_w1730_,
		_w1731_,
		_w1732_
	);
	LUT3 #(
		.INIT('h70)
	) name1270 (
		_w1688_,
		_w1690_,
		_w1695_,
		_w1733_
	);
	LUT3 #(
		.INIT('h70)
	) name1271 (
		_w1697_,
		_w1699_,
		_w1706_,
		_w1734_
	);
	LUT3 #(
		.INIT('h54)
	) name1272 (
		_w1696_,
		_w1733_,
		_w1734_,
		_w1735_
	);
	LUT3 #(
		.INIT('h0d)
	) name1273 (
		_w1708_,
		_w1732_,
		_w1735_,
		_w1736_
	);
	LUT3 #(
		.INIT('h6c)
	) name1274 (
		\P2_reg3_reg[10]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		_w1385_,
		_w1737_
	);
	LUT4 #(
		.INIT('h37f7)
	) name1275 (
		\P2_reg2_reg[11]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1737_,
		_w1738_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1276 (
		\P2_reg0_reg[11]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1739_
	);
	LUT2 #(
		.INIT('h8)
	) name1277 (
		_w1738_,
		_w1739_,
		_w1740_
	);
	LUT2 #(
		.INIT('h7)
	) name1278 (
		_w1738_,
		_w1739_,
		_w1741_
	);
	LUT4 #(
		.INIT('hccc8)
	) name1279 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w1742_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1280 (
		\P2_IR_reg[31]/NET0131 ,
		_w1259_,
		_w1260_,
		_w1742_,
		_w1743_
	);
	LUT2 #(
		.INIT('h9)
	) name1281 (
		\P2_IR_reg[11]/NET0131 ,
		_w1743_,
		_w1744_
	);
	LUT3 #(
		.INIT('h01)
	) name1282 (
		_w1302_,
		_w1305_,
		_w1744_,
		_w1745_
	);
	LUT4 #(
		.INIT('h9565)
	) name1283 (
		\P1_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w568_,
		_w1467_,
		_w1746_
	);
	LUT3 #(
		.INIT('h23)
	) name1284 (
		_w1306_,
		_w1745_,
		_w1746_,
		_w1747_
	);
	LUT4 #(
		.INIT('h8000)
	) name1285 (
		\P2_reg3_reg[10]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		_w1385_,
		_w1748_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1286 (
		\P2_reg3_reg[10]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		_w1385_,
		_w1749_
	);
	LUT4 #(
		.INIT('h37f7)
	) name1287 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1749_,
		_w1750_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1288 (
		\P2_reg0_reg[12]/NET0131 ,
		\P2_reg1_reg[12]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1751_
	);
	LUT2 #(
		.INIT('h8)
	) name1289 (
		_w1750_,
		_w1751_,
		_w1752_
	);
	LUT2 #(
		.INIT('h7)
	) name1290 (
		_w1750_,
		_w1751_,
		_w1753_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1291 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1259_,
		_w1260_,
		_w1754_
	);
	LUT3 #(
		.INIT('h56)
	) name1292 (
		\P2_IR_reg[12]/NET0131 ,
		_w1742_,
		_w1754_,
		_w1755_
	);
	LUT3 #(
		.INIT('h01)
	) name1293 (
		_w1302_,
		_w1305_,
		_w1755_,
		_w1756_
	);
	LUT3 #(
		.INIT('hb0)
	) name1294 (
		_w1413_,
		_w1416_,
		_w1418_,
		_w1757_
	);
	LUT4 #(
		.INIT('h9565)
	) name1295 (
		\P1_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w568_,
		_w1757_,
		_w1758_
	);
	LUT3 #(
		.INIT('h23)
	) name1296 (
		_w1306_,
		_w1756_,
		_w1758_,
		_w1759_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1297 (
		_w1740_,
		_w1747_,
		_w1752_,
		_w1759_,
		_w1760_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1298 (
		\P2_reg0_reg[10]/NET0131 ,
		\P2_reg1_reg[10]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1761_
	);
	LUT2 #(
		.INIT('h6)
	) name1299 (
		\P2_reg3_reg[10]/NET0131 ,
		_w1385_,
		_w1762_
	);
	LUT4 #(
		.INIT('h37f7)
	) name1300 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1762_,
		_w1763_
	);
	LUT2 #(
		.INIT('h8)
	) name1301 (
		_w1761_,
		_w1763_,
		_w1764_
	);
	LUT2 #(
		.INIT('h7)
	) name1302 (
		_w1761_,
		_w1763_,
		_w1765_
	);
	LUT3 #(
		.INIT('ha8)
	) name1303 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w1766_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1304 (
		\P2_IR_reg[31]/NET0131 ,
		_w1259_,
		_w1260_,
		_w1766_,
		_w1767_
	);
	LUT2 #(
		.INIT('h9)
	) name1305 (
		\P2_IR_reg[10]/NET0131 ,
		_w1767_,
		_w1768_
	);
	LUT3 #(
		.INIT('h01)
	) name1306 (
		_w1302_,
		_w1305_,
		_w1768_,
		_w1769_
	);
	LUT2 #(
		.INIT('h2)
	) name1307 (
		\P1_datao_reg[10]/NET0131 ,
		_w568_,
		_w1770_
	);
	LUT2 #(
		.INIT('h6)
	) name1308 (
		\P1_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w1771_
	);
	LUT4 #(
		.INIT('h208a)
	) name1309 (
		_w568_,
		_w1493_,
		_w1495_,
		_w1771_,
		_w1772_
	);
	LUT4 #(
		.INIT('h000e)
	) name1310 (
		_w1302_,
		_w1305_,
		_w1770_,
		_w1772_,
		_w1773_
	);
	LUT2 #(
		.INIT('h1)
	) name1311 (
		_w1769_,
		_w1773_,
		_w1774_
	);
	LUT4 #(
		.INIT('h8880)
	) name1312 (
		_w1761_,
		_w1763_,
		_w1769_,
		_w1773_,
		_w1775_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1313 (
		\P2_reg3_reg[7]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		\P2_reg3_reg[9]/NET0131 ,
		_w1384_,
		_w1776_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1314 (
		\P2_reg1_reg[9]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1776_,
		_w1777_
	);
	LUT4 #(
		.INIT('hff35)
	) name1315 (
		\P2_reg0_reg[9]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1778_
	);
	LUT2 #(
		.INIT('h8)
	) name1316 (
		_w1777_,
		_w1778_,
		_w1779_
	);
	LUT2 #(
		.INIT('h7)
	) name1317 (
		_w1777_,
		_w1778_,
		_w1780_
	);
	LUT4 #(
		.INIT('h7555)
	) name1318 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		_w1259_,
		_w1260_,
		_w1781_
	);
	LUT2 #(
		.INIT('h9)
	) name1319 (
		\P2_IR_reg[9]/NET0131 ,
		_w1781_,
		_w1782_
	);
	LUT3 #(
		.INIT('h01)
	) name1320 (
		_w1302_,
		_w1305_,
		_w1782_,
		_w1783_
	);
	LUT2 #(
		.INIT('h2)
	) name1321 (
		\P1_datao_reg[9]/NET0131 ,
		_w568_,
		_w1784_
	);
	LUT2 #(
		.INIT('h6)
	) name1322 (
		\P1_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w1785_
	);
	LUT4 #(
		.INIT('h208a)
	) name1323 (
		_w568_,
		_w1328_,
		_w1333_,
		_w1785_,
		_w1786_
	);
	LUT4 #(
		.INIT('h000e)
	) name1324 (
		_w1302_,
		_w1305_,
		_w1784_,
		_w1786_,
		_w1787_
	);
	LUT2 #(
		.INIT('h1)
	) name1325 (
		_w1783_,
		_w1787_,
		_w1788_
	);
	LUT4 #(
		.INIT('h8880)
	) name1326 (
		_w1777_,
		_w1778_,
		_w1783_,
		_w1787_,
		_w1789_
	);
	LUT2 #(
		.INIT('h1)
	) name1327 (
		_w1775_,
		_w1789_,
		_w1790_
	);
	LUT2 #(
		.INIT('h8)
	) name1328 (
		_w1760_,
		_w1790_,
		_w1791_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1329 (
		_w1687_,
		_w1729_,
		_w1736_,
		_w1791_,
		_w1792_
	);
	LUT4 #(
		.INIT('h0007)
	) name1330 (
		_w1761_,
		_w1763_,
		_w1769_,
		_w1773_,
		_w1793_
	);
	LUT4 #(
		.INIT('h0007)
	) name1331 (
		_w1777_,
		_w1778_,
		_w1783_,
		_w1787_,
		_w1794_
	);
	LUT3 #(
		.INIT('h23)
	) name1332 (
		_w1775_,
		_w1793_,
		_w1794_,
		_w1795_
	);
	LUT4 #(
		.INIT('h4f04)
	) name1333 (
		_w1740_,
		_w1747_,
		_w1752_,
		_w1759_,
		_w1796_
	);
	LUT3 #(
		.INIT('h0d)
	) name1334 (
		_w1760_,
		_w1795_,
		_w1796_,
		_w1797_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1335 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1798_
	);
	LUT4 #(
		.INIT('h55a6)
	) name1336 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1262_,
		_w1798_,
		_w1799_
	);
	LUT3 #(
		.INIT('h01)
	) name1337 (
		_w1302_,
		_w1305_,
		_w1799_,
		_w1800_
	);
	LUT4 #(
		.INIT('h9565)
	) name1338 (
		\P1_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w568_,
		_w1424_,
		_w1801_
	);
	LUT3 #(
		.INIT('h23)
	) name1339 (
		_w1306_,
		_w1800_,
		_w1801_,
		_w1802_
	);
	LUT3 #(
		.INIT('h6c)
	) name1340 (
		\P2_reg3_reg[15]/NET0131 ,
		\P2_reg3_reg[16]/NET0131 ,
		_w1388_,
		_w1803_
	);
	LUT3 #(
		.INIT('h80)
	) name1341 (
		_w1378_,
		_w1382_,
		_w1803_,
		_w1804_
	);
	LUT3 #(
		.INIT('h20)
	) name1342 (
		\P2_reg1_reg[16]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1805_
	);
	LUT4 #(
		.INIT('hff35)
	) name1343 (
		\P2_reg0_reg[16]/NET0131 ,
		\P2_reg2_reg[16]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1806_
	);
	LUT3 #(
		.INIT('h10)
	) name1344 (
		_w1805_,
		_w1804_,
		_w1806_,
		_w1807_
	);
	LUT3 #(
		.INIT('hef)
	) name1345 (
		_w1805_,
		_w1804_,
		_w1806_,
		_w1808_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1346 (
		\P2_reg0_reg[15]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1809_
	);
	LUT2 #(
		.INIT('h6)
	) name1347 (
		\P2_reg3_reg[15]/NET0131 ,
		_w1388_,
		_w1810_
	);
	LUT4 #(
		.INIT('h37f7)
	) name1348 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1810_,
		_w1811_
	);
	LUT2 #(
		.INIT('h8)
	) name1349 (
		_w1809_,
		_w1811_,
		_w1812_
	);
	LUT2 #(
		.INIT('h7)
	) name1350 (
		_w1809_,
		_w1811_,
		_w1813_
	);
	LUT4 #(
		.INIT('h7333)
	) name1351 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1261_,
		_w1268_,
		_w1814_
	);
	LUT2 #(
		.INIT('h9)
	) name1352 (
		\P2_IR_reg[15]/NET0131 ,
		_w1814_,
		_w1815_
	);
	LUT3 #(
		.INIT('h01)
	) name1353 (
		_w1302_,
		_w1305_,
		_w1815_,
		_w1816_
	);
	LUT2 #(
		.INIT('h2)
	) name1354 (
		\P1_datao_reg[15]/NET0131 ,
		_w568_,
		_w1817_
	);
	LUT2 #(
		.INIT('h6)
	) name1355 (
		\P1_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w1818_
	);
	LUT4 #(
		.INIT('h08a2)
	) name1356 (
		_w568_,
		_w1472_,
		_w1469_,
		_w1818_,
		_w1819_
	);
	LUT4 #(
		.INIT('h3332)
	) name1357 (
		_w1306_,
		_w1816_,
		_w1817_,
		_w1819_,
		_w1820_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name1358 (
		_w1802_,
		_w1807_,
		_w1812_,
		_w1820_,
		_w1821_
	);
	LUT4 #(
		.INIT('hff35)
	) name1359 (
		\P2_reg0_reg[14]/NET0131 ,
		\P2_reg2_reg[14]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1822_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1360 (
		\P2_reg3_reg[10]/NET0131 ,
		\P2_reg3_reg[14]/NET0131 ,
		_w1385_,
		_w1386_,
		_w1823_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1361 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1823_,
		_w1824_
	);
	LUT2 #(
		.INIT('h8)
	) name1362 (
		_w1822_,
		_w1824_,
		_w1825_
	);
	LUT2 #(
		.INIT('h7)
	) name1363 (
		_w1822_,
		_w1824_,
		_w1826_
	);
	LUT4 #(
		.INIT('ha666)
	) name1364 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1261_,
		_w1268_,
		_w1827_
	);
	LUT3 #(
		.INIT('h01)
	) name1365 (
		_w1302_,
		_w1305_,
		_w1827_,
		_w1828_
	);
	LUT4 #(
		.INIT('h9565)
	) name1366 (
		\P1_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w568_,
		_w1557_,
		_w1829_
	);
	LUT3 #(
		.INIT('h23)
	) name1367 (
		_w1306_,
		_w1828_,
		_w1829_,
		_w1830_
	);
	LUT3 #(
		.INIT('h32)
	) name1368 (
		\P2_reg3_reg[13]/NET0131 ,
		_w1387_,
		_w1748_,
		_w1831_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1369 (
		\P2_reg0_reg[13]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1831_,
		_w1832_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1370 (
		\P2_reg1_reg[13]/NET0131 ,
		\P2_reg2_reg[13]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1833_
	);
	LUT2 #(
		.INIT('h8)
	) name1371 (
		_w1832_,
		_w1833_,
		_w1834_
	);
	LUT2 #(
		.INIT('h7)
	) name1372 (
		_w1832_,
		_w1833_,
		_w1835_
	);
	LUT3 #(
		.INIT('h59)
	) name1373 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1262_,
		_w1836_
	);
	LUT3 #(
		.INIT('h10)
	) name1374 (
		_w1302_,
		_w1305_,
		_w1836_,
		_w1837_
	);
	LUT4 #(
		.INIT('h9565)
	) name1375 (
		\P1_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w568_,
		_w1337_,
		_w1838_
	);
	LUT3 #(
		.INIT('h23)
	) name1376 (
		_w1306_,
		_w1837_,
		_w1838_,
		_w1839_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1377 (
		_w1825_,
		_w1830_,
		_w1834_,
		_w1839_,
		_w1840_
	);
	LUT2 #(
		.INIT('h8)
	) name1378 (
		_w1821_,
		_w1840_,
		_w1841_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1379 (
		_w1635_,
		_w1792_,
		_w1797_,
		_w1841_,
		_w1842_
	);
	LUT4 #(
		.INIT('h4d44)
	) name1380 (
		_w1825_,
		_w1830_,
		_w1834_,
		_w1839_,
		_w1843_
	);
	LUT4 #(
		.INIT('hd4dd)
	) name1381 (
		_w1802_,
		_w1807_,
		_w1812_,
		_w1820_,
		_w1844_
	);
	LUT3 #(
		.INIT('h70)
	) name1382 (
		_w1821_,
		_w1843_,
		_w1844_,
		_w1845_
	);
	LUT2 #(
		.INIT('h2)
	) name1383 (
		_w1626_,
		_w1631_,
		_w1846_
	);
	LUT4 #(
		.INIT('h20f2)
	) name1384 (
		_w1612_,
		_w1617_,
		_w1626_,
		_w1631_,
		_w1847_
	);
	LUT3 #(
		.INIT('h10)
	) name1385 (
		_w1594_,
		_w1606_,
		_w1847_,
		_w1848_
	);
	LUT3 #(
		.INIT('h01)
	) name1386 (
		_w1306_,
		_w1586_,
		_w1592_,
		_w1849_
	);
	LUT4 #(
		.INIT('h0023)
	) name1387 (
		_w1306_,
		_w1596_,
		_w1598_,
		_w1604_,
		_w1850_
	);
	LUT3 #(
		.INIT('h23)
	) name1388 (
		_w1594_,
		_w1849_,
		_w1850_,
		_w1851_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1389 (
		_w1635_,
		_w1845_,
		_w1848_,
		_w1851_,
		_w1852_
	);
	LUT3 #(
		.INIT('he0)
	) name1390 (
		_w1306_,
		_w1568_,
		_w1573_,
		_w1853_
	);
	LUT2 #(
		.INIT('h1)
	) name1391 (
		_w1567_,
		_w1853_,
		_w1854_
	);
	LUT3 #(
		.INIT('h40)
	) name1392 (
		_w1451_,
		_w1554_,
		_w1854_,
		_w1855_
	);
	LUT2 #(
		.INIT('h8)
	) name1393 (
		_w1530_,
		_w1855_,
		_w1856_
	);
	LUT4 #(
		.INIT('h1055)
	) name1394 (
		_w1585_,
		_w1842_,
		_w1852_,
		_w1856_,
		_w1857_
	);
	LUT4 #(
		.INIT('hd11d)
	) name1395 (
		\P2_reg2_reg[29]/NET0131 ,
		_w1298_,
		_w1404_,
		_w1857_,
		_w1858_
	);
	LUT2 #(
		.INIT('h6)
	) name1396 (
		\P2_IR_reg[20]/NET0131 ,
		_w1272_,
		_w1859_
	);
	LUT4 #(
		.INIT('h0001)
	) name1397 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_IR_reg[18]/NET0131 ,
		\P2_IR_reg[19]/NET0131 ,
		\P2_IR_reg[20]/NET0131 ,
		_w1860_
	);
	LUT2 #(
		.INIT('h2)
	) name1398 (
		\P2_IR_reg[31]/NET0131 ,
		_w1860_,
		_w1861_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1399 (
		\P2_IR_reg[31]/NET0131 ,
		_w1262_,
		_w1263_,
		_w1861_,
		_w1862_
	);
	LUT2 #(
		.INIT('h9)
	) name1400 (
		\P2_IR_reg[21]/NET0131 ,
		_w1862_,
		_w1863_
	);
	LUT4 #(
		.INIT('h4812)
	) name1401 (
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		_w1272_,
		_w1862_,
		_w1864_
	);
	LUT3 #(
		.INIT('he0)
	) name1402 (
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1865_
	);
	LUT3 #(
		.INIT('h56)
	) name1403 (
		\P2_IR_reg[22]/NET0131 ,
		_w1272_,
		_w1865_,
		_w1866_
	);
	LUT2 #(
		.INIT('h8)
	) name1404 (
		_w1863_,
		_w1866_,
		_w1867_
	);
	LUT2 #(
		.INIT('h1)
	) name1405 (
		_w1863_,
		_w1866_,
		_w1868_
	);
	LUT4 #(
		.INIT('h0530)
	) name1406 (
		_w1595_,
		_w1859_,
		_w1863_,
		_w1866_,
		_w1869_
	);
	LUT2 #(
		.INIT('h4)
	) name1407 (
		_w1858_,
		_w1869_,
		_w1870_
	);
	LUT4 #(
		.INIT('h0777)
	) name1408 (
		_w1740_,
		_w1747_,
		_w1752_,
		_w1759_,
		_w1871_
	);
	LUT4 #(
		.INIT('h0008)
	) name1409 (
		_w1761_,
		_w1763_,
		_w1769_,
		_w1773_,
		_w1872_
	);
	LUT4 #(
		.INIT('h7770)
	) name1410 (
		_w1761_,
		_w1763_,
		_w1769_,
		_w1773_,
		_w1873_
	);
	LUT4 #(
		.INIT('h7770)
	) name1411 (
		_w1777_,
		_w1778_,
		_w1783_,
		_w1787_,
		_w1874_
	);
	LUT3 #(
		.INIT('h54)
	) name1412 (
		_w1872_,
		_w1873_,
		_w1874_,
		_w1875_
	);
	LUT2 #(
		.INIT('h1)
	) name1413 (
		_w1740_,
		_w1747_,
		_w1876_
	);
	LUT4 #(
		.INIT('hfee0)
	) name1414 (
		_w1740_,
		_w1747_,
		_w1752_,
		_w1759_,
		_w1877_
	);
	LUT3 #(
		.INIT('h70)
	) name1415 (
		_w1871_,
		_w1875_,
		_w1877_,
		_w1878_
	);
	LUT3 #(
		.INIT('h80)
	) name1416 (
		_w1688_,
		_w1690_,
		_w1695_,
		_w1879_
	);
	LUT3 #(
		.INIT('h80)
	) name1417 (
		_w1697_,
		_w1699_,
		_w1706_,
		_w1880_
	);
	LUT2 #(
		.INIT('h1)
	) name1418 (
		_w1879_,
		_w1880_,
		_w1881_
	);
	LUT3 #(
		.INIT('h08)
	) name1419 (
		_w1654_,
		_w1655_,
		_w1660_,
		_w1882_
	);
	LUT3 #(
		.INIT('h70)
	) name1420 (
		_w1636_,
		_w1637_,
		_w1643_,
		_w1883_
	);
	LUT4 #(
		.INIT('h00b2)
	) name1421 (
		_w1648_,
		_w1653_,
		_w1882_,
		_w1883_,
		_w1884_
	);
	LUT3 #(
		.INIT('h40)
	) name1422 (
		_w1666_,
		_w1667_,
		_w1669_,
		_w1885_
	);
	LUT3 #(
		.INIT('h08)
	) name1423 (
		_w1673_,
		_w1674_,
		_w1681_,
		_w1886_
	);
	LUT3 #(
		.INIT('h08)
	) name1424 (
		_w1636_,
		_w1637_,
		_w1643_,
		_w1887_
	);
	LUT2 #(
		.INIT('h1)
	) name1425 (
		_w1886_,
		_w1887_,
		_w1888_
	);
	LUT3 #(
		.INIT('h01)
	) name1426 (
		_w1885_,
		_w1886_,
		_w1887_,
		_w1889_
	);
	LUT3 #(
		.INIT('h2a)
	) name1427 (
		_w1666_,
		_w1667_,
		_w1669_,
		_w1890_
	);
	LUT3 #(
		.INIT('h70)
	) name1428 (
		_w1673_,
		_w1674_,
		_w1681_,
		_w1891_
	);
	LUT2 #(
		.INIT('h1)
	) name1429 (
		_w1890_,
		_w1891_,
		_w1892_
	);
	LUT3 #(
		.INIT('h54)
	) name1430 (
		_w1885_,
		_w1890_,
		_w1891_,
		_w1893_
	);
	LUT3 #(
		.INIT('h80)
	) name1431 (
		_w1709_,
		_w1711_,
		_w1717_,
		_w1894_
	);
	LUT3 #(
		.INIT('h80)
	) name1432 (
		_w1720_,
		_w1721_,
		_w1726_,
		_w1895_
	);
	LUT2 #(
		.INIT('h1)
	) name1433 (
		_w1894_,
		_w1895_,
		_w1896_
	);
	LUT4 #(
		.INIT('hf400)
	) name1434 (
		_w1884_,
		_w1889_,
		_w1893_,
		_w1896_,
		_w1897_
	);
	LUT3 #(
		.INIT('h07)
	) name1435 (
		_w1709_,
		_w1711_,
		_w1717_,
		_w1898_
	);
	LUT3 #(
		.INIT('h07)
	) name1436 (
		_w1720_,
		_w1721_,
		_w1726_,
		_w1899_
	);
	LUT2 #(
		.INIT('h1)
	) name1437 (
		_w1898_,
		_w1899_,
		_w1900_
	);
	LUT3 #(
		.INIT('h54)
	) name1438 (
		_w1894_,
		_w1898_,
		_w1899_,
		_w1901_
	);
	LUT3 #(
		.INIT('h07)
	) name1439 (
		_w1688_,
		_w1690_,
		_w1695_,
		_w1902_
	);
	LUT3 #(
		.INIT('h07)
	) name1440 (
		_w1697_,
		_w1699_,
		_w1706_,
		_w1903_
	);
	LUT3 #(
		.INIT('h54)
	) name1441 (
		_w1879_,
		_w1902_,
		_w1903_,
		_w1904_
	);
	LUT4 #(
		.INIT('h0057)
	) name1442 (
		_w1881_,
		_w1897_,
		_w1901_,
		_w1904_,
		_w1905_
	);
	LUT4 #(
		.INIT('h0008)
	) name1443 (
		_w1777_,
		_w1778_,
		_w1783_,
		_w1787_,
		_w1906_
	);
	LUT2 #(
		.INIT('h1)
	) name1444 (
		_w1872_,
		_w1906_,
		_w1907_
	);
	LUT2 #(
		.INIT('h8)
	) name1445 (
		_w1871_,
		_w1907_,
		_w1908_
	);
	LUT3 #(
		.INIT('h10)
	) name1446 (
		_w1306_,
		_w1586_,
		_w1592_,
		_w1909_
	);
	LUT4 #(
		.INIT('h2300)
	) name1447 (
		_w1306_,
		_w1596_,
		_w1598_,
		_w1604_,
		_w1910_
	);
	LUT2 #(
		.INIT('h8)
	) name1448 (
		_w1626_,
		_w1631_,
		_w1911_
	);
	LUT4 #(
		.INIT('h0777)
	) name1449 (
		_w1612_,
		_w1617_,
		_w1626_,
		_w1631_,
		_w1912_
	);
	LUT3 #(
		.INIT('h10)
	) name1450 (
		_w1909_,
		_w1910_,
		_w1912_,
		_w1913_
	);
	LUT4 #(
		.INIT('h0777)
	) name1451 (
		_w1802_,
		_w1807_,
		_w1812_,
		_w1820_,
		_w1914_
	);
	LUT4 #(
		.INIT('h0777)
	) name1452 (
		_w1825_,
		_w1830_,
		_w1834_,
		_w1839_,
		_w1915_
	);
	LUT2 #(
		.INIT('h8)
	) name1453 (
		_w1914_,
		_w1915_,
		_w1916_
	);
	LUT2 #(
		.INIT('h8)
	) name1454 (
		_w1913_,
		_w1916_,
		_w1917_
	);
	LUT4 #(
		.INIT('h7500)
	) name1455 (
		_w1878_,
		_w1905_,
		_w1908_,
		_w1917_,
		_w1918_
	);
	LUT4 #(
		.INIT('heee0)
	) name1456 (
		_w1825_,
		_w1830_,
		_w1834_,
		_w1839_,
		_w1919_
	);
	LUT4 #(
		.INIT('h1117)
	) name1457 (
		_w1825_,
		_w1830_,
		_w1834_,
		_w1839_,
		_w1920_
	);
	LUT2 #(
		.INIT('h1)
	) name1458 (
		_w1812_,
		_w1820_,
		_w1921_
	);
	LUT4 #(
		.INIT('heee8)
	) name1459 (
		_w1802_,
		_w1807_,
		_w1812_,
		_w1820_,
		_w1922_
	);
	LUT3 #(
		.INIT('h70)
	) name1460 (
		_w1914_,
		_w1920_,
		_w1922_,
		_w1923_
	);
	LUT2 #(
		.INIT('h1)
	) name1461 (
		_w1626_,
		_w1631_,
		_w1924_
	);
	LUT4 #(
		.INIT('heee0)
	) name1462 (
		_w1612_,
		_w1617_,
		_w1626_,
		_w1631_,
		_w1925_
	);
	LUT4 #(
		.INIT('h011f)
	) name1463 (
		_w1612_,
		_w1617_,
		_w1626_,
		_w1631_,
		_w1926_
	);
	LUT3 #(
		.INIT('h10)
	) name1464 (
		_w1909_,
		_w1910_,
		_w1926_,
		_w1927_
	);
	LUT3 #(
		.INIT('h0e)
	) name1465 (
		_w1306_,
		_w1586_,
		_w1592_,
		_w1928_
	);
	LUT4 #(
		.INIT('h00dc)
	) name1466 (
		_w1306_,
		_w1596_,
		_w1598_,
		_w1604_,
		_w1929_
	);
	LUT3 #(
		.INIT('h54)
	) name1467 (
		_w1909_,
		_w1928_,
		_w1929_,
		_w1930_
	);
	LUT2 #(
		.INIT('h1)
	) name1468 (
		_w1927_,
		_w1930_,
		_w1931_
	);
	LUT4 #(
		.INIT('h000d)
	) name1469 (
		_w1913_,
		_w1923_,
		_w1927_,
		_w1930_,
		_w1932_
	);
	LUT3 #(
		.INIT('h10)
	) name1470 (
		_w1306_,
		_w1441_,
		_w1449_,
		_w1933_
	);
	LUT4 #(
		.INIT('h5400)
	) name1471 (
		_w1306_,
		_w1452_,
		_w1478_,
		_w1483_,
		_w1934_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1472 (
		_w1306_,
		_w1441_,
		_w1449_,
		_w1934_,
		_w1935_
	);
	LUT3 #(
		.INIT('h10)
	) name1473 (
		_w1306_,
		_w1505_,
		_w1510_,
		_w1936_
	);
	LUT4 #(
		.INIT('h5400)
	) name1474 (
		_w1306_,
		_w1514_,
		_w1521_,
		_w1527_,
		_w1937_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1475 (
		_w1306_,
		_w1505_,
		_w1510_,
		_w1937_,
		_w1938_
	);
	LUT2 #(
		.INIT('h8)
	) name1476 (
		_w1935_,
		_w1938_,
		_w1939_
	);
	LUT3 #(
		.INIT('h10)
	) name1477 (
		_w1306_,
		_w1546_,
		_w1551_,
		_w1940_
	);
	LUT3 #(
		.INIT('h07)
	) name1478 (
		_w1534_,
		_w1542_,
		_w1940_,
		_w1941_
	);
	LUT4 #(
		.INIT('h5400)
	) name1479 (
		_w1306_,
		_w1555_,
		_w1559_,
		_w1564_,
		_w1942_
	);
	LUT3 #(
		.INIT('h10)
	) name1480 (
		_w1306_,
		_w1568_,
		_w1573_,
		_w1943_
	);
	LUT2 #(
		.INIT('h1)
	) name1481 (
		_w1942_,
		_w1943_,
		_w1944_
	);
	LUT2 #(
		.INIT('h8)
	) name1482 (
		_w1941_,
		_w1944_,
		_w1945_
	);
	LUT4 #(
		.INIT('h8000)
	) name1483 (
		_w1935_,
		_w1938_,
		_w1941_,
		_w1944_,
		_w1946_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1484 (
		_w1306_,
		_w1555_,
		_w1559_,
		_w1564_,
		_w1947_
	);
	LUT3 #(
		.INIT('h0e)
	) name1485 (
		_w1306_,
		_w1568_,
		_w1573_,
		_w1948_
	);
	LUT3 #(
		.INIT('h54)
	) name1486 (
		_w1942_,
		_w1947_,
		_w1948_,
		_w1949_
	);
	LUT3 #(
		.INIT('h0e)
	) name1487 (
		_w1306_,
		_w1546_,
		_w1551_,
		_w1950_
	);
	LUT3 #(
		.INIT('h8e)
	) name1488 (
		_w1534_,
		_w1542_,
		_w1950_,
		_w1951_
	);
	LUT3 #(
		.INIT('h70)
	) name1489 (
		_w1941_,
		_w1949_,
		_w1951_,
		_w1952_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1490 (
		_w1306_,
		_w1514_,
		_w1521_,
		_w1527_,
		_w1953_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1491 (
		_w1306_,
		_w1505_,
		_w1510_,
		_w1953_,
		_w1954_
	);
	LUT4 #(
		.INIT('hef0e)
	) name1492 (
		_w1306_,
		_w1505_,
		_w1510_,
		_w1953_,
		_w1955_
	);
	LUT3 #(
		.INIT('h0e)
	) name1493 (
		_w1306_,
		_w1441_,
		_w1449_,
		_w1956_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1494 (
		_w1306_,
		_w1452_,
		_w1478_,
		_w1483_,
		_w1957_
	);
	LUT4 #(
		.INIT('hef0e)
	) name1495 (
		_w1306_,
		_w1441_,
		_w1449_,
		_w1957_,
		_w1958_
	);
	LUT3 #(
		.INIT('h07)
	) name1496 (
		_w1935_,
		_w1955_,
		_w1958_,
		_w1959_
	);
	LUT3 #(
		.INIT('hd0)
	) name1497 (
		_w1939_,
		_w1952_,
		_w1959_,
		_w1960_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1498 (
		_w1918_,
		_w1932_,
		_w1946_,
		_w1960_,
		_w1961_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name1499 (
		\P2_reg2_reg[29]/NET0131 ,
		_w1298_,
		_w1404_,
		_w1961_,
		_w1962_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name1500 (
		_w1595_,
		_w1859_,
		_w1863_,
		_w1866_,
		_w1963_
	);
	LUT3 #(
		.INIT('h8a)
	) name1501 (
		_w1305_,
		_w1445_,
		_w1448_,
		_w1964_
	);
	LUT3 #(
		.INIT('h08)
	) name1502 (
		\P2_reg2_reg[31]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1965_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1503 (
		\P2_reg0_reg[31]/NET0131 ,
		\P2_reg1_reg[31]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1966_
	);
	LUT3 #(
		.INIT('h10)
	) name1504 (
		_w1397_,
		_w1965_,
		_w1966_,
		_w1967_
	);
	LUT3 #(
		.INIT('hef)
	) name1505 (
		_w1397_,
		_w1965_,
		_w1966_,
		_w1968_
	);
	LUT4 #(
		.INIT('h0001)
	) name1506 (
		_w1638_,
		_w1648_,
		_w1656_,
		_w1967_,
		_w1969_
	);
	LUT4 #(
		.INIT('h0777)
	) name1507 (
		_w1697_,
		_w1699_,
		_w1709_,
		_w1711_,
		_w1970_
	);
	LUT2 #(
		.INIT('h4)
	) name1508 (
		_w1722_,
		_w1970_,
		_w1971_
	);
	LUT4 #(
		.INIT('h1000)
	) name1509 (
		_w1670_,
		_w1675_,
		_w1969_,
		_w1971_,
		_w1972_
	);
	LUT4 #(
		.INIT('h0777)
	) name1510 (
		_w1688_,
		_w1690_,
		_w1777_,
		_w1778_,
		_w1973_
	);
	LUT4 #(
		.INIT('h0777)
	) name1511 (
		_w1738_,
		_w1739_,
		_w1750_,
		_w1751_,
		_w1974_
	);
	LUT2 #(
		.INIT('h4)
	) name1512 (
		_w1764_,
		_w1974_,
		_w1975_
	);
	LUT3 #(
		.INIT('h80)
	) name1513 (
		_w1972_,
		_w1973_,
		_w1975_,
		_w1976_
	);
	LUT4 #(
		.INIT('h0777)
	) name1514 (
		_w1822_,
		_w1824_,
		_w1832_,
		_w1833_,
		_w1977_
	);
	LUT4 #(
		.INIT('h8000)
	) name1515 (
		_w1972_,
		_w1973_,
		_w1975_,
		_w1977_,
		_w1978_
	);
	LUT3 #(
		.INIT('h01)
	) name1516 (
		_w1604_,
		_w1631_,
		_w1812_,
		_w1979_
	);
	LUT2 #(
		.INIT('h1)
	) name1517 (
		_w1617_,
		_w1807_,
		_w1980_
	);
	LUT3 #(
		.INIT('h01)
	) name1518 (
		_w1592_,
		_w1617_,
		_w1807_,
		_w1981_
	);
	LUT2 #(
		.INIT('h8)
	) name1519 (
		_w1979_,
		_w1981_,
		_w1982_
	);
	LUT3 #(
		.INIT('h40)
	) name1520 (
		_w1573_,
		_w1979_,
		_w1981_,
		_w1983_
	);
	LUT2 #(
		.INIT('h1)
	) name1521 (
		_w1551_,
		_w1564_,
		_w1984_
	);
	LUT4 #(
		.INIT('h4000)
	) name1522 (
		_w1573_,
		_w1979_,
		_w1981_,
		_w1984_,
		_w1985_
	);
	LUT2 #(
		.INIT('h4)
	) name1523 (
		_w1542_,
		_w1985_,
		_w1986_
	);
	LUT3 #(
		.INIT('h10)
	) name1524 (
		_w1527_,
		_w1542_,
		_w1985_,
		_w1987_
	);
	LUT4 #(
		.INIT('h000b)
	) name1525 (
		_w1445_,
		_w1448_,
		_w1483_,
		_w1510_,
		_w1988_
	);
	LUT2 #(
		.INIT('h4)
	) name1526 (
		_w1400_,
		_w1988_,
		_w1989_
	);
	LUT3 #(
		.INIT('h80)
	) name1527 (
		_w1978_,
		_w1987_,
		_w1989_,
		_w1990_
	);
	LUT3 #(
		.INIT('h20)
	) name1528 (
		\P2_reg1_reg[30]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1991_
	);
	LUT4 #(
		.INIT('hff35)
	) name1529 (
		\P2_reg0_reg[30]/NET0131 ,
		\P2_reg2_reg[30]/NET0131 ,
		_w1378_,
		_w1382_,
		_w1992_
	);
	LUT3 #(
		.INIT('h10)
	) name1530 (
		_w1397_,
		_w1991_,
		_w1992_,
		_w1993_
	);
	LUT3 #(
		.INIT('hef)
	) name1531 (
		_w1397_,
		_w1991_,
		_w1992_,
		_w1994_
	);
	LUT4 #(
		.INIT('h0080)
	) name1532 (
		_w1978_,
		_w1987_,
		_w1989_,
		_w1993_,
		_w1995_
	);
	LUT4 #(
		.INIT('h8828)
	) name1533 (
		\P2_B_reg/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1301_,
		_w1996_
	);
	LUT2 #(
		.INIT('h1)
	) name1534 (
		_w1305_,
		_w1996_,
		_w1997_
	);
	LUT4 #(
		.INIT('h1455)
	) name1535 (
		_w1964_,
		_w1990_,
		_w1993_,
		_w1997_,
		_w1998_
	);
	LUT4 #(
		.INIT('h8421)
	) name1536 (
		\P2_IR_reg[19]/NET0131 ,
		\P2_IR_reg[20]/NET0131 ,
		_w1264_,
		_w1272_,
		_w1999_
	);
	LUT3 #(
		.INIT('h80)
	) name1537 (
		_w1863_,
		_w1866_,
		_w1999_,
		_w2000_
	);
	LUT3 #(
		.INIT('h02)
	) name1538 (
		_w1859_,
		_w1863_,
		_w1866_,
		_w2001_
	);
	LUT3 #(
		.INIT('h10)
	) name1539 (
		_w1306_,
		_w1373_,
		_w2001_,
		_w2002_
	);
	LUT4 #(
		.INIT('h8000)
	) name1540 (
		_w1643_,
		_w1653_,
		_w1660_,
		_w1681_,
		_w2003_
	);
	LUT3 #(
		.INIT('h40)
	) name1541 (
		_w1726_,
		_w1666_,
		_w2003_,
		_w2004_
	);
	LUT4 #(
		.INIT('h1000)
	) name1542 (
		_w1717_,
		_w1726_,
		_w1666_,
		_w2003_,
		_w2005_
	);
	LUT3 #(
		.INIT('h10)
	) name1543 (
		_w1695_,
		_w1706_,
		_w2005_,
		_w2006_
	);
	LUT4 #(
		.INIT('heee0)
	) name1544 (
		_w1769_,
		_w1773_,
		_w1783_,
		_w1787_,
		_w2007_
	);
	LUT2 #(
		.INIT('h4)
	) name1545 (
		_w1747_,
		_w2007_,
		_w2008_
	);
	LUT4 #(
		.INIT('h1000)
	) name1546 (
		_w1695_,
		_w1706_,
		_w2005_,
		_w2008_,
		_w2009_
	);
	LUT2 #(
		.INIT('h1)
	) name1547 (
		_w1759_,
		_w1839_,
		_w2010_
	);
	LUT4 #(
		.INIT('h000e)
	) name1548 (
		_w1306_,
		_w1586_,
		_w1612_,
		_w1626_,
		_w2011_
	);
	LUT2 #(
		.INIT('h4)
	) name1549 (
		_w1599_,
		_w2011_,
		_w2012_
	);
	LUT3 #(
		.INIT('h10)
	) name1550 (
		_w1569_,
		_w1599_,
		_w2011_,
		_w2013_
	);
	LUT4 #(
		.INIT('haaae)
	) name1551 (
		_w1306_,
		_w1546_,
		_w1555_,
		_w1559_,
		_w2014_
	);
	LUT4 #(
		.INIT('h1000)
	) name1552 (
		_w1569_,
		_w1599_,
		_w2011_,
		_w2014_,
		_w2015_
	);
	LUT3 #(
		.INIT('h80)
	) name1553 (
		_w2009_,
		_w2010_,
		_w2015_,
		_w2016_
	);
	LUT3 #(
		.INIT('h01)
	) name1554 (
		_w1802_,
		_w1820_,
		_w1830_,
		_w2017_
	);
	LUT3 #(
		.INIT('h10)
	) name1555 (
		_w1522_,
		_w1534_,
		_w2017_,
		_w2018_
	);
	LUT3 #(
		.INIT('h32)
	) name1556 (
		_w1306_,
		_w1479_,
		_w1505_,
		_w2019_
	);
	LUT2 #(
		.INIT('h8)
	) name1557 (
		_w2018_,
		_w2019_,
		_w2020_
	);
	LUT2 #(
		.INIT('h8)
	) name1558 (
		_w2016_,
		_w2020_,
		_w2021_
	);
	LUT4 #(
		.INIT('h1000)
	) name1559 (
		_w1374_,
		_w1442_,
		_w2016_,
		_w2020_,
		_w2022_
	);
	LUT4 #(
		.INIT('h6555)
	) name1560 (
		_w1374_,
		_w1442_,
		_w2016_,
		_w2020_,
		_w2023_
	);
	LUT2 #(
		.INIT('h4)
	) name1561 (
		_w1863_,
		_w1999_,
		_w2024_
	);
	LUT3 #(
		.INIT('h10)
	) name1562 (
		_w1863_,
		_w1866_,
		_w1999_,
		_w2025_
	);
	LUT3 #(
		.INIT('h15)
	) name1563 (
		_w2002_,
		_w2023_,
		_w2025_,
		_w2026_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1564 (
		_w1298_,
		_w1998_,
		_w2000_,
		_w2026_,
		_w2027_
	);
	LUT4 #(
		.INIT('h4812)
	) name1565 (
		\P2_IR_reg[19]/NET0131 ,
		\P2_IR_reg[20]/NET0131 ,
		_w1264_,
		_w1272_,
		_w2028_
	);
	LUT3 #(
		.INIT('h10)
	) name1566 (
		_w1863_,
		_w1866_,
		_w2028_,
		_w2029_
	);
	LUT2 #(
		.INIT('h8)
	) name1567 (
		_w1396_,
		_w2029_,
		_w2030_
	);
	LUT2 #(
		.INIT('h4)
	) name1568 (
		_w1298_,
		_w2000_,
		_w2031_
	);
	LUT3 #(
		.INIT('h08)
	) name1569 (
		_w1863_,
		_w1866_,
		_w1999_,
		_w2032_
	);
	LUT3 #(
		.INIT('h01)
	) name1570 (
		_w1863_,
		_w1866_,
		_w2028_,
		_w2033_
	);
	LUT4 #(
		.INIT('h1ff2)
	) name1571 (
		_w1595_,
		_w1859_,
		_w1863_,
		_w1866_,
		_w2034_
	);
	LUT3 #(
		.INIT('h0d)
	) name1572 (
		_w1298_,
		_w2032_,
		_w2034_,
		_w2035_
	);
	LUT4 #(
		.INIT('h0a0b)
	) name1573 (
		_w1298_,
		_w2000_,
		_w2032_,
		_w2033_,
		_w2036_
	);
	LUT3 #(
		.INIT('h31)
	) name1574 (
		\P2_reg2_reg[29]/NET0131 ,
		_w2030_,
		_w2036_,
		_w2037_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1575 (
		_w1962_,
		_w1963_,
		_w2027_,
		_w2037_,
		_w2038_
	);
	LUT3 #(
		.INIT('h40)
	) name1576 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w2039_
	);
	LUT4 #(
		.INIT('h2000)
	) name1577 (
		\P2_reg2_reg[29]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w2040_
	);
	LUT4 #(
		.INIT('h0075)
	) name1578 (
		_w1285_,
		_w1870_,
		_w2038_,
		_w2040_,
		_w2041_
	);
	LUT4 #(
		.INIT('h8882)
	) name1579 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1264_,
		_w1266_,
		_w2042_
	);
	LUT2 #(
		.INIT('h2)
	) name1580 (
		\P2_reg2_reg[29]/NET0131 ,
		_w2042_,
		_w2043_
	);
	LUT3 #(
		.INIT('hf2)
	) name1581 (
		\P1_state_reg[0]/NET0131 ,
		_w2041_,
		_w2043_,
		_w2044_
	);
	LUT4 #(
		.INIT('h6669)
	) name1582 (
		\P1_B_reg/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		_w482_,
		_w1250_,
		_w2045_
	);
	LUT4 #(
		.INIT('h1428)
	) name1583 (
		\P1_IR_reg[25]/NET0131 ,
		\P1_IR_reg[26]/NET0131 ,
		_w573_,
		_w1247_,
		_w2046_
	);
	LUT2 #(
		.INIT('h4)
	) name1584 (
		_w2045_,
		_w2046_,
		_w2047_
	);
	LUT3 #(
		.INIT('h1d)
	) name1585 (
		\P1_d_reg[0]/NET0131 ,
		_w1249_,
		_w1251_,
		_w2048_
	);
	LUT2 #(
		.INIT('hb)
	) name1586 (
		_w2047_,
		_w2048_,
		_w2049_
	);
	LUT3 #(
		.INIT('h48)
	) name1587 (
		\P1_IR_reg[26]/NET0131 ,
		\P1_d_reg[1]/NET0131 ,
		_w573_,
		_w2050_
	);
	LUT4 #(
		.INIT('h8241)
	) name1588 (
		\P1_IR_reg[25]/NET0131 ,
		\P1_IR_reg[26]/NET0131 ,
		_w573_,
		_w1247_,
		_w2051_
	);
	LUT2 #(
		.INIT('h1)
	) name1589 (
		_w2050_,
		_w2051_,
		_w2052_
	);
	LUT4 #(
		.INIT('h1d1c)
	) name1590 (
		\P1_d_reg[1]/NET0131 ,
		_w1249_,
		_w1248_,
		_w2045_,
		_w2053_
	);
	LUT4 #(
		.INIT('he2e3)
	) name1591 (
		\P1_d_reg[1]/NET0131 ,
		_w1249_,
		_w1248_,
		_w2045_,
		_w2054_
	);
	LUT3 #(
		.INIT('h0b)
	) name1592 (
		_w2047_,
		_w2048_,
		_w2053_,
		_w2055_
	);
	LUT2 #(
		.INIT('h2)
	) name1593 (
		_w704_,
		_w2055_,
		_w2056_
	);
	LUT3 #(
		.INIT('h80)
	) name1594 (
		_w887_,
		_w888_,
		_w893_,
		_w2057_
	);
	LUT4 #(
		.INIT('h0008)
	) name1595 (
		_w873_,
		_w875_,
		_w881_,
		_w883_,
		_w2058_
	);
	LUT2 #(
		.INIT('h1)
	) name1596 (
		_w2057_,
		_w2058_,
		_w2059_
	);
	LUT3 #(
		.INIT('h07)
	) name1597 (
		_w909_,
		_w910_,
		_w915_,
		_w2060_
	);
	LUT3 #(
		.INIT('h23)
	) name1598 (
		_w1171_,
		_w1172_,
		_w2060_,
		_w2061_
	);
	LUT3 #(
		.INIT('h07)
	) name1599 (
		_w887_,
		_w888_,
		_w893_,
		_w2062_
	);
	LUT4 #(
		.INIT('h7770)
	) name1600 (
		_w873_,
		_w875_,
		_w881_,
		_w883_,
		_w2063_
	);
	LUT3 #(
		.INIT('h54)
	) name1601 (
		_w2058_,
		_w2062_,
		_w2063_,
		_w2064_
	);
	LUT3 #(
		.INIT('h0d)
	) name1602 (
		_w2059_,
		_w2061_,
		_w2064_,
		_w2065_
	);
	LUT3 #(
		.INIT('h80)
	) name1603 (
		_w924_,
		_w926_,
		_w933_,
		_w2066_
	);
	LUT2 #(
		.INIT('h1)
	) name1604 (
		_w1182_,
		_w2066_,
		_w2067_
	);
	LUT3 #(
		.INIT('h07)
	) name1605 (
		_w996_,
		_w997_,
		_w1001_,
		_w2068_
	);
	LUT3 #(
		.INIT('h8e)
	) name1606 (
		_w989_,
		_w993_,
		_w2068_,
		_w2069_
	);
	LUT3 #(
		.INIT('h80)
	) name1607 (
		_w978_,
		_w979_,
		_w984_,
		_w2070_
	);
	LUT2 #(
		.INIT('h1)
	) name1608 (
		_w1185_,
		_w2070_,
		_w2071_
	);
	LUT3 #(
		.INIT('h07)
	) name1609 (
		_w978_,
		_w979_,
		_w984_,
		_w2072_
	);
	LUT3 #(
		.INIT('h54)
	) name1610 (
		_w1185_,
		_w1186_,
		_w2072_,
		_w2073_
	);
	LUT3 #(
		.INIT('h0b)
	) name1611 (
		_w2069_,
		_w2071_,
		_w2073_,
		_w2074_
	);
	LUT3 #(
		.INIT('h80)
	) name1612 (
		_w946_,
		_w948_,
		_w956_,
		_w2075_
	);
	LUT2 #(
		.INIT('h1)
	) name1613 (
		_w1176_,
		_w2075_,
		_w2076_
	);
	LUT4 #(
		.INIT('hf400)
	) name1614 (
		_w2069_,
		_w2071_,
		_w2073_,
		_w2076_,
		_w2077_
	);
	LUT3 #(
		.INIT('h07)
	) name1615 (
		_w946_,
		_w948_,
		_w956_,
		_w2078_
	);
	LUT3 #(
		.INIT('h32)
	) name1616 (
		_w1175_,
		_w2075_,
		_w2078_,
		_w2079_
	);
	LUT3 #(
		.INIT('h07)
	) name1617 (
		_w924_,
		_w926_,
		_w933_,
		_w2080_
	);
	LUT3 #(
		.INIT('h23)
	) name1618 (
		_w1182_,
		_w1183_,
		_w2080_,
		_w2081_
	);
	LUT4 #(
		.INIT('h5700)
	) name1619 (
		_w2067_,
		_w2077_,
		_w2079_,
		_w2081_,
		_w2082_
	);
	LUT3 #(
		.INIT('h80)
	) name1620 (
		_w909_,
		_w910_,
		_w915_,
		_w2083_
	);
	LUT2 #(
		.INIT('h1)
	) name1621 (
		_w1171_,
		_w2083_,
		_w2084_
	);
	LUT4 #(
		.INIT('h0001)
	) name1622 (
		_w1171_,
		_w2057_,
		_w2058_,
		_w2083_,
		_w2085_
	);
	LUT4 #(
		.INIT('h0777)
	) name1623 (
		_w749_,
		_w754_,
		_w759_,
		_w764_,
		_w2086_
	);
	LUT4 #(
		.INIT('h0e00)
	) name1624 (
		_w489_,
		_w717_,
		_w719_,
		_w724_,
		_w2087_
	);
	LUT3 #(
		.INIT('h04)
	) name1625 (
		_w1215_,
		_w2086_,
		_w2087_,
		_w2088_
	);
	LUT4 #(
		.INIT('h0777)
	) name1626 (
		_w827_,
		_w833_,
		_w837_,
		_w842_,
		_w2089_
	);
	LUT4 #(
		.INIT('h0777)
	) name1627 (
		_w847_,
		_w852_,
		_w856_,
		_w864_,
		_w2090_
	);
	LUT2 #(
		.INIT('h8)
	) name1628 (
		_w2089_,
		_w2090_,
		_w2091_
	);
	LUT2 #(
		.INIT('h8)
	) name1629 (
		_w2088_,
		_w2091_,
		_w2092_
	);
	LUT4 #(
		.INIT('h7500)
	) name1630 (
		_w2065_,
		_w2082_,
		_w2085_,
		_w2092_,
		_w2093_
	);
	LUT4 #(
		.INIT('h1117)
	) name1631 (
		_w847_,
		_w852_,
		_w856_,
		_w864_,
		_w2094_
	);
	LUT4 #(
		.INIT('heee8)
	) name1632 (
		_w827_,
		_w833_,
		_w837_,
		_w842_,
		_w2095_
	);
	LUT3 #(
		.INIT('h70)
	) name1633 (
		_w2089_,
		_w2094_,
		_w2095_,
		_w2096_
	);
	LUT4 #(
		.INIT('heee8)
	) name1634 (
		_w749_,
		_w754_,
		_w759_,
		_w764_,
		_w2097_
	);
	LUT3 #(
		.INIT('h01)
	) name1635 (
		_w1215_,
		_w2087_,
		_w2097_,
		_w2098_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1636 (
		_w489_,
		_w717_,
		_w719_,
		_w724_,
		_w2099_
	);
	LUT3 #(
		.INIT('h0d)
	) name1637 (
		_w1214_,
		_w2087_,
		_w2099_,
		_w2100_
	);
	LUT2 #(
		.INIT('h4)
	) name1638 (
		_w2098_,
		_w2100_,
		_w2101_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1639 (
		_w2088_,
		_w2096_,
		_w2098_,
		_w2100_,
		_w2102_
	);
	LUT4 #(
		.INIT('h001f)
	) name1640 (
		_w489_,
		_w1040_,
		_w1047_,
		_w1222_,
		_w2103_
	);
	LUT2 #(
		.INIT('h1)
	) name1641 (
		_w1219_,
		_w1208_,
		_w2104_
	);
	LUT2 #(
		.INIT('h8)
	) name1642 (
		_w2103_,
		_w2104_,
		_w2105_
	);
	LUT2 #(
		.INIT('h1)
	) name1643 (
		_w1199_,
		_w1211_,
		_w2106_
	);
	LUT2 #(
		.INIT('h1)
	) name1644 (
		_w1227_,
		_w1202_,
		_w2107_
	);
	LUT4 #(
		.INIT('h0001)
	) name1645 (
		_w1227_,
		_w1199_,
		_w1202_,
		_w1211_,
		_w2108_
	);
	LUT3 #(
		.INIT('h80)
	) name1646 (
		_w2103_,
		_w2104_,
		_w2108_,
		_w2109_
	);
	LUT3 #(
		.INIT('h0d)
	) name1647 (
		_w1226_,
		_w1202_,
		_w1203_,
		_w2110_
	);
	LUT3 #(
		.INIT('h0d)
	) name1648 (
		_w1200_,
		_w1211_,
		_w1212_,
		_w2111_
	);
	LUT3 #(
		.INIT('hd0)
	) name1649 (
		_w2106_,
		_w2110_,
		_w2111_,
		_w2112_
	);
	LUT3 #(
		.INIT('h23)
	) name1650 (
		_w1219_,
		_w1220_,
		_w1209_,
		_w2113_
	);
	LUT4 #(
		.INIT('h040d)
	) name1651 (
		_w1059_,
		_w1063_,
		_w1223_,
		_w1209_,
		_w2114_
	);
	LUT3 #(
		.INIT('h51)
	) name1652 (
		_w1163_,
		_w2103_,
		_w2114_,
		_w2115_
	);
	LUT3 #(
		.INIT('hd0)
	) name1653 (
		_w2105_,
		_w2112_,
		_w2115_,
		_w2116_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1654 (
		_w2093_,
		_w2102_,
		_w2109_,
		_w2116_,
		_w2117_
	);
	LUT4 #(
		.INIT('h070b)
	) name1655 (
		_w1160_,
		_w2055_,
		_w2056_,
		_w2117_,
		_w2118_
	);
	LUT3 #(
		.INIT('h07)
	) name1656 (
		_w1096_,
		_w1100_,
		_w1111_,
		_w2119_
	);
	LUT2 #(
		.INIT('h6)
	) name1657 (
		_w1096_,
		_w1098_,
		_w2120_
	);
	LUT4 #(
		.INIT('h5202)
	) name1658 (
		_w1096_,
		_w1100_,
		_w1098_,
		_w718_,
		_w2121_
	);
	LUT2 #(
		.INIT('h8)
	) name1659 (
		_w872_,
		_w1023_,
		_w2122_
	);
	LUT4 #(
		.INIT('h1011)
	) name1660 (
		_w768_,
		_w771_,
		_w870_,
		_w1023_,
		_w2123_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1661 (
		_w922_,
		_w1019_,
		_w2122_,
		_w2123_,
		_w2124_
	);
	LUT3 #(
		.INIT('h80)
	) name1662 (
		_w1021_,
		_w1050_,
		_w1082_,
		_w2125_
	);
	LUT3 #(
		.INIT('hb0)
	) name1663 (
		_w817_,
		_w1083_,
		_w1090_,
		_w2126_
	);
	LUT4 #(
		.INIT('h9a55)
	) name1664 (
		_w1160_,
		_w2124_,
		_w2125_,
		_w2126_,
		_w2127_
	);
	LUT4 #(
		.INIT('h0858)
	) name1665 (
		_w1096_,
		_w1100_,
		_w1098_,
		_w718_,
		_w2128_
	);
	LUT4 #(
		.INIT('h2e00)
	) name1666 (
		_w704_,
		_w2055_,
		_w2127_,
		_w2128_,
		_w2129_
	);
	LUT4 #(
		.INIT('h0001)
	) name1667 (
		_w980_,
		_w989_,
		_w998_,
		_w602_,
		_w2130_
	);
	LUT4 #(
		.INIT('h0777)
	) name1668 (
		_w896_,
		_w898_,
		_w909_,
		_w910_,
		_w2131_
	);
	LUT4 #(
		.INIT('h0777)
	) name1669 (
		_w924_,
		_w926_,
		_w935_,
		_w937_,
		_w2132_
	);
	LUT3 #(
		.INIT('h40)
	) name1670 (
		_w949_,
		_w2131_,
		_w2132_,
		_w2133_
	);
	LUT4 #(
		.INIT('h1000)
	) name1671 (
		_w961_,
		_w971_,
		_w2130_,
		_w2133_,
		_w2134_
	);
	LUT4 #(
		.INIT('h0777)
	) name1672 (
		_w834_,
		_w836_,
		_w845_,
		_w846_,
		_w2135_
	);
	LUT4 #(
		.INIT('h0777)
	) name1673 (
		_w824_,
		_w826_,
		_w854_,
		_w855_,
		_w2136_
	);
	LUT3 #(
		.INIT('h40)
	) name1674 (
		_w876_,
		_w2135_,
		_w2136_,
		_w2137_
	);
	LUT3 #(
		.INIT('h40)
	) name1675 (
		_w889_,
		_w2134_,
		_w2137_,
		_w2138_
	);
	LUT4 #(
		.INIT('h1000)
	) name1676 (
		_w764_,
		_w889_,
		_w2134_,
		_w2137_,
		_w2139_
	);
	LUT2 #(
		.INIT('h1)
	) name1677 (
		_w724_,
		_w810_,
		_w2140_
	);
	LUT4 #(
		.INIT('h0001)
	) name1678 (
		_w724_,
		_w780_,
		_w800_,
		_w810_,
		_w2141_
	);
	LUT2 #(
		.INIT('h4)
	) name1679 (
		_w789_,
		_w2141_,
		_w2142_
	);
	LUT3 #(
		.INIT('h45)
	) name1680 (
		_w1063_,
		_w1075_,
		_w1078_,
		_w2143_
	);
	LUT3 #(
		.INIT('h40)
	) name1681 (
		_w789_,
		_w2141_,
		_w2143_,
		_w2144_
	);
	LUT3 #(
		.INIT('h45)
	) name1682 (
		_w1035_,
		_w1043_,
		_w1046_,
		_w2145_
	);
	LUT4 #(
		.INIT('h4000)
	) name1683 (
		_w789_,
		_w2141_,
		_w2143_,
		_w2145_,
		_w2146_
	);
	LUT2 #(
		.INIT('h1)
	) name1684 (
		_w739_,
		_w754_,
		_w2147_
	);
	LUT2 #(
		.INIT('h4)
	) name1685 (
		_w708_,
		_w2147_,
		_w2148_
	);
	LUT2 #(
		.INIT('h8)
	) name1686 (
		_w2146_,
		_w2148_,
		_w2149_
	);
	LUT4 #(
		.INIT('h4111)
	) name1687 (
		_w488_,
		_w677_,
		_w2139_,
		_w2149_,
		_w2150_
	);
	LUT3 #(
		.INIT('h8a)
	) name1688 (
		_w488_,
		_w1043_,
		_w1046_,
		_w2151_
	);
	LUT4 #(
		.INIT('h1113)
	) name1689 (
		_w2055_,
		_w2056_,
		_w2150_,
		_w2151_,
		_w2152_
	);
	LUT3 #(
		.INIT('h80)
	) name1690 (
		_w734_,
		_w749_,
		_w759_,
		_w2153_
	);
	LUT2 #(
		.INIT('h1)
	) name1691 (
		_w776_,
		_w796_,
		_w2154_
	);
	LUT4 #(
		.INIT('h2000)
	) name1692 (
		_w720_,
		_w805_,
		_w2153_,
		_w2154_,
		_w2155_
	);
	LUT4 #(
		.INIT('h8000)
	) name1693 (
		_w976_,
		_w984_,
		_w993_,
		_w1001_,
		_w2156_
	);
	LUT3 #(
		.INIT('h80)
	) name1694 (
		_w956_,
		_w966_,
		_w2156_,
		_w2157_
	);
	LUT2 #(
		.INIT('h8)
	) name1695 (
		_w933_,
		_w943_,
		_w2158_
	);
	LUT4 #(
		.INIT('h8000)
	) name1696 (
		_w956_,
		_w966_,
		_w2156_,
		_w2158_,
		_w2159_
	);
	LUT2 #(
		.INIT('h8)
	) name1697 (
		_w905_,
		_w915_,
		_w2160_
	);
	LUT3 #(
		.INIT('h10)
	) name1698 (
		_w881_,
		_w883_,
		_w893_,
		_w2161_
	);
	LUT4 #(
		.INIT('h8000)
	) name1699 (
		_w833_,
		_w842_,
		_w852_,
		_w864_,
		_w2162_
	);
	LUT4 #(
		.INIT('h8000)
	) name1700 (
		_w2159_,
		_w2160_,
		_w2161_,
		_w2162_,
		_w2163_
	);
	LUT3 #(
		.INIT('h0e)
	) name1701 (
		_w489_,
		_w783_,
		_w1073_,
		_w2164_
	);
	LUT3 #(
		.INIT('hea)
	) name1702 (
		_w489_,
		_w1030_,
		_w1058_,
		_w2165_
	);
	LUT2 #(
		.INIT('h8)
	) name1703 (
		_w2164_,
		_w2165_,
		_w2166_
	);
	LUT4 #(
		.INIT('he000)
	) name1704 (
		_w489_,
		_w1040_,
		_w2164_,
		_w2165_,
		_w2167_
	);
	LUT4 #(
		.INIT('h4000)
	) name1705 (
		_w702_,
		_w2155_,
		_w2163_,
		_w2167_,
		_w2168_
	);
	LUT4 #(
		.INIT('h9555)
	) name1706 (
		_w702_,
		_w2155_,
		_w2163_,
		_w2167_,
		_w2169_
	);
	LUT3 #(
		.INIT('h10)
	) name1707 (
		_w1096_,
		_w1098_,
		_w1122_,
		_w2170_
	);
	LUT3 #(
		.INIT('h08)
	) name1708 (
		_w1096_,
		_w1098_,
		_w1122_,
		_w2171_
	);
	LUT3 #(
		.INIT('h01)
	) name1709 (
		_w1096_,
		_w1098_,
		_w1101_,
		_w2172_
	);
	LUT4 #(
		.INIT('h5400)
	) name1710 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2172_,
		_w2173_
	);
	LUT3 #(
		.INIT('ha8)
	) name1711 (
		_w704_,
		_w2171_,
		_w2173_,
		_w2174_
	);
	LUT4 #(
		.INIT('h1110)
	) name1712 (
		_w1120_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w2175_
	);
	LUT3 #(
		.INIT('h01)
	) name1713 (
		_w1096_,
		_w1098_,
		_w1122_,
		_w2176_
	);
	LUT2 #(
		.INIT('h4)
	) name1714 (
		_w2175_,
		_w2176_,
		_w2177_
	);
	LUT3 #(
		.INIT('h13)
	) name1715 (
		_w702_,
		_w2174_,
		_w2177_,
		_w2178_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1716 (
		_w2055_,
		_w2169_,
		_w2170_,
		_w2178_,
		_w2179_
	);
	LUT3 #(
		.INIT('hd0)
	) name1717 (
		_w1237_,
		_w2152_,
		_w2179_,
		_w2180_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1718 (
		_w2118_,
		_w2121_,
		_w2129_,
		_w2180_,
		_w2181_
	);
	LUT4 #(
		.INIT('h4555)
	) name1719 (
		_w1243_,
		_w1249_,
		_w1251_,
		_w1248_,
		_w2182_
	);
	LUT4 #(
		.INIT('h1000)
	) name1720 (
		_w1243_,
		_w1249_,
		_w1251_,
		_w1248_,
		_w2183_
	);
	LUT2 #(
		.INIT('h8)
	) name1721 (
		_w704_,
		_w2183_,
		_w2184_
	);
	LUT4 #(
		.INIT('haa20)
	) name1722 (
		\P1_state_reg[0]/NET0131 ,
		_w2181_,
		_w2182_,
		_w2184_,
		_w2185_
	);
	LUT2 #(
		.INIT('h2)
	) name1723 (
		\P1_reg3_reg[28]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2186_
	);
	LUT3 #(
		.INIT('h07)
	) name1724 (
		_w704_,
		_w1244_,
		_w2186_,
		_w2187_
	);
	LUT2 #(
		.INIT('hb)
	) name1725 (
		_w2185_,
		_w2187_,
		_w2188_
	);
	LUT3 #(
		.INIT('h04)
	) name1726 (
		_w2047_,
		_w2048_,
		_w2053_,
		_w2189_
	);
	LUT4 #(
		.INIT('h3c55)
	) name1727 (
		\P1_reg2_reg[28]/NET0131 ,
		_w1160_,
		_w2117_,
		_w2189_,
		_w2190_
	);
	LUT4 #(
		.INIT('h30a0)
	) name1728 (
		\P1_reg2_reg[28]/NET0131 ,
		_w2127_,
		_w2128_,
		_w2189_,
		_w2191_
	);
	LUT4 #(
		.INIT('h0355)
	) name1729 (
		\P1_reg2_reg[28]/NET0131 ,
		_w2150_,
		_w2151_,
		_w2189_,
		_w2192_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name1730 (
		\P1_reg2_reg[28]/NET0131 ,
		_w2169_,
		_w2170_,
		_w2189_,
		_w2193_
	);
	LUT3 #(
		.INIT('h04)
	) name1731 (
		_w1096_,
		_w1100_,
		_w1098_,
		_w2194_
	);
	LUT4 #(
		.INIT('h5400)
	) name1732 (
		_w489_,
		_w680_,
		_w701_,
		_w2194_,
		_w2195_
	);
	LUT4 #(
		.INIT('hfb00)
	) name1733 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2194_,
		_w2196_
	);
	LUT3 #(
		.INIT('ha8)
	) name1734 (
		\P1_reg2_reg[28]/NET0131 ,
		_w2171_,
		_w2196_,
		_w2197_
	);
	LUT2 #(
		.INIT('h8)
	) name1735 (
		_w704_,
		_w1120_,
		_w2198_
	);
	LUT4 #(
		.INIT('h0103)
	) name1736 (
		_w2189_,
		_w2197_,
		_w2198_,
		_w2195_,
		_w2199_
	);
	LUT2 #(
		.INIT('h4)
	) name1737 (
		_w2193_,
		_w2199_,
		_w2200_
	);
	LUT3 #(
		.INIT('hd0)
	) name1738 (
		_w1237_,
		_w2192_,
		_w2200_,
		_w2201_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1739 (
		_w2121_,
		_w2190_,
		_w2191_,
		_w2201_,
		_w2202_
	);
	LUT2 #(
		.INIT('h8)
	) name1740 (
		\P1_reg2_reg[28]/NET0131 ,
		_w2183_,
		_w2203_
	);
	LUT4 #(
		.INIT('haa08)
	) name1741 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w2202_,
		_w2203_,
		_w2204_
	);
	LUT3 #(
		.INIT('h84)
	) name1742 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w2205_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1743 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[28]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w2206_
	);
	LUT2 #(
		.INIT('he)
	) name1744 (
		_w2204_,
		_w2206_,
		_w2207_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1745 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[29]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w2208_
	);
	LUT2 #(
		.INIT('h8)
	) name1746 (
		\P1_reg2_reg[29]/NET0131 ,
		_w2183_,
		_w2209_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1747 (
		\P1_reg2_reg[29]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w2210_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1748 (
		_w488_,
		_w585_,
		_w704_,
		_w707_,
		_w2211_
	);
	LUT3 #(
		.INIT('h01)
	) name1749 (
		_w739_,
		_w754_,
		_w764_,
		_w2212_
	);
	LUT4 #(
		.INIT('h4000)
	) name1750 (
		_w889_,
		_w2134_,
		_w2137_,
		_w2212_,
		_w2213_
	);
	LUT4 #(
		.INIT('h1000)
	) name1751 (
		_w677_,
		_w708_,
		_w2146_,
		_w2213_,
		_w2214_
	);
	LUT4 #(
		.INIT('h8828)
	) name1752 (
		\P1_B_reg/NET0131 ,
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w478_,
		_w2215_
	);
	LUT2 #(
		.INIT('h1)
	) name1753 (
		_w488_,
		_w2215_,
		_w2216_
	);
	LUT4 #(
		.INIT('h1233)
	) name1754 (
		_w650_,
		_w2211_,
		_w2214_,
		_w2216_,
		_w2217_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1755 (
		\P1_reg2_reg[29]/NET0131 ,
		_w1237_,
		_w2189_,
		_w2217_,
		_w2218_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1756 (
		_w734_,
		_w739_,
		_w749_,
		_w754_,
		_w2219_
	);
	LUT3 #(
		.INIT('h10)
	) name1757 (
		_w726_,
		_w818_,
		_w2219_,
		_w2220_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1758 (
		_w837_,
		_w842_,
		_w847_,
		_w852_,
		_w2221_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name1759 (
		_w759_,
		_w764_,
		_w827_,
		_w833_,
		_w2222_
	);
	LUT2 #(
		.INIT('h8)
	) name1760 (
		_w2221_,
		_w2222_,
		_w2223_
	);
	LUT2 #(
		.INIT('h8)
	) name1761 (
		_w2220_,
		_w2223_,
		_w2224_
	);
	LUT3 #(
		.INIT('h0d)
	) name1762 (
		_w856_,
		_w864_,
		_w885_,
		_w2225_
	);
	LUT3 #(
		.INIT('h54)
	) name1763 (
		_w894_,
		_w907_,
		_w918_,
		_w2226_
	);
	LUT3 #(
		.INIT('h2b)
	) name1764 (
		_w856_,
		_w864_,
		_w919_,
		_w2227_
	);
	LUT3 #(
		.INIT('h70)
	) name1765 (
		_w2225_,
		_w2226_,
		_w2227_,
		_w2228_
	);
	LUT4 #(
		.INIT('h00b2)
	) name1766 (
		_w989_,
		_w993_,
		_w1002_,
		_w1005_,
		_w2229_
	);
	LUT3 #(
		.INIT('h01)
	) name1767 (
		_w967_,
		_w977_,
		_w985_,
		_w2230_
	);
	LUT3 #(
		.INIT('h54)
	) name1768 (
		_w967_,
		_w1004_,
		_w1009_,
		_w2231_
	);
	LUT3 #(
		.INIT('h0b)
	) name1769 (
		_w2229_,
		_w2230_,
		_w2231_,
		_w2232_
	);
	LUT2 #(
		.INIT('h1)
	) name1770 (
		_w944_,
		_w1016_,
		_w2233_
	);
	LUT2 #(
		.INIT('h1)
	) name1771 (
		_w934_,
		_w957_,
		_w2234_
	);
	LUT4 #(
		.INIT('h0001)
	) name1772 (
		_w934_,
		_w944_,
		_w957_,
		_w1016_,
		_w2235_
	);
	LUT4 #(
		.INIT('hf400)
	) name1773 (
		_w2229_,
		_w2230_,
		_w2231_,
		_w2235_,
		_w2236_
	);
	LUT3 #(
		.INIT('h54)
	) name1774 (
		_w934_,
		_w1008_,
		_w1012_,
		_w2237_
	);
	LUT3 #(
		.INIT('h0e)
	) name1775 (
		_w916_,
		_w1011_,
		_w1016_,
		_w2238_
	);
	LUT3 #(
		.INIT('h07)
	) name1776 (
		_w2233_,
		_w2237_,
		_w2238_,
		_w2239_
	);
	LUT2 #(
		.INIT('h1)
	) name1777 (
		_w894_,
		_w906_,
		_w2240_
	);
	LUT2 #(
		.INIT('h8)
	) name1778 (
		_w2225_,
		_w2240_,
		_w2241_
	);
	LUT3 #(
		.INIT('hb0)
	) name1779 (
		_w2236_,
		_w2239_,
		_w2241_,
		_w2242_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1780 (
		_w2228_,
		_w2236_,
		_w2239_,
		_w2241_,
		_w2243_
	);
	LUT4 #(
		.INIT('h4d44)
	) name1781 (
		_w837_,
		_w842_,
		_w847_,
		_w852_,
		_w2244_
	);
	LUT4 #(
		.INIT('h2b22)
	) name1782 (
		_w759_,
		_w764_,
		_w827_,
		_w833_,
		_w2245_
	);
	LUT3 #(
		.INIT('h07)
	) name1783 (
		_w2222_,
		_w2244_,
		_w2245_,
		_w2246_
	);
	LUT4 #(
		.INIT('h22b2)
	) name1784 (
		_w734_,
		_w739_,
		_w749_,
		_w754_,
		_w2247_
	);
	LUT3 #(
		.INIT('h10)
	) name1785 (
		_w726_,
		_w818_,
		_w2247_,
		_w2248_
	);
	LUT3 #(
		.INIT('h0e)
	) name1786 (
		_w770_,
		_w812_,
		_w818_,
		_w2249_
	);
	LUT2 #(
		.INIT('h1)
	) name1787 (
		_w2248_,
		_w2249_,
		_w2250_
	);
	LUT4 #(
		.INIT('h000d)
	) name1788 (
		_w2220_,
		_w2246_,
		_w2248_,
		_w2249_,
		_w2251_
	);
	LUT4 #(
		.INIT('h0777)
	) name1789 (
		_w776_,
		_w780_,
		_w796_,
		_w800_,
		_w2252_
	);
	LUT3 #(
		.INIT('h10)
	) name1790 (
		_w791_,
		_w1081_,
		_w2252_,
		_w2253_
	);
	LUT2 #(
		.INIT('h1)
	) name1791 (
		_w1037_,
		_w1065_,
		_w2254_
	);
	LUT3 #(
		.INIT('h10)
	) name1792 (
		_w1049_,
		_w1092_,
		_w2254_,
		_w2255_
	);
	LUT4 #(
		.INIT('h1000)
	) name1793 (
		_w1049_,
		_w1092_,
		_w2253_,
		_w2254_,
		_w2256_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1794 (
		_w2224_,
		_w2243_,
		_w2251_,
		_w2256_,
		_w2257_
	);
	LUT4 #(
		.INIT('h1117)
	) name1795 (
		_w776_,
		_w780_,
		_w796_,
		_w800_,
		_w2258_
	);
	LUT3 #(
		.INIT('h10)
	) name1796 (
		_w791_,
		_w1081_,
		_w2258_,
		_w2259_
	);
	LUT3 #(
		.INIT('h32)
	) name1797 (
		_w814_,
		_w1081_,
		_w1087_,
		_w2260_
	);
	LUT2 #(
		.INIT('h1)
	) name1798 (
		_w2259_,
		_w2260_,
		_w2261_
	);
	LUT3 #(
		.INIT('h54)
	) name1799 (
		_w1037_,
		_w1085_,
		_w1086_,
		_w2262_
	);
	LUT4 #(
		.INIT('h0701)
	) name1800 (
		_w1041_,
		_w1047_,
		_w1092_,
		_w2262_,
		_w2263_
	);
	LUT4 #(
		.INIT('h0051)
	) name1801 (
		_w710_,
		_w2255_,
		_w2261_,
		_w2263_,
		_w2264_
	);
	LUT4 #(
		.INIT('h4844)
	) name1802 (
		_w1197_,
		_w2189_,
		_w2257_,
		_w2264_,
		_w2265_
	);
	LUT3 #(
		.INIT('ha8)
	) name1803 (
		_w2128_,
		_w2210_,
		_w2265_,
		_w2266_
	);
	LUT2 #(
		.INIT('h1)
	) name1804 (
		_w1171_,
		_w2057_,
		_w2267_
	);
	LUT3 #(
		.INIT('h07)
	) name1805 (
		_w856_,
		_w864_,
		_w2058_,
		_w2268_
	);
	LUT2 #(
		.INIT('h8)
	) name1806 (
		_w2267_,
		_w2268_,
		_w2269_
	);
	LUT4 #(
		.INIT('h008e)
	) name1807 (
		_w989_,
		_w993_,
		_w2068_,
		_w2072_,
		_w2270_
	);
	LUT2 #(
		.INIT('h1)
	) name1808 (
		_w1186_,
		_w1175_,
		_w2271_
	);
	LUT4 #(
		.INIT('h0455)
	) name1809 (
		_w1176_,
		_w2071_,
		_w2270_,
		_w2271_,
		_w2272_
	);
	LUT2 #(
		.INIT('h1)
	) name1810 (
		_w1182_,
		_w2083_,
		_w2273_
	);
	LUT2 #(
		.INIT('h1)
	) name1811 (
		_w2066_,
		_w2075_,
		_w2274_
	);
	LUT4 #(
		.INIT('h0001)
	) name1812 (
		_w1182_,
		_w2066_,
		_w2075_,
		_w2083_,
		_w2275_
	);
	LUT3 #(
		.INIT('h80)
	) name1813 (
		_w2269_,
		_w2272_,
		_w2275_,
		_w2276_
	);
	LUT3 #(
		.INIT('h54)
	) name1814 (
		_w2066_,
		_w2078_,
		_w2080_,
		_w2277_
	);
	LUT3 #(
		.INIT('h31)
	) name1815 (
		_w1183_,
		_w2060_,
		_w2083_,
		_w2278_
	);
	LUT3 #(
		.INIT('h70)
	) name1816 (
		_w2273_,
		_w2277_,
		_w2278_,
		_w2279_
	);
	LUT3 #(
		.INIT('h32)
	) name1817 (
		_w1172_,
		_w2057_,
		_w2062_,
		_w2280_
	);
	LUT3 #(
		.INIT('h8e)
	) name1818 (
		_w856_,
		_w864_,
		_w2063_,
		_w2281_
	);
	LUT3 #(
		.INIT('h70)
	) name1819 (
		_w2268_,
		_w2280_,
		_w2281_,
		_w2282_
	);
	LUT3 #(
		.INIT('hd0)
	) name1820 (
		_w2269_,
		_w2279_,
		_w2282_,
		_w2283_
	);
	LUT4 #(
		.INIT('h0777)
	) name1821 (
		_w734_,
		_w739_,
		_w749_,
		_w754_,
		_w2284_
	);
	LUT3 #(
		.INIT('h10)
	) name1822 (
		_w1227_,
		_w2087_,
		_w2284_,
		_w2285_
	);
	LUT4 #(
		.INIT('h0777)
	) name1823 (
		_w837_,
		_w842_,
		_w847_,
		_w852_,
		_w2286_
	);
	LUT4 #(
		.INIT('h0777)
	) name1824 (
		_w759_,
		_w764_,
		_w827_,
		_w833_,
		_w2287_
	);
	LUT2 #(
		.INIT('h8)
	) name1825 (
		_w2286_,
		_w2287_,
		_w2288_
	);
	LUT2 #(
		.INIT('h8)
	) name1826 (
		_w2285_,
		_w2288_,
		_w2289_
	);
	LUT4 #(
		.INIT('heee8)
	) name1827 (
		_w837_,
		_w842_,
		_w847_,
		_w852_,
		_w2290_
	);
	LUT4 #(
		.INIT('h1117)
	) name1828 (
		_w759_,
		_w764_,
		_w827_,
		_w833_,
		_w2291_
	);
	LUT3 #(
		.INIT('h0d)
	) name1829 (
		_w2287_,
		_w2290_,
		_w2291_,
		_w2292_
	);
	LUT4 #(
		.INIT('heee8)
	) name1830 (
		_w734_,
		_w739_,
		_w749_,
		_w754_,
		_w2293_
	);
	LUT3 #(
		.INIT('h01)
	) name1831 (
		_w1227_,
		_w2087_,
		_w2293_,
		_w2294_
	);
	LUT3 #(
		.INIT('h45)
	) name1832 (
		_w1226_,
		_w1227_,
		_w2099_,
		_w2295_
	);
	LUT2 #(
		.INIT('h4)
	) name1833 (
		_w2294_,
		_w2295_,
		_w2296_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1834 (
		_w2285_,
		_w2292_,
		_w2294_,
		_w2295_,
		_w2297_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1835 (
		_w2276_,
		_w2283_,
		_w2289_,
		_w2297_,
		_w2298_
	);
	LUT2 #(
		.INIT('h1)
	) name1836 (
		_w1164_,
		_w1158_,
		_w2299_
	);
	LUT2 #(
		.INIT('h1)
	) name1837 (
		_w1219_,
		_w1222_,
		_w2300_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1838 (
		_w776_,
		_w780_,
		_w796_,
		_w800_,
		_w2301_
	);
	LUT3 #(
		.INIT('h10)
	) name1839 (
		_w1208_,
		_w1211_,
		_w2301_,
		_w2302_
	);
	LUT4 #(
		.INIT('h1000)
	) name1840 (
		_w1164_,
		_w1158_,
		_w2300_,
		_w2302_,
		_w2303_
	);
	LUT4 #(
		.INIT('hdd4d)
	) name1841 (
		_w776_,
		_w780_,
		_w796_,
		_w800_,
		_w2304_
	);
	LUT3 #(
		.INIT('h01)
	) name1842 (
		_w1208_,
		_w1211_,
		_w2304_,
		_w2305_
	);
	LUT3 #(
		.INIT('h23)
	) name1843 (
		_w1208_,
		_w1209_,
		_w1212_,
		_w2306_
	);
	LUT2 #(
		.INIT('h4)
	) name1844 (
		_w2305_,
		_w2306_,
		_w2307_
	);
	LUT3 #(
		.INIT('h0d)
	) name1845 (
		_w1220_,
		_w1222_,
		_w1223_,
		_w2308_
	);
	LUT4 #(
		.INIT('h7500)
	) name1846 (
		_w2300_,
		_w2305_,
		_w2306_,
		_w2308_,
		_w2309_
	);
	LUT3 #(
		.INIT('h0d)
	) name1847 (
		_w1163_,
		_w1158_,
		_w1159_,
		_w2310_
	);
	LUT3 #(
		.INIT('hd0)
	) name1848 (
		_w2299_,
		_w2309_,
		_w2310_,
		_w2311_
	);
	LUT4 #(
		.INIT('h9a55)
	) name1849 (
		_w1197_,
		_w2298_,
		_w2303_,
		_w2311_,
		_w2312_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1850 (
		\P1_reg2_reg[29]/NET0131 ,
		_w2121_,
		_w2189_,
		_w2312_,
		_w2313_
	);
	LUT4 #(
		.INIT('h3c55)
	) name1851 (
		\P1_reg2_reg[29]/NET0131 ,
		_w674_,
		_w2168_,
		_w2189_,
		_w2314_
	);
	LUT4 #(
		.INIT('h1000)
	) name1852 (
		_w489_,
		_w673_,
		_w2189_,
		_w2194_,
		_w2315_
	);
	LUT2 #(
		.INIT('h8)
	) name1853 (
		_w599_,
		_w1120_,
		_w2316_
	);
	LUT4 #(
		.INIT('h0057)
	) name1854 (
		\P1_reg2_reg[29]/NET0131 ,
		_w2171_,
		_w2196_,
		_w2316_,
		_w2317_
	);
	LUT2 #(
		.INIT('h4)
	) name1855 (
		_w2315_,
		_w2317_,
		_w2318_
	);
	LUT3 #(
		.INIT('hd0)
	) name1856 (
		_w2170_,
		_w2314_,
		_w2318_,
		_w2319_
	);
	LUT4 #(
		.INIT('h0100)
	) name1857 (
		_w2218_,
		_w2313_,
		_w2266_,
		_w2319_,
		_w2320_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1858 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w2209_,
		_w2320_,
		_w2321_
	);
	LUT2 #(
		.INIT('he)
	) name1859 (
		_w2208_,
		_w2321_,
		_w2322_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1860 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[29]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w2323_
	);
	LUT2 #(
		.INIT('h8)
	) name1861 (
		\P1_reg0_reg[29]/NET0131 ,
		_w2183_,
		_w2324_
	);
	LUT3 #(
		.INIT('h40)
	) name1862 (
		_w2047_,
		_w2048_,
		_w2053_,
		_w2325_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1863 (
		\P1_reg0_reg[29]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w2326_
	);
	LUT4 #(
		.INIT('h0c88)
	) name1864 (
		\P1_reg0_reg[29]/NET0131 ,
		_w1237_,
		_w2217_,
		_w2325_,
		_w2327_
	);
	LUT4 #(
		.INIT('h0c88)
	) name1865 (
		\P1_reg0_reg[29]/NET0131 ,
		_w2121_,
		_w2312_,
		_w2325_,
		_w2328_
	);
	LUT4 #(
		.INIT('h6500)
	) name1866 (
		_w1197_,
		_w2257_,
		_w2264_,
		_w2325_,
		_w2329_
	);
	LUT4 #(
		.INIT('h3c55)
	) name1867 (
		\P1_reg0_reg[29]/NET0131 ,
		_w674_,
		_w2168_,
		_w2325_,
		_w2330_
	);
	LUT4 #(
		.INIT('h1000)
	) name1868 (
		_w489_,
		_w673_,
		_w2194_,
		_w2325_,
		_w2331_
	);
	LUT4 #(
		.INIT('h7f5e)
	) name1869 (
		_w1096_,
		_w1100_,
		_w1098_,
		_w718_,
		_w2332_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1870 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2194_,
		_w2333_
	);
	LUT3 #(
		.INIT('ha2)
	) name1871 (
		\P1_reg0_reg[29]/NET0131 ,
		_w2332_,
		_w2333_,
		_w2334_
	);
	LUT2 #(
		.INIT('h1)
	) name1872 (
		_w2331_,
		_w2334_,
		_w2335_
	);
	LUT3 #(
		.INIT('hd0)
	) name1873 (
		_w2170_,
		_w2330_,
		_w2335_,
		_w2336_
	);
	LUT4 #(
		.INIT('h5700)
	) name1874 (
		_w2128_,
		_w2326_,
		_w2329_,
		_w2336_,
		_w2337_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1875 (
		_w2182_,
		_w2327_,
		_w2328_,
		_w2337_,
		_w2338_
	);
	LUT4 #(
		.INIT('heeec)
	) name1876 (
		\P1_state_reg[0]/NET0131 ,
		_w2323_,
		_w2324_,
		_w2338_,
		_w2339_
	);
	LUT2 #(
		.INIT('h8)
	) name1877 (
		_w1302_,
		_w1305_,
		_w2340_
	);
	LUT4 #(
		.INIT('h7000)
	) name1878 (
		_w1275_,
		_w1283_,
		_w1863_,
		_w1866_,
		_w2341_
	);
	LUT4 #(
		.INIT('h1555)
	) name1879 (
		_w1267_,
		_w1999_,
		_w2341_,
		_w2340_,
		_w2342_
	);
	LUT3 #(
		.INIT('hc4)
	) name1880 (
		\P1_state_reg[0]/NET0131 ,
		\P2_B_reg/NET0131 ,
		_w2342_,
		_w2343_
	);
	LUT4 #(
		.INIT('h2228)
	) name1881 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1264_,
		_w1266_,
		_w2344_
	);
	LUT2 #(
		.INIT('h1)
	) name1882 (
		\P1_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w2345_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1883 (
		\P1_datao_reg[28]/NET0131 ,
		\P1_datao_reg[29]/NET0131 ,
		\si[28]_pad ,
		\si[29]_pad ,
		_w2346_
	);
	LUT3 #(
		.INIT('h10)
	) name1884 (
		_w1356_,
		_w2345_,
		_w2346_,
		_w2347_
	);
	LUT2 #(
		.INIT('h8)
	) name1885 (
		_w1455_,
		_w2347_,
		_w2348_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name1886 (
		_w1307_,
		_w1365_,
		_w2345_,
		_w2346_,
		_w2349_
	);
	LUT2 #(
		.INIT('h8)
	) name1887 (
		\P1_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w2350_
	);
	LUT4 #(
		.INIT('h000b)
	) name1888 (
		_w1454_,
		_w2347_,
		_w2349_,
		_w2350_,
		_w2351_
	);
	LUT3 #(
		.INIT('hb0)
	) name1889 (
		_w1545_,
		_w2348_,
		_w2351_,
		_w2352_
	);
	LUT4 #(
		.INIT('h6a9a)
	) name1890 (
		\P1_datao_reg[31]/NET0131 ,
		\si[31]_pad ,
		_w568_,
		_w2352_,
		_w2353_
	);
	LUT2 #(
		.INIT('h4)
	) name1891 (
		_w1306_,
		_w2353_,
		_w2354_
	);
	LUT3 #(
		.INIT('h23)
	) name1892 (
		_w1306_,
		_w1967_,
		_w2353_,
		_w2355_
	);
	LUT3 #(
		.INIT('h10)
	) name1893 (
		_w1356_,
		_w1357_,
		_w2346_,
		_w2356_
	);
	LUT2 #(
		.INIT('h8)
	) name1894 (
		_w1488_,
		_w2356_,
		_w2357_
	);
	LUT4 #(
		.INIT('h137f)
	) name1895 (
		\P1_datao_reg[28]/NET0131 ,
		\P1_datao_reg[29]/NET0131 ,
		\si[28]_pad ,
		\si[29]_pad ,
		_w2358_
	);
	LUT4 #(
		.INIT('hef00)
	) name1896 (
		_w1356_,
		_w1405_,
		_w2346_,
		_w2358_,
		_w2359_
	);
	LUT3 #(
		.INIT('hb0)
	) name1897 (
		_w1487_,
		_w2356_,
		_w2359_,
		_w2360_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1898 (
		_w1489_,
		_w1558_,
		_w2357_,
		_w2360_,
		_w2361_
	);
	LUT4 #(
		.INIT('h9565)
	) name1899 (
		\P1_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w568_,
		_w2361_,
		_w2362_
	);
	LUT2 #(
		.INIT('h1)
	) name1900 (
		_w1306_,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('h1)
	) name1901 (
		_w1967_,
		_w1993_,
		_w2364_
	);
	LUT3 #(
		.INIT('h01)
	) name1902 (
		_w1306_,
		_w2362_,
		_w2364_,
		_w2365_
	);
	LUT2 #(
		.INIT('h1)
	) name1903 (
		_w2355_,
		_w2365_,
		_w2366_
	);
	LUT4 #(
		.INIT('h0001)
	) name1904 (
		_w1402_,
		_w1933_,
		_w2355_,
		_w2365_,
		_w2367_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1905 (
		_w1306_,
		_w1505_,
		_w1510_,
		_w1957_,
		_w2368_
	);
	LUT3 #(
		.INIT('h0e)
	) name1906 (
		_w1534_,
		_w1542_,
		_w1953_,
		_w2369_
	);
	LUT4 #(
		.INIT('h0f01)
	) name1907 (
		_w1534_,
		_w1542_,
		_w1937_,
		_w1953_,
		_w2370_
	);
	LUT4 #(
		.INIT('h1505)
	) name1908 (
		_w1934_,
		_w1936_,
		_w2368_,
		_w2370_,
		_w2371_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1909 (
		_w1306_,
		_w1505_,
		_w1510_,
		_w1934_,
		_w2372_
	);
	LUT3 #(
		.INIT('h07)
	) name1910 (
		_w1534_,
		_w1542_,
		_w1937_,
		_w2373_
	);
	LUT2 #(
		.INIT('h8)
	) name1911 (
		_w2372_,
		_w2373_,
		_w2374_
	);
	LUT2 #(
		.INIT('h1)
	) name1912 (
		_w1940_,
		_w1942_,
		_w2375_
	);
	LUT3 #(
		.INIT('h0d)
	) name1913 (
		_w1928_,
		_w1943_,
		_w1948_,
		_w2376_
	);
	LUT2 #(
		.INIT('h1)
	) name1914 (
		_w1947_,
		_w1950_,
		_w2377_
	);
	LUT3 #(
		.INIT('h54)
	) name1915 (
		_w1940_,
		_w1947_,
		_w1950_,
		_w2378_
	);
	LUT3 #(
		.INIT('h0d)
	) name1916 (
		_w2375_,
		_w2376_,
		_w2378_,
		_w2379_
	);
	LUT2 #(
		.INIT('h1)
	) name1917 (
		_w1909_,
		_w1943_,
		_w2380_
	);
	LUT4 #(
		.INIT('h0001)
	) name1918 (
		_w1909_,
		_w1940_,
		_w1942_,
		_w1943_,
		_w2381_
	);
	LUT4 #(
		.INIT('heee0)
	) name1919 (
		_w1612_,
		_w1617_,
		_w1802_,
		_w1807_,
		_w2382_
	);
	LUT4 #(
		.INIT('h1117)
	) name1920 (
		_w1612_,
		_w1617_,
		_w1802_,
		_w1807_,
		_w2383_
	);
	LUT3 #(
		.INIT('h10)
	) name1921 (
		_w1910_,
		_w1911_,
		_w2383_,
		_w2384_
	);
	LUT3 #(
		.INIT('h54)
	) name1922 (
		_w1910_,
		_w1924_,
		_w1929_,
		_w2385_
	);
	LUT2 #(
		.INIT('h1)
	) name1923 (
		_w2384_,
		_w2385_,
		_w2386_
	);
	LUT3 #(
		.INIT('ha8)
	) name1924 (
		_w2381_,
		_w2384_,
		_w2385_,
		_w2387_
	);
	LUT2 #(
		.INIT('h2)
	) name1925 (
		_w2379_,
		_w2387_,
		_w2388_
	);
	LUT4 #(
		.INIT('h1151)
	) name1926 (
		_w2371_,
		_w2374_,
		_w2379_,
		_w2387_,
		_w2389_
	);
	LUT2 #(
		.INIT('h2)
	) name1927 (
		_w2367_,
		_w2389_,
		_w2390_
	);
	LUT4 #(
		.INIT('h0777)
	) name1928 (
		_w1812_,
		_w1820_,
		_w1825_,
		_w1830_,
		_w2391_
	);
	LUT4 #(
		.INIT('heee0)
	) name1929 (
		_w1752_,
		_w1759_,
		_w1834_,
		_w1839_,
		_w2392_
	);
	LUT4 #(
		.INIT('h011f)
	) name1930 (
		_w1752_,
		_w1759_,
		_w1834_,
		_w1839_,
		_w2393_
	);
	LUT4 #(
		.INIT('heee0)
	) name1931 (
		_w1812_,
		_w1820_,
		_w1825_,
		_w1830_,
		_w2394_
	);
	LUT4 #(
		.INIT('h1117)
	) name1932 (
		_w1812_,
		_w1820_,
		_w1825_,
		_w1830_,
		_w2395_
	);
	LUT3 #(
		.INIT('h07)
	) name1933 (
		_w2391_,
		_w2393_,
		_w2395_,
		_w2396_
	);
	LUT4 #(
		.INIT('h0777)
	) name1934 (
		_w1752_,
		_w1759_,
		_w1834_,
		_w1839_,
		_w2397_
	);
	LUT2 #(
		.INIT('h8)
	) name1935 (
		_w2391_,
		_w2397_,
		_w2398_
	);
	LUT3 #(
		.INIT('h07)
	) name1936 (
		_w1740_,
		_w1747_,
		_w1872_,
		_w2399_
	);
	LUT3 #(
		.INIT('h0e)
	) name1937 (
		_w1874_,
		_w1902_,
		_w1906_,
		_w2400_
	);
	LUT3 #(
		.INIT('h0e)
	) name1938 (
		_w1740_,
		_w1747_,
		_w1873_,
		_w2401_
	);
	LUT3 #(
		.INIT('h71)
	) name1939 (
		_w1740_,
		_w1747_,
		_w1873_,
		_w2402_
	);
	LUT3 #(
		.INIT('h07)
	) name1940 (
		_w2399_,
		_w2400_,
		_w2402_,
		_w2403_
	);
	LUT3 #(
		.INIT('ha2)
	) name1941 (
		_w2396_,
		_w2398_,
		_w2403_,
		_w2404_
	);
	LUT2 #(
		.INIT('h1)
	) name1942 (
		_w1880_,
		_w1894_,
		_w2405_
	);
	LUT2 #(
		.INIT('h1)
	) name1943 (
		_w1885_,
		_w1895_,
		_w2406_
	);
	LUT3 #(
		.INIT('hb2)
	) name1944 (
		_w1648_,
		_w1653_,
		_w1882_,
		_w2407_
	);
	LUT3 #(
		.INIT('h0d)
	) name1945 (
		_w1883_,
		_w1886_,
		_w1891_,
		_w2408_
	);
	LUT3 #(
		.INIT('hd0)
	) name1946 (
		_w1888_,
		_w2407_,
		_w2408_,
		_w2409_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1947 (
		_w1888_,
		_w2406_,
		_w2407_,
		_w2408_,
		_w2410_
	);
	LUT3 #(
		.INIT('h0d)
	) name1948 (
		_w1890_,
		_w1895_,
		_w1899_,
		_w2411_
	);
	LUT3 #(
		.INIT('h54)
	) name1949 (
		_w1880_,
		_w1898_,
		_w1903_,
		_w2412_
	);
	LUT4 #(
		.INIT('h0075)
	) name1950 (
		_w2405_,
		_w2410_,
		_w2411_,
		_w2412_,
		_w2413_
	);
	LUT2 #(
		.INIT('h1)
	) name1951 (
		_w1879_,
		_w1906_,
		_w2414_
	);
	LUT4 #(
		.INIT('h0e08)
	) name1952 (
		_w1779_,
		_w1788_,
		_w1873_,
		_w1879_,
		_w2415_
	);
	LUT3 #(
		.INIT('h51)
	) name1953 (
		_w1876_,
		_w2399_,
		_w2415_,
		_w2416_
	);
	LUT4 #(
		.INIT('h0323)
	) name1954 (
		_w1919_,
		_w1921_,
		_w2391_,
		_w2397_,
		_w2417_
	);
	LUT3 #(
		.INIT('ha8)
	) name1955 (
		_w2396_,
		_w2416_,
		_w2417_,
		_w2418_
	);
	LUT4 #(
		.INIT('h0777)
	) name1956 (
		_w1612_,
		_w1617_,
		_w1802_,
		_w1807_,
		_w2419_
	);
	LUT3 #(
		.INIT('h10)
	) name1957 (
		_w1910_,
		_w1911_,
		_w2419_,
		_w2420_
	);
	LUT4 #(
		.INIT('h5700)
	) name1958 (
		_w2396_,
		_w2416_,
		_w2417_,
		_w2420_,
		_w2421_
	);
	LUT3 #(
		.INIT('h70)
	) name1959 (
		_w2404_,
		_w2413_,
		_w2421_,
		_w2422_
	);
	LUT3 #(
		.INIT('h80)
	) name1960 (
		_w2372_,
		_w2373_,
		_w2381_,
		_w2423_
	);
	LUT2 #(
		.INIT('h8)
	) name1961 (
		_w2367_,
		_w2423_,
		_w2424_
	);
	LUT3 #(
		.INIT('h54)
	) name1962 (
		_w1402_,
		_w1403_,
		_w1956_,
		_w2425_
	);
	LUT3 #(
		.INIT('h32)
	) name1963 (
		_w1306_,
		_w1993_,
		_w2362_,
		_w2426_
	);
	LUT4 #(
		.INIT('h3031)
	) name1964 (
		_w1306_,
		_w1967_,
		_w1993_,
		_w2362_,
		_w2427_
	);
	LUT2 #(
		.INIT('h2)
	) name1965 (
		_w2354_,
		_w2427_,
		_w2428_
	);
	LUT3 #(
		.INIT('h07)
	) name1966 (
		_w2425_,
		_w2366_,
		_w2428_,
		_w2429_
	);
	LUT3 #(
		.INIT('h70)
	) name1967 (
		_w2422_,
		_w2424_,
		_w2429_,
		_w2430_
	);
	LUT2 #(
		.INIT('h2)
	) name1968 (
		_w1864_,
		_w1866_,
		_w2431_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1969 (
		_w1595_,
		_w2390_,
		_w2430_,
		_w2431_,
		_w2432_
	);
	LUT3 #(
		.INIT('h40)
	) name1970 (
		_w1306_,
		_w1967_,
		_w2353_,
		_w2433_
	);
	LUT3 #(
		.INIT('h04)
	) name1971 (
		_w1306_,
		_w1993_,
		_w2362_,
		_w2434_
	);
	LUT2 #(
		.INIT('h1)
	) name1972 (
		_w2355_,
		_w2434_,
		_w2435_
	);
	LUT4 #(
		.INIT('h00e8)
	) name1973 (
		_w1374_,
		_w1400_,
		_w1933_,
		_w2426_,
		_w2436_
	);
	LUT3 #(
		.INIT('h51)
	) name1974 (
		_w2433_,
		_w2435_,
		_w2436_,
		_w2437_
	);
	LUT2 #(
		.INIT('h1)
	) name1975 (
		_w2433_,
		_w2426_,
		_w2438_
	);
	LUT4 #(
		.INIT('h0001)
	) name1976 (
		_w1403_,
		_w1956_,
		_w2433_,
		_w2426_,
		_w2439_
	);
	LUT2 #(
		.INIT('h8)
	) name1977 (
		_w2368_,
		_w2369_,
		_w2440_
	);
	LUT2 #(
		.INIT('h8)
	) name1978 (
		_w2439_,
		_w2440_,
		_w2441_
	);
	LUT3 #(
		.INIT('h70)
	) name1979 (
		_w1654_,
		_w1655_,
		_w1660_,
		_w2442_
	);
	LUT4 #(
		.INIT('h020b)
	) name1980 (
		_w1648_,
		_w1653_,
		_w1883_,
		_w2442_,
		_w2443_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1981 (
		_w1888_,
		_w1892_,
		_w2406_,
		_w2443_,
		_w2444_
	);
	LUT3 #(
		.INIT('h01)
	) name1982 (
		_w1874_,
		_w1902_,
		_w1903_,
		_w2445_
	);
	LUT4 #(
		.INIT('h8000)
	) name1983 (
		_w2392_,
		_w2394_,
		_w2401_,
		_w2445_,
		_w2446_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1984 (
		_w1900_,
		_w2405_,
		_w2444_,
		_w2446_,
		_w2447_
	);
	LUT3 #(
		.INIT('h01)
	) name1985 (
		_w1928_,
		_w1929_,
		_w1948_,
		_w2448_
	);
	LUT2 #(
		.INIT('h4)
	) name1986 (
		_w1924_,
		_w2382_,
		_w2449_
	);
	LUT3 #(
		.INIT('h80)
	) name1987 (
		_w2377_,
		_w2448_,
		_w2449_,
		_w2450_
	);
	LUT3 #(
		.INIT('he0)
	) name1988 (
		_w2418_,
		_w2447_,
		_w2450_,
		_w2451_
	);
	LUT3 #(
		.INIT('h15)
	) name1989 (
		_w2437_,
		_w2441_,
		_w2451_,
		_w2452_
	);
	LUT4 #(
		.INIT('h00e8)
	) name1990 (
		_w1569_,
		_w1573_,
		_w1909_,
		_w1947_,
		_w2453_
	);
	LUT3 #(
		.INIT('h51)
	) name1991 (
		_w1950_,
		_w2375_,
		_w2453_,
		_w2454_
	);
	LUT4 #(
		.INIT('h1101)
	) name1992 (
		_w1910_,
		_w1911_,
		_w1925_,
		_w2419_,
		_w2455_
	);
	LUT3 #(
		.INIT('h08)
	) name1993 (
		_w2377_,
		_w2448_,
		_w2455_,
		_w2456_
	);
	LUT4 #(
		.INIT('h8880)
	) name1994 (
		_w2439_,
		_w2440_,
		_w2454_,
		_w2456_,
		_w2457_
	);
	LUT3 #(
		.INIT('hc4)
	) name1995 (
		_w1954_,
		_w2372_,
		_w2373_,
		_w2458_
	);
	LUT3 #(
		.INIT('h04)
	) name1996 (
		_w1957_,
		_w2439_,
		_w2458_,
		_w2459_
	);
	LUT2 #(
		.INIT('h1)
	) name1997 (
		_w2457_,
		_w2459_,
		_w2460_
	);
	LUT4 #(
		.INIT('h8421)
	) name1998 (
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		_w1272_,
		_w1862_,
		_w2461_
	);
	LUT2 #(
		.INIT('h4)
	) name1999 (
		_w1866_,
		_w2461_,
		_w2462_
	);
	LUT4 #(
		.INIT('h9500)
	) name2000 (
		_w1595_,
		_w2452_,
		_w2460_,
		_w2462_,
		_w2463_
	);
	LUT2 #(
		.INIT('h8)
	) name2001 (
		_w2381_,
		_w2420_,
		_w2464_
	);
	LUT4 #(
		.INIT('h0080)
	) name2002 (
		_w2399_,
		_w2414_,
		_w2398_,
		_w2413_,
		_w2465_
	);
	LUT4 #(
		.INIT('h22a2)
	) name2003 (
		_w2388_,
		_w2464_,
		_w2404_,
		_w2465_,
		_w2466_
	);
	LUT4 #(
		.INIT('h0001)
	) name2004 (
		_w1402_,
		_w1933_,
		_w2355_,
		_w2434_,
		_w2467_
	);
	LUT2 #(
		.INIT('h8)
	) name2005 (
		_w2467_,
		_w2374_,
		_w2468_
	);
	LUT2 #(
		.INIT('h8)
	) name2006 (
		_w2371_,
		_w2467_,
		_w2469_
	);
	LUT4 #(
		.INIT('h0071)
	) name2007 (
		_w1374_,
		_w1400_,
		_w1956_,
		_w2434_,
		_w2470_
	);
	LUT3 #(
		.INIT('h51)
	) name2008 (
		_w2355_,
		_w2438_,
		_w2470_,
		_w2471_
	);
	LUT2 #(
		.INIT('h1)
	) name2009 (
		_w2469_,
		_w2471_,
		_w2472_
	);
	LUT4 #(
		.INIT('h4500)
	) name2010 (
		\P2_B_reg/NET0131 ,
		_w2466_,
		_w2468_,
		_w2472_,
		_w2473_
	);
	LUT4 #(
		.INIT('h2184)
	) name2011 (
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		_w1272_,
		_w1862_,
		_w2474_
	);
	LUT3 #(
		.INIT('h80)
	) name2012 (
		_w1595_,
		_w1866_,
		_w2474_,
		_w2475_
	);
	LUT4 #(
		.INIT('h0045)
	) name2013 (
		_w2463_,
		_w2473_,
		_w2475_,
		_w2432_,
		_w2476_
	);
	LUT4 #(
		.INIT('h1411)
	) name2014 (
		\P2_B_reg/NET0131 ,
		_w1595_,
		_w2390_,
		_w2430_,
		_w2477_
	);
	LUT3 #(
		.INIT('h80)
	) name2015 (
		_w1859_,
		_w1863_,
		_w1866_,
		_w2478_
	);
	LUT2 #(
		.INIT('h4)
	) name2016 (
		_w2477_,
		_w2478_,
		_w2479_
	);
	LUT4 #(
		.INIT('hc888)
	) name2017 (
		\P2_B_reg/NET0131 ,
		_w1867_,
		_w2452_,
		_w2460_,
		_w2480_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2018 (
		_w1868_,
		_w2466_,
		_w2468_,
		_w2472_,
		_w2481_
	);
	LUT3 #(
		.INIT('ha8)
	) name2019 (
		_w2028_,
		_w2480_,
		_w2481_,
		_w2482_
	);
	LUT4 #(
		.INIT('h7778)
	) name2020 (
		_w1761_,
		_w1763_,
		_w1769_,
		_w1773_,
		_w2483_
	);
	LUT4 #(
		.INIT('h7778)
	) name2021 (
		_w1777_,
		_w1778_,
		_w1783_,
		_w1787_,
		_w2484_
	);
	LUT3 #(
		.INIT('h87)
	) name2022 (
		_w1709_,
		_w1711_,
		_w1717_,
		_w2485_
	);
	LUT3 #(
		.INIT('h87)
	) name2023 (
		_w1673_,
		_w1674_,
		_w1681_,
		_w2486_
	);
	LUT3 #(
		.INIT('h87)
	) name2024 (
		_w1636_,
		_w1637_,
		_w1643_,
		_w2487_
	);
	LUT3 #(
		.INIT('h95)
	) name2025 (
		_w1666_,
		_w1667_,
		_w1669_,
		_w2488_
	);
	LUT4 #(
		.INIT('h4000)
	) name2026 (
		_w2485_,
		_w2486_,
		_w2487_,
		_w2488_,
		_w2489_
	);
	LUT4 #(
		.INIT('h0200)
	) name2027 (
		_w1915_,
		_w2484_,
		_w2483_,
		_w2489_,
		_w2490_
	);
	LUT2 #(
		.INIT('h9)
	) name2028 (
		_w1802_,
		_w1807_,
		_w2491_
	);
	LUT2 #(
		.INIT('h2)
	) name2029 (
		_w1919_,
		_w2491_,
		_w2492_
	);
	LUT2 #(
		.INIT('h9)
	) name2030 (
		_w1812_,
		_w1820_,
		_w2493_
	);
	LUT2 #(
		.INIT('h9)
	) name2031 (
		_w1752_,
		_w1759_,
		_w2494_
	);
	LUT2 #(
		.INIT('h9)
	) name2032 (
		_w1740_,
		_w1747_,
		_w2495_
	);
	LUT3 #(
		.INIT('h87)
	) name2033 (
		_w1697_,
		_w1699_,
		_w1706_,
		_w2496_
	);
	LUT3 #(
		.INIT('h78)
	) name2034 (
		_w1720_,
		_w1721_,
		_w1726_,
		_w2497_
	);
	LUT3 #(
		.INIT('h10)
	) name2035 (
		_w2442_,
		_w2496_,
		_w2497_,
		_w2498_
	);
	LUT3 #(
		.INIT('h87)
	) name2036 (
		_w1688_,
		_w1690_,
		_w1695_,
		_w2499_
	);
	LUT3 #(
		.INIT('h87)
	) name2037 (
		_w1646_,
		_w1647_,
		_w1653_,
		_w2500_
	);
	LUT3 #(
		.INIT('h10)
	) name2038 (
		_w1882_,
		_w2499_,
		_w2500_,
		_w2501_
	);
	LUT4 #(
		.INIT('h1000)
	) name2039 (
		_w2495_,
		_w2494_,
		_w2498_,
		_w2501_,
		_w2502_
	);
	LUT4 #(
		.INIT('h4000)
	) name2040 (
		_w2493_,
		_w2502_,
		_w2490_,
		_w2492_,
		_w2503_
	);
	LUT4 #(
		.INIT('h23dc)
	) name2041 (
		_w1306_,
		_w1596_,
		_w1598_,
		_w1604_,
		_w2504_
	);
	LUT3 #(
		.INIT('h1e)
	) name2042 (
		_w1306_,
		_w1546_,
		_w1551_,
		_w2505_
	);
	LUT2 #(
		.INIT('h1)
	) name2043 (
		_w2504_,
		_w2505_,
		_w2506_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2044 (
		_w1306_,
		_w1555_,
		_w1559_,
		_w1564_,
		_w2507_
	);
	LUT2 #(
		.INIT('h9)
	) name2045 (
		_w1612_,
		_w1617_,
		_w2508_
	);
	LUT3 #(
		.INIT('h1e)
	) name2046 (
		_w1306_,
		_w1568_,
		_w1573_,
		_w2509_
	);
	LUT3 #(
		.INIT('h1e)
	) name2047 (
		_w1306_,
		_w1586_,
		_w1592_,
		_w2510_
	);
	LUT2 #(
		.INIT('h9)
	) name2048 (
		_w1626_,
		_w1631_,
		_w2511_
	);
	LUT4 #(
		.INIT('h0001)
	) name2049 (
		_w2508_,
		_w2509_,
		_w2510_,
		_w2511_,
		_w2512_
	);
	LUT2 #(
		.INIT('h4)
	) name2050 (
		_w2507_,
		_w2512_,
		_w2513_
	);
	LUT3 #(
		.INIT('h1e)
	) name2051 (
		_w1306_,
		_w1505_,
		_w1510_,
		_w2514_
	);
	LUT2 #(
		.INIT('h2)
	) name2052 (
		_w1404_,
		_w2514_,
		_w2515_
	);
	LUT4 #(
		.INIT('h8000)
	) name2053 (
		_w2503_,
		_w2506_,
		_w2513_,
		_w2515_,
		_w2516_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2054 (
		_w1306_,
		_w1452_,
		_w1478_,
		_w1483_,
		_w2517_
	);
	LUT2 #(
		.INIT('h9)
	) name2055 (
		_w1534_,
		_w1542_,
		_w2518_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2056 (
		_w1306_,
		_w1514_,
		_w1521_,
		_w1527_,
		_w2519_
	);
	LUT4 #(
		.INIT('h0006)
	) name2057 (
		_w1534_,
		_w1542_,
		_w2519_,
		_w2517_,
		_w2520_
	);
	LUT3 #(
		.INIT('h10)
	) name2058 (
		_w2355_,
		_w2434_,
		_w2520_,
		_w2521_
	);
	LUT3 #(
		.INIT('h1e)
	) name2059 (
		_w1306_,
		_w1441_,
		_w1449_,
		_w2522_
	);
	LUT3 #(
		.INIT('h01)
	) name2060 (
		_w2433_,
		_w2426_,
		_w2522_,
		_w2523_
	);
	LUT2 #(
		.INIT('h8)
	) name2061 (
		_w2521_,
		_w2523_,
		_w2524_
	);
	LUT4 #(
		.INIT('h4888)
	) name2062 (
		_w1595_,
		_w1859_,
		_w2516_,
		_w2524_,
		_w2525_
	);
	LUT4 #(
		.INIT('h2228)
	) name2063 (
		\P2_B_reg/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		_w1272_,
		_w1865_,
		_w2526_
	);
	LUT2 #(
		.INIT('h4)
	) name2064 (
		_w2028_,
		_w2526_,
		_w2527_
	);
	LUT3 #(
		.INIT('h54)
	) name2065 (
		_w1863_,
		_w2525_,
		_w2527_,
		_w2528_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2066 (
		_w2024_,
		_w2466_,
		_w2468_,
		_w2472_,
		_w2529_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name2067 (
		\P2_B_reg/NET0131 ,
		_w2000_,
		_w2452_,
		_w2460_,
		_w2530_
	);
	LUT3 #(
		.INIT('h01)
	) name2068 (
		_w2528_,
		_w2529_,
		_w2530_,
		_w2531_
	);
	LUT4 #(
		.INIT('h1000)
	) name2069 (
		_w2482_,
		_w2479_,
		_w2531_,
		_w2476_,
		_w2532_
	);
	LUT3 #(
		.INIT('hae)
	) name2070 (
		_w2343_,
		_w2344_,
		_w2532_,
		_w2533_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2071 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[29]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w2534_
	);
	LUT2 #(
		.INIT('h8)
	) name2072 (
		\P1_reg1_reg[29]/NET0131 ,
		_w2183_,
		_w2535_
	);
	LUT3 #(
		.INIT('hb0)
	) name2073 (
		_w2047_,
		_w2048_,
		_w2053_,
		_w2536_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2074 (
		\P1_reg1_reg[29]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w2537_
	);
	LUT4 #(
		.INIT('h0c88)
	) name2075 (
		\P1_reg1_reg[29]/NET0131 ,
		_w1237_,
		_w2217_,
		_w2536_,
		_w2538_
	);
	LUT4 #(
		.INIT('h6500)
	) name2076 (
		_w1197_,
		_w2257_,
		_w2264_,
		_w2536_,
		_w2539_
	);
	LUT3 #(
		.INIT('ha8)
	) name2077 (
		_w2128_,
		_w2537_,
		_w2539_,
		_w2540_
	);
	LUT4 #(
		.INIT('h0c88)
	) name2078 (
		\P1_reg1_reg[29]/NET0131 ,
		_w2121_,
		_w2312_,
		_w2536_,
		_w2541_
	);
	LUT4 #(
		.INIT('h3c55)
	) name2079 (
		\P1_reg1_reg[29]/NET0131 ,
		_w674_,
		_w2168_,
		_w2536_,
		_w2542_
	);
	LUT4 #(
		.INIT('h1000)
	) name2080 (
		_w489_,
		_w673_,
		_w2194_,
		_w2536_,
		_w2543_
	);
	LUT4 #(
		.INIT('hef00)
	) name2081 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2194_,
		_w2544_
	);
	LUT3 #(
		.INIT('ha2)
	) name2082 (
		\P1_reg1_reg[29]/NET0131 ,
		_w2332_,
		_w2544_,
		_w2545_
	);
	LUT2 #(
		.INIT('h1)
	) name2083 (
		_w2543_,
		_w2545_,
		_w2546_
	);
	LUT3 #(
		.INIT('hd0)
	) name2084 (
		_w2170_,
		_w2542_,
		_w2546_,
		_w2547_
	);
	LUT4 #(
		.INIT('h0100)
	) name2085 (
		_w2538_,
		_w2541_,
		_w2540_,
		_w2547_,
		_w2548_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2086 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w2535_,
		_w2548_,
		_w2549_
	);
	LUT2 #(
		.INIT('he)
	) name2087 (
		_w2534_,
		_w2549_,
		_w2550_
	);
	LUT4 #(
		.INIT('h0c84)
	) name2088 (
		_w2022_,
		_w2025_,
		_w2354_,
		_w2363_,
		_w2551_
	);
	LUT3 #(
		.INIT('h40)
	) name2089 (
		_w1306_,
		_w2001_,
		_w2353_,
		_w2552_
	);
	LUT4 #(
		.INIT('hef00)
	) name2090 (
		_w1397_,
		_w1965_,
		_w1966_,
		_w2000_,
		_w2553_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2091 (
		_w1995_,
		_w1997_,
		_w2552_,
		_w2553_,
		_w2554_
	);
	LUT4 #(
		.INIT('h1311)
	) name2092 (
		_w1298_,
		_w2030_,
		_w2551_,
		_w2554_,
		_w2555_
	);
	LUT4 #(
		.INIT('h0222)
	) name2093 (
		\P1_state_reg[0]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w2556_
	);
	LUT4 #(
		.INIT('hce00)
	) name2094 (
		_w1298_,
		_w2029_,
		_w2032_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h2)
	) name2095 (
		\P2_reg2_reg[31]/NET0131 ,
		_w2557_,
		_w2558_
	);
	LUT3 #(
		.INIT('hf4)
	) name2096 (
		_w2555_,
		_w2556_,
		_w2558_,
		_w2559_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2097 (
		\P1_reg3_reg[24]/NET0131 ,
		_w785_,
		_w597_,
		_w2183_,
		_w2560_
	);
	LUT2 #(
		.INIT('h2)
	) name2098 (
		_w1074_,
		_w2055_,
		_w2561_
	);
	LUT3 #(
		.INIT('h40)
	) name2099 (
		_w2082_,
		_w2085_,
		_w2092_,
		_w2562_
	);
	LUT4 #(
		.INIT('h40cc)
	) name2100 (
		_w2065_,
		_w2088_,
		_w2091_,
		_w2096_,
		_w2563_
	);
	LUT2 #(
		.INIT('h2)
	) name2101 (
		_w2101_,
		_w2563_,
		_w2564_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2102 (
		_w2108_,
		_w2112_,
		_w2562_,
		_w2564_,
		_w2565_
	);
	LUT4 #(
		.INIT('h070b)
	) name2103 (
		_w1210_,
		_w2055_,
		_w2561_,
		_w2565_,
		_w2566_
	);
	LUT4 #(
		.INIT('h6555)
	) name2104 (
		_w1063_,
		_w1079_,
		_w2142_,
		_w2213_,
		_w2567_
	);
	LUT4 #(
		.INIT('h7020)
	) name2105 (
		_w488_,
		_w789_,
		_w2055_,
		_w2567_,
		_w2568_
	);
	LUT3 #(
		.INIT('ha8)
	) name2106 (
		_w1237_,
		_w2561_,
		_w2568_,
		_w2569_
	);
	LUT4 #(
		.INIT('h5d00)
	) name2107 (
		_w870_,
		_w872_,
		_w922_,
		_w1023_,
		_w2570_
	);
	LUT3 #(
		.INIT('hc4)
	) name2108 (
		_w772_,
		_w1021_,
		_w2570_,
		_w2571_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2109 (
		_w817_,
		_w872_,
		_w1019_,
		_w1024_,
		_w2572_
	);
	LUT4 #(
		.INIT('h8488)
	) name2110 (
		_w1210_,
		_w2055_,
		_w2571_,
		_w2572_,
		_w2573_
	);
	LUT3 #(
		.INIT('h80)
	) name2111 (
		_w2155_,
		_w2163_,
		_w2164_,
		_w2574_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2112 (
		_w783_,
		_w1073_,
		_w2155_,
		_w2163_,
		_w2575_
	);
	LUT4 #(
		.INIT('h3331)
	) name2113 (
		_w2055_,
		_w2561_,
		_w2574_,
		_w2575_,
		_w2576_
	);
	LUT3 #(
		.INIT('h20)
	) name2114 (
		_w1073_,
		_w2175_,
		_w2176_,
		_w2577_
	);
	LUT4 #(
		.INIT('h5400)
	) name2115 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2194_,
		_w2578_
	);
	LUT3 #(
		.INIT('ha8)
	) name2116 (
		_w1074_,
		_w2171_,
		_w2578_,
		_w2579_
	);
	LUT2 #(
		.INIT('h1)
	) name2117 (
		_w2577_,
		_w2579_,
		_w2580_
	);
	LUT3 #(
		.INIT('hd0)
	) name2118 (
		_w2170_,
		_w2576_,
		_w2580_,
		_w2581_
	);
	LUT4 #(
		.INIT('h5700)
	) name2119 (
		_w2128_,
		_w2561_,
		_w2573_,
		_w2581_,
		_w2582_
	);
	LUT4 #(
		.INIT('h3100)
	) name2120 (
		_w2121_,
		_w2569_,
		_w2566_,
		_w2582_,
		_w2583_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2121 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w2560_,
		_w2583_,
		_w2584_
	);
	LUT2 #(
		.INIT('h2)
	) name2122 (
		\P1_reg3_reg[24]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2585_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2123 (
		\P1_reg3_reg[24]/NET0131 ,
		_w785_,
		_w597_,
		_w1244_,
		_w2586_
	);
	LUT2 #(
		.INIT('h1)
	) name2124 (
		_w2585_,
		_w2586_,
		_w2587_
	);
	LUT2 #(
		.INIT('hb)
	) name2125 (
		_w2584_,
		_w2587_,
		_w2588_
	);
	LUT2 #(
		.INIT('h2)
	) name2126 (
		\P2_reg2_reg[27]/NET0131 ,
		_w1298_,
		_w2589_
	);
	LUT2 #(
		.INIT('h8)
	) name2127 (
		_w1938_,
		_w1941_,
		_w2590_
	);
	LUT4 #(
		.INIT('h0001)
	) name2128 (
		_w1872_,
		_w1879_,
		_w1880_,
		_w1906_,
		_w2591_
	);
	LUT3 #(
		.INIT('h15)
	) name2129 (
		_w1875_,
		_w1904_,
		_w1907_,
		_w2592_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2130 (
		_w1897_,
		_w1901_,
		_w2591_,
		_w2592_,
		_w2593_
	);
	LUT2 #(
		.INIT('h8)
	) name2131 (
		_w1871_,
		_w1915_,
		_w2594_
	);
	LUT3 #(
		.INIT('h0b)
	) name2132 (
		_w1877_,
		_w1915_,
		_w1920_,
		_w2595_
	);
	LUT2 #(
		.INIT('h8)
	) name2133 (
		_w1912_,
		_w1914_,
		_w2596_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2134 (
		_w2593_,
		_w2594_,
		_w2595_,
		_w2596_,
		_w2597_
	);
	LUT3 #(
		.INIT('h0d)
	) name2135 (
		_w1912_,
		_w1922_,
		_w1926_,
		_w2598_
	);
	LUT4 #(
		.INIT('h0001)
	) name2136 (
		_w1909_,
		_w1910_,
		_w1942_,
		_w1943_,
		_w2599_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2137 (
		_w2590_,
		_w2597_,
		_w2598_,
		_w2599_,
		_w2600_
	);
	LUT3 #(
		.INIT('h07)
	) name2138 (
		_w1930_,
		_w1944_,
		_w1949_,
		_w2601_
	);
	LUT3 #(
		.INIT('h0d)
	) name2139 (
		_w1938_,
		_w1951_,
		_w1955_,
		_w2602_
	);
	LUT3 #(
		.INIT('hd0)
	) name2140 (
		_w2590_,
		_w2601_,
		_w2602_,
		_w2603_
	);
	LUT4 #(
		.INIT('h8288)
	) name2141 (
		_w1298_,
		_w2517_,
		_w2600_,
		_w2603_,
		_w2604_
	);
	LUT3 #(
		.INIT('ha8)
	) name2142 (
		_w1963_,
		_w2589_,
		_w2604_,
		_w2605_
	);
	LUT3 #(
		.INIT('h8a)
	) name2143 (
		_w1576_,
		_w1851_,
		_w1854_,
		_w2606_
	);
	LUT3 #(
		.INIT('h45)
	) name2144 (
		_w1529_,
		_w1534_,
		_w1542_,
		_w2607_
	);
	LUT4 #(
		.INIT('h0045)
	) name2145 (
		_w1529_,
		_w1534_,
		_w1542_,
		_w1553_,
		_w2608_
	);
	LUT4 #(
		.INIT('h7500)
	) name2146 (
		_w1576_,
		_w1851_,
		_w1854_,
		_w2608_,
		_w2609_
	);
	LUT4 #(
		.INIT('h4504)
	) name2147 (
		_w1529_,
		_w1534_,
		_w1542_,
		_w1577_,
		_w2610_
	);
	LUT2 #(
		.INIT('h2)
	) name2148 (
		_w1581_,
		_w2610_,
		_w2611_
	);
	LUT3 #(
		.INIT('h45)
	) name2149 (
		_w1512_,
		_w2609_,
		_w2611_,
		_w2612_
	);
	LUT4 #(
		.INIT('h0001)
	) name2150 (
		_w1696_,
		_w1707_,
		_w1775_,
		_w1789_,
		_w2613_
	);
	LUT4 #(
		.INIT('h2f00)
	) name2151 (
		_w1728_,
		_w1687_,
		_w1732_,
		_w2613_,
		_w2614_
	);
	LUT3 #(
		.INIT('h70)
	) name2152 (
		_w1735_,
		_w1790_,
		_w1795_,
		_w2615_
	);
	LUT2 #(
		.INIT('h8)
	) name2153 (
		_w1634_,
		_w1821_,
		_w2616_
	);
	LUT2 #(
		.INIT('h8)
	) name2154 (
		_w1760_,
		_w1840_,
		_w2617_
	);
	LUT4 #(
		.INIT('h8000)
	) name2155 (
		_w1634_,
		_w1760_,
		_w1821_,
		_w1840_,
		_w2618_
	);
	LUT3 #(
		.INIT('h07)
	) name2156 (
		_w1796_,
		_w1840_,
		_w1843_,
		_w2619_
	);
	LUT3 #(
		.INIT('h0d)
	) name2157 (
		_w1634_,
		_w1844_,
		_w1847_,
		_w2620_
	);
	LUT3 #(
		.INIT('hd0)
	) name2158 (
		_w2616_,
		_w2619_,
		_w2620_,
		_w2621_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2159 (
		_w2614_,
		_w2615_,
		_w2618_,
		_w2621_,
		_w2622_
	);
	LUT4 #(
		.INIT('h0001)
	) name2160 (
		_w1567_,
		_w1594_,
		_w1606_,
		_w1853_,
		_w2623_
	);
	LUT3 #(
		.INIT('h40)
	) name2161 (
		_w1512_,
		_w2608_,
		_w2623_,
		_w2624_
	);
	LUT4 #(
		.INIT('h9a99)
	) name2162 (
		_w2517_,
		_w2612_,
		_w2622_,
		_w2624_,
		_w2625_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2163 (
		\P2_reg2_reg[27]/NET0131 ,
		_w1298_,
		_w1869_,
		_w2625_,
		_w2626_
	);
	LUT2 #(
		.INIT('h2)
	) name2164 (
		_w1305_,
		_w1510_,
		_w2627_
	);
	LUT4 #(
		.INIT('h1000)
	) name2165 (
		_w1483_,
		_w1510_,
		_w1978_,
		_w1987_,
		_w2628_
	);
	LUT4 #(
		.INIT('h1555)
	) name2166 (
		_w1305_,
		_w1988_,
		_w1978_,
		_w1987_,
		_w2629_
	);
	LUT4 #(
		.INIT('h0233)
	) name2167 (
		_w1449_,
		_w2627_,
		_w2628_,
		_w2629_,
		_w2630_
	);
	LUT4 #(
		.INIT('h5400)
	) name2168 (
		_w1306_,
		_w1452_,
		_w1478_,
		_w2001_,
		_w2631_
	);
	LUT4 #(
		.INIT('h8000)
	) name2169 (
		_w2009_,
		_w2010_,
		_w2015_,
		_w2018_,
		_w2632_
	);
	LUT3 #(
		.INIT('h8a)
	) name2170 (
		_w1479_,
		_w1506_,
		_w2632_,
		_w2633_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name2171 (
		_w2021_,
		_w2025_,
		_w2631_,
		_w2633_,
		_w2634_
	);
	LUT3 #(
		.INIT('hd0)
	) name2172 (
		_w2000_,
		_w2630_,
		_w2634_,
		_w2635_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2173 (
		_w1298_,
		_w2000_,
		_w2630_,
		_w2634_,
		_w2636_
	);
	LUT2 #(
		.INIT('h8)
	) name2174 (
		_w1480_,
		_w2029_,
		_w2637_
	);
	LUT4 #(
		.INIT('h1ff3)
	) name2175 (
		_w1595_,
		_w1859_,
		_w1863_,
		_w1866_,
		_w2638_
	);
	LUT3 #(
		.INIT('h0d)
	) name2176 (
		_w1298_,
		_w2032_,
		_w2638_,
		_w2639_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2177 (
		_w1298_,
		_w2001_,
		_w2025_,
		_w2032_,
		_w2640_
	);
	LUT4 #(
		.INIT('h0705)
	) name2178 (
		\P2_reg2_reg[27]/NET0131 ,
		_w2031_,
		_w2637_,
		_w2640_,
		_w2641_
	);
	LUT3 #(
		.INIT('h10)
	) name2179 (
		_w2626_,
		_w2636_,
		_w2641_,
		_w2642_
	);
	LUT4 #(
		.INIT('h2000)
	) name2180 (
		\P2_reg2_reg[27]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w2643_
	);
	LUT4 #(
		.INIT('h0075)
	) name2181 (
		_w1285_,
		_w2605_,
		_w2642_,
		_w2643_,
		_w2644_
	);
	LUT2 #(
		.INIT('h2)
	) name2182 (
		\P2_reg2_reg[27]/NET0131 ,
		_w2042_,
		_w2645_
	);
	LUT3 #(
		.INIT('hf2)
	) name2183 (
		\P1_state_reg[0]/NET0131 ,
		_w2644_,
		_w2645_,
		_w2646_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2184 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[26]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w2647_
	);
	LUT2 #(
		.INIT('h8)
	) name2185 (
		\P1_reg2_reg[26]/NET0131 ,
		_w2183_,
		_w2648_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2186 (
		\P1_reg2_reg[26]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w2649_
	);
	LUT3 #(
		.INIT('h15)
	) name2187 (
		_w767_,
		_w869_,
		_w1022_,
		_w2650_
	);
	LUT4 #(
		.INIT('h0001)
	) name2188 (
		_w906_,
		_w934_,
		_w944_,
		_w1016_,
		_w2651_
	);
	LUT3 #(
		.INIT('h15)
	) name2189 (
		_w917_,
		_w1013_,
		_w1017_,
		_w2652_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2190 (
		_w1007_,
		_w1010_,
		_w2651_,
		_w2652_,
		_w2653_
	);
	LUT2 #(
		.INIT('h8)
	) name2191 (
		_w871_,
		_w895_,
		_w2654_
	);
	LUT3 #(
		.INIT('h15)
	) name2192 (
		_w866_,
		_w871_,
		_w921_,
		_w2655_
	);
	LUT2 #(
		.INIT('h8)
	) name2193 (
		_w843_,
		_w1022_,
		_w2656_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2194 (
		_w2653_,
		_w2654_,
		_w2655_,
		_w2656_,
		_w2657_
	);
	LUT4 #(
		.INIT('h0001)
	) name2195 (
		_w782_,
		_w791_,
		_w1065_,
		_w1081_,
		_w2658_
	);
	LUT4 #(
		.INIT('h0001)
	) name2196 (
		_w726_,
		_w741_,
		_w802_,
		_w818_,
		_w2659_
	);
	LUT2 #(
		.INIT('h8)
	) name2197 (
		_w2658_,
		_w2659_,
		_w2660_
	);
	LUT3 #(
		.INIT('h13)
	) name2198 (
		_w771_,
		_w813_,
		_w819_,
		_w2661_
	);
	LUT4 #(
		.INIT('hec00)
	) name2199 (
		_w771_,
		_w813_,
		_w819_,
		_w2658_,
		_w2662_
	);
	LUT3 #(
		.INIT('h70)
	) name2200 (
		_w816_,
		_w1082_,
		_w1088_,
		_w2663_
	);
	LUT2 #(
		.INIT('h4)
	) name2201 (
		_w2662_,
		_w2663_,
		_w2664_
	);
	LUT4 #(
		.INIT('h2f00)
	) name2202 (
		_w2650_,
		_w2657_,
		_w2660_,
		_w2664_,
		_w2665_
	);
	LUT4 #(
		.INIT('hc535)
	) name2203 (
		\P1_reg2_reg[26]/NET0131 ,
		_w1224_,
		_w2189_,
		_w2665_,
		_w2666_
	);
	LUT2 #(
		.INIT('h2)
	) name2204 (
		_w488_,
		_w1063_,
		_w2667_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name2205 (
		_w1035_,
		_w1047_,
		_w2144_,
		_w2213_,
		_w2668_
	);
	LUT3 #(
		.INIT('h15)
	) name2206 (
		_w488_,
		_w2146_,
		_w2213_,
		_w2669_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2207 (
		_w2189_,
		_w2667_,
		_w2668_,
		_w2669_,
		_w2670_
	);
	LUT3 #(
		.INIT('ha8)
	) name2208 (
		_w1237_,
		_w2649_,
		_w2670_,
		_w2671_
	);
	LUT4 #(
		.INIT('h0001)
	) name2209 (
		_w1219_,
		_w1199_,
		_w1208_,
		_w1211_,
		_w2672_
	);
	LUT3 #(
		.INIT('hb0)
	) name2210 (
		_w2100_,
		_w2107_,
		_w2110_,
		_w2673_
	);
	LUT4 #(
		.INIT('h0001)
	) name2211 (
		_w1227_,
		_w1202_,
		_w1215_,
		_w2087_,
		_w2674_
	);
	LUT2 #(
		.INIT('h8)
	) name2212 (
		_w2086_,
		_w2089_,
		_w2675_
	);
	LUT3 #(
		.INIT('h07)
	) name2213 (
		_w2064_,
		_w2090_,
		_w2094_,
		_w2676_
	);
	LUT3 #(
		.INIT('hd0)
	) name2214 (
		_w2086_,
		_w2095_,
		_w2097_,
		_w2677_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2215 (
		_w2674_,
		_w2675_,
		_w2676_,
		_w2677_,
		_w2678_
	);
	LUT3 #(
		.INIT('ha2)
	) name2216 (
		_w2672_,
		_w2673_,
		_w2678_,
		_w2679_
	);
	LUT4 #(
		.INIT('h0001)
	) name2217 (
		_w1182_,
		_w1171_,
		_w2066_,
		_w2083_,
		_w2680_
	);
	LUT3 #(
		.INIT('h8a)
	) name2218 (
		_w2061_,
		_w2081_,
		_w2084_,
		_w2681_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2219 (
		_w2077_,
		_w2079_,
		_w2680_,
		_w2681_,
		_w2682_
	);
	LUT2 #(
		.INIT('h8)
	) name2220 (
		_w2059_,
		_w2090_,
		_w2683_
	);
	LUT3 #(
		.INIT('h80)
	) name2221 (
		_w2672_,
		_w2674_,
		_w2675_,
		_w2684_
	);
	LUT3 #(
		.INIT('hc4)
	) name2222 (
		_w2104_,
		_w2113_,
		_w2111_,
		_w2685_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2223 (
		_w2682_,
		_w2683_,
		_w2684_,
		_w2685_,
		_w2686_
	);
	LUT4 #(
		.INIT('h4844)
	) name2224 (
		_w1224_,
		_w2189_,
		_w2679_,
		_w2686_,
		_w2687_
	);
	LUT4 #(
		.INIT('h4000)
	) name2225 (
		_w1059_,
		_w2155_,
		_w2163_,
		_w2164_,
		_w2688_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2226 (
		\P1_reg2_reg[26]/NET0131 ,
		_w1031_,
		_w2189_,
		_w2688_,
		_w2689_
	);
	LUT3 #(
		.INIT('h10)
	) name2227 (
		_w489_,
		_w1030_,
		_w2194_,
		_w2690_
	);
	LUT4 #(
		.INIT('h1000)
	) name2228 (
		_w489_,
		_w1030_,
		_w2189_,
		_w2194_,
		_w2691_
	);
	LUT2 #(
		.INIT('h8)
	) name2229 (
		_w1032_,
		_w1120_,
		_w2692_
	);
	LUT4 #(
		.INIT('h0057)
	) name2230 (
		\P1_reg2_reg[26]/NET0131 ,
		_w2171_,
		_w2196_,
		_w2692_,
		_w2693_
	);
	LUT2 #(
		.INIT('h4)
	) name2231 (
		_w2691_,
		_w2693_,
		_w2694_
	);
	LUT3 #(
		.INIT('hd0)
	) name2232 (
		_w2170_,
		_w2689_,
		_w2694_,
		_w2695_
	);
	LUT4 #(
		.INIT('h5700)
	) name2233 (
		_w2121_,
		_w2649_,
		_w2687_,
		_w2695_,
		_w2696_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2234 (
		_w2128_,
		_w2666_,
		_w2671_,
		_w2696_,
		_w2697_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2235 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w2648_,
		_w2697_,
		_w2698_
	);
	LUT2 #(
		.INIT('he)
	) name2236 (
		_w2647_,
		_w2698_,
		_w2699_
	);
	LUT2 #(
		.INIT('h8)
	) name2237 (
		_w1060_,
		_w2183_,
		_w2700_
	);
	LUT4 #(
		.INIT('h2220)
	) name2238 (
		_w1060_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w2701_
	);
	LUT4 #(
		.INIT('h8000)
	) name2239 (
		_w2267_,
		_w2268_,
		_w2286_,
		_w2287_,
		_w2702_
	);
	LUT4 #(
		.INIT('h8f00)
	) name2240 (
		_w2272_,
		_w2275_,
		_w2279_,
		_w2702_,
		_w2703_
	);
	LUT3 #(
		.INIT('hb0)
	) name2241 (
		_w2282_,
		_w2288_,
		_w2292_,
		_w2704_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2242 (
		_w2285_,
		_w2296_,
		_w2703_,
		_w2704_,
		_w2705_
	);
	LUT4 #(
		.INIT('h5a9a)
	) name2243 (
		_w1221_,
		_w2302_,
		_w2307_,
		_w2705_,
		_w2706_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2244 (
		_w1060_,
		_w2055_,
		_w2121_,
		_w2706_,
		_w2707_
	);
	LUT4 #(
		.INIT('h1444)
	) name2245 (
		_w488_,
		_w1035_,
		_w2144_,
		_w2213_,
		_w2708_
	);
	LUT3 #(
		.INIT('h20)
	) name2246 (
		_w488_,
		_w1075_,
		_w1078_,
		_w2709_
	);
	LUT4 #(
		.INIT('h3331)
	) name2247 (
		_w2055_,
		_w2701_,
		_w2708_,
		_w2709_,
		_w2710_
	);
	LUT2 #(
		.INIT('h2)
	) name2248 (
		_w1237_,
		_w2710_,
		_w2711_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2249 (
		_w2220_,
		_w2223_,
		_w2228_,
		_w2246_,
		_w2712_
	);
	LUT3 #(
		.INIT('hc4)
	) name2250 (
		_w2250_,
		_w2253_,
		_w2712_,
		_w2713_
	);
	LUT3 #(
		.INIT('h80)
	) name2251 (
		_w2220_,
		_w2223_,
		_w2253_,
		_w2714_
	);
	LUT3 #(
		.INIT('h4c)
	) name2252 (
		_w2242_,
		_w2261_,
		_w2714_,
		_w2715_
	);
	LUT4 #(
		.INIT('h8488)
	) name2253 (
		_w1221_,
		_w2055_,
		_w2713_,
		_w2715_,
		_w2716_
	);
	LUT4 #(
		.INIT('h9555)
	) name2254 (
		_w1059_,
		_w2155_,
		_w2163_,
		_w2164_,
		_w2717_
	);
	LUT4 #(
		.INIT('h5400)
	) name2255 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2170_,
		_w2718_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2256 (
		_w1060_,
		_w2171_,
		_w2578_,
		_w2718_,
		_w2719_
	);
	LUT4 #(
		.INIT('h0100)
	) name2257 (
		_w489_,
		_w1058_,
		_w2175_,
		_w2176_,
		_w2720_
	);
	LUT2 #(
		.INIT('h1)
	) name2258 (
		_w2719_,
		_w2720_,
		_w2721_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2259 (
		_w2055_,
		_w2170_,
		_w2717_,
		_w2721_,
		_w2722_
	);
	LUT4 #(
		.INIT('h5700)
	) name2260 (
		_w2128_,
		_w2701_,
		_w2716_,
		_w2722_,
		_w2723_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2261 (
		_w2182_,
		_w2707_,
		_w2711_,
		_w2723_,
		_w2724_
	);
	LUT2 #(
		.INIT('h2)
	) name2262 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2725_
	);
	LUT4 #(
		.INIT('h6a00)
	) name2263 (
		\P1_reg3_reg[25]/NET0131 ,
		_w593_,
		_w596_,
		_w1244_,
		_w2726_
	);
	LUT2 #(
		.INIT('h1)
	) name2264 (
		_w2725_,
		_w2726_,
		_w2727_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2265 (
		\P1_state_reg[0]/NET0131 ,
		_w2700_,
		_w2724_,
		_w2727_,
		_w2728_
	);
	LUT4 #(
		.INIT('h1000)
	) name2266 (
		_w1290_,
		_w1288_,
		_w1291_,
		_w1295_,
		_w2729_
	);
	LUT4 #(
		.INIT('hc355)
	) name2267 (
		\P2_reg0_reg[29]/NET0131 ,
		_w1404_,
		_w1857_,
		_w2729_,
		_w2730_
	);
	LUT2 #(
		.INIT('h2)
	) name2268 (
		_w1869_,
		_w2730_,
		_w2731_
	);
	LUT4 #(
		.INIT('h3c55)
	) name2269 (
		\P2_reg0_reg[29]/NET0131 ,
		_w1404_,
		_w1961_,
		_w2729_,
		_w2732_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2270 (
		_w1998_,
		_w2000_,
		_w2026_,
		_w2729_,
		_w2733_
	);
	LUT4 #(
		.INIT('h1ffd)
	) name2271 (
		_w1595_,
		_w1859_,
		_w1863_,
		_w1866_,
		_w2734_
	);
	LUT3 #(
		.INIT('hd0)
	) name2272 (
		_w2033_,
		_w2729_,
		_w2734_,
		_w2735_
	);
	LUT2 #(
		.INIT('h2)
	) name2273 (
		_w2000_,
		_w2729_,
		_w2736_
	);
	LUT4 #(
		.INIT('hf100)
	) name2274 (
		_w2000_,
		_w2033_,
		_w2729_,
		_w2734_,
		_w2737_
	);
	LUT2 #(
		.INIT('h2)
	) name2275 (
		\P2_reg0_reg[29]/NET0131 ,
		_w2737_,
		_w2738_
	);
	LUT4 #(
		.INIT('h000d)
	) name2276 (
		_w1963_,
		_w2732_,
		_w2733_,
		_w2738_,
		_w2739_
	);
	LUT4 #(
		.INIT('h2000)
	) name2277 (
		\P2_reg0_reg[29]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w2740_
	);
	LUT4 #(
		.INIT('h0075)
	) name2278 (
		_w1285_,
		_w2731_,
		_w2739_,
		_w2740_,
		_w2741_
	);
	LUT2 #(
		.INIT('h2)
	) name2279 (
		\P2_reg0_reg[29]/NET0131 ,
		_w2042_,
		_w2742_
	);
	LUT3 #(
		.INIT('hf2)
	) name2280 (
		\P1_state_reg[0]/NET0131 ,
		_w2741_,
		_w2742_,
		_w2743_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2281 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[24]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w2744_
	);
	LUT2 #(
		.INIT('h8)
	) name2282 (
		\P1_reg2_reg[24]/NET0131 ,
		_w2183_,
		_w2745_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2283 (
		\P1_reg2_reg[24]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w2746_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2284 (
		\P1_reg2_reg[24]/NET0131 ,
		_w1210_,
		_w2189_,
		_w2565_,
		_w2747_
	);
	LUT4 #(
		.INIT('h7020)
	) name2285 (
		_w488_,
		_w789_,
		_w2189_,
		_w2567_,
		_w2748_
	);
	LUT3 #(
		.INIT('ha8)
	) name2286 (
		_w1237_,
		_w2746_,
		_w2748_,
		_w2749_
	);
	LUT4 #(
		.INIT('h8488)
	) name2287 (
		_w1210_,
		_w2189_,
		_w2571_,
		_w2572_,
		_w2750_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2288 (
		\P1_reg2_reg[24]/NET0131 ,
		_w2189_,
		_w2574_,
		_w2575_,
		_w2751_
	);
	LUT4 #(
		.INIT('h5400)
	) name2289 (
		_w489_,
		_w1066_,
		_w1072_,
		_w2194_,
		_w2752_
	);
	LUT2 #(
		.INIT('h8)
	) name2290 (
		_w2189_,
		_w2752_,
		_w2753_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2291 (
		\P1_reg3_reg[24]/NET0131 ,
		_w785_,
		_w597_,
		_w1120_,
		_w2754_
	);
	LUT4 #(
		.INIT('h0057)
	) name2292 (
		\P1_reg2_reg[24]/NET0131 ,
		_w2171_,
		_w2196_,
		_w2754_,
		_w2755_
	);
	LUT2 #(
		.INIT('h4)
	) name2293 (
		_w2753_,
		_w2755_,
		_w2756_
	);
	LUT3 #(
		.INIT('hd0)
	) name2294 (
		_w2170_,
		_w2751_,
		_w2756_,
		_w2757_
	);
	LUT4 #(
		.INIT('h5700)
	) name2295 (
		_w2128_,
		_w2746_,
		_w2750_,
		_w2757_,
		_w2758_
	);
	LUT4 #(
		.INIT('h3100)
	) name2296 (
		_w2121_,
		_w2749_,
		_w2747_,
		_w2758_,
		_w2759_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2297 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w2745_,
		_w2759_,
		_w2760_
	);
	LUT2 #(
		.INIT('he)
	) name2298 (
		_w2744_,
		_w2760_,
		_w2761_
	);
	LUT4 #(
		.INIT('h0100)
	) name2299 (
		_w1290_,
		_w1288_,
		_w1291_,
		_w1295_,
		_w2762_
	);
	LUT4 #(
		.INIT('hc355)
	) name2300 (
		\P2_reg1_reg[29]/NET0131 ,
		_w1404_,
		_w1857_,
		_w2762_,
		_w2763_
	);
	LUT2 #(
		.INIT('h2)
	) name2301 (
		_w1869_,
		_w2763_,
		_w2764_
	);
	LUT4 #(
		.INIT('h3c55)
	) name2302 (
		\P2_reg1_reg[29]/NET0131 ,
		_w1404_,
		_w1961_,
		_w2762_,
		_w2765_
	);
	LUT4 #(
		.INIT('h30a0)
	) name2303 (
		\P2_reg1_reg[29]/NET0131 ,
		_w1998_,
		_w2000_,
		_w2762_,
		_w2766_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name2304 (
		\P2_reg1_reg[29]/NET0131 ,
		_w2023_,
		_w2025_,
		_w2762_,
		_w2767_
	);
	LUT2 #(
		.INIT('h2)
	) name2305 (
		\P2_reg1_reg[29]/NET0131 ,
		_w2734_,
		_w2768_
	);
	LUT4 #(
		.INIT('hfc55)
	) name2306 (
		\P2_reg1_reg[29]/NET0131 ,
		_w1306_,
		_w1373_,
		_w2762_,
		_w2769_
	);
	LUT3 #(
		.INIT('h31)
	) name2307 (
		_w2001_,
		_w2768_,
		_w2769_,
		_w2770_
	);
	LUT2 #(
		.INIT('h4)
	) name2308 (
		_w2767_,
		_w2770_,
		_w2771_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2309 (
		_w1963_,
		_w2765_,
		_w2766_,
		_w2771_,
		_w2772_
	);
	LUT4 #(
		.INIT('h2000)
	) name2310 (
		\P2_reg1_reg[29]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w2773_
	);
	LUT4 #(
		.INIT('h0075)
	) name2311 (
		_w1285_,
		_w2764_,
		_w2772_,
		_w2773_,
		_w2774_
	);
	LUT2 #(
		.INIT('h2)
	) name2312 (
		\P2_reg1_reg[29]/NET0131 ,
		_w2042_,
		_w2775_
	);
	LUT3 #(
		.INIT('hf2)
	) name2313 (
		\P1_state_reg[0]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2776_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2314 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[28]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w2777_
	);
	LUT4 #(
		.INIT('h3c55)
	) name2315 (
		\P1_reg0_reg[28]/NET0131 ,
		_w1160_,
		_w2117_,
		_w2325_,
		_w2778_
	);
	LUT4 #(
		.INIT('h30a0)
	) name2316 (
		\P1_reg0_reg[28]/NET0131 ,
		_w2127_,
		_w2128_,
		_w2325_,
		_w2779_
	);
	LUT3 #(
		.INIT('h07)
	) name2317 (
		_w2169_,
		_w2170_,
		_w2195_,
		_w2780_
	);
	LUT4 #(
		.INIT('h5700)
	) name2318 (
		_w1237_,
		_w2150_,
		_w2151_,
		_w2780_,
		_w2781_
	);
	LUT3 #(
		.INIT('h90)
	) name2319 (
		_w1096_,
		_w1098_,
		_w1122_,
		_w2782_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2320 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2782_,
		_w2783_
	);
	LUT3 #(
		.INIT('h02)
	) name2321 (
		_w2332_,
		_w2333_,
		_w2783_,
		_w2784_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2322 (
		\P1_reg0_reg[28]/NET0131 ,
		_w2332_,
		_w2333_,
		_w2783_,
		_w2785_
	);
	LUT3 #(
		.INIT('h0d)
	) name2323 (
		_w2325_,
		_w2781_,
		_w2785_,
		_w2786_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2324 (
		_w2121_,
		_w2778_,
		_w2779_,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('h8)
	) name2325 (
		\P1_reg0_reg[28]/NET0131 ,
		_w2183_,
		_w2788_
	);
	LUT4 #(
		.INIT('haa08)
	) name2326 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w2787_,
		_w2788_,
		_w2789_
	);
	LUT2 #(
		.INIT('he)
	) name2327 (
		_w2777_,
		_w2789_,
		_w2790_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2328 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[25]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w2791_
	);
	LUT2 #(
		.INIT('h8)
	) name2329 (
		\P1_reg0_reg[25]/NET0131 ,
		_w2183_,
		_w2792_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2330 (
		\P1_reg0_reg[25]/NET0131 ,
		_w2121_,
		_w2325_,
		_w2706_,
		_w2793_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2331 (
		\P1_reg0_reg[25]/NET0131 ,
		_w2325_,
		_w2708_,
		_w2709_,
		_w2794_
	);
	LUT2 #(
		.INIT('h2)
	) name2332 (
		_w1237_,
		_w2794_,
		_w2795_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2333 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2170_,
		_w2796_
	);
	LUT3 #(
		.INIT('h02)
	) name2334 (
		_w2332_,
		_w2333_,
		_w2796_,
		_w2797_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2335 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2128_,
		_w2798_
	);
	LUT4 #(
		.INIT('h0002)
	) name2336 (
		_w2332_,
		_w2333_,
		_w2796_,
		_w2798_,
		_w2799_
	);
	LUT2 #(
		.INIT('h2)
	) name2337 (
		\P1_reg0_reg[25]/NET0131 ,
		_w2799_,
		_w2800_
	);
	LUT4 #(
		.INIT('h8488)
	) name2338 (
		_w1221_,
		_w2128_,
		_w2713_,
		_w2715_,
		_w2801_
	);
	LUT3 #(
		.INIT('h10)
	) name2339 (
		_w489_,
		_w1058_,
		_w2194_,
		_w2802_
	);
	LUT3 #(
		.INIT('h07)
	) name2340 (
		_w2170_,
		_w2717_,
		_w2802_,
		_w2803_
	);
	LUT4 #(
		.INIT('h1311)
	) name2341 (
		_w2325_,
		_w2800_,
		_w2801_,
		_w2803_,
		_w2804_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2342 (
		_w2182_,
		_w2793_,
		_w2795_,
		_w2804_,
		_w2805_
	);
	LUT4 #(
		.INIT('heeec)
	) name2343 (
		\P1_state_reg[0]/NET0131 ,
		_w2791_,
		_w2792_,
		_w2805_,
		_w2806_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2344 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[26]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w2807_
	);
	LUT2 #(
		.INIT('h8)
	) name2345 (
		\P1_reg1_reg[26]/NET0131 ,
		_w2183_,
		_w2808_
	);
	LUT4 #(
		.INIT('h5455)
	) name2346 (
		\P1_reg1_reg[26]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w2809_
	);
	LUT2 #(
		.INIT('h2)
	) name2347 (
		_w2128_,
		_w2809_,
		_w2810_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2348 (
		_w1224_,
		_w2536_,
		_w2665_,
		_w2810_,
		_w2811_
	);
	LUT4 #(
		.INIT('h4844)
	) name2349 (
		_w1224_,
		_w2121_,
		_w2679_,
		_w2686_,
		_w2812_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2350 (
		_w1237_,
		_w2667_,
		_w2668_,
		_w2669_,
		_w2813_
	);
	LUT4 #(
		.INIT('h007b)
	) name2351 (
		_w1031_,
		_w2170_,
		_w2688_,
		_w2690_,
		_w2814_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2352 (
		_w2536_,
		_w2813_,
		_w2812_,
		_w2814_,
		_w2815_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2353 (
		_w1237_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w2816_
	);
	LUT4 #(
		.INIT('hef00)
	) name2354 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2170_,
		_w2817_
	);
	LUT4 #(
		.INIT('h0002)
	) name2355 (
		_w2332_,
		_w2544_,
		_w2816_,
		_w2817_,
		_w2818_
	);
	LUT4 #(
		.INIT('h7202)
	) name2356 (
		_w1096_,
		_w1100_,
		_w1098_,
		_w718_,
		_w2819_
	);
	LUT4 #(
		.INIT('hef00)
	) name2357 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2819_,
		_w2820_
	);
	LUT2 #(
		.INIT('h4)
	) name2358 (
		_w1236_,
		_w2820_,
		_w2821_
	);
	LUT3 #(
		.INIT('ha2)
	) name2359 (
		\P1_reg1_reg[26]/NET0131 ,
		_w2818_,
		_w2821_,
		_w2822_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2360 (
		_w2182_,
		_w2815_,
		_w2822_,
		_w2811_,
		_w2823_
	);
	LUT4 #(
		.INIT('heeec)
	) name2361 (
		\P1_state_reg[0]/NET0131 ,
		_w2807_,
		_w2808_,
		_w2823_,
		_w2824_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2362 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[28]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w2825_
	);
	LUT4 #(
		.INIT('h3c55)
	) name2363 (
		\P1_reg1_reg[28]/NET0131 ,
		_w1160_,
		_w2117_,
		_w2536_,
		_w2826_
	);
	LUT4 #(
		.INIT('h30a0)
	) name2364 (
		\P1_reg1_reg[28]/NET0131 ,
		_w2127_,
		_w2128_,
		_w2536_,
		_w2827_
	);
	LUT2 #(
		.INIT('h2)
	) name2365 (
		\P1_reg1_reg[28]/NET0131 ,
		_w2818_,
		_w2828_
	);
	LUT3 #(
		.INIT('h0d)
	) name2366 (
		_w2536_,
		_w2781_,
		_w2828_,
		_w2829_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2367 (
		_w2121_,
		_w2826_,
		_w2827_,
		_w2829_,
		_w2830_
	);
	LUT2 #(
		.INIT('h8)
	) name2368 (
		\P1_reg1_reg[28]/NET0131 ,
		_w2183_,
		_w2831_
	);
	LUT4 #(
		.INIT('haa08)
	) name2369 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w2830_,
		_w2831_,
		_w2832_
	);
	LUT2 #(
		.INIT('he)
	) name2370 (
		_w2825_,
		_w2832_,
		_w2833_
	);
	LUT2 #(
		.INIT('h8)
	) name2371 (
		_w760_,
		_w2183_,
		_w2834_
	);
	LUT4 #(
		.INIT('h2220)
	) name2372 (
		_w760_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w2835_
	);
	LUT4 #(
		.INIT('h7500)
	) name2373 (
		_w2065_,
		_w2082_,
		_w2085_,
		_w2091_,
		_w2836_
	);
	LUT4 #(
		.INIT('h8848)
	) name2374 (
		_w1198_,
		_w2055_,
		_w2096_,
		_w2836_,
		_w2837_
	);
	LUT3 #(
		.INIT('ha8)
	) name2375 (
		_w2121_,
		_w2835_,
		_w2837_,
		_w2838_
	);
	LUT3 #(
		.INIT('h80)
	) name2376 (
		_w488_,
		_w824_,
		_w826_,
		_w2839_
	);
	LUT4 #(
		.INIT('h00eb)
	) name2377 (
		_w488_,
		_w754_,
		_w2139_,
		_w2839_,
		_w2840_
	);
	LUT4 #(
		.INIT('hc808)
	) name2378 (
		_w760_,
		_w1237_,
		_w2055_,
		_w2840_,
		_w2841_
	);
	LUT3 #(
		.INIT('h60)
	) name2379 (
		_w759_,
		_w2163_,
		_w2170_,
		_w2842_
	);
	LUT4 #(
		.INIT('h006f)
	) name2380 (
		_w1020_,
		_w1198_,
		_w2128_,
		_w2842_,
		_w2843_
	);
	LUT3 #(
		.INIT('h10)
	) name2381 (
		_w759_,
		_w2175_,
		_w2176_,
		_w2844_
	);
	LUT4 #(
		.INIT('h5400)
	) name2382 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2128_,
		_w2845_
	);
	LUT4 #(
		.INIT('h0001)
	) name2383 (
		_w2171_,
		_w2578_,
		_w2718_,
		_w2845_,
		_w2846_
	);
	LUT3 #(
		.INIT('h31)
	) name2384 (
		_w760_,
		_w2844_,
		_w2846_,
		_w2847_
	);
	LUT4 #(
		.INIT('h3100)
	) name2385 (
		_w2055_,
		_w2841_,
		_w2843_,
		_w2847_,
		_w2848_
	);
	LUT4 #(
		.INIT('h1311)
	) name2386 (
		_w2182_,
		_w2834_,
		_w2838_,
		_w2848_,
		_w2849_
	);
	LUT2 #(
		.INIT('h2)
	) name2387 (
		\P1_reg3_reg[16]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2850_
	);
	LUT3 #(
		.INIT('h07)
	) name2388 (
		_w760_,
		_w1244_,
		_w2850_,
		_w2851_
	);
	LUT3 #(
		.INIT('h2f)
	) name2389 (
		\P1_state_reg[0]/NET0131 ,
		_w2849_,
		_w2851_,
		_w2852_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2390 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w2853_
	);
	LUT2 #(
		.INIT('h8)
	) name2391 (
		\P1_reg2_reg[31]/NET0131 ,
		_w2183_,
		_w2854_
	);
	LUT3 #(
		.INIT('h40)
	) name2392 (
		_w489_,
		_w569_,
		_w2194_,
		_w2855_
	);
	LUT2 #(
		.INIT('h4)
	) name2393 (
		_w602_,
		_w1237_,
		_w2856_
	);
	LUT4 #(
		.INIT('hb000)
	) name2394 (
		_w650_,
		_w2214_,
		_w2216_,
		_w2856_,
		_w2857_
	);
	LUT2 #(
		.INIT('h8)
	) name2395 (
		_w864_,
		_w2161_,
		_w2858_
	);
	LUT4 #(
		.INIT('h8000)
	) name2396 (
		_w852_,
		_w2159_,
		_w2160_,
		_w2858_,
		_w2859_
	);
	LUT4 #(
		.INIT('h8000)
	) name2397 (
		_w833_,
		_w842_,
		_w2155_,
		_w2859_,
		_w2860_
	);
	LUT3 #(
		.INIT('hea)
	) name2398 (
		_w489_,
		_w673_,
		_w646_,
		_w2861_
	);
	LUT2 #(
		.INIT('h4)
	) name2399 (
		_w702_,
		_w2861_,
		_w2862_
	);
	LUT4 #(
		.INIT('h9555)
	) name2400 (
		_w570_,
		_w2167_,
		_w2860_,
		_w2862_,
		_w2863_
	);
	LUT4 #(
		.INIT('h5545)
	) name2401 (
		\P1_reg2_reg[31]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w2864_
	);
	LUT2 #(
		.INIT('h2)
	) name2402 (
		_w2170_,
		_w2864_,
		_w2865_
	);
	LUT4 #(
		.INIT('h5545)
	) name2403 (
		_w1119_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w2866_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2404 (
		\P1_reg2_reg[31]/NET0131 ,
		_w2171_,
		_w2196_,
		_w2866_,
		_w2867_
	);
	LUT2 #(
		.INIT('h1)
	) name2405 (
		_w2316_,
		_w2867_,
		_w2868_
	);
	LUT4 #(
		.INIT('h2f00)
	) name2406 (
		_w2189_,
		_w2863_,
		_w2865_,
		_w2868_,
		_w2869_
	);
	LUT4 #(
		.INIT('h5700)
	) name2407 (
		_w2189_,
		_w2855_,
		_w2857_,
		_w2869_,
		_w2870_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2408 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w2854_,
		_w2870_,
		_w2871_
	);
	LUT2 #(
		.INIT('he)
	) name2409 (
		_w2853_,
		_w2871_,
		_w2872_
	);
	LUT2 #(
		.INIT('h2)
	) name2410 (
		\P2_reg2_reg[25]/NET0131 ,
		_w2042_,
		_w2873_
	);
	LUT4 #(
		.INIT('h2000)
	) name2411 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w2874_
	);
	LUT3 #(
		.INIT('h40)
	) name2412 (
		_w1905_,
		_w1908_,
		_w1917_,
		_w2875_
	);
	LUT4 #(
		.INIT('h40cc)
	) name2413 (
		_w1878_,
		_w1913_,
		_w1916_,
		_w1923_,
		_w2876_
	);
	LUT2 #(
		.INIT('h2)
	) name2414 (
		_w1931_,
		_w2876_,
		_w2877_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2415 (
		_w1945_,
		_w1952_,
		_w2875_,
		_w2877_,
		_w2878_
	);
	LUT4 #(
		.INIT('hd11d)
	) name2416 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1298_,
		_w2519_,
		_w2878_,
		_w2879_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2417 (
		_w1792_,
		_w1797_,
		_w1841_,
		_w1845_,
		_w2880_
	);
	LUT3 #(
		.INIT('h80)
	) name2418 (
		_w1554_,
		_w1635_,
		_w1854_,
		_w2881_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2419 (
		_w1554_,
		_w1848_,
		_w1851_,
		_w1854_,
		_w2882_
	);
	LUT2 #(
		.INIT('h2)
	) name2420 (
		_w1579_,
		_w2882_,
		_w2883_
	);
	LUT4 #(
		.INIT('h65aa)
	) name2421 (
		_w2519_,
		_w2880_,
		_w2881_,
		_w2883_,
		_w2884_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2422 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1298_,
		_w1869_,
		_w2884_,
		_w2885_
	);
	LUT4 #(
		.INIT('h1444)
	) name2423 (
		_w1305_,
		_w1510_,
		_w1978_,
		_w1987_,
		_w2886_
	);
	LUT3 #(
		.INIT('h20)
	) name2424 (
		_w1305_,
		_w1538_,
		_w1541_,
		_w2887_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2425 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1298_,
		_w2886_,
		_w2887_,
		_w2888_
	);
	LUT4 #(
		.INIT('h5400)
	) name2426 (
		_w1306_,
		_w1514_,
		_w1521_,
		_w2001_,
		_w2889_
	);
	LUT4 #(
		.INIT('h8000)
	) name2427 (
		_w2009_,
		_w2010_,
		_w2015_,
		_w2017_,
		_w2890_
	);
	LUT3 #(
		.INIT('h8a)
	) name2428 (
		_w1522_,
		_w1534_,
		_w2890_,
		_w2891_
	);
	LUT2 #(
		.INIT('h2)
	) name2429 (
		_w2025_,
		_w2632_,
		_w2892_
	);
	LUT3 #(
		.INIT('h45)
	) name2430 (
		_w2889_,
		_w2891_,
		_w2892_,
		_w2893_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2431 (
		_w1298_,
		_w2889_,
		_w2891_,
		_w2892_,
		_w2894_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name2432 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1298_,
		_w2032_,
		_w2033_,
		_w2895_
	);
	LUT2 #(
		.INIT('h8)
	) name2433 (
		_w1523_,
		_w2029_,
		_w2896_
	);
	LUT2 #(
		.INIT('h1)
	) name2434 (
		_w2895_,
		_w2896_,
		_w2897_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2435 (
		_w2000_,
		_w2888_,
		_w2894_,
		_w2897_,
		_w2898_
	);
	LUT4 #(
		.INIT('h3100)
	) name2436 (
		_w1963_,
		_w2885_,
		_w2879_,
		_w2898_,
		_w2899_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2437 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w2874_,
		_w2899_,
		_w2900_
	);
	LUT2 #(
		.INIT('he)
	) name2438 (
		_w2873_,
		_w2900_,
		_w2901_
	);
	LUT2 #(
		.INIT('h8)
	) name2439 (
		_w1523_,
		_w2039_,
		_w2902_
	);
	LUT4 #(
		.INIT('heeef)
	) name2440 (
		_w1290_,
		_w1288_,
		_w1291_,
		_w1295_,
		_w2903_
	);
	LUT2 #(
		.INIT('h2)
	) name2441 (
		_w1523_,
		_w2903_,
		_w2904_
	);
	LUT4 #(
		.INIT('h009f)
	) name2442 (
		_w2519_,
		_w2878_,
		_w2903_,
		_w2904_,
		_w2905_
	);
	LUT4 #(
		.INIT('h0c88)
	) name2443 (
		_w1523_,
		_w1869_,
		_w2884_,
		_w2903_,
		_w2906_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2444 (
		_w2886_,
		_w2887_,
		_w2903_,
		_w2904_,
		_w2907_
	);
	LUT4 #(
		.INIT('hba00)
	) name2445 (
		_w2889_,
		_w2891_,
		_w2892_,
		_w2903_,
		_w2908_
	);
	LUT4 #(
		.INIT('h88a8)
	) name2446 (
		_w1523_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w2909_
	);
	LUT4 #(
		.INIT('h5400)
	) name2447 (
		_w1306_,
		_w1514_,
		_w1521_,
		_w2029_,
		_w2910_
	);
	LUT2 #(
		.INIT('h1)
	) name2448 (
		_w2909_,
		_w2910_,
		_w2911_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2449 (
		_w2000_,
		_w2907_,
		_w2908_,
		_w2911_,
		_w2912_
	);
	LUT4 #(
		.INIT('h3100)
	) name2450 (
		_w1963_,
		_w2906_,
		_w2905_,
		_w2912_,
		_w2913_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2451 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w2902_,
		_w2913_,
		_w2914_
	);
	LUT4 #(
		.INIT('h9b3b)
	) name2452 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[25]/NET0131 ,
		_w1267_,
		_w1394_,
		_w2915_
	);
	LUT2 #(
		.INIT('hb)
	) name2453 (
		_w2914_,
		_w2915_,
		_w2916_
	);
	LUT2 #(
		.INIT('h8)
	) name2454 (
		_w1032_,
		_w2183_,
		_w2917_
	);
	LUT4 #(
		.INIT('h2220)
	) name2455 (
		_w1032_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w2918_
	);
	LUT4 #(
		.INIT('h00b7)
	) name2456 (
		_w1224_,
		_w2055_,
		_w2665_,
		_w2918_,
		_w2919_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2457 (
		_w2055_,
		_w2667_,
		_w2668_,
		_w2669_,
		_w2920_
	);
	LUT3 #(
		.INIT('ha8)
	) name2458 (
		_w1237_,
		_w2918_,
		_w2920_,
		_w2921_
	);
	LUT4 #(
		.INIT('h4844)
	) name2459 (
		_w1224_,
		_w2055_,
		_w2679_,
		_w2686_,
		_w2922_
	);
	LUT4 #(
		.INIT('h8040)
	) name2460 (
		_w1031_,
		_w2055_,
		_w2170_,
		_w2688_,
		_w2923_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2461 (
		_w1032_,
		_w2171_,
		_w2578_,
		_w2718_,
		_w2924_
	);
	LUT4 #(
		.INIT('h0100)
	) name2462 (
		_w489_,
		_w1030_,
		_w2175_,
		_w2176_,
		_w2925_
	);
	LUT2 #(
		.INIT('h1)
	) name2463 (
		_w2924_,
		_w2925_,
		_w2926_
	);
	LUT2 #(
		.INIT('h4)
	) name2464 (
		_w2923_,
		_w2926_,
		_w2927_
	);
	LUT4 #(
		.INIT('h5700)
	) name2465 (
		_w2121_,
		_w2918_,
		_w2922_,
		_w2927_,
		_w2928_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2466 (
		_w2128_,
		_w2919_,
		_w2921_,
		_w2928_,
		_w2929_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2467 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w2917_,
		_w2929_,
		_w2930_
	);
	LUT2 #(
		.INIT('h2)
	) name2468 (
		\P1_reg3_reg[26]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2931_
	);
	LUT3 #(
		.INIT('h07)
	) name2469 (
		_w1032_,
		_w1244_,
		_w2931_,
		_w2932_
	);
	LUT2 #(
		.INIT('hb)
	) name2470 (
		_w2930_,
		_w2932_,
		_w2933_
	);
	LUT2 #(
		.INIT('h2)
	) name2471 (
		_w1042_,
		_w2055_,
		_w2934_
	);
	LUT4 #(
		.INIT('hf400)
	) name2472 (
		_w2229_,
		_w2230_,
		_w2231_,
		_w2234_,
		_w2935_
	);
	LUT4 #(
		.INIT('h0001)
	) name2473 (
		_w894_,
		_w906_,
		_w944_,
		_w1016_,
		_w2936_
	);
	LUT3 #(
		.INIT('h15)
	) name2474 (
		_w2226_,
		_w2238_,
		_w2240_,
		_w2937_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2475 (
		_w2237_,
		_w2935_,
		_w2936_,
		_w2937_,
		_w2938_
	);
	LUT2 #(
		.INIT('h8)
	) name2476 (
		_w2221_,
		_w2225_,
		_w2939_
	);
	LUT3 #(
		.INIT('h0d)
	) name2477 (
		_w2221_,
		_w2227_,
		_w2244_,
		_w2940_
	);
	LUT2 #(
		.INIT('h8)
	) name2478 (
		_w2219_,
		_w2222_,
		_w2941_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2479 (
		_w2938_,
		_w2939_,
		_w2940_,
		_w2941_,
		_w2942_
	);
	LUT3 #(
		.INIT('h07)
	) name2480 (
		_w2219_,
		_w2245_,
		_w2247_,
		_w2943_
	);
	LUT4 #(
		.INIT('h0001)
	) name2481 (
		_w791_,
		_w1037_,
		_w1065_,
		_w1081_,
		_w2944_
	);
	LUT3 #(
		.INIT('h10)
	) name2482 (
		_w726_,
		_w818_,
		_w2252_,
		_w2945_
	);
	LUT2 #(
		.INIT('h8)
	) name2483 (
		_w2944_,
		_w2945_,
		_w2946_
	);
	LUT4 #(
		.INIT('h2b00)
	) name2484 (
		_w770_,
		_w805_,
		_w810_,
		_w2252_,
		_w2947_
	);
	LUT2 #(
		.INIT('h1)
	) name2485 (
		_w2258_,
		_w2947_,
		_w2948_
	);
	LUT3 #(
		.INIT('hc8)
	) name2486 (
		_w2258_,
		_w2944_,
		_w2947_,
		_w2949_
	);
	LUT3 #(
		.INIT('h07)
	) name2487 (
		_w2254_,
		_w2260_,
		_w2262_,
		_w2950_
	);
	LUT2 #(
		.INIT('h4)
	) name2488 (
		_w2949_,
		_w2950_,
		_w2951_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2489 (
		_w2942_,
		_w2943_,
		_w2946_,
		_w2951_,
		_w2952_
	);
	LUT4 #(
		.INIT('h0b07)
	) name2490 (
		_w1165_,
		_w2055_,
		_w2934_,
		_w2952_,
		_w2953_
	);
	LUT4 #(
		.INIT('h1444)
	) name2491 (
		_w488_,
		_w708_,
		_w2146_,
		_w2213_,
		_w2954_
	);
	LUT2 #(
		.INIT('h8)
	) name2492 (
		_w488_,
		_w1035_,
		_w2955_
	);
	LUT4 #(
		.INIT('h3331)
	) name2493 (
		_w2055_,
		_w2934_,
		_w2954_,
		_w2955_,
		_w2956_
	);
	LUT2 #(
		.INIT('h2)
	) name2494 (
		_w1237_,
		_w2956_,
		_w2957_
	);
	LUT4 #(
		.INIT('h0001)
	) name2495 (
		_w1219_,
		_w1222_,
		_w1208_,
		_w1211_,
		_w2958_
	);
	LUT3 #(
		.INIT('h10)
	) name2496 (
		_w1227_,
		_w2087_,
		_w2301_,
		_w2959_
	);
	LUT2 #(
		.INIT('h8)
	) name2497 (
		_w2958_,
		_w2959_,
		_w2960_
	);
	LUT4 #(
		.INIT('h0001)
	) name2498 (
		_w1182_,
		_w1171_,
		_w2057_,
		_w2083_,
		_w2961_
	);
	LUT4 #(
		.INIT('hf800)
	) name2499 (
		_w2272_,
		_w2274_,
		_w2277_,
		_w2961_,
		_w2962_
	);
	LUT3 #(
		.INIT('h0d)
	) name2500 (
		_w2267_,
		_w2278_,
		_w2280_,
		_w2963_
	);
	LUT2 #(
		.INIT('h8)
	) name2501 (
		_w2284_,
		_w2287_,
		_w2964_
	);
	LUT2 #(
		.INIT('h8)
	) name2502 (
		_w2268_,
		_w2286_,
		_w2965_
	);
	LUT4 #(
		.INIT('h8000)
	) name2503 (
		_w2268_,
		_w2284_,
		_w2286_,
		_w2287_,
		_w2966_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2504 (
		_w2960_,
		_w2962_,
		_w2963_,
		_w2966_,
		_w2967_
	);
	LUT4 #(
		.INIT('hb200)
	) name2505 (
		_w805_,
		_w810_,
		_w2099_,
		_w2301_,
		_w2968_
	);
	LUT3 #(
		.INIT('hc4)
	) name2506 (
		_w2304_,
		_w2958_,
		_w2968_,
		_w2969_
	);
	LUT3 #(
		.INIT('hb0)
	) name2507 (
		_w2281_,
		_w2286_,
		_w2290_,
		_w2970_
	);
	LUT3 #(
		.INIT('h70)
	) name2508 (
		_w2284_,
		_w2291_,
		_w2293_,
		_w2971_
	);
	LUT3 #(
		.INIT('hd0)
	) name2509 (
		_w2964_,
		_w2970_,
		_w2971_,
		_w2972_
	);
	LUT3 #(
		.INIT('hd0)
	) name2510 (
		_w2300_,
		_w2306_,
		_w2308_,
		_w2973_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2511 (
		_w2960_,
		_w2972_,
		_w2969_,
		_w2973_,
		_w2974_
	);
	LUT4 #(
		.INIT('h4844)
	) name2512 (
		_w1165_,
		_w2055_,
		_w2967_,
		_w2974_,
		_w2975_
	);
	LUT4 #(
		.INIT('h8444)
	) name2513 (
		_w1041_,
		_w2055_,
		_w2166_,
		_w2860_,
		_w2976_
	);
	LUT3 #(
		.INIT('ha8)
	) name2514 (
		_w1042_,
		_w2171_,
		_w2578_,
		_w2977_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2515 (
		_w489_,
		_w1040_,
		_w2177_,
		_w2977_,
		_w2978_
	);
	LUT4 #(
		.INIT('h5700)
	) name2516 (
		_w2170_,
		_w2934_,
		_w2976_,
		_w2978_,
		_w2979_
	);
	LUT4 #(
		.INIT('h5700)
	) name2517 (
		_w2121_,
		_w2934_,
		_w2975_,
		_w2979_,
		_w2980_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2518 (
		_w2128_,
		_w2953_,
		_w2957_,
		_w2980_,
		_w2981_
	);
	LUT3 #(
		.INIT('h60)
	) name2519 (
		\P1_reg3_reg[27]/NET0131 ,
		_w703_,
		_w2183_,
		_w2982_
	);
	LUT4 #(
		.INIT('haa08)
	) name2520 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w2981_,
		_w2982_,
		_w2983_
	);
	LUT4 #(
		.INIT('h95dd)
	) name2521 (
		\P1_reg3_reg[27]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w703_,
		_w1243_,
		_w2984_
	);
	LUT2 #(
		.INIT('hb)
	) name2522 (
		_w2983_,
		_w2984_,
		_w2985_
	);
	LUT2 #(
		.INIT('h2)
	) name2523 (
		_w1480_,
		_w2903_,
		_w2986_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2524 (
		_w2517_,
		_w2600_,
		_w2603_,
		_w2903_,
		_w2987_
	);
	LUT3 #(
		.INIT('ha8)
	) name2525 (
		_w1963_,
		_w2986_,
		_w2987_,
		_w2988_
	);
	LUT4 #(
		.INIT('h0c88)
	) name2526 (
		_w1480_,
		_w1869_,
		_w2625_,
		_w2903_,
		_w2989_
	);
	LUT4 #(
		.INIT('h0c88)
	) name2527 (
		_w1480_,
		_w2000_,
		_w2630_,
		_w2903_,
		_w2990_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2528 (
		_w2021_,
		_w2633_,
		_w2903_,
		_w2986_,
		_w2991_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2529 (
		_w1480_,
		_w2001_,
		_w2032_,
		_w2903_,
		_w2992_
	);
	LUT3 #(
		.INIT('h13)
	) name2530 (
		_w2001_,
		_w2029_,
		_w2903_,
		_w2993_
	);
	LUT3 #(
		.INIT('h31)
	) name2531 (
		_w1479_,
		_w2992_,
		_w2993_,
		_w2994_
	);
	LUT3 #(
		.INIT('hd0)
	) name2532 (
		_w2025_,
		_w2991_,
		_w2994_,
		_w2995_
	);
	LUT3 #(
		.INIT('h10)
	) name2533 (
		_w2989_,
		_w2990_,
		_w2995_,
		_w2996_
	);
	LUT2 #(
		.INIT('h8)
	) name2534 (
		_w1480_,
		_w2039_,
		_w2997_
	);
	LUT4 #(
		.INIT('h0075)
	) name2535 (
		_w1285_,
		_w2988_,
		_w2996_,
		_w2997_,
		_w2998_
	);
	LUT2 #(
		.INIT('h4)
	) name2536 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[27]/NET0131 ,
		_w2999_
	);
	LUT3 #(
		.INIT('h07)
	) name2537 (
		_w1480_,
		_w2344_,
		_w2999_,
		_w3000_
	);
	LUT3 #(
		.INIT('h2f)
	) name2538 (
		\P1_state_reg[0]/NET0131 ,
		_w2998_,
		_w3000_,
		_w3001_
	);
	LUT2 #(
		.INIT('h2)
	) name2539 (
		_w1444_,
		_w2903_,
		_w3002_
	);
	LUT4 #(
		.INIT('hf070)
	) name2540 (
		_w2399_,
		_w2414_,
		_w2403_,
		_w2413_,
		_w3003_
	);
	LUT2 #(
		.INIT('h8)
	) name2541 (
		_w2420_,
		_w2398_,
		_w3004_
	);
	LUT4 #(
		.INIT('h0203)
	) name2542 (
		_w2396_,
		_w2384_,
		_w2385_,
		_w2420_,
		_w3005_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2543 (
		_w2423_,
		_w3003_,
		_w3004_,
		_w3005_,
		_w3006_
	);
	LUT3 #(
		.INIT('h51)
	) name2544 (
		_w2371_,
		_w2374_,
		_w2379_,
		_w3007_
	);
	LUT4 #(
		.INIT('h8488)
	) name2545 (
		_w2522_,
		_w2903_,
		_w3006_,
		_w3007_,
		_w3008_
	);
	LUT3 #(
		.INIT('ha8)
	) name2546 (
		_w1963_,
		_w3002_,
		_w3008_,
		_w3009_
	);
	LUT2 #(
		.INIT('h1)
	) name2547 (
		_w1644_,
		_w1685_,
		_w3010_
	);
	LUT2 #(
		.INIT('h1)
	) name2548 (
		_w1707_,
		_w1718_,
		_w3011_
	);
	LUT2 #(
		.INIT('h1)
	) name2549 (
		_w1727_,
		_w1672_,
		_w3012_
	);
	LUT4 #(
		.INIT('h0001)
	) name2550 (
		_w1707_,
		_w1718_,
		_w1727_,
		_w1672_,
		_w3013_
	);
	LUT4 #(
		.INIT('h2300)
	) name2551 (
		_w1662_,
		_w1682_,
		_w3010_,
		_w3013_,
		_w3014_
	);
	LUT3 #(
		.INIT('h54)
	) name2552 (
		_w1727_,
		_w1684_,
		_w1731_,
		_w3015_
	);
	LUT3 #(
		.INIT('h0b)
	) name2553 (
		_w1707_,
		_w1730_,
		_w1734_,
		_w3016_
	);
	LUT3 #(
		.INIT('h70)
	) name2554 (
		_w3011_,
		_w3015_,
		_w3016_,
		_w3017_
	);
	LUT2 #(
		.INIT('h1)
	) name2555 (
		_w1696_,
		_w1789_,
		_w3018_
	);
	LUT3 #(
		.INIT('h0d)
	) name2556 (
		_w1740_,
		_w1747_,
		_w1775_,
		_w3019_
	);
	LUT2 #(
		.INIT('h8)
	) name2557 (
		_w3018_,
		_w3019_,
		_w3020_
	);
	LUT3 #(
		.INIT('hb0)
	) name2558 (
		_w3014_,
		_w3017_,
		_w3020_,
		_w3021_
	);
	LUT3 #(
		.INIT('h32)
	) name2559 (
		_w1733_,
		_w1789_,
		_w1794_,
		_w3022_
	);
	LUT3 #(
		.INIT('h2b)
	) name2560 (
		_w1740_,
		_w1747_,
		_w1793_,
		_w3023_
	);
	LUT3 #(
		.INIT('h70)
	) name2561 (
		_w3019_,
		_w3022_,
		_w3023_,
		_w3024_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2562 (
		_w3014_,
		_w3017_,
		_w3020_,
		_w3024_,
		_w3025_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name2563 (
		_w1752_,
		_w1759_,
		_w1834_,
		_w1839_,
		_w3026_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name2564 (
		_w1812_,
		_w1820_,
		_w1825_,
		_w1830_,
		_w3027_
	);
	LUT2 #(
		.INIT('h8)
	) name2565 (
		_w3026_,
		_w3027_,
		_w3028_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2566 (
		_w1612_,
		_w1617_,
		_w1802_,
		_w1807_,
		_w3029_
	);
	LUT3 #(
		.INIT('h10)
	) name2567 (
		_w1606_,
		_w1633_,
		_w3029_,
		_w3030_
	);
	LUT2 #(
		.INIT('h8)
	) name2568 (
		_w3028_,
		_w3030_,
		_w3031_
	);
	LUT4 #(
		.INIT('h4f04)
	) name2569 (
		_w1752_,
		_w1759_,
		_w1834_,
		_w1839_,
		_w3032_
	);
	LUT4 #(
		.INIT('hb2bb)
	) name2570 (
		_w1812_,
		_w1820_,
		_w1825_,
		_w1830_,
		_w3033_
	);
	LUT3 #(
		.INIT('h70)
	) name2571 (
		_w3027_,
		_w3032_,
		_w3033_,
		_w3034_
	);
	LUT4 #(
		.INIT('h22b2)
	) name2572 (
		_w1612_,
		_w1617_,
		_w1802_,
		_w1807_,
		_w3035_
	);
	LUT3 #(
		.INIT('h10)
	) name2573 (
		_w1606_,
		_w1633_,
		_w3035_,
		_w3036_
	);
	LUT3 #(
		.INIT('h54)
	) name2574 (
		_w1606_,
		_w1846_,
		_w1850_,
		_w3037_
	);
	LUT2 #(
		.INIT('h1)
	) name2575 (
		_w3036_,
		_w3037_,
		_w3038_
	);
	LUT4 #(
		.INIT('h000d)
	) name2576 (
		_w3030_,
		_w3034_,
		_w3036_,
		_w3037_,
		_w3039_
	);
	LUT3 #(
		.INIT('hb0)
	) name2577 (
		_w3025_,
		_w3031_,
		_w3039_,
		_w3040_
	);
	LUT2 #(
		.INIT('h1)
	) name2578 (
		_w1594_,
		_w1853_,
		_w3041_
	);
	LUT2 #(
		.INIT('h1)
	) name2579 (
		_w1553_,
		_w1567_,
		_w3042_
	);
	LUT4 #(
		.INIT('h0001)
	) name2580 (
		_w1553_,
		_w1567_,
		_w1594_,
		_w1853_,
		_w3043_
	);
	LUT2 #(
		.INIT('h8)
	) name2581 (
		_w1513_,
		_w2607_,
		_w3044_
	);
	LUT3 #(
		.INIT('h80)
	) name2582 (
		_w1513_,
		_w2607_,
		_w3043_,
		_w3045_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2583 (
		_w3025_,
		_w3031_,
		_w3039_,
		_w3045_,
		_w3046_
	);
	LUT3 #(
		.INIT('h51)
	) name2584 (
		_w1575_,
		_w1849_,
		_w1853_,
		_w3047_
	);
	LUT3 #(
		.INIT('h0b)
	) name2585 (
		_w1553_,
		_w1566_,
		_w1577_,
		_w3048_
	);
	LUT3 #(
		.INIT('hd0)
	) name2586 (
		_w3042_,
		_w3047_,
		_w3048_,
		_w3049_
	);
	LUT4 #(
		.INIT('h00fb)
	) name2587 (
		_w1529_,
		_w1534_,
		_w1542_,
		_w1580_,
		_w3050_
	);
	LUT4 #(
		.INIT('h0001)
	) name2588 (
		_w1306_,
		_w1485_,
		_w1505_,
		_w1510_,
		_w3051_
	);
	LUT4 #(
		.INIT('h0031)
	) name2589 (
		_w1513_,
		_w1582_,
		_w3050_,
		_w3051_,
		_w3052_
	);
	LUT3 #(
		.INIT('hd0)
	) name2590 (
		_w3044_,
		_w3049_,
		_w3052_,
		_w3053_
	);
	LUT4 #(
		.INIT('h4844)
	) name2591 (
		_w2522_,
		_w2903_,
		_w3046_,
		_w3053_,
		_w3054_
	);
	LUT3 #(
		.INIT('ha8)
	) name2592 (
		_w1869_,
		_w3002_,
		_w3054_,
		_w3055_
	);
	LUT4 #(
		.INIT('h9555)
	) name2593 (
		_w1400_,
		_w1988_,
		_w1978_,
		_w1987_,
		_w3056_
	);
	LUT4 #(
		.INIT('h7020)
	) name2594 (
		_w1305_,
		_w1483_,
		_w2903_,
		_w3056_,
		_w3057_
	);
	LUT4 #(
		.INIT('h9500)
	) name2595 (
		_w1442_,
		_w2016_,
		_w2020_,
		_w2903_,
		_w3058_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2596 (
		_w1444_,
		_w2001_,
		_w2032_,
		_w2903_,
		_w3059_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2597 (
		_w1306_,
		_w1441_,
		_w2993_,
		_w3059_,
		_w3060_
	);
	LUT4 #(
		.INIT('h5700)
	) name2598 (
		_w2025_,
		_w3002_,
		_w3058_,
		_w3060_,
		_w3061_
	);
	LUT4 #(
		.INIT('h5700)
	) name2599 (
		_w2000_,
		_w3002_,
		_w3057_,
		_w3061_,
		_w3062_
	);
	LUT2 #(
		.INIT('h4)
	) name2600 (
		_w3055_,
		_w3062_,
		_w3063_
	);
	LUT3 #(
		.INIT('h60)
	) name2601 (
		\P2_reg3_reg[28]/NET0131 ,
		_w1443_,
		_w2039_,
		_w3064_
	);
	LUT4 #(
		.INIT('h0075)
	) name2602 (
		_w1285_,
		_w3009_,
		_w3063_,
		_w3064_,
		_w3065_
	);
	LUT4 #(
		.INIT('h9b3b)
	) name2603 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w1267_,
		_w1443_,
		_w3066_
	);
	LUT3 #(
		.INIT('h2f)
	) name2604 (
		\P1_state_reg[0]/NET0131 ,
		_w3065_,
		_w3066_,
		_w3067_
	);
	LUT2 #(
		.INIT('h2)
	) name2605 (
		\P2_reg0_reg[25]/NET0131 ,
		_w2042_,
		_w3068_
	);
	LUT4 #(
		.INIT('h2000)
	) name2606 (
		\P2_reg0_reg[25]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3069_
	);
	LUT4 #(
		.INIT('hc535)
	) name2607 (
		\P2_reg0_reg[25]/NET0131 ,
		_w2519_,
		_w2729_,
		_w2878_,
		_w3070_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2608 (
		\P2_reg0_reg[25]/NET0131 ,
		_w1869_,
		_w2729_,
		_w2884_,
		_w3071_
	);
	LUT3 #(
		.INIT('h02)
	) name2609 (
		_w2000_,
		_w2886_,
		_w2887_,
		_w3072_
	);
	LUT2 #(
		.INIT('h2)
	) name2610 (
		\P2_reg0_reg[25]/NET0131 ,
		_w2737_,
		_w3073_
	);
	LUT4 #(
		.INIT('h005d)
	) name2611 (
		_w2729_,
		_w2893_,
		_w3072_,
		_w3073_,
		_w3074_
	);
	LUT4 #(
		.INIT('h3100)
	) name2612 (
		_w1963_,
		_w3071_,
		_w3070_,
		_w3074_,
		_w3075_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2613 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w3069_,
		_w3075_,
		_w3076_
	);
	LUT2 #(
		.INIT('he)
	) name2614 (
		_w3068_,
		_w3076_,
		_w3077_
	);
	LUT2 #(
		.INIT('h2)
	) name2615 (
		\P2_reg0_reg[27]/NET0131 ,
		_w2729_,
		_w3078_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2616 (
		_w2517_,
		_w2600_,
		_w2603_,
		_w2729_,
		_w3079_
	);
	LUT3 #(
		.INIT('ha8)
	) name2617 (
		_w1963_,
		_w3078_,
		_w3079_,
		_w3080_
	);
	LUT4 #(
		.INIT('h0c88)
	) name2618 (
		\P2_reg0_reg[27]/NET0131 ,
		_w1869_,
		_w2625_,
		_w2729_,
		_w3081_
	);
	LUT3 #(
		.INIT('hd0)
	) name2619 (
		_w2001_,
		_w2729_,
		_w2734_,
		_w3082_
	);
	LUT2 #(
		.INIT('h2)
	) name2620 (
		_w2025_,
		_w2729_,
		_w3083_
	);
	LUT4 #(
		.INIT('hf100)
	) name2621 (
		_w2001_,
		_w2025_,
		_w2729_,
		_w2734_,
		_w3084_
	);
	LUT3 #(
		.INIT('h8a)
	) name2622 (
		\P2_reg0_reg[27]/NET0131 ,
		_w2736_,
		_w3084_,
		_w3085_
	);
	LUT4 #(
		.INIT('h2f00)
	) name2623 (
		_w2000_,
		_w2630_,
		_w2634_,
		_w2729_,
		_w3086_
	);
	LUT3 #(
		.INIT('h01)
	) name2624 (
		_w3081_,
		_w3085_,
		_w3086_,
		_w3087_
	);
	LUT4 #(
		.INIT('h2000)
	) name2625 (
		\P2_reg0_reg[27]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3088_
	);
	LUT4 #(
		.INIT('h0075)
	) name2626 (
		_w1285_,
		_w3080_,
		_w3087_,
		_w3088_,
		_w3089_
	);
	LUT2 #(
		.INIT('h2)
	) name2627 (
		\P2_reg0_reg[27]/NET0131 ,
		_w2042_,
		_w3090_
	);
	LUT3 #(
		.INIT('hf2)
	) name2628 (
		\P1_state_reg[0]/NET0131 ,
		_w3089_,
		_w3090_,
		_w3091_
	);
	LUT4 #(
		.INIT('h2300)
	) name2629 (
		_w1662_,
		_w1682_,
		_w3010_,
		_w3012_,
		_w3092_
	);
	LUT4 #(
		.INIT('h0001)
	) name2630 (
		_w1696_,
		_w1707_,
		_w1718_,
		_w1789_,
		_w3093_
	);
	LUT3 #(
		.INIT('h0b)
	) name2631 (
		_w3016_,
		_w3018_,
		_w3022_,
		_w3094_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2632 (
		_w3015_,
		_w3092_,
		_w3093_,
		_w3094_,
		_w3095_
	);
	LUT2 #(
		.INIT('h8)
	) name2633 (
		_w3019_,
		_w3026_,
		_w3096_
	);
	LUT3 #(
		.INIT('h0b)
	) name2634 (
		_w3023_,
		_w3026_,
		_w3032_,
		_w3097_
	);
	LUT2 #(
		.INIT('h8)
	) name2635 (
		_w3027_,
		_w3029_,
		_w3098_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2636 (
		_w3095_,
		_w3096_,
		_w3097_,
		_w3098_,
		_w3099_
	);
	LUT3 #(
		.INIT('h0d)
	) name2637 (
		_w3029_,
		_w3033_,
		_w3035_,
		_w3100_
	);
	LUT4 #(
		.INIT('h0001)
	) name2638 (
		_w1594_,
		_w1606_,
		_w1633_,
		_w1853_,
		_w3101_
	);
	LUT2 #(
		.INIT('h4)
	) name2639 (
		_w1567_,
		_w2608_,
		_w3102_
	);
	LUT3 #(
		.INIT('h40)
	) name2640 (
		_w1567_,
		_w2608_,
		_w3101_,
		_w3103_
	);
	LUT3 #(
		.INIT('h70)
	) name2641 (
		_w3037_,
		_w3041_,
		_w3047_,
		_w3104_
	);
	LUT3 #(
		.INIT('hd0)
	) name2642 (
		_w2607_,
		_w3048_,
		_w3050_,
		_w3105_
	);
	LUT3 #(
		.INIT('hd0)
	) name2643 (
		_w3102_,
		_w3104_,
		_w3105_,
		_w3106_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2644 (
		_w3099_,
		_w3100_,
		_w3103_,
		_w3106_,
		_w3107_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2645 (
		\P2_reg0_reg[26]/NET0131 ,
		_w2514_,
		_w2729_,
		_w3107_,
		_w3108_
	);
	LUT2 #(
		.INIT('h2)
	) name2646 (
		_w1869_,
		_w3108_,
		_w3109_
	);
	LUT2 #(
		.INIT('h8)
	) name2647 (
		_w2391_,
		_w2419_,
		_w3110_
	);
	LUT2 #(
		.INIT('h8)
	) name2648 (
		_w2399_,
		_w2397_,
		_w3111_
	);
	LUT4 #(
		.INIT('h8000)
	) name2649 (
		_w2391_,
		_w2399_,
		_w2397_,
		_w2419_,
		_w3112_
	);
	LUT4 #(
		.INIT('hce00)
	) name2650 (
		_w2414_,
		_w2400_,
		_w2413_,
		_w3112_,
		_w3113_
	);
	LUT3 #(
		.INIT('h07)
	) name2651 (
		_w2395_,
		_w2419_,
		_w2383_,
		_w3114_
	);
	LUT3 #(
		.INIT('h15)
	) name2652 (
		_w2393_,
		_w2397_,
		_w2402_,
		_w3115_
	);
	LUT3 #(
		.INIT('hc4)
	) name2653 (
		_w3110_,
		_w3114_,
		_w3115_,
		_w3116_
	);
	LUT2 #(
		.INIT('h8)
	) name2654 (
		_w2375_,
		_w2373_,
		_w3117_
	);
	LUT4 #(
		.INIT('h0001)
	) name2655 (
		_w1909_,
		_w1910_,
		_w1911_,
		_w1943_,
		_w3118_
	);
	LUT3 #(
		.INIT('h80)
	) name2656 (
		_w2375_,
		_w2373_,
		_w3118_,
		_w3119_
	);
	LUT3 #(
		.INIT('h4c)
	) name2657 (
		_w2380_,
		_w2376_,
		_w2385_,
		_w3120_
	);
	LUT3 #(
		.INIT('h13)
	) name2658 (
		_w2373_,
		_w2370_,
		_w2378_,
		_w3121_
	);
	LUT3 #(
		.INIT('hd0)
	) name2659 (
		_w3117_,
		_w3120_,
		_w3121_,
		_w3122_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2660 (
		_w3113_,
		_w3116_,
		_w3119_,
		_w3122_,
		_w3123_
	);
	LUT4 #(
		.INIT('hc535)
	) name2661 (
		\P2_reg0_reg[26]/NET0131 ,
		_w2514_,
		_w2729_,
		_w3123_,
		_w3124_
	);
	LUT4 #(
		.INIT('h6555)
	) name2662 (
		_w1483_,
		_w1510_,
		_w1978_,
		_w1987_,
		_w3125_
	);
	LUT4 #(
		.INIT('h7020)
	) name2663 (
		_w1305_,
		_w1527_,
		_w2000_,
		_w3125_,
		_w3126_
	);
	LUT3 #(
		.INIT('h10)
	) name2664 (
		_w1306_,
		_w1505_,
		_w2001_,
		_w3127_
	);
	LUT4 #(
		.INIT('h007b)
	) name2665 (
		_w1506_,
		_w2025_,
		_w2632_,
		_w3127_,
		_w3128_
	);
	LUT3 #(
		.INIT('h8a)
	) name2666 (
		\P2_reg0_reg[26]/NET0131 ,
		_w2736_,
		_w3084_,
		_w3129_
	);
	LUT4 #(
		.INIT('h0075)
	) name2667 (
		_w2729_,
		_w3126_,
		_w3128_,
		_w3129_,
		_w3130_
	);
	LUT3 #(
		.INIT('hd0)
	) name2668 (
		_w1963_,
		_w3124_,
		_w3130_,
		_w3131_
	);
	LUT4 #(
		.INIT('h2000)
	) name2669 (
		\P2_reg0_reg[26]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3132_
	);
	LUT4 #(
		.INIT('h0075)
	) name2670 (
		_w1285_,
		_w3109_,
		_w3131_,
		_w3132_,
		_w3133_
	);
	LUT2 #(
		.INIT('h2)
	) name2671 (
		\P2_reg0_reg[26]/NET0131 ,
		_w2042_,
		_w3134_
	);
	LUT3 #(
		.INIT('hf2)
	) name2672 (
		\P1_state_reg[0]/NET0131 ,
		_w3133_,
		_w3134_,
		_w3135_
	);
	LUT2 #(
		.INIT('h2)
	) name2673 (
		\P2_reg0_reg[28]/NET0131 ,
		_w2729_,
		_w3136_
	);
	LUT4 #(
		.INIT('h8488)
	) name2674 (
		_w2522_,
		_w2729_,
		_w3006_,
		_w3007_,
		_w3137_
	);
	LUT3 #(
		.INIT('ha8)
	) name2675 (
		_w1963_,
		_w3136_,
		_w3137_,
		_w3138_
	);
	LUT4 #(
		.INIT('h7020)
	) name2676 (
		_w1305_,
		_w1483_,
		_w2729_,
		_w3056_,
		_w3139_
	);
	LUT3 #(
		.INIT('ha8)
	) name2677 (
		_w2000_,
		_w3136_,
		_w3139_,
		_w3140_
	);
	LUT4 #(
		.INIT('h4844)
	) name2678 (
		_w2522_,
		_w2729_,
		_w3046_,
		_w3053_,
		_w3141_
	);
	LUT4 #(
		.INIT('h9500)
	) name2679 (
		_w1442_,
		_w2016_,
		_w2020_,
		_w2729_,
		_w3142_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2680 (
		\P2_reg0_reg[28]/NET0131 ,
		_w2001_,
		_w2729_,
		_w2734_,
		_w3143_
	);
	LUT4 #(
		.INIT('h1000)
	) name2681 (
		_w1306_,
		_w1441_,
		_w2001_,
		_w2729_,
		_w3144_
	);
	LUT2 #(
		.INIT('h1)
	) name2682 (
		_w3143_,
		_w3144_,
		_w3145_
	);
	LUT4 #(
		.INIT('h5700)
	) name2683 (
		_w2025_,
		_w3136_,
		_w3142_,
		_w3145_,
		_w3146_
	);
	LUT4 #(
		.INIT('h5700)
	) name2684 (
		_w1869_,
		_w3136_,
		_w3141_,
		_w3146_,
		_w3147_
	);
	LUT2 #(
		.INIT('h4)
	) name2685 (
		_w3140_,
		_w3147_,
		_w3148_
	);
	LUT4 #(
		.INIT('h2000)
	) name2686 (
		\P2_reg0_reg[28]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3149_
	);
	LUT4 #(
		.INIT('h0075)
	) name2687 (
		_w1285_,
		_w3138_,
		_w3148_,
		_w3149_,
		_w3150_
	);
	LUT2 #(
		.INIT('h2)
	) name2688 (
		\P2_reg0_reg[28]/NET0131 ,
		_w2042_,
		_w3151_
	);
	LUT3 #(
		.INIT('hf2)
	) name2689 (
		\P1_state_reg[0]/NET0131 ,
		_w3150_,
		_w3151_,
		_w3152_
	);
	LUT2 #(
		.INIT('h8)
	) name2690 (
		_w2556_,
		_w2729_,
		_w3153_
	);
	LUT3 #(
		.INIT('h09)
	) name2691 (
		_w1863_,
		_w1866_,
		_w1999_,
		_w3154_
	);
	LUT3 #(
		.INIT('ha8)
	) name2692 (
		_w2556_,
		_w2729_,
		_w3154_,
		_w3155_
	);
	LUT3 #(
		.INIT('h2a)
	) name2693 (
		\P2_reg0_reg[31]/NET0131 ,
		_w3082_,
		_w3155_,
		_w3156_
	);
	LUT4 #(
		.INIT('hffb0)
	) name2694 (
		_w2551_,
		_w2554_,
		_w3153_,
		_w3156_,
		_w3157_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2695 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[20]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3158_
	);
	LUT2 #(
		.INIT('h8)
	) name2696 (
		\P1_reg2_reg[20]/NET0131 ,
		_w2183_,
		_w3159_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2697 (
		\P1_reg2_reg[20]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3160_
	);
	LUT4 #(
		.INIT('h6500)
	) name2698 (
		_w1228_,
		_w2093_,
		_w2102_,
		_w2189_,
		_w3161_
	);
	LUT3 #(
		.INIT('ha8)
	) name2699 (
		_w2121_,
		_w3160_,
		_w3161_,
		_w3162_
	);
	LUT4 #(
		.INIT('h1444)
	) name2700 (
		_w488_,
		_w800_,
		_w2140_,
		_w2213_,
		_w3163_
	);
	LUT2 #(
		.INIT('h8)
	) name2701 (
		_w488_,
		_w724_,
		_w3164_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2702 (
		\P1_reg2_reg[20]/NET0131 ,
		_w2189_,
		_w3163_,
		_w3164_,
		_w3165_
	);
	LUT2 #(
		.INIT('h2)
	) name2703 (
		_w1237_,
		_w3165_,
		_w3166_
	);
	LUT3 #(
		.INIT('h10)
	) name2704 (
		_w489_,
		_w804_,
		_w2194_,
		_w3167_
	);
	LUT3 #(
		.INIT('h80)
	) name2705 (
		_w720_,
		_w2153_,
		_w2163_,
		_w3168_
	);
	LUT4 #(
		.INIT('h2000)
	) name2706 (
		_w720_,
		_w805_,
		_w2153_,
		_w2163_,
		_w3169_
	);
	LUT4 #(
		.INIT('h070b)
	) name2707 (
		_w805_,
		_w2170_,
		_w3167_,
		_w3168_,
		_w3170_
	);
	LUT4 #(
		.INIT('h9f00)
	) name2708 (
		_w1228_,
		_w2124_,
		_w2128_,
		_w3170_,
		_w3171_
	);
	LUT2 #(
		.INIT('h8)
	) name2709 (
		_w806_,
		_w1120_,
		_w3172_
	);
	LUT4 #(
		.INIT('hfb00)
	) name2710 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2172_,
		_w3173_
	);
	LUT4 #(
		.INIT('hfb00)
	) name2711 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2128_,
		_w3174_
	);
	LUT3 #(
		.INIT('h01)
	) name2712 (
		_w2171_,
		_w3173_,
		_w3174_,
		_w3175_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2713 (
		\P1_reg2_reg[20]/NET0131 ,
		_w2171_,
		_w3173_,
		_w3174_,
		_w3176_
	);
	LUT2 #(
		.INIT('h1)
	) name2714 (
		_w3172_,
		_w3176_,
		_w3177_
	);
	LUT3 #(
		.INIT('hd0)
	) name2715 (
		_w2189_,
		_w3171_,
		_w3177_,
		_w3178_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2716 (
		_w2182_,
		_w3166_,
		_w3162_,
		_w3178_,
		_w3179_
	);
	LUT4 #(
		.INIT('heeec)
	) name2717 (
		\P1_state_reg[0]/NET0131 ,
		_w3158_,
		_w3159_,
		_w3179_,
		_w3180_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2718 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[25]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3181_
	);
	LUT2 #(
		.INIT('h8)
	) name2719 (
		\P1_reg2_reg[25]/NET0131 ,
		_w2183_,
		_w3182_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2720 (
		\P1_reg2_reg[25]/NET0131 ,
		_w2121_,
		_w2189_,
		_w2706_,
		_w3183_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2721 (
		\P1_reg2_reg[25]/NET0131 ,
		_w2189_,
		_w2708_,
		_w2709_,
		_w3184_
	);
	LUT2 #(
		.INIT('h2)
	) name2722 (
		_w1237_,
		_w3184_,
		_w3185_
	);
	LUT2 #(
		.INIT('h8)
	) name2723 (
		_w1060_,
		_w1120_,
		_w3186_
	);
	LUT4 #(
		.INIT('hfb00)
	) name2724 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2170_,
		_w3187_
	);
	LUT4 #(
		.INIT('h0001)
	) name2725 (
		_w2171_,
		_w2196_,
		_w3174_,
		_w3187_,
		_w3188_
	);
	LUT3 #(
		.INIT('h31)
	) name2726 (
		\P1_reg2_reg[25]/NET0131 ,
		_w3186_,
		_w3188_,
		_w3189_
	);
	LUT4 #(
		.INIT('h7500)
	) name2727 (
		_w2189_,
		_w2801_,
		_w2803_,
		_w3189_,
		_w3190_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2728 (
		_w2182_,
		_w3183_,
		_w3185_,
		_w3190_,
		_w3191_
	);
	LUT4 #(
		.INIT('heeec)
	) name2729 (
		\P1_state_reg[0]/NET0131 ,
		_w3181_,
		_w3182_,
		_w3191_,
		_w3192_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2730 (
		\P1_reg2_reg[27]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3193_
	);
	LUT4 #(
		.INIT('hc535)
	) name2731 (
		\P1_reg2_reg[27]/NET0131 ,
		_w1165_,
		_w2189_,
		_w2952_,
		_w3194_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2732 (
		\P1_reg2_reg[27]/NET0131 ,
		_w2189_,
		_w2954_,
		_w2955_,
		_w3195_
	);
	LUT2 #(
		.INIT('h2)
	) name2733 (
		_w1237_,
		_w3195_,
		_w3196_
	);
	LUT4 #(
		.INIT('h4844)
	) name2734 (
		_w1165_,
		_w2189_,
		_w2967_,
		_w2974_,
		_w3197_
	);
	LUT4 #(
		.INIT('h9050)
	) name2735 (
		_w1041_,
		_w2166_,
		_w2189_,
		_w2860_,
		_w3198_
	);
	LUT4 #(
		.INIT('h1000)
	) name2736 (
		_w489_,
		_w1040_,
		_w2189_,
		_w2194_,
		_w3199_
	);
	LUT3 #(
		.INIT('h60)
	) name2737 (
		\P1_reg3_reg[27]/NET0131 ,
		_w703_,
		_w1120_,
		_w3200_
	);
	LUT4 #(
		.INIT('h0057)
	) name2738 (
		\P1_reg2_reg[27]/NET0131 ,
		_w2171_,
		_w2196_,
		_w3200_,
		_w3201_
	);
	LUT2 #(
		.INIT('h4)
	) name2739 (
		_w3199_,
		_w3201_,
		_w3202_
	);
	LUT4 #(
		.INIT('h5700)
	) name2740 (
		_w2170_,
		_w3193_,
		_w3198_,
		_w3202_,
		_w3203_
	);
	LUT4 #(
		.INIT('h5700)
	) name2741 (
		_w2121_,
		_w3193_,
		_w3197_,
		_w3203_,
		_w3204_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2742 (
		_w2128_,
		_w3194_,
		_w3196_,
		_w3204_,
		_w3205_
	);
	LUT2 #(
		.INIT('h8)
	) name2743 (
		\P1_reg2_reg[27]/NET0131 ,
		_w2183_,
		_w3206_
	);
	LUT4 #(
		.INIT('haa08)
	) name2744 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w3205_,
		_w3206_,
		_w3207_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2745 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[27]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3208_
	);
	LUT2 #(
		.INIT('he)
	) name2746 (
		_w3207_,
		_w3208_,
		_w3209_
	);
	LUT2 #(
		.INIT('h2)
	) name2747 (
		\P2_reg1_reg[24]/NET0131 ,
		_w2042_,
		_w3210_
	);
	LUT4 #(
		.INIT('h2000)
	) name2748 (
		\P2_reg1_reg[24]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3211_
	);
	LUT4 #(
		.INIT('h40f0)
	) name2749 (
		_w3024_,
		_w3028_,
		_w3030_,
		_w3034_,
		_w3212_
	);
	LUT4 #(
		.INIT('h0070)
	) name2750 (
		_w3021_,
		_w3031_,
		_w3038_,
		_w3212_,
		_w3213_
	);
	LUT4 #(
		.INIT('h5a9a)
	) name2751 (
		_w2518_,
		_w3043_,
		_w3049_,
		_w3213_,
		_w3214_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2752 (
		\P2_reg1_reg[24]/NET0131 ,
		_w1869_,
		_w2762_,
		_w3214_,
		_w3215_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2753 (
		_w2396_,
		_w2420_,
		_w2398_,
		_w2403_,
		_w3216_
	);
	LUT4 #(
		.INIT('h22a2)
	) name2754 (
		_w2379_,
		_w2381_,
		_w2386_,
		_w3216_,
		_w3217_
	);
	LUT4 #(
		.INIT('h780f)
	) name2755 (
		_w2464_,
		_w2465_,
		_w2518_,
		_w3217_,
		_w3218_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2756 (
		\P2_reg1_reg[24]/NET0131 ,
		_w1963_,
		_w2762_,
		_w3218_,
		_w3219_
	);
	LUT4 #(
		.INIT('h5400)
	) name2757 (
		_w1306_,
		_w1531_,
		_w1533_,
		_w2001_,
		_w3220_
	);
	LUT4 #(
		.INIT('h1444)
	) name2758 (
		_w1305_,
		_w1527_,
		_w1978_,
		_w1986_,
		_w3221_
	);
	LUT3 #(
		.INIT('h70)
	) name2759 (
		_w1305_,
		_w1551_,
		_w2000_,
		_w3222_
	);
	LUT3 #(
		.INIT('h84)
	) name2760 (
		_w1534_,
		_w2025_,
		_w2890_,
		_w3223_
	);
	LUT4 #(
		.INIT('h0045)
	) name2761 (
		_w3220_,
		_w3221_,
		_w3222_,
		_w3223_,
		_w3224_
	);
	LUT3 #(
		.INIT('hc4)
	) name2762 (
		_w2033_,
		_w2734_,
		_w2762_,
		_w3225_
	);
	LUT4 #(
		.INIT('hf010)
	) name2763 (
		_w2000_,
		_w2033_,
		_w2734_,
		_w2762_,
		_w3226_
	);
	LUT2 #(
		.INIT('h2)
	) name2764 (
		\P2_reg1_reg[24]/NET0131 ,
		_w3226_,
		_w3227_
	);
	LUT3 #(
		.INIT('h0d)
	) name2765 (
		_w2762_,
		_w3224_,
		_w3227_,
		_w3228_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2766 (
		_w1285_,
		_w3219_,
		_w3215_,
		_w3228_,
		_w3229_
	);
	LUT4 #(
		.INIT('heeec)
	) name2767 (
		\P1_state_reg[0]/NET0131 ,
		_w3210_,
		_w3211_,
		_w3229_,
		_w3230_
	);
	LUT2 #(
		.INIT('h2)
	) name2768 (
		\P2_reg1_reg[26]/NET0131 ,
		_w2042_,
		_w3231_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2769 (
		\P2_reg1_reg[26]/NET0131 ,
		_w2514_,
		_w2762_,
		_w3107_,
		_w3232_
	);
	LUT2 #(
		.INIT('h2)
	) name2770 (
		_w1869_,
		_w3232_,
		_w3233_
	);
	LUT4 #(
		.INIT('hc535)
	) name2771 (
		\P2_reg1_reg[26]/NET0131 ,
		_w2514_,
		_w2762_,
		_w3123_,
		_w3234_
	);
	LUT2 #(
		.INIT('h2)
	) name2772 (
		\P2_reg1_reg[26]/NET0131 ,
		_w3226_,
		_w3235_
	);
	LUT4 #(
		.INIT('h0075)
	) name2773 (
		_w2762_,
		_w3126_,
		_w3128_,
		_w3235_,
		_w3236_
	);
	LUT3 #(
		.INIT('hd0)
	) name2774 (
		_w1963_,
		_w3234_,
		_w3236_,
		_w3237_
	);
	LUT4 #(
		.INIT('h2000)
	) name2775 (
		\P2_reg1_reg[26]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3238_
	);
	LUT4 #(
		.INIT('h0075)
	) name2776 (
		_w1285_,
		_w3233_,
		_w3237_,
		_w3238_,
		_w3239_
	);
	LUT3 #(
		.INIT('hce)
	) name2777 (
		\P1_state_reg[0]/NET0131 ,
		_w3231_,
		_w3239_,
		_w3240_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name2778 (
		_w2001_,
		_w2734_,
		_w2762_,
		_w3154_,
		_w3241_
	);
	LUT3 #(
		.INIT('h2a)
	) name2779 (
		\P2_reg1_reg[27]/NET0131 ,
		_w2556_,
		_w3241_,
		_w3242_
	);
	LUT2 #(
		.INIT('h8)
	) name2780 (
		_w1285_,
		_w2762_,
		_w3243_
	);
	LUT3 #(
		.INIT('h80)
	) name2781 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w2762_,
		_w3244_
	);
	LUT4 #(
		.INIT('h8288)
	) name2782 (
		_w1963_,
		_w2517_,
		_w2600_,
		_w2603_,
		_w3245_
	);
	LUT2 #(
		.INIT('h2)
	) name2783 (
		_w1869_,
		_w2625_,
		_w3246_
	);
	LUT4 #(
		.INIT('hccc4)
	) name2784 (
		_w2635_,
		_w3244_,
		_w3246_,
		_w3245_,
		_w3247_
	);
	LUT2 #(
		.INIT('he)
	) name2785 (
		_w3242_,
		_w3247_,
		_w3248_
	);
	LUT2 #(
		.INIT('h2)
	) name2786 (
		\P2_reg1_reg[28]/NET0131 ,
		_w2762_,
		_w3249_
	);
	LUT4 #(
		.INIT('h8488)
	) name2787 (
		_w2522_,
		_w2762_,
		_w3006_,
		_w3007_,
		_w3250_
	);
	LUT3 #(
		.INIT('ha8)
	) name2788 (
		_w1963_,
		_w3249_,
		_w3250_,
		_w3251_
	);
	LUT4 #(
		.INIT('h7020)
	) name2789 (
		_w1305_,
		_w1483_,
		_w2762_,
		_w3056_,
		_w3252_
	);
	LUT3 #(
		.INIT('ha8)
	) name2790 (
		_w2000_,
		_w3249_,
		_w3252_,
		_w3253_
	);
	LUT4 #(
		.INIT('h4844)
	) name2791 (
		_w2522_,
		_w2762_,
		_w3046_,
		_w3053_,
		_w3254_
	);
	LUT4 #(
		.INIT('h9500)
	) name2792 (
		_w1442_,
		_w2016_,
		_w2020_,
		_w2762_,
		_w3255_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2793 (
		\P2_reg1_reg[28]/NET0131 ,
		_w2001_,
		_w2734_,
		_w2762_,
		_w3256_
	);
	LUT4 #(
		.INIT('h1000)
	) name2794 (
		_w1306_,
		_w1441_,
		_w2001_,
		_w2762_,
		_w3257_
	);
	LUT2 #(
		.INIT('h1)
	) name2795 (
		_w3256_,
		_w3257_,
		_w3258_
	);
	LUT4 #(
		.INIT('h5700)
	) name2796 (
		_w2025_,
		_w3249_,
		_w3255_,
		_w3258_,
		_w3259_
	);
	LUT4 #(
		.INIT('h5700)
	) name2797 (
		_w1869_,
		_w3249_,
		_w3254_,
		_w3259_,
		_w3260_
	);
	LUT2 #(
		.INIT('h4)
	) name2798 (
		_w3253_,
		_w3260_,
		_w3261_
	);
	LUT4 #(
		.INIT('h2000)
	) name2799 (
		\P2_reg1_reg[28]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3262_
	);
	LUT4 #(
		.INIT('h0075)
	) name2800 (
		_w1285_,
		_w3251_,
		_w3261_,
		_w3262_,
		_w3263_
	);
	LUT2 #(
		.INIT('h2)
	) name2801 (
		\P2_reg1_reg[28]/NET0131 ,
		_w2042_,
		_w3264_
	);
	LUT3 #(
		.INIT('hf2)
	) name2802 (
		\P1_state_reg[0]/NET0131 ,
		_w3263_,
		_w3264_,
		_w3265_
	);
	LUT3 #(
		.INIT('h19)
	) name2803 (
		_w1863_,
		_w1866_,
		_w1999_,
		_w3266_
	);
	LUT3 #(
		.INIT('ha8)
	) name2804 (
		_w2556_,
		_w2762_,
		_w3266_,
		_w3267_
	);
	LUT3 #(
		.INIT('h2a)
	) name2805 (
		\P2_reg1_reg[31]/NET0131 ,
		_w3225_,
		_w3267_,
		_w3268_
	);
	LUT4 #(
		.INIT('hffb0)
	) name2806 (
		_w2551_,
		_w2554_,
		_w3244_,
		_w3268_,
		_w3269_
	);
	LUT2 #(
		.INIT('h2)
	) name2807 (
		\P2_reg2_reg[28]/NET0131 ,
		_w1298_,
		_w3270_
	);
	LUT4 #(
		.INIT('h8288)
	) name2808 (
		_w1298_,
		_w2522_,
		_w3006_,
		_w3007_,
		_w3271_
	);
	LUT3 #(
		.INIT('ha8)
	) name2809 (
		_w1963_,
		_w3270_,
		_w3271_,
		_w3272_
	);
	LUT4 #(
		.INIT('h2822)
	) name2810 (
		_w1298_,
		_w2522_,
		_w3046_,
		_w3053_,
		_w3273_
	);
	LUT3 #(
		.INIT('ha8)
	) name2811 (
		_w1869_,
		_w3270_,
		_w3273_,
		_w3274_
	);
	LUT4 #(
		.INIT('h2a08)
	) name2812 (
		_w1298_,
		_w1305_,
		_w1483_,
		_w3056_,
		_w3275_
	);
	LUT4 #(
		.INIT('h8222)
	) name2813 (
		_w1298_,
		_w1442_,
		_w2016_,
		_w2020_,
		_w3276_
	);
	LUT4 #(
		.INIT('h0200)
	) name2814 (
		_w1298_,
		_w1306_,
		_w1441_,
		_w2001_,
		_w3277_
	);
	LUT4 #(
		.INIT('haa20)
	) name2815 (
		\P2_reg2_reg[28]/NET0131 ,
		_w1298_,
		_w2001_,
		_w2032_,
		_w3278_
	);
	LUT3 #(
		.INIT('h60)
	) name2816 (
		\P2_reg3_reg[28]/NET0131 ,
		_w1443_,
		_w2029_,
		_w3279_
	);
	LUT2 #(
		.INIT('h1)
	) name2817 (
		_w3278_,
		_w3279_,
		_w3280_
	);
	LUT2 #(
		.INIT('h4)
	) name2818 (
		_w3277_,
		_w3280_,
		_w3281_
	);
	LUT4 #(
		.INIT('h5700)
	) name2819 (
		_w2025_,
		_w3270_,
		_w3276_,
		_w3281_,
		_w3282_
	);
	LUT4 #(
		.INIT('h5700)
	) name2820 (
		_w2000_,
		_w3270_,
		_w3275_,
		_w3282_,
		_w3283_
	);
	LUT2 #(
		.INIT('h4)
	) name2821 (
		_w3274_,
		_w3283_,
		_w3284_
	);
	LUT4 #(
		.INIT('h2000)
	) name2822 (
		\P2_reg2_reg[28]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3285_
	);
	LUT4 #(
		.INIT('h0075)
	) name2823 (
		_w1285_,
		_w3272_,
		_w3284_,
		_w3285_,
		_w3286_
	);
	LUT2 #(
		.INIT('h2)
	) name2824 (
		\P2_reg2_reg[28]/NET0131 ,
		_w2042_,
		_w3287_
	);
	LUT3 #(
		.INIT('hf2)
	) name2825 (
		\P1_state_reg[0]/NET0131 ,
		_w3286_,
		_w3287_,
		_w3288_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2826 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[26]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3289_
	);
	LUT2 #(
		.INIT('h8)
	) name2827 (
		\P1_reg0_reg[26]/NET0131 ,
		_w2183_,
		_w3290_
	);
	LUT4 #(
		.INIT('h4555)
	) name2828 (
		\P1_reg0_reg[26]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3291_
	);
	LUT2 #(
		.INIT('h2)
	) name2829 (
		_w2128_,
		_w3291_,
		_w3292_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2830 (
		_w1224_,
		_w2325_,
		_w2665_,
		_w3292_,
		_w3293_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2831 (
		_w2325_,
		_w2813_,
		_w2812_,
		_w2814_,
		_w3294_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2832 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2819_,
		_w3295_
	);
	LUT4 #(
		.INIT('h0002)
	) name2833 (
		_w2332_,
		_w2333_,
		_w2796_,
		_w3295_,
		_w3296_
	);
	LUT2 #(
		.INIT('h2)
	) name2834 (
		\P1_reg0_reg[26]/NET0131 ,
		_w3296_,
		_w3297_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2835 (
		_w2182_,
		_w3294_,
		_w3297_,
		_w3293_,
		_w3298_
	);
	LUT4 #(
		.INIT('heeec)
	) name2836 (
		\P1_state_reg[0]/NET0131 ,
		_w3289_,
		_w3290_,
		_w3298_,
		_w3299_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name2837 (
		\P1_reg0_reg[27]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3300_
	);
	LUT4 #(
		.INIT('hc535)
	) name2838 (
		\P1_reg0_reg[27]/NET0131 ,
		_w1165_,
		_w2325_,
		_w2952_,
		_w3301_
	);
	LUT4 #(
		.INIT('h4844)
	) name2839 (
		_w1165_,
		_w2325_,
		_w2967_,
		_w2974_,
		_w3302_
	);
	LUT3 #(
		.INIT('ha8)
	) name2840 (
		_w2121_,
		_w3300_,
		_w3302_,
		_w3303_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2841 (
		\P1_reg0_reg[27]/NET0131 ,
		_w2325_,
		_w2954_,
		_w2955_,
		_w3304_
	);
	LUT4 #(
		.INIT('h9050)
	) name2842 (
		_w1041_,
		_w2166_,
		_w2325_,
		_w2860_,
		_w3305_
	);
	LUT3 #(
		.INIT('ha2)
	) name2843 (
		\P1_reg0_reg[27]/NET0131 ,
		_w2332_,
		_w2333_,
		_w3306_
	);
	LUT4 #(
		.INIT('h1000)
	) name2844 (
		_w489_,
		_w1040_,
		_w2194_,
		_w2325_,
		_w3307_
	);
	LUT2 #(
		.INIT('h1)
	) name2845 (
		_w3306_,
		_w3307_,
		_w3308_
	);
	LUT4 #(
		.INIT('h5700)
	) name2846 (
		_w2170_,
		_w3300_,
		_w3305_,
		_w3308_,
		_w3309_
	);
	LUT3 #(
		.INIT('hd0)
	) name2847 (
		_w1237_,
		_w3304_,
		_w3309_,
		_w3310_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2848 (
		_w2128_,
		_w3301_,
		_w3303_,
		_w3310_,
		_w3311_
	);
	LUT2 #(
		.INIT('h8)
	) name2849 (
		\P1_reg0_reg[27]/NET0131 ,
		_w2183_,
		_w3312_
	);
	LUT4 #(
		.INIT('haa08)
	) name2850 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w3311_,
		_w3312_,
		_w3313_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2851 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[27]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3314_
	);
	LUT2 #(
		.INIT('he)
	) name2852 (
		_w3313_,
		_w3314_,
		_w3315_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2853 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[25]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3316_
	);
	LUT2 #(
		.INIT('h8)
	) name2854 (
		\P1_reg1_reg[25]/NET0131 ,
		_w2183_,
		_w3317_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2855 (
		\P1_reg1_reg[25]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3318_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2856 (
		\P1_reg1_reg[25]/NET0131 ,
		_w2121_,
		_w2536_,
		_w2706_,
		_w3319_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2857 (
		\P1_reg1_reg[25]/NET0131 ,
		_w2536_,
		_w2708_,
		_w2709_,
		_w3320_
	);
	LUT2 #(
		.INIT('h2)
	) name2858 (
		_w1237_,
		_w3320_,
		_w3321_
	);
	LUT4 #(
		.INIT('h8488)
	) name2859 (
		_w1221_,
		_w2536_,
		_w2713_,
		_w2715_,
		_w3322_
	);
	LUT4 #(
		.INIT('hc808)
	) name2860 (
		\P1_reg1_reg[25]/NET0131 ,
		_w2170_,
		_w2536_,
		_w2717_,
		_w3323_
	);
	LUT4 #(
		.INIT('h1000)
	) name2861 (
		_w489_,
		_w1058_,
		_w2194_,
		_w2536_,
		_w3324_
	);
	LUT3 #(
		.INIT('ha2)
	) name2862 (
		\P1_reg1_reg[25]/NET0131 ,
		_w2332_,
		_w2544_,
		_w3325_
	);
	LUT2 #(
		.INIT('h1)
	) name2863 (
		_w3324_,
		_w3325_,
		_w3326_
	);
	LUT2 #(
		.INIT('h4)
	) name2864 (
		_w3323_,
		_w3326_,
		_w3327_
	);
	LUT4 #(
		.INIT('h5700)
	) name2865 (
		_w2128_,
		_w3318_,
		_w3322_,
		_w3327_,
		_w3328_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2866 (
		_w2182_,
		_w3319_,
		_w3321_,
		_w3328_,
		_w3329_
	);
	LUT4 #(
		.INIT('heeec)
	) name2867 (
		\P1_state_reg[0]/NET0131 ,
		_w3316_,
		_w3317_,
		_w3329_,
		_w3330_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2868 (
		\P1_reg1_reg[27]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3331_
	);
	LUT4 #(
		.INIT('hc535)
	) name2869 (
		\P1_reg1_reg[27]/NET0131 ,
		_w1165_,
		_w2536_,
		_w2952_,
		_w3332_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2870 (
		\P1_reg1_reg[27]/NET0131 ,
		_w2536_,
		_w2954_,
		_w2955_,
		_w3333_
	);
	LUT2 #(
		.INIT('h2)
	) name2871 (
		_w1237_,
		_w3333_,
		_w3334_
	);
	LUT4 #(
		.INIT('h4844)
	) name2872 (
		_w1165_,
		_w2536_,
		_w2967_,
		_w2974_,
		_w3335_
	);
	LUT4 #(
		.INIT('h9050)
	) name2873 (
		_w1041_,
		_w2166_,
		_w2536_,
		_w2860_,
		_w3336_
	);
	LUT3 #(
		.INIT('ha2)
	) name2874 (
		\P1_reg1_reg[27]/NET0131 ,
		_w2332_,
		_w2544_,
		_w3337_
	);
	LUT4 #(
		.INIT('h1000)
	) name2875 (
		_w489_,
		_w1040_,
		_w2194_,
		_w2536_,
		_w3338_
	);
	LUT2 #(
		.INIT('h1)
	) name2876 (
		_w3337_,
		_w3338_,
		_w3339_
	);
	LUT4 #(
		.INIT('h5700)
	) name2877 (
		_w2170_,
		_w3331_,
		_w3336_,
		_w3339_,
		_w3340_
	);
	LUT4 #(
		.INIT('h5700)
	) name2878 (
		_w2121_,
		_w3331_,
		_w3335_,
		_w3340_,
		_w3341_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2879 (
		_w2128_,
		_w3332_,
		_w3334_,
		_w3341_,
		_w3342_
	);
	LUT2 #(
		.INIT('h8)
	) name2880 (
		\P1_reg1_reg[27]/NET0131 ,
		_w2183_,
		_w3343_
	);
	LUT4 #(
		.INIT('haa08)
	) name2881 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w3342_,
		_w3343_,
		_w3344_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2882 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[27]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3345_
	);
	LUT2 #(
		.INIT('he)
	) name2883 (
		_w3344_,
		_w3345_,
		_w3346_
	);
	LUT2 #(
		.INIT('h8)
	) name2884 (
		_w853_,
		_w2183_,
		_w3347_
	);
	LUT4 #(
		.INIT('h4044)
	) name2885 (
		_w1167_,
		_w2065_,
		_w2082_,
		_w2085_,
		_w3348_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2886 (
		_w1167_,
		_w2065_,
		_w2082_,
		_w2085_,
		_w3349_
	);
	LUT3 #(
		.INIT('h02)
	) name2887 (
		_w2121_,
		_w3349_,
		_w3348_,
		_w3350_
	);
	LUT4 #(
		.INIT('h0100)
	) name2888 (
		_w856_,
		_w876_,
		_w889_,
		_w2134_,
		_w3351_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2889 (
		_w488_,
		_w873_,
		_w875_,
		_w1237_,
		_w3352_
	);
	LUT4 #(
		.INIT('heb00)
	) name2890 (
		_w488_,
		_w847_,
		_w3351_,
		_w3352_,
		_w3353_
	);
	LUT4 #(
		.INIT('hd200)
	) name2891 (
		_w922_,
		_w1019_,
		_w1167_,
		_w2128_,
		_w3354_
	);
	LUT4 #(
		.INIT('h1555)
	) name2892 (
		_w864_,
		_w2159_,
		_w2160_,
		_w2161_,
		_w3355_
	);
	LUT4 #(
		.INIT('h70f0)
	) name2893 (
		_w2159_,
		_w2160_,
		_w2170_,
		_w2858_,
		_w3356_
	);
	LUT2 #(
		.INIT('h4)
	) name2894 (
		_w3355_,
		_w3356_,
		_w3357_
	);
	LUT3 #(
		.INIT('h01)
	) name2895 (
		_w3353_,
		_w3354_,
		_w3357_,
		_w3358_
	);
	LUT3 #(
		.INIT('h10)
	) name2896 (
		_w864_,
		_w2175_,
		_w2176_,
		_w3359_
	);
	LUT3 #(
		.INIT('h09)
	) name2897 (
		_w1096_,
		_w1098_,
		_w1122_,
		_w3360_
	);
	LUT4 #(
		.INIT('h0054)
	) name2898 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w3360_,
		_w3361_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2899 (
		_w853_,
		_w2171_,
		_w2578_,
		_w3361_,
		_w3362_
	);
	LUT2 #(
		.INIT('h1)
	) name2900 (
		_w3359_,
		_w3362_,
		_w3363_
	);
	LUT4 #(
		.INIT('h7500)
	) name2901 (
		_w2055_,
		_w3350_,
		_w3358_,
		_w3363_,
		_w3364_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2902 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w3347_,
		_w3364_,
		_w3365_
	);
	LUT2 #(
		.INIT('h2)
	) name2903 (
		\P1_reg3_reg[12]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3366_
	);
	LUT4 #(
		.INIT('h4080)
	) name2904 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w853_,
		_w1242_,
		_w3367_
	);
	LUT2 #(
		.INIT('h1)
	) name2905 (
		_w3366_,
		_w3367_,
		_w3368_
	);
	LUT2 #(
		.INIT('hb)
	) name2906 (
		_w3365_,
		_w3368_,
		_w3369_
	);
	LUT2 #(
		.INIT('h8)
	) name2907 (
		_w735_,
		_w2183_,
		_w3370_
	);
	LUT4 #(
		.INIT('h2220)
	) name2908 (
		_w735_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3371_
	);
	LUT4 #(
		.INIT('h8848)
	) name2909 (
		_w1216_,
		_w2055_,
		_w2650_,
		_w2657_,
		_w3372_
	);
	LUT3 #(
		.INIT('ha8)
	) name2910 (
		_w2128_,
		_w3371_,
		_w3372_,
		_w3373_
	);
	LUT3 #(
		.INIT('h8a)
	) name2911 (
		_w2676_,
		_w2682_,
		_w2683_,
		_w3374_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2912 (
		_w2675_,
		_w2676_,
		_w2682_,
		_w2683_,
		_w3375_
	);
	LUT4 #(
		.INIT('h4484)
	) name2913 (
		_w1216_,
		_w2055_,
		_w2677_,
		_w3375_,
		_w3376_
	);
	LUT3 #(
		.INIT('ha8)
	) name2914 (
		_w2121_,
		_w3371_,
		_w3376_,
		_w3377_
	);
	LUT2 #(
		.INIT('h8)
	) name2915 (
		_w488_,
		_w754_,
		_w3378_
	);
	LUT4 #(
		.INIT('h00eb)
	) name2916 (
		_w488_,
		_w724_,
		_w2213_,
		_w3378_,
		_w3379_
	);
	LUT4 #(
		.INIT('hc808)
	) name2917 (
		_w735_,
		_w1237_,
		_w2055_,
		_w3379_,
		_w3380_
	);
	LUT4 #(
		.INIT('h1555)
	) name2918 (
		_w734_,
		_w749_,
		_w759_,
		_w2163_,
		_w3381_
	);
	LUT3 #(
		.INIT('h70)
	) name2919 (
		_w2153_,
		_w2163_,
		_w2170_,
		_w3382_
	);
	LUT3 #(
		.INIT('ha8)
	) name2920 (
		_w735_,
		_w2171_,
		_w2173_,
		_w3383_
	);
	LUT3 #(
		.INIT('h10)
	) name2921 (
		_w734_,
		_w2175_,
		_w2176_,
		_w3384_
	);
	LUT2 #(
		.INIT('h1)
	) name2922 (
		_w3383_,
		_w3384_,
		_w3385_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2923 (
		_w2055_,
		_w3381_,
		_w3382_,
		_w3385_,
		_w3386_
	);
	LUT2 #(
		.INIT('h4)
	) name2924 (
		_w3380_,
		_w3386_,
		_w3387_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2925 (
		_w2182_,
		_w3377_,
		_w3373_,
		_w3387_,
		_w3388_
	);
	LUT2 #(
		.INIT('h2)
	) name2926 (
		\P1_reg3_reg[18]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3389_
	);
	LUT3 #(
		.INIT('h07)
	) name2927 (
		_w735_,
		_w1244_,
		_w3389_,
		_w3390_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2928 (
		\P1_state_reg[0]/NET0131 ,
		_w3370_,
		_w3388_,
		_w3390_,
		_w3391_
	);
	LUT4 #(
		.INIT('h4000)
	) name2929 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1613_,
		_w3392_
	);
	LUT2 #(
		.INIT('h2)
	) name2930 (
		_w1613_,
		_w2903_,
		_w3393_
	);
	LUT4 #(
		.INIT('h1000)
	) name2931 (
		_w1631_,
		_w1812_,
		_w1978_,
		_w1980_,
		_w3394_
	);
	LUT4 #(
		.INIT('h6555)
	) name2932 (
		_w1631_,
		_w1812_,
		_w1978_,
		_w1980_,
		_w3395_
	);
	LUT4 #(
		.INIT('h7020)
	) name2933 (
		_w1305_,
		_w1807_,
		_w2903_,
		_w3395_,
		_w3396_
	);
	LUT3 #(
		.INIT('ha8)
	) name2934 (
		_w2000_,
		_w3393_,
		_w3396_,
		_w3397_
	);
	LUT4 #(
		.INIT('h7500)
	) name2935 (
		_w1878_,
		_w1905_,
		_w1908_,
		_w1916_,
		_w3398_
	);
	LUT4 #(
		.INIT('hc060)
	) name2936 (
		_w1923_,
		_w2508_,
		_w2903_,
		_w3398_,
		_w3399_
	);
	LUT3 #(
		.INIT('ha8)
	) name2937 (
		_w1963_,
		_w3393_,
		_w3399_,
		_w3400_
	);
	LUT4 #(
		.INIT('h006f)
	) name2938 (
		_w2508_,
		_w2880_,
		_w2903_,
		_w3393_,
		_w3401_
	);
	LUT3 #(
		.INIT('h80)
	) name2939 (
		_w2009_,
		_w2010_,
		_w2017_,
		_w3402_
	);
	LUT4 #(
		.INIT('h4000)
	) name2940 (
		_w1612_,
		_w2009_,
		_w2010_,
		_w2017_,
		_w3403_
	);
	LUT4 #(
		.INIT('h9555)
	) name2941 (
		_w1612_,
		_w2009_,
		_w2010_,
		_w2017_,
		_w3404_
	);
	LUT4 #(
		.INIT('hc808)
	) name2942 (
		_w1613_,
		_w2025_,
		_w2903_,
		_w3404_,
		_w3405_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name2943 (
		_w1612_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w3406_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2944 (
		_w1613_,
		_w2001_,
		_w2032_,
		_w2903_,
		_w3407_
	);
	LUT2 #(
		.INIT('h1)
	) name2945 (
		_w3406_,
		_w3407_,
		_w3408_
	);
	LUT2 #(
		.INIT('h4)
	) name2946 (
		_w3405_,
		_w3408_,
		_w3409_
	);
	LUT3 #(
		.INIT('hd0)
	) name2947 (
		_w1869_,
		_w3401_,
		_w3409_,
		_w3410_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2948 (
		_w1285_,
		_w3397_,
		_w3400_,
		_w3410_,
		_w3411_
	);
	LUT2 #(
		.INIT('h4)
	) name2949 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[17]/NET0131 ,
		_w3412_
	);
	LUT3 #(
		.INIT('h07)
	) name2950 (
		_w1613_,
		_w2344_,
		_w3412_,
		_w3413_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2951 (
		\P1_state_reg[0]/NET0131 ,
		_w3392_,
		_w3411_,
		_w3413_,
		_w3414_
	);
	LUT4 #(
		.INIT('h4000)
	) name2952 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1627_,
		_w3415_
	);
	LUT2 #(
		.INIT('h2)
	) name2953 (
		_w1627_,
		_w2903_,
		_w3416_
	);
	LUT4 #(
		.INIT('h0200)
	) name2954 (
		_w1305_,
		_w1615_,
		_w1614_,
		_w1616_,
		_w3417_
	);
	LUT4 #(
		.INIT('h00eb)
	) name2955 (
		_w1305_,
		_w1604_,
		_w3394_,
		_w3417_,
		_w3418_
	);
	LUT4 #(
		.INIT('hc808)
	) name2956 (
		_w1627_,
		_w2000_,
		_w2903_,
		_w3418_,
		_w3419_
	);
	LUT4 #(
		.INIT('h4844)
	) name2957 (
		_w2511_,
		_w2903_,
		_w3099_,
		_w3100_,
		_w3420_
	);
	LUT3 #(
		.INIT('ha8)
	) name2958 (
		_w1869_,
		_w3416_,
		_w3420_,
		_w3421_
	);
	LUT4 #(
		.INIT('h8488)
	) name2959 (
		_w2511_,
		_w2903_,
		_w3113_,
		_w3116_,
		_w3422_
	);
	LUT4 #(
		.INIT('h8040)
	) name2960 (
		_w1626_,
		_w2025_,
		_w2903_,
		_w3403_,
		_w3423_
	);
	LUT4 #(
		.INIT('h88a8)
	) name2961 (
		_w1627_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w3424_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name2962 (
		_w1626_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w3425_
	);
	LUT2 #(
		.INIT('h1)
	) name2963 (
		_w3424_,
		_w3425_,
		_w3426_
	);
	LUT2 #(
		.INIT('h4)
	) name2964 (
		_w3423_,
		_w3426_,
		_w3427_
	);
	LUT4 #(
		.INIT('h5700)
	) name2965 (
		_w1963_,
		_w3416_,
		_w3422_,
		_w3427_,
		_w3428_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2966 (
		_w1285_,
		_w3419_,
		_w3421_,
		_w3428_,
		_w3429_
	);
	LUT2 #(
		.INIT('h4)
	) name2967 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		_w3430_
	);
	LUT3 #(
		.INIT('h07)
	) name2968 (
		_w1627_,
		_w2344_,
		_w3430_,
		_w3431_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2969 (
		\P1_state_reg[0]/NET0131 ,
		_w3415_,
		_w3429_,
		_w3431_,
		_w3432_
	);
	LUT4 #(
		.INIT('h4000)
	) name2970 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1600_,
		_w3433_
	);
	LUT4 #(
		.INIT('h6050)
	) name2971 (
		_w1599_,
		_w1626_,
		_w2025_,
		_w3403_,
		_w3434_
	);
	LUT4 #(
		.INIT('h8288)
	) name2972 (
		_w1963_,
		_w2504_,
		_w2597_,
		_w2598_,
		_w3435_
	);
	LUT3 #(
		.INIT('h82)
	) name2973 (
		_w1869_,
		_w2504_,
		_w2622_,
		_w3436_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2974 (
		_w2903_,
		_w3435_,
		_w3436_,
		_w3434_,
		_w3437_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2975 (
		_w1305_,
		_w1629_,
		_w1628_,
		_w1630_,
		_w3438_
	);
	LUT3 #(
		.INIT('h15)
	) name2976 (
		_w1305_,
		_w1978_,
		_w1982_,
		_w3439_
	);
	LUT4 #(
		.INIT('h7500)
	) name2977 (
		_w1592_,
		_w1604_,
		_w3394_,
		_w3439_,
		_w3440_
	);
	LUT3 #(
		.INIT('hc8)
	) name2978 (
		_w1600_,
		_w2000_,
		_w2903_,
		_w3441_
	);
	LUT4 #(
		.INIT('hfd00)
	) name2979 (
		_w2903_,
		_w3438_,
		_w3440_,
		_w3441_,
		_w3442_
	);
	LUT4 #(
		.INIT('hcc03)
	) name2980 (
		_w1595_,
		_w1863_,
		_w1864_,
		_w1866_,
		_w3443_
	);
	LUT4 #(
		.INIT('h5150)
	) name2981 (
		_w2032_,
		_w2033_,
		_w2903_,
		_w3443_,
		_w3444_
	);
	LUT4 #(
		.INIT('hf531)
	) name2982 (
		_w1599_,
		_w1600_,
		_w2993_,
		_w3444_,
		_w3445_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2983 (
		_w1285_,
		_w3442_,
		_w3437_,
		_w3445_,
		_w3446_
	);
	LUT2 #(
		.INIT('h4)
	) name2984 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[19]/NET0131 ,
		_w3447_
	);
	LUT3 #(
		.INIT('h07)
	) name2985 (
		_w1600_,
		_w2344_,
		_w3447_,
		_w3448_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2986 (
		\P1_state_reg[0]/NET0131 ,
		_w3433_,
		_w3446_,
		_w3448_,
		_w3449_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2987 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[17]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3450_
	);
	LUT2 #(
		.INIT('h8)
	) name2988 (
		\P1_reg2_reg[17]/NET0131 ,
		_w2183_,
		_w3451_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2989 (
		\P1_reg2_reg[17]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3452_
	);
	LUT4 #(
		.INIT('h0075)
	) name2990 (
		_w739_,
		_w754_,
		_w2139_,
		_w2213_,
		_w3453_
	);
	LUT4 #(
		.INIT('h7020)
	) name2991 (
		_w488_,
		_w764_,
		_w2189_,
		_w3453_,
		_w3454_
	);
	LUT3 #(
		.INIT('ha8)
	) name2992 (
		_w1237_,
		_w3452_,
		_w3454_,
		_w3455_
	);
	LUT4 #(
		.INIT('h59aa)
	) name2993 (
		_w1225_,
		_w2223_,
		_w2243_,
		_w2246_,
		_w3456_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2994 (
		\P1_reg2_reg[17]/NET0131 ,
		_w2128_,
		_w2189_,
		_w3456_,
		_w3457_
	);
	LUT4 #(
		.INIT('h8488)
	) name2995 (
		_w1225_,
		_w2189_,
		_w2703_,
		_w2704_,
		_w3458_
	);
	LUT4 #(
		.INIT('h6a00)
	) name2996 (
		_w749_,
		_w759_,
		_w2163_,
		_w2189_,
		_w3459_
	);
	LUT2 #(
		.INIT('h4)
	) name2997 (
		_w749_,
		_w2194_,
		_w3460_
	);
	LUT3 #(
		.INIT('h40)
	) name2998 (
		_w749_,
		_w2189_,
		_w2194_,
		_w3461_
	);
	LUT2 #(
		.INIT('h8)
	) name2999 (
		_w751_,
		_w1120_,
		_w3462_
	);
	LUT4 #(
		.INIT('h0057)
	) name3000 (
		\P1_reg2_reg[17]/NET0131 ,
		_w2171_,
		_w2196_,
		_w3462_,
		_w3463_
	);
	LUT2 #(
		.INIT('h4)
	) name3001 (
		_w3461_,
		_w3463_,
		_w3464_
	);
	LUT4 #(
		.INIT('h5700)
	) name3002 (
		_w2170_,
		_w3452_,
		_w3459_,
		_w3464_,
		_w3465_
	);
	LUT4 #(
		.INIT('h5700)
	) name3003 (
		_w2121_,
		_w3452_,
		_w3458_,
		_w3465_,
		_w3466_
	);
	LUT2 #(
		.INIT('h4)
	) name3004 (
		_w3457_,
		_w3466_,
		_w3467_
	);
	LUT4 #(
		.INIT('h1311)
	) name3005 (
		_w2182_,
		_w3451_,
		_w3455_,
		_w3467_,
		_w3468_
	);
	LUT3 #(
		.INIT('hce)
	) name3006 (
		\P1_state_reg[0]/NET0131 ,
		_w3450_,
		_w3468_,
		_w3469_
	);
	LUT2 #(
		.INIT('h8)
	) name3007 (
		_w806_,
		_w2183_,
		_w3470_
	);
	LUT4 #(
		.INIT('h2220)
	) name3008 (
		_w806_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3471_
	);
	LUT4 #(
		.INIT('h4844)
	) name3009 (
		_w1228_,
		_w2055_,
		_w2093_,
		_w2102_,
		_w3472_
	);
	LUT3 #(
		.INIT('ha8)
	) name3010 (
		_w2121_,
		_w3471_,
		_w3472_,
		_w3473_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3011 (
		_w2055_,
		_w3163_,
		_w3164_,
		_w3471_,
		_w3474_
	);
	LUT2 #(
		.INIT('h2)
	) name3012 (
		_w1237_,
		_w3474_,
		_w3475_
	);
	LUT4 #(
		.INIT('h00b7)
	) name3013 (
		_w1228_,
		_w2055_,
		_w2124_,
		_w3471_,
		_w3476_
	);
	LUT4 #(
		.INIT('h8040)
	) name3014 (
		_w805_,
		_w2055_,
		_w2170_,
		_w3168_,
		_w3477_
	);
	LUT3 #(
		.INIT('ha8)
	) name3015 (
		_w806_,
		_w2171_,
		_w2173_,
		_w3478_
	);
	LUT4 #(
		.INIT('h0100)
	) name3016 (
		_w489_,
		_w804_,
		_w2175_,
		_w2176_,
		_w3479_
	);
	LUT2 #(
		.INIT('h1)
	) name3017 (
		_w3478_,
		_w3479_,
		_w3480_
	);
	LUT2 #(
		.INIT('h4)
	) name3018 (
		_w3477_,
		_w3480_,
		_w3481_
	);
	LUT3 #(
		.INIT('hd0)
	) name3019 (
		_w2128_,
		_w3476_,
		_w3481_,
		_w3482_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3020 (
		_w2182_,
		_w3475_,
		_w3473_,
		_w3482_,
		_w3483_
	);
	LUT4 #(
		.INIT('h95dd)
	) name3021 (
		\P1_reg3_reg[20]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w593_,
		_w1243_,
		_w3484_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3022 (
		\P1_state_reg[0]/NET0131 ,
		_w3470_,
		_w3483_,
		_w3484_,
		_w3485_
	);
	LUT2 #(
		.INIT('h2)
	) name3023 (
		\P2_reg0_reg[22]/NET0131 ,
		_w2042_,
		_w3486_
	);
	LUT4 #(
		.INIT('h2000)
	) name3024 (
		\P2_reg0_reg[22]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3487_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3025 (
		_w3099_,
		_w3100_,
		_w3101_,
		_w3104_,
		_w3488_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3026 (
		\P2_reg0_reg[22]/NET0131 ,
		_w2507_,
		_w2729_,
		_w3488_,
		_w3489_
	);
	LUT2 #(
		.INIT('h2)
	) name3027 (
		_w1869_,
		_w3489_,
		_w3490_
	);
	LUT4 #(
		.INIT('hce00)
	) name3028 (
		_w2414_,
		_w2400_,
		_w2413_,
		_w3111_,
		_w3491_
	);
	LUT2 #(
		.INIT('h8)
	) name3029 (
		_w3110_,
		_w3118_,
		_w3492_
	);
	LUT2 #(
		.INIT('h4)
	) name3030 (
		_w3114_,
		_w3118_,
		_w3493_
	);
	LUT2 #(
		.INIT('h2)
	) name3031 (
		_w3120_,
		_w3493_,
		_w3494_
	);
	LUT4 #(
		.INIT('h2f00)
	) name3032 (
		_w3115_,
		_w3491_,
		_w3492_,
		_w3494_,
		_w3495_
	);
	LUT4 #(
		.INIT('hc535)
	) name3033 (
		\P2_reg0_reg[22]/NET0131 ,
		_w2507_,
		_w2729_,
		_w3495_,
		_w3496_
	);
	LUT2 #(
		.INIT('h2)
	) name3034 (
		_w1305_,
		_w1573_,
		_w3497_
	);
	LUT2 #(
		.INIT('h8)
	) name3035 (
		_w1978_,
		_w1985_,
		_w3498_
	);
	LUT2 #(
		.INIT('h1)
	) name3036 (
		_w1305_,
		_w1551_,
		_w3499_
	);
	LUT4 #(
		.INIT('h00bf)
	) name3037 (
		_w1564_,
		_w1978_,
		_w1983_,
		_w3499_,
		_w3500_
	);
	LUT4 #(
		.INIT('h888a)
	) name3038 (
		_w2000_,
		_w3497_,
		_w3498_,
		_w3500_,
		_w3501_
	);
	LUT4 #(
		.INIT('h5400)
	) name3039 (
		_w1306_,
		_w1555_,
		_w1559_,
		_w2001_,
		_w3502_
	);
	LUT4 #(
		.INIT('h8000)
	) name3040 (
		_w2009_,
		_w2010_,
		_w2013_,
		_w2017_,
		_w3503_
	);
	LUT4 #(
		.INIT('h070b)
	) name3041 (
		_w1560_,
		_w2025_,
		_w3502_,
		_w3503_,
		_w3504_
	);
	LUT2 #(
		.INIT('h4)
	) name3042 (
		_w3501_,
		_w3504_,
		_w3505_
	);
	LUT3 #(
		.INIT('h8a)
	) name3043 (
		\P2_reg0_reg[22]/NET0131 ,
		_w2736_,
		_w3084_,
		_w3506_
	);
	LUT4 #(
		.INIT('h0075)
	) name3044 (
		_w2729_,
		_w3501_,
		_w3504_,
		_w3506_,
		_w3507_
	);
	LUT3 #(
		.INIT('hd0)
	) name3045 (
		_w1963_,
		_w3496_,
		_w3507_,
		_w3508_
	);
	LUT4 #(
		.INIT('h1311)
	) name3046 (
		_w1285_,
		_w3487_,
		_w3490_,
		_w3508_,
		_w3509_
	);
	LUT3 #(
		.INIT('hce)
	) name3047 (
		\P1_state_reg[0]/NET0131 ,
		_w3486_,
		_w3509_,
		_w3510_
	);
	LUT4 #(
		.INIT('hbf00)
	) name3048 (
		_w1249_,
		_w1251_,
		_w1248_,
		_w2205_,
		_w3511_
	);
	LUT3 #(
		.INIT('h70)
	) name3049 (
		_w2119_,
		_w2866_,
		_w3511_,
		_w3512_
	);
	LUT3 #(
		.INIT('h2a)
	) name3050 (
		\P1_reg2_reg[16]/NET0131 ,
		_w3175_,
		_w3512_,
		_w3513_
	);
	LUT4 #(
		.INIT('h1000)
	) name3051 (
		_w1096_,
		_w1098_,
		_w760_,
		_w1101_,
		_w3514_
	);
	LUT4 #(
		.INIT('ha060)
	) name3052 (
		_w1198_,
		_w2096_,
		_w2121_,
		_w2836_,
		_w3515_
	);
	LUT2 #(
		.INIT('h8)
	) name3053 (
		_w1237_,
		_w2840_,
		_w3516_
	);
	LUT4 #(
		.INIT('hf100)
	) name3054 (
		_w489_,
		_w756_,
		_w758_,
		_w2194_,
		_w3517_
	);
	LUT4 #(
		.INIT('h0002)
	) name3055 (
		_w2843_,
		_w3517_,
		_w3515_,
		_w3516_,
		_w3518_
	);
	LUT4 #(
		.INIT('hc0c8)
	) name3056 (
		_w2189_,
		_w3511_,
		_w3514_,
		_w3518_,
		_w3519_
	);
	LUT2 #(
		.INIT('he)
	) name3057 (
		_w3513_,
		_w3519_,
		_w3520_
	);
	LUT2 #(
		.INIT('h2)
	) name3058 (
		\P2_reg0_reg[24]/NET0131 ,
		_w2042_,
		_w3521_
	);
	LUT4 #(
		.INIT('h2000)
	) name3059 (
		\P2_reg0_reg[24]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3522_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3060 (
		\P2_reg0_reg[24]/NET0131 ,
		_w1869_,
		_w2729_,
		_w3214_,
		_w3523_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3061 (
		\P2_reg0_reg[24]/NET0131 ,
		_w1963_,
		_w2729_,
		_w3218_,
		_w3524_
	);
	LUT3 #(
		.INIT('h8a)
	) name3062 (
		\P2_reg0_reg[24]/NET0131 ,
		_w2736_,
		_w3084_,
		_w3525_
	);
	LUT3 #(
		.INIT('h0d)
	) name3063 (
		_w2729_,
		_w3224_,
		_w3525_,
		_w3526_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3064 (
		_w1285_,
		_w3524_,
		_w3523_,
		_w3526_,
		_w3527_
	);
	LUT4 #(
		.INIT('heeec)
	) name3065 (
		\P1_state_reg[0]/NET0131 ,
		_w3521_,
		_w3522_,
		_w3527_,
		_w3528_
	);
	LUT2 #(
		.INIT('h2)
	) name3066 (
		\P2_reg1_reg[25]/NET0131 ,
		_w2042_,
		_w3529_
	);
	LUT4 #(
		.INIT('h2000)
	) name3067 (
		\P2_reg1_reg[25]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3530_
	);
	LUT4 #(
		.INIT('hc535)
	) name3068 (
		\P2_reg1_reg[25]/NET0131 ,
		_w2519_,
		_w2762_,
		_w2878_,
		_w3531_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3069 (
		\P2_reg1_reg[25]/NET0131 ,
		_w1869_,
		_w2762_,
		_w2884_,
		_w3532_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3070 (
		\P2_reg1_reg[25]/NET0131 ,
		_w2762_,
		_w2886_,
		_w2887_,
		_w3533_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3071 (
		\P2_reg1_reg[25]/NET0131 ,
		_w2033_,
		_w2734_,
		_w2762_,
		_w3534_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3072 (
		_w2762_,
		_w2889_,
		_w2891_,
		_w2892_,
		_w3535_
	);
	LUT4 #(
		.INIT('h0031)
	) name3073 (
		_w2000_,
		_w3534_,
		_w3533_,
		_w3535_,
		_w3536_
	);
	LUT4 #(
		.INIT('h3100)
	) name3074 (
		_w1963_,
		_w3532_,
		_w3531_,
		_w3536_,
		_w3537_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3075 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w3530_,
		_w3537_,
		_w3538_
	);
	LUT2 #(
		.INIT('he)
	) name3076 (
		_w3529_,
		_w3538_,
		_w3539_
	);
	LUT2 #(
		.INIT('h2)
	) name3077 (
		\P2_reg2_reg[24]/NET0131 ,
		_w2042_,
		_w3540_
	);
	LUT4 #(
		.INIT('h2000)
	) name3078 (
		\P2_reg2_reg[24]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3541_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3079 (
		\P2_reg2_reg[24]/NET0131 ,
		_w1298_,
		_w1869_,
		_w3214_,
		_w3542_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3080 (
		\P2_reg2_reg[24]/NET0131 ,
		_w1298_,
		_w1963_,
		_w3218_,
		_w3543_
	);
	LUT4 #(
		.INIT('h3200)
	) name3081 (
		\P2_reg3_reg[24]/NET0131 ,
		_w1394_,
		_w1536_,
		_w2029_,
		_w3544_
	);
	LUT4 #(
		.INIT('h0075)
	) name3082 (
		\P2_reg2_reg[24]/NET0131 ,
		_w2031_,
		_w2640_,
		_w3544_,
		_w3545_
	);
	LUT3 #(
		.INIT('hd0)
	) name3083 (
		_w1298_,
		_w3224_,
		_w3545_,
		_w3546_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3084 (
		_w1285_,
		_w3543_,
		_w3542_,
		_w3546_,
		_w3547_
	);
	LUT4 #(
		.INIT('heeec)
	) name3085 (
		\P1_state_reg[0]/NET0131 ,
		_w3540_,
		_w3541_,
		_w3547_,
		_w3548_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3086 (
		\P2_reg2_reg[26]/NET0131 ,
		_w1298_,
		_w2514_,
		_w3107_,
		_w3549_
	);
	LUT2 #(
		.INIT('h2)
	) name3087 (
		_w1869_,
		_w3549_,
		_w3550_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3088 (
		\P2_reg2_reg[26]/NET0131 ,
		_w1298_,
		_w2514_,
		_w3123_,
		_w3551_
	);
	LUT2 #(
		.INIT('h8)
	) name3089 (
		_w1507_,
		_w2029_,
		_w3552_
	);
	LUT4 #(
		.INIT('h0075)
	) name3090 (
		\P2_reg2_reg[26]/NET0131 ,
		_w2031_,
		_w2640_,
		_w3552_,
		_w3553_
	);
	LUT4 #(
		.INIT('h7500)
	) name3091 (
		_w1298_,
		_w3126_,
		_w3128_,
		_w3553_,
		_w3554_
	);
	LUT3 #(
		.INIT('hd0)
	) name3092 (
		_w1963_,
		_w3551_,
		_w3554_,
		_w3555_
	);
	LUT4 #(
		.INIT('h2000)
	) name3093 (
		\P2_reg2_reg[26]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3556_
	);
	LUT4 #(
		.INIT('h0075)
	) name3094 (
		_w1285_,
		_w3550_,
		_w3555_,
		_w3556_,
		_w3557_
	);
	LUT2 #(
		.INIT('h2)
	) name3095 (
		\P2_reg2_reg[26]/NET0131 ,
		_w2042_,
		_w3558_
	);
	LUT3 #(
		.INIT('hf2)
	) name3096 (
		\P1_state_reg[0]/NET0131 ,
		_w3557_,
		_w3558_,
		_w3559_
	);
	LUT4 #(
		.INIT('hbf00)
	) name3097 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2172_,
		_w3560_
	);
	LUT4 #(
		.INIT('h0002)
	) name3098 (
		_w2332_,
		_w2798_,
		_w3295_,
		_w3560_,
		_w3561_
	);
	LUT3 #(
		.INIT('h2a)
	) name3099 (
		\P1_reg0_reg[16]/NET0131 ,
		_w3511_,
		_w3561_,
		_w3562_
	);
	LUT4 #(
		.INIT('h4000)
	) name3100 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w3511_,
		_w3563_
	);
	LUT3 #(
		.INIT('hdc)
	) name3101 (
		_w3518_,
		_w3562_,
		_w3563_,
		_w3564_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name3102 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[21]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3565_
	);
	LUT2 #(
		.INIT('h8)
	) name3103 (
		\P1_reg0_reg[21]/NET0131 ,
		_w2183_,
		_w3566_
	);
	LUT4 #(
		.INIT('h00bf)
	) name3104 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w3360_,
		_w3567_
	);
	LUT4 #(
		.INIT('haaa2)
	) name3105 (
		\P1_reg0_reg[21]/NET0131 ,
		_w2332_,
		_w2333_,
		_w3567_,
		_w3568_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3106 (
		_w780_,
		_w800_,
		_w2140_,
		_w2213_,
		_w3569_
	);
	LUT2 #(
		.INIT('h8)
	) name3107 (
		_w2141_,
		_w2213_,
		_w3570_
	);
	LUT4 #(
		.INIT('h0200)
	) name3108 (
		_w488_,
		_w808_,
		_w807_,
		_w809_,
		_w3571_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3109 (
		_w488_,
		_w3569_,
		_w3570_,
		_w3571_,
		_w3572_
	);
	LUT2 #(
		.INIT('h8)
	) name3110 (
		_w1237_,
		_w3572_,
		_w3573_
	);
	LUT3 #(
		.INIT('h84)
	) name3111 (
		_w796_,
		_w2170_,
		_w3169_,
		_w3574_
	);
	LUT4 #(
		.INIT('h5400)
	) name3112 (
		_w489_,
		_w793_,
		_w795_,
		_w2194_,
		_w3575_
	);
	LUT3 #(
		.INIT('h84)
	) name3113 (
		_w1204_,
		_w2121_,
		_w2298_,
		_w3576_
	);
	LUT4 #(
		.INIT('h0455)
	) name3114 (
		_w1204_,
		_w2224_,
		_w2243_,
		_w2251_,
		_w3577_
	);
	LUT4 #(
		.INIT('ha200)
	) name3115 (
		_w1204_,
		_w2224_,
		_w2243_,
		_w2251_,
		_w3578_
	);
	LUT3 #(
		.INIT('h02)
	) name3116 (
		_w2128_,
		_w3578_,
		_w3577_,
		_w3579_
	);
	LUT3 #(
		.INIT('h01)
	) name3117 (
		_w3575_,
		_w3576_,
		_w3579_,
		_w3580_
	);
	LUT4 #(
		.INIT('h0001)
	) name3118 (
		_w3574_,
		_w3575_,
		_w3576_,
		_w3579_,
		_w3581_
	);
	LUT4 #(
		.INIT('h1311)
	) name3119 (
		_w2325_,
		_w3568_,
		_w3573_,
		_w3581_,
		_w3582_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3120 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w3566_,
		_w3582_,
		_w3583_
	);
	LUT2 #(
		.INIT('he)
	) name3121 (
		_w3565_,
		_w3583_,
		_w3584_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name3122 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[24]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3585_
	);
	LUT2 #(
		.INIT('h8)
	) name3123 (
		\P1_reg0_reg[24]/NET0131 ,
		_w2183_,
		_w3586_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3124 (
		\P1_reg0_reg[24]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3587_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3125 (
		\P1_reg0_reg[24]/NET0131 ,
		_w1210_,
		_w2325_,
		_w2565_,
		_w3588_
	);
	LUT4 #(
		.INIT('h7020)
	) name3126 (
		_w488_,
		_w789_,
		_w2325_,
		_w2567_,
		_w3589_
	);
	LUT3 #(
		.INIT('ha8)
	) name3127 (
		_w1237_,
		_w3587_,
		_w3589_,
		_w3590_
	);
	LUT4 #(
		.INIT('h8488)
	) name3128 (
		_w1210_,
		_w2325_,
		_w2571_,
		_w2572_,
		_w3591_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3129 (
		\P1_reg0_reg[24]/NET0131 ,
		_w2325_,
		_w2574_,
		_w2575_,
		_w3592_
	);
	LUT3 #(
		.INIT('ha2)
	) name3130 (
		\P1_reg0_reg[24]/NET0131 ,
		_w2332_,
		_w2333_,
		_w3593_
	);
	LUT2 #(
		.INIT('h8)
	) name3131 (
		_w2325_,
		_w2752_,
		_w3594_
	);
	LUT2 #(
		.INIT('h1)
	) name3132 (
		_w3593_,
		_w3594_,
		_w3595_
	);
	LUT3 #(
		.INIT('hd0)
	) name3133 (
		_w2170_,
		_w3592_,
		_w3595_,
		_w3596_
	);
	LUT4 #(
		.INIT('h5700)
	) name3134 (
		_w2128_,
		_w3587_,
		_w3591_,
		_w3596_,
		_w3597_
	);
	LUT4 #(
		.INIT('h3100)
	) name3135 (
		_w2121_,
		_w3590_,
		_w3588_,
		_w3597_,
		_w3598_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3136 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w3586_,
		_w3598_,
		_w3599_
	);
	LUT2 #(
		.INIT('he)
	) name3137 (
		_w3585_,
		_w3599_,
		_w3600_
	);
	LUT2 #(
		.INIT('h8)
	) name3138 (
		_w2170_,
		_w2863_,
		_w3601_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name3139 (
		_w2855_,
		_w2857_,
		_w3563_,
		_w3601_,
		_w3602_
	);
	LUT3 #(
		.INIT('h2a)
	) name3140 (
		\P1_reg0_reg[31]/NET0131 ,
		_w2332_,
		_w3563_,
		_w3603_
	);
	LUT2 #(
		.INIT('he)
	) name3141 (
		_w3602_,
		_w3603_,
		_w3604_
	);
	LUT4 #(
		.INIT('hef00)
	) name3142 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2128_,
		_w3605_
	);
	LUT4 #(
		.INIT('h0002)
	) name3143 (
		_w2332_,
		_w2544_,
		_w2817_,
		_w3605_,
		_w3606_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3144 (
		\P1_reg1_reg[16]/NET0131 ,
		_w2820_,
		_w3511_,
		_w3606_,
		_w3607_
	);
	LUT4 #(
		.INIT('h1000)
	) name3145 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w3511_,
		_w3608_
	);
	LUT3 #(
		.INIT('hdc)
	) name3146 (
		_w3518_,
		_w3607_,
		_w3608_,
		_w3609_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name3147 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[17]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3610_
	);
	LUT2 #(
		.INIT('h8)
	) name3148 (
		\P1_reg1_reg[17]/NET0131 ,
		_w2183_,
		_w3611_
	);
	LUT4 #(
		.INIT('h7020)
	) name3149 (
		_w488_,
		_w764_,
		_w1237_,
		_w3453_,
		_w3612_
	);
	LUT2 #(
		.INIT('h2)
	) name3150 (
		_w2128_,
		_w3456_,
		_w3613_
	);
	LUT4 #(
		.INIT('h6a00)
	) name3151 (
		_w749_,
		_w759_,
		_w2163_,
		_w2170_,
		_w3614_
	);
	LUT4 #(
		.INIT('h8488)
	) name3152 (
		_w1225_,
		_w2121_,
		_w2703_,
		_w2704_,
		_w3615_
	);
	LUT3 #(
		.INIT('h01)
	) name3153 (
		_w3460_,
		_w3615_,
		_w3614_,
		_w3616_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3154 (
		_w2536_,
		_w3612_,
		_w3613_,
		_w3616_,
		_w3617_
	);
	LUT3 #(
		.INIT('h8a)
	) name3155 (
		\P1_reg1_reg[17]/NET0131 ,
		_w2820_,
		_w3606_,
		_w3618_
	);
	LUT4 #(
		.INIT('h1113)
	) name3156 (
		_w2182_,
		_w3611_,
		_w3617_,
		_w3618_,
		_w3619_
	);
	LUT3 #(
		.INIT('hce)
	) name3157 (
		\P1_state_reg[0]/NET0131 ,
		_w3610_,
		_w3619_,
		_w3620_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name3158 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[21]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3621_
	);
	LUT2 #(
		.INIT('h8)
	) name3159 (
		\P1_reg1_reg[21]/NET0131 ,
		_w2183_,
		_w3622_
	);
	LUT4 #(
		.INIT('h5455)
	) name3160 (
		\P1_reg1_reg[21]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3623_
	);
	LUT2 #(
		.INIT('h2)
	) name3161 (
		_w1237_,
		_w3623_,
		_w3624_
	);
	LUT3 #(
		.INIT('hd0)
	) name3162 (
		_w2536_,
		_w3572_,
		_w3624_,
		_w3625_
	);
	LUT4 #(
		.INIT('hef00)
	) name3163 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2120_,
		_w3626_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3164 (
		_w1123_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3627_
	);
	LUT4 #(
		.INIT('h0002)
	) name3165 (
		_w2332_,
		_w2544_,
		_w3626_,
		_w3627_,
		_w3628_
	);
	LUT2 #(
		.INIT('h2)
	) name3166 (
		\P1_reg1_reg[21]/NET0131 ,
		_w3628_,
		_w3629_
	);
	LUT4 #(
		.INIT('h000d)
	) name3167 (
		_w2536_,
		_w3581_,
		_w3625_,
		_w3629_,
		_w3630_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3168 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w3622_,
		_w3630_,
		_w3631_
	);
	LUT2 #(
		.INIT('he)
	) name3169 (
		_w3621_,
		_w3631_,
		_w3632_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name3170 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[24]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3633_
	);
	LUT2 #(
		.INIT('h8)
	) name3171 (
		\P1_reg1_reg[24]/NET0131 ,
		_w2183_,
		_w3634_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3172 (
		\P1_reg1_reg[24]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3635_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3173 (
		\P1_reg1_reg[24]/NET0131 ,
		_w1210_,
		_w2536_,
		_w2565_,
		_w3636_
	);
	LUT4 #(
		.INIT('h7020)
	) name3174 (
		_w488_,
		_w789_,
		_w2536_,
		_w2567_,
		_w3637_
	);
	LUT3 #(
		.INIT('ha8)
	) name3175 (
		_w1237_,
		_w3635_,
		_w3637_,
		_w3638_
	);
	LUT4 #(
		.INIT('h8488)
	) name3176 (
		_w1210_,
		_w2536_,
		_w2571_,
		_w2572_,
		_w3639_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3177 (
		\P1_reg1_reg[24]/NET0131 ,
		_w2536_,
		_w2574_,
		_w2575_,
		_w3640_
	);
	LUT2 #(
		.INIT('h8)
	) name3178 (
		_w2536_,
		_w2752_,
		_w3641_
	);
	LUT3 #(
		.INIT('ha2)
	) name3179 (
		\P1_reg1_reg[24]/NET0131 ,
		_w2332_,
		_w2544_,
		_w3642_
	);
	LUT2 #(
		.INIT('h1)
	) name3180 (
		_w3641_,
		_w3642_,
		_w3643_
	);
	LUT3 #(
		.INIT('hd0)
	) name3181 (
		_w2170_,
		_w3640_,
		_w3643_,
		_w3644_
	);
	LUT4 #(
		.INIT('h5700)
	) name3182 (
		_w2128_,
		_w3635_,
		_w3639_,
		_w3644_,
		_w3645_
	);
	LUT4 #(
		.INIT('h3100)
	) name3183 (
		_w2121_,
		_w3638_,
		_w3636_,
		_w3645_,
		_w3646_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3184 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w3634_,
		_w3646_,
		_w3647_
	);
	LUT2 #(
		.INIT('he)
	) name3185 (
		_w3633_,
		_w3647_,
		_w3648_
	);
	LUT4 #(
		.INIT('hfe00)
	) name3186 (
		_w2855_,
		_w2857_,
		_w3601_,
		_w3608_,
		_w3649_
	);
	LUT3 #(
		.INIT('h2a)
	) name3187 (
		\P1_reg1_reg[31]/NET0131 ,
		_w2332_,
		_w3608_,
		_w3650_
	);
	LUT2 #(
		.INIT('he)
	) name3188 (
		_w3649_,
		_w3650_,
		_w3651_
	);
	LUT2 #(
		.INIT('h8)
	) name3189 (
		_w751_,
		_w2183_,
		_w3652_
	);
	LUT4 #(
		.INIT('h2220)
	) name3190 (
		_w751_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3653_
	);
	LUT4 #(
		.INIT('h7020)
	) name3191 (
		_w488_,
		_w764_,
		_w2055_,
		_w3453_,
		_w3654_
	);
	LUT3 #(
		.INIT('ha8)
	) name3192 (
		_w1237_,
		_w3653_,
		_w3654_,
		_w3655_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3193 (
		_w751_,
		_w2055_,
		_w2128_,
		_w3456_,
		_w3656_
	);
	LUT4 #(
		.INIT('h8488)
	) name3194 (
		_w1225_,
		_w2055_,
		_w2703_,
		_w2704_,
		_w3657_
	);
	LUT3 #(
		.INIT('ha8)
	) name3195 (
		_w751_,
		_w2171_,
		_w2173_,
		_w3658_
	);
	LUT3 #(
		.INIT('h10)
	) name3196 (
		_w749_,
		_w2175_,
		_w2176_,
		_w3659_
	);
	LUT2 #(
		.INIT('h1)
	) name3197 (
		_w3658_,
		_w3659_,
		_w3660_
	);
	LUT3 #(
		.INIT('h70)
	) name3198 (
		_w2055_,
		_w3614_,
		_w3660_,
		_w3661_
	);
	LUT4 #(
		.INIT('h5700)
	) name3199 (
		_w2121_,
		_w3653_,
		_w3657_,
		_w3661_,
		_w3662_
	);
	LUT2 #(
		.INIT('h4)
	) name3200 (
		_w3656_,
		_w3662_,
		_w3663_
	);
	LUT4 #(
		.INIT('h1311)
	) name3201 (
		_w2182_,
		_w3652_,
		_w3655_,
		_w3663_,
		_w3664_
	);
	LUT4 #(
		.INIT('h3200)
	) name3202 (
		\P1_reg3_reg[17]/NET0131 ,
		_w591_,
		_w750_,
		_w1244_,
		_w3665_
	);
	LUT2 #(
		.INIT('h2)
	) name3203 (
		\P1_reg3_reg[17]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3666_
	);
	LUT2 #(
		.INIT('h1)
	) name3204 (
		_w3665_,
		_w3666_,
		_w3667_
	);
	LUT3 #(
		.INIT('h2f)
	) name3205 (
		\P1_state_reg[0]/NET0131 ,
		_w3664_,
		_w3667_,
		_w3668_
	);
	LUT2 #(
		.INIT('h8)
	) name3206 (
		_w721_,
		_w2183_,
		_w3669_
	);
	LUT4 #(
		.INIT('h2220)
	) name3207 (
		_w721_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3670_
	);
	LUT4 #(
		.INIT('h4150)
	) name3208 (
		_w488_,
		_w724_,
		_w810_,
		_w2213_,
		_w3671_
	);
	LUT4 #(
		.INIT('h0200)
	) name3209 (
		_w488_,
		_w737_,
		_w736_,
		_w738_,
		_w3672_
	);
	LUT4 #(
		.INIT('h3331)
	) name3210 (
		_w2055_,
		_w3670_,
		_w3671_,
		_w3672_,
		_w3673_
	);
	LUT2 #(
		.INIT('h2)
	) name3211 (
		_w1237_,
		_w3673_,
		_w3674_
	);
	LUT4 #(
		.INIT('h4844)
	) name3212 (
		_w1217_,
		_w2055_,
		_w2942_,
		_w2943_,
		_w3675_
	);
	LUT3 #(
		.INIT('ha8)
	) name3213 (
		_w2128_,
		_w3670_,
		_w3675_,
		_w3676_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3214 (
		_w2962_,
		_w2963_,
		_w2966_,
		_w2972_,
		_w3677_
	);
	LUT4 #(
		.INIT('h0b07)
	) name3215 (
		_w1217_,
		_w2055_,
		_w3670_,
		_w3677_,
		_w3678_
	);
	LUT4 #(
		.INIT('h8000)
	) name3216 (
		_w734_,
		_w749_,
		_w759_,
		_w833_,
		_w3679_
	);
	LUT4 #(
		.INIT('h1555)
	) name3217 (
		_w720_,
		_w842_,
		_w2859_,
		_w3679_,
		_w3680_
	);
	LUT4 #(
		.INIT('h0008)
	) name3218 (
		_w2055_,
		_w2170_,
		_w3168_,
		_w3680_,
		_w3681_
	);
	LUT3 #(
		.INIT('ha8)
	) name3219 (
		_w721_,
		_w2171_,
		_w2173_,
		_w3682_
	);
	LUT3 #(
		.INIT('h0b)
	) name3220 (
		_w720_,
		_w2177_,
		_w3682_,
		_w3683_
	);
	LUT2 #(
		.INIT('h4)
	) name3221 (
		_w3681_,
		_w3683_,
		_w3684_
	);
	LUT3 #(
		.INIT('hd0)
	) name3222 (
		_w2121_,
		_w3678_,
		_w3684_,
		_w3685_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3223 (
		_w2182_,
		_w3676_,
		_w3674_,
		_w3685_,
		_w3686_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3224 (
		\P1_reg3_reg[18]/NET0131 ,
		\P1_reg3_reg[19]/NET0131 ,
		_w591_,
		_w1244_,
		_w3687_
	);
	LUT2 #(
		.INIT('h2)
	) name3225 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3688_
	);
	LUT2 #(
		.INIT('h1)
	) name3226 (
		_w3687_,
		_w3688_,
		_w3689_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3227 (
		\P1_state_reg[0]/NET0131 ,
		_w3669_,
		_w3686_,
		_w3689_,
		_w3690_
	);
	LUT2 #(
		.INIT('h2)
	) name3228 (
		_w1749_,
		_w2903_,
		_w3691_
	);
	LUT4 #(
		.INIT('h00b7)
	) name3229 (
		_w2494_,
		_w2903_,
		_w3003_,
		_w3691_,
		_w3692_
	);
	LUT4 #(
		.INIT('h9555)
	) name3230 (
		_w1834_,
		_w1972_,
		_w1973_,
		_w1975_,
		_w3693_
	);
	LUT4 #(
		.INIT('h7020)
	) name3231 (
		_w1305_,
		_w1740_,
		_w2903_,
		_w3693_,
		_w3694_
	);
	LUT3 #(
		.INIT('ha8)
	) name3232 (
		_w2000_,
		_w3691_,
		_w3694_,
		_w3695_
	);
	LUT4 #(
		.INIT('h007b)
	) name3233 (
		_w2494_,
		_w2903_,
		_w3025_,
		_w3691_,
		_w3696_
	);
	LUT4 #(
		.INIT('h9000)
	) name3234 (
		_w1759_,
		_w2009_,
		_w2025_,
		_w2903_,
		_w3697_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3235 (
		_w1749_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w3698_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3236 (
		_w1759_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w3699_
	);
	LUT2 #(
		.INIT('h1)
	) name3237 (
		_w3698_,
		_w3699_,
		_w3700_
	);
	LUT2 #(
		.INIT('h4)
	) name3238 (
		_w3697_,
		_w3700_,
		_w3701_
	);
	LUT3 #(
		.INIT('hd0)
	) name3239 (
		_w1869_,
		_w3696_,
		_w3701_,
		_w3702_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3240 (
		_w1963_,
		_w3692_,
		_w3695_,
		_w3702_,
		_w3703_
	);
	LUT4 #(
		.INIT('h4000)
	) name3241 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1749_,
		_w3704_
	);
	LUT4 #(
		.INIT('haa08)
	) name3242 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w3703_,
		_w3704_,
		_w3705_
	);
	LUT2 #(
		.INIT('h4)
	) name3243 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		_w3706_
	);
	LUT3 #(
		.INIT('h07)
	) name3244 (
		_w1749_,
		_w2344_,
		_w3706_,
		_w3707_
	);
	LUT2 #(
		.INIT('hb)
	) name3245 (
		_w3705_,
		_w3707_,
		_w3708_
	);
	LUT4 #(
		.INIT('h4000)
	) name3246 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1803_,
		_w3709_
	);
	LUT2 #(
		.INIT('h2)
	) name3247 (
		_w1803_,
		_w2903_,
		_w3710_
	);
	LUT4 #(
		.INIT('h5655)
	) name3248 (
		_w1617_,
		_w1807_,
		_w1812_,
		_w1978_,
		_w3711_
	);
	LUT4 #(
		.INIT('h7020)
	) name3249 (
		_w1305_,
		_w1812_,
		_w2903_,
		_w3711_,
		_w3712_
	);
	LUT3 #(
		.INIT('ha8)
	) name3250 (
		_w2000_,
		_w3710_,
		_w3712_,
		_w3713_
	);
	LUT4 #(
		.INIT('hd200)
	) name3251 (
		_w2404_,
		_w2465_,
		_w2491_,
		_w2903_,
		_w3714_
	);
	LUT3 #(
		.INIT('ha8)
	) name3252 (
		_w1963_,
		_w3710_,
		_w3714_,
		_w3715_
	);
	LUT3 #(
		.INIT('h40)
	) name3253 (
		_w1830_,
		_w2009_,
		_w2010_,
		_w3716_
	);
	LUT4 #(
		.INIT('h1000)
	) name3254 (
		_w1820_,
		_w1830_,
		_w2009_,
		_w2010_,
		_w3717_
	);
	LUT4 #(
		.INIT('h0c04)
	) name3255 (
		_w1802_,
		_w2903_,
		_w3402_,
		_w3717_,
		_w3718_
	);
	LUT3 #(
		.INIT('ha8)
	) name3256 (
		_w2025_,
		_w3710_,
		_w3718_,
		_w3719_
	);
	LUT4 #(
		.INIT('h65aa)
	) name3257 (
		_w2491_,
		_w3025_,
		_w3028_,
		_w3034_,
		_w3720_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3258 (
		_w1803_,
		_w1869_,
		_w2903_,
		_w3720_,
		_w3721_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3259 (
		_w1802_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w3722_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3260 (
		_w1803_,
		_w2001_,
		_w2032_,
		_w2903_,
		_w3723_
	);
	LUT2 #(
		.INIT('h1)
	) name3261 (
		_w3722_,
		_w3723_,
		_w3724_
	);
	LUT3 #(
		.INIT('h10)
	) name3262 (
		_w3721_,
		_w3719_,
		_w3724_,
		_w3725_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3263 (
		_w1285_,
		_w3713_,
		_w3715_,
		_w3725_,
		_w3726_
	);
	LUT2 #(
		.INIT('h4)
	) name3264 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[16]/NET0131 ,
		_w3727_
	);
	LUT3 #(
		.INIT('h07)
	) name3265 (
		_w1803_,
		_w2344_,
		_w3727_,
		_w3728_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3266 (
		\P1_state_reg[0]/NET0131 ,
		_w3709_,
		_w3726_,
		_w3728_,
		_w3729_
	);
	LUT2 #(
		.INIT('h8)
	) name3267 (
		_w897_,
		_w2183_,
		_w3730_
	);
	LUT4 #(
		.INIT('h2220)
	) name3268 (
		_w897_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3731_
	);
	LUT3 #(
		.INIT('h80)
	) name3269 (
		_w488_,
		_w909_,
		_w910_,
		_w3732_
	);
	LUT4 #(
		.INIT('h00eb)
	) name3270 (
		_w488_,
		_w889_,
		_w2134_,
		_w3732_,
		_w3733_
	);
	LUT4 #(
		.INIT('hc808)
	) name3271 (
		_w897_,
		_w1237_,
		_w2055_,
		_w3733_,
		_w3734_
	);
	LUT4 #(
		.INIT('h6a55)
	) name3272 (
		_w1173_,
		_w2272_,
		_w2275_,
		_w2279_,
		_w3735_
	);
	LUT4 #(
		.INIT('he020)
	) name3273 (
		_w897_,
		_w2055_,
		_w2121_,
		_w3735_,
		_w3736_
	);
	LUT4 #(
		.INIT('h8488)
	) name3274 (
		_w1173_,
		_w2055_,
		_w2236_,
		_w2239_,
		_w3737_
	);
	LUT4 #(
		.INIT('h6a00)
	) name3275 (
		_w905_,
		_w915_,
		_w2159_,
		_w2170_,
		_w3738_
	);
	LUT3 #(
		.INIT('ha8)
	) name3276 (
		_w897_,
		_w2171_,
		_w2173_,
		_w3739_
	);
	LUT3 #(
		.INIT('h10)
	) name3277 (
		_w905_,
		_w2175_,
		_w2176_,
		_w3740_
	);
	LUT2 #(
		.INIT('h1)
	) name3278 (
		_w3739_,
		_w3740_,
		_w3741_
	);
	LUT3 #(
		.INIT('h70)
	) name3279 (
		_w2055_,
		_w3738_,
		_w3741_,
		_w3742_
	);
	LUT4 #(
		.INIT('h5700)
	) name3280 (
		_w2128_,
		_w3731_,
		_w3737_,
		_w3742_,
		_w3743_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3281 (
		_w2182_,
		_w3734_,
		_w3736_,
		_w3743_,
		_w3744_
	);
	LUT2 #(
		.INIT('h2)
	) name3282 (
		\P1_reg3_reg[9]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3745_
	);
	LUT4 #(
		.INIT('h4080)
	) name3283 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w897_,
		_w1242_,
		_w3746_
	);
	LUT2 #(
		.INIT('h1)
	) name3284 (
		_w3745_,
		_w3746_,
		_w3747_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3285 (
		\P1_state_reg[0]/NET0131 ,
		_w3730_,
		_w3744_,
		_w3747_,
		_w3748_
	);
	LUT2 #(
		.INIT('h2)
	) name3286 (
		\P2_reg2_reg[18]/NET0131 ,
		_w2042_,
		_w3749_
	);
	LUT4 #(
		.INIT('h2000)
	) name3287 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3750_
	);
	LUT2 #(
		.INIT('h2)
	) name3288 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1298_,
		_w3751_
	);
	LUT4 #(
		.INIT('he020)
	) name3289 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1298_,
		_w2000_,
		_w3418_,
		_w3752_
	);
	LUT4 #(
		.INIT('h2822)
	) name3290 (
		_w1298_,
		_w2511_,
		_w3099_,
		_w3100_,
		_w3753_
	);
	LUT3 #(
		.INIT('ha8)
	) name3291 (
		_w1869_,
		_w3751_,
		_w3753_,
		_w3754_
	);
	LUT4 #(
		.INIT('h8288)
	) name3292 (
		_w1298_,
		_w2511_,
		_w3113_,
		_w3116_,
		_w3755_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3293 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1298_,
		_w1626_,
		_w3403_,
		_w3756_
	);
	LUT4 #(
		.INIT('he200)
	) name3294 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1298_,
		_w1626_,
		_w2001_,
		_w3757_
	);
	LUT4 #(
		.INIT('h0200)
	) name3295 (
		_w1627_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w3758_
	);
	LUT4 #(
		.INIT('h0080)
	) name3296 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1863_,
		_w1866_,
		_w1999_,
		_w3759_
	);
	LUT2 #(
		.INIT('h1)
	) name3297 (
		_w3758_,
		_w3759_,
		_w3760_
	);
	LUT2 #(
		.INIT('h4)
	) name3298 (
		_w3757_,
		_w3760_,
		_w3761_
	);
	LUT3 #(
		.INIT('hd0)
	) name3299 (
		_w2025_,
		_w3756_,
		_w3761_,
		_w3762_
	);
	LUT4 #(
		.INIT('h5700)
	) name3300 (
		_w1963_,
		_w3751_,
		_w3755_,
		_w3762_,
		_w3763_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3301 (
		_w1285_,
		_w3752_,
		_w3754_,
		_w3763_,
		_w3764_
	);
	LUT4 #(
		.INIT('heeec)
	) name3302 (
		\P1_state_reg[0]/NET0131 ,
		_w3749_,
		_w3750_,
		_w3764_,
		_w3765_
	);
	LUT2 #(
		.INIT('h8)
	) name3303 (
		_w797_,
		_w2183_,
		_w3766_
	);
	LUT3 #(
		.INIT('h01)
	) name3304 (
		_w3574_,
		_w3576_,
		_w3579_,
		_w3767_
	);
	LUT3 #(
		.INIT('h20)
	) name3305 (
		_w796_,
		_w2175_,
		_w2176_,
		_w3768_
	);
	LUT3 #(
		.INIT('ha8)
	) name3306 (
		_w797_,
		_w2171_,
		_w2175_,
		_w3769_
	);
	LUT2 #(
		.INIT('h1)
	) name3307 (
		_w3768_,
		_w3769_,
		_w3770_
	);
	LUT4 #(
		.INIT('h7500)
	) name3308 (
		_w2055_,
		_w3573_,
		_w3767_,
		_w3770_,
		_w3771_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3309 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w3766_,
		_w3771_,
		_w3772_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3310 (
		\P1_reg3_reg[20]/NET0131 ,
		\P1_reg3_reg[21]/NET0131 ,
		_w593_,
		_w1244_,
		_w3773_
	);
	LUT2 #(
		.INIT('h2)
	) name3311 (
		\P1_reg3_reg[21]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3774_
	);
	LUT2 #(
		.INIT('h1)
	) name3312 (
		_w3773_,
		_w3774_,
		_w3775_
	);
	LUT2 #(
		.INIT('hb)
	) name3313 (
		_w3772_,
		_w3775_,
		_w3776_
	);
	LUT2 #(
		.INIT('h8)
	) name3314 (
		_w777_,
		_w2183_,
		_w3777_
	);
	LUT4 #(
		.INIT('h2220)
	) name3315 (
		_w777_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3778_
	);
	LUT4 #(
		.INIT('h22a2)
	) name3316 (
		_w2673_,
		_w2674_,
		_w2677_,
		_w3375_,
		_w3779_
	);
	LUT4 #(
		.INIT('h070b)
	) name3317 (
		_w1201_,
		_w2055_,
		_w3778_,
		_w3779_,
		_w3780_
	);
	LUT2 #(
		.INIT('h4)
	) name3318 (
		_w2650_,
		_w2659_,
		_w3781_
	);
	LUT2 #(
		.INIT('h2)
	) name3319 (
		_w2661_,
		_w3781_,
		_w3782_
	);
	LUT4 #(
		.INIT('h6a55)
	) name3320 (
		_w1201_,
		_w2657_,
		_w2659_,
		_w3782_,
		_w3783_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3321 (
		_w777_,
		_w2055_,
		_w2128_,
		_w3783_,
		_w3784_
	);
	LUT2 #(
		.INIT('h2)
	) name3322 (
		_w488_,
		_w800_,
		_w3785_
	);
	LUT4 #(
		.INIT('h4111)
	) name3323 (
		_w488_,
		_w789_,
		_w2141_,
		_w2213_,
		_w3786_
	);
	LUT3 #(
		.INIT('h70)
	) name3324 (
		_w2155_,
		_w2163_,
		_w2170_,
		_w3787_
	);
	LUT4 #(
		.INIT('h7500)
	) name3325 (
		_w776_,
		_w796_,
		_w3169_,
		_w3787_,
		_w3788_
	);
	LUT4 #(
		.INIT('h0057)
	) name3326 (
		_w1237_,
		_w3785_,
		_w3786_,
		_w3788_,
		_w3789_
	);
	LUT3 #(
		.INIT('h20)
	) name3327 (
		_w776_,
		_w2175_,
		_w2176_,
		_w3790_
	);
	LUT4 #(
		.INIT('h2220)
	) name3328 (
		_w1237_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3791_
	);
	LUT4 #(
		.INIT('h0001)
	) name3329 (
		_w2171_,
		_w2578_,
		_w2718_,
		_w3791_,
		_w3792_
	);
	LUT3 #(
		.INIT('h31)
	) name3330 (
		_w777_,
		_w3790_,
		_w3792_,
		_w3793_
	);
	LUT3 #(
		.INIT('hd0)
	) name3331 (
		_w2055_,
		_w3789_,
		_w3793_,
		_w3794_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3332 (
		_w2121_,
		_w3780_,
		_w3784_,
		_w3794_,
		_w3795_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3333 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w3777_,
		_w3795_,
		_w3796_
	);
	LUT2 #(
		.INIT('h2)
	) name3334 (
		\P1_reg3_reg[22]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3797_
	);
	LUT4 #(
		.INIT('h6a00)
	) name3335 (
		\P1_reg3_reg[22]/NET0131 ,
		_w593_,
		_w594_,
		_w1244_,
		_w3798_
	);
	LUT2 #(
		.INIT('h1)
	) name3336 (
		_w3797_,
		_w3798_,
		_w3799_
	);
	LUT2 #(
		.INIT('hb)
	) name3337 (
		_w3796_,
		_w3799_,
		_w3800_
	);
	LUT2 #(
		.INIT('h8)
	) name3338 (
		_w1561_,
		_w2039_,
		_w3801_
	);
	LUT2 #(
		.INIT('h2)
	) name3339 (
		_w1561_,
		_w2903_,
		_w3802_
	);
	LUT4 #(
		.INIT('h007b)
	) name3340 (
		_w2507_,
		_w2903_,
		_w3488_,
		_w3802_,
		_w3803_
	);
	LUT2 #(
		.INIT('h2)
	) name3341 (
		_w1869_,
		_w3803_,
		_w3804_
	);
	LUT4 #(
		.INIT('h00b7)
	) name3342 (
		_w2507_,
		_w2903_,
		_w3495_,
		_w3802_,
		_w3805_
	);
	LUT4 #(
		.INIT('h888a)
	) name3343 (
		_w2903_,
		_w3497_,
		_w3498_,
		_w3500_,
		_w3806_
	);
	LUT4 #(
		.INIT('h8040)
	) name3344 (
		_w1560_,
		_w2025_,
		_w2903_,
		_w3503_,
		_w3807_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3345 (
		_w1561_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w3808_
	);
	LUT3 #(
		.INIT('h0d)
	) name3346 (
		_w1560_,
		_w2993_,
		_w3808_,
		_w3809_
	);
	LUT2 #(
		.INIT('h4)
	) name3347 (
		_w3807_,
		_w3809_,
		_w3810_
	);
	LUT4 #(
		.INIT('h5700)
	) name3348 (
		_w2000_,
		_w3802_,
		_w3806_,
		_w3810_,
		_w3811_
	);
	LUT3 #(
		.INIT('hd0)
	) name3349 (
		_w1963_,
		_w3805_,
		_w3811_,
		_w3812_
	);
	LUT4 #(
		.INIT('h1311)
	) name3350 (
		_w1285_,
		_w3801_,
		_w3804_,
		_w3812_,
		_w3813_
	);
	LUT4 #(
		.INIT('h6a00)
	) name3351 (
		\P2_reg3_reg[22]/NET0131 ,
		_w1391_,
		_w1535_,
		_w2344_,
		_w3814_
	);
	LUT2 #(
		.INIT('h4)
	) name3352 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[22]/NET0131 ,
		_w3815_
	);
	LUT2 #(
		.INIT('h1)
	) name3353 (
		_w3814_,
		_w3815_,
		_w3816_
	);
	LUT3 #(
		.INIT('h2f)
	) name3354 (
		\P1_state_reg[0]/NET0131 ,
		_w3813_,
		_w3816_,
		_w3817_
	);
	LUT3 #(
		.INIT('h2a)
	) name3355 (
		\P1_reg2_reg[12]/NET0131 ,
		_w3175_,
		_w3512_,
		_w3818_
	);
	LUT4 #(
		.INIT('h1000)
	) name3356 (
		_w1096_,
		_w1098_,
		_w853_,
		_w1101_,
		_w3819_
	);
	LUT4 #(
		.INIT('hf100)
	) name3357 (
		_w489_,
		_w859_,
		_w863_,
		_w2194_,
		_w3820_
	);
	LUT4 #(
		.INIT('haa8a)
	) name3358 (
		_w2189_,
		_w3350_,
		_w3358_,
		_w3820_,
		_w3821_
	);
	LUT4 #(
		.INIT('heeec)
	) name3359 (
		_w3511_,
		_w3818_,
		_w3819_,
		_w3821_,
		_w3822_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name3360 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[18]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3823_
	);
	LUT2 #(
		.INIT('h8)
	) name3361 (
		\P1_reg2_reg[18]/NET0131 ,
		_w2183_,
		_w3824_
	);
	LUT4 #(
		.INIT('haa8a)
	) name3362 (
		\P1_reg2_reg[18]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3825_
	);
	LUT4 #(
		.INIT('h8848)
	) name3363 (
		_w1216_,
		_w2189_,
		_w2650_,
		_w2657_,
		_w3826_
	);
	LUT3 #(
		.INIT('ha8)
	) name3364 (
		_w2128_,
		_w3825_,
		_w3826_,
		_w3827_
	);
	LUT4 #(
		.INIT('h4484)
	) name3365 (
		_w1216_,
		_w2189_,
		_w2677_,
		_w3375_,
		_w3828_
	);
	LUT3 #(
		.INIT('ha8)
	) name3366 (
		_w2121_,
		_w3825_,
		_w3828_,
		_w3829_
	);
	LUT4 #(
		.INIT('hc808)
	) name3367 (
		\P1_reg2_reg[18]/NET0131 ,
		_w1237_,
		_w2189_,
		_w3379_,
		_w3830_
	);
	LUT2 #(
		.INIT('h4)
	) name3368 (
		_w734_,
		_w2194_,
		_w3831_
	);
	LUT4 #(
		.INIT('haa20)
	) name3369 (
		_w2189_,
		_w3381_,
		_w3382_,
		_w3831_,
		_w3832_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3370 (
		\P1_reg2_reg[18]/NET0131 ,
		_w2171_,
		_w2196_,
		_w3187_,
		_w3833_
	);
	LUT4 #(
		.INIT('h1000)
	) name3371 (
		_w1096_,
		_w1098_,
		_w735_,
		_w1101_,
		_w3834_
	);
	LUT2 #(
		.INIT('h1)
	) name3372 (
		_w3833_,
		_w3834_,
		_w3835_
	);
	LUT2 #(
		.INIT('h4)
	) name3373 (
		_w3832_,
		_w3835_,
		_w3836_
	);
	LUT2 #(
		.INIT('h4)
	) name3374 (
		_w3830_,
		_w3836_,
		_w3837_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3375 (
		_w2182_,
		_w3829_,
		_w3827_,
		_w3837_,
		_w3838_
	);
	LUT4 #(
		.INIT('heeec)
	) name3376 (
		\P1_state_reg[0]/NET0131 ,
		_w3823_,
		_w3824_,
		_w3838_,
		_w3839_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name3377 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[21]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3840_
	);
	LUT2 #(
		.INIT('h8)
	) name3378 (
		\P1_reg2_reg[21]/NET0131 ,
		_w2183_,
		_w3841_
	);
	LUT4 #(
		.INIT('h5545)
	) name3379 (
		\P1_reg2_reg[21]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3842_
	);
	LUT2 #(
		.INIT('h2)
	) name3380 (
		_w2170_,
		_w3842_,
		_w3843_
	);
	LUT4 #(
		.INIT('hb700)
	) name3381 (
		_w796_,
		_w2189_,
		_w3169_,
		_w3843_,
		_w3844_
	);
	LUT2 #(
		.INIT('h8)
	) name3382 (
		_w797_,
		_w1120_,
		_w3845_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3383 (
		\P1_reg2_reg[21]/NET0131 ,
		_w2171_,
		_w2196_,
		_w2866_,
		_w3846_
	);
	LUT2 #(
		.INIT('h1)
	) name3384 (
		_w3845_,
		_w3846_,
		_w3847_
	);
	LUT2 #(
		.INIT('h4)
	) name3385 (
		_w3844_,
		_w3847_,
		_w3848_
	);
	LUT4 #(
		.INIT('h7500)
	) name3386 (
		_w2189_,
		_w3573_,
		_w3580_,
		_w3848_,
		_w3849_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3387 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w3841_,
		_w3849_,
		_w3850_
	);
	LUT2 #(
		.INIT('he)
	) name3388 (
		_w3840_,
		_w3850_,
		_w3851_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name3389 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[22]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3852_
	);
	LUT2 #(
		.INIT('h8)
	) name3390 (
		\P1_reg2_reg[22]/NET0131 ,
		_w2183_,
		_w3853_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3391 (
		\P1_reg2_reg[22]/NET0131 ,
		_w1201_,
		_w2189_,
		_w3779_,
		_w3854_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3392 (
		\P1_reg2_reg[22]/NET0131 ,
		_w2128_,
		_w2189_,
		_w3783_,
		_w3855_
	);
	LUT4 #(
		.INIT('h5400)
	) name3393 (
		_w489_,
		_w773_,
		_w775_,
		_w2194_,
		_w3856_
	);
	LUT4 #(
		.INIT('hfb00)
	) name3394 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2782_,
		_w3857_
	);
	LUT3 #(
		.INIT('h01)
	) name3395 (
		_w2171_,
		_w2196_,
		_w3857_,
		_w3858_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3396 (
		\P1_reg2_reg[22]/NET0131 ,
		_w2171_,
		_w2196_,
		_w3857_,
		_w3859_
	);
	LUT2 #(
		.INIT('h8)
	) name3397 (
		_w777_,
		_w1120_,
		_w3860_
	);
	LUT2 #(
		.INIT('h1)
	) name3398 (
		_w3859_,
		_w3860_,
		_w3861_
	);
	LUT4 #(
		.INIT('h5d00)
	) name3399 (
		_w2189_,
		_w3789_,
		_w3856_,
		_w3861_,
		_w3862_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3400 (
		_w2121_,
		_w3854_,
		_w3855_,
		_w3862_,
		_w3863_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3401 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w3853_,
		_w3863_,
		_w3864_
	);
	LUT2 #(
		.INIT('he)
	) name3402 (
		_w3852_,
		_w3864_,
		_w3865_
	);
	LUT4 #(
		.INIT('h7020)
	) name3403 (
		_w1305_,
		_w1807_,
		_w2000_,
		_w3395_,
		_w3866_
	);
	LUT3 #(
		.INIT('h82)
	) name3404 (
		_w1869_,
		_w2508_,
		_w2880_,
		_w3867_
	);
	LUT4 #(
		.INIT('hc048)
	) name3405 (
		_w1923_,
		_w1963_,
		_w2508_,
		_w3398_,
		_w3868_
	);
	LUT2 #(
		.INIT('h8)
	) name3406 (
		_w1612_,
		_w2001_,
		_w3869_
	);
	LUT3 #(
		.INIT('h07)
	) name3407 (
		_w2025_,
		_w3404_,
		_w3869_,
		_w3870_
	);
	LUT4 #(
		.INIT('h0100)
	) name3408 (
		_w3866_,
		_w3868_,
		_w3867_,
		_w3870_,
		_w3871_
	);
	LUT4 #(
		.INIT('hf010)
	) name3409 (
		_w1963_,
		_w2033_,
		_w2734_,
		_w2762_,
		_w3872_
	);
	LUT4 #(
		.INIT('h1530)
	) name3410 (
		_w1595_,
		_w1859_,
		_w1863_,
		_w1866_,
		_w3873_
	);
	LUT3 #(
		.INIT('h10)
	) name3411 (
		_w1867_,
		_w2762_,
		_w3873_,
		_w3874_
	);
	LUT4 #(
		.INIT('hf2f3)
	) name3412 (
		_w1867_,
		_w2000_,
		_w2762_,
		_w3873_,
		_w3875_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3413 (
		\P2_reg1_reg[17]/NET0131 ,
		_w2556_,
		_w3872_,
		_w3875_,
		_w3876_
	);
	LUT3 #(
		.INIT('hf2)
	) name3414 (
		_w3244_,
		_w3871_,
		_w3876_,
		_w3877_
	);
	LUT2 #(
		.INIT('h2)
	) name3415 (
		\P2_reg1_reg[18]/NET0131 ,
		_w2042_,
		_w3878_
	);
	LUT4 #(
		.INIT('h2000)
	) name3416 (
		\P2_reg1_reg[18]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3879_
	);
	LUT2 #(
		.INIT('h2)
	) name3417 (
		\P2_reg1_reg[18]/NET0131 ,
		_w2762_,
		_w3880_
	);
	LUT4 #(
		.INIT('hc808)
	) name3418 (
		\P2_reg1_reg[18]/NET0131 ,
		_w2000_,
		_w2762_,
		_w3418_,
		_w3881_
	);
	LUT4 #(
		.INIT('h4844)
	) name3419 (
		_w2511_,
		_w2762_,
		_w3099_,
		_w3100_,
		_w3882_
	);
	LUT3 #(
		.INIT('ha8)
	) name3420 (
		_w1869_,
		_w3880_,
		_w3882_,
		_w3883_
	);
	LUT4 #(
		.INIT('h8288)
	) name3421 (
		_w1963_,
		_w2511_,
		_w3113_,
		_w3116_,
		_w3884_
	);
	LUT2 #(
		.INIT('h8)
	) name3422 (
		_w1626_,
		_w2001_,
		_w3885_
	);
	LUT4 #(
		.INIT('h007b)
	) name3423 (
		_w1626_,
		_w2025_,
		_w3403_,
		_w3885_,
		_w3886_
	);
	LUT2 #(
		.INIT('h2)
	) name3424 (
		\P2_reg1_reg[18]/NET0131 ,
		_w3872_,
		_w3887_
	);
	LUT4 #(
		.INIT('h0075)
	) name3425 (
		_w2762_,
		_w3884_,
		_w3886_,
		_w3887_,
		_w3888_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3426 (
		_w1285_,
		_w3881_,
		_w3883_,
		_w3888_,
		_w3889_
	);
	LUT4 #(
		.INIT('heeec)
	) name3427 (
		\P1_state_reg[0]/NET0131 ,
		_w3878_,
		_w3879_,
		_w3889_,
		_w3890_
	);
	LUT3 #(
		.INIT('h45)
	) name3428 (
		_w1284_,
		_w2762_,
		_w3873_,
		_w3891_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3429 (
		\P2_reg1_reg[19]/NET0131 ,
		_w2042_,
		_w3872_,
		_w3891_,
		_w3892_
	);
	LUT3 #(
		.INIT('ha8)
	) name3430 (
		_w2000_,
		_w3438_,
		_w3440_,
		_w3893_
	);
	LUT4 #(
		.INIT('h2300)
	) name3431 (
		_w1306_,
		_w1596_,
		_w1598_,
		_w2001_,
		_w3894_
	);
	LUT4 #(
		.INIT('h0001)
	) name3432 (
		_w3435_,
		_w3436_,
		_w3434_,
		_w3894_,
		_w3895_
	);
	LUT4 #(
		.INIT('hecee)
	) name3433 (
		_w3244_,
		_w3892_,
		_w3893_,
		_w3895_,
		_w3896_
	);
	LUT2 #(
		.INIT('h2)
	) name3434 (
		\P2_reg1_reg[22]/NET0131 ,
		_w2042_,
		_w3897_
	);
	LUT4 #(
		.INIT('h2000)
	) name3435 (
		\P2_reg1_reg[22]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3898_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3436 (
		\P2_reg1_reg[22]/NET0131 ,
		_w2507_,
		_w2762_,
		_w3488_,
		_w3899_
	);
	LUT2 #(
		.INIT('h2)
	) name3437 (
		_w1869_,
		_w3899_,
		_w3900_
	);
	LUT4 #(
		.INIT('hc535)
	) name3438 (
		\P2_reg1_reg[22]/NET0131 ,
		_w2507_,
		_w2762_,
		_w3495_,
		_w3901_
	);
	LUT2 #(
		.INIT('h2)
	) name3439 (
		\P2_reg1_reg[22]/NET0131 ,
		_w3226_,
		_w3902_
	);
	LUT4 #(
		.INIT('h0075)
	) name3440 (
		_w2762_,
		_w3501_,
		_w3504_,
		_w3902_,
		_w3903_
	);
	LUT3 #(
		.INIT('hd0)
	) name3441 (
		_w1963_,
		_w3901_,
		_w3903_,
		_w3904_
	);
	LUT4 #(
		.INIT('h1311)
	) name3442 (
		_w1285_,
		_w3898_,
		_w3900_,
		_w3904_,
		_w3905_
	);
	LUT3 #(
		.INIT('hce)
	) name3443 (
		\P1_state_reg[0]/NET0131 ,
		_w3897_,
		_w3905_,
		_w3906_
	);
	LUT3 #(
		.INIT('h2a)
	) name3444 (
		\P1_reg0_reg[12]/NET0131 ,
		_w3511_,
		_w3561_,
		_w3907_
	);
	LUT4 #(
		.INIT('hf0b0)
	) name3445 (
		_w3350_,
		_w3358_,
		_w3563_,
		_w3820_,
		_w3908_
	);
	LUT2 #(
		.INIT('he)
	) name3446 (
		_w3907_,
		_w3908_,
		_w3909_
	);
	LUT4 #(
		.INIT('h6300)
	) name3447 (
		_w674_,
		_w647_,
		_w2168_,
		_w2170_,
		_w3910_
	);
	LUT3 #(
		.INIT('h10)
	) name3448 (
		_w489_,
		_w646_,
		_w2194_,
		_w3911_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3449 (
		_w2189_,
		_w2857_,
		_w3911_,
		_w3910_,
		_w3912_
	);
	LUT4 #(
		.INIT('h5545)
	) name3450 (
		_w1120_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3913_
	);
	LUT2 #(
		.INIT('h4)
	) name3451 (
		_w2171_,
		_w3511_,
		_w3914_
	);
	LUT3 #(
		.INIT('h8a)
	) name3452 (
		\P1_reg2_reg[30]/NET0131 ,
		_w3913_,
		_w3914_,
		_w3915_
	);
	LUT4 #(
		.INIT('hffc8)
	) name3453 (
		_w2316_,
		_w3511_,
		_w3912_,
		_w3915_,
		_w3916_
	);
	LUT2 #(
		.INIT('h4)
	) name3454 (
		_w1298_,
		_w1869_,
		_w3917_
	);
	LUT2 #(
		.INIT('h4)
	) name3455 (
		_w1298_,
		_w1963_,
		_w3918_
	);
	LUT3 #(
		.INIT('hab)
	) name3456 (
		_w1298_,
		_w1869_,
		_w1963_,
		_w3919_
	);
	LUT4 #(
		.INIT('h4000)
	) name3457 (
		_w2031_,
		_w2556_,
		_w2640_,
		_w3919_,
		_w3920_
	);
	LUT2 #(
		.INIT('h2)
	) name3458 (
		\P2_reg2_reg[17]/NET0131 ,
		_w3920_,
		_w3921_
	);
	LUT4 #(
		.INIT('h0200)
	) name3459 (
		_w1613_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w3922_
	);
	LUT4 #(
		.INIT('hcc08)
	) name3460 (
		_w1298_,
		_w2556_,
		_w3871_,
		_w3922_,
		_w3923_
	);
	LUT2 #(
		.INIT('he)
	) name3461 (
		_w3921_,
		_w3923_,
		_w3924_
	);
	LUT4 #(
		.INIT('h0200)
	) name3462 (
		_w1600_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w3925_
	);
	LUT4 #(
		.INIT('h0075)
	) name3463 (
		_w1298_,
		_w3893_,
		_w3895_,
		_w3925_,
		_w3926_
	);
	LUT3 #(
		.INIT('hc8)
	) name3464 (
		_w1298_,
		_w2556_,
		_w3154_,
		_w3927_
	);
	LUT3 #(
		.INIT('h8a)
	) name3465 (
		\P2_reg2_reg[19]/NET0131 ,
		_w2639_,
		_w3927_,
		_w3928_
	);
	LUT3 #(
		.INIT('hf2)
	) name3466 (
		_w2556_,
		_w3926_,
		_w3928_,
		_w3929_
	);
	LUT2 #(
		.INIT('h2)
	) name3467 (
		\P2_reg2_reg[20]/NET0131 ,
		_w2042_,
		_w3930_
	);
	LUT4 #(
		.INIT('h2000)
	) name3468 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3931_
	);
	LUT4 #(
		.INIT('h65aa)
	) name3469 (
		_w2510_,
		_w3003_,
		_w3004_,
		_w3005_,
		_w3932_
	);
	LUT4 #(
		.INIT('he020)
	) name3470 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1298_,
		_w1963_,
		_w3932_,
		_w3933_
	);
	LUT4 #(
		.INIT('h8000)
	) name3471 (
		_w2009_,
		_w2010_,
		_w2012_,
		_w2017_,
		_w3934_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3472 (
		_w1587_,
		_w1599_,
		_w1626_,
		_w3403_,
		_w3935_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3473 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1298_,
		_w3934_,
		_w3935_,
		_w3936_
	);
	LUT2 #(
		.INIT('h2)
	) name3474 (
		_w2025_,
		_w3936_,
		_w3937_
	);
	LUT4 #(
		.INIT('h1444)
	) name3475 (
		_w1305_,
		_w1573_,
		_w1978_,
		_w1982_,
		_w3938_
	);
	LUT4 #(
		.INIT('h0200)
	) name3476 (
		_w1305_,
		_w1602_,
		_w1601_,
		_w1603_,
		_w3939_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3477 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1298_,
		_w3938_,
		_w3939_,
		_w3940_
	);
	LUT2 #(
		.INIT('h2)
	) name3478 (
		_w2000_,
		_w3940_,
		_w3941_
	);
	LUT3 #(
		.INIT('h10)
	) name3479 (
		_w1306_,
		_w1586_,
		_w2001_,
		_w3942_
	);
	LUT4 #(
		.INIT('h007d)
	) name3480 (
		_w1869_,
		_w2510_,
		_w3040_,
		_w3942_,
		_w3943_
	);
	LUT2 #(
		.INIT('h8)
	) name3481 (
		_w1588_,
		_w2029_,
		_w3944_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3482 (
		_w1298_,
		_w1869_,
		_w2001_,
		_w2032_,
		_w3945_
	);
	LUT3 #(
		.INIT('h31)
	) name3483 (
		\P2_reg2_reg[20]/NET0131 ,
		_w3944_,
		_w3945_,
		_w3946_
	);
	LUT3 #(
		.INIT('hd0)
	) name3484 (
		_w1298_,
		_w3943_,
		_w3946_,
		_w3947_
	);
	LUT4 #(
		.INIT('h0100)
	) name3485 (
		_w3937_,
		_w3933_,
		_w3941_,
		_w3947_,
		_w3948_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3486 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w3931_,
		_w3948_,
		_w3949_
	);
	LUT2 #(
		.INIT('he)
	) name3487 (
		_w3930_,
		_w3949_,
		_w3950_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3488 (
		\P1_reg0_reg[17]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w3951_
	);
	LUT4 #(
		.INIT('h7200)
	) name3489 (
		_w488_,
		_w764_,
		_w3453_,
		_w3563_,
		_w3952_
	);
	LUT3 #(
		.INIT('ha8)
	) name3490 (
		_w1237_,
		_w3951_,
		_w3952_,
		_w3953_
	);
	LUT2 #(
		.INIT('h4)
	) name3491 (
		_w2798_,
		_w3511_,
		_w3954_
	);
	LUT4 #(
		.INIT('h2300)
	) name3492 (
		_w1236_,
		_w2798_,
		_w3295_,
		_w3511_,
		_w3955_
	);
	LUT3 #(
		.INIT('h2a)
	) name3493 (
		\P1_reg0_reg[17]/NET0131 ,
		_w2797_,
		_w3955_,
		_w3956_
	);
	LUT4 #(
		.INIT('h0075)
	) name3494 (
		_w3563_,
		_w3613_,
		_w3616_,
		_w3956_,
		_w3957_
	);
	LUT2 #(
		.INIT('hb)
	) name3495 (
		_w3953_,
		_w3957_,
		_w3958_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name3496 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[20]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3959_
	);
	LUT3 #(
		.INIT('h02)
	) name3497 (
		_w1237_,
		_w3163_,
		_w3164_,
		_w3960_
	);
	LUT4 #(
		.INIT('h6500)
	) name3498 (
		_w1228_,
		_w2093_,
		_w2102_,
		_w2121_,
		_w3961_
	);
	LUT4 #(
		.INIT('h4000)
	) name3499 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2182_,
		_w3962_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3500 (
		_w3171_,
		_w3961_,
		_w3960_,
		_w3962_,
		_w3963_
	);
	LUT3 #(
		.INIT('h84)
	) name3501 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[20]/NET0131 ,
		_w1242_,
		_w3964_
	);
	LUT3 #(
		.INIT('hb0)
	) name3502 (
		_w1252_,
		_w3561_,
		_w3964_,
		_w3965_
	);
	LUT4 #(
		.INIT('heeec)
	) name3503 (
		\P1_state_reg[0]/NET0131 ,
		_w3959_,
		_w3963_,
		_w3965_,
		_w3966_
	);
	LUT3 #(
		.INIT('h2a)
	) name3504 (
		\P1_reg0_reg[30]/NET0131 ,
		_w2332_,
		_w3563_,
		_w3967_
	);
	LUT4 #(
		.INIT('hccc8)
	) name3505 (
		_w2857_,
		_w3563_,
		_w3911_,
		_w3910_,
		_w3968_
	);
	LUT2 #(
		.INIT('he)
	) name3506 (
		_w3967_,
		_w3968_,
		_w3969_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3507 (
		\P1_reg1_reg[12]/NET0131 ,
		_w2820_,
		_w3511_,
		_w3606_,
		_w3970_
	);
	LUT4 #(
		.INIT('hf0b0)
	) name3508 (
		_w3350_,
		_w3358_,
		_w3608_,
		_w3820_,
		_w3971_
	);
	LUT2 #(
		.INIT('he)
	) name3509 (
		_w3970_,
		_w3971_,
		_w3972_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name3510 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[20]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w3973_
	);
	LUT2 #(
		.INIT('h8)
	) name3511 (
		\P1_reg1_reg[20]/NET0131 ,
		_w2183_,
		_w3974_
	);
	LUT4 #(
		.INIT('hef00)
	) name3512 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2172_,
		_w3975_
	);
	LUT4 #(
		.INIT('h0002)
	) name3513 (
		_w2332_,
		_w2820_,
		_w3605_,
		_w3975_,
		_w3976_
	);
	LUT2 #(
		.INIT('h2)
	) name3514 (
		\P1_reg1_reg[20]/NET0131 ,
		_w3976_,
		_w3977_
	);
	LUT4 #(
		.INIT('haaa2)
	) name3515 (
		_w2536_,
		_w3171_,
		_w3961_,
		_w3960_,
		_w3978_
	);
	LUT4 #(
		.INIT('h1113)
	) name3516 (
		_w2182_,
		_w3974_,
		_w3977_,
		_w3978_,
		_w3979_
	);
	LUT3 #(
		.INIT('hce)
	) name3517 (
		\P1_state_reg[0]/NET0131 ,
		_w3973_,
		_w3979_,
		_w3980_
	);
	LUT2 #(
		.INIT('h2)
	) name3518 (
		_w1963_,
		_w2729_,
		_w3981_
	);
	LUT4 #(
		.INIT('hf100)
	) name3519 (
		_w1963_,
		_w2033_,
		_w2729_,
		_w2734_,
		_w3982_
	);
	LUT2 #(
		.INIT('h4)
	) name3520 (
		_w2729_,
		_w3873_,
		_w3983_
	);
	LUT3 #(
		.INIT('h8a)
	) name3521 (
		_w2556_,
		_w2729_,
		_w3873_,
		_w3984_
	);
	LUT3 #(
		.INIT('h2a)
	) name3522 (
		\P2_reg0_reg[17]/NET0131 ,
		_w3982_,
		_w3984_,
		_w3985_
	);
	LUT3 #(
		.INIT('hf2)
	) name3523 (
		_w3153_,
		_w3871_,
		_w3985_,
		_w3986_
	);
	LUT2 #(
		.INIT('h2)
	) name3524 (
		\P2_reg0_reg[18]/NET0131 ,
		_w2042_,
		_w3987_
	);
	LUT4 #(
		.INIT('h2000)
	) name3525 (
		\P2_reg0_reg[18]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w3988_
	);
	LUT2 #(
		.INIT('h2)
	) name3526 (
		\P2_reg0_reg[18]/NET0131 ,
		_w2729_,
		_w3989_
	);
	LUT4 #(
		.INIT('hc808)
	) name3527 (
		\P2_reg0_reg[18]/NET0131 ,
		_w2000_,
		_w2729_,
		_w3418_,
		_w3990_
	);
	LUT4 #(
		.INIT('h4844)
	) name3528 (
		_w2511_,
		_w2729_,
		_w3099_,
		_w3100_,
		_w3991_
	);
	LUT3 #(
		.INIT('ha8)
	) name3529 (
		_w1869_,
		_w3989_,
		_w3991_,
		_w3992_
	);
	LUT2 #(
		.INIT('h2)
	) name3530 (
		\P2_reg0_reg[18]/NET0131 ,
		_w3982_,
		_w3993_
	);
	LUT4 #(
		.INIT('h0075)
	) name3531 (
		_w2729_,
		_w3884_,
		_w3886_,
		_w3993_,
		_w3994_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3532 (
		_w1285_,
		_w3990_,
		_w3992_,
		_w3994_,
		_w3995_
	);
	LUT4 #(
		.INIT('heeec)
	) name3533 (
		\P1_state_reg[0]/NET0131 ,
		_w3987_,
		_w3988_,
		_w3995_,
		_w3996_
	);
	LUT3 #(
		.INIT('h2a)
	) name3534 (
		\P1_reg1_reg[30]/NET0131 ,
		_w2332_,
		_w3608_,
		_w3997_
	);
	LUT4 #(
		.INIT('hccc8)
	) name3535 (
		_w2857_,
		_w3608_,
		_w3911_,
		_w3910_,
		_w3998_
	);
	LUT2 #(
		.INIT('he)
	) name3536 (
		_w3997_,
		_w3998_,
		_w3999_
	);
	LUT3 #(
		.INIT('h2a)
	) name3537 (
		\P2_reg0_reg[19]/NET0131 ,
		_w3982_,
		_w3984_,
		_w4000_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3538 (
		_w3153_,
		_w3893_,
		_w3895_,
		_w4000_,
		_w4001_
	);
	LUT2 #(
		.INIT('h8)
	) name3539 (
		_w874_,
		_w2183_,
		_w4002_
	);
	LUT4 #(
		.INIT('h2220)
	) name3540 (
		_w874_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4003_
	);
	LUT4 #(
		.INIT('h5655)
	) name3541 (
		_w856_,
		_w876_,
		_w889_,
		_w2134_,
		_w4004_
	);
	LUT4 #(
		.INIT('h7020)
	) name3542 (
		_w488_,
		_w889_,
		_w2055_,
		_w4004_,
		_w4005_
	);
	LUT3 #(
		.INIT('ha8)
	) name3543 (
		_w1237_,
		_w4003_,
		_w4005_,
		_w4006_
	);
	LUT4 #(
		.INIT('h8488)
	) name3544 (
		_w1174_,
		_w2055_,
		_w2962_,
		_w2963_,
		_w4007_
	);
	LUT3 #(
		.INIT('ha8)
	) name3545 (
		_w2121_,
		_w4003_,
		_w4007_,
		_w4008_
	);
	LUT3 #(
		.INIT('he0)
	) name3546 (
		_w881_,
		_w883_,
		_w2194_,
		_w4009_
	);
	LUT4 #(
		.INIT('h1555)
	) name3547 (
		_w884_,
		_w893_,
		_w2159_,
		_w2160_,
		_w4010_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3548 (
		_w2159_,
		_w2160_,
		_w2161_,
		_w2170_,
		_w4011_
	);
	LUT3 #(
		.INIT('h45)
	) name3549 (
		_w4009_,
		_w4010_,
		_w4011_,
		_w4012_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3550 (
		_w1174_,
		_w2128_,
		_w2938_,
		_w4012_,
		_w4013_
	);
	LUT3 #(
		.INIT('he0)
	) name3551 (
		_w881_,
		_w883_,
		_w1120_,
		_w4014_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3552 (
		_w874_,
		_w2171_,
		_w2173_,
		_w2845_,
		_w4015_
	);
	LUT2 #(
		.INIT('h1)
	) name3553 (
		_w4014_,
		_w4015_,
		_w4016_
	);
	LUT3 #(
		.INIT('hd0)
	) name3554 (
		_w2055_,
		_w4013_,
		_w4016_,
		_w4017_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3555 (
		_w2182_,
		_w4006_,
		_w4008_,
		_w4017_,
		_w4018_
	);
	LUT2 #(
		.INIT('h2)
	) name3556 (
		\P1_reg3_reg[11]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4019_
	);
	LUT4 #(
		.INIT('h4080)
	) name3557 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w874_,
		_w1242_,
		_w4020_
	);
	LUT2 #(
		.INIT('h1)
	) name3558 (
		_w4019_,
		_w4020_,
		_w4021_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3559 (
		\P1_state_reg[0]/NET0131 ,
		_w4002_,
		_w4018_,
		_w4021_,
		_w4022_
	);
	LUT2 #(
		.INIT('h8)
	) name3560 (
		_w886_,
		_w2183_,
		_w4023_
	);
	LUT4 #(
		.INIT('h2220)
	) name3561 (
		_w886_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4024_
	);
	LUT4 #(
		.INIT('h4144)
	) name3562 (
		_w488_,
		_w876_,
		_w889_,
		_w2134_,
		_w4025_
	);
	LUT3 #(
		.INIT('h80)
	) name3563 (
		_w488_,
		_w896_,
		_w898_,
		_w4026_
	);
	LUT4 #(
		.INIT('h3331)
	) name3564 (
		_w2055_,
		_w4024_,
		_w4025_,
		_w4026_,
		_w4027_
	);
	LUT2 #(
		.INIT('h2)
	) name3565 (
		_w1237_,
		_w4027_,
		_w4028_
	);
	LUT4 #(
		.INIT('h00b7)
	) name3566 (
		_w1178_,
		_w2055_,
		_w2682_,
		_w4024_,
		_w4029_
	);
	LUT2 #(
		.INIT('h2)
	) name3567 (
		_w2121_,
		_w4029_,
		_w4030_
	);
	LUT4 #(
		.INIT('h007b)
	) name3568 (
		_w1178_,
		_w2055_,
		_w2653_,
		_w4024_,
		_w4031_
	);
	LUT2 #(
		.INIT('h4)
	) name3569 (
		_w893_,
		_w2194_,
		_w4032_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3570 (
		_w893_,
		_w2159_,
		_w2160_,
		_w2170_,
		_w4033_
	);
	LUT4 #(
		.INIT('h6a00)
	) name3571 (
		_w893_,
		_w2159_,
		_w2160_,
		_w2170_,
		_w4034_
	);
	LUT2 #(
		.INIT('h4)
	) name3572 (
		_w893_,
		_w1120_,
		_w4035_
	);
	LUT4 #(
		.INIT('h0057)
	) name3573 (
		_w886_,
		_w2171_,
		_w2173_,
		_w4035_,
		_w4036_
	);
	LUT4 #(
		.INIT('h5700)
	) name3574 (
		_w2055_,
		_w4032_,
		_w4034_,
		_w4036_,
		_w4037_
	);
	LUT3 #(
		.INIT('hd0)
	) name3575 (
		_w2128_,
		_w4031_,
		_w4037_,
		_w4038_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3576 (
		_w2182_,
		_w4028_,
		_w4030_,
		_w4038_,
		_w4039_
	);
	LUT2 #(
		.INIT('h2)
	) name3577 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4040_
	);
	LUT4 #(
		.INIT('h4080)
	) name3578 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w886_,
		_w1242_,
		_w4041_
	);
	LUT2 #(
		.INIT('h1)
	) name3579 (
		_w4040_,
		_w4041_,
		_w4042_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3580 (
		\P1_state_reg[0]/NET0131 ,
		_w4023_,
		_w4039_,
		_w4042_,
		_w4043_
	);
	LUT2 #(
		.INIT('h8)
	) name3581 (
		_w835_,
		_w2183_,
		_w4044_
	);
	LUT4 #(
		.INIT('h0d05)
	) name3582 (
		_w827_,
		_w2135_,
		_w2138_,
		_w3351_,
		_w4045_
	);
	LUT4 #(
		.INIT('h80d0)
	) name3583 (
		_w488_,
		_w847_,
		_w2055_,
		_w4045_,
		_w4046_
	);
	LUT4 #(
		.INIT('h1110)
	) name3584 (
		_w835_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4047_
	);
	LUT2 #(
		.INIT('h2)
	) name3585 (
		_w1237_,
		_w4047_,
		_w4048_
	);
	LUT2 #(
		.INIT('h4)
	) name3586 (
		_w4046_,
		_w4048_,
		_w4049_
	);
	LUT4 #(
		.INIT('h4500)
	) name3587 (
		_w1189_,
		_w2653_,
		_w2654_,
		_w2655_,
		_w4050_
	);
	LUT4 #(
		.INIT('h20aa)
	) name3588 (
		_w1189_,
		_w2653_,
		_w2654_,
		_w2655_,
		_w4051_
	);
	LUT3 #(
		.INIT('h02)
	) name3589 (
		_w2128_,
		_w4051_,
		_w4050_,
		_w4052_
	);
	LUT3 #(
		.INIT('h48)
	) name3590 (
		_w842_,
		_w2170_,
		_w2859_,
		_w4053_
	);
	LUT4 #(
		.INIT('h00b7)
	) name3591 (
		_w1189_,
		_w2121_,
		_w3374_,
		_w4053_,
		_w4054_
	);
	LUT3 #(
		.INIT('h10)
	) name3592 (
		_w842_,
		_w2175_,
		_w2176_,
		_w4055_
	);
	LUT4 #(
		.INIT('h5400)
	) name3593 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2120_,
		_w4056_
	);
	LUT4 #(
		.INIT('h0001)
	) name3594 (
		_w2171_,
		_w2578_,
		_w2718_,
		_w4056_,
		_w4057_
	);
	LUT3 #(
		.INIT('h31)
	) name3595 (
		_w835_,
		_w4055_,
		_w4057_,
		_w4058_
	);
	LUT4 #(
		.INIT('h7500)
	) name3596 (
		_w2055_,
		_w4052_,
		_w4054_,
		_w4058_,
		_w4059_
	);
	LUT4 #(
		.INIT('h1311)
	) name3597 (
		_w2182_,
		_w4044_,
		_w4049_,
		_w4059_,
		_w4060_
	);
	LUT2 #(
		.INIT('h2)
	) name3598 (
		\P1_reg3_reg[14]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4061_
	);
	LUT3 #(
		.INIT('h07)
	) name3599 (
		_w835_,
		_w1244_,
		_w4061_,
		_w4062_
	);
	LUT3 #(
		.INIT('h2f)
	) name3600 (
		\P1_state_reg[0]/NET0131 ,
		_w4060_,
		_w4062_,
		_w4063_
	);
	LUT2 #(
		.INIT('h8)
	) name3601 (
		_w825_,
		_w2183_,
		_w4064_
	);
	LUT4 #(
		.INIT('h2220)
	) name3602 (
		_w825_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4065_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3603 (
		_w2962_,
		_w2963_,
		_w2965_,
		_w2970_,
		_w4066_
	);
	LUT4 #(
		.INIT('h070b)
	) name3604 (
		_w1168_,
		_w2055_,
		_w4065_,
		_w4066_,
		_w4067_
	);
	LUT2 #(
		.INIT('h2)
	) name3605 (
		_w2121_,
		_w4067_,
		_w4068_
	);
	LUT4 #(
		.INIT('h9a55)
	) name3606 (
		_w1168_,
		_w2938_,
		_w2939_,
		_w2940_,
		_w4069_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3607 (
		_w825_,
		_w2055_,
		_w2128_,
		_w4069_,
		_w4070_
	);
	LUT4 #(
		.INIT('h6555)
	) name3608 (
		_w764_,
		_w889_,
		_w2134_,
		_w2137_,
		_w4071_
	);
	LUT4 #(
		.INIT('h7020)
	) name3609 (
		_w488_,
		_w837_,
		_w2055_,
		_w4071_,
		_w4072_
	);
	LUT3 #(
		.INIT('ha8)
	) name3610 (
		_w1237_,
		_w4065_,
		_w4072_,
		_w4073_
	);
	LUT4 #(
		.INIT('h0e0a)
	) name3611 (
		_w833_,
		_w842_,
		_w2163_,
		_w2859_,
		_w4074_
	);
	LUT4 #(
		.INIT('he020)
	) name3612 (
		_w825_,
		_w2055_,
		_w2170_,
		_w4074_,
		_w4075_
	);
	LUT3 #(
		.INIT('h10)
	) name3613 (
		_w833_,
		_w2175_,
		_w2176_,
		_w4076_
	);
	LUT3 #(
		.INIT('ha8)
	) name3614 (
		_w825_,
		_w2171_,
		_w2578_,
		_w4077_
	);
	LUT2 #(
		.INIT('h1)
	) name3615 (
		_w4076_,
		_w4077_,
		_w4078_
	);
	LUT2 #(
		.INIT('h4)
	) name3616 (
		_w4075_,
		_w4078_,
		_w4079_
	);
	LUT3 #(
		.INIT('h10)
	) name3617 (
		_w4073_,
		_w4070_,
		_w4079_,
		_w4080_
	);
	LUT4 #(
		.INIT('h1311)
	) name3618 (
		_w2182_,
		_w4064_,
		_w4068_,
		_w4080_,
		_w4081_
	);
	LUT2 #(
		.INIT('h2)
	) name3619 (
		\P1_reg3_reg[15]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4082_
	);
	LUT3 #(
		.INIT('h07)
	) name3620 (
		_w825_,
		_w1244_,
		_w4082_,
		_w4083_
	);
	LUT3 #(
		.INIT('h2f)
	) name3621 (
		\P1_state_reg[0]/NET0131 ,
		_w4081_,
		_w4083_,
		_w4084_
	);
	LUT4 #(
		.INIT('h4000)
	) name3622 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1762_,
		_w4085_
	);
	LUT2 #(
		.INIT('h2)
	) name3623 (
		_w1762_,
		_w2903_,
		_w4086_
	);
	LUT4 #(
		.INIT('h1000)
	) name3624 (
		_w1740_,
		_w1764_,
		_w1972_,
		_w1973_,
		_w4087_
	);
	LUT4 #(
		.INIT('h6555)
	) name3625 (
		_w1740_,
		_w1764_,
		_w1972_,
		_w1973_,
		_w4088_
	);
	LUT4 #(
		.INIT('h7020)
	) name3626 (
		_w1305_,
		_w1779_,
		_w2903_,
		_w4088_,
		_w4089_
	);
	LUT3 #(
		.INIT('ha8)
	) name3627 (
		_w2000_,
		_w4086_,
		_w4089_,
		_w4090_
	);
	LUT4 #(
		.INIT('h31ce)
	) name3628 (
		_w2414_,
		_w2400_,
		_w2413_,
		_w2483_,
		_w4091_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3629 (
		_w1762_,
		_w1963_,
		_w2903_,
		_w4091_,
		_w4092_
	);
	LUT4 #(
		.INIT('h007b)
	) name3630 (
		_w2483_,
		_w2903_,
		_w3095_,
		_w4086_,
		_w4093_
	);
	LUT4 #(
		.INIT('h0100)
	) name3631 (
		_w1695_,
		_w1706_,
		_w1788_,
		_w2005_,
		_w4094_
	);
	LUT4 #(
		.INIT('h8040)
	) name3632 (
		_w1774_,
		_w2025_,
		_w2903_,
		_w4094_,
		_w4095_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3633 (
		_w1762_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w4096_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3634 (
		_w1774_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w4097_
	);
	LUT2 #(
		.INIT('h1)
	) name3635 (
		_w4096_,
		_w4097_,
		_w4098_
	);
	LUT2 #(
		.INIT('h4)
	) name3636 (
		_w4095_,
		_w4098_,
		_w4099_
	);
	LUT3 #(
		.INIT('hd0)
	) name3637 (
		_w1869_,
		_w4093_,
		_w4099_,
		_w4100_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3638 (
		_w1285_,
		_w4092_,
		_w4090_,
		_w4100_,
		_w4101_
	);
	LUT2 #(
		.INIT('h4)
	) name3639 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[10]/NET0131 ,
		_w4102_
	);
	LUT3 #(
		.INIT('h07)
	) name3640 (
		_w1762_,
		_w2344_,
		_w4102_,
		_w4103_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3641 (
		\P1_state_reg[0]/NET0131 ,
		_w4085_,
		_w4101_,
		_w4103_,
		_w4104_
	);
	LUT4 #(
		.INIT('h4000)
	) name3642 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1831_,
		_w4105_
	);
	LUT2 #(
		.INIT('h2)
	) name3643 (
		_w1831_,
		_w2903_,
		_w4106_
	);
	LUT4 #(
		.INIT('h4144)
	) name3644 (
		_w1305_,
		_w1825_,
		_w1834_,
		_w1976_,
		_w4107_
	);
	LUT3 #(
		.INIT('h80)
	) name3645 (
		_w1305_,
		_w1750_,
		_w1751_,
		_w4108_
	);
	LUT4 #(
		.INIT('h3331)
	) name3646 (
		_w2903_,
		_w4106_,
		_w4107_,
		_w4108_,
		_w4109_
	);
	LUT2 #(
		.INIT('h2)
	) name3647 (
		_w2000_,
		_w4109_,
		_w4110_
	);
	LUT2 #(
		.INIT('h9)
	) name3648 (
		_w1834_,
		_w1839_,
		_w4111_
	);
	LUT4 #(
		.INIT('h40b0)
	) name3649 (
		_w1792_,
		_w1797_,
		_w2903_,
		_w4111_,
		_w4112_
	);
	LUT3 #(
		.INIT('ha8)
	) name3650 (
		_w1869_,
		_w4106_,
		_w4112_,
		_w4113_
	);
	LUT4 #(
		.INIT('h8a75)
	) name3651 (
		_w1878_,
		_w1905_,
		_w1908_,
		_w4111_,
		_w4114_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3652 (
		_w1831_,
		_w1963_,
		_w2903_,
		_w4114_,
		_w4115_
	);
	LUT4 #(
		.INIT('h1033)
	) name3653 (
		_w1759_,
		_w1839_,
		_w2009_,
		_w2025_,
		_w4116_
	);
	LUT4 #(
		.INIT('h0023)
	) name3654 (
		_w1306_,
		_w1837_,
		_w1838_,
		_w2001_,
		_w4117_
	);
	LUT4 #(
		.INIT('hbf00)
	) name3655 (
		_w1759_,
		_w2009_,
		_w2025_,
		_w4117_,
		_w4118_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3656 (
		_w1831_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w4119_
	);
	LUT4 #(
		.INIT('h2300)
	) name3657 (
		_w1306_,
		_w1837_,
		_w1838_,
		_w2029_,
		_w4120_
	);
	LUT2 #(
		.INIT('h1)
	) name3658 (
		_w4119_,
		_w4120_,
		_w4121_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3659 (
		_w2903_,
		_w4116_,
		_w4118_,
		_w4121_,
		_w4122_
	);
	LUT3 #(
		.INIT('h10)
	) name3660 (
		_w4115_,
		_w4113_,
		_w4122_,
		_w4123_
	);
	LUT4 #(
		.INIT('h1311)
	) name3661 (
		_w1285_,
		_w4105_,
		_w4110_,
		_w4123_,
		_w4124_
	);
	LUT2 #(
		.INIT('h4)
	) name3662 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[13]/NET0131 ,
		_w4125_
	);
	LUT3 #(
		.INIT('h07)
	) name3663 (
		_w1831_,
		_w2344_,
		_w4125_,
		_w4126_
	);
	LUT3 #(
		.INIT('h2f)
	) name3664 (
		\P1_state_reg[0]/NET0131 ,
		_w4124_,
		_w4126_,
		_w4127_
	);
	LUT4 #(
		.INIT('h4000)
	) name3665 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1810_,
		_w4128_
	);
	LUT2 #(
		.INIT('h2)
	) name3666 (
		_w1810_,
		_w2903_,
		_w4129_
	);
	LUT4 #(
		.INIT('h4144)
	) name3667 (
		_w1305_,
		_w1807_,
		_w1812_,
		_w1978_,
		_w4130_
	);
	LUT3 #(
		.INIT('h80)
	) name3668 (
		_w1305_,
		_w1822_,
		_w1824_,
		_w4131_
	);
	LUT4 #(
		.INIT('h3331)
	) name3669 (
		_w2903_,
		_w4129_,
		_w4130_,
		_w4131_,
		_w4132_
	);
	LUT2 #(
		.INIT('h2)
	) name3670 (
		_w2000_,
		_w4132_,
		_w4133_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3671 (
		_w2614_,
		_w2615_,
		_w2617_,
		_w2619_,
		_w4134_
	);
	LUT4 #(
		.INIT('h070b)
	) name3672 (
		_w2493_,
		_w2903_,
		_w4129_,
		_w4134_,
		_w4135_
	);
	LUT4 #(
		.INIT('h9a55)
	) name3673 (
		_w2493_,
		_w2593_,
		_w2594_,
		_w2595_,
		_w4136_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3674 (
		_w1810_,
		_w1963_,
		_w2903_,
		_w4136_,
		_w4137_
	);
	LUT4 #(
		.INIT('h8040)
	) name3675 (
		_w1820_,
		_w2025_,
		_w2903_,
		_w3716_,
		_w4138_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3676 (
		_w1810_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w4139_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3677 (
		_w1820_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w4140_
	);
	LUT2 #(
		.INIT('h1)
	) name3678 (
		_w4139_,
		_w4140_,
		_w4141_
	);
	LUT2 #(
		.INIT('h4)
	) name3679 (
		_w4138_,
		_w4141_,
		_w4142_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3680 (
		_w1869_,
		_w4135_,
		_w4137_,
		_w4142_,
		_w4143_
	);
	LUT4 #(
		.INIT('h1311)
	) name3681 (
		_w1285_,
		_w4128_,
		_w4133_,
		_w4143_,
		_w4144_
	);
	LUT2 #(
		.INIT('h4)
	) name3682 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[15]/NET0131 ,
		_w4145_
	);
	LUT3 #(
		.INIT('h07)
	) name3683 (
		_w1810_,
		_w2344_,
		_w4145_,
		_w4146_
	);
	LUT3 #(
		.INIT('h2f)
	) name3684 (
		\P1_state_reg[0]/NET0131 ,
		_w4144_,
		_w4146_,
		_w4147_
	);
	LUT4 #(
		.INIT('h4000)
	) name3685 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1776_,
		_w4148_
	);
	LUT2 #(
		.INIT('h2)
	) name3686 (
		_w1776_,
		_w2903_,
		_w4149_
	);
	LUT4 #(
		.INIT('h1444)
	) name3687 (
		_w1305_,
		_w1764_,
		_w1972_,
		_w1973_,
		_w4150_
	);
	LUT3 #(
		.INIT('h80)
	) name3688 (
		_w1305_,
		_w1688_,
		_w1690_,
		_w4151_
	);
	LUT4 #(
		.INIT('h3331)
	) name3689 (
		_w2903_,
		_w4149_,
		_w4150_,
		_w4151_,
		_w4152_
	);
	LUT2 #(
		.INIT('h2)
	) name3690 (
		_w2000_,
		_w4152_,
		_w4153_
	);
	LUT4 #(
		.INIT('h009f)
	) name3691 (
		_w1905_,
		_w2484_,
		_w2903_,
		_w4149_,
		_w4154_
	);
	LUT4 #(
		.INIT('hb04f)
	) name3692 (
		_w1687_,
		_w1729_,
		_w1736_,
		_w2484_,
		_w4155_
	);
	LUT4 #(
		.INIT('hc808)
	) name3693 (
		_w1776_,
		_w1869_,
		_w2903_,
		_w4155_,
		_w4156_
	);
	LUT3 #(
		.INIT('h10)
	) name3694 (
		_w1783_,
		_w1787_,
		_w2001_,
		_w4157_
	);
	LUT4 #(
		.INIT('h006f)
	) name3695 (
		_w1788_,
		_w2006_,
		_w2025_,
		_w4157_,
		_w4158_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3696 (
		_w1776_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w4159_
	);
	LUT3 #(
		.INIT('h10)
	) name3697 (
		_w1783_,
		_w1787_,
		_w2029_,
		_w4160_
	);
	LUT2 #(
		.INIT('h1)
	) name3698 (
		_w4159_,
		_w4160_,
		_w4161_
	);
	LUT3 #(
		.INIT('hd0)
	) name3699 (
		_w2903_,
		_w4158_,
		_w4161_,
		_w4162_
	);
	LUT4 #(
		.INIT('h3100)
	) name3700 (
		_w1963_,
		_w4156_,
		_w4154_,
		_w4162_,
		_w4163_
	);
	LUT4 #(
		.INIT('h1311)
	) name3701 (
		_w1285_,
		_w4148_,
		_w4153_,
		_w4163_,
		_w4164_
	);
	LUT2 #(
		.INIT('h4)
	) name3702 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[9]/NET0131 ,
		_w4165_
	);
	LUT3 #(
		.INIT('h07)
	) name3703 (
		_w1776_,
		_w2344_,
		_w4165_,
		_w4166_
	);
	LUT3 #(
		.INIT('h2f)
	) name3704 (
		\P1_state_reg[0]/NET0131 ,
		_w4164_,
		_w4166_,
		_w4167_
	);
	LUT2 #(
		.INIT('h8)
	) name3705 (
		_w908_,
		_w2183_,
		_w4168_
	);
	LUT4 #(
		.INIT('h0100)
	) name3706 (
		_w949_,
		_w961_,
		_w971_,
		_w2130_,
		_w4169_
	);
	LUT4 #(
		.INIT('h0100)
	) name3707 (
		_w911_,
		_w927_,
		_w938_,
		_w4169_,
		_w4170_
	);
	LUT3 #(
		.INIT('h15)
	) name3708 (
		_w488_,
		_w896_,
		_w898_,
		_w4171_
	);
	LUT3 #(
		.INIT('h2a)
	) name3709 (
		_w488_,
		_w935_,
		_w937_,
		_w4172_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3710 (
		_w2134_,
		_w4170_,
		_w4171_,
		_w4172_,
		_w4173_
	);
	LUT3 #(
		.INIT('h60)
	) name3711 (
		_w915_,
		_w2159_,
		_w2170_,
		_w4174_
	);
	LUT4 #(
		.INIT('h006f)
	) name3712 (
		_w1015_,
		_w1191_,
		_w2128_,
		_w4174_,
		_w4175_
	);
	LUT4 #(
		.INIT('h08cc)
	) name3713 (
		_w1237_,
		_w2055_,
		_w4173_,
		_w4175_,
		_w4176_
	);
	LUT4 #(
		.INIT('h1110)
	) name3714 (
		_w908_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4177_
	);
	LUT2 #(
		.INIT('h2)
	) name3715 (
		_w2121_,
		_w4177_,
		_w4178_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3716 (
		_w1191_,
		_w2055_,
		_w2082_,
		_w4178_,
		_w4179_
	);
	LUT3 #(
		.INIT('h10)
	) name3717 (
		_w915_,
		_w2175_,
		_w2176_,
		_w4180_
	);
	LUT4 #(
		.INIT('h0001)
	) name3718 (
		_w2171_,
		_w2173_,
		_w2845_,
		_w3791_,
		_w4181_
	);
	LUT3 #(
		.INIT('h31)
	) name3719 (
		_w908_,
		_w4180_,
		_w4181_,
		_w4182_
	);
	LUT2 #(
		.INIT('h4)
	) name3720 (
		_w4179_,
		_w4182_,
		_w4183_
	);
	LUT4 #(
		.INIT('h1311)
	) name3721 (
		_w2182_,
		_w4168_,
		_w4176_,
		_w4183_,
		_w4184_
	);
	LUT2 #(
		.INIT('h2)
	) name3722 (
		\P1_reg3_reg[8]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4185_
	);
	LUT4 #(
		.INIT('h4080)
	) name3723 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w908_,
		_w1242_,
		_w4186_
	);
	LUT2 #(
		.INIT('h1)
	) name3724 (
		_w4185_,
		_w4186_,
		_w4187_
	);
	LUT3 #(
		.INIT('h2f)
	) name3725 (
		\P1_state_reg[0]/NET0131 ,
		_w4184_,
		_w4187_,
		_w4188_
	);
	LUT3 #(
		.INIT('h02)
	) name3726 (
		_w2025_,
		_w3934_,
		_w3935_,
		_w4189_
	);
	LUT3 #(
		.INIT('h02)
	) name3727 (
		_w2000_,
		_w3938_,
		_w3939_,
		_w4190_
	);
	LUT4 #(
		.INIT('h0070)
	) name3728 (
		_w1963_,
		_w3932_,
		_w3943_,
		_w4190_,
		_w4191_
	);
	LUT3 #(
		.INIT('h10)
	) name3729 (
		_w1306_,
		_w1586_,
		_w2029_,
		_w4192_
	);
	LUT4 #(
		.INIT('h0075)
	) name3730 (
		_w2903_,
		_w4189_,
		_w4191_,
		_w4192_,
		_w4193_
	);
	LUT3 #(
		.INIT('h45)
	) name3731 (
		_w2029_,
		_w2032_,
		_w2903_,
		_w4194_
	);
	LUT4 #(
		.INIT('h1011)
	) name3732 (
		_w1963_,
		_w2029_,
		_w2032_,
		_w2903_,
		_w4195_
	);
	LUT3 #(
		.INIT('h51)
	) name3733 (
		_w1284_,
		_w1963_,
		_w2903_,
		_w4196_
	);
	LUT3 #(
		.INIT('h12)
	) name3734 (
		\P2_reg3_reg[20]/NET0131 ,
		_w1267_,
		_w1535_,
		_w4197_
	);
	LUT3 #(
		.INIT('hb0)
	) name3735 (
		_w4195_,
		_w4196_,
		_w4197_,
		_w4198_
	);
	LUT4 #(
		.INIT('haa08)
	) name3736 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w4193_,
		_w4198_,
		_w4199_
	);
	LUT4 #(
		.INIT('h9b3b)
	) name3737 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[20]/NET0131 ,
		_w1267_,
		_w1535_,
		_w4200_
	);
	LUT2 #(
		.INIT('hb)
	) name3738 (
		_w4199_,
		_w4200_,
		_w4201_
	);
	LUT4 #(
		.INIT('h2220)
	) name3739 (
		_w786_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4202_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3740 (
		_w2942_,
		_w2943_,
		_w2945_,
		_w2948_,
		_w4203_
	);
	LUT4 #(
		.INIT('h0b07)
	) name3741 (
		_w1213_,
		_w2055_,
		_w4202_,
		_w4203_,
		_w4204_
	);
	LUT2 #(
		.INIT('h8)
	) name3742 (
		_w2959_,
		_w2964_,
		_w4205_
	);
	LUT4 #(
		.INIT('h00a2)
	) name3743 (
		_w2304_,
		_w2959_,
		_w2971_,
		_w2968_,
		_w4206_
	);
	LUT4 #(
		.INIT('h65aa)
	) name3744 (
		_w1213_,
		_w4066_,
		_w4205_,
		_w4206_,
		_w4207_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3745 (
		_w786_,
		_w2055_,
		_w2121_,
		_w4207_,
		_w4208_
	);
	LUT4 #(
		.INIT('h1444)
	) name3746 (
		_w488_,
		_w1079_,
		_w2142_,
		_w2213_,
		_w4209_
	);
	LUT2 #(
		.INIT('h8)
	) name3747 (
		_w488_,
		_w780_,
		_w4210_
	);
	LUT4 #(
		.INIT('h3331)
	) name3748 (
		_w2055_,
		_w4202_,
		_w4209_,
		_w4210_,
		_w4211_
	);
	LUT4 #(
		.INIT('h8040)
	) name3749 (
		_w784_,
		_w2055_,
		_w2170_,
		_w2860_,
		_w4212_
	);
	LUT3 #(
		.INIT('ha8)
	) name3750 (
		_w786_,
		_w2171_,
		_w2173_,
		_w4213_
	);
	LUT4 #(
		.INIT('h0100)
	) name3751 (
		_w489_,
		_w783_,
		_w2175_,
		_w2176_,
		_w4214_
	);
	LUT2 #(
		.INIT('h1)
	) name3752 (
		_w4213_,
		_w4214_,
		_w4215_
	);
	LUT2 #(
		.INIT('h4)
	) name3753 (
		_w4212_,
		_w4215_,
		_w4216_
	);
	LUT3 #(
		.INIT('hd0)
	) name3754 (
		_w1237_,
		_w4211_,
		_w4216_,
		_w4217_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3755 (
		_w2128_,
		_w4204_,
		_w4208_,
		_w4217_,
		_w4218_
	);
	LUT2 #(
		.INIT('h8)
	) name3756 (
		_w786_,
		_w2183_,
		_w4219_
	);
	LUT4 #(
		.INIT('haa08)
	) name3757 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w4218_,
		_w4219_,
		_w4220_
	);
	LUT2 #(
		.INIT('h2)
	) name3758 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4221_
	);
	LUT3 #(
		.INIT('h07)
	) name3759 (
		_w786_,
		_w1244_,
		_w4221_,
		_w4222_
	);
	LUT2 #(
		.INIT('hb)
	) name3760 (
		_w4220_,
		_w4222_,
		_w4223_
	);
	LUT2 #(
		.INIT('h8)
	) name3761 (
		_w1570_,
		_w2039_,
		_w4224_
	);
	LUT2 #(
		.INIT('h2)
	) name3762 (
		_w1570_,
		_w2903_,
		_w4225_
	);
	LUT4 #(
		.INIT('h4b00)
	) name3763 (
		_w1842_,
		_w1852_,
		_w2509_,
		_w2903_,
		_w4226_
	);
	LUT3 #(
		.INIT('ha8)
	) name3764 (
		_w1869_,
		_w4225_,
		_w4226_,
		_w4227_
	);
	LUT4 #(
		.INIT('hb400)
	) name3765 (
		_w1918_,
		_w1932_,
		_w2509_,
		_w2903_,
		_w4228_
	);
	LUT3 #(
		.INIT('ha8)
	) name3766 (
		_w1963_,
		_w4225_,
		_w4228_,
		_w4229_
	);
	LUT4 #(
		.INIT('h1444)
	) name3767 (
		_w1305_,
		_w1564_,
		_w1978_,
		_w1983_,
		_w4230_
	);
	LUT4 #(
		.INIT('h0200)
	) name3768 (
		_w1305_,
		_w1590_,
		_w1589_,
		_w1591_,
		_w4231_
	);
	LUT4 #(
		.INIT('h3331)
	) name3769 (
		_w2903_,
		_w4225_,
		_w4230_,
		_w4231_,
		_w4232_
	);
	LUT4 #(
		.INIT('h9050)
	) name3770 (
		_w1569_,
		_w2012_,
		_w2903_,
		_w3402_,
		_w4233_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3771 (
		_w1570_,
		_w2001_,
		_w2032_,
		_w2903_,
		_w4234_
	);
	LUT3 #(
		.INIT('h0d)
	) name3772 (
		_w1569_,
		_w2993_,
		_w4234_,
		_w4235_
	);
	LUT4 #(
		.INIT('h5700)
	) name3773 (
		_w2025_,
		_w4225_,
		_w4233_,
		_w4235_,
		_w4236_
	);
	LUT3 #(
		.INIT('hd0)
	) name3774 (
		_w2000_,
		_w4232_,
		_w4236_,
		_w4237_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3775 (
		_w1285_,
		_w4227_,
		_w4229_,
		_w4237_,
		_w4238_
	);
	LUT2 #(
		.INIT('h4)
	) name3776 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[21]/NET0131 ,
		_w4239_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3777 (
		\P2_reg3_reg[20]/NET0131 ,
		\P2_reg3_reg[21]/NET0131 ,
		_w1535_,
		_w2344_,
		_w4240_
	);
	LUT2 #(
		.INIT('h1)
	) name3778 (
		_w4239_,
		_w4240_,
		_w4241_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3779 (
		\P1_state_reg[0]/NET0131 ,
		_w4224_,
		_w4238_,
		_w4241_,
		_w4242_
	);
	LUT2 #(
		.INIT('h8)
	) name3780 (
		_w1548_,
		_w2039_,
		_w4243_
	);
	LUT2 #(
		.INIT('h2)
	) name3781 (
		_w1548_,
		_w2903_,
		_w4244_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3782 (
		_w2597_,
		_w2598_,
		_w2599_,
		_w2601_,
		_w4245_
	);
	LUT4 #(
		.INIT('h0b07)
	) name3783 (
		_w2505_,
		_w2903_,
		_w4244_,
		_w4245_,
		_w4246_
	);
	LUT2 #(
		.INIT('h8)
	) name3784 (
		_w2616_,
		_w2623_,
		_w4247_
	);
	LUT2 #(
		.INIT('h4)
	) name3785 (
		_w2620_,
		_w2623_,
		_w4248_
	);
	LUT2 #(
		.INIT('h2)
	) name3786 (
		_w2606_,
		_w4248_,
		_w4249_
	);
	LUT4 #(
		.INIT('h65aa)
	) name3787 (
		_w2505_,
		_w4134_,
		_w4247_,
		_w4249_,
		_w4250_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3788 (
		_w1548_,
		_w1869_,
		_w2903_,
		_w4250_,
		_w4251_
	);
	LUT4 #(
		.INIT('h1444)
	) name3789 (
		_w1305_,
		_w1542_,
		_w1978_,
		_w1985_,
		_w4252_
	);
	LUT2 #(
		.INIT('h8)
	) name3790 (
		_w1305_,
		_w1564_,
		_w4253_
	);
	LUT4 #(
		.INIT('h3331)
	) name3791 (
		_w2903_,
		_w4244_,
		_w4252_,
		_w4253_,
		_w4254_
	);
	LUT3 #(
		.INIT('h8a)
	) name3792 (
		_w1547_,
		_w1560_,
		_w3503_,
		_w4255_
	);
	LUT2 #(
		.INIT('h2)
	) name3793 (
		_w2025_,
		_w2890_,
		_w4256_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3794 (
		_w1548_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w4257_
	);
	LUT3 #(
		.INIT('h0d)
	) name3795 (
		_w1547_,
		_w2993_,
		_w4257_,
		_w4258_
	);
	LUT4 #(
		.INIT('hdf00)
	) name3796 (
		_w2903_,
		_w4255_,
		_w4256_,
		_w4258_,
		_w4259_
	);
	LUT3 #(
		.INIT('hd0)
	) name3797 (
		_w2000_,
		_w4254_,
		_w4259_,
		_w4260_
	);
	LUT4 #(
		.INIT('h3100)
	) name3798 (
		_w1963_,
		_w4251_,
		_w4246_,
		_w4260_,
		_w4261_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3799 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w4243_,
		_w4261_,
		_w4262_
	);
	LUT2 #(
		.INIT('h4)
	) name3800 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		_w4263_
	);
	LUT3 #(
		.INIT('h07)
	) name3801 (
		_w1548_,
		_w2344_,
		_w4263_,
		_w4264_
	);
	LUT2 #(
		.INIT('hb)
	) name3802 (
		_w4262_,
		_w4264_,
		_w4265_
	);
	LUT2 #(
		.INIT('h2)
	) name3803 (
		\P2_reg0_reg[21]/NET0131 ,
		_w2042_,
		_w4266_
	);
	LUT4 #(
		.INIT('h2000)
	) name3804 (
		\P2_reg0_reg[21]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4267_
	);
	LUT2 #(
		.INIT('h2)
	) name3805 (
		\P2_reg0_reg[21]/NET0131 ,
		_w2729_,
		_w4268_
	);
	LUT4 #(
		.INIT('h4b00)
	) name3806 (
		_w1842_,
		_w1852_,
		_w2509_,
		_w2729_,
		_w4269_
	);
	LUT3 #(
		.INIT('ha8)
	) name3807 (
		_w1869_,
		_w4268_,
		_w4269_,
		_w4270_
	);
	LUT4 #(
		.INIT('hb400)
	) name3808 (
		_w1918_,
		_w1932_,
		_w2509_,
		_w2729_,
		_w4271_
	);
	LUT3 #(
		.INIT('ha8)
	) name3809 (
		_w1963_,
		_w4268_,
		_w4271_,
		_w4272_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3810 (
		\P2_reg0_reg[21]/NET0131 ,
		_w2729_,
		_w4230_,
		_w4231_,
		_w4273_
	);
	LUT2 #(
		.INIT('h2)
	) name3811 (
		\P2_reg0_reg[21]/NET0131 ,
		_w3084_,
		_w4274_
	);
	LUT3 #(
		.INIT('h10)
	) name3812 (
		_w1306_,
		_w1568_,
		_w2001_,
		_w4275_
	);
	LUT4 #(
		.INIT('h9050)
	) name3813 (
		_w1569_,
		_w2012_,
		_w2025_,
		_w3402_,
		_w4276_
	);
	LUT4 #(
		.INIT('h1113)
	) name3814 (
		_w2729_,
		_w4274_,
		_w4275_,
		_w4276_,
		_w4277_
	);
	LUT3 #(
		.INIT('hd0)
	) name3815 (
		_w2000_,
		_w4273_,
		_w4277_,
		_w4278_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3816 (
		_w1285_,
		_w4270_,
		_w4272_,
		_w4278_,
		_w4279_
	);
	LUT4 #(
		.INIT('heeec)
	) name3817 (
		\P1_state_reg[0]/NET0131 ,
		_w4266_,
		_w4267_,
		_w4279_,
		_w4280_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3818 (
		\P1_reg1_reg[8]/NET0131 ,
		_w2820_,
		_w3511_,
		_w3606_,
		_w4281_
	);
	LUT2 #(
		.INIT('h4)
	) name3819 (
		_w915_,
		_w2194_,
		_w4282_
	);
	LUT4 #(
		.INIT('h009f)
	) name3820 (
		_w1191_,
		_w2082_,
		_w2121_,
		_w4282_,
		_w4283_
	);
	LUT4 #(
		.INIT('hd000)
	) name3821 (
		_w1237_,
		_w4173_,
		_w4175_,
		_w4283_,
		_w4284_
	);
	LUT3 #(
		.INIT('hce)
	) name3822 (
		_w3608_,
		_w4281_,
		_w4284_,
		_w4285_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name3823 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[9]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4286_
	);
	LUT2 #(
		.INIT('h8)
	) name3824 (
		\P1_reg1_reg[9]/NET0131 ,
		_w2183_,
		_w4287_
	);
	LUT4 #(
		.INIT('hc808)
	) name3825 (
		\P1_reg1_reg[9]/NET0131 ,
		_w1237_,
		_w2536_,
		_w3733_,
		_w4288_
	);
	LUT4 #(
		.INIT('hc808)
	) name3826 (
		\P1_reg1_reg[9]/NET0131 ,
		_w2121_,
		_w2536_,
		_w3735_,
		_w4289_
	);
	LUT2 #(
		.INIT('h2)
	) name3827 (
		\P1_reg1_reg[9]/NET0131 ,
		_w3606_,
		_w4290_
	);
	LUT4 #(
		.INIT('h8488)
	) name3828 (
		_w1173_,
		_w2128_,
		_w2236_,
		_w2239_,
		_w4291_
	);
	LUT2 #(
		.INIT('h4)
	) name3829 (
		_w905_,
		_w2194_,
		_w4292_
	);
	LUT2 #(
		.INIT('h1)
	) name3830 (
		_w3738_,
		_w4292_,
		_w4293_
	);
	LUT4 #(
		.INIT('h1311)
	) name3831 (
		_w2536_,
		_w4290_,
		_w4291_,
		_w4293_,
		_w4294_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3832 (
		_w2182_,
		_w4289_,
		_w4288_,
		_w4294_,
		_w4295_
	);
	LUT4 #(
		.INIT('heeec)
	) name3833 (
		\P1_state_reg[0]/NET0131 ,
		_w4286_,
		_w4287_,
		_w4295_,
		_w4296_
	);
	LUT3 #(
		.INIT('h04)
	) name3834 (
		_w1306_,
		_w2001_,
		_w2362_,
		_w4297_
	);
	LUT4 #(
		.INIT('h00bf)
	) name3835 (
		_w1995_,
		_w1997_,
		_w2553_,
		_w4297_,
		_w4298_
	);
	LUT3 #(
		.INIT('hc8)
	) name3836 (
		\P2_reg0_reg[30]/NET0131 ,
		_w2025_,
		_w2729_,
		_w4299_
	);
	LUT4 #(
		.INIT('h9f00)
	) name3837 (
		_w2022_,
		_w2363_,
		_w2729_,
		_w4299_,
		_w4300_
	);
	LUT4 #(
		.INIT('haa08)
	) name3838 (
		_w2556_,
		_w2729_,
		_w4298_,
		_w4300_,
		_w4301_
	);
	LUT3 #(
		.INIT('ha8)
	) name3839 (
		_w2556_,
		_w2729_,
		_w3266_,
		_w4302_
	);
	LUT3 #(
		.INIT('h2a)
	) name3840 (
		\P2_reg0_reg[30]/NET0131 ,
		_w3082_,
		_w4302_,
		_w4303_
	);
	LUT2 #(
		.INIT('he)
	) name3841 (
		_w4301_,
		_w4303_,
		_w4304_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name3842 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[19]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4305_
	);
	LUT2 #(
		.INIT('h8)
	) name3843 (
		\P1_reg2_reg[19]/NET0131 ,
		_w2183_,
		_w4306_
	);
	LUT4 #(
		.INIT('haa8a)
	) name3844 (
		\P1_reg2_reg[19]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4307_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3845 (
		\P1_reg2_reg[19]/NET0131 ,
		_w2189_,
		_w3671_,
		_w3672_,
		_w4308_
	);
	LUT2 #(
		.INIT('h2)
	) name3846 (
		_w1237_,
		_w4308_,
		_w4309_
	);
	LUT4 #(
		.INIT('h4844)
	) name3847 (
		_w1217_,
		_w2189_,
		_w2942_,
		_w2943_,
		_w4310_
	);
	LUT3 #(
		.INIT('ha8)
	) name3848 (
		_w2128_,
		_w4307_,
		_w4310_,
		_w4311_
	);
	LUT4 #(
		.INIT('hc535)
	) name3849 (
		\P1_reg2_reg[19]/NET0131 ,
		_w1217_,
		_w2189_,
		_w3677_,
		_w4312_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3850 (
		\P1_reg2_reg[19]/NET0131 ,
		_w2189_,
		_w3168_,
		_w3680_,
		_w4313_
	);
	LUT4 #(
		.INIT('hf100)
	) name3851 (
		_w489_,
		_w717_,
		_w719_,
		_w2194_,
		_w4314_
	);
	LUT2 #(
		.INIT('h8)
	) name3852 (
		_w721_,
		_w1120_,
		_w4315_
	);
	LUT4 #(
		.INIT('h0057)
	) name3853 (
		\P1_reg2_reg[19]/NET0131 ,
		_w2171_,
		_w2196_,
		_w4315_,
		_w4316_
	);
	LUT3 #(
		.INIT('h70)
	) name3854 (
		_w2189_,
		_w4314_,
		_w4316_,
		_w4317_
	);
	LUT3 #(
		.INIT('hd0)
	) name3855 (
		_w2170_,
		_w4313_,
		_w4317_,
		_w4318_
	);
	LUT3 #(
		.INIT('hd0)
	) name3856 (
		_w2121_,
		_w4312_,
		_w4318_,
		_w4319_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3857 (
		_w2182_,
		_w4311_,
		_w4309_,
		_w4319_,
		_w4320_
	);
	LUT4 #(
		.INIT('heeec)
	) name3858 (
		\P1_state_reg[0]/NET0131 ,
		_w4305_,
		_w4306_,
		_w4320_,
		_w4321_
	);
	LUT2 #(
		.INIT('h2)
	) name3859 (
		\P2_reg1_reg[12]/NET0131 ,
		_w2762_,
		_w4322_
	);
	LUT4 #(
		.INIT('hc535)
	) name3860 (
		\P2_reg1_reg[12]/NET0131 ,
		_w2494_,
		_w2762_,
		_w3003_,
		_w4323_
	);
	LUT4 #(
		.INIT('h7020)
	) name3861 (
		_w1305_,
		_w1740_,
		_w2762_,
		_w3693_,
		_w4324_
	);
	LUT3 #(
		.INIT('ha8)
	) name3862 (
		_w2000_,
		_w4322_,
		_w4324_,
		_w4325_
	);
	LUT4 #(
		.INIT('h2300)
	) name3863 (
		_w1306_,
		_w1756_,
		_w1758_,
		_w2001_,
		_w4326_
	);
	LUT4 #(
		.INIT('h006f)
	) name3864 (
		_w1759_,
		_w2009_,
		_w2025_,
		_w4326_,
		_w4327_
	);
	LUT4 #(
		.INIT('h7d00)
	) name3865 (
		_w1869_,
		_w2494_,
		_w3025_,
		_w4327_,
		_w4328_
	);
	LUT3 #(
		.INIT('ha2)
	) name3866 (
		\P2_reg1_reg[12]/NET0131 ,
		_w3225_,
		_w3874_,
		_w4329_
	);
	LUT3 #(
		.INIT('h0d)
	) name3867 (
		_w2762_,
		_w4328_,
		_w4329_,
		_w4330_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3868 (
		_w1963_,
		_w4323_,
		_w4325_,
		_w4330_,
		_w4331_
	);
	LUT4 #(
		.INIT('h2000)
	) name3869 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4332_
	);
	LUT4 #(
		.INIT('haa08)
	) name3870 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w4331_,
		_w4332_,
		_w4333_
	);
	LUT2 #(
		.INIT('h2)
	) name3871 (
		\P2_reg1_reg[12]/NET0131 ,
		_w2042_,
		_w4334_
	);
	LUT2 #(
		.INIT('he)
	) name3872 (
		_w4333_,
		_w4334_,
		_w4335_
	);
	LUT2 #(
		.INIT('h8)
	) name3873 (
		\P1_reg2_reg[23]/NET0131 ,
		_w2183_,
		_w4336_
	);
	LUT4 #(
		.INIT('hc535)
	) name3874 (
		\P1_reg2_reg[23]/NET0131 ,
		_w1213_,
		_w2189_,
		_w4203_,
		_w4337_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3875 (
		\P1_reg2_reg[23]/NET0131 ,
		_w2121_,
		_w2189_,
		_w4207_,
		_w4338_
	);
	LUT3 #(
		.INIT('h10)
	) name3876 (
		_w489_,
		_w783_,
		_w2194_,
		_w4339_
	);
	LUT4 #(
		.INIT('h007b)
	) name3877 (
		_w784_,
		_w2170_,
		_w2860_,
		_w4339_,
		_w4340_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3878 (
		_w1237_,
		_w4209_,
		_w4210_,
		_w4340_,
		_w4341_
	);
	LUT2 #(
		.INIT('h8)
	) name3879 (
		_w786_,
		_w1120_,
		_w4342_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3880 (
		\P1_reg2_reg[23]/NET0131 ,
		_w2171_,
		_w2196_,
		_w3857_,
		_w4343_
	);
	LUT2 #(
		.INIT('h1)
	) name3881 (
		_w4342_,
		_w4343_,
		_w4344_
	);
	LUT3 #(
		.INIT('hd0)
	) name3882 (
		_w2189_,
		_w4341_,
		_w4344_,
		_w4345_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3883 (
		_w2128_,
		_w4337_,
		_w4338_,
		_w4345_,
		_w4346_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3884 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w4336_,
		_w4346_,
		_w4347_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name3885 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4348_
	);
	LUT2 #(
		.INIT('he)
	) name3886 (
		_w4347_,
		_w4348_,
		_w4349_
	);
	LUT2 #(
		.INIT('h2)
	) name3887 (
		\P2_reg1_reg[16]/NET0131 ,
		_w2042_,
		_w4350_
	);
	LUT4 #(
		.INIT('h2000)
	) name3888 (
		\P2_reg1_reg[16]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4351_
	);
	LUT3 #(
		.INIT('h2a)
	) name3889 (
		\P2_reg1_reg[16]/NET0131 ,
		_w3872_,
		_w3875_,
		_w4352_
	);
	LUT4 #(
		.INIT('h0c04)
	) name3890 (
		_w1802_,
		_w2025_,
		_w3402_,
		_w3717_,
		_w4353_
	);
	LUT4 #(
		.INIT('h2300)
	) name3891 (
		_w1306_,
		_w1800_,
		_w1801_,
		_w2001_,
		_w4354_
	);
	LUT4 #(
		.INIT('h000d)
	) name3892 (
		_w1869_,
		_w3720_,
		_w4354_,
		_w4353_,
		_w4355_
	);
	LUT4 #(
		.INIT('h7020)
	) name3893 (
		_w1305_,
		_w1812_,
		_w2000_,
		_w3711_,
		_w4356_
	);
	LUT4 #(
		.INIT('ha208)
	) name3894 (
		_w1963_,
		_w2404_,
		_w2465_,
		_w2491_,
		_w4357_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3895 (
		_w2762_,
		_w4356_,
		_w4357_,
		_w4355_,
		_w4358_
	);
	LUT4 #(
		.INIT('h1113)
	) name3896 (
		_w1285_,
		_w4351_,
		_w4352_,
		_w4358_,
		_w4359_
	);
	LUT3 #(
		.INIT('hce)
	) name3897 (
		\P1_state_reg[0]/NET0131 ,
		_w4350_,
		_w4359_,
		_w4360_
	);
	LUT3 #(
		.INIT('h2a)
	) name3898 (
		\P2_reg1_reg[20]/NET0131 ,
		_w3225_,
		_w3267_,
		_w4361_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3899 (
		_w3244_,
		_w4189_,
		_w4191_,
		_w4361_,
		_w4362_
	);
	LUT2 #(
		.INIT('h2)
	) name3900 (
		\P2_reg1_reg[21]/NET0131 ,
		_w2042_,
		_w4363_
	);
	LUT4 #(
		.INIT('h2000)
	) name3901 (
		\P2_reg1_reg[21]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4364_
	);
	LUT2 #(
		.INIT('h2)
	) name3902 (
		\P2_reg1_reg[21]/NET0131 ,
		_w2762_,
		_w4365_
	);
	LUT4 #(
		.INIT('h4b00)
	) name3903 (
		_w1842_,
		_w1852_,
		_w2509_,
		_w2762_,
		_w4366_
	);
	LUT3 #(
		.INIT('ha8)
	) name3904 (
		_w1869_,
		_w4365_,
		_w4366_,
		_w4367_
	);
	LUT4 #(
		.INIT('hb400)
	) name3905 (
		_w1918_,
		_w1932_,
		_w2509_,
		_w2762_,
		_w4368_
	);
	LUT3 #(
		.INIT('ha8)
	) name3906 (
		_w1963_,
		_w4365_,
		_w4368_,
		_w4369_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3907 (
		\P2_reg1_reg[21]/NET0131 ,
		_w2762_,
		_w4230_,
		_w4231_,
		_w4370_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3908 (
		\P2_reg1_reg[21]/NET0131 ,
		_w2033_,
		_w2734_,
		_w2762_,
		_w4371_
	);
	LUT4 #(
		.INIT('h0057)
	) name3909 (
		_w2762_,
		_w4275_,
		_w4276_,
		_w4371_,
		_w4372_
	);
	LUT3 #(
		.INIT('hd0)
	) name3910 (
		_w2000_,
		_w4370_,
		_w4372_,
		_w4373_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3911 (
		_w1285_,
		_w4367_,
		_w4369_,
		_w4373_,
		_w4374_
	);
	LUT4 #(
		.INIT('heeec)
	) name3912 (
		\P1_state_reg[0]/NET0131 ,
		_w4363_,
		_w4364_,
		_w4374_,
		_w4375_
	);
	LUT3 #(
		.INIT('h84)
	) name3913 (
		_w2022_,
		_w2025_,
		_w2363_,
		_w4376_
	);
	LUT3 #(
		.INIT('h2a)
	) name3914 (
		\P2_reg1_reg[30]/NET0131 ,
		_w2556_,
		_w3241_,
		_w4377_
	);
	LUT4 #(
		.INIT('hffa2)
	) name3915 (
		_w3244_,
		_w4298_,
		_w4376_,
		_w4377_,
		_w4378_
	);
	LUT2 #(
		.INIT('h2)
	) name3916 (
		\P2_reg2_reg[12]/NET0131 ,
		_w2042_,
		_w4379_
	);
	LUT2 #(
		.INIT('h2)
	) name3917 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1298_,
		_w4380_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3918 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1298_,
		_w2494_,
		_w3003_,
		_w4381_
	);
	LUT4 #(
		.INIT('h2a08)
	) name3919 (
		_w1298_,
		_w1305_,
		_w1740_,
		_w3693_,
		_w4382_
	);
	LUT3 #(
		.INIT('ha8)
	) name3920 (
		_w2000_,
		_w4380_,
		_w4382_,
		_w4383_
	);
	LUT4 #(
		.INIT('h0200)
	) name3921 (
		_w1749_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w4384_
	);
	LUT4 #(
		.INIT('h005d)
	) name3922 (
		\P2_reg2_reg[12]/NET0131 ,
		_w2640_,
		_w3917_,
		_w4384_,
		_w4385_
	);
	LUT3 #(
		.INIT('hd0)
	) name3923 (
		_w1298_,
		_w4328_,
		_w4385_,
		_w4386_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3924 (
		_w1963_,
		_w4381_,
		_w4383_,
		_w4386_,
		_w4387_
	);
	LUT4 #(
		.INIT('h2000)
	) name3925 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4388_
	);
	LUT4 #(
		.INIT('haa08)
	) name3926 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w4387_,
		_w4388_,
		_w4389_
	);
	LUT2 #(
		.INIT('he)
	) name3927 (
		_w4379_,
		_w4389_,
		_w4390_
	);
	LUT2 #(
		.INIT('h2)
	) name3928 (
		\P2_reg2_reg[16]/NET0131 ,
		_w2042_,
		_w4391_
	);
	LUT4 #(
		.INIT('h2000)
	) name3929 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4392_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3930 (
		_w1298_,
		_w4356_,
		_w4357_,
		_w4355_,
		_w4393_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3931 (
		\P2_reg2_reg[16]/NET0131 ,
		_w2031_,
		_w2640_,
		_w3919_,
		_w4394_
	);
	LUT4 #(
		.INIT('h0200)
	) name3932 (
		_w1803_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w4395_
	);
	LUT2 #(
		.INIT('h1)
	) name3933 (
		_w4394_,
		_w4395_,
		_w4396_
	);
	LUT4 #(
		.INIT('h1311)
	) name3934 (
		_w1285_,
		_w4392_,
		_w4393_,
		_w4396_,
		_w4397_
	);
	LUT3 #(
		.INIT('hce)
	) name3935 (
		\P1_state_reg[0]/NET0131 ,
		_w4391_,
		_w4397_,
		_w4398_
	);
	LUT4 #(
		.INIT('h1000)
	) name3936 (
		_w1096_,
		_w1098_,
		_w908_,
		_w1101_,
		_w4399_
	);
	LUT4 #(
		.INIT('hcc08)
	) name3937 (
		_w2189_,
		_w3511_,
		_w4284_,
		_w4399_,
		_w4400_
	);
	LUT4 #(
		.INIT('h00fb)
	) name3938 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w3360_,
		_w4401_
	);
	LUT4 #(
		.INIT('h0010)
	) name3939 (
		_w2171_,
		_w2196_,
		_w3511_,
		_w4401_,
		_w4402_
	);
	LUT2 #(
		.INIT('h2)
	) name3940 (
		\P1_reg2_reg[8]/NET0131 ,
		_w4402_,
		_w4403_
	);
	LUT2 #(
		.INIT('he)
	) name3941 (
		_w4400_,
		_w4403_,
		_w4404_
	);
	LUT2 #(
		.INIT('h2)
	) name3942 (
		\P2_reg2_reg[21]/NET0131 ,
		_w2042_,
		_w4405_
	);
	LUT4 #(
		.INIT('h2000)
	) name3943 (
		\P2_reg2_reg[21]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4406_
	);
	LUT2 #(
		.INIT('h2)
	) name3944 (
		\P2_reg2_reg[21]/NET0131 ,
		_w1298_,
		_w4407_
	);
	LUT4 #(
		.INIT('h208a)
	) name3945 (
		_w1298_,
		_w1842_,
		_w1852_,
		_w2509_,
		_w4408_
	);
	LUT3 #(
		.INIT('ha8)
	) name3946 (
		_w1869_,
		_w4407_,
		_w4408_,
		_w4409_
	);
	LUT4 #(
		.INIT('h8a20)
	) name3947 (
		_w1298_,
		_w1918_,
		_w1932_,
		_w2509_,
		_w4410_
	);
	LUT3 #(
		.INIT('ha8)
	) name3948 (
		_w1963_,
		_w4407_,
		_w4410_,
		_w4411_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3949 (
		\P2_reg2_reg[21]/NET0131 ,
		_w1298_,
		_w4230_,
		_w4231_,
		_w4412_
	);
	LUT2 #(
		.INIT('h8)
	) name3950 (
		_w1570_,
		_w2029_,
		_w4413_
	);
	LUT3 #(
		.INIT('h0d)
	) name3951 (
		\P2_reg2_reg[21]/NET0131 ,
		_w2640_,
		_w4413_,
		_w4414_
	);
	LUT4 #(
		.INIT('h5700)
	) name3952 (
		_w1298_,
		_w4275_,
		_w4276_,
		_w4414_,
		_w4415_
	);
	LUT3 #(
		.INIT('hd0)
	) name3953 (
		_w2000_,
		_w4412_,
		_w4415_,
		_w4416_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3954 (
		_w1285_,
		_w4409_,
		_w4411_,
		_w4416_,
		_w4417_
	);
	LUT4 #(
		.INIT('heeec)
	) name3955 (
		\P1_state_reg[0]/NET0131 ,
		_w4405_,
		_w4406_,
		_w4417_,
		_w4418_
	);
	LUT2 #(
		.INIT('h2)
	) name3956 (
		\P2_reg2_reg[23]/NET0131 ,
		_w2042_,
		_w4419_
	);
	LUT4 #(
		.INIT('h2000)
	) name3957 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4420_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3958 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1298_,
		_w2505_,
		_w4245_,
		_w4421_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3959 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1298_,
		_w1869_,
		_w4250_,
		_w4422_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3960 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1298_,
		_w4252_,
		_w4253_,
		_w4423_
	);
	LUT3 #(
		.INIT('h10)
	) name3961 (
		_w1306_,
		_w1546_,
		_w2001_,
		_w4424_
	);
	LUT4 #(
		.INIT('haa20)
	) name3962 (
		_w1298_,
		_w4255_,
		_w4256_,
		_w4424_,
		_w4425_
	);
	LUT2 #(
		.INIT('h8)
	) name3963 (
		_w1548_,
		_w2029_,
		_w4426_
	);
	LUT3 #(
		.INIT('h0d)
	) name3964 (
		\P2_reg2_reg[23]/NET0131 ,
		_w2640_,
		_w4426_,
		_w4427_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3965 (
		_w2000_,
		_w4423_,
		_w4425_,
		_w4427_,
		_w4428_
	);
	LUT4 #(
		.INIT('h3100)
	) name3966 (
		_w1963_,
		_w4422_,
		_w4421_,
		_w4428_,
		_w4429_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3967 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w4420_,
		_w4429_,
		_w4430_
	);
	LUT2 #(
		.INIT('he)
	) name3968 (
		_w4419_,
		_w4430_,
		_w4431_
	);
	LUT2 #(
		.INIT('h2)
	) name3969 (
		\P2_reg2_reg[30]/NET0131 ,
		_w2042_,
		_w4432_
	);
	LUT4 #(
		.INIT('h2000)
	) name3970 (
		\P2_reg2_reg[30]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4433_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3971 (
		\P2_reg2_reg[30]/NET0131 ,
		_w1863_,
		_w1866_,
		_w2028_,
		_w4434_
	);
	LUT2 #(
		.INIT('h1)
	) name3972 (
		_w1298_,
		_w4434_,
		_w4435_
	);
	LUT3 #(
		.INIT('ha2)
	) name3973 (
		\P2_reg2_reg[30]/NET0131 ,
		_w1298_,
		_w2032_,
		_w4436_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name3974 (
		_w4298_,
		_w4376_,
		_w4435_,
		_w4436_,
		_w4437_
	);
	LUT4 #(
		.INIT('h0507)
	) name3975 (
		_w1285_,
		_w2030_,
		_w4433_,
		_w4437_,
		_w4438_
	);
	LUT3 #(
		.INIT('hce)
	) name3976 (
		\P1_state_reg[0]/NET0131 ,
		_w4432_,
		_w4438_,
		_w4439_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name3977 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[18]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4440_
	);
	LUT2 #(
		.INIT('h8)
	) name3978 (
		\P1_reg0_reg[18]/NET0131 ,
		_w2183_,
		_w4441_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3979 (
		\P1_reg0_reg[18]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4442_
	);
	LUT4 #(
		.INIT('h8848)
	) name3980 (
		_w1216_,
		_w2325_,
		_w2650_,
		_w2657_,
		_w4443_
	);
	LUT3 #(
		.INIT('ha8)
	) name3981 (
		_w2128_,
		_w4442_,
		_w4443_,
		_w4444_
	);
	LUT4 #(
		.INIT('h4484)
	) name3982 (
		_w1216_,
		_w2325_,
		_w2677_,
		_w3375_,
		_w4445_
	);
	LUT3 #(
		.INIT('ha8)
	) name3983 (
		_w2121_,
		_w4442_,
		_w4445_,
		_w4446_
	);
	LUT4 #(
		.INIT('hc808)
	) name3984 (
		\P1_reg0_reg[18]/NET0131 ,
		_w1237_,
		_w2325_,
		_w3379_,
		_w4447_
	);
	LUT4 #(
		.INIT('haaa2)
	) name3985 (
		\P1_reg0_reg[18]/NET0131 ,
		_w2332_,
		_w2333_,
		_w2796_,
		_w4448_
	);
	LUT4 #(
		.INIT('haa20)
	) name3986 (
		_w2325_,
		_w3381_,
		_w3382_,
		_w3831_,
		_w4449_
	);
	LUT2 #(
		.INIT('h1)
	) name3987 (
		_w4448_,
		_w4449_,
		_w4450_
	);
	LUT2 #(
		.INIT('h4)
	) name3988 (
		_w4447_,
		_w4450_,
		_w4451_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3989 (
		_w2182_,
		_w4446_,
		_w4444_,
		_w4451_,
		_w4452_
	);
	LUT4 #(
		.INIT('heeec)
	) name3990 (
		\P1_state_reg[0]/NET0131 ,
		_w4440_,
		_w4441_,
		_w4452_,
		_w4453_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name3991 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[19]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4454_
	);
	LUT2 #(
		.INIT('h8)
	) name3992 (
		\P1_reg0_reg[19]/NET0131 ,
		_w2183_,
		_w4455_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3993 (
		\P1_reg0_reg[19]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4456_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3994 (
		\P1_reg0_reg[19]/NET0131 ,
		_w2325_,
		_w3671_,
		_w3672_,
		_w4457_
	);
	LUT2 #(
		.INIT('h2)
	) name3995 (
		_w1237_,
		_w4457_,
		_w4458_
	);
	LUT4 #(
		.INIT('h4844)
	) name3996 (
		_w1217_,
		_w2325_,
		_w2942_,
		_w2943_,
		_w4459_
	);
	LUT3 #(
		.INIT('ha8)
	) name3997 (
		_w2128_,
		_w4456_,
		_w4459_,
		_w4460_
	);
	LUT4 #(
		.INIT('hc535)
	) name3998 (
		\P1_reg0_reg[19]/NET0131 ,
		_w1217_,
		_w2325_,
		_w3677_,
		_w4461_
	);
	LUT4 #(
		.INIT('haaa2)
	) name3999 (
		\P1_reg0_reg[19]/NET0131 ,
		_w2332_,
		_w2333_,
		_w2796_,
		_w4462_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4000 (
		_w2170_,
		_w3168_,
		_w3680_,
		_w4314_,
		_w4463_
	);
	LUT3 #(
		.INIT('h31)
	) name4001 (
		_w2325_,
		_w4462_,
		_w4463_,
		_w4464_
	);
	LUT3 #(
		.INIT('hd0)
	) name4002 (
		_w2121_,
		_w4461_,
		_w4464_,
		_w4465_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4003 (
		_w2182_,
		_w4460_,
		_w4458_,
		_w4465_,
		_w4466_
	);
	LUT4 #(
		.INIT('heeec)
	) name4004 (
		\P1_state_reg[0]/NET0131 ,
		_w4454_,
		_w4455_,
		_w4466_,
		_w4467_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4005 (
		\P1_reg0_reg[22]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4468_
	);
	LUT4 #(
		.INIT('h007b)
	) name4006 (
		_w1201_,
		_w3563_,
		_w3779_,
		_w4468_,
		_w4469_
	);
	LUT2 #(
		.INIT('h2)
	) name4007 (
		_w2121_,
		_w4469_,
		_w4470_
	);
	LUT4 #(
		.INIT('h00d0)
	) name4008 (
		_w2128_,
		_w3783_,
		_w3789_,
		_w3856_,
		_w4471_
	);
	LUT3 #(
		.INIT('h2a)
	) name4009 (
		\P1_reg0_reg[22]/NET0131 ,
		_w2784_,
		_w3954_,
		_w4472_
	);
	LUT3 #(
		.INIT('h0d)
	) name4010 (
		_w3563_,
		_w4471_,
		_w4472_,
		_w4473_
	);
	LUT2 #(
		.INIT('hb)
	) name4011 (
		_w4470_,
		_w4473_,
		_w4474_
	);
	LUT4 #(
		.INIT('hc535)
	) name4012 (
		\P1_reg0_reg[23]/NET0131 ,
		_w1213_,
		_w2325_,
		_w4203_,
		_w4475_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4013 (
		\P1_reg0_reg[23]/NET0131 ,
		_w2121_,
		_w2325_,
		_w4207_,
		_w4476_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4014 (
		\P1_reg0_reg[23]/NET0131 ,
		_w2332_,
		_w2333_,
		_w2783_,
		_w4477_
	);
	LUT3 #(
		.INIT('h0d)
	) name4015 (
		_w2325_,
		_w4341_,
		_w4477_,
		_w4478_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4016 (
		_w2128_,
		_w4475_,
		_w4476_,
		_w4478_,
		_w4479_
	);
	LUT2 #(
		.INIT('h8)
	) name4017 (
		\P1_reg0_reg[23]/NET0131 ,
		_w2183_,
		_w4480_
	);
	LUT4 #(
		.INIT('haa08)
	) name4018 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w4479_,
		_w4480_,
		_w4481_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4019 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4482_
	);
	LUT2 #(
		.INIT('he)
	) name4020 (
		_w4481_,
		_w4482_,
		_w4483_
	);
	LUT3 #(
		.INIT('h2a)
	) name4021 (
		\P1_reg0_reg[8]/NET0131 ,
		_w2332_,
		_w3563_,
		_w4484_
	);
	LUT3 #(
		.INIT('hf2)
	) name4022 (
		_w3563_,
		_w4284_,
		_w4484_,
		_w4485_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4023 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[9]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4486_
	);
	LUT2 #(
		.INIT('h8)
	) name4024 (
		\P1_reg0_reg[9]/NET0131 ,
		_w2183_,
		_w4487_
	);
	LUT4 #(
		.INIT('hc808)
	) name4025 (
		\P1_reg0_reg[9]/NET0131 ,
		_w1237_,
		_w2325_,
		_w3733_,
		_w4488_
	);
	LUT4 #(
		.INIT('hc808)
	) name4026 (
		\P1_reg0_reg[9]/NET0131 ,
		_w2121_,
		_w2325_,
		_w3735_,
		_w4489_
	);
	LUT2 #(
		.INIT('h2)
	) name4027 (
		\P1_reg0_reg[9]/NET0131 ,
		_w2799_,
		_w4490_
	);
	LUT4 #(
		.INIT('h0075)
	) name4028 (
		_w2325_,
		_w4291_,
		_w4293_,
		_w4490_,
		_w4491_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4029 (
		_w2182_,
		_w4489_,
		_w4488_,
		_w4491_,
		_w4492_
	);
	LUT4 #(
		.INIT('heeec)
	) name4030 (
		\P1_state_reg[0]/NET0131 ,
		_w4486_,
		_w4487_,
		_w4492_,
		_w4493_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4031 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[18]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4494_
	);
	LUT2 #(
		.INIT('h8)
	) name4032 (
		\P1_reg1_reg[18]/NET0131 ,
		_w2183_,
		_w4495_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4033 (
		\P1_reg1_reg[18]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4496_
	);
	LUT4 #(
		.INIT('h8848)
	) name4034 (
		_w1216_,
		_w2536_,
		_w2650_,
		_w2657_,
		_w4497_
	);
	LUT3 #(
		.INIT('ha8)
	) name4035 (
		_w2128_,
		_w4496_,
		_w4497_,
		_w4498_
	);
	LUT4 #(
		.INIT('h4484)
	) name4036 (
		_w1216_,
		_w2536_,
		_w2677_,
		_w3375_,
		_w4499_
	);
	LUT3 #(
		.INIT('ha8)
	) name4037 (
		_w2121_,
		_w4496_,
		_w4499_,
		_w4500_
	);
	LUT4 #(
		.INIT('hc808)
	) name4038 (
		\P1_reg1_reg[18]/NET0131 ,
		_w1237_,
		_w2536_,
		_w3379_,
		_w4501_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4039 (
		\P1_reg1_reg[18]/NET0131 ,
		_w2332_,
		_w2544_,
		_w2817_,
		_w4502_
	);
	LUT4 #(
		.INIT('haa20)
	) name4040 (
		_w2536_,
		_w3381_,
		_w3382_,
		_w3831_,
		_w4503_
	);
	LUT2 #(
		.INIT('h1)
	) name4041 (
		_w4502_,
		_w4503_,
		_w4504_
	);
	LUT2 #(
		.INIT('h4)
	) name4042 (
		_w4501_,
		_w4504_,
		_w4505_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4043 (
		_w2182_,
		_w4500_,
		_w4498_,
		_w4505_,
		_w4506_
	);
	LUT4 #(
		.INIT('heeec)
	) name4044 (
		\P1_state_reg[0]/NET0131 ,
		_w4494_,
		_w4495_,
		_w4506_,
		_w4507_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4045 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[19]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4508_
	);
	LUT2 #(
		.INIT('h8)
	) name4046 (
		\P1_reg1_reg[19]/NET0131 ,
		_w2183_,
		_w4509_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4047 (
		\P1_reg1_reg[19]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4510_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4048 (
		\P1_reg1_reg[19]/NET0131 ,
		_w2536_,
		_w3671_,
		_w3672_,
		_w4511_
	);
	LUT2 #(
		.INIT('h2)
	) name4049 (
		_w1237_,
		_w4511_,
		_w4512_
	);
	LUT4 #(
		.INIT('h4844)
	) name4050 (
		_w1217_,
		_w2536_,
		_w2942_,
		_w2943_,
		_w4513_
	);
	LUT3 #(
		.INIT('ha8)
	) name4051 (
		_w2128_,
		_w4510_,
		_w4513_,
		_w4514_
	);
	LUT4 #(
		.INIT('hc535)
	) name4052 (
		\P1_reg1_reg[19]/NET0131 ,
		_w1217_,
		_w2536_,
		_w3677_,
		_w4515_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4053 (
		\P1_reg1_reg[19]/NET0131 ,
		_w2332_,
		_w2544_,
		_w2817_,
		_w4516_
	);
	LUT3 #(
		.INIT('h0d)
	) name4054 (
		_w2536_,
		_w4463_,
		_w4516_,
		_w4517_
	);
	LUT3 #(
		.INIT('hd0)
	) name4055 (
		_w2121_,
		_w4515_,
		_w4517_,
		_w4518_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4056 (
		_w2182_,
		_w4514_,
		_w4512_,
		_w4518_,
		_w4519_
	);
	LUT4 #(
		.INIT('heeec)
	) name4057 (
		\P1_state_reg[0]/NET0131 ,
		_w4508_,
		_w4509_,
		_w4519_,
		_w4520_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4058 (
		\P1_reg1_reg[22]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4521_
	);
	LUT4 #(
		.INIT('h007b)
	) name4059 (
		_w1201_,
		_w3608_,
		_w3779_,
		_w4521_,
		_w4522_
	);
	LUT2 #(
		.INIT('h2)
	) name4060 (
		_w2121_,
		_w4522_,
		_w4523_
	);
	LUT4 #(
		.INIT('h0200)
	) name4061 (
		_w2332_,
		_w2544_,
		_w2817_,
		_w3511_,
		_w4524_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4062 (
		\P1_reg1_reg[22]/NET0131 ,
		_w2816_,
		_w3605_,
		_w4524_,
		_w4525_
	);
	LUT3 #(
		.INIT('h0d)
	) name4063 (
		_w3608_,
		_w4471_,
		_w4525_,
		_w4526_
	);
	LUT2 #(
		.INIT('hb)
	) name4064 (
		_w4523_,
		_w4526_,
		_w4527_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4065 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4528_
	);
	LUT4 #(
		.INIT('hc535)
	) name4066 (
		\P1_reg1_reg[23]/NET0131 ,
		_w1213_,
		_w2536_,
		_w4203_,
		_w4529_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4067 (
		\P1_reg1_reg[23]/NET0131 ,
		_w2121_,
		_w2536_,
		_w4207_,
		_w4530_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4068 (
		\P1_reg1_reg[23]/NET0131 ,
		_w2332_,
		_w2816_,
		_w3975_,
		_w4531_
	);
	LUT3 #(
		.INIT('h0d)
	) name4069 (
		_w2536_,
		_w4341_,
		_w4531_,
		_w4532_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4070 (
		_w2128_,
		_w4529_,
		_w4530_,
		_w4532_,
		_w4533_
	);
	LUT2 #(
		.INIT('h8)
	) name4071 (
		\P1_reg1_reg[23]/NET0131 ,
		_w2183_,
		_w4534_
	);
	LUT4 #(
		.INIT('haa08)
	) name4072 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w4533_,
		_w4534_,
		_w4535_
	);
	LUT2 #(
		.INIT('he)
	) name4073 (
		_w4528_,
		_w4535_,
		_w4536_
	);
	LUT2 #(
		.INIT('h2)
	) name4074 (
		\P2_reg0_reg[12]/NET0131 ,
		_w2042_,
		_w4537_
	);
	LUT2 #(
		.INIT('h2)
	) name4075 (
		\P2_reg0_reg[12]/NET0131 ,
		_w2729_,
		_w4538_
	);
	LUT4 #(
		.INIT('hc535)
	) name4076 (
		\P2_reg0_reg[12]/NET0131 ,
		_w2494_,
		_w2729_,
		_w3003_,
		_w4539_
	);
	LUT4 #(
		.INIT('h7020)
	) name4077 (
		_w1305_,
		_w1740_,
		_w2729_,
		_w3693_,
		_w4540_
	);
	LUT3 #(
		.INIT('ha8)
	) name4078 (
		_w2000_,
		_w4538_,
		_w4540_,
		_w4541_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4079 (
		\P2_reg0_reg[12]/NET0131 ,
		_w2494_,
		_w2729_,
		_w3025_,
		_w4542_
	);
	LUT4 #(
		.INIT('h3c55)
	) name4080 (
		\P2_reg0_reg[12]/NET0131 ,
		_w1759_,
		_w2009_,
		_w2729_,
		_w4543_
	);
	LUT2 #(
		.INIT('h2)
	) name4081 (
		\P2_reg0_reg[12]/NET0131 ,
		_w2734_,
		_w4544_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4082 (
		\P2_reg0_reg[12]/NET0131 ,
		_w1759_,
		_w2001_,
		_w2729_,
		_w4545_
	);
	LUT2 #(
		.INIT('h1)
	) name4083 (
		_w4544_,
		_w4545_,
		_w4546_
	);
	LUT3 #(
		.INIT('hd0)
	) name4084 (
		_w2025_,
		_w4543_,
		_w4546_,
		_w4547_
	);
	LUT3 #(
		.INIT('hd0)
	) name4085 (
		_w1869_,
		_w4542_,
		_w4547_,
		_w4548_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4086 (
		_w1963_,
		_w4539_,
		_w4541_,
		_w4548_,
		_w4549_
	);
	LUT4 #(
		.INIT('h2000)
	) name4087 (
		\P2_reg0_reg[12]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4550_
	);
	LUT4 #(
		.INIT('haa08)
	) name4088 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w4549_,
		_w4550_,
		_w4551_
	);
	LUT2 #(
		.INIT('he)
	) name4089 (
		_w4537_,
		_w4551_,
		_w4552_
	);
	LUT2 #(
		.INIT('h2)
	) name4090 (
		\P2_reg0_reg[16]/NET0131 ,
		_w2042_,
		_w4553_
	);
	LUT4 #(
		.INIT('h2000)
	) name4091 (
		\P2_reg0_reg[16]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4554_
	);
	LUT2 #(
		.INIT('h2)
	) name4092 (
		\P2_reg0_reg[16]/NET0131 ,
		_w2729_,
		_w4555_
	);
	LUT4 #(
		.INIT('h7020)
	) name4093 (
		_w1305_,
		_w1812_,
		_w2729_,
		_w3711_,
		_w4556_
	);
	LUT3 #(
		.INIT('ha8)
	) name4094 (
		_w2000_,
		_w4555_,
		_w4556_,
		_w4557_
	);
	LUT4 #(
		.INIT('hd200)
	) name4095 (
		_w2404_,
		_w2465_,
		_w2491_,
		_w2729_,
		_w4558_
	);
	LUT3 #(
		.INIT('ha8)
	) name4096 (
		_w1963_,
		_w4555_,
		_w4558_,
		_w4559_
	);
	LUT2 #(
		.INIT('h2)
	) name4097 (
		_w1869_,
		_w2729_,
		_w4560_
	);
	LUT3 #(
		.INIT('ha2)
	) name4098 (
		\P2_reg0_reg[16]/NET0131 ,
		_w3084_,
		_w4560_,
		_w4561_
	);
	LUT3 #(
		.INIT('h0d)
	) name4099 (
		_w2729_,
		_w4355_,
		_w4561_,
		_w4562_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4100 (
		_w1285_,
		_w4559_,
		_w4557_,
		_w4562_,
		_w4563_
	);
	LUT4 #(
		.INIT('heeec)
	) name4101 (
		\P1_state_reg[0]/NET0131 ,
		_w4553_,
		_w4554_,
		_w4563_,
		_w4564_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4102 (
		\P2_reg0_reg[20]/NET0131 ,
		_w3082_,
		_w3083_,
		_w4302_,
		_w4565_
	);
	LUT4 #(
		.INIT('hff8a)
	) name4103 (
		_w3153_,
		_w4189_,
		_w4191_,
		_w4565_,
		_w4566_
	);
	LUT2 #(
		.INIT('h8)
	) name4104 (
		_w844_,
		_w2183_,
		_w4567_
	);
	LUT4 #(
		.INIT('h4144)
	) name4105 (
		_w488_,
		_w837_,
		_w847_,
		_w3351_,
		_w4568_
	);
	LUT3 #(
		.INIT('h80)
	) name4106 (
		_w488_,
		_w854_,
		_w855_,
		_w4569_
	);
	LUT4 #(
		.INIT('h1110)
	) name4107 (
		_w844_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4570_
	);
	LUT2 #(
		.INIT('h2)
	) name4108 (
		_w1237_,
		_w4570_,
		_w4571_
	);
	LUT4 #(
		.INIT('h5700)
	) name4109 (
		_w2055_,
		_w4568_,
		_w4569_,
		_w4571_,
		_w4572_
	);
	LUT3 #(
		.INIT('h84)
	) name4110 (
		_w1166_,
		_w2128_,
		_w2243_,
		_w4573_
	);
	LUT4 #(
		.INIT('h1555)
	) name4111 (
		_w852_,
		_w2159_,
		_w2160_,
		_w2858_,
		_w4574_
	);
	LUT3 #(
		.INIT('h02)
	) name4112 (
		_w2170_,
		_w2859_,
		_w4574_,
		_w4575_
	);
	LUT4 #(
		.INIT('h8488)
	) name4113 (
		_w1166_,
		_w2121_,
		_w2276_,
		_w2283_,
		_w4576_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4114 (
		_w2055_,
		_w4575_,
		_w4576_,
		_w4573_,
		_w4577_
	);
	LUT3 #(
		.INIT('h10)
	) name4115 (
		_w852_,
		_w2175_,
		_w2176_,
		_w4578_
	);
	LUT3 #(
		.INIT('h0d)
	) name4116 (
		_w844_,
		_w4057_,
		_w4578_,
		_w4579_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4117 (
		_w2182_,
		_w4577_,
		_w4572_,
		_w4579_,
		_w4580_
	);
	LUT2 #(
		.INIT('h2)
	) name4118 (
		\P1_reg3_reg[13]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4581_
	);
	LUT3 #(
		.INIT('h07)
	) name4119 (
		_w844_,
		_w1244_,
		_w4581_,
		_w4582_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4120 (
		\P1_state_reg[0]/NET0131 ,
		_w4567_,
		_w4580_,
		_w4582_,
		_w4583_
	);
	LUT4 #(
		.INIT('h4000)
	) name4121 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1737_,
		_w4584_
	);
	LUT2 #(
		.INIT('h2)
	) name4122 (
		_w1737_,
		_w2903_,
		_w4585_
	);
	LUT4 #(
		.INIT('h5054)
	) name4123 (
		_w1305_,
		_w1752_,
		_w1976_,
		_w4087_,
		_w4586_
	);
	LUT3 #(
		.INIT('h80)
	) name4124 (
		_w1305_,
		_w1761_,
		_w1763_,
		_w4587_
	);
	LUT4 #(
		.INIT('h3331)
	) name4125 (
		_w2903_,
		_w4585_,
		_w4586_,
		_w4587_,
		_w4588_
	);
	LUT4 #(
		.INIT('h6500)
	) name4126 (
		_w2495_,
		_w2614_,
		_w2615_,
		_w2903_,
		_w4589_
	);
	LUT3 #(
		.INIT('ha8)
	) name4127 (
		_w1869_,
		_w4585_,
		_w4589_,
		_w4590_
	);
	LUT4 #(
		.INIT('h009f)
	) name4128 (
		_w2495_,
		_w2593_,
		_w2903_,
		_w4585_,
		_w4591_
	);
	LUT3 #(
		.INIT('h8a)
	) name4129 (
		_w1747_,
		_w1774_,
		_w4094_,
		_w4592_
	);
	LUT2 #(
		.INIT('h4)
	) name4130 (
		_w2009_,
		_w2025_,
		_w4593_
	);
	LUT4 #(
		.INIT('h88a8)
	) name4131 (
		_w1737_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w4594_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name4132 (
		_w1747_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w4595_
	);
	LUT2 #(
		.INIT('h1)
	) name4133 (
		_w4594_,
		_w4595_,
		_w4596_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4134 (
		_w2903_,
		_w4592_,
		_w4593_,
		_w4596_,
		_w4597_
	);
	LUT3 #(
		.INIT('hd0)
	) name4135 (
		_w1963_,
		_w4591_,
		_w4597_,
		_w4598_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4136 (
		_w2000_,
		_w4588_,
		_w4590_,
		_w4598_,
		_w4599_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4137 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w4584_,
		_w4599_,
		_w4600_
	);
	LUT2 #(
		.INIT('h4)
	) name4138 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		_w4601_
	);
	LUT3 #(
		.INIT('h07)
	) name4139 (
		_w1737_,
		_w2344_,
		_w4601_,
		_w4602_
	);
	LUT2 #(
		.INIT('hb)
	) name4140 (
		_w4600_,
		_w4602_,
		_w4603_
	);
	LUT4 #(
		.INIT('h4000)
	) name4141 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1823_,
		_w4604_
	);
	LUT2 #(
		.INIT('h2)
	) name4142 (
		_w1823_,
		_w2903_,
		_w4605_
	);
	LUT2 #(
		.INIT('h9)
	) name4143 (
		_w1825_,
		_w1830_,
		_w4606_
	);
	LUT4 #(
		.INIT('ha208)
	) name4144 (
		_w2903_,
		_w3115_,
		_w3491_,
		_w4606_,
		_w4607_
	);
	LUT3 #(
		.INIT('ha8)
	) name4145 (
		_w1963_,
		_w4605_,
		_w4607_,
		_w4608_
	);
	LUT3 #(
		.INIT('h80)
	) name4146 (
		_w1305_,
		_w1832_,
		_w1833_,
		_w4609_
	);
	LUT4 #(
		.INIT('h00eb)
	) name4147 (
		_w1305_,
		_w1812_,
		_w1978_,
		_w4609_,
		_w4610_
	);
	LUT4 #(
		.INIT('hc808)
	) name4148 (
		_w1823_,
		_w2000_,
		_w2903_,
		_w4610_,
		_w4611_
	);
	LUT4 #(
		.INIT('h4fb0)
	) name4149 (
		_w3095_,
		_w3096_,
		_w3097_,
		_w4606_,
		_w4612_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4150 (
		_w1823_,
		_w1869_,
		_w2903_,
		_w4612_,
		_w4613_
	);
	LUT4 #(
		.INIT('h9500)
	) name4151 (
		_w1830_,
		_w2009_,
		_w2010_,
		_w2025_,
		_w4614_
	);
	LUT4 #(
		.INIT('h88a8)
	) name4152 (
		_w1823_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w4615_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name4153 (
		_w1830_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w4616_
	);
	LUT2 #(
		.INIT('h1)
	) name4154 (
		_w4615_,
		_w4616_,
		_w4617_
	);
	LUT3 #(
		.INIT('h70)
	) name4155 (
		_w2903_,
		_w4614_,
		_w4617_,
		_w4618_
	);
	LUT3 #(
		.INIT('h10)
	) name4156 (
		_w4613_,
		_w4611_,
		_w4618_,
		_w4619_
	);
	LUT4 #(
		.INIT('h1311)
	) name4157 (
		_w1285_,
		_w4604_,
		_w4608_,
		_w4619_,
		_w4620_
	);
	LUT2 #(
		.INIT('h4)
	) name4158 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[14]/NET0131 ,
		_w4621_
	);
	LUT3 #(
		.INIT('h07)
	) name4159 (
		_w1823_,
		_w2344_,
		_w4621_,
		_w4622_
	);
	LUT3 #(
		.INIT('h2f)
	) name4160 (
		\P1_state_reg[0]/NET0131 ,
		_w4620_,
		_w4622_,
		_w4623_
	);
	LUT2 #(
		.INIT('h8)
	) name4161 (
		_w958_,
		_w2183_,
		_w4624_
	);
	LUT4 #(
		.INIT('h5655)
	) name4162 (
		_w949_,
		_w961_,
		_w971_,
		_w2130_,
		_w4625_
	);
	LUT4 #(
		.INIT('h80d0)
	) name4163 (
		_w488_,
		_w971_,
		_w2055_,
		_w4625_,
		_w4626_
	);
	LUT3 #(
		.INIT('h01)
	) name4164 (
		_w2171_,
		_w2173_,
		_w4056_,
		_w4627_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4165 (
		_w958_,
		_w1237_,
		_w4626_,
		_w4627_,
		_w4628_
	);
	LUT4 #(
		.INIT('h7020)
	) name4166 (
		_w488_,
		_w971_,
		_w1237_,
		_w4625_,
		_w4629_
	);
	LUT4 #(
		.INIT('hd000)
	) name4167 (
		_w986_,
		_w1003_,
		_w1006_,
		_w1177_,
		_w4630_
	);
	LUT4 #(
		.INIT('h002f)
	) name4168 (
		_w986_,
		_w1003_,
		_w1006_,
		_w1177_,
		_w4631_
	);
	LUT3 #(
		.INIT('h02)
	) name4169 (
		_w2128_,
		_w4631_,
		_w4630_,
		_w4632_
	);
	LUT2 #(
		.INIT('h4)
	) name4170 (
		_w966_,
		_w2194_,
		_w4633_
	);
	LUT4 #(
		.INIT('h009f)
	) name4171 (
		_w966_,
		_w2156_,
		_w2170_,
		_w4633_,
		_w4634_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4172 (
		_w1177_,
		_w2074_,
		_w2121_,
		_w4634_,
		_w4635_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4173 (
		_w2055_,
		_w4629_,
		_w4632_,
		_w4635_,
		_w4636_
	);
	LUT2 #(
		.INIT('h4)
	) name4174 (
		_w966_,
		_w1120_,
		_w4637_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4175 (
		_w2182_,
		_w4636_,
		_w4628_,
		_w4637_,
		_w4638_
	);
	LUT3 #(
		.INIT('h6c)
	) name4176 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4639_
	);
	LUT4 #(
		.INIT('h7b00)
	) name4177 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4639_,
		_w4640_
	);
	LUT4 #(
		.INIT('hffa8)
	) name4178 (
		\P1_state_reg[0]/NET0131 ,
		_w4624_,
		_w4638_,
		_w4640_,
		_w4641_
	);
	LUT4 #(
		.INIT('h4000)
	) name4179 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1689_,
		_w4642_
	);
	LUT2 #(
		.INIT('h2)
	) name4180 (
		_w1689_,
		_w2903_,
		_w4643_
	);
	LUT3 #(
		.INIT('h2a)
	) name4181 (
		_w1305_,
		_w1697_,
		_w1699_,
		_w4644_
	);
	LUT4 #(
		.INIT('h1405)
	) name4182 (
		_w1305_,
		_w1691_,
		_w1779_,
		_w1972_,
		_w4645_
	);
	LUT4 #(
		.INIT('h1113)
	) name4183 (
		_w2903_,
		_w4643_,
		_w4644_,
		_w4645_,
		_w4646_
	);
	LUT2 #(
		.INIT('h2)
	) name4184 (
		_w2000_,
		_w4646_,
		_w4647_
	);
	LUT4 #(
		.INIT('h009f)
	) name4185 (
		_w2413_,
		_w2499_,
		_w2903_,
		_w4643_,
		_w4648_
	);
	LUT4 #(
		.INIT('h4844)
	) name4186 (
		_w2499_,
		_w2903_,
		_w3014_,
		_w3017_,
		_w4649_
	);
	LUT4 #(
		.INIT('h6500)
	) name4187 (
		_w1695_,
		_w1706_,
		_w2005_,
		_w2025_,
		_w4650_
	);
	LUT4 #(
		.INIT('h88a8)
	) name4188 (
		_w1689_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w4651_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name4189 (
		_w1695_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w4652_
	);
	LUT2 #(
		.INIT('h1)
	) name4190 (
		_w4651_,
		_w4652_,
		_w4653_
	);
	LUT3 #(
		.INIT('h70)
	) name4191 (
		_w2903_,
		_w4650_,
		_w4653_,
		_w4654_
	);
	LUT4 #(
		.INIT('h5700)
	) name4192 (
		_w1869_,
		_w4643_,
		_w4649_,
		_w4654_,
		_w4655_
	);
	LUT3 #(
		.INIT('hd0)
	) name4193 (
		_w1963_,
		_w4648_,
		_w4655_,
		_w4656_
	);
	LUT4 #(
		.INIT('h1311)
	) name4194 (
		_w1285_,
		_w4642_,
		_w4647_,
		_w4656_,
		_w4657_
	);
	LUT2 #(
		.INIT('h4)
	) name4195 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		_w4658_
	);
	LUT3 #(
		.INIT('h07)
	) name4196 (
		_w1689_,
		_w2344_,
		_w4658_,
		_w4659_
	);
	LUT3 #(
		.INIT('h2f)
	) name4197 (
		\P1_state_reg[0]/NET0131 ,
		_w4657_,
		_w4659_,
		_w4660_
	);
	LUT2 #(
		.INIT('h8)
	) name4198 (
		_w947_,
		_w2183_,
		_w4661_
	);
	LUT3 #(
		.INIT('h80)
	) name4199 (
		_w488_,
		_w959_,
		_w960_,
		_w4662_
	);
	LUT4 #(
		.INIT('h00eb)
	) name4200 (
		_w488_,
		_w927_,
		_w4169_,
		_w4662_,
		_w4663_
	);
	LUT4 #(
		.INIT('h50d0)
	) name4201 (
		_w1237_,
		_w2055_,
		_w4627_,
		_w4663_,
		_w4664_
	);
	LUT2 #(
		.INIT('h2)
	) name4202 (
		_w947_,
		_w4664_,
		_w4665_
	);
	LUT3 #(
		.INIT('h84)
	) name4203 (
		_w1192_,
		_w2121_,
		_w2272_,
		_w4666_
	);
	LUT2 #(
		.INIT('h4)
	) name4204 (
		_w956_,
		_w2194_,
		_w4667_
	);
	LUT4 #(
		.INIT('h6a00)
	) name4205 (
		_w956_,
		_w966_,
		_w2156_,
		_w2170_,
		_w4668_
	);
	LUT2 #(
		.INIT('h1)
	) name4206 (
		_w4667_,
		_w4668_,
		_w4669_
	);
	LUT4 #(
		.INIT('h7b00)
	) name4207 (
		_w1192_,
		_w2128_,
		_w2232_,
		_w4669_,
		_w4670_
	);
	LUT4 #(
		.INIT('h0700)
	) name4208 (
		_w1237_,
		_w4663_,
		_w4666_,
		_w4670_,
		_w4671_
	);
	LUT2 #(
		.INIT('h4)
	) name4209 (
		_w956_,
		_w1120_,
		_w4672_
	);
	LUT3 #(
		.INIT('h0d)
	) name4210 (
		_w2055_,
		_w4671_,
		_w4672_,
		_w4673_
	);
	LUT4 #(
		.INIT('h1311)
	) name4211 (
		_w2182_,
		_w4661_,
		_w4665_,
		_w4673_,
		_w4674_
	);
	LUT2 #(
		.INIT('h2)
	) name4212 (
		\P1_reg3_reg[5]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4675_
	);
	LUT4 #(
		.INIT('h4080)
	) name4213 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w947_,
		_w1242_,
		_w4676_
	);
	LUT2 #(
		.INIT('h1)
	) name4214 (
		_w4675_,
		_w4676_,
		_w4677_
	);
	LUT3 #(
		.INIT('h2f)
	) name4215 (
		\P1_state_reg[0]/NET0131 ,
		_w4674_,
		_w4677_,
		_w4678_
	);
	LUT2 #(
		.INIT('h2)
	) name4216 (
		\P2_reg0_reg[23]/NET0131 ,
		_w2042_,
		_w4679_
	);
	LUT4 #(
		.INIT('h2000)
	) name4217 (
		\P2_reg0_reg[23]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4680_
	);
	LUT4 #(
		.INIT('hc535)
	) name4218 (
		\P2_reg0_reg[23]/NET0131 ,
		_w2505_,
		_w2729_,
		_w4245_,
		_w4681_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4219 (
		\P2_reg0_reg[23]/NET0131 ,
		_w1869_,
		_w2729_,
		_w4250_,
		_w4682_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4220 (
		\P2_reg0_reg[23]/NET0131 ,
		_w2729_,
		_w4252_,
		_w4253_,
		_w4683_
	);
	LUT2 #(
		.INIT('h2)
	) name4221 (
		\P2_reg0_reg[23]/NET0131 ,
		_w3084_,
		_w4684_
	);
	LUT4 #(
		.INIT('haa20)
	) name4222 (
		_w2729_,
		_w4255_,
		_w4256_,
		_w4424_,
		_w4685_
	);
	LUT4 #(
		.INIT('h0031)
	) name4223 (
		_w2000_,
		_w4684_,
		_w4683_,
		_w4685_,
		_w4686_
	);
	LUT4 #(
		.INIT('h3100)
	) name4224 (
		_w1963_,
		_w4682_,
		_w4681_,
		_w4686_,
		_w4687_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4225 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w4680_,
		_w4687_,
		_w4688_
	);
	LUT2 #(
		.INIT('he)
	) name4226 (
		_w4679_,
		_w4688_,
		_w4689_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4227 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4690_
	);
	LUT2 #(
		.INIT('h8)
	) name4228 (
		\P1_reg2_reg[10]/NET0131 ,
		_w2183_,
		_w4691_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4229 (
		\P1_reg2_reg[10]/NET0131 ,
		_w2189_,
		_w4025_,
		_w4026_,
		_w4692_
	);
	LUT2 #(
		.INIT('h2)
	) name4230 (
		_w1237_,
		_w4692_,
		_w4693_
	);
	LUT4 #(
		.INIT('hc535)
	) name4231 (
		\P1_reg2_reg[10]/NET0131 ,
		_w1178_,
		_w2189_,
		_w2682_,
		_w4694_
	);
	LUT2 #(
		.INIT('h2)
	) name4232 (
		_w2121_,
		_w4694_,
		_w4695_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4233 (
		\P1_reg2_reg[10]/NET0131 ,
		_w1178_,
		_w2189_,
		_w2653_,
		_w4696_
	);
	LUT4 #(
		.INIT('h1000)
	) name4234 (
		_w1096_,
		_w1098_,
		_w886_,
		_w1101_,
		_w4697_
	);
	LUT4 #(
		.INIT('h0057)
	) name4235 (
		\P1_reg2_reg[10]/NET0131 ,
		_w2171_,
		_w3173_,
		_w4697_,
		_w4698_
	);
	LUT4 #(
		.INIT('h5700)
	) name4236 (
		_w2189_,
		_w4032_,
		_w4034_,
		_w4698_,
		_w4699_
	);
	LUT3 #(
		.INIT('hd0)
	) name4237 (
		_w2128_,
		_w4696_,
		_w4699_,
		_w4700_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4238 (
		_w2182_,
		_w4693_,
		_w4695_,
		_w4700_,
		_w4701_
	);
	LUT4 #(
		.INIT('heeec)
	) name4239 (
		\P1_state_reg[0]/NET0131 ,
		_w4690_,
		_w4691_,
		_w4701_,
		_w4702_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4240 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[11]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4703_
	);
	LUT2 #(
		.INIT('h8)
	) name4241 (
		\P1_reg2_reg[11]/NET0131 ,
		_w2183_,
		_w4704_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4242 (
		\P1_reg2_reg[11]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4705_
	);
	LUT4 #(
		.INIT('h7020)
	) name4243 (
		_w488_,
		_w889_,
		_w2189_,
		_w4004_,
		_w4706_
	);
	LUT3 #(
		.INIT('ha8)
	) name4244 (
		_w1237_,
		_w4705_,
		_w4706_,
		_w4707_
	);
	LUT4 #(
		.INIT('h8488)
	) name4245 (
		_w1174_,
		_w2189_,
		_w2962_,
		_w2963_,
		_w4708_
	);
	LUT3 #(
		.INIT('ha8)
	) name4246 (
		_w2121_,
		_w4705_,
		_w4708_,
		_w4709_
	);
	LUT4 #(
		.INIT('h1555)
	) name4247 (
		_w1100_,
		_w893_,
		_w2159_,
		_w2160_,
		_w4710_
	);
	LUT4 #(
		.INIT('h5f1b)
	) name4248 (
		_w884_,
		_w2172_,
		_w4033_,
		_w4710_,
		_w4711_
	);
	LUT4 #(
		.INIT('h7b00)
	) name4249 (
		_w1174_,
		_w2128_,
		_w2938_,
		_w4711_,
		_w4712_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4250 (
		\P1_reg2_reg[11]/NET0131 ,
		_w2171_,
		_w3173_,
		_w3174_,
		_w4713_
	);
	LUT4 #(
		.INIT('h1000)
	) name4251 (
		_w1096_,
		_w1098_,
		_w874_,
		_w1101_,
		_w4714_
	);
	LUT2 #(
		.INIT('h1)
	) name4252 (
		_w4713_,
		_w4714_,
		_w4715_
	);
	LUT3 #(
		.INIT('hd0)
	) name4253 (
		_w2189_,
		_w4712_,
		_w4715_,
		_w4716_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4254 (
		_w2182_,
		_w4709_,
		_w4707_,
		_w4716_,
		_w4717_
	);
	LUT4 #(
		.INIT('heeec)
	) name4255 (
		\P1_state_reg[0]/NET0131 ,
		_w4703_,
		_w4704_,
		_w4717_,
		_w4718_
	);
	LUT2 #(
		.INIT('h2)
	) name4256 (
		\P1_reg2_reg[13]/NET0131 ,
		_w4402_,
		_w4719_
	);
	LUT4 #(
		.INIT('h1000)
	) name4257 (
		_w1096_,
		_w1098_,
		_w844_,
		_w1101_,
		_w4720_
	);
	LUT3 #(
		.INIT('h02)
	) name4258 (
		_w1237_,
		_w4568_,
		_w4569_,
		_w4721_
	);
	LUT4 #(
		.INIT('hf100)
	) name4259 (
		_w489_,
		_w849_,
		_w851_,
		_w2194_,
		_w4722_
	);
	LUT4 #(
		.INIT('h0001)
	) name4260 (
		_w4575_,
		_w4576_,
		_w4573_,
		_w4722_,
		_w4723_
	);
	LUT4 #(
		.INIT('h1311)
	) name4261 (
		_w2189_,
		_w4720_,
		_w4721_,
		_w4723_,
		_w4724_
	);
	LUT3 #(
		.INIT('hce)
	) name4262 (
		_w3511_,
		_w4719_,
		_w4724_,
		_w4725_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4263 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[14]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4726_
	);
	LUT2 #(
		.INIT('h8)
	) name4264 (
		\P1_reg2_reg[14]/NET0131 ,
		_w2183_,
		_w4727_
	);
	LUT4 #(
		.INIT('hf100)
	) name4265 (
		_w489_,
		_w839_,
		_w841_,
		_w2194_,
		_w4728_
	);
	LUT4 #(
		.INIT('h7020)
	) name4266 (
		_w488_,
		_w847_,
		_w1237_,
		_w4045_,
		_w4729_
	);
	LUT4 #(
		.INIT('h0004)
	) name4267 (
		_w4052_,
		_w4054_,
		_w4728_,
		_w4729_,
		_w4730_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4268 (
		\P1_reg2_reg[14]/NET0131 ,
		_w2171_,
		_w2196_,
		_w4401_,
		_w4731_
	);
	LUT4 #(
		.INIT('h1000)
	) name4269 (
		_w1096_,
		_w1098_,
		_w835_,
		_w1101_,
		_w4732_
	);
	LUT2 #(
		.INIT('h1)
	) name4270 (
		_w4731_,
		_w4732_,
		_w4733_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4271 (
		_w2182_,
		_w2189_,
		_w4730_,
		_w4733_,
		_w4734_
	);
	LUT4 #(
		.INIT('heeec)
	) name4272 (
		\P1_state_reg[0]/NET0131 ,
		_w4726_,
		_w4727_,
		_w4734_,
		_w4735_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4273 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[15]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4736_
	);
	LUT2 #(
		.INIT('h8)
	) name4274 (
		\P1_reg2_reg[15]/NET0131 ,
		_w2183_,
		_w4737_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4275 (
		\P1_reg2_reg[15]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4738_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4276 (
		\P1_reg2_reg[15]/NET0131 ,
		_w1168_,
		_w2189_,
		_w4066_,
		_w4739_
	);
	LUT2 #(
		.INIT('h2)
	) name4277 (
		_w2121_,
		_w4739_,
		_w4740_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4278 (
		\P1_reg2_reg[15]/NET0131 ,
		_w2128_,
		_w2189_,
		_w4069_,
		_w4741_
	);
	LUT4 #(
		.INIT('h7020)
	) name4279 (
		_w488_,
		_w837_,
		_w2189_,
		_w4071_,
		_w4742_
	);
	LUT3 #(
		.INIT('ha8)
	) name4280 (
		_w1237_,
		_w4738_,
		_w4742_,
		_w4743_
	);
	LUT4 #(
		.INIT('hc808)
	) name4281 (
		\P1_reg2_reg[15]/NET0131 ,
		_w2170_,
		_w2189_,
		_w4074_,
		_w4744_
	);
	LUT4 #(
		.INIT('hf100)
	) name4282 (
		_w489_,
		_w829_,
		_w832_,
		_w2194_,
		_w4745_
	);
	LUT2 #(
		.INIT('h8)
	) name4283 (
		_w2189_,
		_w4745_,
		_w4746_
	);
	LUT4 #(
		.INIT('h1000)
	) name4284 (
		_w1096_,
		_w1098_,
		_w825_,
		_w1101_,
		_w4747_
	);
	LUT4 #(
		.INIT('h0057)
	) name4285 (
		\P1_reg2_reg[15]/NET0131 ,
		_w2171_,
		_w2196_,
		_w4747_,
		_w4748_
	);
	LUT2 #(
		.INIT('h4)
	) name4286 (
		_w4746_,
		_w4748_,
		_w4749_
	);
	LUT2 #(
		.INIT('h4)
	) name4287 (
		_w4744_,
		_w4749_,
		_w4750_
	);
	LUT3 #(
		.INIT('h10)
	) name4288 (
		_w4743_,
		_w4741_,
		_w4750_,
		_w4751_
	);
	LUT4 #(
		.INIT('h1311)
	) name4289 (
		_w2182_,
		_w4737_,
		_w4740_,
		_w4751_,
		_w4752_
	);
	LUT3 #(
		.INIT('hce)
	) name4290 (
		\P1_state_reg[0]/NET0131 ,
		_w4736_,
		_w4752_,
		_w4753_
	);
	LUT2 #(
		.INIT('h2)
	) name4291 (
		\P2_reg0_reg[9]/NET0131 ,
		_w2042_,
		_w4754_
	);
	LUT4 #(
		.INIT('h2000)
	) name4292 (
		\P2_reg0_reg[9]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4755_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4293 (
		\P2_reg0_reg[9]/NET0131 ,
		_w2729_,
		_w4150_,
		_w4151_,
		_w4756_
	);
	LUT2 #(
		.INIT('h2)
	) name4294 (
		_w2000_,
		_w4756_,
		_w4757_
	);
	LUT4 #(
		.INIT('hc355)
	) name4295 (
		\P2_reg0_reg[9]/NET0131 ,
		_w1905_,
		_w2484_,
		_w2729_,
		_w4758_
	);
	LUT4 #(
		.INIT('hc808)
	) name4296 (
		\P2_reg0_reg[9]/NET0131 ,
		_w1869_,
		_w2729_,
		_w4155_,
		_w4759_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4297 (
		\P2_reg0_reg[9]/NET0131 ,
		_w2033_,
		_w2729_,
		_w2734_,
		_w4760_
	);
	LUT3 #(
		.INIT('h0d)
	) name4298 (
		_w2729_,
		_w4158_,
		_w4760_,
		_w4761_
	);
	LUT4 #(
		.INIT('h3100)
	) name4299 (
		_w1963_,
		_w4759_,
		_w4758_,
		_w4761_,
		_w4762_
	);
	LUT4 #(
		.INIT('h1311)
	) name4300 (
		_w1285_,
		_w4755_,
		_w4757_,
		_w4762_,
		_w4763_
	);
	LUT3 #(
		.INIT('hce)
	) name4301 (
		\P1_state_reg[0]/NET0131 ,
		_w4754_,
		_w4763_,
		_w4764_
	);
	LUT2 #(
		.INIT('h2)
	) name4302 (
		\P2_reg1_reg[10]/NET0131 ,
		_w2042_,
		_w4765_
	);
	LUT4 #(
		.INIT('h2000)
	) name4303 (
		\P2_reg1_reg[10]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4766_
	);
	LUT2 #(
		.INIT('h2)
	) name4304 (
		\P2_reg1_reg[10]/NET0131 ,
		_w2762_,
		_w4767_
	);
	LUT4 #(
		.INIT('h7020)
	) name4305 (
		_w1305_,
		_w1779_,
		_w2762_,
		_w4088_,
		_w4768_
	);
	LUT3 #(
		.INIT('ha8)
	) name4306 (
		_w2000_,
		_w4767_,
		_w4768_,
		_w4769_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4307 (
		\P2_reg1_reg[10]/NET0131 ,
		_w1963_,
		_w2762_,
		_w4091_,
		_w4770_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4308 (
		\P2_reg1_reg[10]/NET0131 ,
		_w2483_,
		_w2762_,
		_w3095_,
		_w4771_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4309 (
		\P2_reg1_reg[10]/NET0131 ,
		_w2033_,
		_w2734_,
		_w2762_,
		_w4772_
	);
	LUT3 #(
		.INIT('h10)
	) name4310 (
		_w1769_,
		_w1773_,
		_w2001_,
		_w4773_
	);
	LUT4 #(
		.INIT('h007b)
	) name4311 (
		_w1774_,
		_w2025_,
		_w4094_,
		_w4773_,
		_w4774_
	);
	LUT3 #(
		.INIT('h31)
	) name4312 (
		_w2762_,
		_w4772_,
		_w4774_,
		_w4775_
	);
	LUT3 #(
		.INIT('hd0)
	) name4313 (
		_w1869_,
		_w4771_,
		_w4775_,
		_w4776_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4314 (
		_w1285_,
		_w4770_,
		_w4769_,
		_w4776_,
		_w4777_
	);
	LUT4 #(
		.INIT('heeec)
	) name4315 (
		\P1_state_reg[0]/NET0131 ,
		_w4765_,
		_w4766_,
		_w4777_,
		_w4778_
	);
	LUT2 #(
		.INIT('h2)
	) name4316 (
		\P2_reg1_reg[13]/NET0131 ,
		_w2042_,
		_w4779_
	);
	LUT4 #(
		.INIT('h2000)
	) name4317 (
		\P2_reg1_reg[13]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4780_
	);
	LUT2 #(
		.INIT('h2)
	) name4318 (
		\P2_reg1_reg[13]/NET0131 ,
		_w2762_,
		_w4781_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4319 (
		\P2_reg1_reg[13]/NET0131 ,
		_w2762_,
		_w4107_,
		_w4108_,
		_w4782_
	);
	LUT2 #(
		.INIT('h2)
	) name4320 (
		_w2000_,
		_w4782_,
		_w4783_
	);
	LUT4 #(
		.INIT('h40b0)
	) name4321 (
		_w1792_,
		_w1797_,
		_w2762_,
		_w4111_,
		_w4784_
	);
	LUT3 #(
		.INIT('ha8)
	) name4322 (
		_w1869_,
		_w4781_,
		_w4784_,
		_w4785_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4323 (
		\P2_reg1_reg[13]/NET0131 ,
		_w1963_,
		_w2762_,
		_w4114_,
		_w4786_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4324 (
		\P2_reg1_reg[13]/NET0131 ,
		_w2033_,
		_w2734_,
		_w2762_,
		_w4787_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4325 (
		_w2762_,
		_w4116_,
		_w4118_,
		_w4787_,
		_w4788_
	);
	LUT3 #(
		.INIT('h10)
	) name4326 (
		_w4786_,
		_w4785_,
		_w4788_,
		_w4789_
	);
	LUT4 #(
		.INIT('h1311)
	) name4327 (
		_w1285_,
		_w4780_,
		_w4783_,
		_w4789_,
		_w4790_
	);
	LUT3 #(
		.INIT('hce)
	) name4328 (
		\P1_state_reg[0]/NET0131 ,
		_w4779_,
		_w4790_,
		_w4791_
	);
	LUT2 #(
		.INIT('h2)
	) name4329 (
		\P2_reg1_reg[15]/NET0131 ,
		_w2042_,
		_w4792_
	);
	LUT4 #(
		.INIT('h2000)
	) name4330 (
		\P2_reg1_reg[15]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4793_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4331 (
		\P2_reg1_reg[15]/NET0131 ,
		_w2762_,
		_w4130_,
		_w4131_,
		_w4794_
	);
	LUT2 #(
		.INIT('h2)
	) name4332 (
		_w2000_,
		_w4794_,
		_w4795_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4333 (
		\P2_reg1_reg[15]/NET0131 ,
		_w2493_,
		_w2762_,
		_w4134_,
		_w4796_
	);
	LUT2 #(
		.INIT('h8)
	) name4334 (
		_w1820_,
		_w2001_,
		_w4797_
	);
	LUT4 #(
		.INIT('h007b)
	) name4335 (
		_w1820_,
		_w2025_,
		_w3716_,
		_w4797_,
		_w4798_
	);
	LUT4 #(
		.INIT('h08cc)
	) name4336 (
		_w1963_,
		_w2762_,
		_w4136_,
		_w4798_,
		_w4799_
	);
	LUT2 #(
		.INIT('h2)
	) name4337 (
		\P2_reg1_reg[15]/NET0131 ,
		_w3872_,
		_w4800_
	);
	LUT4 #(
		.INIT('h0301)
	) name4338 (
		_w1869_,
		_w4799_,
		_w4800_,
		_w4796_,
		_w4801_
	);
	LUT4 #(
		.INIT('h1311)
	) name4339 (
		_w1285_,
		_w4793_,
		_w4795_,
		_w4801_,
		_w4802_
	);
	LUT3 #(
		.INIT('hce)
	) name4340 (
		\P1_state_reg[0]/NET0131 ,
		_w4792_,
		_w4802_,
		_w4803_
	);
	LUT2 #(
		.INIT('h2)
	) name4341 (
		\P2_reg1_reg[23]/NET0131 ,
		_w2042_,
		_w4804_
	);
	LUT4 #(
		.INIT('h2000)
	) name4342 (
		\P2_reg1_reg[23]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4805_
	);
	LUT4 #(
		.INIT('hc535)
	) name4343 (
		\P2_reg1_reg[23]/NET0131 ,
		_w2505_,
		_w2762_,
		_w4245_,
		_w4806_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4344 (
		\P2_reg1_reg[23]/NET0131 ,
		_w1869_,
		_w2762_,
		_w4250_,
		_w4807_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4345 (
		\P2_reg1_reg[23]/NET0131 ,
		_w2762_,
		_w4252_,
		_w4253_,
		_w4808_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4346 (
		\P2_reg1_reg[23]/NET0131 ,
		_w2033_,
		_w2734_,
		_w2762_,
		_w4809_
	);
	LUT4 #(
		.INIT('haa20)
	) name4347 (
		_w2762_,
		_w4255_,
		_w4256_,
		_w4424_,
		_w4810_
	);
	LUT4 #(
		.INIT('h0031)
	) name4348 (
		_w2000_,
		_w4809_,
		_w4808_,
		_w4810_,
		_w4811_
	);
	LUT4 #(
		.INIT('h3100)
	) name4349 (
		_w1963_,
		_w4807_,
		_w4806_,
		_w4811_,
		_w4812_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4350 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w4805_,
		_w4812_,
		_w4813_
	);
	LUT2 #(
		.INIT('he)
	) name4351 (
		_w4804_,
		_w4813_,
		_w4814_
	);
	LUT2 #(
		.INIT('h2)
	) name4352 (
		\P2_reg1_reg[9]/NET0131 ,
		_w2042_,
		_w4815_
	);
	LUT4 #(
		.INIT('h2000)
	) name4353 (
		\P2_reg1_reg[9]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4816_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4354 (
		\P2_reg1_reg[9]/NET0131 ,
		_w2762_,
		_w4150_,
		_w4151_,
		_w4817_
	);
	LUT2 #(
		.INIT('h2)
	) name4355 (
		_w2000_,
		_w4817_,
		_w4818_
	);
	LUT4 #(
		.INIT('hc355)
	) name4356 (
		\P2_reg1_reg[9]/NET0131 ,
		_w1905_,
		_w2484_,
		_w2762_,
		_w4819_
	);
	LUT4 #(
		.INIT('hc808)
	) name4357 (
		\P2_reg1_reg[9]/NET0131 ,
		_w1869_,
		_w2762_,
		_w4155_,
		_w4820_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4358 (
		\P2_reg1_reg[9]/NET0131 ,
		_w2033_,
		_w2734_,
		_w2762_,
		_w4821_
	);
	LUT3 #(
		.INIT('h0d)
	) name4359 (
		_w2762_,
		_w4158_,
		_w4821_,
		_w4822_
	);
	LUT4 #(
		.INIT('h3100)
	) name4360 (
		_w1963_,
		_w4820_,
		_w4819_,
		_w4822_,
		_w4823_
	);
	LUT4 #(
		.INIT('h1311)
	) name4361 (
		_w1285_,
		_w4816_,
		_w4818_,
		_w4823_,
		_w4824_
	);
	LUT3 #(
		.INIT('hce)
	) name4362 (
		\P1_state_reg[0]/NET0131 ,
		_w4815_,
		_w4824_,
		_w4825_
	);
	LUT2 #(
		.INIT('h2)
	) name4363 (
		\P2_reg2_reg[10]/NET0131 ,
		_w2042_,
		_w4826_
	);
	LUT4 #(
		.INIT('h2000)
	) name4364 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4827_
	);
	LUT2 #(
		.INIT('h2)
	) name4365 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1298_,
		_w4828_
	);
	LUT4 #(
		.INIT('h2a08)
	) name4366 (
		_w1298_,
		_w1305_,
		_w1779_,
		_w4088_,
		_w4829_
	);
	LUT3 #(
		.INIT('ha8)
	) name4367 (
		_w2000_,
		_w4828_,
		_w4829_,
		_w4830_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4368 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1298_,
		_w1963_,
		_w4091_,
		_w4831_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4369 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1298_,
		_w2483_,
		_w3095_,
		_w4832_
	);
	LUT4 #(
		.INIT('h0200)
	) name4370 (
		_w1762_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w4833_
	);
	LUT3 #(
		.INIT('h0d)
	) name4371 (
		\P2_reg2_reg[10]/NET0131 ,
		_w2640_,
		_w4833_,
		_w4834_
	);
	LUT3 #(
		.INIT('hd0)
	) name4372 (
		_w1298_,
		_w4774_,
		_w4834_,
		_w4835_
	);
	LUT3 #(
		.INIT('hd0)
	) name4373 (
		_w1869_,
		_w4832_,
		_w4835_,
		_w4836_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4374 (
		_w1285_,
		_w4831_,
		_w4830_,
		_w4836_,
		_w4837_
	);
	LUT4 #(
		.INIT('heeec)
	) name4375 (
		\P1_state_reg[0]/NET0131 ,
		_w4826_,
		_w4827_,
		_w4837_,
		_w4838_
	);
	LUT2 #(
		.INIT('h2)
	) name4376 (
		\P2_reg2_reg[13]/NET0131 ,
		_w2042_,
		_w4839_
	);
	LUT4 #(
		.INIT('h2000)
	) name4377 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4840_
	);
	LUT2 #(
		.INIT('h2)
	) name4378 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1298_,
		_w4841_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4379 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1298_,
		_w4107_,
		_w4108_,
		_w4842_
	);
	LUT2 #(
		.INIT('h2)
	) name4380 (
		_w2000_,
		_w4842_,
		_w4843_
	);
	LUT4 #(
		.INIT('h208a)
	) name4381 (
		_w1298_,
		_w1792_,
		_w1797_,
		_w4111_,
		_w4844_
	);
	LUT3 #(
		.INIT('ha8)
	) name4382 (
		_w1869_,
		_w4841_,
		_w4844_,
		_w4845_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4383 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1298_,
		_w1963_,
		_w4114_,
		_w4846_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name4384 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1298_,
		_w2032_,
		_w2033_,
		_w4847_
	);
	LUT4 #(
		.INIT('h0200)
	) name4385 (
		_w1831_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w4848_
	);
	LUT2 #(
		.INIT('h1)
	) name4386 (
		_w4847_,
		_w4848_,
		_w4849_
	);
	LUT4 #(
		.INIT('hfd00)
	) name4387 (
		_w1298_,
		_w4116_,
		_w4118_,
		_w4849_,
		_w4850_
	);
	LUT3 #(
		.INIT('h10)
	) name4388 (
		_w4846_,
		_w4845_,
		_w4850_,
		_w4851_
	);
	LUT4 #(
		.INIT('h1311)
	) name4389 (
		_w1285_,
		_w4840_,
		_w4843_,
		_w4851_,
		_w4852_
	);
	LUT3 #(
		.INIT('hce)
	) name4390 (
		\P1_state_reg[0]/NET0131 ,
		_w4839_,
		_w4852_,
		_w4853_
	);
	LUT2 #(
		.INIT('h2)
	) name4391 (
		\P2_reg2_reg[15]/NET0131 ,
		_w2042_,
		_w4854_
	);
	LUT4 #(
		.INIT('h2000)
	) name4392 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4855_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4393 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1298_,
		_w4130_,
		_w4131_,
		_w4856_
	);
	LUT2 #(
		.INIT('h2)
	) name4394 (
		_w2000_,
		_w4856_,
		_w4857_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4395 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1298_,
		_w2493_,
		_w4134_,
		_w4858_
	);
	LUT2 #(
		.INIT('h2)
	) name4396 (
		_w1869_,
		_w4858_,
		_w4859_
	);
	LUT2 #(
		.INIT('h2)
	) name4397 (
		_w1298_,
		_w4798_,
		_w4860_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4398 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1298_,
		_w1963_,
		_w4136_,
		_w4861_
	);
	LUT4 #(
		.INIT('h0200)
	) name4399 (
		_w1810_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w4862_
	);
	LUT3 #(
		.INIT('h0d)
	) name4400 (
		\P2_reg2_reg[15]/NET0131 ,
		_w2640_,
		_w4862_,
		_w4863_
	);
	LUT3 #(
		.INIT('h10)
	) name4401 (
		_w4861_,
		_w4860_,
		_w4863_,
		_w4864_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4402 (
		_w1285_,
		_w4859_,
		_w4857_,
		_w4864_,
		_w4865_
	);
	LUT4 #(
		.INIT('heeec)
	) name4403 (
		\P1_state_reg[0]/NET0131 ,
		_w4854_,
		_w4855_,
		_w4865_,
		_w4866_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4404 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[9]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4867_
	);
	LUT2 #(
		.INIT('h8)
	) name4405 (
		\P1_reg2_reg[9]/NET0131 ,
		_w2183_,
		_w4868_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4406 (
		\P1_reg2_reg[9]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4869_
	);
	LUT4 #(
		.INIT('hc808)
	) name4407 (
		\P1_reg2_reg[9]/NET0131 ,
		_w1237_,
		_w2189_,
		_w3733_,
		_w4870_
	);
	LUT4 #(
		.INIT('hc808)
	) name4408 (
		\P1_reg2_reg[9]/NET0131 ,
		_w2121_,
		_w2189_,
		_w3735_,
		_w4871_
	);
	LUT4 #(
		.INIT('h8488)
	) name4409 (
		_w1173_,
		_w2189_,
		_w2236_,
		_w2239_,
		_w4872_
	);
	LUT4 #(
		.INIT('h2a00)
	) name4410 (
		_w905_,
		_w915_,
		_w2159_,
		_w2170_,
		_w4873_
	);
	LUT2 #(
		.INIT('h4)
	) name4411 (
		_w905_,
		_w2172_,
		_w4874_
	);
	LUT4 #(
		.INIT('hea00)
	) name4412 (
		_w1100_,
		_w915_,
		_w2159_,
		_w4874_,
		_w4875_
	);
	LUT4 #(
		.INIT('h1000)
	) name4413 (
		_w1096_,
		_w1098_,
		_w897_,
		_w1101_,
		_w4876_
	);
	LUT4 #(
		.INIT('h0057)
	) name4414 (
		\P1_reg2_reg[9]/NET0131 ,
		_w2171_,
		_w3173_,
		_w4876_,
		_w4877_
	);
	LUT4 #(
		.INIT('h5700)
	) name4415 (
		_w2189_,
		_w4873_,
		_w4875_,
		_w4877_,
		_w4878_
	);
	LUT4 #(
		.INIT('h5700)
	) name4416 (
		_w2128_,
		_w4869_,
		_w4872_,
		_w4878_,
		_w4879_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4417 (
		_w2182_,
		_w4870_,
		_w4871_,
		_w4879_,
		_w4880_
	);
	LUT4 #(
		.INIT('heeec)
	) name4418 (
		\P1_state_reg[0]/NET0131 ,
		_w4867_,
		_w4868_,
		_w4880_,
		_w4881_
	);
	LUT2 #(
		.INIT('h2)
	) name4419 (
		\P2_reg2_reg[9]/NET0131 ,
		_w2042_,
		_w4882_
	);
	LUT4 #(
		.INIT('h2000)
	) name4420 (
		\P2_reg2_reg[9]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4883_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4421 (
		\P2_reg2_reg[9]/NET0131 ,
		_w1298_,
		_w4150_,
		_w4151_,
		_w4884_
	);
	LUT2 #(
		.INIT('h2)
	) name4422 (
		_w2000_,
		_w4884_,
		_w4885_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4423 (
		\P2_reg2_reg[9]/NET0131 ,
		_w1298_,
		_w1905_,
		_w2484_,
		_w4886_
	);
	LUT4 #(
		.INIT('he020)
	) name4424 (
		\P2_reg2_reg[9]/NET0131 ,
		_w1298_,
		_w1869_,
		_w4155_,
		_w4887_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name4425 (
		\P2_reg2_reg[9]/NET0131 ,
		_w1298_,
		_w2032_,
		_w2033_,
		_w4888_
	);
	LUT4 #(
		.INIT('h0200)
	) name4426 (
		_w1776_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w4889_
	);
	LUT2 #(
		.INIT('h1)
	) name4427 (
		_w4888_,
		_w4889_,
		_w4890_
	);
	LUT3 #(
		.INIT('hd0)
	) name4428 (
		_w1298_,
		_w4158_,
		_w4890_,
		_w4891_
	);
	LUT4 #(
		.INIT('h3100)
	) name4429 (
		_w1963_,
		_w4887_,
		_w4886_,
		_w4891_,
		_w4892_
	);
	LUT4 #(
		.INIT('h1311)
	) name4430 (
		_w1285_,
		_w4883_,
		_w4885_,
		_w4892_,
		_w4893_
	);
	LUT3 #(
		.INIT('hce)
	) name4431 (
		\P1_state_reg[0]/NET0131 ,
		_w4882_,
		_w4893_,
		_w4894_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4432 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[15]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4895_
	);
	LUT2 #(
		.INIT('h8)
	) name4433 (
		\P1_reg0_reg[15]/NET0131 ,
		_w2183_,
		_w4896_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4434 (
		\P1_reg0_reg[15]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4897_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4435 (
		\P1_reg0_reg[15]/NET0131 ,
		_w1168_,
		_w2325_,
		_w4066_,
		_w4898_
	);
	LUT2 #(
		.INIT('h2)
	) name4436 (
		_w2121_,
		_w4898_,
		_w4899_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4437 (
		\P1_reg0_reg[15]/NET0131 ,
		_w2128_,
		_w2325_,
		_w4069_,
		_w4900_
	);
	LUT4 #(
		.INIT('h7020)
	) name4438 (
		_w488_,
		_w837_,
		_w2325_,
		_w4071_,
		_w4901_
	);
	LUT3 #(
		.INIT('ha8)
	) name4439 (
		_w1237_,
		_w4897_,
		_w4901_,
		_w4902_
	);
	LUT4 #(
		.INIT('hc808)
	) name4440 (
		\P1_reg0_reg[15]/NET0131 ,
		_w2170_,
		_w2325_,
		_w4074_,
		_w4903_
	);
	LUT2 #(
		.INIT('h8)
	) name4441 (
		_w2325_,
		_w4745_,
		_w4904_
	);
	LUT3 #(
		.INIT('ha2)
	) name4442 (
		\P1_reg0_reg[15]/NET0131 ,
		_w2332_,
		_w2333_,
		_w4905_
	);
	LUT2 #(
		.INIT('h1)
	) name4443 (
		_w4904_,
		_w4905_,
		_w4906_
	);
	LUT2 #(
		.INIT('h4)
	) name4444 (
		_w4903_,
		_w4906_,
		_w4907_
	);
	LUT3 #(
		.INIT('h10)
	) name4445 (
		_w4902_,
		_w4900_,
		_w4907_,
		_w4908_
	);
	LUT4 #(
		.INIT('h1311)
	) name4446 (
		_w2182_,
		_w4896_,
		_w4899_,
		_w4908_,
		_w4909_
	);
	LUT3 #(
		.INIT('hce)
	) name4447 (
		\P1_state_reg[0]/NET0131 ,
		_w4895_,
		_w4909_,
		_w4910_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4448 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[15]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4911_
	);
	LUT2 #(
		.INIT('h8)
	) name4449 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2183_,
		_w4912_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4450 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4913_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4451 (
		\P1_reg1_reg[15]/NET0131 ,
		_w1168_,
		_w2536_,
		_w4066_,
		_w4914_
	);
	LUT2 #(
		.INIT('h2)
	) name4452 (
		_w2121_,
		_w4914_,
		_w4915_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4453 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2128_,
		_w2536_,
		_w4069_,
		_w4916_
	);
	LUT4 #(
		.INIT('h7020)
	) name4454 (
		_w488_,
		_w837_,
		_w2536_,
		_w4071_,
		_w4917_
	);
	LUT3 #(
		.INIT('ha8)
	) name4455 (
		_w1237_,
		_w4913_,
		_w4917_,
		_w4918_
	);
	LUT4 #(
		.INIT('hc808)
	) name4456 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2170_,
		_w2536_,
		_w4074_,
		_w4919_
	);
	LUT3 #(
		.INIT('ha2)
	) name4457 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2332_,
		_w2544_,
		_w4920_
	);
	LUT2 #(
		.INIT('h8)
	) name4458 (
		_w2536_,
		_w4745_,
		_w4921_
	);
	LUT2 #(
		.INIT('h1)
	) name4459 (
		_w4920_,
		_w4921_,
		_w4922_
	);
	LUT2 #(
		.INIT('h4)
	) name4460 (
		_w4919_,
		_w4922_,
		_w4923_
	);
	LUT3 #(
		.INIT('h10)
	) name4461 (
		_w4918_,
		_w4916_,
		_w4923_,
		_w4924_
	);
	LUT4 #(
		.INIT('h1311)
	) name4462 (
		_w2182_,
		_w4912_,
		_w4915_,
		_w4924_,
		_w4925_
	);
	LUT3 #(
		.INIT('hce)
	) name4463 (
		\P1_state_reg[0]/NET0131 ,
		_w4911_,
		_w4925_,
		_w4926_
	);
	LUT2 #(
		.INIT('h2)
	) name4464 (
		\P2_reg0_reg[10]/NET0131 ,
		_w2042_,
		_w4927_
	);
	LUT4 #(
		.INIT('h2000)
	) name4465 (
		\P2_reg0_reg[10]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4928_
	);
	LUT2 #(
		.INIT('h2)
	) name4466 (
		\P2_reg0_reg[10]/NET0131 ,
		_w2729_,
		_w4929_
	);
	LUT4 #(
		.INIT('h7020)
	) name4467 (
		_w1305_,
		_w1779_,
		_w2729_,
		_w4088_,
		_w4930_
	);
	LUT3 #(
		.INIT('ha8)
	) name4468 (
		_w2000_,
		_w4929_,
		_w4930_,
		_w4931_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4469 (
		\P2_reg0_reg[10]/NET0131 ,
		_w1963_,
		_w2729_,
		_w4091_,
		_w4932_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4470 (
		\P2_reg0_reg[10]/NET0131 ,
		_w2483_,
		_w2729_,
		_w3095_,
		_w4933_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4471 (
		\P2_reg0_reg[10]/NET0131 ,
		_w2033_,
		_w2729_,
		_w2734_,
		_w4934_
	);
	LUT3 #(
		.INIT('h0d)
	) name4472 (
		_w2729_,
		_w4774_,
		_w4934_,
		_w4935_
	);
	LUT3 #(
		.INIT('hd0)
	) name4473 (
		_w1869_,
		_w4933_,
		_w4935_,
		_w4936_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4474 (
		_w1285_,
		_w4932_,
		_w4931_,
		_w4936_,
		_w4937_
	);
	LUT4 #(
		.INIT('heeec)
	) name4475 (
		\P1_state_reg[0]/NET0131 ,
		_w4927_,
		_w4928_,
		_w4937_,
		_w4938_
	);
	LUT2 #(
		.INIT('h2)
	) name4476 (
		\P2_reg0_reg[13]/NET0131 ,
		_w2042_,
		_w4939_
	);
	LUT4 #(
		.INIT('h2000)
	) name4477 (
		\P2_reg0_reg[13]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4940_
	);
	LUT2 #(
		.INIT('h2)
	) name4478 (
		\P2_reg0_reg[13]/NET0131 ,
		_w2729_,
		_w4941_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4479 (
		\P2_reg0_reg[13]/NET0131 ,
		_w2729_,
		_w4107_,
		_w4108_,
		_w4942_
	);
	LUT2 #(
		.INIT('h2)
	) name4480 (
		_w2000_,
		_w4942_,
		_w4943_
	);
	LUT4 #(
		.INIT('h40b0)
	) name4481 (
		_w1792_,
		_w1797_,
		_w2729_,
		_w4111_,
		_w4944_
	);
	LUT3 #(
		.INIT('ha8)
	) name4482 (
		_w1869_,
		_w4941_,
		_w4944_,
		_w4945_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4483 (
		\P2_reg0_reg[13]/NET0131 ,
		_w1963_,
		_w2729_,
		_w4114_,
		_w4946_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4484 (
		\P2_reg0_reg[13]/NET0131 ,
		_w2033_,
		_w2729_,
		_w2734_,
		_w4947_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4485 (
		_w2729_,
		_w4116_,
		_w4118_,
		_w4947_,
		_w4948_
	);
	LUT3 #(
		.INIT('h10)
	) name4486 (
		_w4946_,
		_w4945_,
		_w4948_,
		_w4949_
	);
	LUT4 #(
		.INIT('h1311)
	) name4487 (
		_w1285_,
		_w4940_,
		_w4943_,
		_w4949_,
		_w4950_
	);
	LUT3 #(
		.INIT('hce)
	) name4488 (
		\P1_state_reg[0]/NET0131 ,
		_w4939_,
		_w4950_,
		_w4951_
	);
	LUT2 #(
		.INIT('h2)
	) name4489 (
		\P2_reg0_reg[15]/NET0131 ,
		_w2042_,
		_w4952_
	);
	LUT4 #(
		.INIT('h2000)
	) name4490 (
		\P2_reg0_reg[15]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w4953_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4491 (
		\P2_reg0_reg[15]/NET0131 ,
		_w2729_,
		_w4130_,
		_w4131_,
		_w4954_
	);
	LUT2 #(
		.INIT('h2)
	) name4492 (
		_w2000_,
		_w4954_,
		_w4955_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4493 (
		\P2_reg0_reg[15]/NET0131 ,
		_w2493_,
		_w2729_,
		_w4134_,
		_w4956_
	);
	LUT2 #(
		.INIT('h2)
	) name4494 (
		\P2_reg0_reg[15]/NET0131 ,
		_w3982_,
		_w4957_
	);
	LUT4 #(
		.INIT('h08cc)
	) name4495 (
		_w1963_,
		_w2729_,
		_w4136_,
		_w4798_,
		_w4958_
	);
	LUT4 #(
		.INIT('h0301)
	) name4496 (
		_w1869_,
		_w4957_,
		_w4958_,
		_w4956_,
		_w4959_
	);
	LUT4 #(
		.INIT('h1311)
	) name4497 (
		_w1285_,
		_w4953_,
		_w4955_,
		_w4959_,
		_w4960_
	);
	LUT3 #(
		.INIT('hce)
	) name4498 (
		\P1_state_reg[0]/NET0131 ,
		_w4952_,
		_w4960_,
		_w4961_
	);
	LUT3 #(
		.INIT('h2a)
	) name4499 (
		\P1_reg1_reg[4]/NET0131 ,
		_w3511_,
		_w3976_,
		_w4962_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4500 (
		_w3608_,
		_w4629_,
		_w4632_,
		_w4635_,
		_w4963_
	);
	LUT2 #(
		.INIT('he)
	) name4501 (
		_w4962_,
		_w4963_,
		_w4964_
	);
	LUT2 #(
		.INIT('h4)
	) name4502 (
		\P1_reg3_reg[3]/NET0131 ,
		_w2183_,
		_w4965_
	);
	LUT4 #(
		.INIT('h4144)
	) name4503 (
		_w488_,
		_w961_,
		_w971_,
		_w2130_,
		_w4966_
	);
	LUT3 #(
		.INIT('h80)
	) name4504 (
		_w488_,
		_w978_,
		_w979_,
		_w4967_
	);
	LUT4 #(
		.INIT('h2220)
	) name4505 (
		\P1_reg3_reg[3]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w4968_
	);
	LUT2 #(
		.INIT('h2)
	) name4506 (
		_w1237_,
		_w4968_,
		_w4969_
	);
	LUT4 #(
		.INIT('h5700)
	) name4507 (
		_w2055_,
		_w4966_,
		_w4967_,
		_w4969_,
		_w4970_
	);
	LUT3 #(
		.INIT('h04)
	) name4508 (
		_w1186_,
		_w2071_,
		_w2270_,
		_w4971_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name4509 (
		_w1187_,
		_w2070_,
		_w2121_,
		_w2270_,
		_w4972_
	);
	LUT4 #(
		.INIT('h3060)
	) name4510 (
		_w985_,
		_w1187_,
		_w2128_,
		_w2229_,
		_w4973_
	);
	LUT4 #(
		.INIT('h1555)
	) name4511 (
		_w976_,
		_w984_,
		_w993_,
		_w1001_,
		_w4974_
	);
	LUT3 #(
		.INIT('h04)
	) name4512 (
		_w2156_,
		_w2170_,
		_w4974_,
		_w4975_
	);
	LUT4 #(
		.INIT('h0045)
	) name4513 (
		_w4973_,
		_w4971_,
		_w4972_,
		_w4975_,
		_w4976_
	);
	LUT3 #(
		.INIT('h10)
	) name4514 (
		_w976_,
		_w2175_,
		_w2176_,
		_w4977_
	);
	LUT4 #(
		.INIT('h5554)
	) name4515 (
		\P1_reg3_reg[3]/NET0131 ,
		_w2171_,
		_w2173_,
		_w4056_,
		_w4978_
	);
	LUT2 #(
		.INIT('h1)
	) name4516 (
		_w4977_,
		_w4978_,
		_w4979_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4517 (
		_w2055_,
		_w4976_,
		_w4970_,
		_w4979_,
		_w4980_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4518 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w4965_,
		_w4980_,
		_w4981_
	);
	LUT2 #(
		.INIT('h2)
	) name4519 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4982_
	);
	LUT4 #(
		.INIT('he3d3)
	) name4520 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg3_reg[3]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w4983_
	);
	LUT2 #(
		.INIT('hb)
	) name4521 (
		_w4981_,
		_w4983_,
		_w4984_
	);
	LUT4 #(
		.INIT('h4000)
	) name4522 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1668_,
		_w4985_
	);
	LUT4 #(
		.INIT('h0100)
	) name4523 (
		_w1722_,
		_w1670_,
		_w1675_,
		_w1969_,
		_w4986_
	);
	LUT4 #(
		.INIT('h5655)
	) name4524 (
		_w1722_,
		_w1670_,
		_w1675_,
		_w1969_,
		_w4987_
	);
	LUT4 #(
		.INIT('h80d0)
	) name4525 (
		_w1305_,
		_w1675_,
		_w2903_,
		_w4987_,
		_w4988_
	);
	LUT3 #(
		.INIT('hc8)
	) name4526 (
		_w1668_,
		_w2000_,
		_w2903_,
		_w4989_
	);
	LUT2 #(
		.INIT('h4)
	) name4527 (
		_w4988_,
		_w4989_,
		_w4990_
	);
	LUT4 #(
		.INIT('h0203)
	) name4528 (
		_w1662_,
		_w1682_,
		_w2488_,
		_w3010_,
		_w4991_
	);
	LUT4 #(
		.INIT('hd0c0)
	) name4529 (
		_w1662_,
		_w1682_,
		_w2488_,
		_w3010_,
		_w4992_
	);
	LUT3 #(
		.INIT('h02)
	) name4530 (
		_w1869_,
		_w4992_,
		_w4991_,
		_w4993_
	);
	LUT3 #(
		.INIT('h60)
	) name4531 (
		_w1666_,
		_w2003_,
		_w2025_,
		_w4994_
	);
	LUT4 #(
		.INIT('h007d)
	) name4532 (
		_w1963_,
		_w2409_,
		_w2488_,
		_w4994_,
		_w4995_
	);
	LUT4 #(
		.INIT('h5450)
	) name4533 (
		_w1666_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w4996_
	);
	LUT3 #(
		.INIT('h0d)
	) name4534 (
		_w1668_,
		_w3444_,
		_w4996_,
		_w4997_
	);
	LUT4 #(
		.INIT('h7500)
	) name4535 (
		_w2903_,
		_w4993_,
		_w4995_,
		_w4997_,
		_w4998_
	);
	LUT4 #(
		.INIT('h1311)
	) name4536 (
		_w1285_,
		_w4985_,
		_w4990_,
		_w4998_,
		_w4999_
	);
	LUT2 #(
		.INIT('h4)
	) name4537 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		_w5000_
	);
	LUT3 #(
		.INIT('h07)
	) name4538 (
		_w1668_,
		_w2344_,
		_w5000_,
		_w5001_
	);
	LUT3 #(
		.INIT('h2f)
	) name4539 (
		\P1_state_reg[0]/NET0131 ,
		_w4999_,
		_w5001_,
		_w5002_
	);
	LUT2 #(
		.INIT('h2)
	) name4540 (
		_w1719_,
		_w2903_,
		_w5003_
	);
	LUT3 #(
		.INIT('h80)
	) name4541 (
		_w1305_,
		_w1667_,
		_w1669_,
		_w5004_
	);
	LUT4 #(
		.INIT('h00eb)
	) name4542 (
		_w1305_,
		_w1712_,
		_w4986_,
		_w5004_,
		_w5005_
	);
	LUT4 #(
		.INIT('hc808)
	) name4543 (
		_w1719_,
		_w2000_,
		_w2903_,
		_w5005_,
		_w5006_
	);
	LUT4 #(
		.INIT('h009f)
	) name4544 (
		_w1687_,
		_w2497_,
		_w2903_,
		_w5003_,
		_w5007_
	);
	LUT4 #(
		.INIT('h0bf4)
	) name4545 (
		_w1884_,
		_w1889_,
		_w1893_,
		_w2497_,
		_w5008_
	);
	LUT4 #(
		.INIT('hc808)
	) name4546 (
		_w1719_,
		_w1963_,
		_w2903_,
		_w5008_,
		_w5009_
	);
	LUT4 #(
		.INIT('h9500)
	) name4547 (
		_w1726_,
		_w1666_,
		_w2003_,
		_w2025_,
		_w5010_
	);
	LUT4 #(
		.INIT('h88a8)
	) name4548 (
		_w1719_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w5011_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name4549 (
		_w1726_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w5012_
	);
	LUT4 #(
		.INIT('h0013)
	) name4550 (
		_w2903_,
		_w5011_,
		_w5010_,
		_w5012_,
		_w5013_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4551 (
		_w1869_,
		_w5007_,
		_w5009_,
		_w5013_,
		_w5014_
	);
	LUT4 #(
		.INIT('h4000)
	) name4552 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1719_,
		_w5015_
	);
	LUT4 #(
		.INIT('h0075)
	) name4553 (
		_w1285_,
		_w5006_,
		_w5014_,
		_w5015_,
		_w5016_
	);
	LUT2 #(
		.INIT('h4)
	) name4554 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		_w5017_
	);
	LUT3 #(
		.INIT('h07)
	) name4555 (
		_w1719_,
		_w2344_,
		_w5017_,
		_w5018_
	);
	LUT3 #(
		.INIT('h2f)
	) name4556 (
		\P1_state_reg[0]/NET0131 ,
		_w5016_,
		_w5018_,
		_w5019_
	);
	LUT4 #(
		.INIT('h4000)
	) name4557 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1698_,
		_w5020_
	);
	LUT2 #(
		.INIT('h2)
	) name4558 (
		_w1698_,
		_w2903_,
		_w5021_
	);
	LUT3 #(
		.INIT('h80)
	) name4559 (
		_w1305_,
		_w1709_,
		_w1711_,
		_w5022_
	);
	LUT4 #(
		.INIT('h00eb)
	) name4560 (
		_w1305_,
		_w1691_,
		_w1972_,
		_w5022_,
		_w5023_
	);
	LUT4 #(
		.INIT('hc808)
	) name4561 (
		_w1698_,
		_w2000_,
		_w2903_,
		_w5023_,
		_w5024_
	);
	LUT4 #(
		.INIT('hd02f)
	) name4562 (
		_w1728_,
		_w1687_,
		_w1732_,
		_w2496_,
		_w5025_
	);
	LUT4 #(
		.INIT('hc808)
	) name4563 (
		_w1698_,
		_w1869_,
		_w2903_,
		_w5025_,
		_w5026_
	);
	LUT4 #(
		.INIT('he100)
	) name4564 (
		_w1897_,
		_w1901_,
		_w2496_,
		_w2903_,
		_w5027_
	);
	LUT4 #(
		.INIT('h9000)
	) name4565 (
		_w1706_,
		_w2005_,
		_w2025_,
		_w2903_,
		_w5028_
	);
	LUT4 #(
		.INIT('h88a8)
	) name4566 (
		_w1698_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w5029_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name4567 (
		_w1706_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w5030_
	);
	LUT2 #(
		.INIT('h1)
	) name4568 (
		_w5029_,
		_w5030_,
		_w5031_
	);
	LUT2 #(
		.INIT('h4)
	) name4569 (
		_w5028_,
		_w5031_,
		_w5032_
	);
	LUT4 #(
		.INIT('h5700)
	) name4570 (
		_w1963_,
		_w5021_,
		_w5027_,
		_w5032_,
		_w5033_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4571 (
		_w1285_,
		_w5026_,
		_w5024_,
		_w5033_,
		_w5034_
	);
	LUT2 #(
		.INIT('h4)
	) name4572 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[7]/NET0131 ,
		_w5035_
	);
	LUT3 #(
		.INIT('h07)
	) name4573 (
		_w1698_,
		_w2344_,
		_w5035_,
		_w5036_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4574 (
		\P1_state_reg[0]/NET0131 ,
		_w5020_,
		_w5034_,
		_w5036_,
		_w5037_
	);
	LUT2 #(
		.INIT('h8)
	) name4575 (
		_w925_,
		_w2183_,
		_w5038_
	);
	LUT4 #(
		.INIT('h4150)
	) name4576 (
		_w488_,
		_w927_,
		_w938_,
		_w4169_,
		_w5039_
	);
	LUT3 #(
		.INIT('h80)
	) name4577 (
		_w488_,
		_w946_,
		_w948_,
		_w5040_
	);
	LUT4 #(
		.INIT('h222a)
	) name4578 (
		_w1237_,
		_w2055_,
		_w5039_,
		_w5040_,
		_w5041_
	);
	LUT3 #(
		.INIT('ha2)
	) name4579 (
		_w925_,
		_w4627_,
		_w5041_,
		_w5042_
	);
	LUT3 #(
		.INIT('h02)
	) name4580 (
		_w1237_,
		_w5039_,
		_w5040_,
		_w5043_
	);
	LUT4 #(
		.INIT('ha900)
	) name4581 (
		_w1181_,
		_w2077_,
		_w2079_,
		_w2121_,
		_w5044_
	);
	LUT4 #(
		.INIT('h4b00)
	) name4582 (
		_w1007_,
		_w1010_,
		_w1181_,
		_w2128_,
		_w5045_
	);
	LUT2 #(
		.INIT('h4)
	) name4583 (
		_w933_,
		_w2194_,
		_w5046_
	);
	LUT4 #(
		.INIT('h8000)
	) name4584 (
		_w933_,
		_w956_,
		_w966_,
		_w2156_,
		_w5047_
	);
	LUT4 #(
		.INIT('h009f)
	) name4585 (
		_w933_,
		_w2157_,
		_w2170_,
		_w5046_,
		_w5048_
	);
	LUT3 #(
		.INIT('h10)
	) name4586 (
		_w5045_,
		_w5044_,
		_w5048_,
		_w5049_
	);
	LUT2 #(
		.INIT('h4)
	) name4587 (
		_w933_,
		_w1120_,
		_w5050_
	);
	LUT4 #(
		.INIT('h0075)
	) name4588 (
		_w2055_,
		_w5043_,
		_w5049_,
		_w5050_,
		_w5051_
	);
	LUT4 #(
		.INIT('h1311)
	) name4589 (
		_w2182_,
		_w5038_,
		_w5042_,
		_w5051_,
		_w5052_
	);
	LUT2 #(
		.INIT('h2)
	) name4590 (
		\P1_reg3_reg[6]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5053_
	);
	LUT4 #(
		.INIT('h4080)
	) name4591 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w925_,
		_w1242_,
		_w5054_
	);
	LUT2 #(
		.INIT('h1)
	) name4592 (
		_w5053_,
		_w5054_,
		_w5055_
	);
	LUT3 #(
		.INIT('h2f)
	) name4593 (
		\P1_state_reg[0]/NET0131 ,
		_w5052_,
		_w5055_,
		_w5056_
	);
	LUT2 #(
		.INIT('h8)
	) name4594 (
		_w936_,
		_w2183_,
		_w5057_
	);
	LUT4 #(
		.INIT('h5655)
	) name4595 (
		_w911_,
		_w927_,
		_w938_,
		_w4169_,
		_w5058_
	);
	LUT4 #(
		.INIT('h7020)
	) name4596 (
		_w488_,
		_w927_,
		_w1237_,
		_w5058_,
		_w5059_
	);
	LUT4 #(
		.INIT('h0015)
	) name4597 (
		_w1184_,
		_w2272_,
		_w2274_,
		_w2277_,
		_w5060_
	);
	LUT4 #(
		.INIT('haa80)
	) name4598 (
		_w1184_,
		_w2272_,
		_w2274_,
		_w2277_,
		_w5061_
	);
	LUT3 #(
		.INIT('h02)
	) name4599 (
		_w2121_,
		_w5061_,
		_w5060_,
		_w5062_
	);
	LUT4 #(
		.INIT('h8884)
	) name4600 (
		_w1184_,
		_w2128_,
		_w2237_,
		_w2935_,
		_w5063_
	);
	LUT4 #(
		.INIT('hab27)
	) name4601 (
		_w943_,
		_w2170_,
		_w2194_,
		_w5047_,
		_w5064_
	);
	LUT2 #(
		.INIT('h4)
	) name4602 (
		_w5063_,
		_w5064_,
		_w5065_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4603 (
		_w2055_,
		_w5059_,
		_w5062_,
		_w5065_,
		_w5066_
	);
	LUT4 #(
		.INIT('h0001)
	) name4604 (
		_w2171_,
		_w2173_,
		_w3791_,
		_w4056_,
		_w5067_
	);
	LUT2 #(
		.INIT('h4)
	) name4605 (
		_w943_,
		_w1120_,
		_w5068_
	);
	LUT3 #(
		.INIT('h0d)
	) name4606 (
		_w936_,
		_w5067_,
		_w5068_,
		_w5069_
	);
	LUT4 #(
		.INIT('h1311)
	) name4607 (
		_w2182_,
		_w5057_,
		_w5066_,
		_w5069_,
		_w5070_
	);
	LUT2 #(
		.INIT('h2)
	) name4608 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5071_
	);
	LUT4 #(
		.INIT('h4080)
	) name4609 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w936_,
		_w1242_,
		_w5072_
	);
	LUT2 #(
		.INIT('h1)
	) name4610 (
		_w5071_,
		_w5072_,
		_w5073_
	);
	LUT3 #(
		.INIT('h2f)
	) name4611 (
		\P1_state_reg[0]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5074_
	);
	LUT2 #(
		.INIT('h2)
	) name4612 (
		\P2_reg0_reg[4]/NET0131 ,
		_w2042_,
		_w5075_
	);
	LUT4 #(
		.INIT('h2000)
	) name4613 (
		\P2_reg0_reg[4]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5076_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4614 (
		\P2_reg0_reg[4]/NET0131 ,
		_w3084_,
		_w3981_,
		_w3983_,
		_w5077_
	);
	LUT2 #(
		.INIT('h4)
	) name4615 (
		_w1666_,
		_w2001_,
		_w5078_
	);
	LUT4 #(
		.INIT('h7020)
	) name4616 (
		_w1305_,
		_w1675_,
		_w2000_,
		_w4987_,
		_w5079_
	);
	LUT4 #(
		.INIT('h0004)
	) name4617 (
		_w4993_,
		_w4995_,
		_w5078_,
		_w5079_,
		_w5080_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4618 (
		_w1285_,
		_w2729_,
		_w5077_,
		_w5080_,
		_w5081_
	);
	LUT4 #(
		.INIT('heeec)
	) name4619 (
		\P1_state_reg[0]/NET0131 ,
		_w5075_,
		_w5076_,
		_w5081_,
		_w5082_
	);
	LUT2 #(
		.INIT('h2)
	) name4620 (
		\P2_reg1_reg[4]/NET0131 ,
		_w2042_,
		_w5083_
	);
	LUT4 #(
		.INIT('h2000)
	) name4621 (
		\P2_reg1_reg[4]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5084_
	);
	LUT3 #(
		.INIT('h2a)
	) name4622 (
		\P2_reg1_reg[4]/NET0131 ,
		_w3872_,
		_w3875_,
		_w5085_
	);
	LUT4 #(
		.INIT('haa08)
	) name4623 (
		_w1285_,
		_w2762_,
		_w5080_,
		_w5085_,
		_w5086_
	);
	LUT4 #(
		.INIT('heeec)
	) name4624 (
		\P1_state_reg[0]/NET0131 ,
		_w5083_,
		_w5084_,
		_w5086_,
		_w5087_
	);
	LUT4 #(
		.INIT('h5545)
	) name4625 (
		\P1_reg2_reg[4]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w5088_
	);
	LUT4 #(
		.INIT('h80d0)
	) name4626 (
		_w488_,
		_w971_,
		_w2189_,
		_w4625_,
		_w5089_
	);
	LUT2 #(
		.INIT('h2)
	) name4627 (
		_w1237_,
		_w5089_,
		_w5090_
	);
	LUT4 #(
		.INIT('h4c44)
	) name4628 (
		_w2189_,
		_w3511_,
		_w4632_,
		_w4635_,
		_w5091_
	);
	LUT4 #(
		.INIT('h1000)
	) name4629 (
		_w1096_,
		_w1098_,
		_w958_,
		_w1101_,
		_w5092_
	);
	LUT4 #(
		.INIT('hfb00)
	) name4630 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w2120_,
		_w5093_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4631 (
		\P1_reg2_reg[4]/NET0131 ,
		_w2171_,
		_w3173_,
		_w5093_,
		_w5094_
	);
	LUT2 #(
		.INIT('h1)
	) name4632 (
		_w5092_,
		_w5094_,
		_w5095_
	);
	LUT4 #(
		.INIT('hba00)
	) name4633 (
		_w5088_,
		_w5090_,
		_w5091_,
		_w5095_,
		_w5096_
	);
	LUT2 #(
		.INIT('h1)
	) name4634 (
		\P1_reg2_reg[4]/NET0131 ,
		_w3511_,
		_w5097_
	);
	LUT2 #(
		.INIT('h1)
	) name4635 (
		_w5096_,
		_w5097_,
		_w5098_
	);
	LUT2 #(
		.INIT('h2)
	) name4636 (
		\P2_reg2_reg[8]/NET0131 ,
		_w2042_,
		_w5099_
	);
	LUT4 #(
		.INIT('h2000)
	) name4637 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5100_
	);
	LUT2 #(
		.INIT('h2)
	) name4638 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1298_,
		_w5101_
	);
	LUT4 #(
		.INIT('h111d)
	) name4639 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1298_,
		_w4644_,
		_w4645_,
		_w5102_
	);
	LUT2 #(
		.INIT('h2)
	) name4640 (
		_w2000_,
		_w5102_,
		_w5103_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4641 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1298_,
		_w2413_,
		_w2499_,
		_w5104_
	);
	LUT4 #(
		.INIT('h2822)
	) name4642 (
		_w1298_,
		_w2499_,
		_w3014_,
		_w3017_,
		_w5105_
	);
	LUT2 #(
		.INIT('h8)
	) name4643 (
		_w1695_,
		_w2001_,
		_w5106_
	);
	LUT4 #(
		.INIT('h0200)
	) name4644 (
		_w1689_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w5107_
	);
	LUT3 #(
		.INIT('h0d)
	) name4645 (
		\P2_reg2_reg[8]/NET0131 ,
		_w2640_,
		_w5107_,
		_w5108_
	);
	LUT4 #(
		.INIT('h5700)
	) name4646 (
		_w1298_,
		_w4650_,
		_w5106_,
		_w5108_,
		_w5109_
	);
	LUT4 #(
		.INIT('h5700)
	) name4647 (
		_w1869_,
		_w5101_,
		_w5105_,
		_w5109_,
		_w5110_
	);
	LUT3 #(
		.INIT('hd0)
	) name4648 (
		_w1963_,
		_w5104_,
		_w5110_,
		_w5111_
	);
	LUT4 #(
		.INIT('h1311)
	) name4649 (
		_w1285_,
		_w5100_,
		_w5103_,
		_w5111_,
		_w5112_
	);
	LUT3 #(
		.INIT('hce)
	) name4650 (
		\P1_state_reg[0]/NET0131 ,
		_w5099_,
		_w5112_,
		_w5113_
	);
	LUT3 #(
		.INIT('h2a)
	) name4651 (
		\P1_reg1_reg[5]/NET0131 ,
		_w3511_,
		_w3976_,
		_w5114_
	);
	LUT3 #(
		.INIT('hf2)
	) name4652 (
		_w3608_,
		_w4671_,
		_w5114_,
		_w5115_
	);
	LUT2 #(
		.INIT('h2)
	) name4653 (
		\P2_reg0_reg[8]/NET0131 ,
		_w2042_,
		_w5116_
	);
	LUT4 #(
		.INIT('h2000)
	) name4654 (
		\P2_reg0_reg[8]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5117_
	);
	LUT2 #(
		.INIT('h2)
	) name4655 (
		\P2_reg0_reg[8]/NET0131 ,
		_w2729_,
		_w5118_
	);
	LUT4 #(
		.INIT('h111d)
	) name4656 (
		\P2_reg0_reg[8]/NET0131 ,
		_w2729_,
		_w4644_,
		_w4645_,
		_w5119_
	);
	LUT2 #(
		.INIT('h2)
	) name4657 (
		_w2000_,
		_w5119_,
		_w5120_
	);
	LUT4 #(
		.INIT('hc355)
	) name4658 (
		\P2_reg0_reg[8]/NET0131 ,
		_w2413_,
		_w2499_,
		_w2729_,
		_w5121_
	);
	LUT4 #(
		.INIT('h4844)
	) name4659 (
		_w2499_,
		_w2729_,
		_w3014_,
		_w3017_,
		_w5122_
	);
	LUT2 #(
		.INIT('h2)
	) name4660 (
		\P2_reg0_reg[8]/NET0131 ,
		_w3084_,
		_w5123_
	);
	LUT4 #(
		.INIT('h0057)
	) name4661 (
		_w2729_,
		_w4650_,
		_w5106_,
		_w5123_,
		_w5124_
	);
	LUT4 #(
		.INIT('h5700)
	) name4662 (
		_w1869_,
		_w5118_,
		_w5122_,
		_w5124_,
		_w5125_
	);
	LUT3 #(
		.INIT('hd0)
	) name4663 (
		_w1963_,
		_w5121_,
		_w5125_,
		_w5126_
	);
	LUT4 #(
		.INIT('h1311)
	) name4664 (
		_w1285_,
		_w5117_,
		_w5120_,
		_w5126_,
		_w5127_
	);
	LUT3 #(
		.INIT('hce)
	) name4665 (
		\P1_state_reg[0]/NET0131 ,
		_w5116_,
		_w5127_,
		_w5128_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4666 (
		\P2_reg1_reg[11]/NET0131 ,
		_w2042_,
		_w3872_,
		_w3891_,
		_w5129_
	);
	LUT3 #(
		.INIT('h02)
	) name4667 (
		_w2000_,
		_w4586_,
		_w4587_,
		_w5130_
	);
	LUT4 #(
		.INIT('h2822)
	) name4668 (
		_w1869_,
		_w2495_,
		_w2614_,
		_w2615_,
		_w5131_
	);
	LUT3 #(
		.INIT('h28)
	) name4669 (
		_w1963_,
		_w2495_,
		_w2593_,
		_w5132_
	);
	LUT4 #(
		.INIT('h2300)
	) name4670 (
		_w1306_,
		_w1745_,
		_w1746_,
		_w2001_,
		_w5133_
	);
	LUT3 #(
		.INIT('h0b)
	) name4671 (
		_w4592_,
		_w4593_,
		_w5133_,
		_w5134_
	);
	LUT3 #(
		.INIT('h10)
	) name4672 (
		_w5131_,
		_w5132_,
		_w5134_,
		_w5135_
	);
	LUT4 #(
		.INIT('hecee)
	) name4673 (
		_w3244_,
		_w5129_,
		_w5130_,
		_w5135_,
		_w5136_
	);
	LUT2 #(
		.INIT('h2)
	) name4674 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2042_,
		_w5137_
	);
	LUT4 #(
		.INIT('h2000)
	) name4675 (
		\P2_reg1_reg[8]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5138_
	);
	LUT2 #(
		.INIT('h2)
	) name4676 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2762_,
		_w5139_
	);
	LUT4 #(
		.INIT('h111d)
	) name4677 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2762_,
		_w4644_,
		_w4645_,
		_w5140_
	);
	LUT2 #(
		.INIT('h2)
	) name4678 (
		_w2000_,
		_w5140_,
		_w5141_
	);
	LUT4 #(
		.INIT('hc355)
	) name4679 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2413_,
		_w2499_,
		_w2762_,
		_w5142_
	);
	LUT4 #(
		.INIT('h4844)
	) name4680 (
		_w2499_,
		_w2762_,
		_w3014_,
		_w3017_,
		_w5143_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4681 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2033_,
		_w2734_,
		_w2762_,
		_w5144_
	);
	LUT4 #(
		.INIT('h0057)
	) name4682 (
		_w2762_,
		_w4650_,
		_w5106_,
		_w5144_,
		_w5145_
	);
	LUT4 #(
		.INIT('h5700)
	) name4683 (
		_w1869_,
		_w5139_,
		_w5143_,
		_w5145_,
		_w5146_
	);
	LUT3 #(
		.INIT('hd0)
	) name4684 (
		_w1963_,
		_w5142_,
		_w5146_,
		_w5147_
	);
	LUT4 #(
		.INIT('h1311)
	) name4685 (
		_w1285_,
		_w5138_,
		_w5141_,
		_w5147_,
		_w5148_
	);
	LUT3 #(
		.INIT('hce)
	) name4686 (
		\P1_state_reg[0]/NET0131 ,
		_w5137_,
		_w5148_,
		_w5149_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4687 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[10]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w5150_
	);
	LUT2 #(
		.INIT('h8)
	) name4688 (
		\P1_reg0_reg[10]/NET0131 ,
		_w2183_,
		_w5151_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4689 (
		\P1_reg0_reg[10]/NET0131 ,
		_w2325_,
		_w4025_,
		_w4026_,
		_w5152_
	);
	LUT2 #(
		.INIT('h2)
	) name4690 (
		_w1237_,
		_w5152_,
		_w5153_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4691 (
		\P1_reg0_reg[10]/NET0131 ,
		_w1178_,
		_w2325_,
		_w2653_,
		_w5154_
	);
	LUT2 #(
		.INIT('h2)
	) name4692 (
		_w2128_,
		_w5154_,
		_w5155_
	);
	LUT4 #(
		.INIT('hc535)
	) name4693 (
		\P1_reg0_reg[10]/NET0131 ,
		_w1178_,
		_w2325_,
		_w2682_,
		_w5156_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4694 (
		\P1_reg0_reg[10]/NET0131 ,
		_w2332_,
		_w2333_,
		_w2796_,
		_w5157_
	);
	LUT4 #(
		.INIT('h0057)
	) name4695 (
		_w2325_,
		_w4032_,
		_w4034_,
		_w5157_,
		_w5158_
	);
	LUT3 #(
		.INIT('hd0)
	) name4696 (
		_w2121_,
		_w5156_,
		_w5158_,
		_w5159_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4697 (
		_w2182_,
		_w5153_,
		_w5155_,
		_w5159_,
		_w5160_
	);
	LUT4 #(
		.INIT('heeec)
	) name4698 (
		\P1_state_reg[0]/NET0131 ,
		_w5150_,
		_w5151_,
		_w5160_,
		_w5161_
	);
	LUT4 #(
		.INIT('h5545)
	) name4699 (
		\P1_reg2_reg[5]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w5162_
	);
	LUT3 #(
		.INIT('ha2)
	) name4700 (
		_w1237_,
		_w2189_,
		_w4663_,
		_w5163_
	);
	LUT4 #(
		.INIT('h4c44)
	) name4701 (
		_w2189_,
		_w3511_,
		_w4666_,
		_w4670_,
		_w5164_
	);
	LUT4 #(
		.INIT('h1000)
	) name4702 (
		_w1096_,
		_w1098_,
		_w947_,
		_w1101_,
		_w5165_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4703 (
		\P1_reg2_reg[5]/NET0131 ,
		_w2171_,
		_w3173_,
		_w5093_,
		_w5166_
	);
	LUT2 #(
		.INIT('h1)
	) name4704 (
		_w5165_,
		_w5166_,
		_w5167_
	);
	LUT4 #(
		.INIT('hba00)
	) name4705 (
		_w5162_,
		_w5163_,
		_w5164_,
		_w5167_,
		_w5168_
	);
	LUT2 #(
		.INIT('h1)
	) name4706 (
		\P1_reg2_reg[5]/NET0131 ,
		_w3511_,
		_w5169_
	);
	LUT2 #(
		.INIT('h1)
	) name4707 (
		_w5168_,
		_w5169_,
		_w5170_
	);
	LUT4 #(
		.INIT('h0200)
	) name4708 (
		_w1737_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w5171_
	);
	LUT4 #(
		.INIT('h0075)
	) name4709 (
		_w1298_,
		_w5130_,
		_w5135_,
		_w5171_,
		_w5172_
	);
	LUT2 #(
		.INIT('h2)
	) name4710 (
		\P2_reg2_reg[11]/NET0131 ,
		_w3920_,
		_w5173_
	);
	LUT3 #(
		.INIT('hf2)
	) name4711 (
		_w2556_,
		_w5172_,
		_w5173_,
		_w5174_
	);
	LUT2 #(
		.INIT('h2)
	) name4712 (
		\P2_reg2_reg[14]/NET0131 ,
		_w2042_,
		_w5175_
	);
	LUT4 #(
		.INIT('h2000)
	) name4713 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5176_
	);
	LUT2 #(
		.INIT('h2)
	) name4714 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1298_,
		_w5177_
	);
	LUT4 #(
		.INIT('ha208)
	) name4715 (
		_w1298_,
		_w3115_,
		_w3491_,
		_w4606_,
		_w5178_
	);
	LUT3 #(
		.INIT('ha8)
	) name4716 (
		_w1963_,
		_w5177_,
		_w5178_,
		_w5179_
	);
	LUT4 #(
		.INIT('he020)
	) name4717 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1298_,
		_w2000_,
		_w4610_,
		_w5180_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4718 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1298_,
		_w1869_,
		_w4612_,
		_w5181_
	);
	LUT4 #(
		.INIT('h2300)
	) name4719 (
		_w1306_,
		_w1828_,
		_w1829_,
		_w2001_,
		_w5182_
	);
	LUT4 #(
		.INIT('h0200)
	) name4720 (
		_w1823_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w5183_
	);
	LUT3 #(
		.INIT('h0d)
	) name4721 (
		\P2_reg2_reg[14]/NET0131 ,
		_w2640_,
		_w5183_,
		_w5184_
	);
	LUT4 #(
		.INIT('h5700)
	) name4722 (
		_w1298_,
		_w4614_,
		_w5182_,
		_w5184_,
		_w5185_
	);
	LUT3 #(
		.INIT('h10)
	) name4723 (
		_w5181_,
		_w5180_,
		_w5185_,
		_w5186_
	);
	LUT4 #(
		.INIT('h1311)
	) name4724 (
		_w1285_,
		_w5176_,
		_w5179_,
		_w5186_,
		_w5187_
	);
	LUT3 #(
		.INIT('hce)
	) name4725 (
		\P1_state_reg[0]/NET0131 ,
		_w5175_,
		_w5187_,
		_w5188_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4726 (
		\P1_reg0_reg[11]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w5189_
	);
	LUT4 #(
		.INIT('h7020)
	) name4727 (
		_w488_,
		_w889_,
		_w2325_,
		_w4004_,
		_w5190_
	);
	LUT3 #(
		.INIT('ha8)
	) name4728 (
		_w1237_,
		_w5189_,
		_w5190_,
		_w5191_
	);
	LUT4 #(
		.INIT('h8488)
	) name4729 (
		_w1174_,
		_w2325_,
		_w2962_,
		_w2963_,
		_w5192_
	);
	LUT3 #(
		.INIT('ha8)
	) name4730 (
		_w2121_,
		_w5189_,
		_w5192_,
		_w5193_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4731 (
		\P1_reg0_reg[11]/NET0131 ,
		_w2332_,
		_w2798_,
		_w3560_,
		_w5194_
	);
	LUT3 #(
		.INIT('h0d)
	) name4732 (
		_w2325_,
		_w4013_,
		_w5194_,
		_w5195_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4733 (
		_w2182_,
		_w5191_,
		_w5193_,
		_w5195_,
		_w5196_
	);
	LUT2 #(
		.INIT('h8)
	) name4734 (
		\P1_reg0_reg[11]/NET0131 ,
		_w2183_,
		_w5197_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4735 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[11]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w5198_
	);
	LUT4 #(
		.INIT('hffa8)
	) name4736 (
		\P1_state_reg[0]/NET0131 ,
		_w5196_,
		_w5197_,
		_w5198_,
		_w5199_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4737 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[13]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w5200_
	);
	LUT2 #(
		.INIT('h8)
	) name4738 (
		\P1_reg0_reg[13]/NET0131 ,
		_w2183_,
		_w5201_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4739 (
		\P1_reg0_reg[13]/NET0131 ,
		_w2332_,
		_w2333_,
		_w3567_,
		_w5202_
	);
	LUT4 #(
		.INIT('h0075)
	) name4740 (
		_w2325_,
		_w4721_,
		_w4723_,
		_w5202_,
		_w5203_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4741 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w5201_,
		_w5203_,
		_w5204_
	);
	LUT2 #(
		.INIT('he)
	) name4742 (
		_w5200_,
		_w5204_,
		_w5205_
	);
	LUT4 #(
		.INIT('h0020)
	) name4743 (
		_w2332_,
		_w2333_,
		_w3511_,
		_w3567_,
		_w5206_
	);
	LUT2 #(
		.INIT('h2)
	) name4744 (
		\P1_reg0_reg[14]/NET0131 ,
		_w5206_,
		_w5207_
	);
	LUT3 #(
		.INIT('hf2)
	) name4745 (
		_w3563_,
		_w4730_,
		_w5207_,
		_w5208_
	);
	LUT3 #(
		.INIT('h2a)
	) name4746 (
		\P1_reg0_reg[4]/NET0131 ,
		_w3511_,
		_w3561_,
		_w5209_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4747 (
		_w3563_,
		_w4629_,
		_w4632_,
		_w4635_,
		_w5210_
	);
	LUT2 #(
		.INIT('he)
	) name4748 (
		_w5209_,
		_w5210_,
		_w5211_
	);
	LUT3 #(
		.INIT('h2a)
	) name4749 (
		\P1_reg0_reg[5]/NET0131 ,
		_w3511_,
		_w3561_,
		_w5212_
	);
	LUT3 #(
		.INIT('hf2)
	) name4750 (
		_w3563_,
		_w4671_,
		_w5212_,
		_w5213_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4751 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[10]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w5214_
	);
	LUT2 #(
		.INIT('h8)
	) name4752 (
		\P1_reg1_reg[10]/NET0131 ,
		_w2183_,
		_w5215_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4753 (
		\P1_reg1_reg[10]/NET0131 ,
		_w2536_,
		_w4025_,
		_w4026_,
		_w5216_
	);
	LUT2 #(
		.INIT('h2)
	) name4754 (
		_w1237_,
		_w5216_,
		_w5217_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4755 (
		\P1_reg1_reg[10]/NET0131 ,
		_w1178_,
		_w2536_,
		_w2653_,
		_w5218_
	);
	LUT2 #(
		.INIT('h2)
	) name4756 (
		_w2128_,
		_w5218_,
		_w5219_
	);
	LUT4 #(
		.INIT('hc535)
	) name4757 (
		\P1_reg1_reg[10]/NET0131 ,
		_w1178_,
		_w2536_,
		_w2682_,
		_w5220_
	);
	LUT3 #(
		.INIT('ha2)
	) name4758 (
		\P1_reg1_reg[10]/NET0131 ,
		_w2332_,
		_w3975_,
		_w5221_
	);
	LUT4 #(
		.INIT('h0057)
	) name4759 (
		_w2536_,
		_w4032_,
		_w4034_,
		_w5221_,
		_w5222_
	);
	LUT3 #(
		.INIT('hd0)
	) name4760 (
		_w2121_,
		_w5220_,
		_w5222_,
		_w5223_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4761 (
		_w2182_,
		_w5217_,
		_w5219_,
		_w5223_,
		_w5224_
	);
	LUT4 #(
		.INIT('heeec)
	) name4762 (
		\P1_state_reg[0]/NET0131 ,
		_w5214_,
		_w5215_,
		_w5224_,
		_w5225_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4763 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg1_reg[11]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w5226_
	);
	LUT2 #(
		.INIT('h8)
	) name4764 (
		\P1_reg1_reg[11]/NET0131 ,
		_w2183_,
		_w5227_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4765 (
		\P1_reg1_reg[11]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w5228_
	);
	LUT4 #(
		.INIT('h7020)
	) name4766 (
		_w488_,
		_w889_,
		_w2536_,
		_w4004_,
		_w5229_
	);
	LUT3 #(
		.INIT('ha8)
	) name4767 (
		_w1237_,
		_w5228_,
		_w5229_,
		_w5230_
	);
	LUT4 #(
		.INIT('h8488)
	) name4768 (
		_w1174_,
		_w2536_,
		_w2962_,
		_w2963_,
		_w5231_
	);
	LUT3 #(
		.INIT('ha8)
	) name4769 (
		_w2121_,
		_w5228_,
		_w5231_,
		_w5232_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4770 (
		\P1_reg1_reg[11]/NET0131 ,
		_w2332_,
		_w3605_,
		_w3975_,
		_w5233_
	);
	LUT3 #(
		.INIT('h0d)
	) name4771 (
		_w2536_,
		_w4013_,
		_w5233_,
		_w5234_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4772 (
		_w2182_,
		_w5230_,
		_w5232_,
		_w5234_,
		_w5235_
	);
	LUT4 #(
		.INIT('heeec)
	) name4773 (
		\P1_state_reg[0]/NET0131 ,
		_w5226_,
		_w5227_,
		_w5235_,
		_w5236_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4774 (
		\P1_reg1_reg[13]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w5237_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4775 (
		_w3608_,
		_w4568_,
		_w4569_,
		_w5237_,
		_w5238_
	);
	LUT2 #(
		.INIT('h2)
	) name4776 (
		_w1237_,
		_w5238_,
		_w5239_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4777 (
		\P1_reg1_reg[13]/NET0131 ,
		_w2821_,
		_w3605_,
		_w4524_,
		_w5240_
	);
	LUT3 #(
		.INIT('h0d)
	) name4778 (
		_w3608_,
		_w4723_,
		_w5240_,
		_w5241_
	);
	LUT2 #(
		.INIT('hb)
	) name4779 (
		_w5239_,
		_w5241_,
		_w5242_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4780 (
		\P1_reg1_reg[14]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w5243_
	);
	LUT4 #(
		.INIT('h7020)
	) name4781 (
		_w488_,
		_w847_,
		_w3608_,
		_w4045_,
		_w5244_
	);
	LUT3 #(
		.INIT('ha8)
	) name4782 (
		_w1237_,
		_w5243_,
		_w5244_,
		_w5245_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4783 (
		_w3608_,
		_w4052_,
		_w4054_,
		_w4728_,
		_w5246_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4784 (
		\P1_reg1_reg[14]/NET0131 ,
		_w2821_,
		_w3605_,
		_w4524_,
		_w5247_
	);
	LUT3 #(
		.INIT('hfe)
	) name4785 (
		_w5246_,
		_w5245_,
		_w5247_,
		_w5248_
	);
	LUT3 #(
		.INIT('h2a)
	) name4786 (
		\P2_reg0_reg[11]/NET0131 ,
		_w2735_,
		_w4302_,
		_w5249_
	);
	LUT4 #(
		.INIT('hff8a)
	) name4787 (
		_w3153_,
		_w5130_,
		_w5135_,
		_w5249_,
		_w5250_
	);
	LUT2 #(
		.INIT('h1)
	) name4788 (
		\P2_reg3_reg[3]/NET0131 ,
		_w2903_,
		_w5251_
	);
	LUT4 #(
		.INIT('h4144)
	) name4789 (
		_w1305_,
		_w1670_,
		_w1675_,
		_w1969_,
		_w5252_
	);
	LUT3 #(
		.INIT('h80)
	) name4790 (
		_w1305_,
		_w1636_,
		_w1637_,
		_w5253_
	);
	LUT4 #(
		.INIT('heee2)
	) name4791 (
		\P2_reg3_reg[3]/NET0131 ,
		_w2903_,
		_w5252_,
		_w5253_,
		_w5254_
	);
	LUT4 #(
		.INIT('he100)
	) name4792 (
		_w1644_,
		_w1662_,
		_w2486_,
		_w2903_,
		_w5255_
	);
	LUT3 #(
		.INIT('ha8)
	) name4793 (
		_w1869_,
		_w5251_,
		_w5255_,
		_w5256_
	);
	LUT4 #(
		.INIT('he100)
	) name4794 (
		_w1884_,
		_w1887_,
		_w2486_,
		_w2903_,
		_w5257_
	);
	LUT4 #(
		.INIT('h7f80)
	) name4795 (
		_w1643_,
		_w1653_,
		_w1660_,
		_w1681_,
		_w5258_
	);
	LUT3 #(
		.INIT('h80)
	) name4796 (
		_w2025_,
		_w2903_,
		_w5258_,
		_w5259_
	);
	LUT4 #(
		.INIT('h4454)
	) name4797 (
		\P2_reg3_reg[3]/NET0131 ,
		_w2032_,
		_w2033_,
		_w2903_,
		_w5260_
	);
	LUT4 #(
		.INIT('h5450)
	) name4798 (
		_w1681_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w5261_
	);
	LUT3 #(
		.INIT('h01)
	) name4799 (
		_w5260_,
		_w5259_,
		_w5261_,
		_w5262_
	);
	LUT4 #(
		.INIT('h5700)
	) name4800 (
		_w1963_,
		_w5251_,
		_w5257_,
		_w5262_,
		_w5263_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4801 (
		_w2000_,
		_w5254_,
		_w5256_,
		_w5263_,
		_w5264_
	);
	LUT4 #(
		.INIT('h1000)
	) name4802 (
		\P2_reg3_reg[3]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5265_
	);
	LUT4 #(
		.INIT('haa08)
	) name4803 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w5264_,
		_w5265_,
		_w5266_
	);
	LUT2 #(
		.INIT('h4)
	) name4804 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[3]/NET0131 ,
		_w5267_
	);
	LUT3 #(
		.INIT('h9b)
	) name4805 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[3]/NET0131 ,
		_w1267_,
		_w5268_
	);
	LUT2 #(
		.INIT('hb)
	) name4806 (
		_w5266_,
		_w5268_,
		_w5269_
	);
	LUT2 #(
		.INIT('h2)
	) name4807 (
		_w1710_,
		_w2903_,
		_w5270_
	);
	LUT3 #(
		.INIT('h2a)
	) name4808 (
		_w1305_,
		_w1720_,
		_w1721_,
		_w5271_
	);
	LUT3 #(
		.INIT('h8a)
	) name4809 (
		_w1700_,
		_w1712_,
		_w4986_,
		_w5272_
	);
	LUT2 #(
		.INIT('h1)
	) name4810 (
		_w1305_,
		_w1972_,
		_w5273_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4811 (
		_w2903_,
		_w5271_,
		_w5272_,
		_w5273_,
		_w5274_
	);
	LUT3 #(
		.INIT('ha8)
	) name4812 (
		_w2000_,
		_w5270_,
		_w5274_,
		_w5275_
	);
	LUT4 #(
		.INIT('h4448)
	) name4813 (
		_w2485_,
		_w2903_,
		_w3015_,
		_w3092_,
		_w5276_
	);
	LUT3 #(
		.INIT('ha8)
	) name4814 (
		_w1869_,
		_w5270_,
		_w5276_,
		_w5277_
	);
	LUT4 #(
		.INIT('hb400)
	) name4815 (
		_w2410_,
		_w2411_,
		_w2485_,
		_w2903_,
		_w5278_
	);
	LUT4 #(
		.INIT('h9000)
	) name4816 (
		_w1717_,
		_w2004_,
		_w2025_,
		_w2903_,
		_w5279_
	);
	LUT4 #(
		.INIT('h88a8)
	) name4817 (
		_w1710_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w5280_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name4818 (
		_w1717_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w5281_
	);
	LUT2 #(
		.INIT('h1)
	) name4819 (
		_w5280_,
		_w5281_,
		_w5282_
	);
	LUT2 #(
		.INIT('h4)
	) name4820 (
		_w5279_,
		_w5282_,
		_w5283_
	);
	LUT4 #(
		.INIT('h5700)
	) name4821 (
		_w1963_,
		_w5270_,
		_w5278_,
		_w5283_,
		_w5284_
	);
	LUT2 #(
		.INIT('h4)
	) name4822 (
		_w5277_,
		_w5284_,
		_w5285_
	);
	LUT4 #(
		.INIT('h4000)
	) name4823 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1710_,
		_w5286_
	);
	LUT4 #(
		.INIT('h0075)
	) name4824 (
		_w1285_,
		_w5275_,
		_w5285_,
		_w5286_,
		_w5287_
	);
	LUT2 #(
		.INIT('h4)
	) name4825 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[6]/NET0131 ,
		_w5288_
	);
	LUT3 #(
		.INIT('h07)
	) name4826 (
		_w1710_,
		_w2344_,
		_w5288_,
		_w5289_
	);
	LUT3 #(
		.INIT('h2f)
	) name4827 (
		\P1_state_reg[0]/NET0131 ,
		_w5287_,
		_w5289_,
		_w5290_
	);
	LUT2 #(
		.INIT('h2)
	) name4828 (
		\P2_reg2_reg[5]/NET0131 ,
		_w2042_,
		_w5291_
	);
	LUT4 #(
		.INIT('he020)
	) name4829 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1298_,
		_w2000_,
		_w5005_,
		_w5292_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4830 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1298_,
		_w1687_,
		_w2497_,
		_w5293_
	);
	LUT2 #(
		.INIT('h8)
	) name4831 (
		_w1726_,
		_w2001_,
		_w5294_
	);
	LUT2 #(
		.INIT('h1)
	) name4832 (
		_w5010_,
		_w5294_,
		_w5295_
	);
	LUT4 #(
		.INIT('h80aa)
	) name4833 (
		_w1298_,
		_w1963_,
		_w5008_,
		_w5295_,
		_w5296_
	);
	LUT4 #(
		.INIT('h0200)
	) name4834 (
		_w1719_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w5297_
	);
	LUT4 #(
		.INIT('h005d)
	) name4835 (
		\P2_reg2_reg[5]/NET0131 ,
		_w2640_,
		_w3918_,
		_w5297_,
		_w5298_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4836 (
		_w1869_,
		_w5293_,
		_w5296_,
		_w5298_,
		_w5299_
	);
	LUT4 #(
		.INIT('h2000)
	) name4837 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5300_
	);
	LUT4 #(
		.INIT('h0075)
	) name4838 (
		_w1285_,
		_w5292_,
		_w5299_,
		_w5300_,
		_w5301_
	);
	LUT3 #(
		.INIT('hce)
	) name4839 (
		\P1_state_reg[0]/NET0131 ,
		_w5291_,
		_w5301_,
		_w5302_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4840 (
		\P1_reg1_reg[7]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w5303_
	);
	LUT4 #(
		.INIT('h7020)
	) name4841 (
		_w488_,
		_w927_,
		_w3608_,
		_w5058_,
		_w5304_
	);
	LUT3 #(
		.INIT('ha8)
	) name4842 (
		_w1237_,
		_w5303_,
		_w5304_,
		_w5305_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4843 (
		\P1_reg1_reg[7]/NET0131 ,
		_w2821_,
		_w3605_,
		_w4524_,
		_w5306_
	);
	LUT4 #(
		.INIT('h0075)
	) name4844 (
		_w3608_,
		_w5062_,
		_w5065_,
		_w5306_,
		_w5307_
	);
	LUT2 #(
		.INIT('hb)
	) name4845 (
		_w5305_,
		_w5307_,
		_w5308_
	);
	LUT2 #(
		.INIT('h2)
	) name4846 (
		\P2_reg0_reg[5]/NET0131 ,
		_w2042_,
		_w5309_
	);
	LUT4 #(
		.INIT('hc808)
	) name4847 (
		\P2_reg0_reg[5]/NET0131 ,
		_w2000_,
		_w2729_,
		_w5005_,
		_w5310_
	);
	LUT4 #(
		.INIT('hc355)
	) name4848 (
		\P2_reg0_reg[5]/NET0131 ,
		_w1687_,
		_w2497_,
		_w2729_,
		_w5311_
	);
	LUT3 #(
		.INIT('ha2)
	) name4849 (
		\P2_reg0_reg[5]/NET0131 ,
		_w3084_,
		_w3981_,
		_w5312_
	);
	LUT4 #(
		.INIT('h80cc)
	) name4850 (
		_w1963_,
		_w2729_,
		_w5008_,
		_w5295_,
		_w5313_
	);
	LUT4 #(
		.INIT('h0031)
	) name4851 (
		_w1869_,
		_w5312_,
		_w5311_,
		_w5313_,
		_w5314_
	);
	LUT4 #(
		.INIT('h2000)
	) name4852 (
		\P2_reg0_reg[5]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5315_
	);
	LUT4 #(
		.INIT('h0075)
	) name4853 (
		_w1285_,
		_w5310_,
		_w5314_,
		_w5315_,
		_w5316_
	);
	LUT3 #(
		.INIT('hce)
	) name4854 (
		\P1_state_reg[0]/NET0131 ,
		_w5309_,
		_w5316_,
		_w5317_
	);
	LUT2 #(
		.INIT('h2)
	) name4855 (
		\P2_reg0_reg[7]/NET0131 ,
		_w2042_,
		_w5318_
	);
	LUT4 #(
		.INIT('h2000)
	) name4856 (
		\P2_reg0_reg[7]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5319_
	);
	LUT4 #(
		.INIT('hc808)
	) name4857 (
		\P2_reg0_reg[7]/NET0131 ,
		_w2000_,
		_w2729_,
		_w5023_,
		_w5320_
	);
	LUT4 #(
		.INIT('hc808)
	) name4858 (
		\P2_reg0_reg[7]/NET0131 ,
		_w1869_,
		_w2729_,
		_w5025_,
		_w5321_
	);
	LUT3 #(
		.INIT('ha2)
	) name4859 (
		\P2_reg0_reg[7]/NET0131 ,
		_w3084_,
		_w3981_,
		_w5322_
	);
	LUT4 #(
		.INIT('he010)
	) name4860 (
		_w1897_,
		_w1901_,
		_w1963_,
		_w2496_,
		_w5323_
	);
	LUT2 #(
		.INIT('h8)
	) name4861 (
		_w1706_,
		_w2001_,
		_w5324_
	);
	LUT4 #(
		.INIT('h006f)
	) name4862 (
		_w1706_,
		_w2005_,
		_w2025_,
		_w5324_,
		_w5325_
	);
	LUT4 #(
		.INIT('h1311)
	) name4863 (
		_w2729_,
		_w5322_,
		_w5323_,
		_w5325_,
		_w5326_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4864 (
		_w1285_,
		_w5321_,
		_w5320_,
		_w5326_,
		_w5327_
	);
	LUT4 #(
		.INIT('heeec)
	) name4865 (
		\P1_state_reg[0]/NET0131 ,
		_w5318_,
		_w5319_,
		_w5327_,
		_w5328_
	);
	LUT2 #(
		.INIT('h2)
	) name4866 (
		\P2_reg1_reg[14]/NET0131 ,
		_w2042_,
		_w5329_
	);
	LUT4 #(
		.INIT('h2000)
	) name4867 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5330_
	);
	LUT2 #(
		.INIT('h2)
	) name4868 (
		\P2_reg1_reg[14]/NET0131 ,
		_w2762_,
		_w5331_
	);
	LUT4 #(
		.INIT('ha208)
	) name4869 (
		_w2762_,
		_w3115_,
		_w3491_,
		_w4606_,
		_w5332_
	);
	LUT3 #(
		.INIT('ha8)
	) name4870 (
		_w1963_,
		_w5331_,
		_w5332_,
		_w5333_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4871 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1869_,
		_w2762_,
		_w4612_,
		_w5334_
	);
	LUT4 #(
		.INIT('hc808)
	) name4872 (
		\P2_reg1_reg[14]/NET0131 ,
		_w2000_,
		_w2762_,
		_w4610_,
		_w5335_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4873 (
		\P2_reg1_reg[14]/NET0131 ,
		_w2033_,
		_w2734_,
		_w2762_,
		_w5336_
	);
	LUT4 #(
		.INIT('h0057)
	) name4874 (
		_w2762_,
		_w4614_,
		_w5182_,
		_w5336_,
		_w5337_
	);
	LUT3 #(
		.INIT('h10)
	) name4875 (
		_w5335_,
		_w5334_,
		_w5337_,
		_w5338_
	);
	LUT4 #(
		.INIT('h1311)
	) name4876 (
		_w1285_,
		_w5330_,
		_w5333_,
		_w5338_,
		_w5339_
	);
	LUT3 #(
		.INIT('hce)
	) name4877 (
		\P1_state_reg[0]/NET0131 ,
		_w5329_,
		_w5339_,
		_w5340_
	);
	LUT2 #(
		.INIT('h2)
	) name4878 (
		\P2_reg1_reg[5]/NET0131 ,
		_w2042_,
		_w5341_
	);
	LUT4 #(
		.INIT('hc808)
	) name4879 (
		\P2_reg1_reg[5]/NET0131 ,
		_w2000_,
		_w2762_,
		_w5005_,
		_w5342_
	);
	LUT4 #(
		.INIT('hc355)
	) name4880 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1687_,
		_w2497_,
		_w2762_,
		_w5343_
	);
	LUT2 #(
		.INIT('h2)
	) name4881 (
		\P2_reg1_reg[5]/NET0131 ,
		_w3872_,
		_w5344_
	);
	LUT4 #(
		.INIT('h80cc)
	) name4882 (
		_w1963_,
		_w2762_,
		_w5008_,
		_w5295_,
		_w5345_
	);
	LUT4 #(
		.INIT('h0031)
	) name4883 (
		_w1869_,
		_w5344_,
		_w5343_,
		_w5345_,
		_w5346_
	);
	LUT4 #(
		.INIT('h2000)
	) name4884 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5347_
	);
	LUT4 #(
		.INIT('h0075)
	) name4885 (
		_w1285_,
		_w5342_,
		_w5346_,
		_w5347_,
		_w5348_
	);
	LUT3 #(
		.INIT('hce)
	) name4886 (
		\P1_state_reg[0]/NET0131 ,
		_w5341_,
		_w5348_,
		_w5349_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name4887 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w5350_
	);
	LUT2 #(
		.INIT('h8)
	) name4888 (
		\P1_reg2_reg[3]/NET0131 ,
		_w2183_,
		_w5351_
	);
	LUT2 #(
		.INIT('h4)
	) name4889 (
		_w976_,
		_w2194_,
		_w5352_
	);
	LUT3 #(
		.INIT('h02)
	) name4890 (
		_w1237_,
		_w4966_,
		_w4967_,
		_w5353_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4891 (
		_w2189_,
		_w4976_,
		_w5352_,
		_w5353_,
		_w5354_
	);
	LUT4 #(
		.INIT('h0100)
	) name4892 (
		\P1_reg3_reg[3]/NET0131 ,
		_w1096_,
		_w1098_,
		_w1101_,
		_w5355_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4893 (
		_w1237_,
		_w2047_,
		_w2048_,
		_w2052_,
		_w5356_
	);
	LUT4 #(
		.INIT('h0001)
	) name4894 (
		_w2171_,
		_w3173_,
		_w5093_,
		_w5356_,
		_w5357_
	);
	LUT3 #(
		.INIT('h31)
	) name4895 (
		\P1_reg2_reg[3]/NET0131 ,
		_w5355_,
		_w5357_,
		_w5358_
	);
	LUT4 #(
		.INIT('h1311)
	) name4896 (
		_w2182_,
		_w5351_,
		_w5354_,
		_w5358_,
		_w5359_
	);
	LUT3 #(
		.INIT('hce)
	) name4897 (
		\P1_state_reg[0]/NET0131 ,
		_w5350_,
		_w5359_,
		_w5360_
	);
	LUT2 #(
		.INIT('h2)
	) name4898 (
		\P2_reg1_reg[7]/NET0131 ,
		_w2042_,
		_w5361_
	);
	LUT4 #(
		.INIT('h2000)
	) name4899 (
		\P2_reg1_reg[7]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5362_
	);
	LUT4 #(
		.INIT('hc808)
	) name4900 (
		\P2_reg1_reg[7]/NET0131 ,
		_w2000_,
		_w2762_,
		_w5023_,
		_w5363_
	);
	LUT4 #(
		.INIT('hc808)
	) name4901 (
		\P2_reg1_reg[7]/NET0131 ,
		_w1869_,
		_w2762_,
		_w5025_,
		_w5364_
	);
	LUT2 #(
		.INIT('h2)
	) name4902 (
		\P2_reg1_reg[7]/NET0131 ,
		_w3872_,
		_w5365_
	);
	LUT4 #(
		.INIT('h0075)
	) name4903 (
		_w2762_,
		_w5323_,
		_w5325_,
		_w5365_,
		_w5366_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4904 (
		_w1285_,
		_w5364_,
		_w5363_,
		_w5366_,
		_w5367_
	);
	LUT4 #(
		.INIT('heeec)
	) name4905 (
		\P1_state_reg[0]/NET0131 ,
		_w5361_,
		_w5362_,
		_w5367_,
		_w5368_
	);
	LUT4 #(
		.INIT('h5545)
	) name4906 (
		\P1_reg2_reg[6]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w5369_
	);
	LUT4 #(
		.INIT('h222a)
	) name4907 (
		_w1237_,
		_w2189_,
		_w5039_,
		_w5040_,
		_w5370_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4908 (
		_w2189_,
		_w5045_,
		_w5044_,
		_w5048_,
		_w5371_
	);
	LUT4 #(
		.INIT('h3331)
	) name4909 (
		_w3511_,
		_w5369_,
		_w5370_,
		_w5371_,
		_w5372_
	);
	LUT4 #(
		.INIT('h1000)
	) name4910 (
		_w1096_,
		_w1098_,
		_w925_,
		_w1101_,
		_w5373_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4911 (
		\P1_reg2_reg[6]/NET0131 ,
		_w2171_,
		_w3173_,
		_w5093_,
		_w5374_
	);
	LUT2 #(
		.INIT('h1)
	) name4912 (
		_w5373_,
		_w5374_,
		_w5375_
	);
	LUT2 #(
		.INIT('h1)
	) name4913 (
		\P1_reg2_reg[6]/NET0131 ,
		_w3511_,
		_w5376_
	);
	LUT3 #(
		.INIT('h0b)
	) name4914 (
		_w5372_,
		_w5375_,
		_w5376_,
		_w5377_
	);
	LUT4 #(
		.INIT('h1000)
	) name4915 (
		_w1096_,
		_w1098_,
		_w936_,
		_w1101_,
		_w5378_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4916 (
		_w2189_,
		_w5059_,
		_w5062_,
		_w5065_,
		_w5379_
	);
	LUT3 #(
		.INIT('h2a)
	) name4917 (
		\P1_reg2_reg[7]/NET0131 ,
		_w3175_,
		_w3512_,
		_w5380_
	);
	LUT4 #(
		.INIT('hffa8)
	) name4918 (
		_w3511_,
		_w5378_,
		_w5379_,
		_w5380_,
		_w5381_
	);
	LUT2 #(
		.INIT('h2)
	) name4919 (
		\P2_reg2_reg[4]/NET0131 ,
		_w2042_,
		_w5382_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4920 (
		_w1298_,
		_w4993_,
		_w4995_,
		_w5079_,
		_w5383_
	);
	LUT4 #(
		.INIT('h2e00)
	) name4921 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1298_,
		_w1666_,
		_w2001_,
		_w5384_
	);
	LUT4 #(
		.INIT('h0200)
	) name4922 (
		_w1668_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w5385_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name4923 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1298_,
		_w2032_,
		_w3154_,
		_w5386_
	);
	LUT3 #(
		.INIT('h01)
	) name4924 (
		_w5385_,
		_w5386_,
		_w5384_,
		_w5387_
	);
	LUT4 #(
		.INIT('h2000)
	) name4925 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5388_
	);
	LUT4 #(
		.INIT('h0075)
	) name4926 (
		_w1285_,
		_w5383_,
		_w5387_,
		_w5388_,
		_w5389_
	);
	LUT3 #(
		.INIT('hce)
	) name4927 (
		\P1_state_reg[0]/NET0131 ,
		_w5382_,
		_w5389_,
		_w5390_
	);
	LUT2 #(
		.INIT('h2)
	) name4928 (
		\P2_reg2_reg[7]/NET0131 ,
		_w2042_,
		_w5391_
	);
	LUT4 #(
		.INIT('h2000)
	) name4929 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5392_
	);
	LUT2 #(
		.INIT('h2)
	) name4930 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1298_,
		_w5393_
	);
	LUT4 #(
		.INIT('he020)
	) name4931 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1298_,
		_w2000_,
		_w5023_,
		_w5394_
	);
	LUT4 #(
		.INIT('he020)
	) name4932 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1298_,
		_w1869_,
		_w5025_,
		_w5395_
	);
	LUT4 #(
		.INIT('ha802)
	) name4933 (
		_w1298_,
		_w1897_,
		_w1901_,
		_w2496_,
		_w5396_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4934 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1298_,
		_w1706_,
		_w2005_,
		_w5397_
	);
	LUT4 #(
		.INIT('he200)
	) name4935 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1298_,
		_w1706_,
		_w2001_,
		_w5398_
	);
	LUT4 #(
		.INIT('h0200)
	) name4936 (
		_w1698_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w5399_
	);
	LUT4 #(
		.INIT('h0080)
	) name4937 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1863_,
		_w1866_,
		_w1999_,
		_w5400_
	);
	LUT2 #(
		.INIT('h1)
	) name4938 (
		_w5399_,
		_w5400_,
		_w5401_
	);
	LUT2 #(
		.INIT('h4)
	) name4939 (
		_w5398_,
		_w5401_,
		_w5402_
	);
	LUT3 #(
		.INIT('hd0)
	) name4940 (
		_w2025_,
		_w5397_,
		_w5402_,
		_w5403_
	);
	LUT4 #(
		.INIT('h5700)
	) name4941 (
		_w1963_,
		_w5393_,
		_w5396_,
		_w5403_,
		_w5404_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4942 (
		_w1285_,
		_w5395_,
		_w5394_,
		_w5404_,
		_w5405_
	);
	LUT4 #(
		.INIT('heeec)
	) name4943 (
		\P1_state_reg[0]/NET0131 ,
		_w5391_,
		_w5392_,
		_w5405_,
		_w5406_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4944 (
		_w3563_,
		_w4976_,
		_w5352_,
		_w5353_,
		_w5407_
	);
	LUT3 #(
		.INIT('h2a)
	) name4945 (
		\P1_reg0_reg[3]/NET0131 ,
		_w2332_,
		_w3563_,
		_w5408_
	);
	LUT2 #(
		.INIT('he)
	) name4946 (
		_w5407_,
		_w5408_,
		_w5409_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4947 (
		_w3563_,
		_w5059_,
		_w5062_,
		_w5065_,
		_w5410_
	);
	LUT3 #(
		.INIT('h2a)
	) name4948 (
		\P1_reg0_reg[7]/NET0131 ,
		_w3511_,
		_w3561_,
		_w5411_
	);
	LUT2 #(
		.INIT('he)
	) name4949 (
		_w5410_,
		_w5411_,
		_w5412_
	);
	LUT2 #(
		.INIT('h2)
	) name4950 (
		\P2_reg0_reg[14]/NET0131 ,
		_w2042_,
		_w5413_
	);
	LUT4 #(
		.INIT('h2000)
	) name4951 (
		\P2_reg0_reg[14]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5414_
	);
	LUT2 #(
		.INIT('h2)
	) name4952 (
		\P2_reg0_reg[14]/NET0131 ,
		_w2729_,
		_w5415_
	);
	LUT4 #(
		.INIT('ha208)
	) name4953 (
		_w2729_,
		_w3115_,
		_w3491_,
		_w4606_,
		_w5416_
	);
	LUT3 #(
		.INIT('ha8)
	) name4954 (
		_w1963_,
		_w5415_,
		_w5416_,
		_w5417_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4955 (
		\P2_reg0_reg[14]/NET0131 ,
		_w1869_,
		_w2729_,
		_w4612_,
		_w5418_
	);
	LUT4 #(
		.INIT('hc808)
	) name4956 (
		\P2_reg0_reg[14]/NET0131 ,
		_w2000_,
		_w2729_,
		_w4610_,
		_w5419_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4957 (
		\P2_reg0_reg[14]/NET0131 ,
		_w2033_,
		_w2729_,
		_w2734_,
		_w5420_
	);
	LUT4 #(
		.INIT('h0057)
	) name4958 (
		_w2729_,
		_w4614_,
		_w5182_,
		_w5420_,
		_w5421_
	);
	LUT3 #(
		.INIT('h10)
	) name4959 (
		_w5419_,
		_w5418_,
		_w5421_,
		_w5422_
	);
	LUT4 #(
		.INIT('h1311)
	) name4960 (
		_w1285_,
		_w5414_,
		_w5417_,
		_w5422_,
		_w5423_
	);
	LUT3 #(
		.INIT('hce)
	) name4961 (
		\P1_state_reg[0]/NET0131 ,
		_w5413_,
		_w5423_,
		_w5424_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4962 (
		\P1_reg1_reg[3]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w5425_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4963 (
		_w3608_,
		_w4966_,
		_w4967_,
		_w5425_,
		_w5426_
	);
	LUT2 #(
		.INIT('h2)
	) name4964 (
		_w1237_,
		_w5426_,
		_w5427_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4965 (
		\P1_reg1_reg[3]/NET0131 ,
		_w2821_,
		_w3605_,
		_w4524_,
		_w5428_
	);
	LUT4 #(
		.INIT('h005d)
	) name4966 (
		_w3608_,
		_w4976_,
		_w5352_,
		_w5428_,
		_w5429_
	);
	LUT2 #(
		.INIT('hb)
	) name4967 (
		_w5427_,
		_w5429_,
		_w5430_
	);
	LUT3 #(
		.INIT('h80)
	) name4968 (
		_w488_,
		_w987_,
		_w988_,
		_w5431_
	);
	LUT4 #(
		.INIT('h00eb)
	) name4969 (
		_w488_,
		_w971_,
		_w2130_,
		_w5431_,
		_w5432_
	);
	LUT4 #(
		.INIT('h4d00)
	) name4970 (
		_w989_,
		_w993_,
		_w1002_,
		_w1193_,
		_w5433_
	);
	LUT4 #(
		.INIT('h00b2)
	) name4971 (
		_w989_,
		_w993_,
		_w1002_,
		_w1193_,
		_w5434_
	);
	LUT3 #(
		.INIT('h02)
	) name4972 (
		_w2128_,
		_w5434_,
		_w5433_,
		_w5435_
	);
	LUT2 #(
		.INIT('h4)
	) name4973 (
		_w984_,
		_w2194_,
		_w5436_
	);
	LUT4 #(
		.INIT('h6a00)
	) name4974 (
		_w984_,
		_w993_,
		_w1001_,
		_w2170_,
		_w5437_
	);
	LUT2 #(
		.INIT('h1)
	) name4975 (
		_w5436_,
		_w5437_,
		_w5438_
	);
	LUT4 #(
		.INIT('h9f00)
	) name4976 (
		_w1193_,
		_w2069_,
		_w2121_,
		_w5438_,
		_w5439_
	);
	LUT4 #(
		.INIT('h0700)
	) name4977 (
		_w1237_,
		_w5432_,
		_w5435_,
		_w5439_,
		_w5440_
	);
	LUT2 #(
		.INIT('h4)
	) name4978 (
		_w984_,
		_w1120_,
		_w5441_
	);
	LUT4 #(
		.INIT('hcc08)
	) name4979 (
		_w2055_,
		_w3511_,
		_w5440_,
		_w5441_,
		_w5442_
	);
	LUT4 #(
		.INIT('h0010)
	) name4980 (
		_w2171_,
		_w2173_,
		_w3511_,
		_w4056_,
		_w5443_
	);
	LUT4 #(
		.INIT('h5d00)
	) name4981 (
		_w1237_,
		_w2055_,
		_w5432_,
		_w5443_,
		_w5444_
	);
	LUT2 #(
		.INIT('h2)
	) name4982 (
		\P1_reg3_reg[2]/NET0131 ,
		_w5444_,
		_w5445_
	);
	LUT2 #(
		.INIT('he)
	) name4983 (
		_w5442_,
		_w5445_,
		_w5446_
	);
	LUT3 #(
		.INIT('he6)
	) name4984 (
		_w1096_,
		_w1098_,
		_w1122_,
		_w5447_
	);
	LUT4 #(
		.INIT('hef00)
	) name4985 (
		_w2047_,
		_w2048_,
		_w2052_,
		_w5447_,
		_w5448_
	);
	LUT4 #(
		.INIT('h0008)
	) name4986 (
		_w2332_,
		_w3511_,
		_w3975_,
		_w5448_,
		_w5449_
	);
	LUT2 #(
		.INIT('h2)
	) name4987 (
		\P1_reg1_reg[6]/NET0131 ,
		_w5449_,
		_w5450_
	);
	LUT4 #(
		.INIT('hff8a)
	) name4988 (
		_w3608_,
		_w5043_,
		_w5049_,
		_w5450_,
		_w5451_
	);
	LUT2 #(
		.INIT('h2)
	) name4989 (
		\P2_reg0_reg[3]/NET0131 ,
		_w2729_,
		_w5452_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4990 (
		\P2_reg0_reg[3]/NET0131 ,
		_w2729_,
		_w5252_,
		_w5253_,
		_w5453_
	);
	LUT4 #(
		.INIT('he100)
	) name4991 (
		_w1644_,
		_w1662_,
		_w2486_,
		_w2729_,
		_w5454_
	);
	LUT3 #(
		.INIT('ha8)
	) name4992 (
		_w1869_,
		_w5452_,
		_w5454_,
		_w5455_
	);
	LUT3 #(
		.INIT('ha2)
	) name4993 (
		\P2_reg0_reg[3]/NET0131 ,
		_w3084_,
		_w3981_,
		_w5456_
	);
	LUT4 #(
		.INIT('he010)
	) name4994 (
		_w1884_,
		_w1887_,
		_w1963_,
		_w2486_,
		_w5457_
	);
	LUT2 #(
		.INIT('h4)
	) name4995 (
		_w1681_,
		_w2001_,
		_w5458_
	);
	LUT3 #(
		.INIT('h07)
	) name4996 (
		_w2025_,
		_w5258_,
		_w5458_,
		_w5459_
	);
	LUT4 #(
		.INIT('h1311)
	) name4997 (
		_w2729_,
		_w5456_,
		_w5457_,
		_w5459_,
		_w5460_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4998 (
		_w2000_,
		_w5453_,
		_w5455_,
		_w5460_,
		_w5461_
	);
	LUT4 #(
		.INIT('h2000)
	) name4999 (
		\P2_reg0_reg[3]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5462_
	);
	LUT4 #(
		.INIT('haa08)
	) name5000 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w5461_,
		_w5462_,
		_w5463_
	);
	LUT2 #(
		.INIT('h2)
	) name5001 (
		\P2_reg0_reg[3]/NET0131 ,
		_w2042_,
		_w5464_
	);
	LUT2 #(
		.INIT('he)
	) name5002 (
		_w5463_,
		_w5464_,
		_w5465_
	);
	LUT2 #(
		.INIT('h2)
	) name5003 (
		\P2_reg1_reg[3]/NET0131 ,
		_w2042_,
		_w5466_
	);
	LUT2 #(
		.INIT('h2)
	) name5004 (
		\P2_reg1_reg[3]/NET0131 ,
		_w2762_,
		_w5467_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5005 (
		\P2_reg1_reg[3]/NET0131 ,
		_w2762_,
		_w5252_,
		_w5253_,
		_w5468_
	);
	LUT4 #(
		.INIT('he100)
	) name5006 (
		_w1644_,
		_w1662_,
		_w2486_,
		_w2762_,
		_w5469_
	);
	LUT3 #(
		.INIT('ha8)
	) name5007 (
		_w1869_,
		_w5467_,
		_w5469_,
		_w5470_
	);
	LUT2 #(
		.INIT('h2)
	) name5008 (
		\P2_reg1_reg[3]/NET0131 ,
		_w3872_,
		_w5471_
	);
	LUT4 #(
		.INIT('h0075)
	) name5009 (
		_w2762_,
		_w5457_,
		_w5459_,
		_w5471_,
		_w5472_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5010 (
		_w2000_,
		_w5468_,
		_w5470_,
		_w5472_,
		_w5473_
	);
	LUT4 #(
		.INIT('h2000)
	) name5011 (
		\P2_reg1_reg[3]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5474_
	);
	LUT4 #(
		.INIT('haa08)
	) name5012 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w5473_,
		_w5474_,
		_w5475_
	);
	LUT2 #(
		.INIT('he)
	) name5013 (
		_w5466_,
		_w5475_,
		_w5476_
	);
	LUT2 #(
		.INIT('h2)
	) name5014 (
		\P2_reg2_reg[3]/NET0131 ,
		_w1298_,
		_w5477_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5015 (
		\P2_reg2_reg[3]/NET0131 ,
		_w1298_,
		_w5252_,
		_w5253_,
		_w5478_
	);
	LUT4 #(
		.INIT('ha802)
	) name5016 (
		_w1298_,
		_w1644_,
		_w1662_,
		_w2486_,
		_w5479_
	);
	LUT3 #(
		.INIT('ha8)
	) name5017 (
		_w1869_,
		_w5477_,
		_w5479_,
		_w5480_
	);
	LUT4 #(
		.INIT('ha802)
	) name5018 (
		_w1298_,
		_w1884_,
		_w1887_,
		_w2486_,
		_w5481_
	);
	LUT4 #(
		.INIT('he020)
	) name5019 (
		\P2_reg2_reg[3]/NET0131 ,
		_w1298_,
		_w2025_,
		_w5258_,
		_w5482_
	);
	LUT4 #(
		.INIT('h2e00)
	) name5020 (
		\P2_reg2_reg[3]/NET0131 ,
		_w1298_,
		_w1681_,
		_w2001_,
		_w5483_
	);
	LUT4 #(
		.INIT('h0100)
	) name5021 (
		\P2_reg3_reg[3]/NET0131 ,
		_w1863_,
		_w1866_,
		_w2028_,
		_w5484_
	);
	LUT4 #(
		.INIT('h0080)
	) name5022 (
		\P2_reg2_reg[3]/NET0131 ,
		_w1863_,
		_w1866_,
		_w1999_,
		_w5485_
	);
	LUT2 #(
		.INIT('h1)
	) name5023 (
		_w5484_,
		_w5485_,
		_w5486_
	);
	LUT3 #(
		.INIT('h10)
	) name5024 (
		_w5482_,
		_w5483_,
		_w5486_,
		_w5487_
	);
	LUT4 #(
		.INIT('h5700)
	) name5025 (
		_w1963_,
		_w5477_,
		_w5481_,
		_w5487_,
		_w5488_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5026 (
		_w2000_,
		_w5478_,
		_w5480_,
		_w5488_,
		_w5489_
	);
	LUT4 #(
		.INIT('h2000)
	) name5027 (
		\P2_reg2_reg[3]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5490_
	);
	LUT4 #(
		.INIT('haa08)
	) name5028 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w5489_,
		_w5490_,
		_w5491_
	);
	LUT2 #(
		.INIT('h2)
	) name5029 (
		\P2_reg2_reg[3]/NET0131 ,
		_w2042_,
		_w5492_
	);
	LUT2 #(
		.INIT('he)
	) name5030 (
		_w5491_,
		_w5492_,
		_w5493_
	);
	LUT2 #(
		.INIT('h2)
	) name5031 (
		\P2_reg2_reg[6]/NET0131 ,
		_w2042_,
		_w5494_
	);
	LUT4 #(
		.INIT('h2000)
	) name5032 (
		\P2_reg2_reg[6]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5495_
	);
	LUT2 #(
		.INIT('h2)
	) name5033 (
		\P2_reg2_reg[6]/NET0131 ,
		_w1298_,
		_w5496_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5034 (
		_w1298_,
		_w5271_,
		_w5272_,
		_w5273_,
		_w5497_
	);
	LUT3 #(
		.INIT('ha8)
	) name5035 (
		_w2000_,
		_w5496_,
		_w5497_,
		_w5498_
	);
	LUT4 #(
		.INIT('h2228)
	) name5036 (
		_w1298_,
		_w2485_,
		_w3015_,
		_w3092_,
		_w5499_
	);
	LUT3 #(
		.INIT('ha8)
	) name5037 (
		_w1869_,
		_w5496_,
		_w5499_,
		_w5500_
	);
	LUT4 #(
		.INIT('h8a20)
	) name5038 (
		_w1963_,
		_w2410_,
		_w2411_,
		_w2485_,
		_w5501_
	);
	LUT2 #(
		.INIT('h8)
	) name5039 (
		_w1717_,
		_w2001_,
		_w5502_
	);
	LUT4 #(
		.INIT('h006f)
	) name5040 (
		_w1717_,
		_w2004_,
		_w2025_,
		_w5502_,
		_w5503_
	);
	LUT4 #(
		.INIT('h0200)
	) name5041 (
		_w1710_,
		_w1863_,
		_w1866_,
		_w2028_,
		_w5504_
	);
	LUT4 #(
		.INIT('h005d)
	) name5042 (
		\P2_reg2_reg[6]/NET0131 ,
		_w2640_,
		_w3918_,
		_w5504_,
		_w5505_
	);
	LUT4 #(
		.INIT('h7500)
	) name5043 (
		_w1298_,
		_w5501_,
		_w5503_,
		_w5505_,
		_w5506_
	);
	LUT2 #(
		.INIT('h4)
	) name5044 (
		_w5500_,
		_w5506_,
		_w5507_
	);
	LUT4 #(
		.INIT('h1311)
	) name5045 (
		_w1285_,
		_w5495_,
		_w5498_,
		_w5507_,
		_w5508_
	);
	LUT3 #(
		.INIT('hce)
	) name5046 (
		\P1_state_reg[0]/NET0131 ,
		_w5494_,
		_w5508_,
		_w5509_
	);
	LUT3 #(
		.INIT('h2a)
	) name5047 (
		\P1_reg0_reg[6]/NET0131 ,
		_w3511_,
		_w3561_,
		_w5510_
	);
	LUT4 #(
		.INIT('hff8a)
	) name5048 (
		_w3563_,
		_w5043_,
		_w5049_,
		_w5510_,
		_w5511_
	);
	LUT2 #(
		.INIT('h2)
	) name5049 (
		\P2_reg0_reg[6]/NET0131 ,
		_w2729_,
		_w5512_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5050 (
		_w2729_,
		_w5271_,
		_w5272_,
		_w5273_,
		_w5513_
	);
	LUT3 #(
		.INIT('ha8)
	) name5051 (
		_w2000_,
		_w5512_,
		_w5513_,
		_w5514_
	);
	LUT4 #(
		.INIT('h4448)
	) name5052 (
		_w2485_,
		_w2729_,
		_w3015_,
		_w3092_,
		_w5515_
	);
	LUT3 #(
		.INIT('ha8)
	) name5053 (
		_w1869_,
		_w5512_,
		_w5515_,
		_w5516_
	);
	LUT3 #(
		.INIT('ha2)
	) name5054 (
		\P2_reg0_reg[6]/NET0131 ,
		_w3084_,
		_w3981_,
		_w5517_
	);
	LUT4 #(
		.INIT('h0075)
	) name5055 (
		_w2729_,
		_w5501_,
		_w5503_,
		_w5517_,
		_w5518_
	);
	LUT2 #(
		.INIT('h4)
	) name5056 (
		_w5516_,
		_w5518_,
		_w5519_
	);
	LUT4 #(
		.INIT('h2000)
	) name5057 (
		\P2_reg0_reg[6]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5520_
	);
	LUT4 #(
		.INIT('h0075)
	) name5058 (
		_w1285_,
		_w5514_,
		_w5519_,
		_w5520_,
		_w5521_
	);
	LUT2 #(
		.INIT('h2)
	) name5059 (
		\P2_reg0_reg[6]/NET0131 ,
		_w2042_,
		_w5522_
	);
	LUT3 #(
		.INIT('hf2)
	) name5060 (
		\P1_state_reg[0]/NET0131 ,
		_w5521_,
		_w5522_,
		_w5523_
	);
	LUT4 #(
		.INIT('h5545)
	) name5061 (
		\P1_reg2_reg[2]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w5524_
	);
	LUT3 #(
		.INIT('ha2)
	) name5062 (
		_w1237_,
		_w2189_,
		_w5432_,
		_w5525_
	);
	LUT4 #(
		.INIT('h4c44)
	) name5063 (
		_w2189_,
		_w3511_,
		_w5435_,
		_w5439_,
		_w5526_
	);
	LUT4 #(
		.INIT('h0200)
	) name5064 (
		\P1_reg3_reg[2]/NET0131 ,
		_w1096_,
		_w1098_,
		_w1101_,
		_w5527_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5065 (
		\P1_reg2_reg[2]/NET0131 ,
		_w2171_,
		_w3173_,
		_w5093_,
		_w5528_
	);
	LUT2 #(
		.INIT('h1)
	) name5066 (
		_w5527_,
		_w5528_,
		_w5529_
	);
	LUT4 #(
		.INIT('hba00)
	) name5067 (
		_w5524_,
		_w5525_,
		_w5526_,
		_w5529_,
		_w5530_
	);
	LUT2 #(
		.INIT('h1)
	) name5068 (
		\P1_reg2_reg[2]/NET0131 ,
		_w3511_,
		_w5531_
	);
	LUT2 #(
		.INIT('h1)
	) name5069 (
		_w5530_,
		_w5531_,
		_w5532_
	);
	LUT2 #(
		.INIT('h2)
	) name5070 (
		\P2_reg1_reg[6]/NET0131 ,
		_w2762_,
		_w5533_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5071 (
		_w2762_,
		_w5271_,
		_w5272_,
		_w5273_,
		_w5534_
	);
	LUT3 #(
		.INIT('ha8)
	) name5072 (
		_w2000_,
		_w5533_,
		_w5534_,
		_w5535_
	);
	LUT4 #(
		.INIT('h4448)
	) name5073 (
		_w2485_,
		_w2762_,
		_w3015_,
		_w3092_,
		_w5536_
	);
	LUT3 #(
		.INIT('ha8)
	) name5074 (
		_w1869_,
		_w5533_,
		_w5536_,
		_w5537_
	);
	LUT2 #(
		.INIT('h2)
	) name5075 (
		\P2_reg1_reg[6]/NET0131 ,
		_w3872_,
		_w5538_
	);
	LUT4 #(
		.INIT('h0075)
	) name5076 (
		_w2762_,
		_w5501_,
		_w5503_,
		_w5538_,
		_w5539_
	);
	LUT2 #(
		.INIT('h4)
	) name5077 (
		_w5537_,
		_w5539_,
		_w5540_
	);
	LUT4 #(
		.INIT('h2000)
	) name5078 (
		\P2_reg1_reg[6]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5541_
	);
	LUT4 #(
		.INIT('h0075)
	) name5079 (
		_w1285_,
		_w5535_,
		_w5540_,
		_w5541_,
		_w5542_
	);
	LUT2 #(
		.INIT('h2)
	) name5080 (
		\P2_reg1_reg[6]/NET0131 ,
		_w2042_,
		_w5543_
	);
	LUT3 #(
		.INIT('hf2)
	) name5081 (
		\P1_state_reg[0]/NET0131 ,
		_w5542_,
		_w5543_,
		_w5544_
	);
	LUT3 #(
		.INIT('h2a)
	) name5082 (
		\P1_reg0_reg[2]/NET0131 ,
		_w3511_,
		_w3561_,
		_w5545_
	);
	LUT3 #(
		.INIT('hf2)
	) name5083 (
		_w3563_,
		_w5440_,
		_w5545_,
		_w5546_
	);
	LUT3 #(
		.INIT('h2a)
	) name5084 (
		\P1_reg1_reg[2]/NET0131 ,
		_w3511_,
		_w3976_,
		_w5547_
	);
	LUT3 #(
		.INIT('hf2)
	) name5085 (
		_w3608_,
		_w5440_,
		_w5547_,
		_w5548_
	);
	LUT3 #(
		.INIT('h10)
	) name5086 (
		_w993_,
		_w2175_,
		_w2176_,
		_w5549_
	);
	LUT4 #(
		.INIT('h5556)
	) name5087 (
		_w980_,
		_w989_,
		_w998_,
		_w602_,
		_w5550_
	);
	LUT4 #(
		.INIT('h7020)
	) name5088 (
		_w488_,
		_w998_,
		_w1237_,
		_w5550_,
		_w5551_
	);
	LUT3 #(
		.INIT('h90)
	) name5089 (
		_w1002_,
		_w1190_,
		_w2128_,
		_w5552_
	);
	LUT3 #(
		.INIT('h60)
	) name5090 (
		_w993_,
		_w1001_,
		_w2170_,
		_w5553_
	);
	LUT4 #(
		.INIT('h006f)
	) name5091 (
		_w1190_,
		_w2068_,
		_w2121_,
		_w5553_,
		_w5554_
	);
	LUT2 #(
		.INIT('h4)
	) name5092 (
		_w5552_,
		_w5554_,
		_w5555_
	);
	LUT4 #(
		.INIT('h1311)
	) name5093 (
		_w2055_,
		_w5549_,
		_w5551_,
		_w5555_,
		_w5556_
	);
	LUT2 #(
		.INIT('h2)
	) name5094 (
		_w3511_,
		_w3791_,
		_w5557_
	);
	LUT3 #(
		.INIT('h2a)
	) name5095 (
		\P1_reg3_reg[1]/NET0131 ,
		_w4057_,
		_w5557_,
		_w5558_
	);
	LUT3 #(
		.INIT('hf2)
	) name5096 (
		_w3511_,
		_w5556_,
		_w5558_,
		_w5559_
	);
	LUT2 #(
		.INIT('h1)
	) name5097 (
		\P2_reg3_reg[1]/NET0131 ,
		_w2903_,
		_w5560_
	);
	LUT4 #(
		.INIT('h5556)
	) name5098 (
		_w1638_,
		_w1648_,
		_w1656_,
		_w1967_,
		_w5561_
	);
	LUT4 #(
		.INIT('h80d0)
	) name5099 (
		_w1305_,
		_w1656_,
		_w2903_,
		_w5561_,
		_w5562_
	);
	LUT2 #(
		.INIT('h6)
	) name5100 (
		_w1653_,
		_w1660_,
		_w5563_
	);
	LUT3 #(
		.INIT('h60)
	) name5101 (
		_w1653_,
		_w1660_,
		_w2025_,
		_w5564_
	);
	LUT3 #(
		.INIT('h84)
	) name5102 (
		_w1882_,
		_w1963_,
		_w2500_,
		_w5565_
	);
	LUT3 #(
		.INIT('h84)
	) name5103 (
		_w1661_,
		_w1869_,
		_w2500_,
		_w5566_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5104 (
		_w2903_,
		_w5564_,
		_w5565_,
		_w5566_,
		_w5567_
	);
	LUT4 #(
		.INIT('h00c4)
	) name5105 (
		_w2000_,
		_w2556_,
		_w5562_,
		_w5567_,
		_w5568_
	);
	LUT4 #(
		.INIT('h5450)
	) name5106 (
		_w1653_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w5569_
	);
	LUT4 #(
		.INIT('haa02)
	) name5107 (
		_w2556_,
		_w5560_,
		_w5568_,
		_w5569_,
		_w5570_
	);
	LUT3 #(
		.INIT('h89)
	) name5108 (
		_w1863_,
		_w1866_,
		_w1999_,
		_w5571_
	);
	LUT4 #(
		.INIT('h3130)
	) name5109 (
		_w2001_,
		_w2032_,
		_w2903_,
		_w5571_,
		_w5572_
	);
	LUT4 #(
		.INIT('h0e00)
	) name5110 (
		_w5560_,
		_w5568_,
		_w5569_,
		_w5572_,
		_w5573_
	);
	LUT3 #(
		.INIT('h0e)
	) name5111 (
		\P2_reg3_reg[1]/NET0131 ,
		_w5570_,
		_w5573_,
		_w5574_
	);
	LUT2 #(
		.INIT('h1)
	) name5112 (
		\P2_reg3_reg[2]/NET0131 ,
		_w2903_,
		_w5575_
	);
	LUT3 #(
		.INIT('h80)
	) name5113 (
		_w1305_,
		_w1646_,
		_w1647_,
		_w5576_
	);
	LUT4 #(
		.INIT('h00eb)
	) name5114 (
		_w1305_,
		_w1675_,
		_w1969_,
		_w5576_,
		_w5577_
	);
	LUT3 #(
		.INIT('ha2)
	) name5115 (
		_w2000_,
		_w2903_,
		_w5577_,
		_w5578_
	);
	LUT4 #(
		.INIT('h0071)
	) name5116 (
		_w1648_,
		_w1653_,
		_w1661_,
		_w2487_,
		_w5579_
	);
	LUT4 #(
		.INIT('h8e00)
	) name5117 (
		_w1648_,
		_w1653_,
		_w1661_,
		_w2487_,
		_w5580_
	);
	LUT3 #(
		.INIT('h02)
	) name5118 (
		_w1869_,
		_w5580_,
		_w5579_,
		_w5581_
	);
	LUT4 #(
		.INIT('h6a00)
	) name5119 (
		_w1643_,
		_w1653_,
		_w1660_,
		_w2025_,
		_w5582_
	);
	LUT4 #(
		.INIT('h007d)
	) name5120 (
		_w1963_,
		_w2407_,
		_w2487_,
		_w5582_,
		_w5583_
	);
	LUT4 #(
		.INIT('h2a22)
	) name5121 (
		_w2556_,
		_w2903_,
		_w5581_,
		_w5583_,
		_w5584_
	);
	LUT4 #(
		.INIT('h5450)
	) name5122 (
		_w1643_,
		_w2001_,
		_w2029_,
		_w2903_,
		_w5585_
	);
	LUT4 #(
		.INIT('h00ba)
	) name5123 (
		_w5575_,
		_w5578_,
		_w5584_,
		_w5585_,
		_w5586_
	);
	LUT4 #(
		.INIT('h0aee)
	) name5124 (
		\P2_reg3_reg[2]/NET0131 ,
		_w2556_,
		_w5572_,
		_w5586_,
		_w5587_
	);
	LUT2 #(
		.INIT('h4)
	) name5125 (
		_w1643_,
		_w2001_,
		_w5588_
	);
	LUT3 #(
		.INIT('h04)
	) name5126 (
		_w5581_,
		_w5583_,
		_w5588_,
		_w5589_
	);
	LUT2 #(
		.INIT('h8)
	) name5127 (
		_w2000_,
		_w5577_,
		_w5590_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name5128 (
		\P2_reg0_reg[2]/NET0131 ,
		_w3082_,
		_w3083_,
		_w4302_,
		_w5591_
	);
	LUT4 #(
		.INIT('hffa2)
	) name5129 (
		_w3153_,
		_w5589_,
		_w5590_,
		_w5591_,
		_w5592_
	);
	LUT2 #(
		.INIT('h2)
	) name5130 (
		\P2_reg1_reg[2]/NET0131 ,
		_w2042_,
		_w5593_
	);
	LUT4 #(
		.INIT('h2000)
	) name5131 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5594_
	);
	LUT2 #(
		.INIT('h2)
	) name5132 (
		\P2_reg1_reg[2]/NET0131 ,
		_w3241_,
		_w5595_
	);
	LUT4 #(
		.INIT('h005d)
	) name5133 (
		_w2762_,
		_w5589_,
		_w5590_,
		_w5595_,
		_w5596_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5134 (
		\P1_state_reg[0]/NET0131 ,
		_w1285_,
		_w5594_,
		_w5596_,
		_w5597_
	);
	LUT2 #(
		.INIT('he)
	) name5135 (
		_w5593_,
		_w5597_,
		_w5598_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name5136 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_reg0_reg[1]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1242_,
		_w5599_
	);
	LUT2 #(
		.INIT('h8)
	) name5137 (
		\P1_reg0_reg[1]/NET0131 ,
		_w2183_,
		_w5600_
	);
	LUT2 #(
		.INIT('h4)
	) name5138 (
		_w993_,
		_w2194_,
		_w5601_
	);
	LUT3 #(
		.INIT('h04)
	) name5139 (
		_w5552_,
		_w5554_,
		_w5601_,
		_w5602_
	);
	LUT4 #(
		.INIT('haaa2)
	) name5140 (
		\P1_reg0_reg[1]/NET0131 ,
		_w2332_,
		_w2333_,
		_w3567_,
		_w5603_
	);
	LUT4 #(
		.INIT('h0075)
	) name5141 (
		_w2325_,
		_w5551_,
		_w5602_,
		_w5603_,
		_w5604_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5142 (
		\P1_state_reg[0]/NET0131 ,
		_w2182_,
		_w5600_,
		_w5604_,
		_w5605_
	);
	LUT2 #(
		.INIT('he)
	) name5143 (
		_w5599_,
		_w5605_,
		_w5606_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5144 (
		\P1_reg1_reg[1]/NET0131 ,
		_w2047_,
		_w2048_,
		_w2052_,
		_w5607_
	);
	LUT4 #(
		.INIT('h7020)
	) name5145 (
		_w488_,
		_w998_,
		_w3608_,
		_w5550_,
		_w5608_
	);
	LUT3 #(
		.INIT('ha8)
	) name5146 (
		_w1237_,
		_w5607_,
		_w5608_,
		_w5609_
	);
	LUT4 #(
		.INIT('haa8a)
	) name5147 (
		_w3608_,
		_w5552_,
		_w5554_,
		_w5601_,
		_w5610_
	);
	LUT3 #(
		.INIT('h8a)
	) name5148 (
		\P1_reg1_reg[1]/NET0131 ,
		_w3626_,
		_w4524_,
		_w5611_
	);
	LUT2 #(
		.INIT('h1)
	) name5149 (
		_w5610_,
		_w5611_,
		_w5612_
	);
	LUT2 #(
		.INIT('hb)
	) name5150 (
		_w5609_,
		_w5612_,
		_w5613_
	);
	LUT2 #(
		.INIT('h2)
	) name5151 (
		\P2_reg2_reg[1]/NET0131 ,
		_w2042_,
		_w5614_
	);
	LUT4 #(
		.INIT('h2000)
	) name5152 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w5615_
	);
	LUT2 #(
		.INIT('h2)
	) name5153 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1298_,
		_w5616_
	);
	LUT4 #(
		.INIT('h2a08)
	) name5154 (
		_w1298_,
		_w1305_,
		_w1656_,
		_w5561_,
		_w5617_
	);
	LUT3 #(
		.INIT('ha8)
	) name5155 (
		_w2000_,
		_w5616_,
		_w5617_,
		_w5618_
	);
	LUT2 #(
		.INIT('h4)
	) name5156 (
		_w1653_,
		_w2001_,
		_w5619_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5157 (
		_w1298_,
		_w5565_,
		_w5566_,
		_w5619_,
		_w5620_
	);
	LUT4 #(
		.INIT('he020)
	) name5158 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1298_,
		_w2025_,
		_w5563_,
		_w5621_
	);
	LUT4 #(
		.INIT('h0200)
	) name5159 (
		\P2_reg3_reg[1]/NET0131 ,
		_w1863_,
		_w1866_,
		_w2028_,
		_w5622_
	);
	LUT4 #(
		.INIT('h0075)
	) name5160 (
		\P2_reg2_reg[1]/NET0131 ,
		_w2639_,
		_w3919_,
		_w5622_,
		_w5623_
	);
	LUT3 #(
		.INIT('h10)
	) name5161 (
		_w5620_,
		_w5621_,
		_w5623_,
		_w5624_
	);
	LUT4 #(
		.INIT('h1311)
	) name5162 (
		_w1285_,
		_w5615_,
		_w5618_,
		_w5624_,
		_w5625_
	);
	LUT3 #(
		.INIT('hce)
	) name5163 (
		\P1_state_reg[0]/NET0131 ,
		_w5614_,
		_w5625_,
		_w5626_
	);
	LUT4 #(
		.INIT('h0200)
	) name5164 (
		\P1_reg3_reg[1]/NET0131 ,
		_w1096_,
		_w1098_,
		_w1101_,
		_w5627_
	);
	LUT4 #(
		.INIT('h0075)
	) name5165 (
		_w2189_,
		_w5551_,
		_w5602_,
		_w5627_,
		_w5628_
	);
	LUT4 #(
		.INIT('h1030)
	) name5166 (
		_w2119_,
		_w3174_,
		_w3511_,
		_w5093_,
		_w5629_
	);
	LUT3 #(
		.INIT('h2a)
	) name5167 (
		\P1_reg2_reg[1]/NET0131 ,
		_w3858_,
		_w5629_,
		_w5630_
	);
	LUT3 #(
		.INIT('hf2)
	) name5168 (
		_w3511_,
		_w5628_,
		_w5630_,
		_w5631_
	);
	LUT2 #(
		.INIT('h2)
	) name5169 (
		\P2_reg1_reg[1]/NET0131 ,
		_w2042_,
		_w5632_
	);
	LUT4 #(
		.INIT('h7020)
	) name5170 (
		_w1305_,
		_w1656_,
		_w2000_,
		_w5561_,
		_w5633_
	);
	LUT4 #(
		.INIT('h0001)
	) name5171 (
		_w5564_,
		_w5565_,
		_w5566_,
		_w5619_,
		_w5634_
	);
	LUT4 #(
		.INIT('h8884)
	) name5172 (
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[1]/NET0131 ,
		_w1264_,
		_w1266_,
		_w5635_
	);
	LUT3 #(
		.INIT('h70)
	) name5173 (
		_w3872_,
		_w3891_,
		_w5635_,
		_w5636_
	);
	LUT4 #(
		.INIT('h0075)
	) name5174 (
		_w3243_,
		_w5633_,
		_w5634_,
		_w5636_,
		_w5637_
	);
	LUT3 #(
		.INIT('hce)
	) name5175 (
		\P1_state_reg[0]/NET0131 ,
		_w5632_,
		_w5637_,
		_w5638_
	);
	LUT2 #(
		.INIT('h1)
	) name5176 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1298_,
		_w5639_
	);
	LUT3 #(
		.INIT('hc4)
	) name5177 (
		_w1298_,
		_w2000_,
		_w5577_,
		_w5640_
	);
	LUT4 #(
		.INIT('haa8a)
	) name5178 (
		_w1298_,
		_w5581_,
		_w5583_,
		_w5588_,
		_w5641_
	);
	LUT4 #(
		.INIT('h3331)
	) name5179 (
		_w2556_,
		_w5639_,
		_w5641_,
		_w5640_,
		_w5642_
	);
	LUT4 #(
		.INIT('h0200)
	) name5180 (
		\P2_reg3_reg[2]/NET0131 ,
		_w1863_,
		_w1866_,
		_w2028_,
		_w5643_
	);
	LUT4 #(
		.INIT('h1115)
	) name5181 (
		\P2_reg2_reg[2]/NET0131 ,
		_w2556_,
		_w5642_,
		_w5643_,
		_w5644_
	);
	LUT2 #(
		.INIT('h4)
	) name5182 (
		_w2035_,
		_w3919_,
		_w5645_
	);
	LUT3 #(
		.INIT('h10)
	) name5183 (
		_w5642_,
		_w5643_,
		_w5645_,
		_w5646_
	);
	LUT2 #(
		.INIT('h1)
	) name5184 (
		_w5644_,
		_w5646_,
		_w5647_
	);
	LUT2 #(
		.INIT('h2)
	) name5185 (
		\P2_reg0_reg[1]/NET0131 ,
		_w2729_,
		_w5648_
	);
	LUT4 #(
		.INIT('h7020)
	) name5186 (
		_w1305_,
		_w1656_,
		_w3153_,
		_w5561_,
		_w5649_
	);
	LUT3 #(
		.INIT('ha8)
	) name5187 (
		_w2000_,
		_w5648_,
		_w5649_,
		_w5650_
	);
	LUT3 #(
		.INIT('hc4)
	) name5188 (
		_w1869_,
		_w2556_,
		_w2729_,
		_w5651_
	);
	LUT3 #(
		.INIT('h2a)
	) name5189 (
		\P2_reg0_reg[1]/NET0131 ,
		_w3982_,
		_w5651_,
		_w5652_
	);
	LUT3 #(
		.INIT('h0d)
	) name5190 (
		_w3153_,
		_w5634_,
		_w5652_,
		_w5653_
	);
	LUT2 #(
		.INIT('hb)
	) name5191 (
		_w5650_,
		_w5653_,
		_w5654_
	);
	LUT4 #(
		.INIT('h1114)
	) name5192 (
		_w488_,
		_w989_,
		_w998_,
		_w602_,
		_w5655_
	);
	LUT2 #(
		.INIT('h4)
	) name5193 (
		_w1001_,
		_w2172_,
		_w5656_
	);
	LUT4 #(
		.INIT('h7800)
	) name5194 (
		_w996_,
		_w997_,
		_w1001_,
		_w2120_,
		_w5657_
	);
	LUT2 #(
		.INIT('h1)
	) name5195 (
		_w5656_,
		_w5657_,
		_w5658_
	);
	LUT4 #(
		.INIT('h80cc)
	) name5196 (
		_w1237_,
		_w2055_,
		_w5655_,
		_w5658_,
		_w5659_
	);
	LUT2 #(
		.INIT('h4)
	) name5197 (
		_w1001_,
		_w1120_,
		_w5660_
	);
	LUT3 #(
		.INIT('ha8)
	) name5198 (
		_w3511_,
		_w5659_,
		_w5660_,
		_w5661_
	);
	LUT4 #(
		.INIT('h50d0)
	) name5199 (
		_w1237_,
		_w2055_,
		_w5443_,
		_w5655_,
		_w5662_
	);
	LUT2 #(
		.INIT('h2)
	) name5200 (
		\P1_reg3_reg[0]/NET0131 ,
		_w5662_,
		_w5663_
	);
	LUT2 #(
		.INIT('he)
	) name5201 (
		_w5661_,
		_w5663_,
		_w5664_
	);
	LUT4 #(
		.INIT('h4000)
	) name5202 (
		_w1305_,
		_w1863_,
		_w1866_,
		_w1999_,
		_w5665_
	);
	LUT4 #(
		.INIT('h5600)
	) name5203 (
		_w1648_,
		_w1656_,
		_w1967_,
		_w5665_,
		_w5666_
	);
	LUT2 #(
		.INIT('h4)
	) name5204 (
		_w1660_,
		_w2033_,
		_w5667_
	);
	LUT4 #(
		.INIT('h0078)
	) name5205 (
		_w1654_,
		_w1655_,
		_w1660_,
		_w3443_,
		_w5668_
	);
	LUT2 #(
		.INIT('h1)
	) name5206 (
		_w5667_,
		_w5668_,
		_w5669_
	);
	LUT2 #(
		.INIT('h4)
	) name5207 (
		_w1660_,
		_w2029_,
		_w5670_
	);
	LUT4 #(
		.INIT('h0075)
	) name5208 (
		_w2903_,
		_w5666_,
		_w5669_,
		_w5670_,
		_w5671_
	);
	LUT4 #(
		.INIT('haaa2)
	) name5209 (
		\P2_reg3_reg[0]/NET0131 ,
		_w2556_,
		_w4194_,
		_w5666_,
		_w5672_
	);
	LUT3 #(
		.INIT('hf2)
	) name5210 (
		_w2556_,
		_w5671_,
		_w5672_,
		_w5673_
	);
	LUT4 #(
		.INIT('h80cc)
	) name5211 (
		_w1237_,
		_w2189_,
		_w5655_,
		_w5658_,
		_w5674_
	);
	LUT4 #(
		.INIT('h0200)
	) name5212 (
		\P1_reg3_reg[0]/NET0131 ,
		_w1096_,
		_w1098_,
		_w1101_,
		_w5675_
	);
	LUT3 #(
		.INIT('ha8)
	) name5213 (
		_w3511_,
		_w5674_,
		_w5675_,
		_w5676_
	);
	LUT4 #(
		.INIT('h0010)
	) name5214 (
		_w2171_,
		_w3173_,
		_w3511_,
		_w5093_,
		_w5677_
	);
	LUT4 #(
		.INIT('h5d00)
	) name5215 (
		_w1237_,
		_w2189_,
		_w5655_,
		_w5677_,
		_w5678_
	);
	LUT2 #(
		.INIT('h2)
	) name5216 (
		\P1_reg2_reg[0]/NET0131 ,
		_w5678_,
		_w5679_
	);
	LUT2 #(
		.INIT('he)
	) name5217 (
		_w5676_,
		_w5679_,
		_w5680_
	);
	LUT3 #(
		.INIT('h8a)
	) name5218 (
		_w3244_,
		_w5666_,
		_w5669_,
		_w5681_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name5219 (
		\P2_reg1_reg[0]/NET0131 ,
		_w2042_,
		_w3872_,
		_w3891_,
		_w5682_
	);
	LUT2 #(
		.INIT('he)
	) name5220 (
		_w5681_,
		_w5682_,
		_w5683_
	);
	LUT3 #(
		.INIT('h2a)
	) name5221 (
		\P1_reg0_reg[0]/NET0131 ,
		_w2332_,
		_w3563_,
		_w5684_
	);
	LUT4 #(
		.INIT('h80cc)
	) name5222 (
		_w1237_,
		_w3563_,
		_w5655_,
		_w5658_,
		_w5685_
	);
	LUT2 #(
		.INIT('he)
	) name5223 (
		_w5684_,
		_w5685_,
		_w5686_
	);
	LUT4 #(
		.INIT('h0200)
	) name5224 (
		\P2_reg3_reg[0]/NET0131 ,
		_w1863_,
		_w1866_,
		_w2028_,
		_w5687_
	);
	LUT4 #(
		.INIT('h0075)
	) name5225 (
		_w1298_,
		_w5666_,
		_w5669_,
		_w5687_,
		_w5688_
	);
	LUT4 #(
		.INIT('h2322)
	) name5226 (
		_w1298_,
		_w2032_,
		_w2033_,
		_w3266_,
		_w5689_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name5227 (
		\P2_reg2_reg[0]/NET0131 ,
		_w2556_,
		_w5666_,
		_w5689_,
		_w5690_
	);
	LUT3 #(
		.INIT('hf2)
	) name5228 (
		_w2556_,
		_w5688_,
		_w5690_,
		_w5691_
	);
	LUT2 #(
		.INIT('h2)
	) name5229 (
		\P1_reg1_reg[0]/NET0131 ,
		_w5449_,
		_w5692_
	);
	LUT4 #(
		.INIT('h80cc)
	) name5230 (
		_w1237_,
		_w3608_,
		_w5655_,
		_w5658_,
		_w5693_
	);
	LUT2 #(
		.INIT('he)
	) name5231 (
		_w5692_,
		_w5693_,
		_w5694_
	);
	LUT3 #(
		.INIT('h8a)
	) name5232 (
		_w3153_,
		_w5666_,
		_w5669_,
		_w5695_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5233 (
		\P2_reg0_reg[0]/NET0131 ,
		_w2736_,
		_w3982_,
		_w5651_,
		_w5696_
	);
	LUT2 #(
		.INIT('he)
	) name5234 (
		_w5695_,
		_w5696_,
		_w5697_
	);
	LUT3 #(
		.INIT('h48)
	) name5235 (
		\P1_IR_reg[25]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1247_,
		_w5698_
	);
	LUT3 #(
		.INIT('h0b)
	) name5236 (
		\P1_state_reg[0]/NET0131 ,
		_w1058_,
		_w5698_,
		_w5699_
	);
	LUT4 #(
		.INIT('ha060)
	) name5237 (
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w478_,
		_w5700_
	);
	LUT3 #(
		.INIT('hf1)
	) name5238 (
		\P1_state_reg[0]/NET0131 ,
		_w1040_,
		_w5700_,
		_w5701_
	);
	LUT2 #(
		.INIT('h2)
	) name5239 (
		\P1_state_reg[0]/NET0131 ,
		_w1279_,
		_w5702_
	);
	LUT4 #(
		.INIT('hff54)
	) name5240 (
		\P1_state_reg[0]/NET0131 ,
		_w1514_,
		_w1521_,
		_w5702_,
		_w5703_
	);
	LUT4 #(
		.INIT('h8828)
	) name5241 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1301_,
		_w5704_
	);
	LUT4 #(
		.INIT('hff54)
	) name5242 (
		\P1_state_reg[0]/NET0131 ,
		_w1452_,
		_w1478_,
		_w5704_,
		_w5705_
	);
	LUT3 #(
		.INIT('h48)
	) name5243 (
		\P1_IR_reg[26]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w573_,
		_w5706_
	);
	LUT3 #(
		.INIT('hf1)
	) name5244 (
		\P1_state_reg[0]/NET0131 ,
		_w1030_,
		_w5706_,
		_w5707_
	);
	LUT4 #(
		.INIT('h8828)
	) name5245 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1281_,
		_w5708_
	);
	LUT3 #(
		.INIT('hf1)
	) name5246 (
		\P1_state_reg[0]/NET0131 ,
		_w1505_,
		_w5708_,
		_w5709_
	);
	LUT4 #(
		.INIT('h2228)
	) name5247 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		_w1272_,
		_w1274_,
		_w5710_
	);
	LUT4 #(
		.INIT('hff54)
	) name5248 (
		\P1_state_reg[0]/NET0131 ,
		_w1531_,
		_w1533_,
		_w5710_,
		_w5711_
	);
	LUT3 #(
		.INIT('h28)
	) name5249 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[10]/NET0131 ,
		_w1767_,
		_w5712_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5250 (
		\P1_state_reg[0]/NET0131 ,
		_w1770_,
		_w1772_,
		_w5712_,
		_w5713_
	);
	LUT3 #(
		.INIT('h28)
	) name5251 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[11]/NET0131 ,
		_w1743_,
		_w5714_
	);
	LUT3 #(
		.INIT('h0b)
	) name5252 (
		\P1_state_reg[0]/NET0131 ,
		_w1746_,
		_w5714_,
		_w5715_
	);
	LUT4 #(
		.INIT('h8882)
	) name5253 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[12]/NET0131 ,
		_w1742_,
		_w1754_,
		_w5716_
	);
	LUT3 #(
		.INIT('h0b)
	) name5254 (
		\P1_state_reg[0]/NET0131 ,
		_w1758_,
		_w5716_,
		_w5717_
	);
	LUT4 #(
		.INIT('h8828)
	) name5255 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1262_,
		_w5718_
	);
	LUT3 #(
		.INIT('hf1)
	) name5256 (
		\P1_state_reg[0]/NET0131 ,
		_w1838_,
		_w5718_,
		_w5719_
	);
	LUT2 #(
		.INIT('h8)
	) name5257 (
		\P1_state_reg[0]/NET0131 ,
		_w1827_,
		_w5720_
	);
	LUT3 #(
		.INIT('hf1)
	) name5258 (
		\P1_state_reg[0]/NET0131 ,
		_w1829_,
		_w5720_,
		_w5721_
	);
	LUT3 #(
		.INIT('h28)
	) name5259 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[15]/NET0131 ,
		_w1814_,
		_w5722_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5260 (
		\P1_state_reg[0]/NET0131 ,
		_w1817_,
		_w1819_,
		_w5722_,
		_w5723_
	);
	LUT2 #(
		.INIT('h2)
	) name5261 (
		\P1_state_reg[0]/NET0131 ,
		_w1799_,
		_w5724_
	);
	LUT3 #(
		.INIT('h0b)
	) name5262 (
		\P1_state_reg[0]/NET0131 ,
		_w1801_,
		_w5724_,
		_w5725_
	);
	LUT2 #(
		.INIT('h8)
	) name5263 (
		\P1_state_reg[0]/NET0131 ,
		_w1607_,
		_w5726_
	);
	LUT4 #(
		.INIT('hff54)
	) name5264 (
		\P1_state_reg[0]/NET0131 ,
		_w1609_,
		_w1611_,
		_w5726_,
		_w5727_
	);
	LUT3 #(
		.INIT('h28)
	) name5265 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[18]/NET0131 ,
		_w1620_,
		_w5728_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5266 (
		\P1_state_reg[0]/NET0131 ,
		_w1623_,
		_w1625_,
		_w5728_,
		_w5729_
	);
	LUT3 #(
		.INIT('h28)
	) name5267 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[19]/NET0131 ,
		_w1264_,
		_w5730_
	);
	LUT3 #(
		.INIT('hf1)
	) name5268 (
		\P1_state_reg[0]/NET0131 ,
		_w1598_,
		_w5730_,
		_w5731_
	);
	LUT4 #(
		.INIT('h28a0)
	) name5269 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w5732_
	);
	LUT3 #(
		.INIT('hf4)
	) name5270 (
		\P1_state_reg[0]/NET0131 ,
		_w1650_,
		_w5732_,
		_w5733_
	);
	LUT3 #(
		.INIT('h82)
	) name5271 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[20]/NET0131 ,
		_w1272_,
		_w5734_
	);
	LUT3 #(
		.INIT('h0b)
	) name5272 (
		\P1_state_reg[0]/NET0131 ,
		_w1586_,
		_w5734_,
		_w5735_
	);
	LUT3 #(
		.INIT('h28)
	) name5273 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		_w1862_,
		_w5736_
	);
	LUT3 #(
		.INIT('h0b)
	) name5274 (
		\P1_state_reg[0]/NET0131 ,
		_w1568_,
		_w5736_,
		_w5737_
	);
	LUT4 #(
		.INIT('h8882)
	) name5275 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		_w1272_,
		_w1865_,
		_w5738_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5276 (
		\P1_state_reg[0]/NET0131 ,
		_w1555_,
		_w1559_,
		_w5738_,
		_w5739_
	);
	LUT3 #(
		.INIT('hf1)
	) name5277 (
		\P1_state_reg[0]/NET0131 ,
		_w1546_,
		_w2344_,
		_w5740_
	);
	LUT2 #(
		.INIT('h8)
	) name5278 (
		\P1_state_reg[0]/NET0131 ,
		_w1305_,
		_w5741_
	);
	LUT3 #(
		.INIT('hf1)
	) name5279 (
		\P1_state_reg[0]/NET0131 ,
		_w1441_,
		_w5741_,
		_w5742_
	);
	LUT3 #(
		.INIT('h28)
	) name5280 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[29]/NET0131 ,
		_w1381_,
		_w5743_
	);
	LUT3 #(
		.INIT('h0b)
	) name5281 (
		\P1_state_reg[0]/NET0131 ,
		_w1373_,
		_w5743_,
		_w5744_
	);
	LUT2 #(
		.INIT('h8)
	) name5282 (
		\P1_state_reg[0]/NET0131 ,
		_w1641_,
		_w5745_
	);
	LUT3 #(
		.INIT('hf1)
	) name5283 (
		\P1_state_reg[0]/NET0131 ,
		_w1640_,
		_w5745_,
		_w5746_
	);
	LUT2 #(
		.INIT('h8)
	) name5284 (
		\P1_state_reg[0]/NET0131 ,
		_w1378_,
		_w5747_
	);
	LUT3 #(
		.INIT('hf1)
	) name5285 (
		\P1_state_reg[0]/NET0131 ,
		_w2362_,
		_w5747_,
		_w5748_
	);
	LUT3 #(
		.INIT('h28)
	) name5286 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[3]/NET0131 ,
		_w1677_,
		_w5749_
	);
	LUT3 #(
		.INIT('hf1)
	) name5287 (
		\P1_state_reg[0]/NET0131 ,
		_w1680_,
		_w5749_,
		_w5750_
	);
	LUT4 #(
		.INIT('ha028)
	) name5288 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		_w1259_,
		_w5751_
	);
	LUT3 #(
		.INIT('hf4)
	) name5289 (
		\P1_state_reg[0]/NET0131 ,
		_w1663_,
		_w5751_,
		_w5752_
	);
	LUT2 #(
		.INIT('h2)
	) name5290 (
		\P1_state_reg[0]/NET0131 ,
		_w1724_,
		_w5753_
	);
	LUT3 #(
		.INIT('hf1)
	) name5291 (
		\P1_state_reg[0]/NET0131 ,
		_w1725_,
		_w5753_,
		_w5754_
	);
	LUT3 #(
		.INIT('h28)
	) name5292 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[6]/NET0131 ,
		_w1714_,
		_w5755_
	);
	LUT3 #(
		.INIT('h0b)
	) name5293 (
		\P1_state_reg[0]/NET0131 ,
		_w1716_,
		_w5755_,
		_w5756_
	);
	LUT3 #(
		.INIT('h28)
	) name5294 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		_w1703_,
		_w5757_
	);
	LUT3 #(
		.INIT('h0b)
	) name5295 (
		\P1_state_reg[0]/NET0131 ,
		_w1705_,
		_w5757_,
		_w5758_
	);
	LUT2 #(
		.INIT('h8)
	) name5296 (
		\P1_state_reg[0]/NET0131 ,
		_w1693_,
		_w5759_
	);
	LUT3 #(
		.INIT('hf1)
	) name5297 (
		\P1_state_reg[0]/NET0131 ,
		_w1694_,
		_w5759_,
		_w5760_
	);
	LUT3 #(
		.INIT('h28)
	) name5298 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w1781_,
		_w5761_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5299 (
		\P1_state_reg[0]/NET0131 ,
		_w1784_,
		_w1786_,
		_w5761_,
		_w5762_
	);
	LUT4 #(
		.INIT('ha060)
	) name5300 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w860_,
		_w5763_
	);
	LUT3 #(
		.INIT('hf1)
	) name5301 (
		\P1_state_reg[0]/NET0131 ,
		_w891_,
		_w5763_,
		_w5764_
	);
	LUT4 #(
		.INIT('ha060)
	) name5302 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w469_,
		_w5765_
	);
	LUT4 #(
		.INIT('hff54)
	) name5303 (
		\P1_state_reg[0]/NET0131 ,
		_w878_,
		_w880_,
		_w5765_,
		_w5766_
	);
	LUT2 #(
		.INIT('h8)
	) name5304 (
		\P1_state_reg[0]/NET0131 ,
		_w862_,
		_w5767_
	);
	LUT3 #(
		.INIT('hf1)
	) name5305 (
		\P1_state_reg[0]/NET0131 ,
		_w859_,
		_w5767_,
		_w5768_
	);
	LUT2 #(
		.INIT('h8)
	) name5306 (
		\P1_state_reg[0]/NET0131 ,
		_w850_,
		_w5769_
	);
	LUT3 #(
		.INIT('hf1)
	) name5307 (
		\P1_state_reg[0]/NET0131 ,
		_w849_,
		_w5769_,
		_w5770_
	);
	LUT2 #(
		.INIT('h2)
	) name5308 (
		\P1_state_reg[0]/NET0131 ,
		_w840_,
		_w5771_
	);
	LUT3 #(
		.INIT('hf1)
	) name5309 (
		\P1_state_reg[0]/NET0131 ,
		_w839_,
		_w5771_,
		_w5772_
	);
	LUT2 #(
		.INIT('h8)
	) name5310 (
		\P1_state_reg[0]/NET0131 ,
		_w831_,
		_w5773_
	);
	LUT3 #(
		.INIT('hf1)
	) name5311 (
		\P1_state_reg[0]/NET0131 ,
		_w829_,
		_w5773_,
		_w5774_
	);
	LUT3 #(
		.INIT('h48)
	) name5312 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w482_,
		_w5775_
	);
	LUT3 #(
		.INIT('hf1)
	) name5313 (
		\P1_state_reg[0]/NET0131 ,
		_w756_,
		_w5775_,
		_w5776_
	);
	LUT3 #(
		.INIT('h48)
	) name5314 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w746_,
		_w5777_
	);
	LUT4 #(
		.INIT('hff54)
	) name5315 (
		\P1_state_reg[0]/NET0131 ,
		_w742_,
		_w745_,
		_w5777_,
		_w5778_
	);
	LUT4 #(
		.INIT('h4448)
	) name5316 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w482_,
		_w731_,
		_w5779_
	);
	LUT4 #(
		.INIT('hff54)
	) name5317 (
		\P1_state_reg[0]/NET0131 ,
		_w727_,
		_w730_,
		_w5779_,
		_w5780_
	);
	LUT2 #(
		.INIT('h2)
	) name5318 (
		\P1_state_reg[0]/NET0131 ,
		_w718_,
		_w5781_
	);
	LUT3 #(
		.INIT('hf1)
	) name5319 (
		\P1_state_reg[0]/NET0131 ,
		_w717_,
		_w5781_,
		_w5782_
	);
	LUT4 #(
		.INIT('h6c00)
	) name5320 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5783_
	);
	LUT3 #(
		.INIT('hf4)
	) name5321 (
		\P1_state_reg[0]/NET0131 ,
		_w992_,
		_w5783_,
		_w5784_
	);
	LUT4 #(
		.INIT('h8884)
	) name5322 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w482_,
		_w1099_,
		_w5785_
	);
	LUT3 #(
		.INIT('h0b)
	) name5323 (
		\P1_state_reg[0]/NET0131 ,
		_w804_,
		_w5785_,
		_w5786_
	);
	LUT4 #(
		.INIT('h8884)
	) name5324 (
		\P1_IR_reg[21]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w746_,
		_w1095_,
		_w5787_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5325 (
		\P1_state_reg[0]/NET0131 ,
		_w793_,
		_w795_,
		_w5787_,
		_w5788_
	);
	LUT4 #(
		.INIT('h8884)
	) name5326 (
		\P1_IR_reg[22]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w482_,
		_w1097_,
		_w5789_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5327 (
		\P1_state_reg[0]/NET0131 ,
		_w773_,
		_w775_,
		_w5789_,
		_w5790_
	);
	LUT3 #(
		.INIT('hf1)
	) name5328 (
		\P1_state_reg[0]/NET0131 ,
		_w783_,
		_w1244_,
		_w5791_
	);
	LUT4 #(
		.INIT('h8884)
	) name5329 (
		\P1_IR_reg[24]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w482_,
		_w1250_,
		_w5792_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5330 (
		\P1_state_reg[0]/NET0131 ,
		_w1066_,
		_w1072_,
		_w5792_,
		_w5793_
	);
	LUT4 #(
		.INIT('h4448)
	) name5331 (
		\P1_IR_reg[28]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w482_,
		_w487_,
		_w5794_
	);
	LUT4 #(
		.INIT('hff54)
	) name5332 (
		\P1_state_reg[0]/NET0131 ,
		_w680_,
		_w701_,
		_w5794_,
		_w5795_
	);
	LUT3 #(
		.INIT('h84)
	) name5333 (
		\P1_IR_reg[29]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w583_,
		_w5796_
	);
	LUT3 #(
		.INIT('hf1)
	) name5334 (
		\P1_state_reg[0]/NET0131 ,
		_w673_,
		_w5796_,
		_w5797_
	);
	LUT2 #(
		.INIT('h8)
	) name5335 (
		\P1_state_reg[0]/NET0131 ,
		_w983_,
		_w5798_
	);
	LUT3 #(
		.INIT('hf1)
	) name5336 (
		\P1_state_reg[0]/NET0131 ,
		_w982_,
		_w5798_,
		_w5799_
	);
	LUT4 #(
		.INIT('h4448)
	) name5337 (
		\P1_IR_reg[30]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w573_,
		_w576_,
		_w5800_
	);
	LUT3 #(
		.INIT('hf1)
	) name5338 (
		\P1_state_reg[0]/NET0131 ,
		_w646_,
		_w5800_,
		_w5801_
	);
	LUT4 #(
		.INIT('h1000)
	) name5339 (
		\P1_IR_reg[29]/NET0131 ,
		\P1_IR_reg[30]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5802_
	);
	LUT2 #(
		.INIT('h8)
	) name5340 (
		_w574_,
		_w5802_,
		_w5803_
	);
	LUT2 #(
		.INIT('h8)
	) name5341 (
		_w478_,
		_w5803_,
		_w5804_
	);
	LUT3 #(
		.INIT('hf4)
	) name5342 (
		\P1_state_reg[0]/NET0131 ,
		_w569_,
		_w5804_,
		_w5805_
	);
	LUT3 #(
		.INIT('h48)
	) name5343 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w974_,
		_w5806_
	);
	LUT3 #(
		.INIT('hf1)
	) name5344 (
		\P1_state_reg[0]/NET0131 ,
		_w973_,
		_w5806_,
		_w5807_
	);
	LUT4 #(
		.INIT('hc060)
	) name5345 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w466_,
		_w5808_
	);
	LUT3 #(
		.INIT('hf4)
	) name5346 (
		\P1_state_reg[0]/NET0131 ,
		_w965_,
		_w5808_,
		_w5809_
	);
	LUT2 #(
		.INIT('h2)
	) name5347 (
		\P1_state_reg[0]/NET0131 ,
		_w955_,
		_w5810_
	);
	LUT4 #(
		.INIT('hff54)
	) name5348 (
		\P1_state_reg[0]/NET0131 ,
		_w951_,
		_w953_,
		_w5810_,
		_w5811_
	);
	LUT3 #(
		.INIT('h48)
	) name5349 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w931_,
		_w5812_
	);
	LUT3 #(
		.INIT('hf1)
	) name5350 (
		\P1_state_reg[0]/NET0131 ,
		_w930_,
		_w5812_,
		_w5813_
	);
	LUT4 #(
		.INIT('h4448)
	) name5351 (
		\P1_IR_reg[7]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w931_,
		_w941_,
		_w5814_
	);
	LUT3 #(
		.INIT('hf1)
	) name5352 (
		\P1_state_reg[0]/NET0131 ,
		_w940_,
		_w5814_,
		_w5815_
	);
	LUT3 #(
		.INIT('h48)
	) name5353 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w902_,
		_w5816_
	);
	LUT3 #(
		.INIT('hf1)
	) name5354 (
		\P1_state_reg[0]/NET0131 ,
		_w913_,
		_w5816_,
		_w5817_
	);
	LUT4 #(
		.INIT('h4448)
	) name5355 (
		\P1_IR_reg[9]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w902_,
		_w903_,
		_w5818_
	);
	LUT3 #(
		.INIT('hf1)
	) name5356 (
		\P1_state_reg[0]/NET0131 ,
		_w901_,
		_w5818_,
		_w5819_
	);
	LUT4 #(
		.INIT('h0200)
	) name5357 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[29]/NET0131 ,
		\P2_IR_reg[30]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w5820_
	);
	LUT2 #(
		.INIT('h8)
	) name5358 (
		_w1375_,
		_w5820_,
		_w5821_
	);
	LUT2 #(
		.INIT('h8)
	) name5359 (
		_w1301_,
		_w5821_,
		_w5822_
	);
	LUT3 #(
		.INIT('hf4)
	) name5360 (
		\P1_state_reg[0]/NET0131 ,
		_w2353_,
		_w5822_,
		_w5823_
	);
	LUT3 #(
		.INIT('h84)
	) name5361 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg1_reg[6]/NET0131 ,
		_w1714_,
		_w5824_
	);
	LUT3 #(
		.INIT('h12)
	) name5362 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg1_reg[6]/NET0131 ,
		_w1714_,
		_w5825_
	);
	LUT3 #(
		.INIT('h69)
	) name5363 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg1_reg[6]/NET0131 ,
		_w1714_,
		_w5826_
	);
	LUT3 #(
		.INIT('h48)
	) name5364 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg1_reg[3]/NET0131 ,
		_w1677_,
		_w5827_
	);
	LUT3 #(
		.INIT('h21)
	) name5365 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg1_reg[3]/NET0131 ,
		_w1677_,
		_w5828_
	);
	LUT2 #(
		.INIT('h8)
	) name5366 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w5829_
	);
	LUT3 #(
		.INIT('h4d)
	) name5367 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1651_,
		_w5829_,
		_w5830_
	);
	LUT4 #(
		.INIT('h080e)
	) name5368 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1641_,
		_w5828_,
		_w5830_,
		_w5831_
	);
	LUT4 #(
		.INIT('h444d)
	) name5369 (
		\P2_reg1_reg[4]/NET0131 ,
		_w1664_,
		_w5827_,
		_w5831_,
		_w5832_
	);
	LUT4 #(
		.INIT('h0d04)
	) name5370 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1724_,
		_w5826_,
		_w5832_,
		_w5833_
	);
	LUT2 #(
		.INIT('h4)
	) name5371 (
		_w1302_,
		_w1305_,
		_w5834_
	);
	LUT4 #(
		.INIT('h20b0)
	) name5372 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1724_,
		_w5826_,
		_w5832_,
		_w5835_
	);
	LUT3 #(
		.INIT('h02)
	) name5373 (
		_w5834_,
		_w5835_,
		_w5833_,
		_w5836_
	);
	LUT3 #(
		.INIT('h84)
	) name5374 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w1714_,
		_w5837_
	);
	LUT3 #(
		.INIT('h12)
	) name5375 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w1714_,
		_w5838_
	);
	LUT3 #(
		.INIT('h69)
	) name5376 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w1714_,
		_w5839_
	);
	LUT3 #(
		.INIT('h48)
	) name5377 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w1677_,
		_w5840_
	);
	LUT3 #(
		.INIT('h21)
	) name5378 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w1677_,
		_w5841_
	);
	LUT2 #(
		.INIT('h8)
	) name5379 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w5842_
	);
	LUT3 #(
		.INIT('h4d)
	) name5380 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1651_,
		_w5842_,
		_w5843_
	);
	LUT4 #(
		.INIT('h080e)
	) name5381 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1641_,
		_w5841_,
		_w5843_,
		_w5844_
	);
	LUT4 #(
		.INIT('h444d)
	) name5382 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1664_,
		_w5840_,
		_w5844_,
		_w5845_
	);
	LUT4 #(
		.INIT('h20b0)
	) name5383 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1724_,
		_w5839_,
		_w5845_,
		_w5846_
	);
	LUT4 #(
		.INIT('h0d04)
	) name5384 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1724_,
		_w5839_,
		_w5845_,
		_w5847_
	);
	LUT3 #(
		.INIT('h02)
	) name5385 (
		_w2340_,
		_w5847_,
		_w5846_,
		_w5848_
	);
	LUT4 #(
		.INIT('h00bf)
	) name5386 (
		_w1267_,
		_w1275_,
		_w1283_,
		_w1302_,
		_w5849_
	);
	LUT2 #(
		.INIT('h4)
	) name5387 (
		_w1305_,
		_w1715_,
		_w5850_
	);
	LUT2 #(
		.INIT('h4)
	) name5388 (
		_w5849_,
		_w5850_,
		_w5851_
	);
	LUT4 #(
		.INIT('h0777)
	) name5389 (
		_w1275_,
		_w1283_,
		_w1863_,
		_w1866_,
		_w5852_
	);
	LUT4 #(
		.INIT('h0c0d)
	) name5390 (
		_w1267_,
		_w1306_,
		_w2039_,
		_w5852_,
		_w5853_
	);
	LUT4 #(
		.INIT('h0013)
	) name5391 (
		\P2_addr_reg[6]/NET0131 ,
		_w5851_,
		_w5853_,
		_w5848_,
		_w5854_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5392 (
		\P1_state_reg[0]/NET0131 ,
		\P2_addr_reg[6]/NET0131 ,
		_w1267_,
		_w2341_,
		_w5855_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5393 (
		_w5288_,
		_w5836_,
		_w5854_,
		_w5855_,
		_w5856_
	);
	LUT4 #(
		.INIT('h2221)
	) name5394 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg1_reg[12]/NET0131 ,
		_w1742_,
		_w1754_,
		_w5857_
	);
	LUT3 #(
		.INIT('h12)
	) name5395 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w1743_,
		_w5858_
	);
	LUT3 #(
		.INIT('h12)
	) name5396 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg1_reg[10]/NET0131 ,
		_w1767_,
		_w5859_
	);
	LUT2 #(
		.INIT('h1)
	) name5397 (
		_w5858_,
		_w5859_,
		_w5860_
	);
	LUT3 #(
		.INIT('h12)
	) name5398 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg1_reg[9]/NET0131 ,
		_w1781_,
		_w5861_
	);
	LUT2 #(
		.INIT('h1)
	) name5399 (
		\P2_reg1_reg[8]/NET0131 ,
		_w1693_,
		_w5862_
	);
	LUT4 #(
		.INIT('h0d04)
	) name5400 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1724_,
		_w5824_,
		_w5832_,
		_w5863_
	);
	LUT3 #(
		.INIT('h12)
	) name5401 (
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg1_reg[7]/NET0131 ,
		_w1703_,
		_w5864_
	);
	LUT2 #(
		.INIT('h1)
	) name5402 (
		_w5825_,
		_w5864_,
		_w5865_
	);
	LUT3 #(
		.INIT('h84)
	) name5403 (
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg1_reg[7]/NET0131 ,
		_w1703_,
		_w5866_
	);
	LUT2 #(
		.INIT('h8)
	) name5404 (
		\P2_reg1_reg[8]/NET0131 ,
		_w1693_,
		_w5867_
	);
	LUT2 #(
		.INIT('h1)
	) name5405 (
		_w5866_,
		_w5867_,
		_w5868_
	);
	LUT4 #(
		.INIT('h1055)
	) name5406 (
		_w5862_,
		_w5863_,
		_w5865_,
		_w5868_,
		_w5869_
	);
	LUT3 #(
		.INIT('h84)
	) name5407 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg1_reg[9]/NET0131 ,
		_w1781_,
		_w5870_
	);
	LUT3 #(
		.INIT('h84)
	) name5408 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg1_reg[10]/NET0131 ,
		_w1767_,
		_w5871_
	);
	LUT2 #(
		.INIT('h1)
	) name5409 (
		_w5870_,
		_w5871_,
		_w5872_
	);
	LUT4 #(
		.INIT('h20aa)
	) name5410 (
		_w5860_,
		_w5861_,
		_w5869_,
		_w5872_,
		_w5873_
	);
	LUT4 #(
		.INIT('h4448)
	) name5411 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg1_reg[12]/NET0131 ,
		_w1742_,
		_w1754_,
		_w5874_
	);
	LUT3 #(
		.INIT('h84)
	) name5412 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w1743_,
		_w5875_
	);
	LUT2 #(
		.INIT('h1)
	) name5413 (
		_w5874_,
		_w5875_,
		_w5876_
	);
	LUT4 #(
		.INIT('ha060)
	) name5414 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[13]/NET0131 ,
		_w1262_,
		_w5877_
	);
	LUT4 #(
		.INIT('h0509)
	) name5415 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[13]/NET0131 ,
		_w1262_,
		_w5878_
	);
	LUT4 #(
		.INIT('h5a96)
	) name5416 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[13]/NET0131 ,
		_w1262_,
		_w5879_
	);
	LUT4 #(
		.INIT('h00ba)
	) name5417 (
		_w5857_,
		_w5873_,
		_w5876_,
		_w5879_,
		_w5880_
	);
	LUT4 #(
		.INIT('h4500)
	) name5418 (
		_w5857_,
		_w5873_,
		_w5876_,
		_w5879_,
		_w5881_
	);
	LUT3 #(
		.INIT('h02)
	) name5419 (
		_w5834_,
		_w5881_,
		_w5880_,
		_w5882_
	);
	LUT4 #(
		.INIT('ha060)
	) name5420 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[13]/NET0131 ,
		_w1262_,
		_w5883_
	);
	LUT4 #(
		.INIT('h0509)
	) name5421 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[13]/NET0131 ,
		_w1262_,
		_w5884_
	);
	LUT4 #(
		.INIT('h5a96)
	) name5422 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[13]/NET0131 ,
		_w1262_,
		_w5885_
	);
	LUT4 #(
		.INIT('h2221)
	) name5423 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg2_reg[12]/NET0131 ,
		_w1742_,
		_w1754_,
		_w5886_
	);
	LUT3 #(
		.INIT('h12)
	) name5424 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w1743_,
		_w5887_
	);
	LUT3 #(
		.INIT('h12)
	) name5425 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg2_reg[10]/NET0131 ,
		_w1767_,
		_w5888_
	);
	LUT2 #(
		.INIT('h1)
	) name5426 (
		_w5887_,
		_w5888_,
		_w5889_
	);
	LUT3 #(
		.INIT('h12)
	) name5427 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w1781_,
		_w5890_
	);
	LUT2 #(
		.INIT('h1)
	) name5428 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1693_,
		_w5891_
	);
	LUT4 #(
		.INIT('h0d04)
	) name5429 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1724_,
		_w5837_,
		_w5845_,
		_w5892_
	);
	LUT3 #(
		.INIT('h12)
	) name5430 (
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg2_reg[7]/NET0131 ,
		_w1703_,
		_w5893_
	);
	LUT2 #(
		.INIT('h1)
	) name5431 (
		_w5838_,
		_w5893_,
		_w5894_
	);
	LUT3 #(
		.INIT('h84)
	) name5432 (
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg2_reg[7]/NET0131 ,
		_w1703_,
		_w5895_
	);
	LUT2 #(
		.INIT('h8)
	) name5433 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1693_,
		_w5896_
	);
	LUT2 #(
		.INIT('h1)
	) name5434 (
		_w5895_,
		_w5896_,
		_w5897_
	);
	LUT4 #(
		.INIT('h1055)
	) name5435 (
		_w5891_,
		_w5892_,
		_w5894_,
		_w5897_,
		_w5898_
	);
	LUT3 #(
		.INIT('h84)
	) name5436 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w1781_,
		_w5899_
	);
	LUT3 #(
		.INIT('h84)
	) name5437 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg2_reg[10]/NET0131 ,
		_w1767_,
		_w5900_
	);
	LUT2 #(
		.INIT('h1)
	) name5438 (
		_w5899_,
		_w5900_,
		_w5901_
	);
	LUT4 #(
		.INIT('h20aa)
	) name5439 (
		_w5889_,
		_w5890_,
		_w5898_,
		_w5901_,
		_w5902_
	);
	LUT3 #(
		.INIT('h84)
	) name5440 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w1743_,
		_w5903_
	);
	LUT4 #(
		.INIT('h4448)
	) name5441 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg2_reg[12]/NET0131 ,
		_w1742_,
		_w1754_,
		_w5904_
	);
	LUT2 #(
		.INIT('h1)
	) name5442 (
		_w5903_,
		_w5904_,
		_w5905_
	);
	LUT3 #(
		.INIT('h45)
	) name5443 (
		_w5886_,
		_w5902_,
		_w5905_,
		_w5906_
	);
	LUT3 #(
		.INIT('h54)
	) name5444 (
		\P2_addr_reg[13]/NET0131 ,
		_w1267_,
		_w5852_,
		_w5907_
	);
	LUT2 #(
		.INIT('h1)
	) name5445 (
		_w1305_,
		_w1836_,
		_w5908_
	);
	LUT4 #(
		.INIT('h50f3)
	) name5446 (
		_w1302_,
		_w5853_,
		_w5907_,
		_w5908_,
		_w5909_
	);
	LUT4 #(
		.INIT('hd700)
	) name5447 (
		_w2340_,
		_w5885_,
		_w5906_,
		_w5909_,
		_w5910_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5448 (
		\P1_state_reg[0]/NET0131 ,
		\P2_addr_reg[13]/NET0131 ,
		_w1267_,
		_w2341_,
		_w5911_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5449 (
		_w4125_,
		_w5882_,
		_w5910_,
		_w5911_,
		_w5912_
	);
	LUT2 #(
		.INIT('h6)
	) name5450 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w5913_
	);
	LUT3 #(
		.INIT('h80)
	) name5451 (
		_w1302_,
		_w1305_,
		_w5913_,
		_w5914_
	);
	LUT4 #(
		.INIT('hf95f)
	) name5452 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w1302_,
		_w1305_,
		_w5915_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name5453 (
		_w1267_,
		_w2341_,
		_w5914_,
		_w5915_,
		_w5916_
	);
	LUT3 #(
		.INIT('h08)
	) name5454 (
		\P2_addr_reg[0]/NET0131 ,
		_w1306_,
		_w2039_,
		_w5917_
	);
	LUT4 #(
		.INIT('h1d3f)
	) name5455 (
		\P2_addr_reg[0]/NET0131 ,
		_w1284_,
		_w1659_,
		_w1867_,
		_w5918_
	);
	LUT4 #(
		.INIT('h0032)
	) name5456 (
		_w1267_,
		_w5917_,
		_w5918_,
		_w5916_,
		_w5919_
	);
	LUT3 #(
		.INIT('h4e)
	) name5457 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[0]/NET0131 ,
		_w5919_,
		_w5920_
	);
	LUT3 #(
		.INIT('h69)
	) name5458 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg2_reg[10]/NET0131 ,
		_w1767_,
		_w5921_
	);
	LUT4 #(
		.INIT('h5510)
	) name5459 (
		_w5891_,
		_w5892_,
		_w5894_,
		_w5895_,
		_w5922_
	);
	LUT2 #(
		.INIT('h1)
	) name5460 (
		_w5896_,
		_w5899_,
		_w5923_
	);
	LUT4 #(
		.INIT('h4044)
	) name5461 (
		_w5890_,
		_w5921_,
		_w5922_,
		_w5923_,
		_w5924_
	);
	LUT4 #(
		.INIT('h2322)
	) name5462 (
		_w5890_,
		_w5921_,
		_w5922_,
		_w5923_,
		_w5925_
	);
	LUT3 #(
		.INIT('h02)
	) name5463 (
		_w2340_,
		_w5925_,
		_w5924_,
		_w5926_
	);
	LUT3 #(
		.INIT('h69)
	) name5464 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg1_reg[10]/NET0131 ,
		_w1767_,
		_w5927_
	);
	LUT4 #(
		.INIT('h5510)
	) name5465 (
		_w5862_,
		_w5863_,
		_w5865_,
		_w5866_,
		_w5928_
	);
	LUT2 #(
		.INIT('h1)
	) name5466 (
		_w5867_,
		_w5870_,
		_w5929_
	);
	LUT3 #(
		.INIT('h45)
	) name5467 (
		_w5861_,
		_w5928_,
		_w5929_,
		_w5930_
	);
	LUT3 #(
		.INIT('h54)
	) name5468 (
		\P2_addr_reg[10]/NET0131 ,
		_w1267_,
		_w5852_,
		_w5931_
	);
	LUT2 #(
		.INIT('h4)
	) name5469 (
		_w1305_,
		_w1768_,
		_w5932_
	);
	LUT4 #(
		.INIT('h50f3)
	) name5470 (
		_w1302_,
		_w5853_,
		_w5931_,
		_w5932_,
		_w5933_
	);
	LUT4 #(
		.INIT('hd700)
	) name5471 (
		_w5834_,
		_w5927_,
		_w5930_,
		_w5933_,
		_w5934_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5472 (
		\P1_state_reg[0]/NET0131 ,
		\P2_addr_reg[10]/NET0131 ,
		_w1267_,
		_w2341_,
		_w5935_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5473 (
		_w4102_,
		_w5926_,
		_w5934_,
		_w5935_,
		_w5936_
	);
	LUT2 #(
		.INIT('h2)
	) name5474 (
		_w5873_,
		_w5875_,
		_w5937_
	);
	LUT3 #(
		.INIT('h69)
	) name5475 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w1743_,
		_w5938_
	);
	LUT4 #(
		.INIT('h1055)
	) name5476 (
		_w5859_,
		_w5861_,
		_w5869_,
		_w5872_,
		_w5939_
	);
	LUT3 #(
		.INIT('ha8)
	) name5477 (
		_w5834_,
		_w5938_,
		_w5939_,
		_w5940_
	);
	LUT2 #(
		.INIT('h4)
	) name5478 (
		_w5937_,
		_w5940_,
		_w5941_
	);
	LUT2 #(
		.INIT('h2)
	) name5479 (
		_w5902_,
		_w5903_,
		_w5942_
	);
	LUT3 #(
		.INIT('h69)
	) name5480 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w1743_,
		_w5943_
	);
	LUT4 #(
		.INIT('h1055)
	) name5481 (
		_w5888_,
		_w5890_,
		_w5898_,
		_w5901_,
		_w5944_
	);
	LUT3 #(
		.INIT('ha8)
	) name5482 (
		_w2340_,
		_w5943_,
		_w5944_,
		_w5945_
	);
	LUT3 #(
		.INIT('h54)
	) name5483 (
		\P2_addr_reg[11]/NET0131 ,
		_w1267_,
		_w5852_,
		_w5946_
	);
	LUT2 #(
		.INIT('h4)
	) name5484 (
		_w1305_,
		_w1744_,
		_w5947_
	);
	LUT4 #(
		.INIT('h50f3)
	) name5485 (
		_w1302_,
		_w5853_,
		_w5946_,
		_w5947_,
		_w5948_
	);
	LUT3 #(
		.INIT('hb0)
	) name5486 (
		_w5942_,
		_w5945_,
		_w5948_,
		_w5949_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5487 (
		\P1_state_reg[0]/NET0131 ,
		\P2_addr_reg[11]/NET0131 ,
		_w1267_,
		_w2341_,
		_w5950_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5488 (
		_w4601_,
		_w5941_,
		_w5949_,
		_w5950_,
		_w5951_
	);
	LUT4 #(
		.INIT('h9996)
	) name5489 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg1_reg[12]/NET0131 ,
		_w1742_,
		_w1754_,
		_w5952_
	);
	LUT4 #(
		.INIT('h2322)
	) name5490 (
		_w5861_,
		_w5871_,
		_w5928_,
		_w5929_,
		_w5953_
	);
	LUT4 #(
		.INIT('h0301)
	) name5491 (
		_w5860_,
		_w5875_,
		_w5952_,
		_w5953_,
		_w5954_
	);
	LUT4 #(
		.INIT('hc0e0)
	) name5492 (
		_w5860_,
		_w5875_,
		_w5952_,
		_w5953_,
		_w5955_
	);
	LUT3 #(
		.INIT('h02)
	) name5493 (
		_w5834_,
		_w5955_,
		_w5954_,
		_w5956_
	);
	LUT4 #(
		.INIT('h9996)
	) name5494 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg2_reg[12]/NET0131 ,
		_w1742_,
		_w1754_,
		_w5957_
	);
	LUT4 #(
		.INIT('h2322)
	) name5495 (
		_w5890_,
		_w5900_,
		_w5922_,
		_w5923_,
		_w5958_
	);
	LUT3 #(
		.INIT('h31)
	) name5496 (
		_w5889_,
		_w5903_,
		_w5958_,
		_w5959_
	);
	LUT3 #(
		.INIT('h54)
	) name5497 (
		\P2_addr_reg[12]/NET0131 ,
		_w1267_,
		_w5852_,
		_w5960_
	);
	LUT2 #(
		.INIT('h4)
	) name5498 (
		_w1305_,
		_w1755_,
		_w5961_
	);
	LUT4 #(
		.INIT('h50f3)
	) name5499 (
		_w1302_,
		_w5853_,
		_w5960_,
		_w5961_,
		_w5962_
	);
	LUT4 #(
		.INIT('h7d00)
	) name5500 (
		_w2340_,
		_w5957_,
		_w5959_,
		_w5962_,
		_w5963_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5501 (
		\P1_state_reg[0]/NET0131 ,
		\P2_addr_reg[12]/NET0131 ,
		_w1267_,
		_w2341_,
		_w5964_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5502 (
		_w3706_,
		_w5956_,
		_w5963_,
		_w5964_,
		_w5965_
	);
	LUT2 #(
		.INIT('h8)
	) name5503 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1827_,
		_w5966_
	);
	LUT2 #(
		.INIT('h1)
	) name5504 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1827_,
		_w5967_
	);
	LUT2 #(
		.INIT('h6)
	) name5505 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1827_,
		_w5968_
	);
	LUT4 #(
		.INIT('h5054)
	) name5506 (
		_w5857_,
		_w5860_,
		_w5875_,
		_w5953_,
		_w5969_
	);
	LUT2 #(
		.INIT('h1)
	) name5507 (
		_w5874_,
		_w5877_,
		_w5970_
	);
	LUT4 #(
		.INIT('h4044)
	) name5508 (
		_w5878_,
		_w5968_,
		_w5969_,
		_w5970_,
		_w5971_
	);
	LUT4 #(
		.INIT('h2322)
	) name5509 (
		_w5878_,
		_w5968_,
		_w5969_,
		_w5970_,
		_w5972_
	);
	LUT3 #(
		.INIT('h02)
	) name5510 (
		_w5834_,
		_w5972_,
		_w5971_,
		_w5973_
	);
	LUT2 #(
		.INIT('h8)
	) name5511 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1827_,
		_w5974_
	);
	LUT2 #(
		.INIT('h1)
	) name5512 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1827_,
		_w5975_
	);
	LUT2 #(
		.INIT('h6)
	) name5513 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1827_,
		_w5976_
	);
	LUT4 #(
		.INIT('h5054)
	) name5514 (
		_w5886_,
		_w5889_,
		_w5903_,
		_w5958_,
		_w5977_
	);
	LUT2 #(
		.INIT('h1)
	) name5515 (
		_w5883_,
		_w5904_,
		_w5978_
	);
	LUT3 #(
		.INIT('h45)
	) name5516 (
		_w5884_,
		_w5977_,
		_w5978_,
		_w5979_
	);
	LUT3 #(
		.INIT('h54)
	) name5517 (
		\P2_addr_reg[14]/NET0131 ,
		_w1267_,
		_w5852_,
		_w5980_
	);
	LUT2 #(
		.INIT('h4)
	) name5518 (
		_w1305_,
		_w1827_,
		_w5981_
	);
	LUT4 #(
		.INIT('h50f3)
	) name5519 (
		_w1302_,
		_w5853_,
		_w5980_,
		_w5981_,
		_w5982_
	);
	LUT4 #(
		.INIT('hd700)
	) name5520 (
		_w2340_,
		_w5976_,
		_w5979_,
		_w5982_,
		_w5983_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5521 (
		\P1_state_reg[0]/NET0131 ,
		\P2_addr_reg[14]/NET0131 ,
		_w1267_,
		_w2341_,
		_w5984_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5522 (
		_w4621_,
		_w5973_,
		_w5983_,
		_w5984_,
		_w5985_
	);
	LUT3 #(
		.INIT('h84)
	) name5523 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w1814_,
		_w5986_
	);
	LUT3 #(
		.INIT('h12)
	) name5524 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w1814_,
		_w5987_
	);
	LUT3 #(
		.INIT('h69)
	) name5525 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w1814_,
		_w5988_
	);
	LUT4 #(
		.INIT('h0045)
	) name5526 (
		_w5857_,
		_w5873_,
		_w5876_,
		_w5878_,
		_w5989_
	);
	LUT3 #(
		.INIT('h07)
	) name5527 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1827_,
		_w5877_,
		_w5990_
	);
	LUT4 #(
		.INIT('h4044)
	) name5528 (
		_w5967_,
		_w5988_,
		_w5989_,
		_w5990_,
		_w5991_
	);
	LUT4 #(
		.INIT('h2322)
	) name5529 (
		_w5967_,
		_w5988_,
		_w5989_,
		_w5990_,
		_w5992_
	);
	LUT3 #(
		.INIT('h02)
	) name5530 (
		_w5834_,
		_w5992_,
		_w5991_,
		_w5993_
	);
	LUT3 #(
		.INIT('h12)
	) name5531 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w1814_,
		_w5994_
	);
	LUT3 #(
		.INIT('h84)
	) name5532 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w1814_,
		_w5995_
	);
	LUT3 #(
		.INIT('h69)
	) name5533 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w1814_,
		_w5996_
	);
	LUT4 #(
		.INIT('h1011)
	) name5534 (
		_w5884_,
		_w5886_,
		_w5902_,
		_w5905_,
		_w5997_
	);
	LUT3 #(
		.INIT('h07)
	) name5535 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1827_,
		_w5883_,
		_w5998_
	);
	LUT3 #(
		.INIT('h45)
	) name5536 (
		_w5975_,
		_w5997_,
		_w5998_,
		_w5999_
	);
	LUT3 #(
		.INIT('h54)
	) name5537 (
		\P2_addr_reg[15]/NET0131 ,
		_w1267_,
		_w5852_,
		_w6000_
	);
	LUT2 #(
		.INIT('h4)
	) name5538 (
		_w1305_,
		_w1815_,
		_w6001_
	);
	LUT4 #(
		.INIT('h50f3)
	) name5539 (
		_w1302_,
		_w5853_,
		_w6000_,
		_w6001_,
		_w6002_
	);
	LUT4 #(
		.INIT('hd700)
	) name5540 (
		_w2340_,
		_w5996_,
		_w5999_,
		_w6002_,
		_w6003_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5541 (
		\P1_state_reg[0]/NET0131 ,
		\P2_addr_reg[15]/NET0131 ,
		_w1267_,
		_w2341_,
		_w6004_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5542 (
		_w4145_,
		_w5993_,
		_w6003_,
		_w6004_,
		_w6005_
	);
	LUT2 #(
		.INIT('h8)
	) name5543 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1799_,
		_w6006_
	);
	LUT2 #(
		.INIT('h1)
	) name5544 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1799_,
		_w6007_
	);
	LUT2 #(
		.INIT('h6)
	) name5545 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1799_,
		_w6008_
	);
	LUT4 #(
		.INIT('h1011)
	) name5546 (
		_w5884_,
		_w5975_,
		_w5977_,
		_w5978_,
		_w6009_
	);
	LUT2 #(
		.INIT('h1)
	) name5547 (
		_w5974_,
		_w5995_,
		_w6010_
	);
	LUT4 #(
		.INIT('h2322)
	) name5548 (
		_w5994_,
		_w6008_,
		_w6009_,
		_w6010_,
		_w6011_
	);
	LUT4 #(
		.INIT('h4044)
	) name5549 (
		_w5994_,
		_w6008_,
		_w6009_,
		_w6010_,
		_w6012_
	);
	LUT3 #(
		.INIT('h02)
	) name5550 (
		_w2340_,
		_w6012_,
		_w6011_,
		_w6013_
	);
	LUT2 #(
		.INIT('h8)
	) name5551 (
		\P2_reg1_reg[16]/NET0131 ,
		_w1799_,
		_w6014_
	);
	LUT2 #(
		.INIT('h1)
	) name5552 (
		\P2_reg1_reg[16]/NET0131 ,
		_w1799_,
		_w6015_
	);
	LUT2 #(
		.INIT('h6)
	) name5553 (
		\P2_reg1_reg[16]/NET0131 ,
		_w1799_,
		_w6016_
	);
	LUT2 #(
		.INIT('h1)
	) name5554 (
		_w5967_,
		_w5987_,
		_w6017_
	);
	LUT4 #(
		.INIT('h4500)
	) name5555 (
		_w5878_,
		_w5969_,
		_w5970_,
		_w6017_,
		_w6018_
	);
	LUT3 #(
		.INIT('he8)
	) name5556 (
		\P2_reg1_reg[15]/NET0131 ,
		_w1815_,
		_w5966_,
		_w6019_
	);
	LUT4 #(
		.INIT('h2228)
	) name5557 (
		_w5834_,
		_w6016_,
		_w6018_,
		_w6019_,
		_w6020_
	);
	LUT3 #(
		.INIT('h54)
	) name5558 (
		\P2_addr_reg[16]/NET0131 ,
		_w1267_,
		_w5852_,
		_w6021_
	);
	LUT2 #(
		.INIT('h4)
	) name5559 (
		_w1305_,
		_w1799_,
		_w6022_
	);
	LUT4 #(
		.INIT('h50f3)
	) name5560 (
		_w1302_,
		_w5853_,
		_w6021_,
		_w6022_,
		_w6023_
	);
	LUT2 #(
		.INIT('h4)
	) name5561 (
		_w6020_,
		_w6023_,
		_w6024_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5562 (
		\P1_state_reg[0]/NET0131 ,
		\P2_addr_reg[16]/NET0131 ,
		_w1267_,
		_w2341_,
		_w6025_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5563 (
		_w3727_,
		_w6013_,
		_w6024_,
		_w6025_,
		_w6026_
	);
	LUT2 #(
		.INIT('h1)
	) name5564 (
		\P2_reg2_reg[17]/NET0131 ,
		_w1607_,
		_w6027_
	);
	LUT2 #(
		.INIT('h8)
	) name5565 (
		\P2_reg2_reg[17]/NET0131 ,
		_w1607_,
		_w6028_
	);
	LUT2 #(
		.INIT('h6)
	) name5566 (
		\P2_reg2_reg[17]/NET0131 ,
		_w1607_,
		_w6029_
	);
	LUT4 #(
		.INIT('h1011)
	) name5567 (
		_w5975_,
		_w5994_,
		_w5997_,
		_w5998_,
		_w6030_
	);
	LUT2 #(
		.INIT('h1)
	) name5568 (
		_w5995_,
		_w6006_,
		_w6031_
	);
	LUT4 #(
		.INIT('h4044)
	) name5569 (
		_w6007_,
		_w6029_,
		_w6030_,
		_w6031_,
		_w6032_
	);
	LUT4 #(
		.INIT('h2322)
	) name5570 (
		_w6007_,
		_w6029_,
		_w6030_,
		_w6031_,
		_w6033_
	);
	LUT3 #(
		.INIT('h02)
	) name5571 (
		_w2340_,
		_w6033_,
		_w6032_,
		_w6034_
	);
	LUT2 #(
		.INIT('h1)
	) name5572 (
		\P2_reg1_reg[17]/NET0131 ,
		_w1607_,
		_w6035_
	);
	LUT2 #(
		.INIT('h8)
	) name5573 (
		\P2_reg1_reg[17]/NET0131 ,
		_w1607_,
		_w6036_
	);
	LUT2 #(
		.INIT('h6)
	) name5574 (
		\P2_reg1_reg[17]/NET0131 ,
		_w1607_,
		_w6037_
	);
	LUT2 #(
		.INIT('h1)
	) name5575 (
		_w5986_,
		_w6014_,
		_w6038_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5576 (
		_w5989_,
		_w5990_,
		_w6017_,
		_w6038_,
		_w6039_
	);
	LUT4 #(
		.INIT('ha082)
	) name5577 (
		_w5834_,
		_w6015_,
		_w6037_,
		_w6039_,
		_w6040_
	);
	LUT3 #(
		.INIT('h54)
	) name5578 (
		\P2_addr_reg[17]/NET0131 ,
		_w1267_,
		_w5852_,
		_w6041_
	);
	LUT2 #(
		.INIT('h4)
	) name5579 (
		_w1305_,
		_w1607_,
		_w6042_
	);
	LUT4 #(
		.INIT('h50f3)
	) name5580 (
		_w1302_,
		_w5853_,
		_w6041_,
		_w6042_,
		_w6043_
	);
	LUT2 #(
		.INIT('h4)
	) name5581 (
		_w6040_,
		_w6043_,
		_w6044_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5582 (
		\P1_state_reg[0]/NET0131 ,
		\P2_addr_reg[17]/NET0131 ,
		_w1267_,
		_w2341_,
		_w6045_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5583 (
		_w3412_,
		_w6034_,
		_w6044_,
		_w6045_,
		_w6046_
	);
	LUT4 #(
		.INIT('h936c)
	) name5584 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[1]/NET0131 ,
		_w6047_
	);
	LUT2 #(
		.INIT('h6)
	) name5585 (
		_w5842_,
		_w6047_,
		_w6048_
	);
	LUT3 #(
		.INIT('h80)
	) name5586 (
		_w1302_,
		_w1305_,
		_w6048_,
		_w6049_
	);
	LUT4 #(
		.INIT('h936c)
	) name5587 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[1]/NET0131 ,
		_w6050_
	);
	LUT2 #(
		.INIT('h6)
	) name5588 (
		_w5829_,
		_w6050_,
		_w6051_
	);
	LUT4 #(
		.INIT('hb9fd)
	) name5589 (
		_w1302_,
		_w1305_,
		_w1651_,
		_w6051_,
		_w6052_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name5590 (
		_w1267_,
		_w2341_,
		_w6049_,
		_w6052_,
		_w6053_
	);
	LUT3 #(
		.INIT('h08)
	) name5591 (
		\P2_addr_reg[1]/NET0131 ,
		_w1306_,
		_w2039_,
		_w6054_
	);
	LUT4 #(
		.INIT('h1d3f)
	) name5592 (
		\P2_addr_reg[1]/NET0131 ,
		_w1284_,
		_w1652_,
		_w1867_,
		_w6055_
	);
	LUT4 #(
		.INIT('h0032)
	) name5593 (
		_w1267_,
		_w6054_,
		_w6055_,
		_w6053_,
		_w6056_
	);
	LUT3 #(
		.INIT('h4e)
	) name5594 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[1]/NET0131 ,
		_w6056_,
		_w6057_
	);
	LUT2 #(
		.INIT('h6)
	) name5595 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1641_,
		_w6058_
	);
	LUT2 #(
		.INIT('h9)
	) name5596 (
		_w5843_,
		_w6058_,
		_w6059_
	);
	LUT3 #(
		.INIT('h80)
	) name5597 (
		_w1302_,
		_w1305_,
		_w6059_,
		_w6060_
	);
	LUT2 #(
		.INIT('h6)
	) name5598 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1641_,
		_w6061_
	);
	LUT2 #(
		.INIT('h9)
	) name5599 (
		_w5830_,
		_w6061_,
		_w6062_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name5600 (
		_w1302_,
		_w1305_,
		_w1641_,
		_w6062_,
		_w6063_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name5601 (
		_w1267_,
		_w2341_,
		_w6060_,
		_w6063_,
		_w6064_
	);
	LUT3 #(
		.INIT('h08)
	) name5602 (
		\P2_addr_reg[2]/NET0131 ,
		_w1306_,
		_w2039_,
		_w6065_
	);
	LUT4 #(
		.INIT('h1d3f)
	) name5603 (
		\P2_addr_reg[2]/NET0131 ,
		_w1284_,
		_w1642_,
		_w1867_,
		_w6066_
	);
	LUT4 #(
		.INIT('h0032)
	) name5604 (
		_w1267_,
		_w6065_,
		_w6066_,
		_w6064_,
		_w6067_
	);
	LUT3 #(
		.INIT('h4e)
	) name5605 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[2]/NET0131 ,
		_w6067_,
		_w6068_
	);
	LUT3 #(
		.INIT('h96)
	) name5606 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w1677_,
		_w6069_
	);
	LUT4 #(
		.INIT('h718e)
	) name5607 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1641_,
		_w5843_,
		_w6069_,
		_w6070_
	);
	LUT3 #(
		.INIT('h80)
	) name5608 (
		_w1302_,
		_w1305_,
		_w6070_,
		_w6071_
	);
	LUT3 #(
		.INIT('h96)
	) name5609 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg1_reg[3]/NET0131 ,
		_w1677_,
		_w6072_
	);
	LUT4 #(
		.INIT('h718e)
	) name5610 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1641_,
		_w5830_,
		_w6072_,
		_w6073_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name5611 (
		_w1302_,
		_w1305_,
		_w1678_,
		_w6073_,
		_w6074_
	);
	LUT3 #(
		.INIT('h45)
	) name5612 (
		_w2341_,
		_w6071_,
		_w6074_,
		_w6075_
	);
	LUT4 #(
		.INIT('h0007)
	) name5613 (
		_w1275_,
		_w1283_,
		_w1302_,
		_w1305_,
		_w6076_
	);
	LUT3 #(
		.INIT('ha8)
	) name5614 (
		\P2_addr_reg[3]/NET0131 ,
		_w2341_,
		_w6076_,
		_w6077_
	);
	LUT3 #(
		.INIT('h15)
	) name5615 (
		_w1267_,
		_w1284_,
		_w1679_,
		_w6078_
	);
	LUT4 #(
		.INIT('hccc4)
	) name5616 (
		\P2_addr_reg[3]/NET0131 ,
		_w1267_,
		_w1302_,
		_w1305_,
		_w6079_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5617 (
		\P1_state_reg[0]/NET0131 ,
		_w6071_,
		_w6074_,
		_w6079_,
		_w6080_
	);
	LUT4 #(
		.INIT('hef00)
	) name5618 (
		_w6077_,
		_w6075_,
		_w6078_,
		_w6080_,
		_w6081_
	);
	LUT2 #(
		.INIT('he)
	) name5619 (
		_w5267_,
		_w6081_,
		_w6082_
	);
	LUT4 #(
		.INIT('h3c96)
	) name5620 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_reg2_reg[4]/NET0131 ,
		_w1259_,
		_w6083_
	);
	LUT3 #(
		.INIT('he0)
	) name5621 (
		_w5840_,
		_w5844_,
		_w6083_,
		_w6084_
	);
	LUT3 #(
		.INIT('h01)
	) name5622 (
		_w5840_,
		_w5844_,
		_w6083_,
		_w6085_
	);
	LUT4 #(
		.INIT('h0008)
	) name5623 (
		_w1302_,
		_w1305_,
		_w6085_,
		_w6084_,
		_w6086_
	);
	LUT3 #(
		.INIT('h02)
	) name5624 (
		_w1302_,
		_w1305_,
		_w1664_,
		_w6087_
	);
	LUT4 #(
		.INIT('h3c96)
	) name5625 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_reg1_reg[4]/NET0131 ,
		_w1259_,
		_w6088_
	);
	LUT3 #(
		.INIT('he0)
	) name5626 (
		_w5827_,
		_w5831_,
		_w6088_,
		_w6089_
	);
	LUT3 #(
		.INIT('h01)
	) name5627 (
		_w5827_,
		_w5831_,
		_w6088_,
		_w6090_
	);
	LUT4 #(
		.INIT('h0004)
	) name5628 (
		_w1302_,
		_w1305_,
		_w6090_,
		_w6089_,
		_w6091_
	);
	LUT4 #(
		.INIT('h5554)
	) name5629 (
		_w2341_,
		_w6087_,
		_w6091_,
		_w6086_,
		_w6092_
	);
	LUT3 #(
		.INIT('ha8)
	) name5630 (
		\P2_addr_reg[4]/NET0131 ,
		_w2341_,
		_w6076_,
		_w6093_
	);
	LUT3 #(
		.INIT('h15)
	) name5631 (
		_w1267_,
		_w1284_,
		_w1665_,
		_w6094_
	);
	LUT3 #(
		.INIT('h10)
	) name5632 (
		_w6092_,
		_w6093_,
		_w6094_,
		_w6095_
	);
	LUT4 #(
		.INIT('hccc4)
	) name5633 (
		\P2_addr_reg[4]/NET0131 ,
		_w1267_,
		_w1302_,
		_w1305_,
		_w6096_
	);
	LUT4 #(
		.INIT('h0100)
	) name5634 (
		_w6087_,
		_w6091_,
		_w6086_,
		_w6096_,
		_w6097_
	);
	LUT2 #(
		.INIT('h2)
	) name5635 (
		\P1_state_reg[0]/NET0131 ,
		_w6097_,
		_w6098_
	);
	LUT3 #(
		.INIT('hba)
	) name5636 (
		_w5000_,
		_w6095_,
		_w6098_,
		_w6099_
	);
	LUT2 #(
		.INIT('h9)
	) name5637 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1724_,
		_w6100_
	);
	LUT4 #(
		.INIT('h4004)
	) name5638 (
		_w1302_,
		_w1305_,
		_w5832_,
		_w6100_,
		_w6101_
	);
	LUT3 #(
		.INIT('h54)
	) name5639 (
		\P2_addr_reg[5]/NET0131 ,
		_w1267_,
		_w5852_,
		_w6102_
	);
	LUT3 #(
		.INIT('h31)
	) name5640 (
		_w5853_,
		_w6101_,
		_w6102_,
		_w6103_
	);
	LUT2 #(
		.INIT('h9)
	) name5641 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1724_,
		_w6104_
	);
	LUT4 #(
		.INIT('h8008)
	) name5642 (
		_w1302_,
		_w1305_,
		_w5845_,
		_w6104_,
		_w6105_
	);
	LUT4 #(
		.INIT('h0504)
	) name5643 (
		\P2_addr_reg[5]/NET0131 ,
		_w1267_,
		_w1302_,
		_w5852_,
		_w6106_
	);
	LUT2 #(
		.INIT('h1)
	) name5644 (
		_w1305_,
		_w1724_,
		_w6107_
	);
	LUT3 #(
		.INIT('h45)
	) name5645 (
		_w6105_,
		_w6106_,
		_w6107_,
		_w6108_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5646 (
		\P1_state_reg[0]/NET0131 ,
		\P2_addr_reg[5]/NET0131 ,
		_w1267_,
		_w2341_,
		_w6109_
	);
	LUT4 #(
		.INIT('hbfaa)
	) name5647 (
		_w5017_,
		_w6103_,
		_w6108_,
		_w6109_,
		_w6110_
	);
	LUT3 #(
		.INIT('h69)
	) name5648 (
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg1_reg[7]/NET0131 ,
		_w1703_,
		_w6111_
	);
	LUT4 #(
		.INIT('ha802)
	) name5649 (
		_w5834_,
		_w5825_,
		_w5863_,
		_w6111_,
		_w6112_
	);
	LUT3 #(
		.INIT('h69)
	) name5650 (
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg2_reg[7]/NET0131 ,
		_w1703_,
		_w6113_
	);
	LUT4 #(
		.INIT('ha802)
	) name5651 (
		_w2340_,
		_w5838_,
		_w5892_,
		_w6113_,
		_w6114_
	);
	LUT3 #(
		.INIT('h54)
	) name5652 (
		\P2_addr_reg[7]/NET0131 ,
		_w1267_,
		_w5852_,
		_w6115_
	);
	LUT2 #(
		.INIT('h4)
	) name5653 (
		_w1305_,
		_w1704_,
		_w6116_
	);
	LUT4 #(
		.INIT('h50f3)
	) name5654 (
		_w1302_,
		_w5853_,
		_w6115_,
		_w6116_,
		_w6117_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5655 (
		\P1_state_reg[0]/NET0131 ,
		\P2_addr_reg[7]/NET0131 ,
		_w1267_,
		_w2341_,
		_w6118_
	);
	LUT4 #(
		.INIT('hef00)
	) name5656 (
		_w6114_,
		_w6112_,
		_w6117_,
		_w6118_,
		_w6119_
	);
	LUT2 #(
		.INIT('he)
	) name5657 (
		_w5035_,
		_w6119_,
		_w6120_
	);
	LUT2 #(
		.INIT('h6)
	) name5658 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1693_,
		_w6121_
	);
	LUT4 #(
		.INIT('hf400)
	) name5659 (
		_w5892_,
		_w5894_,
		_w5895_,
		_w6121_,
		_w6122_
	);
	LUT4 #(
		.INIT('h000b)
	) name5660 (
		_w5892_,
		_w5894_,
		_w5895_,
		_w6121_,
		_w6123_
	);
	LUT3 #(
		.INIT('h02)
	) name5661 (
		_w2340_,
		_w6123_,
		_w6122_,
		_w6124_
	);
	LUT2 #(
		.INIT('h6)
	) name5662 (
		\P2_reg1_reg[8]/NET0131 ,
		_w1693_,
		_w6125_
	);
	LUT4 #(
		.INIT('hf400)
	) name5663 (
		_w5863_,
		_w5865_,
		_w5866_,
		_w6125_,
		_w6126_
	);
	LUT4 #(
		.INIT('h000b)
	) name5664 (
		_w5863_,
		_w5865_,
		_w5866_,
		_w6125_,
		_w6127_
	);
	LUT3 #(
		.INIT('h02)
	) name5665 (
		_w5834_,
		_w6127_,
		_w6126_,
		_w6128_
	);
	LUT3 #(
		.INIT('h54)
	) name5666 (
		\P2_addr_reg[8]/NET0131 ,
		_w1267_,
		_w5852_,
		_w6129_
	);
	LUT2 #(
		.INIT('h4)
	) name5667 (
		_w1305_,
		_w1693_,
		_w6130_
	);
	LUT4 #(
		.INIT('h50f3)
	) name5668 (
		_w1302_,
		_w5853_,
		_w6129_,
		_w6130_,
		_w6131_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5669 (
		\P1_state_reg[0]/NET0131 ,
		\P2_addr_reg[8]/NET0131 ,
		_w1267_,
		_w2341_,
		_w6132_
	);
	LUT4 #(
		.INIT('hef00)
	) name5670 (
		_w6128_,
		_w6124_,
		_w6131_,
		_w6132_,
		_w6133_
	);
	LUT2 #(
		.INIT('he)
	) name5671 (
		_w4658_,
		_w6133_,
		_w6134_
	);
	LUT3 #(
		.INIT('h69)
	) name5672 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg1_reg[9]/NET0131 ,
		_w1781_,
		_w6135_
	);
	LUT3 #(
		.INIT('h28)
	) name5673 (
		_w5834_,
		_w5869_,
		_w6135_,
		_w6136_
	);
	LUT3 #(
		.INIT('h69)
	) name5674 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w1781_,
		_w6137_
	);
	LUT3 #(
		.INIT('h28)
	) name5675 (
		_w2340_,
		_w5898_,
		_w6137_,
		_w6138_
	);
	LUT3 #(
		.INIT('h54)
	) name5676 (
		\P2_addr_reg[9]/NET0131 ,
		_w1267_,
		_w5852_,
		_w6139_
	);
	LUT2 #(
		.INIT('h4)
	) name5677 (
		_w1305_,
		_w1782_,
		_w6140_
	);
	LUT4 #(
		.INIT('h50f3)
	) name5678 (
		_w1302_,
		_w5853_,
		_w6139_,
		_w6140_,
		_w6141_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5679 (
		\P1_state_reg[0]/NET0131 ,
		\P2_addr_reg[9]/NET0131 ,
		_w1267_,
		_w2341_,
		_w6142_
	);
	LUT4 #(
		.INIT('hef00)
	) name5680 (
		_w6138_,
		_w6136_,
		_w6141_,
		_w6142_,
		_w6143_
	);
	LUT2 #(
		.INIT('he)
	) name5681 (
		_w4165_,
		_w6143_,
		_w6144_
	);
	LUT3 #(
		.INIT('h84)
	) name5682 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w1620_,
		_w6145_
	);
	LUT3 #(
		.INIT('h12)
	) name5683 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w1620_,
		_w6146_
	);
	LUT3 #(
		.INIT('h69)
	) name5684 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w1620_,
		_w6147_
	);
	LUT4 #(
		.INIT('h1011)
	) name5685 (
		_w5994_,
		_w6007_,
		_w6009_,
		_w6010_,
		_w6148_
	);
	LUT4 #(
		.INIT('h153f)
	) name5686 (
		\P2_reg2_reg[16]/NET0131 ,
		\P2_reg2_reg[17]/NET0131 ,
		_w1607_,
		_w1799_,
		_w6149_
	);
	LUT4 #(
		.INIT('h4044)
	) name5687 (
		_w6027_,
		_w6147_,
		_w6148_,
		_w6149_,
		_w6150_
	);
	LUT4 #(
		.INIT('h2322)
	) name5688 (
		_w6027_,
		_w6147_,
		_w6148_,
		_w6149_,
		_w6151_
	);
	LUT3 #(
		.INIT('h02)
	) name5689 (
		_w2340_,
		_w6151_,
		_w6150_,
		_w6152_
	);
	LUT3 #(
		.INIT('h84)
	) name5690 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg1_reg[18]/NET0131 ,
		_w1620_,
		_w6153_
	);
	LUT3 #(
		.INIT('h12)
	) name5691 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg1_reg[18]/NET0131 ,
		_w1620_,
		_w6154_
	);
	LUT3 #(
		.INIT('h69)
	) name5692 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg1_reg[18]/NET0131 ,
		_w1620_,
		_w6155_
	);
	LUT4 #(
		.INIT('h153f)
	) name5693 (
		\P2_reg1_reg[16]/NET0131 ,
		\P2_reg1_reg[17]/NET0131 ,
		_w1607_,
		_w1799_,
		_w6156_
	);
	LUT4 #(
		.INIT('hab00)
	) name5694 (
		_w6015_,
		_w6018_,
		_w6019_,
		_w6156_,
		_w6157_
	);
	LUT4 #(
		.INIT('ha082)
	) name5695 (
		_w5834_,
		_w6035_,
		_w6155_,
		_w6157_,
		_w6158_
	);
	LUT3 #(
		.INIT('h54)
	) name5696 (
		\P2_addr_reg[18]/NET0131 ,
		_w1267_,
		_w5852_,
		_w6159_
	);
	LUT2 #(
		.INIT('h4)
	) name5697 (
		_w1305_,
		_w1621_,
		_w6160_
	);
	LUT4 #(
		.INIT('h50f3)
	) name5698 (
		_w1302_,
		_w5853_,
		_w6159_,
		_w6160_,
		_w6161_
	);
	LUT2 #(
		.INIT('h4)
	) name5699 (
		_w6158_,
		_w6161_,
		_w6162_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5700 (
		\P1_state_reg[0]/NET0131 ,
		\P2_addr_reg[18]/NET0131 ,
		_w1267_,
		_w2341_,
		_w6163_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5701 (
		_w3430_,
		_w6152_,
		_w6162_,
		_w6163_,
		_w6164_
	);
	LUT2 #(
		.INIT('h1)
	) name5702 (
		_w6035_,
		_w6154_,
		_w6165_
	);
	LUT4 #(
		.INIT('hcd00)
	) name5703 (
		_w6015_,
		_w6036_,
		_w6039_,
		_w6165_,
		_w6166_
	);
	LUT4 #(
		.INIT('h2221)
	) name5704 (
		\P2_reg1_reg[19]/NET0131 ,
		_w1595_,
		_w6153_,
		_w6166_,
		_w6167_
	);
	LUT4 #(
		.INIT('h4448)
	) name5705 (
		\P2_reg1_reg[19]/NET0131 ,
		_w1595_,
		_w6153_,
		_w6166_,
		_w6168_
	);
	LUT3 #(
		.INIT('h02)
	) name5706 (
		_w5834_,
		_w6168_,
		_w6167_,
		_w6169_
	);
	LUT4 #(
		.INIT('h2322)
	) name5707 (
		_w6007_,
		_w6028_,
		_w6030_,
		_w6031_,
		_w6170_
	);
	LUT2 #(
		.INIT('h1)
	) name5708 (
		_w6027_,
		_w6146_,
		_w6171_
	);
	LUT3 #(
		.INIT('h45)
	) name5709 (
		_w6145_,
		_w6170_,
		_w6171_,
		_w6172_
	);
	LUT3 #(
		.INIT('h96)
	) name5710 (
		\P2_IR_reg[19]/NET0131 ,
		\P2_reg2_reg[19]/NET0131 ,
		_w1264_,
		_w6173_
	);
	LUT3 #(
		.INIT('h54)
	) name5711 (
		\P2_addr_reg[19]/NET0131 ,
		_w1267_,
		_w5852_,
		_w6174_
	);
	LUT2 #(
		.INIT('h4)
	) name5712 (
		_w1305_,
		_w1595_,
		_w6175_
	);
	LUT4 #(
		.INIT('h50f3)
	) name5713 (
		_w1302_,
		_w5853_,
		_w6174_,
		_w6175_,
		_w6176_
	);
	LUT4 #(
		.INIT('h7d00)
	) name5714 (
		_w2340_,
		_w6172_,
		_w6173_,
		_w6176_,
		_w6177_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5715 (
		\P1_state_reg[0]/NET0131 ,
		\P2_addr_reg[19]/NET0131 ,
		_w1267_,
		_w2341_,
		_w6178_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5716 (
		_w3447_,
		_w6169_,
		_w6177_,
		_w6178_,
		_w6179_
	);
	LUT2 #(
		.INIT('h8)
	) name5717 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg2_reg[0]/NET0131 ,
		_w6180_
	);
	LUT2 #(
		.INIT('h6)
	) name5718 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg2_reg[0]/NET0131 ,
		_w6181_
	);
	LUT2 #(
		.INIT('h8)
	) name5719 (
		_w479_,
		_w488_,
		_w6182_
	);
	LUT2 #(
		.INIT('h8)
	) name5720 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg1_reg[0]/NET0131 ,
		_w6183_
	);
	LUT2 #(
		.INIT('h6)
	) name5721 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg1_reg[0]/NET0131 ,
		_w6184_
	);
	LUT4 #(
		.INIT('h37bf)
	) name5722 (
		_w479_,
		_w488_,
		_w6181_,
		_w6184_,
		_w6185_
	);
	LUT4 #(
		.INIT('h8882)
	) name5723 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[28]/NET0131 ,
		_w482_,
		_w487_,
		_w6186_
	);
	LUT3 #(
		.INIT('h40)
	) name5724 (
		\P1_addr_reg[2]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6187_
	);
	LUT4 #(
		.INIT('h8adf)
	) name5725 (
		_w1252_,
		_w6186_,
		_w6185_,
		_w6187_,
		_w6188_
	);
	LUT2 #(
		.INIT('h1)
	) name5726 (
		_w1236_,
		_w1252_,
		_w6189_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5727 (
		\P1_addr_reg[2]/NET0131 ,
		_w479_,
		_w488_,
		_w983_,
		_w6190_
	);
	LUT2 #(
		.INIT('h6)
	) name5728 (
		\P1_reg1_reg[2]/NET0131 ,
		_w983_,
		_w6191_
	);
	LUT3 #(
		.INIT('hb2)
	) name5729 (
		\P1_reg1_reg[1]/NET0131 ,
		_w991_,
		_w6183_,
		_w6192_
	);
	LUT2 #(
		.INIT('h6)
	) name5730 (
		_w6191_,
		_w6192_,
		_w6193_
	);
	LUT2 #(
		.INIT('h6)
	) name5731 (
		\P1_reg2_reg[2]/NET0131 ,
		_w983_,
		_w6194_
	);
	LUT3 #(
		.INIT('hb2)
	) name5732 (
		\P1_reg2_reg[1]/NET0131 ,
		_w991_,
		_w6180_,
		_w6195_
	);
	LUT2 #(
		.INIT('h6)
	) name5733 (
		_w6194_,
		_w6195_,
		_w6196_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name5734 (
		_w479_,
		_w488_,
		_w6193_,
		_w6196_,
		_w6197_
	);
	LUT2 #(
		.INIT('h8)
	) name5735 (
		_w6190_,
		_w6197_,
		_w6198_
	);
	LUT4 #(
		.INIT('h04ee)
	) name5736 (
		_w1243_,
		_w6188_,
		_w6189_,
		_w6198_,
		_w6199_
	);
	LUT3 #(
		.INIT('he2)
	) name5737 (
		\P1_reg3_reg[2]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6199_,
		_w6200_
	);
	LUT3 #(
		.INIT('h40)
	) name5738 (
		\P1_addr_reg[4]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6201_
	);
	LUT4 #(
		.INIT('h8adf)
	) name5739 (
		_w1252_,
		_w6186_,
		_w6185_,
		_w6201_,
		_w6202_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5740 (
		\P1_addr_reg[4]/NET0131 ,
		_w479_,
		_w488_,
		_w963_,
		_w6203_
	);
	LUT4 #(
		.INIT('h3c96)
	) name5741 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_reg2_reg[4]/NET0131 ,
		_w466_,
		_w6204_
	);
	LUT3 #(
		.INIT('h21)
	) name5742 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w974_,
		_w6205_
	);
	LUT3 #(
		.INIT('h48)
	) name5743 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w974_,
		_w6206_
	);
	LUT4 #(
		.INIT('h0017)
	) name5744 (
		\P1_reg2_reg[2]/NET0131 ,
		_w983_,
		_w6195_,
		_w6206_,
		_w6207_
	);
	LUT3 #(
		.INIT('ha9)
	) name5745 (
		_w6204_,
		_w6205_,
		_w6207_,
		_w6208_
	);
	LUT4 #(
		.INIT('h3c96)
	) name5746 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_reg1_reg[4]/NET0131 ,
		_w466_,
		_w6209_
	);
	LUT3 #(
		.INIT('h21)
	) name5747 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg1_reg[3]/NET0131 ,
		_w974_,
		_w6210_
	);
	LUT3 #(
		.INIT('h48)
	) name5748 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg1_reg[3]/NET0131 ,
		_w974_,
		_w6211_
	);
	LUT4 #(
		.INIT('h0017)
	) name5749 (
		\P1_reg1_reg[2]/NET0131 ,
		_w983_,
		_w6192_,
		_w6211_,
		_w6212_
	);
	LUT3 #(
		.INIT('ha9)
	) name5750 (
		_w6209_,
		_w6210_,
		_w6212_,
		_w6213_
	);
	LUT4 #(
		.INIT('h37bf)
	) name5751 (
		_w479_,
		_w488_,
		_w6208_,
		_w6213_,
		_w6214_
	);
	LUT2 #(
		.INIT('h8)
	) name5752 (
		_w6203_,
		_w6214_,
		_w6215_
	);
	LUT4 #(
		.INIT('h10fa)
	) name5753 (
		_w1243_,
		_w6189_,
		_w6202_,
		_w6215_,
		_w6216_
	);
	LUT3 #(
		.INIT('he2)
	) name5754 (
		\P1_reg3_reg[4]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6216_,
		_w6217_
	);
	LUT4 #(
		.INIT('h5f5d)
	) name5755 (
		\P1_state_reg[0]/NET0131 ,
		_w1267_,
		_w1306_,
		_w5852_,
		_w6218_
	);
	LUT4 #(
		.INIT('h5051)
	) name5756 (
		_w489_,
		_w1236_,
		_w1243_,
		_w1252_,
		_w6219_
	);
	LUT2 #(
		.INIT('hd)
	) name5757 (
		\P1_state_reg[0]/NET0131 ,
		_w6219_,
		_w6220_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name5758 (
		\P1_state_reg[0]/NET0131 ,
		_w1236_,
		_w1243_,
		_w1252_,
		_w6221_
	);
	LUT3 #(
		.INIT('h48)
	) name5759 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg1_reg[8]/NET0131 ,
		_w902_,
		_w6222_
	);
	LUT3 #(
		.INIT('h21)
	) name5760 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg1_reg[8]/NET0131 ,
		_w902_,
		_w6223_
	);
	LUT3 #(
		.INIT('h96)
	) name5761 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg1_reg[8]/NET0131 ,
		_w902_,
		_w6224_
	);
	LUT3 #(
		.INIT('h21)
	) name5762 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_reg1_reg[6]/NET0131 ,
		_w931_,
		_w6225_
	);
	LUT3 #(
		.INIT('h48)
	) name5763 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_reg1_reg[6]/NET0131 ,
		_w931_,
		_w6226_
	);
	LUT4 #(
		.INIT('h888e)
	) name5764 (
		\P1_reg1_reg[4]/NET0131 ,
		_w963_,
		_w6210_,
		_w6212_,
		_w6227_
	);
	LUT3 #(
		.INIT('hb2)
	) name5765 (
		\P1_reg1_reg[5]/NET0131 ,
		_w955_,
		_w6227_,
		_w6228_
	);
	LUT4 #(
		.INIT('h040d)
	) name5766 (
		\P1_reg1_reg[5]/NET0131 ,
		_w955_,
		_w6226_,
		_w6227_,
		_w6229_
	);
	LUT4 #(
		.INIT('h7771)
	) name5767 (
		\P1_reg1_reg[7]/NET0131 ,
		_w942_,
		_w6225_,
		_w6229_,
		_w6230_
	);
	LUT3 #(
		.INIT('h82)
	) name5768 (
		_w6182_,
		_w6224_,
		_w6230_,
		_w6231_
	);
	LUT3 #(
		.INIT('h48)
	) name5769 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg2_reg[8]/NET0131 ,
		_w902_,
		_w6232_
	);
	LUT3 #(
		.INIT('h21)
	) name5770 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg2_reg[8]/NET0131 ,
		_w902_,
		_w6233_
	);
	LUT3 #(
		.INIT('h96)
	) name5771 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg2_reg[8]/NET0131 ,
		_w902_,
		_w6234_
	);
	LUT4 #(
		.INIT('h4448)
	) name5772 (
		\P1_IR_reg[7]/NET0131 ,
		\P1_reg2_reg[7]/NET0131 ,
		_w931_,
		_w941_,
		_w6235_
	);
	LUT4 #(
		.INIT('h2221)
	) name5773 (
		\P1_IR_reg[7]/NET0131 ,
		\P1_reg2_reg[7]/NET0131 ,
		_w931_,
		_w941_,
		_w6236_
	);
	LUT3 #(
		.INIT('h21)
	) name5774 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_reg2_reg[6]/NET0131 ,
		_w931_,
		_w6237_
	);
	LUT3 #(
		.INIT('h48)
	) name5775 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_reg2_reg[6]/NET0131 ,
		_w931_,
		_w6238_
	);
	LUT4 #(
		.INIT('h888e)
	) name5776 (
		\P1_reg2_reg[4]/NET0131 ,
		_w963_,
		_w6205_,
		_w6207_,
		_w6239_
	);
	LUT4 #(
		.INIT('h040d)
	) name5777 (
		\P1_reg2_reg[5]/NET0131 ,
		_w955_,
		_w6238_,
		_w6239_,
		_w6240_
	);
	LUT4 #(
		.INIT('h7771)
	) name5778 (
		\P1_reg2_reg[7]/NET0131 ,
		_w942_,
		_w6237_,
		_w6240_,
		_w6241_
	);
	LUT4 #(
		.INIT('hf7f4)
	) name5779 (
		\P1_addr_reg[8]/NET0131 ,
		_w479_,
		_w488_,
		_w914_,
		_w6242_
	);
	LUT4 #(
		.INIT('h7d00)
	) name5780 (
		_w1245_,
		_w6234_,
		_w6241_,
		_w6242_,
		_w6243_
	);
	LUT4 #(
		.INIT('h007f)
	) name5781 (
		\P1_addr_reg[8]/NET0131 ,
		_w1236_,
		_w3511_,
		_w4185_,
		_w6244_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5782 (
		_w6221_,
		_w6231_,
		_w6243_,
		_w6244_,
		_w6245_
	);
	LUT3 #(
		.INIT('h96)
	) name5783 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_reg2_reg[6]/NET0131 ,
		_w931_,
		_w6246_
	);
	LUT4 #(
		.INIT('hb200)
	) name5784 (
		\P1_reg2_reg[5]/NET0131 ,
		_w955_,
		_w6239_,
		_w6246_,
		_w6247_
	);
	LUT4 #(
		.INIT('h004d)
	) name5785 (
		\P1_reg2_reg[5]/NET0131 ,
		_w955_,
		_w6239_,
		_w6246_,
		_w6248_
	);
	LUT3 #(
		.INIT('h02)
	) name5786 (
		_w1245_,
		_w6248_,
		_w6247_,
		_w6249_
	);
	LUT3 #(
		.INIT('h96)
	) name5787 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_reg1_reg[6]/NET0131 ,
		_w931_,
		_w6250_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5788 (
		\P1_addr_reg[6]/NET0131 ,
		_w479_,
		_w488_,
		_w932_,
		_w6251_
	);
	LUT4 #(
		.INIT('hd700)
	) name5789 (
		_w6182_,
		_w6228_,
		_w6250_,
		_w6251_,
		_w6252_
	);
	LUT4 #(
		.INIT('h007f)
	) name5790 (
		\P1_addr_reg[6]/NET0131 ,
		_w1236_,
		_w3511_,
		_w5053_,
		_w6253_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5791 (
		_w6221_,
		_w6249_,
		_w6252_,
		_w6253_,
		_w6254_
	);
	LUT4 #(
		.INIT('h0006)
	) name5792 (
		\P1_reg1_reg[7]/NET0131 ,
		_w942_,
		_w6225_,
		_w6229_,
		_w6255_
	);
	LUT4 #(
		.INIT('h9996)
	) name5793 (
		\P1_IR_reg[7]/NET0131 ,
		\P1_reg1_reg[7]/NET0131 ,
		_w931_,
		_w941_,
		_w6256_
	);
	LUT4 #(
		.INIT('haa02)
	) name5794 (
		_w6182_,
		_w6225_,
		_w6229_,
		_w6256_,
		_w6257_
	);
	LUT2 #(
		.INIT('h4)
	) name5795 (
		_w6255_,
		_w6257_,
		_w6258_
	);
	LUT4 #(
		.INIT('h0006)
	) name5796 (
		\P1_reg2_reg[7]/NET0131 ,
		_w942_,
		_w6237_,
		_w6240_,
		_w6259_
	);
	LUT4 #(
		.INIT('h9996)
	) name5797 (
		\P1_IR_reg[7]/NET0131 ,
		\P1_reg2_reg[7]/NET0131 ,
		_w931_,
		_w941_,
		_w6260_
	);
	LUT4 #(
		.INIT('haa02)
	) name5798 (
		_w1245_,
		_w6237_,
		_w6240_,
		_w6260_,
		_w6261_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5799 (
		\P1_addr_reg[7]/NET0131 ,
		_w479_,
		_w488_,
		_w942_,
		_w6262_
	);
	LUT3 #(
		.INIT('hb0)
	) name5800 (
		_w6259_,
		_w6261_,
		_w6262_,
		_w6263_
	);
	LUT3 #(
		.INIT('h40)
	) name5801 (
		\P1_addr_reg[7]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6264_
	);
	LUT2 #(
		.INIT('h2)
	) name5802 (
		_w3511_,
		_w6264_,
		_w6265_
	);
	LUT4 #(
		.INIT('hef00)
	) name5803 (
		_w1236_,
		_w6258_,
		_w6263_,
		_w6265_,
		_w6266_
	);
	LUT4 #(
		.INIT('h1311)
	) name5804 (
		_w1244_,
		_w5071_,
		_w6258_,
		_w6263_,
		_w6267_
	);
	LUT2 #(
		.INIT('hb)
	) name5805 (
		_w6266_,
		_w6267_,
		_w6268_
	);
	LUT3 #(
		.INIT('h40)
	) name5806 (
		\P1_addr_reg[3]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6269_
	);
	LUT3 #(
		.INIT('h51)
	) name5807 (
		_w1244_,
		_w3511_,
		_w6269_,
		_w6270_
	);
	LUT3 #(
		.INIT('h15)
	) name5808 (
		_w489_,
		_w1236_,
		_w3511_,
		_w6271_
	);
	LUT4 #(
		.INIT('ha888)
	) name5809 (
		\P1_addr_reg[3]/NET0131 ,
		_w489_,
		_w1236_,
		_w3511_,
		_w6272_
	);
	LUT3 #(
		.INIT('h96)
	) name5810 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w974_,
		_w6273_
	);
	LUT4 #(
		.INIT('h17e8)
	) name5811 (
		\P1_reg2_reg[2]/NET0131 ,
		_w983_,
		_w6195_,
		_w6273_,
		_w6274_
	);
	LUT3 #(
		.INIT('h40)
	) name5812 (
		_w479_,
		_w488_,
		_w6274_,
		_w6275_
	);
	LUT3 #(
		.INIT('h96)
	) name5813 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg1_reg[3]/NET0131 ,
		_w974_,
		_w6276_
	);
	LUT4 #(
		.INIT('h17e8)
	) name5814 (
		\P1_reg1_reg[2]/NET0131 ,
		_w983_,
		_w6192_,
		_w6276_,
		_w6277_
	);
	LUT4 #(
		.INIT('h67ef)
	) name5815 (
		_w479_,
		_w488_,
		_w975_,
		_w6277_,
		_w6278_
	);
	LUT2 #(
		.INIT('h4)
	) name5816 (
		_w6275_,
		_w6278_,
		_w6279_
	);
	LUT4 #(
		.INIT('hbabb)
	) name5817 (
		_w4982_,
		_w6270_,
		_w6272_,
		_w6279_,
		_w6280_
	);
	LUT2 #(
		.INIT('h2)
	) name5818 (
		\P1_reg3_reg[0]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6281_
	);
	LUT3 #(
		.INIT('h40)
	) name5819 (
		\P1_addr_reg[0]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6282_
	);
	LUT3 #(
		.INIT('h51)
	) name5820 (
		_w1244_,
		_w3511_,
		_w6282_,
		_w6283_
	);
	LUT4 #(
		.INIT('ha888)
	) name5821 (
		\P1_addr_reg[0]/NET0131 ,
		_w489_,
		_w1236_,
		_w3511_,
		_w6284_
	);
	LUT2 #(
		.INIT('h4)
	) name5822 (
		_w479_,
		_w6186_,
		_w6285_
	);
	LUT2 #(
		.INIT('h2)
	) name5823 (
		_w6185_,
		_w6285_,
		_w6286_
	);
	LUT4 #(
		.INIT('hbabb)
	) name5824 (
		_w6281_,
		_w6283_,
		_w6284_,
		_w6286_,
		_w6287_
	);
	LUT3 #(
		.INIT('h40)
	) name5825 (
		\P1_addr_reg[10]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6288_
	);
	LUT3 #(
		.INIT('h51)
	) name5826 (
		_w1244_,
		_w3511_,
		_w6288_,
		_w6289_
	);
	LUT4 #(
		.INIT('ha060)
	) name5827 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[10]/NET0131 ,
		_w860_,
		_w6290_
	);
	LUT4 #(
		.INIT('h0509)
	) name5828 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[10]/NET0131 ,
		_w860_,
		_w6291_
	);
	LUT4 #(
		.INIT('h5a96)
	) name5829 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[10]/NET0131 ,
		_w860_,
		_w6292_
	);
	LUT4 #(
		.INIT('h2221)
	) name5830 (
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg1_reg[9]/NET0131 ,
		_w902_,
		_w903_,
		_w6293_
	);
	LUT4 #(
		.INIT('h4448)
	) name5831 (
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg1_reg[9]/NET0131 ,
		_w902_,
		_w903_,
		_w6294_
	);
	LUT4 #(
		.INIT('h00d4)
	) name5832 (
		\P1_reg1_reg[8]/NET0131 ,
		_w914_,
		_w6230_,
		_w6294_,
		_w6295_
	);
	LUT4 #(
		.INIT('h8882)
	) name5833 (
		_w6182_,
		_w6292_,
		_w6293_,
		_w6295_,
		_w6296_
	);
	LUT4 #(
		.INIT('ha060)
	) name5834 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w860_,
		_w6297_
	);
	LUT4 #(
		.INIT('h0509)
	) name5835 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w860_,
		_w6298_
	);
	LUT4 #(
		.INIT('h5a96)
	) name5836 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w860_,
		_w6299_
	);
	LUT4 #(
		.INIT('h2221)
	) name5837 (
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg2_reg[9]/NET0131 ,
		_w902_,
		_w903_,
		_w6300_
	);
	LUT4 #(
		.INIT('h4448)
	) name5838 (
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg2_reg[9]/NET0131 ,
		_w902_,
		_w903_,
		_w6301_
	);
	LUT2 #(
		.INIT('h1)
	) name5839 (
		_w6232_,
		_w6301_,
		_w6302_
	);
	LUT4 #(
		.INIT('h010f)
	) name5840 (
		_w6233_,
		_w6241_,
		_w6300_,
		_w6302_,
		_w6303_
	);
	LUT4 #(
		.INIT('ha888)
	) name5841 (
		\P1_addr_reg[10]/NET0131 ,
		_w489_,
		_w1236_,
		_w3511_,
		_w6304_
	);
	LUT3 #(
		.INIT('h01)
	) name5842 (
		_w479_,
		_w488_,
		_w892_,
		_w6305_
	);
	LUT2 #(
		.INIT('h1)
	) name5843 (
		_w6304_,
		_w6305_,
		_w6306_
	);
	LUT4 #(
		.INIT('hd700)
	) name5844 (
		_w1245_,
		_w6299_,
		_w6303_,
		_w6306_,
		_w6307_
	);
	LUT4 #(
		.INIT('hbabb)
	) name5845 (
		_w4040_,
		_w6289_,
		_w6296_,
		_w6307_,
		_w6308_
	);
	LUT4 #(
		.INIT('h0509)
	) name5846 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[11]/NET0131 ,
		_w469_,
		_w6309_
	);
	LUT4 #(
		.INIT('ha060)
	) name5847 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[11]/NET0131 ,
		_w469_,
		_w6310_
	);
	LUT4 #(
		.INIT('h5a96)
	) name5848 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[11]/NET0131 ,
		_w469_,
		_w6311_
	);
	LUT2 #(
		.INIT('h1)
	) name5849 (
		_w6232_,
		_w6235_,
		_w6312_
	);
	LUT4 #(
		.INIT('hfe00)
	) name5850 (
		_w6236_,
		_w6237_,
		_w6240_,
		_w6312_,
		_w6313_
	);
	LUT2 #(
		.INIT('h1)
	) name5851 (
		_w6298_,
		_w6300_,
		_w6314_
	);
	LUT3 #(
		.INIT('h4d)
	) name5852 (
		\P1_reg2_reg[10]/NET0131 ,
		_w892_,
		_w6301_,
		_w6315_
	);
	LUT4 #(
		.INIT('hef00)
	) name5853 (
		_w6233_,
		_w6313_,
		_w6314_,
		_w6315_,
		_w6316_
	);
	LUT3 #(
		.INIT('h82)
	) name5854 (
		_w1245_,
		_w6311_,
		_w6316_,
		_w6317_
	);
	LUT4 #(
		.INIT('h0509)
	) name5855 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[11]/NET0131 ,
		_w469_,
		_w6318_
	);
	LUT4 #(
		.INIT('ha060)
	) name5856 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[11]/NET0131 ,
		_w469_,
		_w6319_
	);
	LUT4 #(
		.INIT('h5a96)
	) name5857 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[11]/NET0131 ,
		_w469_,
		_w6320_
	);
	LUT3 #(
		.INIT('h01)
	) name5858 (
		_w6223_,
		_w6291_,
		_w6293_,
		_w6321_
	);
	LUT3 #(
		.INIT('h4d)
	) name5859 (
		\P1_reg1_reg[10]/NET0131 ,
		_w892_,
		_w6294_,
		_w6322_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5860 (
		_w6222_,
		_w6230_,
		_w6321_,
		_w6322_,
		_w6323_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5861 (
		\P1_addr_reg[11]/NET0131 ,
		_w479_,
		_w488_,
		_w882_,
		_w6324_
	);
	LUT4 #(
		.INIT('h7d00)
	) name5862 (
		_w6182_,
		_w6320_,
		_w6323_,
		_w6324_,
		_w6325_
	);
	LUT4 #(
		.INIT('h007f)
	) name5863 (
		\P1_addr_reg[11]/NET0131 ,
		_w1236_,
		_w3511_,
		_w4019_,
		_w6326_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5864 (
		_w6221_,
		_w6317_,
		_w6325_,
		_w6326_,
		_w6327_
	);
	LUT3 #(
		.INIT('h40)
	) name5865 (
		\P1_addr_reg[12]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6328_
	);
	LUT3 #(
		.INIT('h51)
	) name5866 (
		_w1244_,
		_w3511_,
		_w6328_,
		_w6329_
	);
	LUT2 #(
		.INIT('h1)
	) name5867 (
		\P1_reg1_reg[12]/NET0131 ,
		_w862_,
		_w6330_
	);
	LUT2 #(
		.INIT('h6)
	) name5868 (
		\P1_reg1_reg[12]/NET0131 ,
		_w862_,
		_w6331_
	);
	LUT2 #(
		.INIT('h1)
	) name5869 (
		_w6290_,
		_w6319_,
		_w6332_
	);
	LUT4 #(
		.INIT('hfe00)
	) name5870 (
		_w6291_,
		_w6293_,
		_w6295_,
		_w6332_,
		_w6333_
	);
	LUT4 #(
		.INIT('ha082)
	) name5871 (
		_w6182_,
		_w6318_,
		_w6331_,
		_w6333_,
		_w6334_
	);
	LUT2 #(
		.INIT('h1)
	) name5872 (
		\P1_reg2_reg[12]/NET0131 ,
		_w862_,
		_w6335_
	);
	LUT2 #(
		.INIT('h6)
	) name5873 (
		\P1_reg2_reg[12]/NET0131 ,
		_w862_,
		_w6336_
	);
	LUT2 #(
		.INIT('h1)
	) name5874 (
		_w6297_,
		_w6310_,
		_w6337_
	);
	LUT4 #(
		.INIT('h040f)
	) name5875 (
		_w6298_,
		_w6303_,
		_w6309_,
		_w6337_,
		_w6338_
	);
	LUT3 #(
		.INIT('h10)
	) name5876 (
		_w479_,
		_w488_,
		_w862_,
		_w6339_
	);
	LUT4 #(
		.INIT('ha888)
	) name5877 (
		\P1_addr_reg[12]/NET0131 ,
		_w489_,
		_w1236_,
		_w3511_,
		_w6340_
	);
	LUT2 #(
		.INIT('h1)
	) name5878 (
		_w6339_,
		_w6340_,
		_w6341_
	);
	LUT4 #(
		.INIT('hd700)
	) name5879 (
		_w1245_,
		_w6336_,
		_w6338_,
		_w6341_,
		_w6342_
	);
	LUT4 #(
		.INIT('hbabb)
	) name5880 (
		_w3366_,
		_w6329_,
		_w6334_,
		_w6342_,
		_w6343_
	);
	LUT3 #(
		.INIT('h40)
	) name5881 (
		\P1_addr_reg[13]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6344_
	);
	LUT3 #(
		.INIT('h51)
	) name5882 (
		_w1244_,
		_w3511_,
		_w6344_,
		_w6345_
	);
	LUT2 #(
		.INIT('h1)
	) name5883 (
		\P1_reg2_reg[13]/NET0131 ,
		_w850_,
		_w6346_
	);
	LUT2 #(
		.INIT('h6)
	) name5884 (
		\P1_reg2_reg[13]/NET0131 ,
		_w850_,
		_w6347_
	);
	LUT3 #(
		.INIT('h07)
	) name5885 (
		\P1_reg2_reg[12]/NET0131 ,
		_w862_,
		_w6310_,
		_w6348_
	);
	LUT4 #(
		.INIT('h010f)
	) name5886 (
		_w6309_,
		_w6316_,
		_w6335_,
		_w6348_,
		_w6349_
	);
	LUT3 #(
		.INIT('h28)
	) name5887 (
		_w1245_,
		_w6347_,
		_w6349_,
		_w6350_
	);
	LUT3 #(
		.INIT('h07)
	) name5888 (
		\P1_reg1_reg[12]/NET0131 ,
		_w862_,
		_w6319_,
		_w6351_
	);
	LUT4 #(
		.INIT('h010f)
	) name5889 (
		_w6318_,
		_w6323_,
		_w6330_,
		_w6351_,
		_w6352_
	);
	LUT2 #(
		.INIT('h1)
	) name5890 (
		\P1_reg1_reg[13]/NET0131 ,
		_w850_,
		_w6353_
	);
	LUT2 #(
		.INIT('h6)
	) name5891 (
		\P1_reg1_reg[13]/NET0131 ,
		_w850_,
		_w6354_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5892 (
		\P1_addr_reg[13]/NET0131 ,
		_w479_,
		_w488_,
		_w850_,
		_w6355_
	);
	LUT4 #(
		.INIT('hd700)
	) name5893 (
		_w6182_,
		_w6352_,
		_w6354_,
		_w6355_,
		_w6356_
	);
	LUT4 #(
		.INIT('h007f)
	) name5894 (
		\P1_addr_reg[13]/NET0131 ,
		_w1236_,
		_w3511_,
		_w4581_,
		_w6357_
	);
	LUT4 #(
		.INIT('h45ff)
	) name5895 (
		_w6345_,
		_w6350_,
		_w6356_,
		_w6357_,
		_w6358_
	);
	LUT3 #(
		.INIT('h40)
	) name5896 (
		\P1_addr_reg[14]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6359_
	);
	LUT3 #(
		.INIT('h51)
	) name5897 (
		_w1244_,
		_w3511_,
		_w6359_,
		_w6360_
	);
	LUT2 #(
		.INIT('h4)
	) name5898 (
		\P1_reg1_reg[14]/NET0131 ,
		_w840_,
		_w6361_
	);
	LUT2 #(
		.INIT('h9)
	) name5899 (
		\P1_reg1_reg[14]/NET0131 ,
		_w840_,
		_w6362_
	);
	LUT4 #(
		.INIT('h153f)
	) name5900 (
		\P1_reg1_reg[12]/NET0131 ,
		\P1_reg1_reg[13]/NET0131 ,
		_w850_,
		_w862_,
		_w6363_
	);
	LUT4 #(
		.INIT('hfe00)
	) name5901 (
		_w6318_,
		_w6330_,
		_w6333_,
		_w6363_,
		_w6364_
	);
	LUT4 #(
		.INIT('ha082)
	) name5902 (
		_w6182_,
		_w6353_,
		_w6362_,
		_w6364_,
		_w6365_
	);
	LUT2 #(
		.INIT('h4)
	) name5903 (
		\P1_reg2_reg[14]/NET0131 ,
		_w840_,
		_w6366_
	);
	LUT2 #(
		.INIT('h9)
	) name5904 (
		\P1_reg2_reg[14]/NET0131 ,
		_w840_,
		_w6367_
	);
	LUT4 #(
		.INIT('h153f)
	) name5905 (
		\P1_reg2_reg[12]/NET0131 ,
		\P1_reg2_reg[13]/NET0131 ,
		_w850_,
		_w862_,
		_w6368_
	);
	LUT4 #(
		.INIT('h040f)
	) name5906 (
		_w6335_,
		_w6338_,
		_w6346_,
		_w6368_,
		_w6369_
	);
	LUT3 #(
		.INIT('h01)
	) name5907 (
		_w479_,
		_w488_,
		_w840_,
		_w6370_
	);
	LUT4 #(
		.INIT('ha888)
	) name5908 (
		\P1_addr_reg[14]/NET0131 ,
		_w489_,
		_w1236_,
		_w3511_,
		_w6371_
	);
	LUT2 #(
		.INIT('h1)
	) name5909 (
		_w6370_,
		_w6371_,
		_w6372_
	);
	LUT4 #(
		.INIT('hd700)
	) name5910 (
		_w1245_,
		_w6367_,
		_w6369_,
		_w6372_,
		_w6373_
	);
	LUT4 #(
		.INIT('hbabb)
	) name5911 (
		_w4061_,
		_w6360_,
		_w6365_,
		_w6373_,
		_w6374_
	);
	LUT3 #(
		.INIT('h40)
	) name5912 (
		\P1_addr_reg[16]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6375_
	);
	LUT3 #(
		.INIT('h51)
	) name5913 (
		_w1244_,
		_w3511_,
		_w6375_,
		_w6376_
	);
	LUT3 #(
		.INIT('h48)
	) name5914 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_reg1_reg[16]/NET0131 ,
		_w482_,
		_w6377_
	);
	LUT3 #(
		.INIT('h21)
	) name5915 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_reg1_reg[16]/NET0131 ,
		_w482_,
		_w6378_
	);
	LUT3 #(
		.INIT('h96)
	) name5916 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_reg1_reg[16]/NET0131 ,
		_w482_,
		_w6379_
	);
	LUT2 #(
		.INIT('h1)
	) name5917 (
		\P1_reg1_reg[15]/NET0131 ,
		_w831_,
		_w6380_
	);
	LUT2 #(
		.INIT('h8)
	) name5918 (
		\P1_reg1_reg[15]/NET0131 ,
		_w831_,
		_w6381_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5919 (
		\P1_reg1_reg[14]/NET0131 ,
		\P1_reg1_reg[15]/NET0131 ,
		_w831_,
		_w840_,
		_w6382_
	);
	LUT4 #(
		.INIT('hfe00)
	) name5920 (
		_w6353_,
		_w6361_,
		_w6364_,
		_w6382_,
		_w6383_
	);
	LUT4 #(
		.INIT('h8882)
	) name5921 (
		_w6182_,
		_w6379_,
		_w6380_,
		_w6383_,
		_w6384_
	);
	LUT3 #(
		.INIT('h48)
	) name5922 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_reg2_reg[16]/NET0131 ,
		_w482_,
		_w6385_
	);
	LUT3 #(
		.INIT('h21)
	) name5923 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_reg2_reg[16]/NET0131 ,
		_w482_,
		_w6386_
	);
	LUT3 #(
		.INIT('h96)
	) name5924 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_reg2_reg[16]/NET0131 ,
		_w482_,
		_w6387_
	);
	LUT2 #(
		.INIT('h1)
	) name5925 (
		\P1_reg2_reg[15]/NET0131 ,
		_w831_,
		_w6388_
	);
	LUT2 #(
		.INIT('h8)
	) name5926 (
		\P1_reg2_reg[15]/NET0131 ,
		_w831_,
		_w6389_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5927 (
		\P1_reg2_reg[14]/NET0131 ,
		\P1_reg2_reg[15]/NET0131 ,
		_w831_,
		_w840_,
		_w6390_
	);
	LUT4 #(
		.INIT('h040f)
	) name5928 (
		_w6366_,
		_w6369_,
		_w6388_,
		_w6390_,
		_w6391_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5929 (
		\P1_addr_reg[16]/NET0131 ,
		_w479_,
		_w488_,
		_w757_,
		_w6392_
	);
	LUT4 #(
		.INIT('hd700)
	) name5930 (
		_w1245_,
		_w6387_,
		_w6391_,
		_w6392_,
		_w6393_
	);
	LUT4 #(
		.INIT('h070f)
	) name5931 (
		\P1_addr_reg[16]/NET0131 ,
		_w1236_,
		_w2850_,
		_w3511_,
		_w6394_
	);
	LUT4 #(
		.INIT('h45ff)
	) name5932 (
		_w6376_,
		_w6384_,
		_w6393_,
		_w6394_,
		_w6395_
	);
	LUT3 #(
		.INIT('h40)
	) name5933 (
		\P1_addr_reg[17]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6396_
	);
	LUT3 #(
		.INIT('h51)
	) name5934 (
		_w1244_,
		_w3511_,
		_w6396_,
		_w6397_
	);
	LUT3 #(
		.INIT('h48)
	) name5935 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_reg1_reg[17]/NET0131 ,
		_w746_,
		_w6398_
	);
	LUT3 #(
		.INIT('h21)
	) name5936 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_reg1_reg[17]/NET0131 ,
		_w746_,
		_w6399_
	);
	LUT3 #(
		.INIT('h96)
	) name5937 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_reg1_reg[17]/NET0131 ,
		_w746_,
		_w6400_
	);
	LUT4 #(
		.INIT('h51f3)
	) name5938 (
		\P1_reg1_reg[13]/NET0131 ,
		\P1_reg1_reg[14]/NET0131 ,
		_w840_,
		_w850_,
		_w6401_
	);
	LUT4 #(
		.INIT('h020f)
	) name5939 (
		_w6352_,
		_w6353_,
		_w6361_,
		_w6401_,
		_w6402_
	);
	LUT2 #(
		.INIT('h1)
	) name5940 (
		_w6377_,
		_w6381_,
		_w6403_
	);
	LUT4 #(
		.INIT('h1055)
	) name5941 (
		_w6378_,
		_w6380_,
		_w6402_,
		_w6403_,
		_w6404_
	);
	LUT3 #(
		.INIT('h28)
	) name5942 (
		_w6182_,
		_w6400_,
		_w6404_,
		_w6405_
	);
	LUT3 #(
		.INIT('h48)
	) name5943 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_reg2_reg[17]/NET0131 ,
		_w746_,
		_w6406_
	);
	LUT3 #(
		.INIT('h21)
	) name5944 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_reg2_reg[17]/NET0131 ,
		_w746_,
		_w6407_
	);
	LUT3 #(
		.INIT('h96)
	) name5945 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_reg2_reg[17]/NET0131 ,
		_w746_,
		_w6408_
	);
	LUT4 #(
		.INIT('hfca8)
	) name5946 (
		\P1_reg2_reg[12]/NET0131 ,
		\P1_reg2_reg[13]/NET0131 ,
		_w850_,
		_w862_,
		_w6409_
	);
	LUT4 #(
		.INIT('h1f00)
	) name5947 (
		_w6309_,
		_w6316_,
		_w6348_,
		_w6409_,
		_w6410_
	);
	LUT4 #(
		.INIT('h51f3)
	) name5948 (
		\P1_reg2_reg[13]/NET0131 ,
		\P1_reg2_reg[14]/NET0131 ,
		_w840_,
		_w850_,
		_w6411_
	);
	LUT3 #(
		.INIT('h45)
	) name5949 (
		_w6366_,
		_w6410_,
		_w6411_,
		_w6412_
	);
	LUT4 #(
		.INIT('h1011)
	) name5950 (
		_w6366_,
		_w6388_,
		_w6410_,
		_w6411_,
		_w6413_
	);
	LUT2 #(
		.INIT('h1)
	) name5951 (
		_w6385_,
		_w6389_,
		_w6414_
	);
	LUT3 #(
		.INIT('h45)
	) name5952 (
		_w6386_,
		_w6413_,
		_w6414_,
		_w6415_
	);
	LUT3 #(
		.INIT('h10)
	) name5953 (
		_w479_,
		_w488_,
		_w747_,
		_w6416_
	);
	LUT4 #(
		.INIT('ha888)
	) name5954 (
		\P1_addr_reg[17]/NET0131 ,
		_w489_,
		_w1236_,
		_w3511_,
		_w6417_
	);
	LUT2 #(
		.INIT('h1)
	) name5955 (
		_w6416_,
		_w6417_,
		_w6418_
	);
	LUT4 #(
		.INIT('hd700)
	) name5956 (
		_w1245_,
		_w6408_,
		_w6415_,
		_w6418_,
		_w6419_
	);
	LUT4 #(
		.INIT('hbabb)
	) name5957 (
		_w3666_,
		_w6397_,
		_w6405_,
		_w6419_,
		_w6420_
	);
	LUT3 #(
		.INIT('h40)
	) name5958 (
		\P1_addr_reg[18]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6421_
	);
	LUT3 #(
		.INIT('h51)
	) name5959 (
		_w1244_,
		_w3511_,
		_w6421_,
		_w6422_
	);
	LUT4 #(
		.INIT('h4448)
	) name5960 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_reg1_reg[18]/NET0131 ,
		_w482_,
		_w731_,
		_w6423_
	);
	LUT4 #(
		.INIT('h2221)
	) name5961 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_reg1_reg[18]/NET0131 ,
		_w482_,
		_w731_,
		_w6424_
	);
	LUT4 #(
		.INIT('h9996)
	) name5962 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_reg1_reg[18]/NET0131 ,
		_w482_,
		_w731_,
		_w6425_
	);
	LUT2 #(
		.INIT('h1)
	) name5963 (
		_w6378_,
		_w6399_,
		_w6426_
	);
	LUT3 #(
		.INIT('h17)
	) name5964 (
		\P1_reg1_reg[17]/NET0131 ,
		_w747_,
		_w6377_,
		_w6427_
	);
	LUT4 #(
		.INIT('hef00)
	) name5965 (
		_w6380_,
		_w6383_,
		_w6426_,
		_w6427_,
		_w6428_
	);
	LUT3 #(
		.INIT('h82)
	) name5966 (
		_w6182_,
		_w6425_,
		_w6428_,
		_w6429_
	);
	LUT4 #(
		.INIT('h4448)
	) name5967 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_reg2_reg[18]/NET0131 ,
		_w482_,
		_w731_,
		_w6430_
	);
	LUT4 #(
		.INIT('h2221)
	) name5968 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_reg2_reg[18]/NET0131 ,
		_w482_,
		_w731_,
		_w6431_
	);
	LUT4 #(
		.INIT('h9996)
	) name5969 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_reg2_reg[18]/NET0131 ,
		_w482_,
		_w731_,
		_w6432_
	);
	LUT2 #(
		.INIT('h1)
	) name5970 (
		_w6386_,
		_w6407_,
		_w6433_
	);
	LUT3 #(
		.INIT('h17)
	) name5971 (
		\P1_reg2_reg[17]/NET0131 ,
		_w747_,
		_w6385_,
		_w6434_
	);
	LUT3 #(
		.INIT('h70)
	) name5972 (
		_w6391_,
		_w6433_,
		_w6434_,
		_w6435_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5973 (
		\P1_addr_reg[18]/NET0131 ,
		_w479_,
		_w488_,
		_w732_,
		_w6436_
	);
	LUT4 #(
		.INIT('h7d00)
	) name5974 (
		_w1245_,
		_w6432_,
		_w6435_,
		_w6436_,
		_w6437_
	);
	LUT4 #(
		.INIT('h070f)
	) name5975 (
		\P1_addr_reg[18]/NET0131 ,
		_w1236_,
		_w3389_,
		_w3511_,
		_w6438_
	);
	LUT4 #(
		.INIT('h45ff)
	) name5976 (
		_w6422_,
		_w6429_,
		_w6437_,
		_w6438_,
		_w6439_
	);
	LUT3 #(
		.INIT('h40)
	) name5977 (
		\P1_addr_reg[19]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6440_
	);
	LUT3 #(
		.INIT('h51)
	) name5978 (
		_w1244_,
		_w3511_,
		_w6440_,
		_w6441_
	);
	LUT2 #(
		.INIT('h1)
	) name5979 (
		_w6399_,
		_w6424_,
		_w6442_
	);
	LUT4 #(
		.INIT('h010f)
	) name5980 (
		_w6398_,
		_w6404_,
		_w6423_,
		_w6442_,
		_w6443_
	);
	LUT2 #(
		.INIT('h6)
	) name5981 (
		\P1_reg1_reg[19]/NET0131 ,
		_w718_,
		_w6444_
	);
	LUT3 #(
		.INIT('h28)
	) name5982 (
		_w6182_,
		_w6443_,
		_w6444_,
		_w6445_
	);
	LUT4 #(
		.INIT('h2322)
	) name5983 (
		_w6386_,
		_w6406_,
		_w6413_,
		_w6414_,
		_w6446_
	);
	LUT2 #(
		.INIT('h1)
	) name5984 (
		_w6407_,
		_w6431_,
		_w6447_
	);
	LUT3 #(
		.INIT('h45)
	) name5985 (
		_w6430_,
		_w6446_,
		_w6447_,
		_w6448_
	);
	LUT2 #(
		.INIT('h6)
	) name5986 (
		\P1_reg2_reg[19]/NET0131 ,
		_w718_,
		_w6449_
	);
	LUT4 #(
		.INIT('hff5c)
	) name5987 (
		\P1_addr_reg[19]/NET0131 ,
		_w718_,
		_w479_,
		_w488_,
		_w6450_
	);
	LUT4 #(
		.INIT('hd700)
	) name5988 (
		_w1245_,
		_w6448_,
		_w6449_,
		_w6450_,
		_w6451_
	);
	LUT4 #(
		.INIT('h007f)
	) name5989 (
		\P1_addr_reg[19]/NET0131 ,
		_w1236_,
		_w3511_,
		_w3688_,
		_w6452_
	);
	LUT4 #(
		.INIT('h45ff)
	) name5990 (
		_w6441_,
		_w6445_,
		_w6451_,
		_w6452_,
		_w6453_
	);
	LUT3 #(
		.INIT('h40)
	) name5991 (
		\P1_addr_reg[15]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6454_
	);
	LUT3 #(
		.INIT('h51)
	) name5992 (
		_w1244_,
		_w3511_,
		_w6454_,
		_w6455_
	);
	LUT2 #(
		.INIT('h6)
	) name5993 (
		\P1_reg1_reg[15]/NET0131 ,
		_w831_,
		_w6456_
	);
	LUT3 #(
		.INIT('h28)
	) name5994 (
		_w6182_,
		_w6402_,
		_w6456_,
		_w6457_
	);
	LUT2 #(
		.INIT('h6)
	) name5995 (
		\P1_reg2_reg[15]/NET0131 ,
		_w831_,
		_w6458_
	);
	LUT3 #(
		.INIT('h10)
	) name5996 (
		_w479_,
		_w488_,
		_w831_,
		_w6459_
	);
	LUT4 #(
		.INIT('ha888)
	) name5997 (
		\P1_addr_reg[15]/NET0131 ,
		_w489_,
		_w1236_,
		_w3511_,
		_w6460_
	);
	LUT2 #(
		.INIT('h1)
	) name5998 (
		_w6459_,
		_w6460_,
		_w6461_
	);
	LUT4 #(
		.INIT('hd700)
	) name5999 (
		_w1245_,
		_w6412_,
		_w6458_,
		_w6461_,
		_w6462_
	);
	LUT4 #(
		.INIT('hbabb)
	) name6000 (
		_w4082_,
		_w6455_,
		_w6457_,
		_w6462_,
		_w6463_
	);
	LUT2 #(
		.INIT('h2)
	) name6001 (
		\P1_reg3_reg[1]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6464_
	);
	LUT3 #(
		.INIT('h40)
	) name6002 (
		\P1_addr_reg[1]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6465_
	);
	LUT3 #(
		.INIT('h51)
	) name6003 (
		_w1244_,
		_w3511_,
		_w6465_,
		_w6466_
	);
	LUT4 #(
		.INIT('ha888)
	) name6004 (
		\P1_addr_reg[1]/NET0131 ,
		_w489_,
		_w1236_,
		_w3511_,
		_w6467_
	);
	LUT4 #(
		.INIT('h936c)
	) name6005 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[1]/NET0131 ,
		_w6468_
	);
	LUT2 #(
		.INIT('h6)
	) name6006 (
		_w6180_,
		_w6468_,
		_w6469_
	);
	LUT3 #(
		.INIT('h40)
	) name6007 (
		_w479_,
		_w488_,
		_w6469_,
		_w6470_
	);
	LUT4 #(
		.INIT('h936c)
	) name6008 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[1]/NET0131 ,
		_w6471_
	);
	LUT2 #(
		.INIT('h6)
	) name6009 (
		_w6183_,
		_w6471_,
		_w6472_
	);
	LUT4 #(
		.INIT('h76fe)
	) name6010 (
		_w479_,
		_w488_,
		_w991_,
		_w6472_,
		_w6473_
	);
	LUT2 #(
		.INIT('h4)
	) name6011 (
		_w6470_,
		_w6473_,
		_w6474_
	);
	LUT4 #(
		.INIT('hbabb)
	) name6012 (
		_w6464_,
		_w6466_,
		_w6467_,
		_w6474_,
		_w6475_
	);
	LUT2 #(
		.INIT('h9)
	) name6013 (
		\P1_reg1_reg[5]/NET0131 ,
		_w955_,
		_w6476_
	);
	LUT4 #(
		.INIT('h0880)
	) name6014 (
		_w479_,
		_w488_,
		_w6227_,
		_w6476_,
		_w6477_
	);
	LUT3 #(
		.INIT('h01)
	) name6015 (
		_w479_,
		_w488_,
		_w955_,
		_w6478_
	);
	LUT2 #(
		.INIT('h9)
	) name6016 (
		\P1_reg2_reg[5]/NET0131 ,
		_w955_,
		_w6479_
	);
	LUT4 #(
		.INIT('h0440)
	) name6017 (
		_w479_,
		_w488_,
		_w6239_,
		_w6479_,
		_w6480_
	);
	LUT3 #(
		.INIT('h01)
	) name6018 (
		_w6478_,
		_w6480_,
		_w6477_,
		_w6481_
	);
	LUT2 #(
		.INIT('h2)
	) name6019 (
		_w6221_,
		_w6481_,
		_w6482_
	);
	LUT2 #(
		.INIT('h8)
	) name6020 (
		\P1_addr_reg[5]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6483_
	);
	LUT2 #(
		.INIT('h4)
	) name6021 (
		_w2183_,
		_w6483_,
		_w6484_
	);
	LUT3 #(
		.INIT('h45)
	) name6022 (
		_w4675_,
		_w6271_,
		_w6484_,
		_w6485_
	);
	LUT2 #(
		.INIT('hb)
	) name6023 (
		_w6482_,
		_w6485_,
		_w6486_
	);
	LUT3 #(
		.INIT('h40)
	) name6024 (
		\P1_addr_reg[9]/NET0131 ,
		_w1096_,
		_w1098_,
		_w6487_
	);
	LUT3 #(
		.INIT('h51)
	) name6025 (
		_w1244_,
		_w3511_,
		_w6487_,
		_w6488_
	);
	LUT4 #(
		.INIT('h9996)
	) name6026 (
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg1_reg[9]/NET0131 ,
		_w902_,
		_w903_,
		_w6489_
	);
	LUT4 #(
		.INIT('h00d4)
	) name6027 (
		\P1_reg1_reg[8]/NET0131 ,
		_w914_,
		_w6230_,
		_w6489_,
		_w6490_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6028 (
		\P1_reg1_reg[8]/NET0131 ,
		_w914_,
		_w6230_,
		_w6489_,
		_w6491_
	);
	LUT3 #(
		.INIT('h02)
	) name6029 (
		_w6182_,
		_w6491_,
		_w6490_,
		_w6492_
	);
	LUT4 #(
		.INIT('h9996)
	) name6030 (
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg2_reg[9]/NET0131 ,
		_w902_,
		_w903_,
		_w6493_
	);
	LUT4 #(
		.INIT('ha802)
	) name6031 (
		_w1245_,
		_w6233_,
		_w6313_,
		_w6493_,
		_w6494_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name6032 (
		\P1_addr_reg[9]/NET0131 ,
		_w479_,
		_w488_,
		_w904_,
		_w6495_
	);
	LUT2 #(
		.INIT('h4)
	) name6033 (
		_w6494_,
		_w6495_,
		_w6496_
	);
	LUT4 #(
		.INIT('h007f)
	) name6034 (
		\P1_addr_reg[9]/NET0131 ,
		_w1236_,
		_w3511_,
		_w3745_,
		_w6497_
	);
	LUT4 #(
		.INIT('h45ff)
	) name6035 (
		_w6488_,
		_w6492_,
		_w6496_,
		_w6497_,
		_w6498_
	);
	LUT4 #(
		.INIT('h2000)
	) name6036 (
		\P1_state_reg[0]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w6499_
	);
	LUT2 #(
		.INIT('h8)
	) name6037 (
		\P1_state_reg[0]/NET0131 ,
		_w2183_,
		_w6500_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6038 (
		_w1537_,
		_w1963_,
		_w2903_,
		_w3218_,
		_w6501_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6039 (
		_w1537_,
		_w1869_,
		_w2903_,
		_w3214_,
		_w6502_
	);
	LUT4 #(
		.INIT('haa20)
	) name6040 (
		_w2903_,
		_w3221_,
		_w3222_,
		_w3223_,
		_w6503_
	);
	LUT3 #(
		.INIT('h90)
	) name6041 (
		_w1863_,
		_w1866_,
		_w1999_,
		_w6504_
	);
	LUT4 #(
		.INIT('h3031)
	) name6042 (
		_w2001_,
		_w2032_,
		_w2903_,
		_w6504_,
		_w6505_
	);
	LUT4 #(
		.INIT('hf531)
	) name6043 (
		_w1534_,
		_w1537_,
		_w2993_,
		_w6505_,
		_w6506_
	);
	LUT2 #(
		.INIT('h4)
	) name6044 (
		_w6503_,
		_w6506_,
		_w6507_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6045 (
		_w2556_,
		_w6502_,
		_w6501_,
		_w6507_,
		_w6508_
	);
	LUT2 #(
		.INIT('h4)
	) name6046 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[24]/NET0131 ,
		_w6509_
	);
	LUT4 #(
		.INIT('ha888)
	) name6047 (
		\P1_state_reg[0]/NET0131 ,
		_w1267_,
		_w1275_,
		_w1283_,
		_w6510_
	);
	LUT4 #(
		.INIT('h3200)
	) name6048 (
		\P2_reg3_reg[24]/NET0131 ,
		_w1394_,
		_w1536_,
		_w6510_,
		_w6511_
	);
	LUT2 #(
		.INIT('h1)
	) name6049 (
		_w6509_,
		_w6511_,
		_w6512_
	);
	LUT2 #(
		.INIT('hb)
	) name6050 (
		_w6508_,
		_w6512_,
		_w6513_
	);
	LUT2 #(
		.INIT('h2)
	) name6051 (
		_w1507_,
		_w2903_,
		_w6514_
	);
	LUT4 #(
		.INIT('h007b)
	) name6052 (
		_w2514_,
		_w2903_,
		_w3107_,
		_w6514_,
		_w6515_
	);
	LUT2 #(
		.INIT('h2)
	) name6053 (
		_w1869_,
		_w6515_,
		_w6516_
	);
	LUT4 #(
		.INIT('h00b7)
	) name6054 (
		_w2514_,
		_w2903_,
		_w3123_,
		_w6514_,
		_w6517_
	);
	LUT4 #(
		.INIT('h7020)
	) name6055 (
		_w1305_,
		_w1527_,
		_w2903_,
		_w3125_,
		_w6518_
	);
	LUT4 #(
		.INIT('h8400)
	) name6056 (
		_w1506_,
		_w2025_,
		_w2632_,
		_w2903_,
		_w6519_
	);
	LUT4 #(
		.INIT('h88a8)
	) name6057 (
		_w1507_,
		_w2032_,
		_w2033_,
		_w2903_,
		_w6520_
	);
	LUT4 #(
		.INIT('h00fe)
	) name6058 (
		_w1306_,
		_w1505_,
		_w2993_,
		_w6520_,
		_w6521_
	);
	LUT2 #(
		.INIT('h4)
	) name6059 (
		_w6519_,
		_w6521_,
		_w6522_
	);
	LUT4 #(
		.INIT('h5700)
	) name6060 (
		_w2000_,
		_w6514_,
		_w6518_,
		_w6522_,
		_w6523_
	);
	LUT3 #(
		.INIT('hd0)
	) name6061 (
		_w1963_,
		_w6517_,
		_w6523_,
		_w6524_
	);
	LUT2 #(
		.INIT('h4)
	) name6062 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		_w6525_
	);
	LUT3 #(
		.INIT('h07)
	) name6063 (
		_w1507_,
		_w6510_,
		_w6525_,
		_w6526_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6064 (
		_w2556_,
		_w6516_,
		_w6524_,
		_w6526_,
		_w6527_
	);
	LUT3 #(
		.INIT('h28)
	) name6065 (
		_w1963_,
		_w2507_,
		_w3495_,
		_w6528_
	);
	LUT2 #(
		.INIT('h2)
	) name6066 (
		\P2_reg2_reg[22]/NET0131 ,
		_w1298_,
		_w6529_
	);
	LUT2 #(
		.INIT('h8)
	) name6067 (
		_w1561_,
		_w2029_,
		_w6530_
	);
	LUT4 #(
		.INIT('h00df)
	) name6068 (
		\P2_reg2_reg[22]/NET0131 ,
		_w1298_,
		_w2033_,
		_w6530_,
		_w6531_
	);
	LUT4 #(
		.INIT('h5d00)
	) name6069 (
		_w1298_,
		_w3505_,
		_w6528_,
		_w6531_,
		_w6532_
	);
	LUT2 #(
		.INIT('h8)
	) name6070 (
		_w1298_,
		_w2556_,
		_w6533_
	);
	LUT4 #(
		.INIT('h060f)
	) name6071 (
		_w2507_,
		_w3488_,
		_w6529_,
		_w6533_,
		_w6534_
	);
	LUT2 #(
		.INIT('h4)
	) name6072 (
		_w2032_,
		_w2556_,
		_w6535_
	);
	LUT4 #(
		.INIT('hab00)
	) name6073 (
		_w1298_,
		_w1963_,
		_w2000_,
		_w6535_,
		_w6536_
	);
	LUT2 #(
		.INIT('h2)
	) name6074 (
		\P2_reg2_reg[22]/NET0131 ,
		_w6536_,
		_w6537_
	);
	LUT3 #(
		.INIT('h0d)
	) name6075 (
		_w1869_,
		_w6534_,
		_w6537_,
		_w6538_
	);
	LUT3 #(
		.INIT('h2f)
	) name6076 (
		_w2556_,
		_w6532_,
		_w6538_,
		_w6539_
	);
	LUT2 #(
		.INIT('h9)
	) name6077 (
		\P1_rd_reg/NET0131 ,
		\P2_rd_reg/NET0131 ,
		_w6540_
	);
	LUT2 #(
		.INIT('h6)
	) name6078 (
		\P1_addr_reg[0]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		_w6541_
	);
	LUT2 #(
		.INIT('h6)
	) name6079 (
		\P1_addr_reg[10]/NET0131 ,
		\P2_addr_reg[10]/NET0131 ,
		_w6542_
	);
	LUT2 #(
		.INIT('h1)
	) name6080 (
		\P1_addr_reg[9]/NET0131 ,
		\P2_addr_reg[9]/NET0131 ,
		_w6543_
	);
	LUT2 #(
		.INIT('h8)
	) name6081 (
		\P1_addr_reg[9]/NET0131 ,
		\P2_addr_reg[9]/NET0131 ,
		_w6544_
	);
	LUT2 #(
		.INIT('h1)
	) name6082 (
		\P1_addr_reg[6]/NET0131 ,
		\P2_addr_reg[6]/NET0131 ,
		_w6545_
	);
	LUT2 #(
		.INIT('h8)
	) name6083 (
		\P1_addr_reg[6]/NET0131 ,
		\P2_addr_reg[6]/NET0131 ,
		_w6546_
	);
	LUT2 #(
		.INIT('h1)
	) name6084 (
		\P1_addr_reg[3]/NET0131 ,
		\P2_addr_reg[3]/NET0131 ,
		_w6547_
	);
	LUT2 #(
		.INIT('h8)
	) name6085 (
		\P1_addr_reg[3]/NET0131 ,
		\P2_addr_reg[3]/NET0131 ,
		_w6548_
	);
	LUT4 #(
		.INIT('hec80)
	) name6086 (
		\P1_addr_reg[0]/NET0131 ,
		\P1_addr_reg[1]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		\P2_addr_reg[1]/NET0131 ,
		_w6549_
	);
	LUT4 #(
		.INIT('h0107)
	) name6087 (
		\P1_addr_reg[2]/NET0131 ,
		\P2_addr_reg[2]/NET0131 ,
		_w6548_,
		_w6549_,
		_w6550_
	);
	LUT4 #(
		.INIT('h888e)
	) name6088 (
		\P1_addr_reg[4]/NET0131 ,
		\P2_addr_reg[4]/NET0131 ,
		_w6547_,
		_w6550_,
		_w6551_
	);
	LUT4 #(
		.INIT('h0107)
	) name6089 (
		\P1_addr_reg[5]/NET0131 ,
		\P2_addr_reg[5]/NET0131 ,
		_w6546_,
		_w6551_,
		_w6552_
	);
	LUT4 #(
		.INIT('h888e)
	) name6090 (
		\P1_addr_reg[7]/NET0131 ,
		\P2_addr_reg[7]/NET0131 ,
		_w6545_,
		_w6552_,
		_w6553_
	);
	LUT4 #(
		.INIT('h0107)
	) name6091 (
		\P1_addr_reg[8]/NET0131 ,
		\P2_addr_reg[8]/NET0131 ,
		_w6544_,
		_w6553_,
		_w6554_
	);
	LUT3 #(
		.INIT('ha9)
	) name6092 (
		_w6542_,
		_w6543_,
		_w6554_,
		_w6555_
	);
	LUT2 #(
		.INIT('h6)
	) name6093 (
		\P1_addr_reg[11]/NET0131 ,
		\P2_addr_reg[11]/NET0131 ,
		_w6556_
	);
	LUT4 #(
		.INIT('h888e)
	) name6094 (
		\P1_addr_reg[10]/NET0131 ,
		\P2_addr_reg[10]/NET0131 ,
		_w6543_,
		_w6554_,
		_w6557_
	);
	LUT2 #(
		.INIT('h6)
	) name6095 (
		_w6556_,
		_w6557_,
		_w6558_
	);
	LUT2 #(
		.INIT('h8)
	) name6096 (
		\P1_addr_reg[12]/NET0131 ,
		\P2_addr_reg[12]/NET0131 ,
		_w6559_
	);
	LUT2 #(
		.INIT('h1)
	) name6097 (
		\P1_addr_reg[12]/NET0131 ,
		\P2_addr_reg[12]/NET0131 ,
		_w6560_
	);
	LUT2 #(
		.INIT('h6)
	) name6098 (
		\P1_addr_reg[12]/NET0131 ,
		\P2_addr_reg[12]/NET0131 ,
		_w6561_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6099 (
		\P1_addr_reg[11]/NET0131 ,
		\P2_addr_reg[11]/NET0131 ,
		_w6557_,
		_w6561_,
		_w6562_
	);
	LUT2 #(
		.INIT('h6)
	) name6100 (
		\P1_addr_reg[13]/NET0131 ,
		\P2_addr_reg[13]/NET0131 ,
		_w6563_
	);
	LUT4 #(
		.INIT('h0017)
	) name6101 (
		\P1_addr_reg[11]/NET0131 ,
		\P2_addr_reg[11]/NET0131 ,
		_w6557_,
		_w6559_,
		_w6564_
	);
	LUT3 #(
		.INIT('hc9)
	) name6102 (
		_w6560_,
		_w6563_,
		_w6564_,
		_w6565_
	);
	LUT2 #(
		.INIT('h6)
	) name6103 (
		\P1_addr_reg[14]/NET0131 ,
		\P2_addr_reg[14]/NET0131 ,
		_w6566_
	);
	LUT4 #(
		.INIT('h888e)
	) name6104 (
		\P1_addr_reg[13]/NET0131 ,
		\P2_addr_reg[13]/NET0131 ,
		_w6560_,
		_w6564_,
		_w6567_
	);
	LUT2 #(
		.INIT('h6)
	) name6105 (
		_w6566_,
		_w6567_,
		_w6568_
	);
	LUT2 #(
		.INIT('h8)
	) name6106 (
		\P1_addr_reg[15]/NET0131 ,
		\P2_addr_reg[15]/NET0131 ,
		_w6569_
	);
	LUT2 #(
		.INIT('h1)
	) name6107 (
		\P1_addr_reg[15]/NET0131 ,
		\P2_addr_reg[15]/NET0131 ,
		_w6570_
	);
	LUT2 #(
		.INIT('h6)
	) name6108 (
		\P1_addr_reg[15]/NET0131 ,
		\P2_addr_reg[15]/NET0131 ,
		_w6571_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6109 (
		\P1_addr_reg[14]/NET0131 ,
		\P2_addr_reg[14]/NET0131 ,
		_w6567_,
		_w6571_,
		_w6572_
	);
	LUT2 #(
		.INIT('h6)
	) name6110 (
		\P1_addr_reg[16]/NET0131 ,
		\P2_addr_reg[16]/NET0131 ,
		_w6573_
	);
	LUT4 #(
		.INIT('h0017)
	) name6111 (
		\P1_addr_reg[14]/NET0131 ,
		\P2_addr_reg[14]/NET0131 ,
		_w6567_,
		_w6569_,
		_w6574_
	);
	LUT3 #(
		.INIT('hc9)
	) name6112 (
		_w6570_,
		_w6573_,
		_w6574_,
		_w6575_
	);
	LUT2 #(
		.INIT('h6)
	) name6113 (
		\P1_addr_reg[17]/NET0131 ,
		\P2_addr_reg[17]/NET0131 ,
		_w6576_
	);
	LUT4 #(
		.INIT('h888e)
	) name6114 (
		\P1_addr_reg[16]/NET0131 ,
		\P2_addr_reg[16]/NET0131 ,
		_w6570_,
		_w6574_,
		_w6577_
	);
	LUT2 #(
		.INIT('h6)
	) name6115 (
		_w6576_,
		_w6577_,
		_w6578_
	);
	LUT2 #(
		.INIT('h8)
	) name6116 (
		\P1_addr_reg[18]/NET0131 ,
		\P2_addr_reg[18]/NET0131 ,
		_w6579_
	);
	LUT2 #(
		.INIT('h1)
	) name6117 (
		\P1_addr_reg[18]/NET0131 ,
		\P2_addr_reg[18]/NET0131 ,
		_w6580_
	);
	LUT2 #(
		.INIT('h6)
	) name6118 (
		\P1_addr_reg[18]/NET0131 ,
		\P2_addr_reg[18]/NET0131 ,
		_w6581_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6119 (
		\P1_addr_reg[17]/NET0131 ,
		\P2_addr_reg[17]/NET0131 ,
		_w6577_,
		_w6581_,
		_w6582_
	);
	LUT2 #(
		.INIT('h6)
	) name6120 (
		\P1_addr_reg[19]/NET0131 ,
		\P2_addr_reg[19]/NET0131 ,
		_w6583_
	);
	LUT4 #(
		.INIT('h0017)
	) name6121 (
		\P1_addr_reg[17]/NET0131 ,
		\P2_addr_reg[17]/NET0131 ,
		_w6577_,
		_w6579_,
		_w6584_
	);
	LUT3 #(
		.INIT('hc9)
	) name6122 (
		_w6580_,
		_w6583_,
		_w6584_,
		_w6585_
	);
	LUT4 #(
		.INIT('h936c)
	) name6123 (
		\P1_addr_reg[0]/NET0131 ,
		\P1_addr_reg[1]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		\P2_addr_reg[1]/NET0131 ,
		_w6586_
	);
	LUT2 #(
		.INIT('h6)
	) name6124 (
		\P1_addr_reg[2]/NET0131 ,
		\P2_addr_reg[2]/NET0131 ,
		_w6587_
	);
	LUT2 #(
		.INIT('h6)
	) name6125 (
		_w6549_,
		_w6587_,
		_w6588_
	);
	LUT2 #(
		.INIT('h6)
	) name6126 (
		\P1_addr_reg[3]/NET0131 ,
		\P2_addr_reg[3]/NET0131 ,
		_w6589_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6127 (
		\P1_addr_reg[2]/NET0131 ,
		\P2_addr_reg[2]/NET0131 ,
		_w6549_,
		_w6589_,
		_w6590_
	);
	LUT2 #(
		.INIT('h6)
	) name6128 (
		\P1_addr_reg[4]/NET0131 ,
		\P2_addr_reg[4]/NET0131 ,
		_w6591_
	);
	LUT3 #(
		.INIT('he1)
	) name6129 (
		_w6547_,
		_w6550_,
		_w6591_,
		_w6592_
	);
	LUT2 #(
		.INIT('h6)
	) name6130 (
		\P1_addr_reg[5]/NET0131 ,
		\P2_addr_reg[5]/NET0131 ,
		_w6593_
	);
	LUT2 #(
		.INIT('h6)
	) name6131 (
		_w6551_,
		_w6593_,
		_w6594_
	);
	LUT2 #(
		.INIT('h6)
	) name6132 (
		\P1_addr_reg[6]/NET0131 ,
		\P2_addr_reg[6]/NET0131 ,
		_w6595_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6133 (
		\P1_addr_reg[5]/NET0131 ,
		\P2_addr_reg[5]/NET0131 ,
		_w6551_,
		_w6595_,
		_w6596_
	);
	LUT2 #(
		.INIT('h6)
	) name6134 (
		\P1_addr_reg[7]/NET0131 ,
		\P2_addr_reg[7]/NET0131 ,
		_w6597_
	);
	LUT3 #(
		.INIT('he1)
	) name6135 (
		_w6545_,
		_w6552_,
		_w6597_,
		_w6598_
	);
	LUT2 #(
		.INIT('h6)
	) name6136 (
		\P1_addr_reg[8]/NET0131 ,
		\P2_addr_reg[8]/NET0131 ,
		_w6599_
	);
	LUT2 #(
		.INIT('h6)
	) name6137 (
		_w6553_,
		_w6599_,
		_w6600_
	);
	LUT2 #(
		.INIT('h6)
	) name6138 (
		\P1_addr_reg[9]/NET0131 ,
		\P2_addr_reg[9]/NET0131 ,
		_w6601_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6139 (
		\P1_addr_reg[8]/NET0131 ,
		\P2_addr_reg[8]/NET0131 ,
		_w6553_,
		_w6601_,
		_w6602_
	);
	LUT2 #(
		.INIT('h9)
	) name6140 (
		\P1_wr_reg/NET0131 ,
		\P2_wr_reg/NET0131 ,
		_w6603_
	);
	assign \P1_state_reg[0]/NET0131_syn_2  = _w216_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g70791/_0_  = _w1255_ ;
	assign \g70792/_0_  = _w2044_ ;
	assign \g70793/_0_  = _w2188_ ;
	assign \g70794/_0_  = _w2207_ ;
	assign \g70795/_0_  = _w2322_ ;
	assign \g70796/_0_  = _w2339_ ;
	assign \g70813/_0_  = _w2533_ ;
	assign \g70814/_0_  = _w2550_ ;
	assign \g70848/_0_  = _w2559_ ;
	assign \g70849/_0_  = _w2588_ ;
	assign \g70850/_0_  = _w2646_ ;
	assign \g70851/_0_  = _w2699_ ;
	assign \g70852/_0_  = _w2728_ ;
	assign \g70856/_0_  = _w2743_ ;
	assign \g70857/_0_  = _w2761_ ;
	assign \g70858/_0_  = _w2776_ ;
	assign \g70859/_0_  = _w2790_ ;
	assign \g70860/_0_  = _w2806_ ;
	assign \g70861/_0_  = _w2824_ ;
	assign \g70862/_0_  = _w2833_ ;
	assign \g70896/_0_  = _w2852_ ;
	assign \g70902/_0_  = _w2872_ ;
	assign \g70903/_0_  = _w2901_ ;
	assign \g70904/_0_  = _w2916_ ;
	assign \g70906/_0_  = _w2933_ ;
	assign \g70907/_0_  = _w2985_ ;
	assign \g70908/_0_  = _w3001_ ;
	assign \g70909/_0_  = _w3067_ ;
	assign \g70910/_0_  = _w3077_ ;
	assign \g70911/_0_  = _w3091_ ;
	assign \g70912/_0_  = _w3135_ ;
	assign \g70913/_0_  = _w3152_ ;
	assign \g70914/_0_  = _w3157_ ;
	assign \g70915/_0_  = _w3180_ ;
	assign \g70916/_0_  = _w3192_ ;
	assign \g70917/_0_  = _w3209_ ;
	assign \g70918/_0_  = _w3230_ ;
	assign \g70919/_0_  = _w3240_ ;
	assign \g70920/_0_  = _w3248_ ;
	assign \g70921/_0_  = _w3265_ ;
	assign \g70922/_0_  = _w3269_ ;
	assign \g70923/_0_  = _w3288_ ;
	assign \g70924/_0_  = _w3299_ ;
	assign \g70925/_0_  = _w3315_ ;
	assign \g70926/_0_  = _w3330_ ;
	assign \g70927/_0_  = _w3346_ ;
	assign \g70987/_0_  = _w3369_ ;
	assign \g70988/_0_  = _w3391_ ;
	assign \g70989/_0_  = _w3414_ ;
	assign \g70990/_0_  = _w3432_ ;
	assign \g70991/_0_  = _w3449_ ;
	assign \g71006/_0_  = _w3469_ ;
	assign \g71007/_0_  = _w3485_ ;
	assign \g71009/_0_  = _w3510_ ;
	assign \g71010/_0_  = _w3520_ ;
	assign \g71011/_0_  = _w3528_ ;
	assign \g71012/_0_  = _w3539_ ;
	assign \g71013/_0_  = _w3548_ ;
	assign \g71014/_0_  = _w3559_ ;
	assign \g71015/_0_  = _w3564_ ;
	assign \g71016/_0_  = _w3584_ ;
	assign \g71017/_0_  = _w3600_ ;
	assign \g71018/_0_  = _w3604_ ;
	assign \g71019/_0_  = _w3609_ ;
	assign \g71020/_0_  = _w3620_ ;
	assign \g71021/_0_  = _w3632_ ;
	assign \g71022/_0_  = _w3648_ ;
	assign \g71023/_0_  = _w3651_ ;
	assign \g71090/_0_  = _w3668_ ;
	assign \g71091/_0_  = _w3690_ ;
	assign \g71092/_0_  = _w3708_ ;
	assign \g71093/_0_  = _w3729_ ;
	assign \g71094/_0_  = _w3748_ ;
	assign \g71125/_0_  = _w3765_ ;
	assign \g71130/_0_  = _w3776_ ;
	assign \g71131/_0_  = _w3800_ ;
	assign \g71132/_0_  = _w3817_ ;
	assign \g71133/_0_  = _w3822_ ;
	assign \g71134/_0_  = _w3839_ ;
	assign \g71135/_0_  = _w3851_ ;
	assign \g71136/_0_  = _w3865_ ;
	assign \g71137/_0_  = _w3877_ ;
	assign \g71138/_0_  = _w3890_ ;
	assign \g71139/_0_  = _w3896_ ;
	assign \g71140/_0_  = _w3906_ ;
	assign \g71141/_0_  = _w3909_ ;
	assign \g71142/_0_  = _w3916_ ;
	assign \g71143/_0_  = _w3924_ ;
	assign \g71144/_0_  = _w3929_ ;
	assign \g71145/_0_  = _w3950_ ;
	assign \g71150/_0_  = _w3958_ ;
	assign \g71151/_0_  = _w3966_ ;
	assign \g71152/_0_  = _w3969_ ;
	assign \g71153/_0_  = _w3972_ ;
	assign \g71154/_0_  = _w3980_ ;
	assign \g71155/_0_  = _w3986_ ;
	assign \g71156/_0_  = _w3996_ ;
	assign \g71157/_0_  = _w3999_ ;
	assign \g71158/_0_  = _w4001_ ;
	assign \g71230/_0_  = _w4022_ ;
	assign \g71231/_0_  = _w4043_ ;
	assign \g71232/_0_  = _w4063_ ;
	assign \g71233/_0_  = _w4084_ ;
	assign \g71234/_0_  = _w4104_ ;
	assign \g71235/_0_  = _w4127_ ;
	assign \g71236/_0_  = _w4147_ ;
	assign \g71238/_0_  = _w4167_ ;
	assign \g71239/_0_  = _w4188_ ;
	assign \g71270/_0_  = _w4201_ ;
	assign \g71275/_0_  = _w4223_ ;
	assign \g71276/_0_  = _w4242_ ;
	assign \g71277/_0_  = _w4265_ ;
	assign \g71278/_0_  = _w4280_ ;
	assign \g71279/_0_  = _w4285_ ;
	assign \g71280/_0_  = _w4296_ ;
	assign \g71281/_0_  = _w4304_ ;
	assign \g71282/_0_  = _w4321_ ;
	assign \g71283/_0_  = _w4335_ ;
	assign \g71284/_0_  = _w4349_ ;
	assign \g71285/_0_  = _w4360_ ;
	assign \g71286/_0_  = _w4362_ ;
	assign \g71287/_0_  = _w4375_ ;
	assign \g71288/_0_  = _w4378_ ;
	assign \g71289/_0_  = _w4390_ ;
	assign \g71290/_0_  = _w4398_ ;
	assign \g71291/_0_  = _w4404_ ;
	assign \g71292/_0_  = _w4418_ ;
	assign \g71293/_0_  = _w4431_ ;
	assign \g71294/_0_  = _w4439_ ;
	assign \g71295/_0_  = _w4453_ ;
	assign \g71296/_0_  = _w4467_ ;
	assign \g71297/_0_  = _w4474_ ;
	assign \g71298/_0_  = _w4483_ ;
	assign \g71299/_0_  = _w4485_ ;
	assign \g71300/_0_  = _w4493_ ;
	assign \g71301/_0_  = _w4507_ ;
	assign \g71302/_0_  = _w4520_ ;
	assign \g71303/_0_  = _w4527_ ;
	assign \g71304/_0_  = _w4536_ ;
	assign \g71305/_0_  = _w4552_ ;
	assign \g71306/_0_  = _w4564_ ;
	assign \g71307/_0_  = _w4566_ ;
	assign \g71382/_0_  = _w4583_ ;
	assign \g71384/_0_  = _w4603_ ;
	assign \g71385/_0_  = _w4623_ ;
	assign \g71387/_0_  = _w4641_ ;
	assign \g71388/_0_  = _w4660_ ;
	assign \g71389/_0_  = _w4678_ ;
	assign \g71439/_0_  = _w4689_ ;
	assign \g71440/_0_  = _w4702_ ;
	assign \g71441/_0_  = _w4718_ ;
	assign \g71442/_0_  = _w4725_ ;
	assign \g71443/_0_  = _w4735_ ;
	assign \g71444/_0_  = _w4753_ ;
	assign \g71445/_0_  = _w4764_ ;
	assign \g71446/_0_  = _w4778_ ;
	assign \g71447/_0_  = _w4791_ ;
	assign \g71448/_0_  = _w4803_ ;
	assign \g71449/_0_  = _w4814_ ;
	assign \g71450/_0_  = _w4825_ ;
	assign \g71451/_0_  = _w4838_ ;
	assign \g71452/_0_  = _w4853_ ;
	assign \g71453/_0_  = _w4866_ ;
	assign \g71454/_0_  = _w4881_ ;
	assign \g71455/_0_  = _w4894_ ;
	assign \g71456/_0_  = _w4910_ ;
	assign \g71457/_0_  = _w4926_ ;
	assign \g71458/_0_  = _w4938_ ;
	assign \g71459/_0_  = _w4951_ ;
	assign \g71460/_0_  = _w4961_ ;
	assign \g71461/_0_  = _w4964_ ;
	assign \g71536/_0_  = _w4984_ ;
	assign \g71537/_0_  = _w5002_ ;
	assign \g71538/_0_  = _w5019_ ;
	assign \g71540/_0_  = _w5037_ ;
	assign \g71541/_0_  = _w5056_ ;
	assign \g71542/_0_  = _w5074_ ;
	assign \g71602/_0_  = _w5082_ ;
	assign \g71604/_0_  = _w5087_ ;
	assign \g71610/_0_  = _w5098_ ;
	assign \g71611/_0_  = _w5113_ ;
	assign \g71618/_0_  = _w5115_ ;
	assign \g71619/_0_  = _w5128_ ;
	assign \g71620/_0_  = _w5136_ ;
	assign \g71621/_0_  = _w5149_ ;
	assign \g71622/_0_  = _w5161_ ;
	assign \g71623/_0_  = _w5170_ ;
	assign \g71624/_0_  = _w5174_ ;
	assign \g71625/_0_  = _w5188_ ;
	assign \g71626/_0_  = _w5199_ ;
	assign \g71627/_0_  = _w5205_ ;
	assign \g71629/_0_  = _w5208_ ;
	assign \g71630/_0_  = _w5211_ ;
	assign \g71631/_0_  = _w5213_ ;
	assign \g71632/_0_  = _w5225_ ;
	assign \g71633/_0_  = _w5236_ ;
	assign \g71634/_0_  = _w5242_ ;
	assign \g71635/_0_  = _w5248_ ;
	assign \g71636/_0_  = _w5250_ ;
	assign \g71710/_0_  = _w5269_ ;
	assign \g71711/_0_  = _w5290_ ;
	assign \g71782/_0_  = _w5302_ ;
	assign \g71785/_0_  = _w5308_ ;
	assign \g71786/_0_  = _w5317_ ;
	assign \g71787/_0_  = _w5328_ ;
	assign \g71788/_0_  = _w5340_ ;
	assign \g71789/_0_  = _w5349_ ;
	assign \g71790/_0_  = _w5360_ ;
	assign \g71791/_0_  = _w5368_ ;
	assign \g71792/_0_  = _w5377_ ;
	assign \g71793/_0_  = _w5381_ ;
	assign \g71794/_0_  = _w5390_ ;
	assign \g71795/_0_  = _w5406_ ;
	assign \g71796/_0_  = _w5409_ ;
	assign \g71797/_0_  = _w5412_ ;
	assign \g71798/_0_  = _w5424_ ;
	assign \g71799/_0_  = _w5430_ ;
	assign \g71883/_0_  = _w5446_ ;
	assign \g72000/_0_  = _w5451_ ;
	assign \g72001/_0_  = _w5465_ ;
	assign \g72002/_0_  = _w5476_ ;
	assign \g72003/_0_  = _w5493_ ;
	assign \g72004/_0_  = _w5509_ ;
	assign \g72005/_0_  = _w5511_ ;
	assign \g72236/_0_  = _w5523_ ;
	assign \g72237/_0_  = _w5532_ ;
	assign \g72238/_0_  = _w5544_ ;
	assign \g72239/_0_  = _w5546_ ;
	assign \g72240/_0_  = _w5548_ ;
	assign \g72372/_0_  = _w5559_ ;
	assign \g72376/_0_  = _w5574_ ;
	assign \g72383/_0_  = _w5587_ ;
	assign \g72561/_0_  = _w5592_ ;
	assign \g72562/_0_  = _w5598_ ;
	assign \g72563/_0_  = _w5606_ ;
	assign \g72564/_0_  = _w5613_ ;
	assign \g72970/_0_  = _w5626_ ;
	assign \g72980/_0_  = _w5631_ ;
	assign \g72981/_0_  = _w5638_ ;
	assign \g72982/_0_  = _w5647_ ;
	assign \g72983/_0_  = _w5654_ ;
	assign \g74234/_0_  = _w5664_ ;
	assign \g74260/_0_  = _w5673_ ;
	assign \g75086/_0_  = _w5680_ ;
	assign \g75087/_0_  = _w5683_ ;
	assign \g75088/_0_  = _w5686_ ;
	assign \g75089/_0_  = _w5691_ ;
	assign \g75091/_0_  = _w5694_ ;
	assign \g75092/_0_  = _w5697_ ;
	assign \g80304/_3_  = _w5699_ ;
	assign \g80305/_3_  = _w5701_ ;
	assign \g80306/_3_  = _w5703_ ;
	assign \g80307/_3_  = _w5705_ ;
	assign \g80308/_0_  = _w5707_ ;
	assign \g80309/_0_  = _w5709_ ;
	assign \g80815/_0_  = _w5711_ ;
	assign \g80816/_0_  = _w5713_ ;
	assign \g80817/_0_  = _w5715_ ;
	assign \g80818/_0_  = _w5717_ ;
	assign \g80819/_0_  = _w5719_ ;
	assign \g80820/_0_  = _w5721_ ;
	assign \g80821/_0_  = _w5723_ ;
	assign \g80822/_0_  = _w5725_ ;
	assign \g80823/_0_  = _w5727_ ;
	assign \g80824/_0_  = _w5729_ ;
	assign \g80825/_0_  = _w5731_ ;
	assign \g80826/_3_  = _w5733_ ;
	assign \g80827/_0_  = _w5735_ ;
	assign \g80828/_0_  = _w5737_ ;
	assign \g80829/_0_  = _w5739_ ;
	assign \g80830/_0_  = _w5740_ ;
	assign \g80831/_0_  = _w5742_ ;
	assign \g80832/_0_  = _w5744_ ;
	assign \g80833/_0_  = _w5746_ ;
	assign \g80834/_0_  = _w5748_ ;
	assign \g80835/_0_  = _w5750_ ;
	assign \g80836/_0_  = _w5752_ ;
	assign \g80837/_0_  = _w5754_ ;
	assign \g80838/_3_  = _w5756_ ;
	assign \g80839/_0_  = _w5758_ ;
	assign \g80840/_3_  = _w5760_ ;
	assign \g80841/_0_  = _w5762_ ;
	assign \g80859/_3_  = _w5764_ ;
	assign \g80860/_3_  = _w5766_ ;
	assign \g80861/_3_  = _w5768_ ;
	assign \g80862/_3_  = _w5770_ ;
	assign \g80863/_3_  = _w5772_ ;
	assign \g80864/_3_  = _w5774_ ;
	assign \g80865/_3_  = _w5776_ ;
	assign \g80866/_3_  = _w5778_ ;
	assign \g80867/_3_  = _w5780_ ;
	assign \g80868/_3_  = _w5782_ ;
	assign \g80869/_3_  = _w5784_ ;
	assign \g80870/_3_  = _w5786_ ;
	assign \g80871/_3_  = _w5788_ ;
	assign \g80872/_3_  = _w5790_ ;
	assign \g80873/_3_  = _w5791_ ;
	assign \g80874/_3_  = _w5793_ ;
	assign \g80875/_3_  = _w5795_ ;
	assign \g80876/_3_  = _w5797_ ;
	assign \g80877/_3_  = _w5799_ ;
	assign \g80878/_3_  = _w5801_ ;
	assign \g80879/_0_  = _w5805_ ;
	assign \g80880/_3_  = _w5807_ ;
	assign \g80881/_3_  = _w5809_ ;
	assign \g80882/_3_  = _w5811_ ;
	assign \g80883/_3_  = _w5813_ ;
	assign \g80884/_3_  = _w5815_ ;
	assign \g80885/_3_  = _w5817_ ;
	assign \g80886/_3_  = _w5819_ ;
	assign \g80888/_0_  = _w5823_ ;
	assign \g81262/_0_  = _w1658_ ;
	assign \g81278/_0_  = _w1000_ ;
	assign \g81884/_0_  = _w5856_ ;
	assign \g81893/_0_  = _w5912_ ;
	assign \g81896/_0_  = _w5920_ ;
	assign \g81897/_0_  = _w5936_ ;
	assign \g81898/_0_  = _w5951_ ;
	assign \g81899/_0_  = _w5965_ ;
	assign \g81900/_0_  = _w5985_ ;
	assign \g81901/_0_  = _w6005_ ;
	assign \g81902/_0_  = _w6026_ ;
	assign \g81903/_0_  = _w6046_ ;
	assign \g81904/_0_  = _w6057_ ;
	assign \g81905/_0_  = _w6068_ ;
	assign \g81906/_0_  = _w6082_ ;
	assign \g81907/_0_  = _w6099_ ;
	assign \g81908/_0_  = _w6110_ ;
	assign \g81909/_0_  = _w6120_ ;
	assign \g81910/_0_  = _w6134_ ;
	assign \g81911/_0_  = _w6144_ ;
	assign \g81923/_0_  = _w6164_ ;
	assign \g81924/_0_  = _w6179_ ;
	assign \g81925/_0_  = _w6200_ ;
	assign \g81926/_0_  = _w6217_ ;
	assign \g82414/_0_  = _w6218_ ;
	assign \g82532/_0_  = _w6220_ ;
	assign \g83134/_0_  = _w6245_ ;
	assign \g83135/_0_  = _w6254_ ;
	assign \g83141/_0_  = _w6268_ ;
	assign \g83142/_0_  = _w6280_ ;
	assign \g83145/_0_  = _w6287_ ;
	assign \g83146/_0_  = _w6308_ ;
	assign \g83147/_0_  = _w6327_ ;
	assign \g83148/_0_  = _w6343_ ;
	assign \g83152/_0_  = _w6358_ ;
	assign \g83153/_0_  = _w6374_ ;
	assign \g83154/_0_  = _w6395_ ;
	assign \g83155/_0_  = _w6420_ ;
	assign \g83156/_0_  = _w6439_ ;
	assign \g83157/_0_  = _w6453_ ;
	assign \g83158/_0_  = _w6463_ ;
	assign \g83159/_0_  = _w6475_ ;
	assign \g83164/_0_  = _w6486_ ;
	assign \g83165/_0_  = _w6498_ ;
	assign \g83177/_0_  = _w1292_ ;
	assign \g83178/_0_  = _w2049_ ;
	assign \g83409/_0_  = _w1297_ ;
	assign \g83411/_0_  = _w2054_ ;
	assign \g83807/u3_syn_4  = _w6499_ ;
	assign \g84138/u3_syn_4  = _w6500_ ;
	assign \g85062/_0_  = _w1994_ ;
	assign \g85079/_2_  = _w1484_ ;
	assign \g85113/_0_  = _w1401_ ;
	assign \g85121/_0_  = _w1968_ ;
	assign \g85594/_0_  = _w1808_ ;
	assign \g85663/_0_  = _w603_ ;
	assign \g85669/_0_  = _w678_ ;
	assign \g85749/_0_  = _w1649_ ;
	assign \g85784/_0_  = _w1723_ ;
	assign \g85809/_0_  = _w1753_ ;
	assign \g85817/_0_  = _w1835_ ;
	assign \g85828/_0_  = _w1813_ ;
	assign \g85845/_0_  = _w1618_ ;
	assign \g85851/_0_  = _w1632_ ;
	assign \g85858/_0_  = _w1605_ ;
	assign \g85871/_0_  = _w1450_ ;
	assign \g85882_dup/_0_  = _w1593_ ;
	assign \g85891/_0_  = _w1574_ ;
	assign \g85900/_0_  = _w1565_ ;
	assign \g85905/_0_  = _w1552_ ;
	assign \g85917/_0_  = _w1511_ ;
	assign \g85934/_0_  = _w1692_ ;
	assign \g85949/_0_  = _w1741_ ;
	assign \g85971/_0_  = _w651_ ;
	assign \g85997/_0_  = _w1657_ ;
	assign \g86044/_0_  = _w725_ ;
	assign \g86053/_0_  = _w1064_ ;
	assign \g86063/_0_  = _w981_ ;
	assign \g86082/_0_  = _w709_ ;
	assign \g86088/_0_  = _w790_ ;
	assign \g86098/_0_  = _w765_ ;
	assign \g86105/_0_  = _w838_ ;
	assign \g86179/_0_  = _w828_ ;
	assign \g86256_dup/_0_  = _w857_ ;
	assign \g86264/_0_  = _w848_ ;
	assign \g86273/_0_  = _w950_ ;
	assign \g86281/_0_  = _w781_ ;
	assign \g86288/_0_  = _w877_ ;
	assign \g86297/_0_  = _w890_ ;
	assign \g86304/_0_  = _w912_ ;
	assign \g86310/_0_  = _w900_ ;
	assign \g86320/_0_  = _w801_ ;
	assign \g86328/_0_  = _w811_ ;
	assign \g86339/_0_  = _w755_ ;
	assign \g86353/_0_  = _w928_ ;
	assign \g86360/_0_  = _w939_ ;
	assign \g86368/_0_  = _w740_ ;
	assign \g86373/_0_  = _w962_ ;
	assign \g86385/_0_  = _w972_ ;
	assign \g86392/_0_  = _w999_ ;
	assign \g86399/_0_  = _w990_ ;
	assign \g86421/_0_  = _w1080_ ;
	assign \g86432/_0_  = _w1048_ ;
	assign \g87592/_1__syn_2  = _w2042_ ;
	assign \g87632/_1_  = _w2205_ ;
	assign \g92847/_0_  = _w1826_ ;
	assign \g92957/_0_  = _w6513_ ;
	assign \g93056/_0_  = _w1036_ ;
	assign \g93289/_0_  = _w6527_ ;
	assign \g93538_dup95061/_0_  = _w1765_ ;
	assign \g93856/_0_  = _w6539_ ;
	assign \g93870/_0_  = _w1713_ ;
	assign \g94004/_0_  = _w1543_ ;
	assign \g94128/_0_  = _w1701_ ;
	assign \g94173/_0_  = _w1780_ ;
	assign \g94187/_0_  = _w1676_ ;
	assign \g94191/_0_  = _w1671_ ;
	assign \g94318/_0_  = _w1528_ ;
	assign \g94505/_0_  = _w1639_ ;
	assign rd_pad = _w6540_ ;
	assign \so[0]_pad  = _w6541_ ;
	assign \so[10]_pad  = _w6555_ ;
	assign \so[11]_pad  = _w6558_ ;
	assign \so[12]_pad  = _w6562_ ;
	assign \so[13]_pad  = _w6565_ ;
	assign \so[14]_pad  = _w6568_ ;
	assign \so[15]_pad  = _w6572_ ;
	assign \so[16]_pad  = _w6575_ ;
	assign \so[17]_pad  = _w6578_ ;
	assign \so[18]_pad  = _w6582_ ;
	assign \so[19]_pad  = _w6585_ ;
	assign \so[1]_pad  = _w6586_ ;
	assign \so[2]_pad  = _w6588_ ;
	assign \so[3]_pad  = _w6590_ ;
	assign \so[4]_pad  = _w6592_ ;
	assign \so[5]_pad  = _w6594_ ;
	assign \so[6]_pad  = _w6596_ ;
	assign \so[7]_pad  = _w6598_ ;
	assign \so[8]_pad  = _w6600_ ;
	assign \so[9]_pad  = _w6602_ ;
	assign wr_pad = _w6603_ ;
endmodule;