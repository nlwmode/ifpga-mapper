module top (\G0_pad , \G10_pad , \G11_pad , \G12_pad , \G13_pad , \G14_pad , \G15_pad , \G16_pad , \G18_pad , \G1_pad , \G2_pad , \G38_reg/NET0131 , \G39_reg/NET0131 , \G3_pad , \G40_reg/NET0131 , \G41_reg/NET0131 , \G42_reg/NET0131 , \G4_pad , \G5_pad , \G6_pad , \G7_pad , \G8_pad , \G9_pad , \G288_pad , \G290_pad , \G296_pad , \G302_pad , \G310_pad , \G312_pad , \G315_pad , \G327_pad , \G45_pad , \G47_pad , \G49_pad , \G53_pad , \G55_pad , \_al_n0 , \_al_n1 , \g1452/_0_ , \g1456/_1_ , \g1462/_0_ , \g1463/_0_ , \g1504/_3_ , \g1524/_1_ , \g1524/_2_ , \g1527/_3_ , \g31/_0_ , \g45/_1_ );
	input \G0_pad  ;
	input \G10_pad  ;
	input \G11_pad  ;
	input \G12_pad  ;
	input \G13_pad  ;
	input \G14_pad  ;
	input \G15_pad  ;
	input \G16_pad  ;
	input \G18_pad  ;
	input \G1_pad  ;
	input \G2_pad  ;
	input \G38_reg/NET0131  ;
	input \G39_reg/NET0131  ;
	input \G3_pad  ;
	input \G40_reg/NET0131  ;
	input \G41_reg/NET0131  ;
	input \G42_reg/NET0131  ;
	input \G4_pad  ;
	input \G5_pad  ;
	input \G6_pad  ;
	input \G7_pad  ;
	input \G8_pad  ;
	input \G9_pad  ;
	output \G288_pad  ;
	output \G290_pad  ;
	output \G296_pad  ;
	output \G302_pad  ;
	output \G310_pad  ;
	output \G312_pad  ;
	output \G315_pad  ;
	output \G327_pad  ;
	output \G45_pad  ;
	output \G47_pad  ;
	output \G49_pad  ;
	output \G53_pad  ;
	output \G55_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1452/_0_  ;
	output \g1456/_1_  ;
	output \g1462/_0_  ;
	output \g1463/_0_  ;
	output \g1504/_3_  ;
	output \g1524/_1_  ;
	output \g1524/_2_  ;
	output \g1527/_3_  ;
	output \g31/_0_  ;
	output \g45/_1_  ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w25_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w26_
	);
	LUT3 #(
		.INIT('h40)
	) name2 (
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w27_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		_w25_,
		_w27_,
		_w28_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\G15_pad ,
		\G42_reg/NET0131 ,
		_w29_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w30_
	);
	LUT3 #(
		.INIT('h02)
	) name6 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w31_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		_w29_,
		_w31_,
		_w32_
	);
	LUT3 #(
		.INIT('h08)
	) name8 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w33_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		_w26_,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w35_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		\G16_pad ,
		\G4_pad ,
		_w36_
	);
	LUT3 #(
		.INIT('hc4)
	) name12 (
		\G16_pad ,
		\G40_reg/NET0131 ,
		\G4_pad ,
		_w37_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		\G16_pad ,
		\G40_reg/NET0131 ,
		_w38_
	);
	LUT3 #(
		.INIT('h01)
	) name14 (
		\G1_pad ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w39_
	);
	LUT4 #(
		.INIT('ha888)
	) name15 (
		_w35_,
		_w37_,
		_w38_,
		_w39_,
		_w40_
	);
	LUT3 #(
		.INIT('h02)
	) name16 (
		\G38_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w41_
	);
	LUT4 #(
		.INIT('hccc4)
	) name17 (
		\G38_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w42_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w43_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		_w42_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w46_
	);
	LUT3 #(
		.INIT('h15)
	) name22 (
		\G16_pad ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w47_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w45_,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		\G39_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w49_
	);
	LUT3 #(
		.INIT('hd0)
	) name25 (
		\G38_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		_w49_,
		_w50_,
		_w51_
	);
	LUT3 #(
		.INIT('h40)
	) name27 (
		_w36_,
		_w49_,
		_w50_,
		_w52_
	);
	LUT4 #(
		.INIT('hfffe)
	) name28 (
		_w48_,
		_w40_,
		_w52_,
		_w44_,
		_w53_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w27_,
		_w54_,
		_w55_
	);
	LUT3 #(
		.INIT('h40)
	) name31 (
		\G38_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w57_
	);
	LUT3 #(
		.INIT('h80)
	) name33 (
		\G16_pad ,
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w56_,
		_w58_,
		_w59_
	);
	LUT4 #(
		.INIT('h0001)
	) name35 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w60_
	);
	LUT3 #(
		.INIT('h80)
	) name36 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w61_
	);
	LUT4 #(
		.INIT('h7ffe)
	) name37 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w62_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		\G38_reg/NET0131 ,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\G15_pad ,
		\G42_reg/NET0131 ,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		_w31_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		_w33_,
		_w36_,
		_w66_
	);
	LUT3 #(
		.INIT('h07)
	) name42 (
		\G10_pad ,
		\G11_pad ,
		\G12_pad ,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\G10_pad ,
		\G11_pad ,
		_w68_
	);
	LUT3 #(
		.INIT('h02)
	) name44 (
		\G15_pad ,
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w69_
	);
	LUT3 #(
		.INIT('h10)
	) name45 (
		_w67_,
		_w68_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w66_,
		_w70_,
		_w71_
	);
	LUT3 #(
		.INIT('h40)
	) name47 (
		\G5_pad ,
		_w25_,
		_w27_,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w73_
	);
	LUT2 #(
		.INIT('h6)
	) name49 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w74_
	);
	LUT3 #(
		.INIT('h32)
	) name50 (
		_w41_,
		_w73_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('he)
	) name51 (
		_w51_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w77_
	);
	LUT3 #(
		.INIT('h04)
	) name53 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		_w35_,
		_w78_,
		_w79_
	);
	LUT3 #(
		.INIT('h80)
	) name55 (
		\G5_pad ,
		_w25_,
		_w27_,
		_w80_
	);
	LUT4 #(
		.INIT('h88f3)
	) name56 (
		\G13_pad ,
		\G15_pad ,
		\G38_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w81_
	);
	LUT3 #(
		.INIT('h51)
	) name57 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w81_,
		_w82_
	);
	LUT4 #(
		.INIT('h8000)
	) name58 (
		\G6_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w84_
	);
	LUT3 #(
		.INIT('he0)
	) name60 (
		\G15_pad ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w85_
	);
	LUT4 #(
		.INIT('h1f00)
	) name61 (
		\G40_reg/NET0131 ,
		_w83_,
		_w84_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		_w82_,
		_w86_,
		_w87_
	);
	LUT3 #(
		.INIT('h10)
	) name63 (
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w88_
	);
	LUT4 #(
		.INIT('h0800)
	) name64 (
		\G15_pad ,
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		\G6_pad ,
		_w89_
	);
	LUT3 #(
		.INIT('h01)
	) name65 (
		\G1_pad ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w90_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		\G15_pad ,
		\G42_reg/NET0131 ,
		_w91_
	);
	LUT4 #(
		.INIT('h0111)
	) name67 (
		_w90_,
		_w91_,
		_w88_,
		_w89_,
		_w92_
	);
	LUT4 #(
		.INIT('hb877)
	) name68 (
		\G15_pad ,
		\G39_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w93_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		\G40_reg/NET0131 ,
		_w93_,
		_w94_
	);
	LUT3 #(
		.INIT('h0d)
	) name70 (
		_w35_,
		_w92_,
		_w94_,
		_w95_
	);
	LUT3 #(
		.INIT('h23)
	) name71 (
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		\G5_pad ,
		_w96_
	);
	LUT4 #(
		.INIT('h0100)
	) name72 (
		\G1_pad ,
		\G3_pad ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w97_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name73 (
		\G2_pad ,
		_w57_,
		_w96_,
		_w97_,
		_w98_
	);
	LUT4 #(
		.INIT('hea00)
	) name74 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		\G4_pad ,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		\G14_pad ,
		\G15_pad ,
		_w100_
	);
	LUT4 #(
		.INIT('h5450)
	) name76 (
		\G39_reg/NET0131 ,
		_w78_,
		_w99_,
		_w100_,
		_w101_
	);
	LUT3 #(
		.INIT('h40)
	) name77 (
		\G0_pad ,
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w102_
	);
	LUT4 #(
		.INIT('hb0bf)
	) name78 (
		\G0_pad ,
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w103_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name79 (
		_w42_,
		_w43_,
		_w61_,
		_w103_,
		_w104_
	);
	LUT4 #(
		.INIT('hab00)
	) name80 (
		\G38_reg/NET0131 ,
		_w98_,
		_w101_,
		_w104_,
		_w105_
	);
	LUT4 #(
		.INIT('h7500)
	) name81 (
		\G16_pad ,
		_w87_,
		_w95_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		\G18_pad ,
		_w106_,
		_w107_
	);
	LUT4 #(
		.INIT('h5150)
	) name83 (
		\G38_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		\G5_pad ,
		_w108_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		_w97_,
		_w108_,
		_w109_
	);
	LUT3 #(
		.INIT('h01)
	) name85 (
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		\G4_pad ,
		_w110_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name86 (
		\G0_pad ,
		\G38_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w111_
	);
	LUT3 #(
		.INIT('h8a)
	) name87 (
		_w57_,
		_w110_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		_w109_,
		_w112_,
		_w113_
	);
	LUT3 #(
		.INIT('h04)
	) name89 (
		\G1_pad ,
		\G2_pad ,
		\G3_pad ,
		_w114_
	);
	LUT4 #(
		.INIT('h0010)
	) name90 (
		\G16_pad ,
		\G1_pad ,
		\G2_pad ,
		\G3_pad ,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		\G41_reg/NET0131 ,
		_w115_,
		_w116_
	);
	LUT3 #(
		.INIT('hb0)
	) name92 (
		\G14_pad ,
		\G15_pad ,
		\G41_reg/NET0131 ,
		_w117_
	);
	LUT3 #(
		.INIT('h08)
	) name93 (
		_w35_,
		_w77_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		_w116_,
		_w118_,
		_w119_
	);
	LUT3 #(
		.INIT('h2a)
	) name95 (
		\G38_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w120_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w121_
	);
	LUT3 #(
		.INIT('hc8)
	) name97 (
		\G15_pad ,
		\G16_pad ,
		\G40_reg/NET0131 ,
		_w122_
	);
	LUT3 #(
		.INIT('h40)
	) name98 (
		_w120_,
		_w121_,
		_w122_,
		_w123_
	);
	LUT4 #(
		.INIT('h2333)
	) name99 (
		\G38_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w124_
	);
	LUT3 #(
		.INIT('h0e)
	) name100 (
		\G10_pad ,
		\G11_pad ,
		\G42_reg/NET0131 ,
		_w125_
	);
	LUT3 #(
		.INIT('h80)
	) name101 (
		\G15_pad ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w126_
	);
	LUT3 #(
		.INIT('h45)
	) name102 (
		_w124_,
		_w125_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		\G15_pad ,
		\G38_reg/NET0131 ,
		_w128_
	);
	LUT3 #(
		.INIT('h2a)
	) name104 (
		\G16_pad ,
		_w83_,
		_w128_,
		_w129_
	);
	LUT3 #(
		.INIT('h02)
	) name105 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G4_pad ,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w46_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name107 (
		_w129_,
		_w131_,
		_w132_
	);
	LUT4 #(
		.INIT('h7077)
	) name108 (
		_w123_,
		_w127_,
		_w129_,
		_w131_,
		_w133_
	);
	LUT4 #(
		.INIT('h5455)
	) name109 (
		\G18_pad ,
		_w113_,
		_w119_,
		_w133_,
		_w134_
	);
	LUT3 #(
		.INIT('h40)
	) name110 (
		\G38_reg/NET0131 ,
		_w60_,
		_w115_,
		_w135_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		_w47_,
		_w130_,
		_w136_
	);
	LUT4 #(
		.INIT('h0006)
	) name112 (
		\G10_pad ,
		\G11_pad ,
		\G12_pad ,
		\G42_reg/NET0131 ,
		_w137_
	);
	LUT4 #(
		.INIT('h0020)
	) name113 (
		\G16_pad ,
		\G39_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G4_pad ,
		_w138_
	);
	LUT4 #(
		.INIT('ha020)
	) name114 (
		\G15_pad ,
		\G38_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w139_
	);
	LUT3 #(
		.INIT('h40)
	) name115 (
		_w137_,
		_w138_,
		_w139_,
		_w140_
	);
	LUT3 #(
		.INIT('h01)
	) name116 (
		_w136_,
		_w140_,
		_w135_,
		_w141_
	);
	LUT3 #(
		.INIT('h45)
	) name117 (
		\G18_pad ,
		_w113_,
		_w141_,
		_w142_
	);
	LUT3 #(
		.INIT('h01)
	) name118 (
		\G16_pad ,
		\G1_pad ,
		\G38_reg/NET0131 ,
		_w143_
	);
	LUT4 #(
		.INIT('hc05f)
	) name119 (
		\G0_pad ,
		\G16_pad ,
		\G38_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w144_
	);
	LUT3 #(
		.INIT('h20)
	) name120 (
		_w30_,
		_w143_,
		_w144_,
		_w145_
	);
	LUT3 #(
		.INIT('h13)
	) name121 (
		\G10_pad ,
		\G11_pad ,
		\G12_pad ,
		_w146_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		\G15_pad ,
		\G38_reg/NET0131 ,
		_w147_
	);
	LUT4 #(
		.INIT('h0800)
	) name123 (
		_w33_,
		_w36_,
		_w146_,
		_w147_,
		_w148_
	);
	LUT3 #(
		.INIT('h54)
	) name124 (
		\G39_reg/NET0131 ,
		_w145_,
		_w148_,
		_w149_
	);
	LUT3 #(
		.INIT('hb0)
	) name125 (
		\G0_pad ,
		\G38_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w150_
	);
	LUT2 #(
		.INIT('h2)
	) name126 (
		\G1_pad ,
		\G38_reg/NET0131 ,
		_w151_
	);
	LUT3 #(
		.INIT('h0d)
	) name127 (
		\G1_pad ,
		\G38_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w152_
	);
	LUT3 #(
		.INIT('h80)
	) name128 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w153_
	);
	LUT3 #(
		.INIT('h04)
	) name129 (
		_w152_,
		_w153_,
		_w150_,
		_w154_
	);
	LUT3 #(
		.INIT('h0e)
	) name130 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G4_pad ,
		_w155_
	);
	LUT4 #(
		.INIT('h8880)
	) name131 (
		\G16_pad ,
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w156_
	);
	LUT4 #(
		.INIT('h773f)
	) name132 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w157_
	);
	LUT3 #(
		.INIT('h80)
	) name133 (
		_w155_,
		_w156_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		_w154_,
		_w158_,
		_w159_
	);
	LUT3 #(
		.INIT('h45)
	) name135 (
		\G18_pad ,
		_w149_,
		_w159_,
		_w160_
	);
	LUT3 #(
		.INIT('h31)
	) name136 (
		\G39_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w161_
	);
	LUT3 #(
		.INIT('h74)
	) name137 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w162_
	);
	LUT3 #(
		.INIT('h20)
	) name138 (
		_w151_,
		_w162_,
		_w161_,
		_w163_
	);
	LUT3 #(
		.INIT('h80)
	) name139 (
		\G15_pad ,
		_w35_,
		_w78_,
		_w164_
	);
	LUT3 #(
		.INIT('h80)
	) name140 (
		_w35_,
		_w78_,
		_w100_,
		_w165_
	);
	LUT3 #(
		.INIT('h80)
	) name141 (
		\G3_pad ,
		_w60_,
		_w143_,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		\G39_reg/NET0131 ,
		_w99_,
		_w167_
	);
	LUT4 #(
		.INIT('h0800)
	) name143 (
		\G15_pad ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w168_
	);
	LUT4 #(
		.INIT('hf3d1)
	) name144 (
		\G16_pad ,
		_w77_,
		_w117_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		\G41_reg/NET0131 ,
		\G5_pad ,
		_w170_
	);
	LUT3 #(
		.INIT('h8c)
	) name146 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G4_pad ,
		_w171_
	);
	LUT4 #(
		.INIT('h40fc)
	) name147 (
		\G16_pad ,
		\G39_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w172_
	);
	LUT3 #(
		.INIT('h40)
	) name148 (
		_w170_,
		_w171_,
		_w172_,
		_w173_
	);
	LUT3 #(
		.INIT('hc1)
	) name149 (
		\G16_pad ,
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w174_
	);
	LUT3 #(
		.INIT('h80)
	) name150 (
		_w114_,
		_w161_,
		_w174_,
		_w175_
	);
	LUT4 #(
		.INIT('h0111)
	) name151 (
		_w173_,
		_w175_,
		_w167_,
		_w169_,
		_w176_
	);
	LUT3 #(
		.INIT('h80)
	) name152 (
		\G15_pad ,
		\G39_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w177_
	);
	LUT4 #(
		.INIT('h7100)
	) name153 (
		\G15_pad ,
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w178_
	);
	LUT3 #(
		.INIT('h02)
	) name154 (
		\G16_pad ,
		\G40_reg/NET0131 ,
		\G4_pad ,
		_w179_
	);
	LUT4 #(
		.INIT('hf400)
	) name155 (
		_w83_,
		_w177_,
		_w178_,
		_w179_,
		_w180_
	);
	LUT3 #(
		.INIT('h80)
	) name156 (
		\G13_pad ,
		\G15_pad ,
		\G16_pad ,
		_w181_
	);
	LUT4 #(
		.INIT('h88a8)
	) name157 (
		_w61_,
		_w102_,
		_w121_,
		_w181_,
		_w182_
	);
	LUT4 #(
		.INIT('h040c)
	) name158 (
		\G15_pad ,
		\G16_pad ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w183_
	);
	LUT3 #(
		.INIT('h04)
	) name159 (
		_w46_,
		_w130_,
		_w183_,
		_w184_
	);
	LUT3 #(
		.INIT('h01)
	) name160 (
		_w182_,
		_w184_,
		_w180_,
		_w185_
	);
	LUT4 #(
		.INIT('h0155)
	) name161 (
		\G18_pad ,
		\G38_reg/NET0131 ,
		_w176_,
		_w185_,
		_w186_
	);
	assign \G288_pad  = _w28_ ;
	assign \G290_pad  = _w32_ ;
	assign \G296_pad  = _w34_ ;
	assign \G302_pad  = _w53_ ;
	assign \G310_pad  = _w55_ ;
	assign \G312_pad  = _w59_ ;
	assign \G315_pad  = _w63_ ;
	assign \G327_pad  = _w65_ ;
	assign \G45_pad  = _w71_ ;
	assign \G47_pad  = _w72_ ;
	assign \G49_pad  = _w76_ ;
	assign \G53_pad  = _w79_ ;
	assign \G55_pad  = _w80_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g1452/_0_  = _w107_ ;
	assign \g1456/_1_  = _w134_ ;
	assign \g1462/_0_  = _w142_ ;
	assign \g1463/_0_  = _w160_ ;
	assign \g1504/_3_  = _w163_ ;
	assign \g1524/_1_  = _w164_ ;
	assign \g1524/_2_  = _w165_ ;
	assign \g1527/_3_  = _w166_ ;
	assign \g31/_0_  = _w186_ ;
	assign \g45/_1_  = _w132_ ;
endmodule;