module top( \IN_R_reg[0]/NET0131  , \IN_R_reg[1]/NET0131  , \IN_R_reg[2]/NET0131  , \IN_R_reg[3]/NET0131  , \IN_R_reg[4]/NET0131  , \IN_R_reg[5]/NET0131  , \IN_R_reg[6]/NET0131  , \IN_R_reg[7]/NET0131  , \I[0]_pad  , \I[1]_pad  , \I[2]_pad  , \I[3]_pad  , \I[4]_pad  , \I[5]_pad  , \I[6]_pad  , \I[7]_pad  , \MAR_reg[0]/NET0131  , \MAR_reg[1]/NET0131  , \MAR_reg[2]/NET0131  , \OUT_R_reg[0]/NET0131  , \OUT_R_reg[1]/NET0131  , \OUT_R_reg[2]/NET0131  , \OUT_R_reg[3]/NET0131  , \O[0]_pad  , \O[1]_pad  , \O[2]_pad  , \O[3]_pad  , START_pad , \STATO_reg[0]/NET0131  , \STATO_reg[1]/NET0131  , \_al_n0  , \_al_n1  , \g1016/_0_  , \g1017/_0_  , \g1018/_0_  , \g1019/_0_  , \g1041/_0_  , \g1052/_0_  , \g1053/_0_  , \g1054/_0_  , \g1058/_0_  , \g1059/_0_  , \g1060/_0_  , \g1061/_0_  , \g1063/_0_  , \g1090/_0_  , \g1093/_0_  , \g1095/_0_  , \g1098/_0_  , \g1099/_0_  , \g1100/_0_  , \g1101/_0_  , \g1102/_0_  );
  input \IN_R_reg[0]/NET0131  ;
  input \IN_R_reg[1]/NET0131  ;
  input \IN_R_reg[2]/NET0131  ;
  input \IN_R_reg[3]/NET0131  ;
  input \IN_R_reg[4]/NET0131  ;
  input \IN_R_reg[5]/NET0131  ;
  input \IN_R_reg[6]/NET0131  ;
  input \IN_R_reg[7]/NET0131  ;
  input \I[0]_pad  ;
  input \I[1]_pad  ;
  input \I[2]_pad  ;
  input \I[3]_pad  ;
  input \I[4]_pad  ;
  input \I[5]_pad  ;
  input \I[6]_pad  ;
  input \I[7]_pad  ;
  input \MAR_reg[0]/NET0131  ;
  input \MAR_reg[1]/NET0131  ;
  input \MAR_reg[2]/NET0131  ;
  input \OUT_R_reg[0]/NET0131  ;
  input \OUT_R_reg[1]/NET0131  ;
  input \OUT_R_reg[2]/NET0131  ;
  input \OUT_R_reg[3]/NET0131  ;
  input \O[0]_pad  ;
  input \O[1]_pad  ;
  input \O[2]_pad  ;
  input \O[3]_pad  ;
  input START_pad ;
  input \STATO_reg[0]/NET0131  ;
  input \STATO_reg[1]/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1016/_0_  ;
  output \g1017/_0_  ;
  output \g1018/_0_  ;
  output \g1019/_0_  ;
  output \g1041/_0_  ;
  output \g1052/_0_  ;
  output \g1053/_0_  ;
  output \g1054/_0_  ;
  output \g1058/_0_  ;
  output \g1059/_0_  ;
  output \g1060/_0_  ;
  output \g1061/_0_  ;
  output \g1063/_0_  ;
  output \g1090/_0_  ;
  output \g1093/_0_  ;
  output \g1095/_0_  ;
  output \g1098/_0_  ;
  output \g1099/_0_  ;
  output \g1100/_0_  ;
  output \g1101/_0_  ;
  output \g1102/_0_  ;
  wire n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 ;
  assign n31 = \MAR_reg[0]/NET0131  & \MAR_reg[1]/NET0131  ;
  assign n32 = ~\MAR_reg[0]/NET0131  & ~\MAR_reg[1]/NET0131  ;
  assign n33 = ~n31 & ~n32 ;
  assign n34 = \MAR_reg[1]/NET0131  & \MAR_reg[2]/NET0131  ;
  assign n35 = ~\IN_R_reg[1]/NET0131  & ~n34 ;
  assign n36 = \IN_R_reg[1]/NET0131  & \MAR_reg[2]/NET0131  ;
  assign n37 = ~n35 & ~n36 ;
  assign n38 = n33 & n37 ;
  assign n39 = \MAR_reg[0]/NET0131  & \MAR_reg[2]/NET0131  ;
  assign n40 = \IN_R_reg[2]/NET0131  & ~n39 ;
  assign n41 = n33 & n40 ;
  assign n42 = \MAR_reg[1]/NET0131  & ~\MAR_reg[2]/NET0131  ;
  assign n43 = ~\MAR_reg[1]/NET0131  & \MAR_reg[2]/NET0131  ;
  assign n44 = ~n42 & ~n43 ;
  assign n45 = ~\IN_R_reg[2]/NET0131  & \MAR_reg[0]/NET0131  ;
  assign n46 = ~n44 & n45 ;
  assign n47 = ~n41 & ~n46 ;
  assign n48 = ~n38 & n47 ;
  assign n49 = ~\IN_R_reg[3]/NET0131  & ~n42 ;
  assign n50 = ~\MAR_reg[0]/NET0131  & ~\MAR_reg[2]/NET0131  ;
  assign n51 = ~\IN_R_reg[7]/NET0131  & \MAR_reg[1]/NET0131  ;
  assign n52 = ~n50 & n51 ;
  assign n53 = ~n49 & ~n52 ;
  assign n54 = ~n39 & ~n53 ;
  assign n55 = n48 & ~n54 ;
  assign n56 = \IN_R_reg[5]/NET0131  & \MAR_reg[2]/NET0131  ;
  assign n57 = ~\IN_R_reg[0]/NET0131  & ~n56 ;
  assign n58 = ~\MAR_reg[0]/NET0131  & ~n57 ;
  assign n59 = \MAR_reg[0]/NET0131  & ~\MAR_reg[2]/NET0131  ;
  assign n60 = \IN_R_reg[4]/NET0131  & ~n59 ;
  assign n61 = ~\IN_R_reg[4]/NET0131  & n59 ;
  assign n62 = ~n60 & ~n61 ;
  assign n63 = ~n58 & n62 ;
  assign n64 = \MAR_reg[1]/NET0131  & ~n63 ;
  assign n65 = ~\IN_R_reg[5]/NET0131  & ~\MAR_reg[2]/NET0131  ;
  assign n66 = ~\MAR_reg[1]/NET0131  & n65 ;
  assign n67 = ~\IN_R_reg[0]/NET0131  & ~\MAR_reg[1]/NET0131  ;
  assign n68 = ~n50 & n67 ;
  assign n69 = ~n66 & ~n68 ;
  assign n70 = ~n64 & n69 ;
  assign n71 = n55 & n70 ;
  assign n72 = ~\STATO_reg[0]/NET0131  & \STATO_reg[1]/NET0131  ;
  assign n73 = \STATO_reg[0]/NET0131  & ~\STATO_reg[1]/NET0131  ;
  assign n74 = ~n72 & ~n73 ;
  assign n75 = ~\MAR_reg[0]/NET0131  & \MAR_reg[2]/NET0131  ;
  assign n76 = \MAR_reg[0]/NET0131  & n42 ;
  assign n77 = ~\MAR_reg[1]/NET0131  & ~n59 ;
  assign n78 = \IN_R_reg[6]/NET0131  & ~n77 ;
  assign n79 = ~n76 & n78 ;
  assign n80 = ~\IN_R_reg[6]/NET0131  & ~\MAR_reg[1]/NET0131  ;
  assign n81 = ~n59 & n80 ;
  assign n82 = \IN_R_reg[7]/NET0131  & n44 ;
  assign n83 = ~n81 & ~n82 ;
  assign n84 = ~n79 & n83 ;
  assign n85 = ~n75 & ~n84 ;
  assign n86 = ~n74 & ~n85 ;
  assign n87 = n71 & n86 ;
  assign n88 = \OUT_R_reg[3]/NET0131  & ~n73 ;
  assign n89 = ~n87 & n88 ;
  assign n90 = \MAR_reg[0]/NET0131  & ~\OUT_R_reg[3]/NET0131  ;
  assign n91 = n44 & n90 ;
  assign n92 = n72 & ~n91 ;
  assign n93 = ~n85 & n92 ;
  assign n94 = n71 & n93 ;
  assign n95 = ~n89 & ~n94 ;
  assign n96 = \OUT_R_reg[1]/NET0131  & ~n73 ;
  assign n97 = ~n87 & n96 ;
  assign n98 = ~\OUT_R_reg[1]/NET0131  & n39 ;
  assign n99 = n72 & ~n98 ;
  assign n100 = ~n85 & n99 ;
  assign n101 = n71 & n100 ;
  assign n102 = ~n97 & ~n101 ;
  assign n103 = \OUT_R_reg[0]/NET0131  & ~n73 ;
  assign n104 = ~n87 & n103 ;
  assign n105 = ~\MAR_reg[0]/NET0131  & \MAR_reg[1]/NET0131  ;
  assign n106 = ~\OUT_R_reg[0]/NET0131  & ~n105 ;
  assign n107 = n72 & ~n106 ;
  assign n108 = ~n85 & n107 ;
  assign n109 = n71 & n108 ;
  assign n110 = ~n104 & ~n109 ;
  assign n111 = \OUT_R_reg[2]/NET0131  & ~n73 ;
  assign n112 = ~n87 & n111 ;
  assign n113 = ~\MAR_reg[0]/NET0131  & ~n44 ;
  assign n114 = \MAR_reg[2]/NET0131  & n31 ;
  assign n115 = ~\OUT_R_reg[2]/NET0131  & ~n114 ;
  assign n116 = ~n113 & n115 ;
  assign n117 = n72 & ~n116 ;
  assign n118 = ~n85 & n117 ;
  assign n119 = n71 & n118 ;
  assign n120 = ~n112 & ~n119 ;
  assign n121 = \STATO_reg[0]/NET0131  & \STATO_reg[1]/NET0131  ;
  assign n122 = n31 & n121 ;
  assign n123 = \MAR_reg[2]/NET0131  & ~n73 ;
  assign n124 = ~n122 & ~n123 ;
  assign n125 = \MAR_reg[1]/NET0131  & ~\STATO_reg[0]/NET0131  ;
  assign n126 = ~n32 & n121 ;
  assign n127 = ~n76 & n126 ;
  assign n128 = ~n125 & ~n127 ;
  assign n129 = \MAR_reg[1]/NET0131  & \STATO_reg[1]/NET0131  ;
  assign n130 = n39 & n129 ;
  assign n131 = \STATO_reg[0]/NET0131  & ~n130 ;
  assign n132 = ~START_pad & ~n72 ;
  assign n133 = ~n131 & ~n132 ;
  assign n134 = \MAR_reg[0]/NET0131  & ~START_pad ;
  assign n135 = n34 & n134 ;
  assign n136 = n121 & ~n135 ;
  assign n137 = n74 & ~n136 ;
  assign n138 = n121 & n135 ;
  assign n139 = \O[0]_pad  & ~n138 ;
  assign n140 = \OUT_R_reg[0]/NET0131  & n121 ;
  assign n141 = n135 & n140 ;
  assign n142 = ~n139 & ~n141 ;
  assign n143 = \O[1]_pad  & ~n138 ;
  assign n144 = \OUT_R_reg[1]/NET0131  & n121 ;
  assign n145 = n135 & n144 ;
  assign n146 = ~n143 & ~n145 ;
  assign n147 = \O[2]_pad  & ~n138 ;
  assign n148 = \OUT_R_reg[2]/NET0131  & n121 ;
  assign n149 = n135 & n148 ;
  assign n150 = ~n147 & ~n149 ;
  assign n151 = \O[3]_pad  & ~n138 ;
  assign n152 = \OUT_R_reg[3]/NET0131  & n121 ;
  assign n153 = n135 & n152 ;
  assign n154 = ~n151 & ~n153 ;
  assign n155 = \MAR_reg[0]/NET0131  & \STATO_reg[0]/NET0131  ;
  assign n156 = ~n34 & n155 ;
  assign n157 = ~\MAR_reg[0]/NET0131  & ~\STATO_reg[0]/NET0131  ;
  assign n158 = ~n73 & ~n157 ;
  assign n159 = ~n156 & n158 ;
  assign n160 = \IN_R_reg[2]/NET0131  & ~n73 ;
  assign n161 = \I[2]_pad  & n73 ;
  assign n162 = ~n160 & ~n161 ;
  assign n163 = \IN_R_reg[6]/NET0131  & ~n73 ;
  assign n164 = \I[6]_pad  & n73 ;
  assign n165 = ~n163 & ~n164 ;
  assign n166 = \IN_R_reg[7]/NET0131  & ~n73 ;
  assign n167 = \I[7]_pad  & n73 ;
  assign n168 = ~n166 & ~n167 ;
  assign n169 = \IN_R_reg[3]/NET0131  & ~n73 ;
  assign n170 = \I[3]_pad  & n73 ;
  assign n171 = ~n169 & ~n170 ;
  assign n172 = \IN_R_reg[0]/NET0131  & ~n73 ;
  assign n173 = \I[0]_pad  & n73 ;
  assign n174 = ~n172 & ~n173 ;
  assign n175 = \IN_R_reg[4]/NET0131  & ~n73 ;
  assign n176 = \I[4]_pad  & n73 ;
  assign n177 = ~n175 & ~n176 ;
  assign n178 = \IN_R_reg[5]/NET0131  & ~n73 ;
  assign n179 = \I[5]_pad  & n73 ;
  assign n180 = ~n178 & ~n179 ;
  assign n181 = \IN_R_reg[1]/NET0131  & ~n73 ;
  assign n182 = \I[1]_pad  & n73 ;
  assign n183 = ~n181 & ~n182 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1016/_0_  = ~n95 ;
  assign \g1017/_0_  = ~n102 ;
  assign \g1018/_0_  = ~n110 ;
  assign \g1019/_0_  = ~n120 ;
  assign \g1041/_0_  = ~n124 ;
  assign \g1052/_0_  = ~n128 ;
  assign \g1053/_0_  = n133 ;
  assign \g1054/_0_  = ~n137 ;
  assign \g1058/_0_  = ~n142 ;
  assign \g1059/_0_  = ~n146 ;
  assign \g1060/_0_  = ~n150 ;
  assign \g1061/_0_  = ~n154 ;
  assign \g1063/_0_  = n159 ;
  assign \g1090/_0_  = ~n162 ;
  assign \g1093/_0_  = ~n165 ;
  assign \g1095/_0_  = ~n168 ;
  assign \g1098/_0_  = ~n171 ;
  assign \g1099/_0_  = ~n174 ;
  assign \g1100/_0_  = ~n177 ;
  assign \g1101/_0_  = ~n180 ;
  assign \g1102/_0_  = ~n183 ;
endmodule
