module top( \ACVQN0_reg/NET0131  , \ACVQN1_reg/NET0131  , \ACVQN2_reg/NET0131  , \ACVQN3_reg/NET0131  , \AX0_reg/NET0131  , \AX1_reg/NET0131  , \AX2_reg/NET0131  , \AX3_reg/NET0131  , \B0_pad  , \B1_pad  , \B2_pad  , \B3_pad  , \CT0_reg/NET0131  , \CT1_reg/NET0131  , \CT2_reg/NET0131  , \MRVQN0_reg/NET0131  , \MRVQN1_reg/NET0131  , \MRVQN2_reg/NET0131  , \MRVQN3_reg/NET0131  , START_pad , \ACVQN0_reg/P0001  , \ACVQN1_reg/P0001  , \ACVQN2_reg/P0001  , \ACVQN3_reg/P0001  , \CNTVCON2_pad  , \MRVQN0_reg/P0001  , \P1_pad  , \P2_pad  , \P3_pad  , \_al_n0  , \_al_n1  , \g12/_0_  , \g20/_0_  , \g31/_0_  , \g616/_0_  , \g630/_0_  , \g632/_0_  , \g633/_0_  , \g636/_0_  , \g637/_0_  , \g638/_0_  , \g673/_1__syn_2  , \g675/_1_  , \g795/_0_  , \g810/_0_  );
  input \ACVQN0_reg/NET0131  ;
  input \ACVQN1_reg/NET0131  ;
  input \ACVQN2_reg/NET0131  ;
  input \ACVQN3_reg/NET0131  ;
  input \AX0_reg/NET0131  ;
  input \AX1_reg/NET0131  ;
  input \AX2_reg/NET0131  ;
  input \AX3_reg/NET0131  ;
  input \B0_pad  ;
  input \B1_pad  ;
  input \B2_pad  ;
  input \B3_pad  ;
  input \CT0_reg/NET0131  ;
  input \CT1_reg/NET0131  ;
  input \CT2_reg/NET0131  ;
  input \MRVQN0_reg/NET0131  ;
  input \MRVQN1_reg/NET0131  ;
  input \MRVQN2_reg/NET0131  ;
  input \MRVQN3_reg/NET0131  ;
  input START_pad ;
  output \ACVQN0_reg/P0001  ;
  output \ACVQN1_reg/P0001  ;
  output \ACVQN2_reg/P0001  ;
  output \ACVQN3_reg/P0001  ;
  output \CNTVCON2_pad  ;
  output \MRVQN0_reg/P0001  ;
  output \P1_pad  ;
  output \P2_pad  ;
  output \P3_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g12/_0_  ;
  output \g20/_0_  ;
  output \g31/_0_  ;
  output \g616/_0_  ;
  output \g630/_0_  ;
  output \g632/_0_  ;
  output \g633/_0_  ;
  output \g636/_0_  ;
  output \g637/_0_  ;
  output \g638/_0_  ;
  output \g673/_1__syn_2  ;
  output \g675/_1_  ;
  output \g795/_0_  ;
  output \g810/_0_  ;
  wire n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 ;
  assign n21 = \CT0_reg/NET0131  & \CT2_reg/NET0131  ;
  assign n22 = \CT1_reg/NET0131  & n21 ;
  assign n23 = ~\CT1_reg/NET0131  & n21 ;
  assign n28 = \AX3_reg/NET0131  & ~\MRVQN0_reg/NET0131  ;
  assign n29 = \ACVQN3_reg/NET0131  & ~n28 ;
  assign n30 = ~\ACVQN3_reg/NET0131  & n28 ;
  assign n31 = ~n29 & ~n30 ;
  assign n32 = \AX2_reg/NET0131  & ~\MRVQN0_reg/NET0131  ;
  assign n33 = \ACVQN2_reg/NET0131  & ~n32 ;
  assign n34 = ~\ACVQN2_reg/NET0131  & n32 ;
  assign n35 = ~\ACVQN0_reg/NET0131  & \AX0_reg/NET0131  ;
  assign n36 = ~\MRVQN0_reg/NET0131  & n35 ;
  assign n37 = \ACVQN1_reg/NET0131  & ~n36 ;
  assign n38 = ~\ACVQN1_reg/NET0131  & n36 ;
  assign n39 = \AX1_reg/NET0131  & ~\MRVQN0_reg/NET0131  ;
  assign n40 = ~n38 & ~n39 ;
  assign n41 = ~n37 & ~n40 ;
  assign n42 = ~n34 & ~n41 ;
  assign n43 = ~n33 & ~n42 ;
  assign n45 = n31 & ~n43 ;
  assign n24 = ~\CT0_reg/NET0131  & ~\CT1_reg/NET0131  ;
  assign n25 = ~\CT2_reg/NET0131  & n24 ;
  assign n26 = ~n23 & ~n25 ;
  assign n44 = ~n31 & n43 ;
  assign n46 = n26 & ~n44 ;
  assign n47 = ~n45 & n46 ;
  assign n27 = \ACVQN2_reg/NET0131  & ~n26 ;
  assign n48 = ~START_pad & ~n27 ;
  assign n49 = ~n47 & n48 ;
  assign n51 = ~n29 & n43 ;
  assign n52 = n26 & ~n30 ;
  assign n53 = ~n51 & n52 ;
  assign n50 = \ACVQN3_reg/NET0131  & ~n26 ;
  assign n54 = ~START_pad & ~n50 ;
  assign n55 = ~n53 & n54 ;
  assign n57 = \CT0_reg/NET0131  & ~n23 ;
  assign n58 = ~\CT1_reg/NET0131  & ~n57 ;
  assign n56 = \CT0_reg/NET0131  & \CT1_reg/NET0131  ;
  assign n59 = ~START_pad & ~n56 ;
  assign n60 = ~n58 & n59 ;
  assign n61 = ~\CT2_reg/NET0131  & ~n56 ;
  assign n62 = ~START_pad & ~n22 ;
  assign n63 = ~n61 & n62 ;
  assign n64 = \AX0_reg/NET0131  & ~\MRVQN0_reg/NET0131  ;
  assign n65 = \ACVQN0_reg/NET0131  & ~n64 ;
  assign n66 = ~n36 & ~n65 ;
  assign n67 = n26 & ~n66 ;
  assign n69 = \B3_pad  & ~n23 ;
  assign n68 = ~\MRVQN3_reg/NET0131  & n23 ;
  assign n70 = ~n26 & ~n68 ;
  assign n71 = ~n69 & n70 ;
  assign n72 = ~n67 & ~n71 ;
  assign n73 = ~START_pad & ~n57 ;
  assign n74 = ~\B2_pad  & ~n23 ;
  assign n75 = \MRVQN2_reg/NET0131  & n23 ;
  assign n76 = ~n74 & ~n75 ;
  assign n77 = ~n26 & ~n76 ;
  assign n78 = \MRVQN3_reg/NET0131  & n26 ;
  assign n79 = ~n77 & ~n78 ;
  assign n80 = ~\B0_pad  & ~n23 ;
  assign n81 = \MRVQN0_reg/NET0131  & n23 ;
  assign n82 = ~n80 & ~n81 ;
  assign n83 = ~n26 & ~n82 ;
  assign n84 = \MRVQN1_reg/NET0131  & n26 ;
  assign n85 = ~n83 & ~n84 ;
  assign n86 = ~\B1_pad  & ~n23 ;
  assign n87 = \MRVQN1_reg/NET0131  & n23 ;
  assign n88 = ~n86 & ~n87 ;
  assign n89 = ~n26 & ~n88 ;
  assign n90 = \MRVQN2_reg/NET0131  & n26 ;
  assign n91 = ~n89 & ~n90 ;
  assign n94 = n37 & ~n39 ;
  assign n95 = ~n41 & ~n94 ;
  assign n93 = \AX1_reg/NET0131  & n38 ;
  assign n96 = n26 & ~n93 ;
  assign n97 = ~n95 & n96 ;
  assign n92 = \ACVQN0_reg/NET0131  & ~n26 ;
  assign n98 = ~START_pad & ~n92 ;
  assign n99 = ~n97 & n98 ;
  assign n102 = n33 & ~n41 ;
  assign n103 = ~n43 & ~n102 ;
  assign n101 = n34 & n41 ;
  assign n104 = n26 & ~n101 ;
  assign n105 = ~n103 & n104 ;
  assign n100 = \ACVQN1_reg/NET0131  & ~n26 ;
  assign n106 = ~START_pad & ~n100 ;
  assign n107 = ~n105 & n106 ;
  assign \ACVQN0_reg/P0001  = ~\ACVQN0_reg/NET0131  ;
  assign \ACVQN1_reg/P0001  = ~\ACVQN1_reg/NET0131  ;
  assign \ACVQN2_reg/P0001  = ~\ACVQN2_reg/NET0131  ;
  assign \ACVQN3_reg/P0001  = ~\ACVQN3_reg/NET0131  ;
  assign \CNTVCON2_pad  = ~n22 ;
  assign \MRVQN0_reg/P0001  = ~\MRVQN0_reg/NET0131  ;
  assign \P1_pad  = ~\MRVQN1_reg/NET0131  ;
  assign \P2_pad  = ~\MRVQN2_reg/NET0131  ;
  assign \P3_pad  = ~\MRVQN3_reg/NET0131  ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g12/_0_  = n23 ;
  assign \g20/_0_  = ~n49 ;
  assign \g31/_0_  = ~n55 ;
  assign \g616/_0_  = n60 ;
  assign \g630/_0_  = n63 ;
  assign \g632/_0_  = ~n72 ;
  assign \g633/_0_  = n73 ;
  assign \g636/_0_  = ~n79 ;
  assign \g637/_0_  = ~n85 ;
  assign \g638/_0_  = ~n91 ;
  assign \g673/_1__syn_2  = n25 ;
  assign \g675/_1_  = n22 ;
  assign \g795/_0_  = ~n99 ;
  assign \g810/_0_  = ~n107 ;
endmodule
