module top (\100(38)_pad , \103(39)_pad , \106(40)_pad , \109(41)_pad , \11(2)_pad , \112(42)_pad , \113(43)_pad , \114(44)_pad , \115(45)_pad , \116(46)_pad , \117(47)_pad , \118(48)_pad , \119(49)_pad , \120(50)_pad , \121(51)_pad , \122(52)_pad , \123(53)_pad , \126(54)_pad , \127(55)_pad , \128(56)_pad , \129(57)_pad , \130(58)_pad , \131(59)_pad , \132(60)_pad , \135(61)_pad , \136(62)_pad , \14(3)_pad , \140(64)_pad , \144(354)_pad , \145(66)_pad , \146(67)_pad , \149(68)_pad , \1497(156)_pad , \152(69)_pad , \155(70)_pad , \158(71)_pad , \161(72)_pad , \164(73)_pad , \167(74)_pad , \1689(157)_pad , \1690(158)_pad , \1691(159)_pad , \1694(160)_pad , \17(4)_pad , \170(75)_pad , \173(76)_pad , \176(77)_pad , \179(78)_pad , \182(79)_pad , \185(80)_pad , \188(81)_pad , \191(82)_pad , \194(83)_pad , \197(84)_pad , \20(5)_pad , \200(85)_pad , \203(86)_pad , \206(87)_pad , \209(88)_pad , \210(89)_pad , \217(90)_pad , \2174(161)_pad , \218(91)_pad , \225(92)_pad , \226(93)_pad , \23(6)_pad , \233(94)_pad , \234(95)_pad , \2358(162)_pad , \24(7)_pad , \241(96)_pad , \242(97)_pad , \245(98)_pad , \248(99)_pad , \25(8)_pad , \251(100)_pad , \254(101)_pad , \257(102)_pad , \26(9)_pad , \264(103)_pad , \265(104)_pad , \27(10)_pad , \272(105)_pad , \273(106)_pad , \280(107)_pad , \281(108)_pad , \2824(163)_pad , \288(109)_pad , \289(110)_pad , \292(111)_pad , \298(299)_pad , \302(114)_pad , \307(115)_pad , \308(116)_pad , \31(11)_pad , \315(117)_pad , \316(118)_pad , \323(119)_pad , \324(120)_pad , \331(121)_pad , \332(122)_pad , \335(123)_pad , \338(124)_pad , \34(12)_pad , \341(125)_pad , \348(126)_pad , \351(127)_pad , \3546(165)_pad , \3548(166)_pad , \3550(167)_pad , \3552(168)_pad , \358(128)_pad , \361(129)_pad , \366(130)_pad , \369(131)_pad , \37(13)_pad , \3717(169)_pad , \372(132)_pad , \3724(170)_pad , \373(133)_pad , \374(134)_pad , \386(135)_pad , \389(136)_pad , \4(1)_pad , \40(14)_pad , \400(137)_pad , \4087(171)_pad , \4088(172)_pad , \4089(173)_pad , \4090(174)_pad , \4091(175)_pad , \4092(176)_pad , \411(138)_pad , \4115(177)_pad , \422(139)_pad , \43(15)_pad , \435(140)_pad , \446(141)_pad , \457(142)_pad , \46(16)_pad , \468(143)_pad , \479(144)_pad , \49(17)_pad , \490(145)_pad , \503(146)_pad , \514(147)_pad , \52(18)_pad , \523(148)_pad , \53(19)_pad , \534(149)_pad , \54(20)_pad , \545(150)_pad , \552(152)_pad , \556(153)_pad , \559(154)_pad , \562(155)_pad , \61(21)_pad , \64(22)_pad , \67(23)_pad , \70(24)_pad , \73(25)_pad , \76(26)_pad , \79(27)_pad , \80(28)_pad , \81(29)_pad , \82(30)_pad , \83(31)_pad , \86(32)_pad , \87(33)_pad , \88(34)_pad , \889(734)_pad , \892(408)_pad , \91(35)_pad , \926(624)_pad , \94(36)_pad , \97(37)_pad , \973(202)_pad , \993(850)_pad , \1000(2168)_pad , \1002(1920)_pad , \1004(1977)_pad , \588(1696)_pad , \593(733)_pad , \598(1623)_pad , \599(269)_pad , \600(259)_pad , \601(220)_pad , \604(223)_pad , \606(407)_pad , \611(275)_pad , \612(263)_pad , \615(1750)_pad , \618(1925)_pad , \621(1893)_pad , \626(1752)_pad , \632(1692)_pad , \634(665)_pad , \636(1280)_pad , \639(1275)_pad , \642(2222)_pad , \645(2271)_pad , \648(2295)_pad , \651(2314)_pad , \654(2315)_pad , \656(621)_pad , \658(2483)_pad , \661(2178)_pad , \664(2223)_pad , \667(2224)_pad , \670(2225)_pad , \673(1276)_pad , \676(2229)_pad , \679(2272)_pad , \682(2296)_pad , \685(2316)_pad , \688(2317)_pad , \690(2484)_pad , \693(2179)_pad , \696(2226)_pad , \699(2227)_pad , \702(2228)_pad , \704(1281)_pad , \707(1277)_pad , \712(2297)_pad , \715(1278)_pad , \722(2131)_pad , \727(2298)_pad , \732(2300)_pad , \737(2279)_pad , \742(2238)_pad , \747(2187)_pad , \752(2189)_pad , \757(2190)_pad , \762(2184)_pad , \767(2479)_pad , \772(2299)_pad , \777(2278)_pad , \782(2239)_pad , \787(2186)_pad , \792(2188)_pad , \797(2191)_pad , \802(2183)_pad , \807(2480)_pad , \809(655)_pad , \810(356)_pad , \813(2260)_pad , \815(627)_pad , \820(1283)_pad , \822(1933)_pad , \824(2274)_pad , \826(2275)_pad , \828(2233)_pad , \830(2182)_pad , \832(2133)_pad , \834(2123)_pad , \836(2128)_pad , \838(2064)_pad , \843(2455)_pad , \845(845)_pad , \847(465)_pad , \848(330)_pad , \849(219)_pad , \850(217)_pad , \851(218)_pad , \854(2268)_pad , \859(2132)_pad , \861(2070)_pad , \863(2276)_pad , \865(2277)_pad , \867(2237)_pad , \869(2181)_pad , \871(2127)_pad , \873(2124)_pad , \875(2125)_pad , \877(2126)_pad , \882(2456)_pad , \998(2163)_pad , \u2023_syn_3 , \u2095_syn_3 , \u2109_syn_3 , \u2318_syn_3 , \u3086_syn_3 );
	input \100(38)_pad  ;
	input \103(39)_pad  ;
	input \106(40)_pad  ;
	input \109(41)_pad  ;
	input \11(2)_pad  ;
	input \112(42)_pad  ;
	input \113(43)_pad  ;
	input \114(44)_pad  ;
	input \115(45)_pad  ;
	input \116(46)_pad  ;
	input \117(47)_pad  ;
	input \118(48)_pad  ;
	input \119(49)_pad  ;
	input \120(50)_pad  ;
	input \121(51)_pad  ;
	input \122(52)_pad  ;
	input \123(53)_pad  ;
	input \126(54)_pad  ;
	input \127(55)_pad  ;
	input \128(56)_pad  ;
	input \129(57)_pad  ;
	input \130(58)_pad  ;
	input \131(59)_pad  ;
	input \132(60)_pad  ;
	input \135(61)_pad  ;
	input \136(62)_pad  ;
	input \14(3)_pad  ;
	input \140(64)_pad  ;
	input \144(354)_pad  ;
	input \145(66)_pad  ;
	input \146(67)_pad  ;
	input \149(68)_pad  ;
	input \1497(156)_pad  ;
	input \152(69)_pad  ;
	input \155(70)_pad  ;
	input \158(71)_pad  ;
	input \161(72)_pad  ;
	input \164(73)_pad  ;
	input \167(74)_pad  ;
	input \1689(157)_pad  ;
	input \1690(158)_pad  ;
	input \1691(159)_pad  ;
	input \1694(160)_pad  ;
	input \17(4)_pad  ;
	input \170(75)_pad  ;
	input \173(76)_pad  ;
	input \176(77)_pad  ;
	input \179(78)_pad  ;
	input \182(79)_pad  ;
	input \185(80)_pad  ;
	input \188(81)_pad  ;
	input \191(82)_pad  ;
	input \194(83)_pad  ;
	input \197(84)_pad  ;
	input \20(5)_pad  ;
	input \200(85)_pad  ;
	input \203(86)_pad  ;
	input \206(87)_pad  ;
	input \209(88)_pad  ;
	input \210(89)_pad  ;
	input \217(90)_pad  ;
	input \2174(161)_pad  ;
	input \218(91)_pad  ;
	input \225(92)_pad  ;
	input \226(93)_pad  ;
	input \23(6)_pad  ;
	input \233(94)_pad  ;
	input \234(95)_pad  ;
	input \2358(162)_pad  ;
	input \24(7)_pad  ;
	input \241(96)_pad  ;
	input \242(97)_pad  ;
	input \245(98)_pad  ;
	input \248(99)_pad  ;
	input \25(8)_pad  ;
	input \251(100)_pad  ;
	input \254(101)_pad  ;
	input \257(102)_pad  ;
	input \26(9)_pad  ;
	input \264(103)_pad  ;
	input \265(104)_pad  ;
	input \27(10)_pad  ;
	input \272(105)_pad  ;
	input \273(106)_pad  ;
	input \280(107)_pad  ;
	input \281(108)_pad  ;
	input \2824(163)_pad  ;
	input \288(109)_pad  ;
	input \289(110)_pad  ;
	input \292(111)_pad  ;
	input \298(299)_pad  ;
	input \302(114)_pad  ;
	input \307(115)_pad  ;
	input \308(116)_pad  ;
	input \31(11)_pad  ;
	input \315(117)_pad  ;
	input \316(118)_pad  ;
	input \323(119)_pad  ;
	input \324(120)_pad  ;
	input \331(121)_pad  ;
	input \332(122)_pad  ;
	input \335(123)_pad  ;
	input \338(124)_pad  ;
	input \34(12)_pad  ;
	input \341(125)_pad  ;
	input \348(126)_pad  ;
	input \351(127)_pad  ;
	input \3546(165)_pad  ;
	input \3548(166)_pad  ;
	input \3550(167)_pad  ;
	input \3552(168)_pad  ;
	input \358(128)_pad  ;
	input \361(129)_pad  ;
	input \366(130)_pad  ;
	input \369(131)_pad  ;
	input \37(13)_pad  ;
	input \3717(169)_pad  ;
	input \372(132)_pad  ;
	input \3724(170)_pad  ;
	input \373(133)_pad  ;
	input \374(134)_pad  ;
	input \386(135)_pad  ;
	input \389(136)_pad  ;
	input \4(1)_pad  ;
	input \40(14)_pad  ;
	input \400(137)_pad  ;
	input \4087(171)_pad  ;
	input \4088(172)_pad  ;
	input \4089(173)_pad  ;
	input \4090(174)_pad  ;
	input \4091(175)_pad  ;
	input \4092(176)_pad  ;
	input \411(138)_pad  ;
	input \4115(177)_pad  ;
	input \422(139)_pad  ;
	input \43(15)_pad  ;
	input \435(140)_pad  ;
	input \446(141)_pad  ;
	input \457(142)_pad  ;
	input \46(16)_pad  ;
	input \468(143)_pad  ;
	input \479(144)_pad  ;
	input \49(17)_pad  ;
	input \490(145)_pad  ;
	input \503(146)_pad  ;
	input \514(147)_pad  ;
	input \52(18)_pad  ;
	input \523(148)_pad  ;
	input \53(19)_pad  ;
	input \534(149)_pad  ;
	input \54(20)_pad  ;
	input \545(150)_pad  ;
	input \552(152)_pad  ;
	input \556(153)_pad  ;
	input \559(154)_pad  ;
	input \562(155)_pad  ;
	input \61(21)_pad  ;
	input \64(22)_pad  ;
	input \67(23)_pad  ;
	input \70(24)_pad  ;
	input \73(25)_pad  ;
	input \76(26)_pad  ;
	input \79(27)_pad  ;
	input \80(28)_pad  ;
	input \81(29)_pad  ;
	input \82(30)_pad  ;
	input \83(31)_pad  ;
	input \86(32)_pad  ;
	input \87(33)_pad  ;
	input \88(34)_pad  ;
	input \889(734)_pad  ;
	input \892(408)_pad  ;
	input \91(35)_pad  ;
	input \926(624)_pad  ;
	input \94(36)_pad  ;
	input \97(37)_pad  ;
	input \973(202)_pad  ;
	input \993(850)_pad  ;
	output \1000(2168)_pad  ;
	output \1002(1920)_pad  ;
	output \1004(1977)_pad  ;
	output \588(1696)_pad  ;
	output \593(733)_pad  ;
	output \598(1623)_pad  ;
	output \599(269)_pad  ;
	output \600(259)_pad  ;
	output \601(220)_pad  ;
	output \604(223)_pad  ;
	output \606(407)_pad  ;
	output \611(275)_pad  ;
	output \612(263)_pad  ;
	output \615(1750)_pad  ;
	output \618(1925)_pad  ;
	output \621(1893)_pad  ;
	output \626(1752)_pad  ;
	output \632(1692)_pad  ;
	output \634(665)_pad  ;
	output \636(1280)_pad  ;
	output \639(1275)_pad  ;
	output \642(2222)_pad  ;
	output \645(2271)_pad  ;
	output \648(2295)_pad  ;
	output \651(2314)_pad  ;
	output \654(2315)_pad  ;
	output \656(621)_pad  ;
	output \658(2483)_pad  ;
	output \661(2178)_pad  ;
	output \664(2223)_pad  ;
	output \667(2224)_pad  ;
	output \670(2225)_pad  ;
	output \673(1276)_pad  ;
	output \676(2229)_pad  ;
	output \679(2272)_pad  ;
	output \682(2296)_pad  ;
	output \685(2316)_pad  ;
	output \688(2317)_pad  ;
	output \690(2484)_pad  ;
	output \693(2179)_pad  ;
	output \696(2226)_pad  ;
	output \699(2227)_pad  ;
	output \702(2228)_pad  ;
	output \704(1281)_pad  ;
	output \707(1277)_pad  ;
	output \712(2297)_pad  ;
	output \715(1278)_pad  ;
	output \722(2131)_pad  ;
	output \727(2298)_pad  ;
	output \732(2300)_pad  ;
	output \737(2279)_pad  ;
	output \742(2238)_pad  ;
	output \747(2187)_pad  ;
	output \752(2189)_pad  ;
	output \757(2190)_pad  ;
	output \762(2184)_pad  ;
	output \767(2479)_pad  ;
	output \772(2299)_pad  ;
	output \777(2278)_pad  ;
	output \782(2239)_pad  ;
	output \787(2186)_pad  ;
	output \792(2188)_pad  ;
	output \797(2191)_pad  ;
	output \802(2183)_pad  ;
	output \807(2480)_pad  ;
	output \809(655)_pad  ;
	output \810(356)_pad  ;
	output \813(2260)_pad  ;
	output \815(627)_pad  ;
	output \820(1283)_pad  ;
	output \822(1933)_pad  ;
	output \824(2274)_pad  ;
	output \826(2275)_pad  ;
	output \828(2233)_pad  ;
	output \830(2182)_pad  ;
	output \832(2133)_pad  ;
	output \834(2123)_pad  ;
	output \836(2128)_pad  ;
	output \838(2064)_pad  ;
	output \843(2455)_pad  ;
	output \845(845)_pad  ;
	output \847(465)_pad  ;
	output \848(330)_pad  ;
	output \849(219)_pad  ;
	output \850(217)_pad  ;
	output \851(218)_pad  ;
	output \854(2268)_pad  ;
	output \859(2132)_pad  ;
	output \861(2070)_pad  ;
	output \863(2276)_pad  ;
	output \865(2277)_pad  ;
	output \867(2237)_pad  ;
	output \869(2181)_pad  ;
	output \871(2127)_pad  ;
	output \873(2124)_pad  ;
	output \875(2125)_pad  ;
	output \877(2126)_pad  ;
	output \882(2456)_pad  ;
	output \998(2163)_pad  ;
	output \u2023_syn_3  ;
	output \u2095_syn_3  ;
	output \u2109_syn_3  ;
	output \u2318_syn_3  ;
	output \u3086_syn_3  ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\233(94)_pad ,
		\335(123)_pad ,
		_w179_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		\226(93)_pad ,
		\335(123)_pad ,
		_w180_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w179_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\264(103)_pad ,
		\335(123)_pad ,
		_w182_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\257(102)_pad ,
		\335(123)_pad ,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		_w182_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		\280(107)_pad ,
		\335(123)_pad ,
		_w185_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		\273(106)_pad ,
		\335(123)_pad ,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w185_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w184_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		_w184_,
		_w187_,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		_w188_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		_w181_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		_w181_,
		_w190_,
		_w192_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w191_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\241(96)_pad ,
		\335(123)_pad ,
		_w194_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\234(95)_pad ,
		\335(123)_pad ,
		_w195_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w194_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		\288(109)_pad ,
		\335(123)_pad ,
		_w197_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		\281(108)_pad ,
		\335(123)_pad ,
		_w198_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w197_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		_w196_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		_w196_,
		_w199_,
		_w201_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w200_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\272(105)_pad ,
		\335(123)_pad ,
		_w203_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		\265(104)_pad ,
		\335(123)_pad ,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w203_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		\217(90)_pad ,
		\335(123)_pad ,
		_w206_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		\210(89)_pad ,
		\335(123)_pad ,
		_w207_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		_w206_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w205_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w205_,
		_w208_,
		_w210_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		_w209_,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		\292(111)_pad ,
		\335(123)_pad ,
		_w212_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		\289(110)_pad ,
		\335(123)_pad ,
		_w213_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		_w212_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h2)
	) name36 (
		_w211_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		_w211_,
		_w214_,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		_w215_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w202_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		_w202_,
		_w217_,
		_w219_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w218_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		\225(92)_pad ,
		\335(123)_pad ,
		_w221_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		\218(91)_pad ,
		\335(123)_pad ,
		_w222_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w221_,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		\209(88)_pad ,
		\335(123)_pad ,
		_w224_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		\206(87)_pad ,
		\335(123)_pad ,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w224_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		_w223_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		_w223_,
		_w226_,
		_w228_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		_w227_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h2)
	) name51 (
		_w220_,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		_w220_,
		_w229_,
		_w231_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		_w230_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		_w193_,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w193_,
		_w232_,
		_w234_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		_w233_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		\316(118)_pad ,
		\369(131)_pad ,
		_w236_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		\316(118)_pad ,
		\369(131)_pad ,
		_w237_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w236_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		\324(120)_pad ,
		\341(125)_pad ,
		_w239_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		\324(120)_pad ,
		\341(125)_pad ,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		_w239_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		_w238_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		_w238_,
		_w241_,
		_w243_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		_w242_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\308(116)_pad ,
		\361(129)_pad ,
		_w245_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		\308(116)_pad ,
		\361(129)_pad ,
		_w246_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		_w245_,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		\298(299)_pad ,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		\298(299)_pad ,
		_w247_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w248_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		\302(114)_pad ,
		\351(127)_pad ,
		_w251_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		\302(114)_pad ,
		\351(127)_pad ,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w251_,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h2)
	) name75 (
		_w250_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		_w250_,
		_w253_,
		_w255_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		_w254_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w244_,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		_w244_,
		_w256_,
		_w258_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		_w257_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		\218(91)_pad ,
		\281(108)_pad ,
		_w260_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		\218(91)_pad ,
		\281(108)_pad ,
		_w261_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w260_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		\206(87)_pad ,
		\289(110)_pad ,
		_w263_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		\206(87)_pad ,
		\289(110)_pad ,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		_w263_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h2)
	) name87 (
		_w262_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		_w262_,
		_w265_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		_w266_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		\257(102)_pad ,
		\265(104)_pad ,
		_w269_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		\257(102)_pad ,
		\265(104)_pad ,
		_w270_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		_w269_,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		\210(89)_pad ,
		\273(106)_pad ,
		_w272_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		\210(89)_pad ,
		\273(106)_pad ,
		_w273_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w272_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		_w271_,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w271_,
		_w274_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		_w275_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h2)
	) name99 (
		\226(93)_pad ,
		\234(95)_pad ,
		_w278_
	);
	LUT2 #(
		.INIT('h4)
	) name100 (
		\226(93)_pad ,
		\234(95)_pad ,
		_w279_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w278_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		_w277_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		_w277_,
		_w280_,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		_w281_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		_w268_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w268_,
		_w283_,
		_w285_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		_w284_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h2)
	) name108 (
		\422(139)_pad ,
		_w181_,
		_w287_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		\468(143)_pad ,
		_w223_,
		_w288_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		\468(143)_pad ,
		_w223_,
		_w289_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		_w288_,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		\422(139)_pad ,
		_w181_,
		_w291_
	);
	LUT2 #(
		.INIT('h2)
	) name113 (
		_w290_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h4)
	) name114 (
		_w287_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		\374(134)_pad ,
		_w199_,
		_w294_
	);
	LUT2 #(
		.INIT('h4)
	) name116 (
		\374(134)_pad ,
		_w199_,
		_w295_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		_w294_,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h2)
	) name118 (
		\411(138)_pad ,
		_w187_,
		_w297_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		\411(138)_pad ,
		_w187_,
		_w298_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		_w297_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h2)
	) name121 (
		\400(137)_pad ,
		_w205_,
		_w300_
	);
	LUT2 #(
		.INIT('h4)
	) name122 (
		\400(137)_pad ,
		_w205_,
		_w301_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w300_,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w299_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		_w296_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h2)
	) name126 (
		\435(140)_pad ,
		_w196_,
		_w305_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		\435(140)_pad ,
		_w196_,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		_w305_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h2)
	) name129 (
		\389(136)_pad ,
		_w184_,
		_w308_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		\389(136)_pad ,
		_w184_,
		_w309_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w308_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w307_,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		_w304_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h2)
	) name134 (
		\446(141)_pad ,
		_w226_,
		_w313_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		\446(141)_pad ,
		_w226_,
		_w314_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		_w313_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h2)
	) name137 (
		\457(142)_pad ,
		_w208_,
		_w316_
	);
	LUT2 #(
		.INIT('h4)
	) name138 (
		\457(142)_pad ,
		_w208_,
		_w317_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		_w316_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		_w315_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		_w293_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		_w312_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		\251(100)_pad ,
		\316(118)_pad ,
		_w322_
	);
	LUT2 #(
		.INIT('h4)
	) name144 (
		\248(99)_pad ,
		\316(118)_pad ,
		_w323_
	);
	LUT2 #(
		.INIT('h2)
	) name145 (
		\490(145)_pad ,
		_w322_,
		_w324_
	);
	LUT2 #(
		.INIT('h4)
	) name146 (
		_w323_,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h2)
	) name147 (
		\254(101)_pad ,
		\316(118)_pad ,
		_w326_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\242(97)_pad ,
		\316(118)_pad ,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		\490(145)_pad ,
		_w326_,
		_w328_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		_w327_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w325_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		\251(100)_pad ,
		\308(116)_pad ,
		_w331_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		\248(99)_pad ,
		\308(116)_pad ,
		_w332_
	);
	LUT2 #(
		.INIT('h2)
	) name154 (
		\479(144)_pad ,
		_w331_,
		_w333_
	);
	LUT2 #(
		.INIT('h4)
	) name155 (
		_w332_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h2)
	) name156 (
		\254(101)_pad ,
		\308(116)_pad ,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		\242(97)_pad ,
		\308(116)_pad ,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		\479(144)_pad ,
		_w335_,
		_w337_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		_w336_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		_w334_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		_w330_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h2)
	) name162 (
		\251(100)_pad ,
		\361(129)_pad ,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		\248(99)_pad ,
		\361(129)_pad ,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		_w341_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h4)
	) name165 (
		\341(125)_pad ,
		\3550(167)_pad ,
		_w344_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		\341(125)_pad ,
		\3552(168)_pad ,
		_w345_
	);
	LUT2 #(
		.INIT('h2)
	) name167 (
		\523(148)_pad ,
		_w344_,
		_w346_
	);
	LUT2 #(
		.INIT('h4)
	) name168 (
		_w345_,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		\341(125)_pad ,
		\3548(166)_pad ,
		_w348_
	);
	LUT2 #(
		.INIT('h2)
	) name170 (
		\341(125)_pad ,
		\3546(165)_pad ,
		_w349_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		\523(148)_pad ,
		_w348_,
		_w350_
	);
	LUT2 #(
		.INIT('h4)
	) name172 (
		_w349_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		_w347_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h4)
	) name174 (
		\324(120)_pad ,
		\3550(167)_pad ,
		_w353_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		\324(120)_pad ,
		\3552(168)_pad ,
		_w354_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		\503(146)_pad ,
		_w353_,
		_w355_
	);
	LUT2 #(
		.INIT('h4)
	) name177 (
		_w354_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		\324(120)_pad ,
		\3548(166)_pad ,
		_w357_
	);
	LUT2 #(
		.INIT('h2)
	) name179 (
		\324(120)_pad ,
		\3546(165)_pad ,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		\503(146)_pad ,
		_w357_,
		_w359_
	);
	LUT2 #(
		.INIT('h4)
	) name181 (
		_w358_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		_w356_,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h4)
	) name183 (
		\351(127)_pad ,
		\3550(167)_pad ,
		_w362_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		\351(127)_pad ,
		\3552(168)_pad ,
		_w363_
	);
	LUT2 #(
		.INIT('h2)
	) name185 (
		\534(149)_pad ,
		_w362_,
		_w364_
	);
	LUT2 #(
		.INIT('h4)
	) name186 (
		_w363_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		\351(127)_pad ,
		\3548(166)_pad ,
		_w366_
	);
	LUT2 #(
		.INIT('h2)
	) name188 (
		\351(127)_pad ,
		\3546(165)_pad ,
		_w367_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		\534(149)_pad ,
		_w366_,
		_w368_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		_w367_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		_w365_,
		_w369_,
		_w370_
	);
	LUT2 #(
		.INIT('h2)
	) name192 (
		\254(101)_pad ,
		\298(299)_pad ,
		_w371_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		\242(97)_pad ,
		\298(299)_pad ,
		_w372_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		_w371_,
		_w372_,
		_w373_
	);
	LUT2 #(
		.INIT('h2)
	) name195 (
		\251(100)_pad ,
		\302(114)_pad ,
		_w374_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\248(99)_pad ,
		\302(114)_pad ,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		_w374_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h2)
	) name198 (
		_w373_,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		\3552(168)_pad ,
		\514(147)_pad ,
		_w378_
	);
	LUT2 #(
		.INIT('h2)
	) name200 (
		\3546(165)_pad ,
		\514(147)_pad ,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		_w378_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		_w343_,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		_w377_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		_w352_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		_w361_,
		_w370_,
		_w384_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		_w383_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		_w340_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		\552(152)_pad ,
		\562(155)_pad ,
		_w387_
	);
	LUT2 #(
		.INIT('h2)
	) name209 (
		\332(122)_pad ,
		\338(124)_pad ,
		_w388_
	);
	LUT2 #(
		.INIT('h4)
	) name210 (
		\514(147)_pad ,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		\514(147)_pad ,
		_w388_,
		_w390_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		_w389_,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		\332(122)_pad ,
		\348(126)_pad ,
		_w392_
	);
	LUT2 #(
		.INIT('h4)
	) name214 (
		\332(122)_pad ,
		\341(125)_pad ,
		_w393_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		_w392_,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h2)
	) name216 (
		\523(148)_pad ,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		\523(148)_pad ,
		_w394_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w395_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		\332(122)_pad ,
		\358(128)_pad ,
		_w398_
	);
	LUT2 #(
		.INIT('h4)
	) name220 (
		\332(122)_pad ,
		\351(127)_pad ,
		_w399_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		_w398_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		\534(149)_pad ,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h4)
	) name223 (
		\534(149)_pad ,
		_w400_,
		_w402_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w401_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		_w397_,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		\332(122)_pad ,
		\366(130)_pad ,
		_w405_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		\332(122)_pad ,
		\361(129)_pad ,
		_w406_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		_w405_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		_w404_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w391_,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		\324(120)_pad ,
		\332(122)_pad ,
		_w410_
	);
	LUT2 #(
		.INIT('h4)
	) name232 (
		\331(121)_pad ,
		\332(122)_pad ,
		_w411_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		_w410_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		\503(146)_pad ,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		\503(146)_pad ,
		_w412_,
		_w414_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		_w413_,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		_w409_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		\332(122)_pad ,
		\889(734)_pad ,
		_w417_
	);
	LUT2 #(
		.INIT('h2)
	) name239 (
		\298(299)_pad ,
		\332(122)_pad ,
		_w418_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		_w417_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		\307(115)_pad ,
		\332(122)_pad ,
		_w420_
	);
	LUT2 #(
		.INIT('h2)
	) name242 (
		\302(114)_pad ,
		\332(122)_pad ,
		_w421_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		_w420_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		_w419_,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		\315(117)_pad ,
		\332(122)_pad ,
		_w424_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		\308(116)_pad ,
		\332(122)_pad ,
		_w425_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		_w424_,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h2)
	) name248 (
		\479(144)_pad ,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h4)
	) name249 (
		\479(144)_pad ,
		_w426_,
		_w428_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		_w427_,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h8)
	) name251 (
		\323(119)_pad ,
		\332(122)_pad ,
		_w430_
	);
	LUT2 #(
		.INIT('h2)
	) name252 (
		\316(118)_pad ,
		\332(122)_pad ,
		_w431_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w430_,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h2)
	) name254 (
		\490(145)_pad ,
		_w432_,
		_w433_
	);
	LUT2 #(
		.INIT('h4)
	) name255 (
		\490(145)_pad ,
		_w432_,
		_w434_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		_w433_,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		_w429_,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		_w423_,
		_w436_,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		_w416_,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		_w429_,
		_w433_,
		_w439_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w427_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w402_,
		_w407_,
		_w441_
	);
	LUT2 #(
		.INIT('h1)
	) name263 (
		_w395_,
		_w401_,
		_w442_
	);
	LUT2 #(
		.INIT('h4)
	) name264 (
		_w441_,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		_w396_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h1)
	) name266 (
		_w390_,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		_w389_,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w413_,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		_w414_,
		_w447_,
		_w448_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		_w437_,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		_w423_,
		_w440_,
		_w450_
	);
	LUT2 #(
		.INIT('h4)
	) name272 (
		_w449_,
		_w450_,
		_w451_
	);
	LUT2 #(
		.INIT('h8)
	) name273 (
		_w287_,
		_w290_,
		_w452_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		_w288_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h4)
	) name275 (
		_w316_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h2)
	) name276 (
		_w294_,
		_w298_,
		_w455_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		_w297_,
		_w300_,
		_w456_
	);
	LUT2 #(
		.INIT('h4)
	) name278 (
		_w455_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		_w301_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h4)
	) name280 (
		_w309_,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w308_,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		_w305_,
		_w460_,
		_w461_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		_w306_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h8)
	) name284 (
		_w293_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h2)
	) name285 (
		_w454_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		_w314_,
		_w317_,
		_w465_
	);
	LUT2 #(
		.INIT('h4)
	) name287 (
		_w464_,
		_w465_,
		_w466_
	);
	LUT2 #(
		.INIT('h1)
	) name288 (
		_w313_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h8)
	) name289 (
		\373(133)_pad ,
		\993(850)_pad ,
		_w468_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		\27(10)_pad ,
		\31(11)_pad ,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		\2358(162)_pad ,
		\86(32)_pad ,
		_w470_
	);
	LUT2 #(
		.INIT('h2)
	) name292 (
		\2358(162)_pad ,
		\87(33)_pad ,
		_w471_
	);
	LUT2 #(
		.INIT('h2)
	) name293 (
		_w469_,
		_w470_,
		_w472_
	);
	LUT2 #(
		.INIT('h4)
	) name294 (
		_w471_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h4)
	) name295 (
		\2358(162)_pad ,
		\24(7)_pad ,
		_w474_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		\2358(162)_pad ,
		\25(8)_pad ,
		_w475_
	);
	LUT2 #(
		.INIT('h2)
	) name297 (
		_w469_,
		_w474_,
		_w476_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		_w475_,
		_w476_,
		_w477_
	);
	LUT2 #(
		.INIT('h2)
	) name299 (
		\144(354)_pad ,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h2)
	) name300 (
		\1689(157)_pad ,
		\1690(158)_pad ,
		_w479_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w480_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		\234(95)_pad ,
		\3550(167)_pad ,
		_w481_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		\234(95)_pad ,
		\3552(168)_pad ,
		_w482_
	);
	LUT2 #(
		.INIT('h2)
	) name304 (
		\435(140)_pad ,
		_w481_,
		_w483_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		_w482_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		\234(95)_pad ,
		\3548(166)_pad ,
		_w485_
	);
	LUT2 #(
		.INIT('h2)
	) name307 (
		\234(95)_pad ,
		\3546(165)_pad ,
		_w486_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		\435(140)_pad ,
		_w485_,
		_w487_
	);
	LUT2 #(
		.INIT('h4)
	) name309 (
		_w486_,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		_w484_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h8)
	) name311 (
		_w480_,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('h2)
	) name312 (
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w491_
	);
	LUT2 #(
		.INIT('h8)
	) name313 (
		\4(1)_pad ,
		_w304_,
		_w492_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		_w310_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h2)
	) name315 (
		_w460_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		_w307_,
		_w494_,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w307_,
		_w494_,
		_w496_
	);
	LUT2 #(
		.INIT('h1)
	) name318 (
		_w495_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h2)
	) name319 (
		_w491_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h4)
	) name320 (
		\4091(175)_pad ,
		\4092(176)_pad ,
		_w499_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		\122(52)_pad ,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h1)
	) name322 (
		_w490_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h4)
	) name323 (
		_w498_,
		_w501_,
		_w502_
	);
	LUT2 #(
		.INIT('h2)
	) name324 (
		_w479_,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		\1689(157)_pad ,
		\1690(158)_pad ,
		_w504_
	);
	LUT2 #(
		.INIT('h8)
	) name326 (
		\170(75)_pad ,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h4)
	) name327 (
		\1689(157)_pad ,
		\1690(158)_pad ,
		_w506_
	);
	LUT2 #(
		.INIT('h8)
	) name328 (
		\200(85)_pad ,
		_w506_,
		_w507_
	);
	LUT2 #(
		.INIT('h1)
	) name329 (
		\1689(157)_pad ,
		\1690(158)_pad ,
		_w508_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		_w361_,
		_w480_,
		_w509_
	);
	LUT2 #(
		.INIT('h8)
	) name331 (
		\54(20)_pad ,
		_w408_,
		_w510_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		_w391_,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h1)
	) name333 (
		_w446_,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h2)
	) name334 (
		_w415_,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		_w415_,
		_w512_,
		_w514_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w513_,
		_w514_,
		_w515_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		_w491_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h8)
	) name338 (
		\52(18)_pad ,
		_w499_,
		_w517_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		_w509_,
		_w517_,
		_w518_
	);
	LUT2 #(
		.INIT('h4)
	) name340 (
		_w516_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h2)
	) name341 (
		_w508_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h1)
	) name342 (
		_w505_,
		_w507_,
		_w521_
	);
	LUT2 #(
		.INIT('h4)
	) name343 (
		_w503_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h4)
	) name344 (
		_w520_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h2)
	) name345 (
		\926(624)_pad ,
		_w523_,
		_w524_
	);
	LUT2 #(
		.INIT('h4)
	) name346 (
		\226(93)_pad ,
		\3550(167)_pad ,
		_w525_
	);
	LUT2 #(
		.INIT('h8)
	) name347 (
		\226(93)_pad ,
		\3552(168)_pad ,
		_w526_
	);
	LUT2 #(
		.INIT('h2)
	) name348 (
		\422(139)_pad ,
		_w525_,
		_w527_
	);
	LUT2 #(
		.INIT('h4)
	) name349 (
		_w526_,
		_w527_,
		_w528_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		\226(93)_pad ,
		\3548(166)_pad ,
		_w529_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		\226(93)_pad ,
		\3546(165)_pad ,
		_w530_
	);
	LUT2 #(
		.INIT('h1)
	) name352 (
		\422(139)_pad ,
		_w529_,
		_w531_
	);
	LUT2 #(
		.INIT('h4)
	) name353 (
		_w530_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h1)
	) name354 (
		_w528_,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h8)
	) name355 (
		_w480_,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w287_,
		_w291_,
		_w535_
	);
	LUT2 #(
		.INIT('h2)
	) name357 (
		_w461_,
		_w493_,
		_w536_
	);
	LUT2 #(
		.INIT('h1)
	) name358 (
		_w306_,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h4)
	) name359 (
		_w535_,
		_w537_,
		_w538_
	);
	LUT2 #(
		.INIT('h2)
	) name360 (
		_w535_,
		_w537_,
		_w539_
	);
	LUT2 #(
		.INIT('h1)
	) name361 (
		_w538_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h2)
	) name362 (
		_w491_,
		_w540_,
		_w541_
	);
	LUT2 #(
		.INIT('h8)
	) name363 (
		\113(43)_pad ,
		_w499_,
		_w542_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		_w534_,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w541_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h2)
	) name366 (
		_w479_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h8)
	) name367 (
		\173(76)_pad ,
		_w504_,
		_w546_
	);
	LUT2 #(
		.INIT('h8)
	) name368 (
		\203(86)_pad ,
		_w506_,
		_w547_
	);
	LUT2 #(
		.INIT('h8)
	) name369 (
		_w330_,
		_w480_,
		_w548_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		_w413_,
		_w513_,
		_w549_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w435_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h8)
	) name372 (
		_w435_,
		_w549_,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name373 (
		_w550_,
		_w551_,
		_w552_
	);
	LUT2 #(
		.INIT('h2)
	) name374 (
		_w491_,
		_w552_,
		_w553_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		\112(42)_pad ,
		_w499_,
		_w554_
	);
	LUT2 #(
		.INIT('h1)
	) name376 (
		_w548_,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h4)
	) name377 (
		_w553_,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h2)
	) name378 (
		_w508_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		_w546_,
		_w547_,
		_w558_
	);
	LUT2 #(
		.INIT('h4)
	) name380 (
		_w545_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h4)
	) name381 (
		_w557_,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h2)
	) name382 (
		\926(624)_pad ,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h4)
	) name383 (
		\218(91)_pad ,
		\3550(167)_pad ,
		_w562_
	);
	LUT2 #(
		.INIT('h8)
	) name384 (
		\218(91)_pad ,
		\3552(168)_pad ,
		_w563_
	);
	LUT2 #(
		.INIT('h2)
	) name385 (
		\468(143)_pad ,
		_w562_,
		_w564_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		_w563_,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		\218(91)_pad ,
		\3548(166)_pad ,
		_w566_
	);
	LUT2 #(
		.INIT('h2)
	) name388 (
		\218(91)_pad ,
		\3546(165)_pad ,
		_w567_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		\468(143)_pad ,
		_w566_,
		_w568_
	);
	LUT2 #(
		.INIT('h4)
	) name390 (
		_w567_,
		_w568_,
		_w569_
	);
	LUT2 #(
		.INIT('h1)
	) name391 (
		_w565_,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		_w480_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h8)
	) name393 (
		\53(19)_pad ,
		_w499_,
		_w572_
	);
	LUT2 #(
		.INIT('h4)
	) name394 (
		_w290_,
		_w291_,
		_w573_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		_w292_,
		_w573_,
		_w574_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		_w539_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h8)
	) name397 (
		_w539_,
		_w574_,
		_w576_
	);
	LUT2 #(
		.INIT('h2)
	) name398 (
		_w491_,
		_w575_,
		_w577_
	);
	LUT2 #(
		.INIT('h4)
	) name399 (
		_w576_,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		_w571_,
		_w572_,
		_w579_
	);
	LUT2 #(
		.INIT('h4)
	) name401 (
		_w578_,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h2)
	) name402 (
		_w479_,
		_w580_,
		_w581_
	);
	LUT2 #(
		.INIT('h8)
	) name403 (
		\167(74)_pad ,
		_w504_,
		_w582_
	);
	LUT2 #(
		.INIT('h8)
	) name404 (
		\197(84)_pad ,
		_w506_,
		_w583_
	);
	LUT2 #(
		.INIT('h8)
	) name405 (
		_w339_,
		_w480_,
		_w584_
	);
	LUT2 #(
		.INIT('h8)
	) name406 (
		\116(46)_pad ,
		_w499_,
		_w585_
	);
	LUT2 #(
		.INIT('h2)
	) name407 (
		_w429_,
		_w434_,
		_w586_
	);
	LUT2 #(
		.INIT('h4)
	) name408 (
		_w429_,
		_w434_,
		_w587_
	);
	LUT2 #(
		.INIT('h1)
	) name409 (
		_w586_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		_w551_,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h4)
	) name411 (
		_w429_,
		_w551_,
		_w590_
	);
	LUT2 #(
		.INIT('h2)
	) name412 (
		_w491_,
		_w589_,
		_w591_
	);
	LUT2 #(
		.INIT('h4)
	) name413 (
		_w590_,
		_w591_,
		_w592_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		_w584_,
		_w585_,
		_w593_
	);
	LUT2 #(
		.INIT('h4)
	) name415 (
		_w592_,
		_w593_,
		_w594_
	);
	LUT2 #(
		.INIT('h2)
	) name416 (
		_w508_,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h1)
	) name417 (
		_w582_,
		_w583_,
		_w596_
	);
	LUT2 #(
		.INIT('h4)
	) name418 (
		_w581_,
		_w596_,
		_w597_
	);
	LUT2 #(
		.INIT('h4)
	) name419 (
		_w595_,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h2)
	) name420 (
		\926(624)_pad ,
		_w598_,
		_w599_
	);
	LUT2 #(
		.INIT('h4)
	) name421 (
		\210(89)_pad ,
		\3550(167)_pad ,
		_w600_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		\210(89)_pad ,
		\3552(168)_pad ,
		_w601_
	);
	LUT2 #(
		.INIT('h2)
	) name423 (
		\457(142)_pad ,
		_w600_,
		_w602_
	);
	LUT2 #(
		.INIT('h4)
	) name424 (
		_w601_,
		_w602_,
		_w603_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		\210(89)_pad ,
		\3548(166)_pad ,
		_w604_
	);
	LUT2 #(
		.INIT('h2)
	) name426 (
		\210(89)_pad ,
		\3546(165)_pad ,
		_w605_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		\457(142)_pad ,
		_w604_,
		_w606_
	);
	LUT2 #(
		.INIT('h4)
	) name428 (
		_w605_,
		_w606_,
		_w607_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		_w603_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h8)
	) name430 (
		_w480_,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('h2)
	) name431 (
		_w453_,
		_w537_,
		_w610_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w288_,
		_w292_,
		_w611_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		_w610_,
		_w611_,
		_w612_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		_w318_,
		_w612_,
		_w613_
	);
	LUT2 #(
		.INIT('h1)
	) name435 (
		_w318_,
		_w612_,
		_w614_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		_w613_,
		_w614_,
		_w615_
	);
	LUT2 #(
		.INIT('h8)
	) name437 (
		_w491_,
		_w615_,
		_w616_
	);
	LUT2 #(
		.INIT('h8)
	) name438 (
		\114(44)_pad ,
		_w499_,
		_w617_
	);
	LUT2 #(
		.INIT('h1)
	) name439 (
		_w609_,
		_w617_,
		_w618_
	);
	LUT2 #(
		.INIT('h4)
	) name440 (
		_w616_,
		_w618_,
		_w619_
	);
	LUT2 #(
		.INIT('h2)
	) name441 (
		_w479_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h8)
	) name442 (
		\164(73)_pad ,
		_w504_,
		_w621_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		\194(83)_pad ,
		_w506_,
		_w622_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		_w376_,
		_w480_,
		_w623_
	);
	LUT2 #(
		.INIT('h2)
	) name445 (
		_w436_,
		_w549_,
		_w624_
	);
	LUT2 #(
		.INIT('h2)
	) name446 (
		_w440_,
		_w624_,
		_w625_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		_w422_,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		_w422_,
		_w625_,
		_w627_
	);
	LUT2 #(
		.INIT('h1)
	) name449 (
		_w626_,
		_w627_,
		_w628_
	);
	LUT2 #(
		.INIT('h2)
	) name450 (
		_w491_,
		_w628_,
		_w629_
	);
	LUT2 #(
		.INIT('h8)
	) name451 (
		\121(51)_pad ,
		_w499_,
		_w630_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		_w623_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h4)
	) name453 (
		_w629_,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h2)
	) name454 (
		_w508_,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h1)
	) name455 (
		_w621_,
		_w622_,
		_w634_
	);
	LUT2 #(
		.INIT('h4)
	) name456 (
		_w620_,
		_w634_,
		_w635_
	);
	LUT2 #(
		.INIT('h4)
	) name457 (
		_w633_,
		_w635_,
		_w636_
	);
	LUT2 #(
		.INIT('h2)
	) name458 (
		\926(624)_pad ,
		_w636_,
		_w637_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		\206(87)_pad ,
		\251(100)_pad ,
		_w638_
	);
	LUT2 #(
		.INIT('h2)
	) name460 (
		\206(87)_pad ,
		\248(99)_pad ,
		_w639_
	);
	LUT2 #(
		.INIT('h2)
	) name461 (
		\446(141)_pad ,
		_w638_,
		_w640_
	);
	LUT2 #(
		.INIT('h4)
	) name462 (
		_w639_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h4)
	) name463 (
		\206(87)_pad ,
		\254(101)_pad ,
		_w642_
	);
	LUT2 #(
		.INIT('h8)
	) name464 (
		\206(87)_pad ,
		\242(97)_pad ,
		_w643_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		\446(141)_pad ,
		_w642_,
		_w644_
	);
	LUT2 #(
		.INIT('h4)
	) name466 (
		_w643_,
		_w644_,
		_w645_
	);
	LUT2 #(
		.INIT('h1)
	) name467 (
		_w641_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('h8)
	) name468 (
		_w480_,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h4)
	) name469 (
		_w293_,
		_w454_,
		_w648_
	);
	LUT2 #(
		.INIT('h1)
	) name470 (
		_w317_,
		_w648_,
		_w649_
	);
	LUT2 #(
		.INIT('h2)
	) name471 (
		_w454_,
		_w537_,
		_w650_
	);
	LUT2 #(
		.INIT('h2)
	) name472 (
		_w649_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		_w315_,
		_w651_,
		_w652_
	);
	LUT2 #(
		.INIT('h1)
	) name474 (
		_w315_,
		_w651_,
		_w653_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w652_,
		_w653_,
		_w654_
	);
	LUT2 #(
		.INIT('h8)
	) name476 (
		_w491_,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		\115(45)_pad ,
		_w499_,
		_w656_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		_w647_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h4)
	) name479 (
		_w655_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h2)
	) name480 (
		_w479_,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h8)
	) name481 (
		\161(72)_pad ,
		_w504_,
		_w660_
	);
	LUT2 #(
		.INIT('h8)
	) name482 (
		\191(82)_pad ,
		_w506_,
		_w661_
	);
	LUT2 #(
		.INIT('h4)
	) name483 (
		_w373_,
		_w480_,
		_w662_
	);
	LUT2 #(
		.INIT('h8)
	) name484 (
		\123(53)_pad ,
		_w499_,
		_w663_
	);
	LUT2 #(
		.INIT('h4)
	) name485 (
		_w419_,
		_w627_,
		_w664_
	);
	LUT2 #(
		.INIT('h2)
	) name486 (
		_w419_,
		_w627_,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name487 (
		_w664_,
		_w665_,
		_w666_
	);
	LUT2 #(
		.INIT('h8)
	) name488 (
		_w491_,
		_w666_,
		_w667_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		_w662_,
		_w663_,
		_w668_
	);
	LUT2 #(
		.INIT('h4)
	) name490 (
		_w667_,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h2)
	) name491 (
		_w508_,
		_w669_,
		_w670_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		_w660_,
		_w661_,
		_w671_
	);
	LUT2 #(
		.INIT('h4)
	) name493 (
		_w659_,
		_w671_,
		_w672_
	);
	LUT2 #(
		.INIT('h4)
	) name494 (
		_w670_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h2)
	) name495 (
		\926(624)_pad ,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h8)
	) name496 (
		\140(64)_pad ,
		_w469_,
		_w675_
	);
	LUT2 #(
		.INIT('h8)
	) name497 (
		\4092(176)_pad ,
		\97(37)_pad ,
		_w676_
	);
	LUT2 #(
		.INIT('h1)
	) name498 (
		_w307_,
		_w310_,
		_w677_
	);
	LUT2 #(
		.INIT('h1)
	) name499 (
		_w311_,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		_w294_,
		_w297_,
		_w679_
	);
	LUT2 #(
		.INIT('h1)
	) name501 (
		_w455_,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		_w308_,
		_w458_,
		_w681_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		_w459_,
		_w681_,
		_w682_
	);
	LUT2 #(
		.INIT('h2)
	) name504 (
		_w680_,
		_w682_,
		_w683_
	);
	LUT2 #(
		.INIT('h4)
	) name505 (
		_w680_,
		_w682_,
		_w684_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w683_,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h1)
	) name507 (
		_w296_,
		_w685_,
		_w686_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		_w304_,
		_w458_,
		_w687_
	);
	LUT2 #(
		.INIT('h1)
	) name509 (
		_w309_,
		_w687_,
		_w688_
	);
	LUT2 #(
		.INIT('h4)
	) name510 (
		_w308_,
		_w687_,
		_w689_
	);
	LUT2 #(
		.INIT('h1)
	) name511 (
		_w688_,
		_w689_,
		_w690_
	);
	LUT2 #(
		.INIT('h2)
	) name512 (
		_w295_,
		_w297_,
		_w691_
	);
	LUT2 #(
		.INIT('h1)
	) name513 (
		_w295_,
		_w298_,
		_w692_
	);
	LUT2 #(
		.INIT('h1)
	) name514 (
		_w691_,
		_w692_,
		_w693_
	);
	LUT2 #(
		.INIT('h2)
	) name515 (
		_w690_,
		_w693_,
		_w694_
	);
	LUT2 #(
		.INIT('h4)
	) name516 (
		_w690_,
		_w693_,
		_w695_
	);
	LUT2 #(
		.INIT('h2)
	) name517 (
		_w296_,
		_w694_,
		_w696_
	);
	LUT2 #(
		.INIT('h4)
	) name518 (
		_w695_,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		_w686_,
		_w697_,
		_w698_
	);
	LUT2 #(
		.INIT('h2)
	) name520 (
		\1497(156)_pad ,
		_w698_,
		_w699_
	);
	LUT2 #(
		.INIT('h8)
	) name521 (
		_w296_,
		_w685_,
		_w700_
	);
	LUT2 #(
		.INIT('h1)
	) name522 (
		\1497(156)_pad ,
		_w686_,
		_w701_
	);
	LUT2 #(
		.INIT('h4)
	) name523 (
		_w700_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		_w699_,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h2)
	) name525 (
		_w678_,
		_w703_,
		_w704_
	);
	LUT2 #(
		.INIT('h4)
	) name526 (
		_w678_,
		_w703_,
		_w705_
	);
	LUT2 #(
		.INIT('h1)
	) name527 (
		_w704_,
		_w705_,
		_w706_
	);
	LUT2 #(
		.INIT('h1)
	) name528 (
		_w299_,
		_w302_,
		_w707_
	);
	LUT2 #(
		.INIT('h1)
	) name529 (
		_w303_,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h8)
	) name530 (
		\1497(156)_pad ,
		_w312_,
		_w709_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w462_,
		_w709_,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w317_,
		_w453_,
		_w711_
	);
	LUT2 #(
		.INIT('h1)
	) name533 (
		_w454_,
		_w711_,
		_w712_
	);
	LUT2 #(
		.INIT('h4)
	) name534 (
		_w315_,
		_w712_,
		_w713_
	);
	LUT2 #(
		.INIT('h1)
	) name535 (
		_w315_,
		_w318_,
		_w714_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w319_,
		_w714_,
		_w715_
	);
	LUT2 #(
		.INIT('h4)
	) name537 (
		_w712_,
		_w715_,
		_w716_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		_w713_,
		_w716_,
		_w717_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		_w574_,
		_w717_,
		_w718_
	);
	LUT2 #(
		.INIT('h8)
	) name540 (
		_w574_,
		_w717_,
		_w719_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		_w718_,
		_w719_,
		_w720_
	);
	LUT2 #(
		.INIT('h2)
	) name542 (
		_w710_,
		_w720_,
		_w721_
	);
	LUT2 #(
		.INIT('h1)
	) name543 (
		_w287_,
		_w290_,
		_w722_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		_w452_,
		_w722_,
		_w723_
	);
	LUT2 #(
		.INIT('h8)
	) name545 (
		_w715_,
		_w723_,
		_w724_
	);
	LUT2 #(
		.INIT('h1)
	) name546 (
		_w715_,
		_w723_,
		_w725_
	);
	LUT2 #(
		.INIT('h1)
	) name547 (
		_w724_,
		_w725_,
		_w726_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		_w611_,
		_w649_,
		_w727_
	);
	LUT2 #(
		.INIT('h4)
	) name549 (
		_w293_,
		_w316_,
		_w728_
	);
	LUT2 #(
		.INIT('h8)
	) name550 (
		_w453_,
		_w728_,
		_w729_
	);
	LUT2 #(
		.INIT('h1)
	) name551 (
		_w727_,
		_w729_,
		_w730_
	);
	LUT2 #(
		.INIT('h1)
	) name552 (
		_w726_,
		_w730_,
		_w731_
	);
	LUT2 #(
		.INIT('h8)
	) name553 (
		_w726_,
		_w730_,
		_w732_
	);
	LUT2 #(
		.INIT('h1)
	) name554 (
		_w710_,
		_w731_,
		_w733_
	);
	LUT2 #(
		.INIT('h4)
	) name555 (
		_w732_,
		_w733_,
		_w734_
	);
	LUT2 #(
		.INIT('h1)
	) name556 (
		_w721_,
		_w734_,
		_w735_
	);
	LUT2 #(
		.INIT('h2)
	) name557 (
		_w708_,
		_w735_,
		_w736_
	);
	LUT2 #(
		.INIT('h4)
	) name558 (
		_w708_,
		_w735_,
		_w737_
	);
	LUT2 #(
		.INIT('h1)
	) name559 (
		_w736_,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h4)
	) name560 (
		_w706_,
		_w738_,
		_w739_
	);
	LUT2 #(
		.INIT('h2)
	) name561 (
		_w706_,
		_w738_,
		_w740_
	);
	LUT2 #(
		.INIT('h1)
	) name562 (
		_w739_,
		_w740_,
		_w741_
	);
	LUT2 #(
		.INIT('h8)
	) name563 (
		\4091(175)_pad ,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		\234(95)_pad ,
		\251(100)_pad ,
		_w743_
	);
	LUT2 #(
		.INIT('h2)
	) name565 (
		\234(95)_pad ,
		\248(99)_pad ,
		_w744_
	);
	LUT2 #(
		.INIT('h2)
	) name566 (
		\435(140)_pad ,
		_w743_,
		_w745_
	);
	LUT2 #(
		.INIT('h4)
	) name567 (
		_w744_,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h4)
	) name568 (
		\234(95)_pad ,
		\254(101)_pad ,
		_w747_
	);
	LUT2 #(
		.INIT('h8)
	) name569 (
		\234(95)_pad ,
		\242(97)_pad ,
		_w748_
	);
	LUT2 #(
		.INIT('h1)
	) name570 (
		\435(140)_pad ,
		_w747_,
		_w749_
	);
	LUT2 #(
		.INIT('h4)
	) name571 (
		_w748_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		_w746_,
		_w750_,
		_w751_
	);
	LUT2 #(
		.INIT('h1)
	) name573 (
		\226(93)_pad ,
		\251(100)_pad ,
		_w752_
	);
	LUT2 #(
		.INIT('h2)
	) name574 (
		\226(93)_pad ,
		\248(99)_pad ,
		_w753_
	);
	LUT2 #(
		.INIT('h2)
	) name575 (
		\422(139)_pad ,
		_w752_,
		_w754_
	);
	LUT2 #(
		.INIT('h4)
	) name576 (
		_w753_,
		_w754_,
		_w755_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		\226(93)_pad ,
		\254(101)_pad ,
		_w756_
	);
	LUT2 #(
		.INIT('h8)
	) name578 (
		\226(93)_pad ,
		\242(97)_pad ,
		_w757_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		\422(139)_pad ,
		_w756_,
		_w758_
	);
	LUT2 #(
		.INIT('h4)
	) name580 (
		_w757_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h1)
	) name581 (
		_w755_,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h2)
	) name582 (
		_w751_,
		_w760_,
		_w761_
	);
	LUT2 #(
		.INIT('h4)
	) name583 (
		_w751_,
		_w760_,
		_w762_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		_w761_,
		_w762_,
		_w763_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		\210(89)_pad ,
		\251(100)_pad ,
		_w764_
	);
	LUT2 #(
		.INIT('h2)
	) name586 (
		\210(89)_pad ,
		\248(99)_pad ,
		_w765_
	);
	LUT2 #(
		.INIT('h2)
	) name587 (
		\457(142)_pad ,
		_w764_,
		_w766_
	);
	LUT2 #(
		.INIT('h4)
	) name588 (
		_w765_,
		_w766_,
		_w767_
	);
	LUT2 #(
		.INIT('h4)
	) name589 (
		\210(89)_pad ,
		\254(101)_pad ,
		_w768_
	);
	LUT2 #(
		.INIT('h8)
	) name590 (
		\210(89)_pad ,
		\242(97)_pad ,
		_w769_
	);
	LUT2 #(
		.INIT('h1)
	) name591 (
		\457(142)_pad ,
		_w768_,
		_w770_
	);
	LUT2 #(
		.INIT('h4)
	) name592 (
		_w769_,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('h1)
	) name593 (
		_w767_,
		_w771_,
		_w772_
	);
	LUT2 #(
		.INIT('h4)
	) name594 (
		_w646_,
		_w772_,
		_w773_
	);
	LUT2 #(
		.INIT('h2)
	) name595 (
		_w646_,
		_w772_,
		_w774_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		_w773_,
		_w774_,
		_w775_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		\218(91)_pad ,
		\251(100)_pad ,
		_w776_
	);
	LUT2 #(
		.INIT('h2)
	) name598 (
		\218(91)_pad ,
		\248(99)_pad ,
		_w777_
	);
	LUT2 #(
		.INIT('h2)
	) name599 (
		\468(143)_pad ,
		_w776_,
		_w778_
	);
	LUT2 #(
		.INIT('h4)
	) name600 (
		_w777_,
		_w778_,
		_w779_
	);
	LUT2 #(
		.INIT('h4)
	) name601 (
		\218(91)_pad ,
		\254(101)_pad ,
		_w780_
	);
	LUT2 #(
		.INIT('h8)
	) name602 (
		\218(91)_pad ,
		\242(97)_pad ,
		_w781_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		\468(143)_pad ,
		_w780_,
		_w782_
	);
	LUT2 #(
		.INIT('h4)
	) name604 (
		_w781_,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h1)
	) name605 (
		_w779_,
		_w783_,
		_w784_
	);
	LUT2 #(
		.INIT('h2)
	) name606 (
		_w775_,
		_w784_,
		_w785_
	);
	LUT2 #(
		.INIT('h4)
	) name607 (
		_w775_,
		_w784_,
		_w786_
	);
	LUT2 #(
		.INIT('h1)
	) name608 (
		_w785_,
		_w786_,
		_w787_
	);
	LUT2 #(
		.INIT('h8)
	) name609 (
		_w763_,
		_w787_,
		_w788_
	);
	LUT2 #(
		.INIT('h1)
	) name610 (
		_w763_,
		_w787_,
		_w789_
	);
	LUT2 #(
		.INIT('h1)
	) name611 (
		_w788_,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('h1)
	) name612 (
		\251(100)_pad ,
		\257(102)_pad ,
		_w791_
	);
	LUT2 #(
		.INIT('h4)
	) name613 (
		\248(99)_pad ,
		\257(102)_pad ,
		_w792_
	);
	LUT2 #(
		.INIT('h2)
	) name614 (
		\389(136)_pad ,
		_w791_,
		_w793_
	);
	LUT2 #(
		.INIT('h4)
	) name615 (
		_w792_,
		_w793_,
		_w794_
	);
	LUT2 #(
		.INIT('h2)
	) name616 (
		\254(101)_pad ,
		\257(102)_pad ,
		_w795_
	);
	LUT2 #(
		.INIT('h8)
	) name617 (
		\242(97)_pad ,
		\257(102)_pad ,
		_w796_
	);
	LUT2 #(
		.INIT('h1)
	) name618 (
		\389(136)_pad ,
		_w795_,
		_w797_
	);
	LUT2 #(
		.INIT('h4)
	) name619 (
		_w796_,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('h1)
	) name620 (
		_w794_,
		_w798_,
		_w799_
	);
	LUT2 #(
		.INIT('h1)
	) name621 (
		\251(100)_pad ,
		\281(108)_pad ,
		_w800_
	);
	LUT2 #(
		.INIT('h4)
	) name622 (
		\248(99)_pad ,
		\281(108)_pad ,
		_w801_
	);
	LUT2 #(
		.INIT('h2)
	) name623 (
		\374(134)_pad ,
		_w800_,
		_w802_
	);
	LUT2 #(
		.INIT('h4)
	) name624 (
		_w801_,
		_w802_,
		_w803_
	);
	LUT2 #(
		.INIT('h2)
	) name625 (
		\254(101)_pad ,
		\281(108)_pad ,
		_w804_
	);
	LUT2 #(
		.INIT('h8)
	) name626 (
		\242(97)_pad ,
		\281(108)_pad ,
		_w805_
	);
	LUT2 #(
		.INIT('h1)
	) name627 (
		\374(134)_pad ,
		_w804_,
		_w806_
	);
	LUT2 #(
		.INIT('h4)
	) name628 (
		_w805_,
		_w806_,
		_w807_
	);
	LUT2 #(
		.INIT('h1)
	) name629 (
		_w803_,
		_w807_,
		_w808_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		\251(100)_pad ,
		\273(106)_pad ,
		_w809_
	);
	LUT2 #(
		.INIT('h4)
	) name631 (
		\248(99)_pad ,
		\273(106)_pad ,
		_w810_
	);
	LUT2 #(
		.INIT('h2)
	) name632 (
		\411(138)_pad ,
		_w809_,
		_w811_
	);
	LUT2 #(
		.INIT('h4)
	) name633 (
		_w810_,
		_w811_,
		_w812_
	);
	LUT2 #(
		.INIT('h2)
	) name634 (
		\254(101)_pad ,
		\273(106)_pad ,
		_w813_
	);
	LUT2 #(
		.INIT('h8)
	) name635 (
		\242(97)_pad ,
		\273(106)_pad ,
		_w814_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		\411(138)_pad ,
		_w813_,
		_w815_
	);
	LUT2 #(
		.INIT('h4)
	) name637 (
		_w814_,
		_w815_,
		_w816_
	);
	LUT2 #(
		.INIT('h1)
	) name638 (
		_w812_,
		_w816_,
		_w817_
	);
	LUT2 #(
		.INIT('h4)
	) name639 (
		_w808_,
		_w817_,
		_w818_
	);
	LUT2 #(
		.INIT('h2)
	) name640 (
		_w808_,
		_w817_,
		_w819_
	);
	LUT2 #(
		.INIT('h1)
	) name641 (
		_w818_,
		_w819_,
		_w820_
	);
	LUT2 #(
		.INIT('h1)
	) name642 (
		\251(100)_pad ,
		\265(104)_pad ,
		_w821_
	);
	LUT2 #(
		.INIT('h4)
	) name643 (
		\248(99)_pad ,
		\265(104)_pad ,
		_w822_
	);
	LUT2 #(
		.INIT('h2)
	) name644 (
		\400(137)_pad ,
		_w821_,
		_w823_
	);
	LUT2 #(
		.INIT('h4)
	) name645 (
		_w822_,
		_w823_,
		_w824_
	);
	LUT2 #(
		.INIT('h2)
	) name646 (
		\254(101)_pad ,
		\265(104)_pad ,
		_w825_
	);
	LUT2 #(
		.INIT('h8)
	) name647 (
		\242(97)_pad ,
		\265(104)_pad ,
		_w826_
	);
	LUT2 #(
		.INIT('h1)
	) name648 (
		\400(137)_pad ,
		_w825_,
		_w827_
	);
	LUT2 #(
		.INIT('h4)
	) name649 (
		_w826_,
		_w827_,
		_w828_
	);
	LUT2 #(
		.INIT('h1)
	) name650 (
		_w824_,
		_w828_,
		_w829_
	);
	LUT2 #(
		.INIT('h2)
	) name651 (
		_w820_,
		_w829_,
		_w830_
	);
	LUT2 #(
		.INIT('h4)
	) name652 (
		_w820_,
		_w829_,
		_w831_
	);
	LUT2 #(
		.INIT('h1)
	) name653 (
		_w830_,
		_w831_,
		_w832_
	);
	LUT2 #(
		.INIT('h8)
	) name654 (
		_w799_,
		_w832_,
		_w833_
	);
	LUT2 #(
		.INIT('h1)
	) name655 (
		_w799_,
		_w832_,
		_w834_
	);
	LUT2 #(
		.INIT('h1)
	) name656 (
		_w833_,
		_w834_,
		_w835_
	);
	LUT2 #(
		.INIT('h2)
	) name657 (
		_w790_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h4)
	) name658 (
		_w790_,
		_w835_,
		_w837_
	);
	LUT2 #(
		.INIT('h1)
	) name659 (
		\4091(175)_pad ,
		_w836_,
		_w838_
	);
	LUT2 #(
		.INIT('h4)
	) name660 (
		_w837_,
		_w838_,
		_w839_
	);
	LUT2 #(
		.INIT('h1)
	) name661 (
		\4092(176)_pad ,
		_w839_,
		_w840_
	);
	LUT2 #(
		.INIT('h4)
	) name662 (
		_w742_,
		_w840_,
		_w841_
	);
	LUT2 #(
		.INIT('h1)
	) name663 (
		_w676_,
		_w841_,
		_w842_
	);
	LUT2 #(
		.INIT('h2)
	) name664 (
		_w479_,
		_w842_,
		_w843_
	);
	LUT2 #(
		.INIT('h8)
	) name665 (
		\4092(176)_pad ,
		\94(36)_pad ,
		_w844_
	);
	LUT2 #(
		.INIT('h1)
	) name666 (
		_w397_,
		_w403_,
		_w845_
	);
	LUT2 #(
		.INIT('h1)
	) name667 (
		_w404_,
		_w845_,
		_w846_
	);
	LUT2 #(
		.INIT('h2)
	) name668 (
		_w391_,
		_w415_,
		_w847_
	);
	LUT2 #(
		.INIT('h4)
	) name669 (
		_w391_,
		_w415_,
		_w848_
	);
	LUT2 #(
		.INIT('h1)
	) name670 (
		_w847_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h8)
	) name671 (
		_w846_,
		_w849_,
		_w850_
	);
	LUT2 #(
		.INIT('h1)
	) name672 (
		_w846_,
		_w849_,
		_w851_
	);
	LUT2 #(
		.INIT('h1)
	) name673 (
		_w850_,
		_w851_,
		_w852_
	);
	LUT2 #(
		.INIT('h4)
	) name674 (
		_w395_,
		_w402_,
		_w853_
	);
	LUT2 #(
		.INIT('h1)
	) name675 (
		_w396_,
		_w402_,
		_w854_
	);
	LUT2 #(
		.INIT('h1)
	) name676 (
		_w853_,
		_w854_,
		_w855_
	);
	LUT2 #(
		.INIT('h1)
	) name677 (
		_w409_,
		_w855_,
		_w856_
	);
	LUT2 #(
		.INIT('h1)
	) name678 (
		_w446_,
		_w856_,
		_w857_
	);
	LUT2 #(
		.INIT('h2)
	) name679 (
		_w446_,
		_w855_,
		_w858_
	);
	LUT2 #(
		.INIT('h1)
	) name680 (
		_w857_,
		_w858_,
		_w859_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		_w407_,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('h8)
	) name682 (
		_w407_,
		_w859_,
		_w861_
	);
	LUT2 #(
		.INIT('h1)
	) name683 (
		_w860_,
		_w861_,
		_w862_
	);
	LUT2 #(
		.INIT('h2)
	) name684 (
		\2174(161)_pad ,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h4)
	) name685 (
		_w389_,
		_w444_,
		_w864_
	);
	LUT2 #(
		.INIT('h1)
	) name686 (
		_w445_,
		_w864_,
		_w865_
	);
	LUT2 #(
		.INIT('h1)
	) name687 (
		_w401_,
		_w865_,
		_w866_
	);
	LUT2 #(
		.INIT('h8)
	) name688 (
		_w401_,
		_w865_,
		_w867_
	);
	LUT2 #(
		.INIT('h2)
	) name689 (
		_w407_,
		_w866_,
		_w868_
	);
	LUT2 #(
		.INIT('h4)
	) name690 (
		_w867_,
		_w868_,
		_w869_
	);
	LUT2 #(
		.INIT('h1)
	) name691 (
		\2174(161)_pad ,
		_w860_,
		_w870_
	);
	LUT2 #(
		.INIT('h4)
	) name692 (
		_w869_,
		_w870_,
		_w871_
	);
	LUT2 #(
		.INIT('h1)
	) name693 (
		_w863_,
		_w871_,
		_w872_
	);
	LUT2 #(
		.INIT('h8)
	) name694 (
		\2174(161)_pad ,
		_w416_,
		_w873_
	);
	LUT2 #(
		.INIT('h1)
	) name695 (
		_w448_,
		_w873_,
		_w874_
	);
	LUT2 #(
		.INIT('h1)
	) name696 (
		_w422_,
		_w440_,
		_w875_
	);
	LUT2 #(
		.INIT('h2)
	) name697 (
		_w419_,
		_w875_,
		_w876_
	);
	LUT2 #(
		.INIT('h4)
	) name698 (
		_w419_,
		_w875_,
		_w877_
	);
	LUT2 #(
		.INIT('h1)
	) name699 (
		_w876_,
		_w877_,
		_w878_
	);
	LUT2 #(
		.INIT('h2)
	) name700 (
		_w588_,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('h4)
	) name701 (
		_w588_,
		_w878_,
		_w880_
	);
	LUT2 #(
		.INIT('h1)
	) name702 (
		_w879_,
		_w880_,
		_w881_
	);
	LUT2 #(
		.INIT('h2)
	) name703 (
		_w874_,
		_w881_,
		_w882_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		_w429_,
		_w433_,
		_w883_
	);
	LUT2 #(
		.INIT('h1)
	) name705 (
		_w439_,
		_w883_,
		_w884_
	);
	LUT2 #(
		.INIT('h1)
	) name706 (
		_w427_,
		_w586_,
		_w885_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w422_,
		_w885_,
		_w886_
	);
	LUT2 #(
		.INIT('h2)
	) name708 (
		_w419_,
		_w886_,
		_w887_
	);
	LUT2 #(
		.INIT('h4)
	) name709 (
		_w419_,
		_w886_,
		_w888_
	);
	LUT2 #(
		.INIT('h1)
	) name710 (
		_w887_,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h8)
	) name711 (
		_w884_,
		_w889_,
		_w890_
	);
	LUT2 #(
		.INIT('h1)
	) name712 (
		_w884_,
		_w889_,
		_w891_
	);
	LUT2 #(
		.INIT('h1)
	) name713 (
		_w890_,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h1)
	) name714 (
		_w874_,
		_w892_,
		_w893_
	);
	LUT2 #(
		.INIT('h1)
	) name715 (
		_w882_,
		_w893_,
		_w894_
	);
	LUT2 #(
		.INIT('h2)
	) name716 (
		_w872_,
		_w894_,
		_w895_
	);
	LUT2 #(
		.INIT('h4)
	) name717 (
		_w872_,
		_w894_,
		_w896_
	);
	LUT2 #(
		.INIT('h1)
	) name718 (
		_w895_,
		_w896_,
		_w897_
	);
	LUT2 #(
		.INIT('h8)
	) name719 (
		_w852_,
		_w897_,
		_w898_
	);
	LUT2 #(
		.INIT('h1)
	) name720 (
		_w852_,
		_w897_,
		_w899_
	);
	LUT2 #(
		.INIT('h1)
	) name721 (
		_w898_,
		_w899_,
		_w900_
	);
	LUT2 #(
		.INIT('h8)
	) name722 (
		\4091(175)_pad ,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h4)
	) name723 (
		\248(99)_pad ,
		\514(147)_pad ,
		_w902_
	);
	LUT2 #(
		.INIT('h2)
	) name724 (
		\242(97)_pad ,
		\514(147)_pad ,
		_w903_
	);
	LUT2 #(
		.INIT('h1)
	) name725 (
		_w902_,
		_w903_,
		_w904_
	);
	LUT2 #(
		.INIT('h4)
	) name726 (
		_w373_,
		_w376_,
		_w905_
	);
	LUT2 #(
		.INIT('h1)
	) name727 (
		_w377_,
		_w905_,
		_w906_
	);
	LUT2 #(
		.INIT('h8)
	) name728 (
		_w330_,
		_w339_,
		_w907_
	);
	LUT2 #(
		.INIT('h1)
	) name729 (
		_w340_,
		_w907_,
		_w908_
	);
	LUT2 #(
		.INIT('h2)
	) name730 (
		_w906_,
		_w908_,
		_w909_
	);
	LUT2 #(
		.INIT('h4)
	) name731 (
		_w906_,
		_w908_,
		_w910_
	);
	LUT2 #(
		.INIT('h1)
	) name732 (
		_w909_,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h8)
	) name733 (
		_w904_,
		_w911_,
		_w912_
	);
	LUT2 #(
		.INIT('h1)
	) name734 (
		_w904_,
		_w911_,
		_w913_
	);
	LUT2 #(
		.INIT('h1)
	) name735 (
		_w912_,
		_w913_,
		_w914_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		\251(100)_pad ,
		\324(120)_pad ,
		_w915_
	);
	LUT2 #(
		.INIT('h4)
	) name737 (
		\248(99)_pad ,
		\324(120)_pad ,
		_w916_
	);
	LUT2 #(
		.INIT('h2)
	) name738 (
		\503(146)_pad ,
		_w915_,
		_w917_
	);
	LUT2 #(
		.INIT('h4)
	) name739 (
		_w916_,
		_w917_,
		_w918_
	);
	LUT2 #(
		.INIT('h2)
	) name740 (
		\254(101)_pad ,
		\324(120)_pad ,
		_w919_
	);
	LUT2 #(
		.INIT('h8)
	) name741 (
		\242(97)_pad ,
		\324(120)_pad ,
		_w920_
	);
	LUT2 #(
		.INIT('h1)
	) name742 (
		\503(146)_pad ,
		_w919_,
		_w921_
	);
	LUT2 #(
		.INIT('h4)
	) name743 (
		_w920_,
		_w921_,
		_w922_
	);
	LUT2 #(
		.INIT('h1)
	) name744 (
		_w918_,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('h2)
	) name745 (
		_w343_,
		_w923_,
		_w924_
	);
	LUT2 #(
		.INIT('h4)
	) name746 (
		_w343_,
		_w923_,
		_w925_
	);
	LUT2 #(
		.INIT('h1)
	) name747 (
		_w924_,
		_w925_,
		_w926_
	);
	LUT2 #(
		.INIT('h1)
	) name748 (
		\251(100)_pad ,
		\341(125)_pad ,
		_w927_
	);
	LUT2 #(
		.INIT('h4)
	) name749 (
		\248(99)_pad ,
		\341(125)_pad ,
		_w928_
	);
	LUT2 #(
		.INIT('h2)
	) name750 (
		\523(148)_pad ,
		_w927_,
		_w929_
	);
	LUT2 #(
		.INIT('h4)
	) name751 (
		_w928_,
		_w929_,
		_w930_
	);
	LUT2 #(
		.INIT('h2)
	) name752 (
		\254(101)_pad ,
		\341(125)_pad ,
		_w931_
	);
	LUT2 #(
		.INIT('h8)
	) name753 (
		\242(97)_pad ,
		\341(125)_pad ,
		_w932_
	);
	LUT2 #(
		.INIT('h1)
	) name754 (
		\523(148)_pad ,
		_w931_,
		_w933_
	);
	LUT2 #(
		.INIT('h4)
	) name755 (
		_w932_,
		_w933_,
		_w934_
	);
	LUT2 #(
		.INIT('h1)
	) name756 (
		_w930_,
		_w934_,
		_w935_
	);
	LUT2 #(
		.INIT('h1)
	) name757 (
		\251(100)_pad ,
		\351(127)_pad ,
		_w936_
	);
	LUT2 #(
		.INIT('h4)
	) name758 (
		\248(99)_pad ,
		\351(127)_pad ,
		_w937_
	);
	LUT2 #(
		.INIT('h2)
	) name759 (
		\534(149)_pad ,
		_w936_,
		_w938_
	);
	LUT2 #(
		.INIT('h4)
	) name760 (
		_w937_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h2)
	) name761 (
		\254(101)_pad ,
		\351(127)_pad ,
		_w940_
	);
	LUT2 #(
		.INIT('h8)
	) name762 (
		\242(97)_pad ,
		\351(127)_pad ,
		_w941_
	);
	LUT2 #(
		.INIT('h1)
	) name763 (
		\534(149)_pad ,
		_w940_,
		_w942_
	);
	LUT2 #(
		.INIT('h4)
	) name764 (
		_w941_,
		_w942_,
		_w943_
	);
	LUT2 #(
		.INIT('h1)
	) name765 (
		_w939_,
		_w943_,
		_w944_
	);
	LUT2 #(
		.INIT('h2)
	) name766 (
		_w935_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h4)
	) name767 (
		_w935_,
		_w944_,
		_w946_
	);
	LUT2 #(
		.INIT('h1)
	) name768 (
		_w945_,
		_w946_,
		_w947_
	);
	LUT2 #(
		.INIT('h8)
	) name769 (
		_w926_,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h1)
	) name770 (
		_w926_,
		_w947_,
		_w949_
	);
	LUT2 #(
		.INIT('h1)
	) name771 (
		_w948_,
		_w949_,
		_w950_
	);
	LUT2 #(
		.INIT('h1)
	) name772 (
		_w914_,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h8)
	) name773 (
		_w914_,
		_w950_,
		_w952_
	);
	LUT2 #(
		.INIT('h1)
	) name774 (
		\4091(175)_pad ,
		_w951_,
		_w953_
	);
	LUT2 #(
		.INIT('h4)
	) name775 (
		_w952_,
		_w953_,
		_w954_
	);
	LUT2 #(
		.INIT('h1)
	) name776 (
		\4092(176)_pad ,
		_w954_,
		_w955_
	);
	LUT2 #(
		.INIT('h4)
	) name777 (
		_w901_,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h1)
	) name778 (
		_w844_,
		_w956_,
		_w957_
	);
	LUT2 #(
		.INIT('h2)
	) name779 (
		_w508_,
		_w957_,
		_w958_
	);
	LUT2 #(
		.INIT('h8)
	) name780 (
		\179(78)_pad ,
		_w504_,
		_w959_
	);
	LUT2 #(
		.INIT('h8)
	) name781 (
		\176(77)_pad ,
		_w506_,
		_w960_
	);
	LUT2 #(
		.INIT('h1)
	) name782 (
		_w959_,
		_w960_,
		_w961_
	);
	LUT2 #(
		.INIT('h4)
	) name783 (
		_w958_,
		_w961_,
		_w962_
	);
	LUT2 #(
		.INIT('h4)
	) name784 (
		_w843_,
		_w962_,
		_w963_
	);
	LUT2 #(
		.INIT('h2)
	) name785 (
		\926(624)_pad ,
		_w963_,
		_w964_
	);
	LUT2 #(
		.INIT('h8)
	) name786 (
		_w343_,
		_w480_,
		_w965_
	);
	LUT2 #(
		.INIT('h2)
	) name787 (
		\54(20)_pad ,
		_w407_,
		_w966_
	);
	LUT2 #(
		.INIT('h4)
	) name788 (
		\54(20)_pad ,
		_w407_,
		_w967_
	);
	LUT2 #(
		.INIT('h1)
	) name789 (
		_w966_,
		_w967_,
		_w968_
	);
	LUT2 #(
		.INIT('h2)
	) name790 (
		_w491_,
		_w968_,
		_w969_
	);
	LUT2 #(
		.INIT('h8)
	) name791 (
		\131(59)_pad ,
		_w499_,
		_w970_
	);
	LUT2 #(
		.INIT('h1)
	) name792 (
		_w965_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h4)
	) name793 (
		_w969_,
		_w971_,
		_w972_
	);
	LUT2 #(
		.INIT('h2)
	) name794 (
		_w508_,
		_w972_,
		_w973_
	);
	LUT2 #(
		.INIT('h8)
	) name795 (
		\185(80)_pad ,
		_w504_,
		_w974_
	);
	LUT2 #(
		.INIT('h8)
	) name796 (
		\182(79)_pad ,
		_w506_,
		_w975_
	);
	LUT2 #(
		.INIT('h4)
	) name797 (
		\281(108)_pad ,
		\3550(167)_pad ,
		_w976_
	);
	LUT2 #(
		.INIT('h8)
	) name798 (
		\281(108)_pad ,
		\3552(168)_pad ,
		_w977_
	);
	LUT2 #(
		.INIT('h2)
	) name799 (
		\374(134)_pad ,
		_w976_,
		_w978_
	);
	LUT2 #(
		.INIT('h4)
	) name800 (
		_w977_,
		_w978_,
		_w979_
	);
	LUT2 #(
		.INIT('h1)
	) name801 (
		\281(108)_pad ,
		\3548(166)_pad ,
		_w980_
	);
	LUT2 #(
		.INIT('h2)
	) name802 (
		\281(108)_pad ,
		\3546(165)_pad ,
		_w981_
	);
	LUT2 #(
		.INIT('h1)
	) name803 (
		\374(134)_pad ,
		_w980_,
		_w982_
	);
	LUT2 #(
		.INIT('h4)
	) name804 (
		_w981_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h1)
	) name805 (
		_w979_,
		_w983_,
		_w984_
	);
	LUT2 #(
		.INIT('h8)
	) name806 (
		_w480_,
		_w984_,
		_w985_
	);
	LUT2 #(
		.INIT('h8)
	) name807 (
		\4(1)_pad ,
		_w296_,
		_w986_
	);
	LUT2 #(
		.INIT('h1)
	) name808 (
		\4(1)_pad ,
		_w296_,
		_w987_
	);
	LUT2 #(
		.INIT('h1)
	) name809 (
		_w986_,
		_w987_,
		_w988_
	);
	LUT2 #(
		.INIT('h8)
	) name810 (
		_w491_,
		_w988_,
		_w989_
	);
	LUT2 #(
		.INIT('h8)
	) name811 (
		\117(47)_pad ,
		_w499_,
		_w990_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		_w985_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h4)
	) name813 (
		_w989_,
		_w991_,
		_w992_
	);
	LUT2 #(
		.INIT('h2)
	) name814 (
		_w479_,
		_w992_,
		_w993_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w974_,
		_w975_,
		_w994_
	);
	LUT2 #(
		.INIT('h4)
	) name816 (
		_w973_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h4)
	) name817 (
		_w993_,
		_w995_,
		_w996_
	);
	LUT2 #(
		.INIT('h2)
	) name818 (
		\926(624)_pad ,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h8)
	) name819 (
		_w370_,
		_w480_,
		_w998_
	);
	LUT2 #(
		.INIT('h8)
	) name820 (
		\129(57)_pad ,
		_w499_,
		_w999_
	);
	LUT2 #(
		.INIT('h4)
	) name821 (
		_w403_,
		_w967_,
		_w1000_
	);
	LUT2 #(
		.INIT('h1)
	) name822 (
		_w402_,
		_w967_,
		_w1001_
	);
	LUT2 #(
		.INIT('h4)
	) name823 (
		_w401_,
		_w1001_,
		_w1002_
	);
	LUT2 #(
		.INIT('h2)
	) name824 (
		_w491_,
		_w1000_,
		_w1003_
	);
	LUT2 #(
		.INIT('h4)
	) name825 (
		_w1002_,
		_w1003_,
		_w1004_
	);
	LUT2 #(
		.INIT('h1)
	) name826 (
		_w998_,
		_w999_,
		_w1005_
	);
	LUT2 #(
		.INIT('h4)
	) name827 (
		_w1004_,
		_w1005_,
		_w1006_
	);
	LUT2 #(
		.INIT('h2)
	) name828 (
		_w508_,
		_w1006_,
		_w1007_
	);
	LUT2 #(
		.INIT('h8)
	) name829 (
		\158(71)_pad ,
		_w504_,
		_w1008_
	);
	LUT2 #(
		.INIT('h8)
	) name830 (
		\188(81)_pad ,
		_w506_,
		_w1009_
	);
	LUT2 #(
		.INIT('h4)
	) name831 (
		\273(106)_pad ,
		\3550(167)_pad ,
		_w1010_
	);
	LUT2 #(
		.INIT('h8)
	) name832 (
		\273(106)_pad ,
		\3552(168)_pad ,
		_w1011_
	);
	LUT2 #(
		.INIT('h2)
	) name833 (
		\411(138)_pad ,
		_w1010_,
		_w1012_
	);
	LUT2 #(
		.INIT('h4)
	) name834 (
		_w1011_,
		_w1012_,
		_w1013_
	);
	LUT2 #(
		.INIT('h1)
	) name835 (
		\273(106)_pad ,
		\3548(166)_pad ,
		_w1014_
	);
	LUT2 #(
		.INIT('h2)
	) name836 (
		\273(106)_pad ,
		\3546(165)_pad ,
		_w1015_
	);
	LUT2 #(
		.INIT('h1)
	) name837 (
		\411(138)_pad ,
		_w1014_,
		_w1016_
	);
	LUT2 #(
		.INIT('h4)
	) name838 (
		_w1015_,
		_w1016_,
		_w1017_
	);
	LUT2 #(
		.INIT('h1)
	) name839 (
		_w1013_,
		_w1017_,
		_w1018_
	);
	LUT2 #(
		.INIT('h8)
	) name840 (
		_w480_,
		_w1018_,
		_w1019_
	);
	LUT2 #(
		.INIT('h2)
	) name841 (
		\4(1)_pad ,
		_w295_,
		_w1020_
	);
	LUT2 #(
		.INIT('h1)
	) name842 (
		_w294_,
		_w1020_,
		_w1021_
	);
	LUT2 #(
		.INIT('h2)
	) name843 (
		_w299_,
		_w1021_,
		_w1022_
	);
	LUT2 #(
		.INIT('h4)
	) name844 (
		_w299_,
		_w1021_,
		_w1023_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		_w1022_,
		_w1023_,
		_w1024_
	);
	LUT2 #(
		.INIT('h8)
	) name846 (
		_w491_,
		_w1024_,
		_w1025_
	);
	LUT2 #(
		.INIT('h8)
	) name847 (
		\126(54)_pad ,
		_w499_,
		_w1026_
	);
	LUT2 #(
		.INIT('h1)
	) name848 (
		_w1019_,
		_w1026_,
		_w1027_
	);
	LUT2 #(
		.INIT('h4)
	) name849 (
		_w1025_,
		_w1027_,
		_w1028_
	);
	LUT2 #(
		.INIT('h2)
	) name850 (
		_w479_,
		_w1028_,
		_w1029_
	);
	LUT2 #(
		.INIT('h1)
	) name851 (
		_w1008_,
		_w1009_,
		_w1030_
	);
	LUT2 #(
		.INIT('h4)
	) name852 (
		_w1007_,
		_w1030_,
		_w1031_
	);
	LUT2 #(
		.INIT('h4)
	) name853 (
		_w1029_,
		_w1031_,
		_w1032_
	);
	LUT2 #(
		.INIT('h2)
	) name854 (
		\926(624)_pad ,
		_w1032_,
		_w1033_
	);
	LUT2 #(
		.INIT('h8)
	) name855 (
		_w352_,
		_w480_,
		_w1034_
	);
	LUT2 #(
		.INIT('h1)
	) name856 (
		_w401_,
		_w1001_,
		_w1035_
	);
	LUT2 #(
		.INIT('h8)
	) name857 (
		_w397_,
		_w1035_,
		_w1036_
	);
	LUT2 #(
		.INIT('h1)
	) name858 (
		_w397_,
		_w1035_,
		_w1037_
	);
	LUT2 #(
		.INIT('h1)
	) name859 (
		_w1036_,
		_w1037_,
		_w1038_
	);
	LUT2 #(
		.INIT('h2)
	) name860 (
		_w491_,
		_w1038_,
		_w1039_
	);
	LUT2 #(
		.INIT('h8)
	) name861 (
		\119(49)_pad ,
		_w499_,
		_w1040_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		_w1034_,
		_w1040_,
		_w1041_
	);
	LUT2 #(
		.INIT('h4)
	) name863 (
		_w1039_,
		_w1041_,
		_w1042_
	);
	LUT2 #(
		.INIT('h2)
	) name864 (
		_w508_,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('h8)
	) name865 (
		\152(69)_pad ,
		_w504_,
		_w1044_
	);
	LUT2 #(
		.INIT('h8)
	) name866 (
		\155(70)_pad ,
		_w506_,
		_w1045_
	);
	LUT2 #(
		.INIT('h4)
	) name867 (
		\265(104)_pad ,
		\3550(167)_pad ,
		_w1046_
	);
	LUT2 #(
		.INIT('h8)
	) name868 (
		\265(104)_pad ,
		\3552(168)_pad ,
		_w1047_
	);
	LUT2 #(
		.INIT('h2)
	) name869 (
		\400(137)_pad ,
		_w1046_,
		_w1048_
	);
	LUT2 #(
		.INIT('h4)
	) name870 (
		_w1047_,
		_w1048_,
		_w1049_
	);
	LUT2 #(
		.INIT('h1)
	) name871 (
		\265(104)_pad ,
		\3548(166)_pad ,
		_w1050_
	);
	LUT2 #(
		.INIT('h2)
	) name872 (
		\265(104)_pad ,
		\3546(165)_pad ,
		_w1051_
	);
	LUT2 #(
		.INIT('h1)
	) name873 (
		\400(137)_pad ,
		_w1050_,
		_w1052_
	);
	LUT2 #(
		.INIT('h4)
	) name874 (
		_w1051_,
		_w1052_,
		_w1053_
	);
	LUT2 #(
		.INIT('h1)
	) name875 (
		_w1049_,
		_w1053_,
		_w1054_
	);
	LUT2 #(
		.INIT('h8)
	) name876 (
		_w480_,
		_w1054_,
		_w1055_
	);
	LUT2 #(
		.INIT('h1)
	) name877 (
		_w298_,
		_w1021_,
		_w1056_
	);
	LUT2 #(
		.INIT('h1)
	) name878 (
		_w297_,
		_w1056_,
		_w1057_
	);
	LUT2 #(
		.INIT('h2)
	) name879 (
		_w302_,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h4)
	) name880 (
		_w302_,
		_w1057_,
		_w1059_
	);
	LUT2 #(
		.INIT('h1)
	) name881 (
		_w1058_,
		_w1059_,
		_w1060_
	);
	LUT2 #(
		.INIT('h8)
	) name882 (
		_w491_,
		_w1060_,
		_w1061_
	);
	LUT2 #(
		.INIT('h8)
	) name883 (
		\127(55)_pad ,
		_w499_,
		_w1062_
	);
	LUT2 #(
		.INIT('h1)
	) name884 (
		_w1055_,
		_w1062_,
		_w1063_
	);
	LUT2 #(
		.INIT('h4)
	) name885 (
		_w1061_,
		_w1063_,
		_w1064_
	);
	LUT2 #(
		.INIT('h2)
	) name886 (
		_w479_,
		_w1064_,
		_w1065_
	);
	LUT2 #(
		.INIT('h1)
	) name887 (
		_w1044_,
		_w1045_,
		_w1066_
	);
	LUT2 #(
		.INIT('h4)
	) name888 (
		_w1043_,
		_w1066_,
		_w1067_
	);
	LUT2 #(
		.INIT('h4)
	) name889 (
		_w1065_,
		_w1067_,
		_w1068_
	);
	LUT2 #(
		.INIT('h2)
	) name890 (
		\926(624)_pad ,
		_w1068_,
		_w1069_
	);
	LUT2 #(
		.INIT('h8)
	) name891 (
		_w380_,
		_w480_,
		_w1070_
	);
	LUT2 #(
		.INIT('h1)
	) name892 (
		_w444_,
		_w510_,
		_w1071_
	);
	LUT2 #(
		.INIT('h8)
	) name893 (
		_w391_,
		_w1071_,
		_w1072_
	);
	LUT2 #(
		.INIT('h1)
	) name894 (
		_w391_,
		_w1071_,
		_w1073_
	);
	LUT2 #(
		.INIT('h1)
	) name895 (
		_w1072_,
		_w1073_,
		_w1074_
	);
	LUT2 #(
		.INIT('h2)
	) name896 (
		_w491_,
		_w1074_,
		_w1075_
	);
	LUT2 #(
		.INIT('h8)
	) name897 (
		\130(58)_pad ,
		_w499_,
		_w1076_
	);
	LUT2 #(
		.INIT('h1)
	) name898 (
		_w1070_,
		_w1076_,
		_w1077_
	);
	LUT2 #(
		.INIT('h4)
	) name899 (
		_w1075_,
		_w1077_,
		_w1078_
	);
	LUT2 #(
		.INIT('h2)
	) name900 (
		_w508_,
		_w1078_,
		_w1079_
	);
	LUT2 #(
		.INIT('h8)
	) name901 (
		\146(67)_pad ,
		_w504_,
		_w1080_
	);
	LUT2 #(
		.INIT('h8)
	) name902 (
		\149(68)_pad ,
		_w506_,
		_w1081_
	);
	LUT2 #(
		.INIT('h4)
	) name903 (
		\257(102)_pad ,
		\3550(167)_pad ,
		_w1082_
	);
	LUT2 #(
		.INIT('h8)
	) name904 (
		\257(102)_pad ,
		\3552(168)_pad ,
		_w1083_
	);
	LUT2 #(
		.INIT('h2)
	) name905 (
		\389(136)_pad ,
		_w1082_,
		_w1084_
	);
	LUT2 #(
		.INIT('h4)
	) name906 (
		_w1083_,
		_w1084_,
		_w1085_
	);
	LUT2 #(
		.INIT('h1)
	) name907 (
		\257(102)_pad ,
		\3548(166)_pad ,
		_w1086_
	);
	LUT2 #(
		.INIT('h2)
	) name908 (
		\257(102)_pad ,
		\3546(165)_pad ,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name909 (
		\389(136)_pad ,
		_w1086_,
		_w1088_
	);
	LUT2 #(
		.INIT('h4)
	) name910 (
		_w1087_,
		_w1088_,
		_w1089_
	);
	LUT2 #(
		.INIT('h1)
	) name911 (
		_w1085_,
		_w1089_,
		_w1090_
	);
	LUT2 #(
		.INIT('h8)
	) name912 (
		_w480_,
		_w1090_,
		_w1091_
	);
	LUT2 #(
		.INIT('h1)
	) name913 (
		_w458_,
		_w492_,
		_w1092_
	);
	LUT2 #(
		.INIT('h8)
	) name914 (
		_w310_,
		_w1092_,
		_w1093_
	);
	LUT2 #(
		.INIT('h1)
	) name915 (
		_w310_,
		_w1092_,
		_w1094_
	);
	LUT2 #(
		.INIT('h1)
	) name916 (
		_w1093_,
		_w1094_,
		_w1095_
	);
	LUT2 #(
		.INIT('h2)
	) name917 (
		_w491_,
		_w1095_,
		_w1096_
	);
	LUT2 #(
		.INIT('h8)
	) name918 (
		\128(56)_pad ,
		_w499_,
		_w1097_
	);
	LUT2 #(
		.INIT('h1)
	) name919 (
		_w1091_,
		_w1097_,
		_w1098_
	);
	LUT2 #(
		.INIT('h4)
	) name920 (
		_w1096_,
		_w1098_,
		_w1099_
	);
	LUT2 #(
		.INIT('h2)
	) name921 (
		_w479_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h1)
	) name922 (
		_w1080_,
		_w1081_,
		_w1101_
	);
	LUT2 #(
		.INIT('h4)
	) name923 (
		_w1079_,
		_w1101_,
		_w1102_
	);
	LUT2 #(
		.INIT('h4)
	) name924 (
		_w1100_,
		_w1102_,
		_w1103_
	);
	LUT2 #(
		.INIT('h2)
	) name925 (
		\926(624)_pad ,
		_w1103_,
		_w1104_
	);
	LUT2 #(
		.INIT('h4)
	) name926 (
		\2358(162)_pad ,
		\26(9)_pad ,
		_w1105_
	);
	LUT2 #(
		.INIT('h8)
	) name927 (
		\2358(162)_pad ,
		\81(29)_pad ,
		_w1106_
	);
	LUT2 #(
		.INIT('h2)
	) name928 (
		_w469_,
		_w1105_,
		_w1107_
	);
	LUT2 #(
		.INIT('h4)
	) name929 (
		_w1106_,
		_w1107_,
		_w1108_
	);
	LUT2 #(
		.INIT('h2)
	) name930 (
		\144(354)_pad ,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h2)
	) name931 (
		\1691(159)_pad ,
		\1694(160)_pad ,
		_w1110_
	);
	LUT2 #(
		.INIT('h4)
	) name932 (
		_w502_,
		_w1110_,
		_w1111_
	);
	LUT2 #(
		.INIT('h8)
	) name933 (
		\1691(159)_pad ,
		\1694(160)_pad ,
		_w1112_
	);
	LUT2 #(
		.INIT('h8)
	) name934 (
		\170(75)_pad ,
		_w1112_,
		_w1113_
	);
	LUT2 #(
		.INIT('h4)
	) name935 (
		\1691(159)_pad ,
		\1694(160)_pad ,
		_w1114_
	);
	LUT2 #(
		.INIT('h8)
	) name936 (
		\200(85)_pad ,
		_w1114_,
		_w1115_
	);
	LUT2 #(
		.INIT('h1)
	) name937 (
		\1691(159)_pad ,
		\1694(160)_pad ,
		_w1116_
	);
	LUT2 #(
		.INIT('h4)
	) name938 (
		_w519_,
		_w1116_,
		_w1117_
	);
	LUT2 #(
		.INIT('h1)
	) name939 (
		_w1113_,
		_w1115_,
		_w1118_
	);
	LUT2 #(
		.INIT('h4)
	) name940 (
		_w1111_,
		_w1118_,
		_w1119_
	);
	LUT2 #(
		.INIT('h4)
	) name941 (
		_w1117_,
		_w1119_,
		_w1120_
	);
	LUT2 #(
		.INIT('h2)
	) name942 (
		\926(624)_pad ,
		_w1120_,
		_w1121_
	);
	LUT2 #(
		.INIT('h4)
	) name943 (
		_w544_,
		_w1110_,
		_w1122_
	);
	LUT2 #(
		.INIT('h8)
	) name944 (
		\173(76)_pad ,
		_w1112_,
		_w1123_
	);
	LUT2 #(
		.INIT('h8)
	) name945 (
		\203(86)_pad ,
		_w1114_,
		_w1124_
	);
	LUT2 #(
		.INIT('h4)
	) name946 (
		_w556_,
		_w1116_,
		_w1125_
	);
	LUT2 #(
		.INIT('h1)
	) name947 (
		_w1123_,
		_w1124_,
		_w1126_
	);
	LUT2 #(
		.INIT('h4)
	) name948 (
		_w1122_,
		_w1126_,
		_w1127_
	);
	LUT2 #(
		.INIT('h4)
	) name949 (
		_w1125_,
		_w1127_,
		_w1128_
	);
	LUT2 #(
		.INIT('h2)
	) name950 (
		\926(624)_pad ,
		_w1128_,
		_w1129_
	);
	LUT2 #(
		.INIT('h4)
	) name951 (
		_w580_,
		_w1110_,
		_w1130_
	);
	LUT2 #(
		.INIT('h8)
	) name952 (
		\167(74)_pad ,
		_w1112_,
		_w1131_
	);
	LUT2 #(
		.INIT('h8)
	) name953 (
		\197(84)_pad ,
		_w1114_,
		_w1132_
	);
	LUT2 #(
		.INIT('h4)
	) name954 (
		_w594_,
		_w1116_,
		_w1133_
	);
	LUT2 #(
		.INIT('h1)
	) name955 (
		_w1131_,
		_w1132_,
		_w1134_
	);
	LUT2 #(
		.INIT('h4)
	) name956 (
		_w1130_,
		_w1134_,
		_w1135_
	);
	LUT2 #(
		.INIT('h4)
	) name957 (
		_w1133_,
		_w1135_,
		_w1136_
	);
	LUT2 #(
		.INIT('h2)
	) name958 (
		\926(624)_pad ,
		_w1136_,
		_w1137_
	);
	LUT2 #(
		.INIT('h4)
	) name959 (
		_w619_,
		_w1110_,
		_w1138_
	);
	LUT2 #(
		.INIT('h8)
	) name960 (
		\164(73)_pad ,
		_w1112_,
		_w1139_
	);
	LUT2 #(
		.INIT('h8)
	) name961 (
		\194(83)_pad ,
		_w1114_,
		_w1140_
	);
	LUT2 #(
		.INIT('h4)
	) name962 (
		_w632_,
		_w1116_,
		_w1141_
	);
	LUT2 #(
		.INIT('h1)
	) name963 (
		_w1139_,
		_w1140_,
		_w1142_
	);
	LUT2 #(
		.INIT('h4)
	) name964 (
		_w1138_,
		_w1142_,
		_w1143_
	);
	LUT2 #(
		.INIT('h4)
	) name965 (
		_w1141_,
		_w1143_,
		_w1144_
	);
	LUT2 #(
		.INIT('h2)
	) name966 (
		\926(624)_pad ,
		_w1144_,
		_w1145_
	);
	LUT2 #(
		.INIT('h4)
	) name967 (
		_w658_,
		_w1110_,
		_w1146_
	);
	LUT2 #(
		.INIT('h8)
	) name968 (
		\161(72)_pad ,
		_w1112_,
		_w1147_
	);
	LUT2 #(
		.INIT('h8)
	) name969 (
		\191(82)_pad ,
		_w1114_,
		_w1148_
	);
	LUT2 #(
		.INIT('h4)
	) name970 (
		_w669_,
		_w1116_,
		_w1149_
	);
	LUT2 #(
		.INIT('h1)
	) name971 (
		_w1147_,
		_w1148_,
		_w1150_
	);
	LUT2 #(
		.INIT('h4)
	) name972 (
		_w1146_,
		_w1150_,
		_w1151_
	);
	LUT2 #(
		.INIT('h4)
	) name973 (
		_w1149_,
		_w1151_,
		_w1152_
	);
	LUT2 #(
		.INIT('h2)
	) name974 (
		\926(624)_pad ,
		_w1152_,
		_w1153_
	);
	LUT2 #(
		.INIT('h4)
	) name975 (
		_w842_,
		_w1110_,
		_w1154_
	);
	LUT2 #(
		.INIT('h4)
	) name976 (
		_w957_,
		_w1116_,
		_w1155_
	);
	LUT2 #(
		.INIT('h8)
	) name977 (
		\179(78)_pad ,
		_w1112_,
		_w1156_
	);
	LUT2 #(
		.INIT('h8)
	) name978 (
		\176(77)_pad ,
		_w1114_,
		_w1157_
	);
	LUT2 #(
		.INIT('h1)
	) name979 (
		_w1156_,
		_w1157_,
		_w1158_
	);
	LUT2 #(
		.INIT('h4)
	) name980 (
		_w1155_,
		_w1158_,
		_w1159_
	);
	LUT2 #(
		.INIT('h4)
	) name981 (
		_w1154_,
		_w1159_,
		_w1160_
	);
	LUT2 #(
		.INIT('h2)
	) name982 (
		\926(624)_pad ,
		_w1160_,
		_w1161_
	);
	LUT2 #(
		.INIT('h4)
	) name983 (
		_w972_,
		_w1116_,
		_w1162_
	);
	LUT2 #(
		.INIT('h8)
	) name984 (
		\185(80)_pad ,
		_w1112_,
		_w1163_
	);
	LUT2 #(
		.INIT('h8)
	) name985 (
		\182(79)_pad ,
		_w1114_,
		_w1164_
	);
	LUT2 #(
		.INIT('h4)
	) name986 (
		_w992_,
		_w1110_,
		_w1165_
	);
	LUT2 #(
		.INIT('h1)
	) name987 (
		_w1163_,
		_w1164_,
		_w1166_
	);
	LUT2 #(
		.INIT('h4)
	) name988 (
		_w1162_,
		_w1166_,
		_w1167_
	);
	LUT2 #(
		.INIT('h4)
	) name989 (
		_w1165_,
		_w1167_,
		_w1168_
	);
	LUT2 #(
		.INIT('h2)
	) name990 (
		\926(624)_pad ,
		_w1168_,
		_w1169_
	);
	LUT2 #(
		.INIT('h4)
	) name991 (
		_w1006_,
		_w1116_,
		_w1170_
	);
	LUT2 #(
		.INIT('h8)
	) name992 (
		\158(71)_pad ,
		_w1112_,
		_w1171_
	);
	LUT2 #(
		.INIT('h8)
	) name993 (
		\188(81)_pad ,
		_w1114_,
		_w1172_
	);
	LUT2 #(
		.INIT('h4)
	) name994 (
		_w1028_,
		_w1110_,
		_w1173_
	);
	LUT2 #(
		.INIT('h1)
	) name995 (
		_w1171_,
		_w1172_,
		_w1174_
	);
	LUT2 #(
		.INIT('h4)
	) name996 (
		_w1170_,
		_w1174_,
		_w1175_
	);
	LUT2 #(
		.INIT('h4)
	) name997 (
		_w1173_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h2)
	) name998 (
		\926(624)_pad ,
		_w1176_,
		_w1177_
	);
	LUT2 #(
		.INIT('h4)
	) name999 (
		_w1042_,
		_w1116_,
		_w1178_
	);
	LUT2 #(
		.INIT('h8)
	) name1000 (
		\152(69)_pad ,
		_w1112_,
		_w1179_
	);
	LUT2 #(
		.INIT('h8)
	) name1001 (
		\155(70)_pad ,
		_w1114_,
		_w1180_
	);
	LUT2 #(
		.INIT('h4)
	) name1002 (
		_w1064_,
		_w1110_,
		_w1181_
	);
	LUT2 #(
		.INIT('h1)
	) name1003 (
		_w1179_,
		_w1180_,
		_w1182_
	);
	LUT2 #(
		.INIT('h4)
	) name1004 (
		_w1178_,
		_w1182_,
		_w1183_
	);
	LUT2 #(
		.INIT('h4)
	) name1005 (
		_w1181_,
		_w1183_,
		_w1184_
	);
	LUT2 #(
		.INIT('h2)
	) name1006 (
		\926(624)_pad ,
		_w1184_,
		_w1185_
	);
	LUT2 #(
		.INIT('h4)
	) name1007 (
		_w1078_,
		_w1116_,
		_w1186_
	);
	LUT2 #(
		.INIT('h8)
	) name1008 (
		\146(67)_pad ,
		_w1112_,
		_w1187_
	);
	LUT2 #(
		.INIT('h8)
	) name1009 (
		\149(68)_pad ,
		_w1114_,
		_w1188_
	);
	LUT2 #(
		.INIT('h4)
	) name1010 (
		_w1099_,
		_w1110_,
		_w1189_
	);
	LUT2 #(
		.INIT('h1)
	) name1011 (
		_w1187_,
		_w1188_,
		_w1190_
	);
	LUT2 #(
		.INIT('h4)
	) name1012 (
		_w1186_,
		_w1190_,
		_w1191_
	);
	LUT2 #(
		.INIT('h4)
	) name1013 (
		_w1189_,
		_w1191_,
		_w1192_
	);
	LUT2 #(
		.INIT('h2)
	) name1014 (
		\926(624)_pad ,
		_w1192_,
		_w1193_
	);
	LUT2 #(
		.INIT('h1)
	) name1015 (
		\2358(162)_pad ,
		\88(34)_pad ,
		_w1194_
	);
	LUT2 #(
		.INIT('h2)
	) name1016 (
		\2358(162)_pad ,
		\34(12)_pad ,
		_w1195_
	);
	LUT2 #(
		.INIT('h2)
	) name1017 (
		_w469_,
		_w1194_,
		_w1196_
	);
	LUT2 #(
		.INIT('h4)
	) name1018 (
		_w1195_,
		_w1196_,
		_w1197_
	);
	LUT2 #(
		.INIT('h4)
	) name1019 (
		\2358(162)_pad ,
		\79(27)_pad ,
		_w1198_
	);
	LUT2 #(
		.INIT('h8)
	) name1020 (
		\23(6)_pad ,
		\2358(162)_pad ,
		_w1199_
	);
	LUT2 #(
		.INIT('h2)
	) name1021 (
		_w469_,
		_w1198_,
		_w1200_
	);
	LUT2 #(
		.INIT('h4)
	) name1022 (
		_w1199_,
		_w1200_,
		_w1201_
	);
	LUT2 #(
		.INIT('h2)
	) name1023 (
		\144(354)_pad ,
		_w1201_,
		_w1202_
	);
	LUT2 #(
		.INIT('h2)
	) name1024 (
		\4089(173)_pad ,
		\4090(174)_pad ,
		_w1203_
	);
	LUT2 #(
		.INIT('h4)
	) name1025 (
		_w658_,
		_w1203_,
		_w1204_
	);
	LUT2 #(
		.INIT('h8)
	) name1026 (
		\4089(173)_pad ,
		\4090(174)_pad ,
		_w1205_
	);
	LUT2 #(
		.INIT('h8)
	) name1027 (
		\106(40)_pad ,
		_w1205_,
		_w1206_
	);
	LUT2 #(
		.INIT('h4)
	) name1028 (
		\4089(173)_pad ,
		\4090(174)_pad ,
		_w1207_
	);
	LUT2 #(
		.INIT('h8)
	) name1029 (
		\109(41)_pad ,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h1)
	) name1030 (
		\4089(173)_pad ,
		\4090(174)_pad ,
		_w1209_
	);
	LUT2 #(
		.INIT('h4)
	) name1031 (
		_w669_,
		_w1209_,
		_w1210_
	);
	LUT2 #(
		.INIT('h1)
	) name1032 (
		_w1206_,
		_w1208_,
		_w1211_
	);
	LUT2 #(
		.INIT('h4)
	) name1033 (
		_w1204_,
		_w1211_,
		_w1212_
	);
	LUT2 #(
		.INIT('h4)
	) name1034 (
		_w1210_,
		_w1212_,
		_w1213_
	);
	LUT2 #(
		.INIT('h4)
	) name1035 (
		\2358(162)_pad ,
		\82(30)_pad ,
		_w1214_
	);
	LUT2 #(
		.INIT('h8)
	) name1036 (
		\2358(162)_pad ,
		\80(28)_pad ,
		_w1215_
	);
	LUT2 #(
		.INIT('h2)
	) name1037 (
		_w469_,
		_w1214_,
		_w1216_
	);
	LUT2 #(
		.INIT('h4)
	) name1038 (
		_w1215_,
		_w1216_,
		_w1217_
	);
	LUT2 #(
		.INIT('h2)
	) name1039 (
		\144(354)_pad ,
		_w1217_,
		_w1218_
	);
	LUT2 #(
		.INIT('h1)
	) name1040 (
		\4087(171)_pad ,
		\4088(172)_pad ,
		_w1219_
	);
	LUT2 #(
		.INIT('h4)
	) name1041 (
		_w972_,
		_w1219_,
		_w1220_
	);
	LUT2 #(
		.INIT('h8)
	) name1042 (
		\4087(171)_pad ,
		\4088(172)_pad ,
		_w1221_
	);
	LUT2 #(
		.INIT('h8)
	) name1043 (
		\61(21)_pad ,
		_w1221_,
		_w1222_
	);
	LUT2 #(
		.INIT('h2)
	) name1044 (
		\4087(171)_pad ,
		\4088(172)_pad ,
		_w1223_
	);
	LUT2 #(
		.INIT('h8)
	) name1045 (
		\11(2)_pad ,
		_w1223_,
		_w1224_
	);
	LUT2 #(
		.INIT('h4)
	) name1046 (
		\4087(171)_pad ,
		\4088(172)_pad ,
		_w1225_
	);
	LUT2 #(
		.INIT('h4)
	) name1047 (
		_w992_,
		_w1225_,
		_w1226_
	);
	LUT2 #(
		.INIT('h1)
	) name1048 (
		_w1222_,
		_w1224_,
		_w1227_
	);
	LUT2 #(
		.INIT('h4)
	) name1049 (
		_w1220_,
		_w1227_,
		_w1228_
	);
	LUT2 #(
		.INIT('h4)
	) name1050 (
		_w1226_,
		_w1228_,
		_w1229_
	);
	LUT2 #(
		.INIT('h4)
	) name1051 (
		_w658_,
		_w1225_,
		_w1230_
	);
	LUT2 #(
		.INIT('h8)
	) name1052 (
		\106(40)_pad ,
		_w1221_,
		_w1231_
	);
	LUT2 #(
		.INIT('h8)
	) name1053 (
		\109(41)_pad ,
		_w1223_,
		_w1232_
	);
	LUT2 #(
		.INIT('h4)
	) name1054 (
		_w669_,
		_w1219_,
		_w1233_
	);
	LUT2 #(
		.INIT('h1)
	) name1055 (
		_w1231_,
		_w1232_,
		_w1234_
	);
	LUT2 #(
		.INIT('h4)
	) name1056 (
		_w1230_,
		_w1234_,
		_w1235_
	);
	LUT2 #(
		.INIT('h4)
	) name1057 (
		_w1233_,
		_w1235_,
		_w1236_
	);
	LUT2 #(
		.INIT('h4)
	) name1058 (
		_w619_,
		_w1225_,
		_w1237_
	);
	LUT2 #(
		.INIT('h8)
	) name1059 (
		\49(17)_pad ,
		_w1221_,
		_w1238_
	);
	LUT2 #(
		.INIT('h8)
	) name1060 (
		\46(16)_pad ,
		_w1223_,
		_w1239_
	);
	LUT2 #(
		.INIT('h4)
	) name1061 (
		_w632_,
		_w1219_,
		_w1240_
	);
	LUT2 #(
		.INIT('h1)
	) name1062 (
		_w1238_,
		_w1239_,
		_w1241_
	);
	LUT2 #(
		.INIT('h4)
	) name1063 (
		_w1237_,
		_w1241_,
		_w1242_
	);
	LUT2 #(
		.INIT('h4)
	) name1064 (
		_w1240_,
		_w1242_,
		_w1243_
	);
	LUT2 #(
		.INIT('h4)
	) name1065 (
		_w580_,
		_w1225_,
		_w1244_
	);
	LUT2 #(
		.INIT('h8)
	) name1066 (
		\103(39)_pad ,
		_w1221_,
		_w1245_
	);
	LUT2 #(
		.INIT('h8)
	) name1067 (
		\100(38)_pad ,
		_w1223_,
		_w1246_
	);
	LUT2 #(
		.INIT('h4)
	) name1068 (
		_w594_,
		_w1219_,
		_w1247_
	);
	LUT2 #(
		.INIT('h1)
	) name1069 (
		_w1245_,
		_w1246_,
		_w1248_
	);
	LUT2 #(
		.INIT('h4)
	) name1070 (
		_w1244_,
		_w1248_,
		_w1249_
	);
	LUT2 #(
		.INIT('h4)
	) name1071 (
		_w1247_,
		_w1249_,
		_w1250_
	);
	LUT2 #(
		.INIT('h4)
	) name1072 (
		_w544_,
		_w1225_,
		_w1251_
	);
	LUT2 #(
		.INIT('h8)
	) name1073 (
		\40(14)_pad ,
		_w1221_,
		_w1252_
	);
	LUT2 #(
		.INIT('h8)
	) name1074 (
		\91(35)_pad ,
		_w1223_,
		_w1253_
	);
	LUT2 #(
		.INIT('h4)
	) name1075 (
		_w556_,
		_w1219_,
		_w1254_
	);
	LUT2 #(
		.INIT('h1)
	) name1076 (
		_w1252_,
		_w1253_,
		_w1255_
	);
	LUT2 #(
		.INIT('h4)
	) name1077 (
		_w1251_,
		_w1255_,
		_w1256_
	);
	LUT2 #(
		.INIT('h4)
	) name1078 (
		_w1254_,
		_w1256_,
		_w1257_
	);
	LUT2 #(
		.INIT('h4)
	) name1079 (
		_w502_,
		_w1225_,
		_w1258_
	);
	LUT2 #(
		.INIT('h8)
	) name1080 (
		\37(13)_pad ,
		_w1221_,
		_w1259_
	);
	LUT2 #(
		.INIT('h8)
	) name1081 (
		\43(15)_pad ,
		_w1223_,
		_w1260_
	);
	LUT2 #(
		.INIT('h4)
	) name1082 (
		_w519_,
		_w1219_,
		_w1261_
	);
	LUT2 #(
		.INIT('h1)
	) name1083 (
		_w1259_,
		_w1260_,
		_w1262_
	);
	LUT2 #(
		.INIT('h4)
	) name1084 (
		_w1258_,
		_w1262_,
		_w1263_
	);
	LUT2 #(
		.INIT('h4)
	) name1085 (
		_w1261_,
		_w1263_,
		_w1264_
	);
	LUT2 #(
		.INIT('h4)
	) name1086 (
		_w1078_,
		_w1219_,
		_w1265_
	);
	LUT2 #(
		.INIT('h8)
	) name1087 (
		\20(5)_pad ,
		_w1221_,
		_w1266_
	);
	LUT2 #(
		.INIT('h8)
	) name1088 (
		\76(26)_pad ,
		_w1223_,
		_w1267_
	);
	LUT2 #(
		.INIT('h4)
	) name1089 (
		_w1099_,
		_w1225_,
		_w1268_
	);
	LUT2 #(
		.INIT('h1)
	) name1090 (
		_w1266_,
		_w1267_,
		_w1269_
	);
	LUT2 #(
		.INIT('h4)
	) name1091 (
		_w1265_,
		_w1269_,
		_w1270_
	);
	LUT2 #(
		.INIT('h4)
	) name1092 (
		_w1268_,
		_w1270_,
		_w1271_
	);
	LUT2 #(
		.INIT('h4)
	) name1093 (
		_w1042_,
		_w1219_,
		_w1272_
	);
	LUT2 #(
		.INIT('h8)
	) name1094 (
		\17(4)_pad ,
		_w1221_,
		_w1273_
	);
	LUT2 #(
		.INIT('h8)
	) name1095 (
		\73(25)_pad ,
		_w1223_,
		_w1274_
	);
	LUT2 #(
		.INIT('h4)
	) name1096 (
		_w1064_,
		_w1225_,
		_w1275_
	);
	LUT2 #(
		.INIT('h1)
	) name1097 (
		_w1273_,
		_w1274_,
		_w1276_
	);
	LUT2 #(
		.INIT('h4)
	) name1098 (
		_w1272_,
		_w1276_,
		_w1277_
	);
	LUT2 #(
		.INIT('h4)
	) name1099 (
		_w1275_,
		_w1277_,
		_w1278_
	);
	LUT2 #(
		.INIT('h4)
	) name1100 (
		_w1006_,
		_w1219_,
		_w1279_
	);
	LUT2 #(
		.INIT('h8)
	) name1101 (
		\70(24)_pad ,
		_w1221_,
		_w1280_
	);
	LUT2 #(
		.INIT('h8)
	) name1102 (
		\67(23)_pad ,
		_w1223_,
		_w1281_
	);
	LUT2 #(
		.INIT('h4)
	) name1103 (
		_w1028_,
		_w1225_,
		_w1282_
	);
	LUT2 #(
		.INIT('h1)
	) name1104 (
		_w1280_,
		_w1281_,
		_w1283_
	);
	LUT2 #(
		.INIT('h4)
	) name1105 (
		_w1279_,
		_w1283_,
		_w1284_
	);
	LUT2 #(
		.INIT('h4)
	) name1106 (
		_w1282_,
		_w1284_,
		_w1285_
	);
	LUT2 #(
		.INIT('h4)
	) name1107 (
		_w957_,
		_w1219_,
		_w1286_
	);
	LUT2 #(
		.INIT('h8)
	) name1108 (
		\64(22)_pad ,
		_w1221_,
		_w1287_
	);
	LUT2 #(
		.INIT('h8)
	) name1109 (
		\14(3)_pad ,
		_w1223_,
		_w1288_
	);
	LUT2 #(
		.INIT('h4)
	) name1110 (
		_w842_,
		_w1225_,
		_w1289_
	);
	LUT2 #(
		.INIT('h1)
	) name1111 (
		_w1287_,
		_w1288_,
		_w1290_
	);
	LUT2 #(
		.INIT('h4)
	) name1112 (
		_w1286_,
		_w1290_,
		_w1291_
	);
	LUT2 #(
		.INIT('h4)
	) name1113 (
		_w1289_,
		_w1291_,
		_w1292_
	);
	LUT2 #(
		.INIT('h4)
	) name1114 (
		_w619_,
		_w1203_,
		_w1293_
	);
	LUT2 #(
		.INIT('h8)
	) name1115 (
		\49(17)_pad ,
		_w1205_,
		_w1294_
	);
	LUT2 #(
		.INIT('h8)
	) name1116 (
		\46(16)_pad ,
		_w1207_,
		_w1295_
	);
	LUT2 #(
		.INIT('h4)
	) name1117 (
		_w632_,
		_w1209_,
		_w1296_
	);
	LUT2 #(
		.INIT('h1)
	) name1118 (
		_w1294_,
		_w1295_,
		_w1297_
	);
	LUT2 #(
		.INIT('h4)
	) name1119 (
		_w1293_,
		_w1297_,
		_w1298_
	);
	LUT2 #(
		.INIT('h4)
	) name1120 (
		_w1296_,
		_w1298_,
		_w1299_
	);
	LUT2 #(
		.INIT('h4)
	) name1121 (
		_w580_,
		_w1203_,
		_w1300_
	);
	LUT2 #(
		.INIT('h8)
	) name1122 (
		\103(39)_pad ,
		_w1205_,
		_w1301_
	);
	LUT2 #(
		.INIT('h8)
	) name1123 (
		\100(38)_pad ,
		_w1207_,
		_w1302_
	);
	LUT2 #(
		.INIT('h4)
	) name1124 (
		_w594_,
		_w1209_,
		_w1303_
	);
	LUT2 #(
		.INIT('h1)
	) name1125 (
		_w1301_,
		_w1302_,
		_w1304_
	);
	LUT2 #(
		.INIT('h4)
	) name1126 (
		_w1300_,
		_w1304_,
		_w1305_
	);
	LUT2 #(
		.INIT('h4)
	) name1127 (
		_w1303_,
		_w1305_,
		_w1306_
	);
	LUT2 #(
		.INIT('h4)
	) name1128 (
		_w544_,
		_w1203_,
		_w1307_
	);
	LUT2 #(
		.INIT('h8)
	) name1129 (
		\40(14)_pad ,
		_w1205_,
		_w1308_
	);
	LUT2 #(
		.INIT('h8)
	) name1130 (
		\91(35)_pad ,
		_w1207_,
		_w1309_
	);
	LUT2 #(
		.INIT('h4)
	) name1131 (
		_w556_,
		_w1209_,
		_w1310_
	);
	LUT2 #(
		.INIT('h1)
	) name1132 (
		_w1308_,
		_w1309_,
		_w1311_
	);
	LUT2 #(
		.INIT('h4)
	) name1133 (
		_w1307_,
		_w1311_,
		_w1312_
	);
	LUT2 #(
		.INIT('h4)
	) name1134 (
		_w1310_,
		_w1312_,
		_w1313_
	);
	LUT2 #(
		.INIT('h4)
	) name1135 (
		_w502_,
		_w1203_,
		_w1314_
	);
	LUT2 #(
		.INIT('h8)
	) name1136 (
		\37(13)_pad ,
		_w1205_,
		_w1315_
	);
	LUT2 #(
		.INIT('h8)
	) name1137 (
		\43(15)_pad ,
		_w1207_,
		_w1316_
	);
	LUT2 #(
		.INIT('h4)
	) name1138 (
		_w519_,
		_w1209_,
		_w1317_
	);
	LUT2 #(
		.INIT('h1)
	) name1139 (
		_w1315_,
		_w1316_,
		_w1318_
	);
	LUT2 #(
		.INIT('h4)
	) name1140 (
		_w1314_,
		_w1318_,
		_w1319_
	);
	LUT2 #(
		.INIT('h4)
	) name1141 (
		_w1317_,
		_w1319_,
		_w1320_
	);
	LUT2 #(
		.INIT('h4)
	) name1142 (
		_w1078_,
		_w1209_,
		_w1321_
	);
	LUT2 #(
		.INIT('h8)
	) name1143 (
		\20(5)_pad ,
		_w1205_,
		_w1322_
	);
	LUT2 #(
		.INIT('h8)
	) name1144 (
		\76(26)_pad ,
		_w1207_,
		_w1323_
	);
	LUT2 #(
		.INIT('h4)
	) name1145 (
		_w1099_,
		_w1203_,
		_w1324_
	);
	LUT2 #(
		.INIT('h1)
	) name1146 (
		_w1322_,
		_w1323_,
		_w1325_
	);
	LUT2 #(
		.INIT('h4)
	) name1147 (
		_w1321_,
		_w1325_,
		_w1326_
	);
	LUT2 #(
		.INIT('h4)
	) name1148 (
		_w1324_,
		_w1326_,
		_w1327_
	);
	LUT2 #(
		.INIT('h4)
	) name1149 (
		_w1042_,
		_w1209_,
		_w1328_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		\17(4)_pad ,
		_w1205_,
		_w1329_
	);
	LUT2 #(
		.INIT('h8)
	) name1151 (
		\73(25)_pad ,
		_w1207_,
		_w1330_
	);
	LUT2 #(
		.INIT('h4)
	) name1152 (
		_w1064_,
		_w1203_,
		_w1331_
	);
	LUT2 #(
		.INIT('h1)
	) name1153 (
		_w1329_,
		_w1330_,
		_w1332_
	);
	LUT2 #(
		.INIT('h4)
	) name1154 (
		_w1328_,
		_w1332_,
		_w1333_
	);
	LUT2 #(
		.INIT('h4)
	) name1155 (
		_w1331_,
		_w1333_,
		_w1334_
	);
	LUT2 #(
		.INIT('h4)
	) name1156 (
		_w1006_,
		_w1209_,
		_w1335_
	);
	LUT2 #(
		.INIT('h8)
	) name1157 (
		\70(24)_pad ,
		_w1205_,
		_w1336_
	);
	LUT2 #(
		.INIT('h8)
	) name1158 (
		\67(23)_pad ,
		_w1207_,
		_w1337_
	);
	LUT2 #(
		.INIT('h4)
	) name1159 (
		_w1028_,
		_w1203_,
		_w1338_
	);
	LUT2 #(
		.INIT('h1)
	) name1160 (
		_w1336_,
		_w1337_,
		_w1339_
	);
	LUT2 #(
		.INIT('h4)
	) name1161 (
		_w1335_,
		_w1339_,
		_w1340_
	);
	LUT2 #(
		.INIT('h4)
	) name1162 (
		_w1338_,
		_w1340_,
		_w1341_
	);
	LUT2 #(
		.INIT('h4)
	) name1163 (
		_w957_,
		_w1209_,
		_w1342_
	);
	LUT2 #(
		.INIT('h8)
	) name1164 (
		\64(22)_pad ,
		_w1205_,
		_w1343_
	);
	LUT2 #(
		.INIT('h8)
	) name1165 (
		\14(3)_pad ,
		_w1207_,
		_w1344_
	);
	LUT2 #(
		.INIT('h4)
	) name1166 (
		_w842_,
		_w1203_,
		_w1345_
	);
	LUT2 #(
		.INIT('h1)
	) name1167 (
		_w1343_,
		_w1344_,
		_w1346_
	);
	LUT2 #(
		.INIT('h4)
	) name1168 (
		_w1342_,
		_w1346_,
		_w1347_
	);
	LUT2 #(
		.INIT('h4)
	) name1169 (
		_w1345_,
		_w1347_,
		_w1348_
	);
	LUT2 #(
		.INIT('h8)
	) name1170 (
		\144(354)_pad ,
		\145(66)_pad ,
		_w1349_
	);
	LUT2 #(
		.INIT('h2)
	) name1171 (
		\132(60)_pad ,
		_w627_,
		_w1350_
	);
	LUT2 #(
		.INIT('h4)
	) name1172 (
		\132(60)_pad ,
		_w627_,
		_w1351_
	);
	LUT2 #(
		.INIT('h1)
	) name1173 (
		_w1350_,
		_w1351_,
		_w1352_
	);
	LUT2 #(
		.INIT('h2)
	) name1174 (
		\136(62)_pad ,
		\973(202)_pad ,
		_w1353_
	);
	LUT2 #(
		.INIT('h8)
	) name1175 (
		\83(31)_pad ,
		_w469_,
		_w1354_
	);
	LUT2 #(
		.INIT('h8)
	) name1176 (
		_w491_,
		_w900_,
		_w1355_
	);
	LUT2 #(
		.INIT('h1)
	) name1177 (
		_w499_,
		_w955_,
		_w1356_
	);
	LUT2 #(
		.INIT('h8)
	) name1178 (
		\120(50)_pad ,
		_w499_,
		_w1357_
	);
	LUT2 #(
		.INIT('h1)
	) name1179 (
		_w1356_,
		_w1357_,
		_w1358_
	);
	LUT2 #(
		.INIT('h4)
	) name1180 (
		_w1355_,
		_w1358_,
		_w1359_
	);
	LUT2 #(
		.INIT('h2)
	) name1181 (
		\27(10)_pad ,
		\2824(163)_pad ,
		_w1360_
	);
	LUT2 #(
		.INIT('h8)
	) name1182 (
		\386(135)_pad ,
		\556(153)_pad ,
		_w1361_
	);
	LUT2 #(
		.INIT('h2)
	) name1183 (
		_w394_,
		_w422_,
		_w1362_
	);
	LUT2 #(
		.INIT('h4)
	) name1184 (
		_w394_,
		_w422_,
		_w1363_
	);
	LUT2 #(
		.INIT('h1)
	) name1185 (
		_w1362_,
		_w1363_,
		_w1364_
	);
	LUT2 #(
		.INIT('h4)
	) name1186 (
		\332(122)_pad ,
		\369(131)_pad ,
		_w1365_
	);
	LUT2 #(
		.INIT('h8)
	) name1187 (
		\332(122)_pad ,
		\372(132)_pad ,
		_w1366_
	);
	LUT2 #(
		.INIT('h1)
	) name1188 (
		_w1365_,
		_w1366_,
		_w1367_
	);
	LUT2 #(
		.INIT('h2)
	) name1189 (
		_w426_,
		_w1367_,
		_w1368_
	);
	LUT2 #(
		.INIT('h4)
	) name1190 (
		_w426_,
		_w1367_,
		_w1369_
	);
	LUT2 #(
		.INIT('h1)
	) name1191 (
		_w1368_,
		_w1369_,
		_w1370_
	);
	LUT2 #(
		.INIT('h2)
	) name1192 (
		_w1364_,
		_w1370_,
		_w1371_
	);
	LUT2 #(
		.INIT('h4)
	) name1193 (
		_w1364_,
		_w1370_,
		_w1372_
	);
	LUT2 #(
		.INIT('h1)
	) name1194 (
		_w1371_,
		_w1372_,
		_w1373_
	);
	LUT2 #(
		.INIT('h1)
	) name1195 (
		_w407_,
		_w419_,
		_w1374_
	);
	LUT2 #(
		.INIT('h8)
	) name1196 (
		_w407_,
		_w419_,
		_w1375_
	);
	LUT2 #(
		.INIT('h1)
	) name1197 (
		_w1374_,
		_w1375_,
		_w1376_
	);
	LUT2 #(
		.INIT('h2)
	) name1198 (
		_w400_,
		_w1376_,
		_w1377_
	);
	LUT2 #(
		.INIT('h4)
	) name1199 (
		_w400_,
		_w1376_,
		_w1378_
	);
	LUT2 #(
		.INIT('h1)
	) name1200 (
		_w1377_,
		_w1378_,
		_w1379_
	);
	LUT2 #(
		.INIT('h8)
	) name1201 (
		_w432_,
		_w1379_,
		_w1380_
	);
	LUT2 #(
		.INIT('h1)
	) name1202 (
		_w432_,
		_w1379_,
		_w1381_
	);
	LUT2 #(
		.INIT('h1)
	) name1203 (
		_w1380_,
		_w1381_,
		_w1382_
	);
	LUT2 #(
		.INIT('h4)
	) name1204 (
		_w388_,
		_w412_,
		_w1383_
	);
	LUT2 #(
		.INIT('h4)
	) name1205 (
		\331(121)_pad ,
		_w388_,
		_w1384_
	);
	LUT2 #(
		.INIT('h1)
	) name1206 (
		_w1383_,
		_w1384_,
		_w1385_
	);
	LUT2 #(
		.INIT('h2)
	) name1207 (
		_w1382_,
		_w1385_,
		_w1386_
	);
	LUT2 #(
		.INIT('h4)
	) name1208 (
		_w1382_,
		_w1385_,
		_w1387_
	);
	LUT2 #(
		.INIT('h1)
	) name1209 (
		_w1386_,
		_w1387_,
		_w1388_
	);
	LUT2 #(
		.INIT('h8)
	) name1210 (
		_w1373_,
		_w1388_,
		_w1389_
	);
	LUT2 #(
		.INIT('h1)
	) name1211 (
		_w1373_,
		_w1388_,
		_w1390_
	);
	LUT2 #(
		.INIT('h1)
	) name1212 (
		_w1389_,
		_w1390_,
		_w1391_
	);
	LUT2 #(
		.INIT('h8)
	) name1213 (
		\245(98)_pad ,
		\559(154)_pad ,
		_w1392_
	);
	LUT2 #(
		.INIT('h8)
	) name1214 (
		_w387_,
		_w1392_,
		_w1393_
	);
	LUT2 #(
		.INIT('h8)
	) name1215 (
		_w1361_,
		_w1393_,
		_w1394_
	);
	LUT2 #(
		.INIT('h8)
	) name1216 (
		_w259_,
		_w1394_,
		_w1395_
	);
	LUT2 #(
		.INIT('h8)
	) name1217 (
		_w286_,
		_w1395_,
		_w1396_
	);
	LUT2 #(
		.INIT('h4)
	) name1218 (
		_w235_,
		_w1396_,
		_w1397_
	);
	LUT2 #(
		.INIT('h8)
	) name1219 (
		_w1391_,
		_w1397_,
		_w1398_
	);
	LUT2 #(
		.INIT('h4)
	) name1220 (
		_w972_,
		_w1209_,
		_w1399_
	);
	LUT2 #(
		.INIT('h8)
	) name1221 (
		\61(21)_pad ,
		_w1205_,
		_w1400_
	);
	LUT2 #(
		.INIT('h8)
	) name1222 (
		\11(2)_pad ,
		_w1207_,
		_w1401_
	);
	LUT2 #(
		.INIT('h4)
	) name1223 (
		_w992_,
		_w1203_,
		_w1402_
	);
	LUT2 #(
		.INIT('h1)
	) name1224 (
		_w1400_,
		_w1401_,
		_w1403_
	);
	LUT2 #(
		.INIT('h4)
	) name1225 (
		_w1399_,
		_w1403_,
		_w1404_
	);
	LUT2 #(
		.INIT('h4)
	) name1226 (
		_w1402_,
		_w1404_,
		_w1405_
	);
	LUT2 #(
		.INIT('h8)
	) name1227 (
		_w491_,
		_w741_,
		_w1406_
	);
	LUT2 #(
		.INIT('h1)
	) name1228 (
		_w499_,
		_w840_,
		_w1407_
	);
	LUT2 #(
		.INIT('h8)
	) name1229 (
		\118(48)_pad ,
		_w499_,
		_w1408_
	);
	LUT2 #(
		.INIT('h1)
	) name1230 (
		_w1407_,
		_w1408_,
		_w1409_
	);
	LUT2 #(
		.INIT('h4)
	) name1231 (
		_w1406_,
		_w1409_,
		_w1410_
	);
	LUT2 #(
		.INIT('h8)
	) name1232 (
		\135(61)_pad ,
		\4115(177)_pad ,
		_w1411_
	);
	LUT2 #(
		.INIT('h1)
	) name1233 (
		\3724(170)_pad ,
		_w373_,
		_w1412_
	);
	LUT2 #(
		.INIT('h2)
	) name1234 (
		\132(60)_pad ,
		_w419_,
		_w1413_
	);
	LUT2 #(
		.INIT('h4)
	) name1235 (
		\132(60)_pad ,
		_w419_,
		_w1414_
	);
	LUT2 #(
		.INIT('h1)
	) name1236 (
		_w1413_,
		_w1414_,
		_w1415_
	);
	LUT2 #(
		.INIT('h2)
	) name1237 (
		\3724(170)_pad ,
		_w1415_,
		_w1416_
	);
	LUT2 #(
		.INIT('h1)
	) name1238 (
		\3717(169)_pad ,
		_w1412_,
		_w1417_
	);
	LUT2 #(
		.INIT('h4)
	) name1239 (
		_w1416_,
		_w1417_,
		_w1418_
	);
	LUT2 #(
		.INIT('h2)
	) name1240 (
		\123(53)_pad ,
		\3724(170)_pad ,
		_w1419_
	);
	LUT2 #(
		.INIT('h8)
	) name1241 (
		\3724(170)_pad ,
		_w666_,
		_w1420_
	);
	LUT2 #(
		.INIT('h2)
	) name1242 (
		\3717(169)_pad ,
		_w1419_,
		_w1421_
	);
	LUT2 #(
		.INIT('h4)
	) name1243 (
		_w1420_,
		_w1421_,
		_w1422_
	);
	LUT2 #(
		.INIT('h1)
	) name1244 (
		_w1411_,
		_w1418_,
		_w1423_
	);
	LUT2 #(
		.INIT('h4)
	) name1245 (
		_w1422_,
		_w1423_,
		_w1424_
	);
	LUT2 #(
		.INIT('h1)
	) name1246 (
		_w574_,
		_w988_,
		_w1425_
	);
	LUT2 #(
		.INIT('h4)
	) name1247 (
		_w1024_,
		_w1425_,
		_w1426_
	);
	LUT2 #(
		.INIT('h4)
	) name1248 (
		_w1060_,
		_w1426_,
		_w1427_
	);
	LUT2 #(
		.INIT('h8)
	) name1249 (
		_w1095_,
		_w1427_,
		_w1428_
	);
	LUT2 #(
		.INIT('h8)
	) name1250 (
		_w497_,
		_w1428_,
		_w1429_
	);
	LUT2 #(
		.INIT('h8)
	) name1251 (
		_w540_,
		_w1429_,
		_w1430_
	);
	LUT2 #(
		.INIT('h4)
	) name1252 (
		_w615_,
		_w1430_,
		_w1431_
	);
	LUT2 #(
		.INIT('h4)
	) name1253 (
		_w654_,
		_w1431_,
		_w1432_
	);
	LUT2 #(
		.INIT('h8)
	) name1254 (
		_w403_,
		_w968_,
		_w1433_
	);
	LUT2 #(
		.INIT('h4)
	) name1255 (
		_w588_,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('h8)
	) name1256 (
		_w1038_,
		_w1434_,
		_w1435_
	);
	LUT2 #(
		.INIT('h8)
	) name1257 (
		_w1074_,
		_w1435_,
		_w1436_
	);
	LUT2 #(
		.INIT('h4)
	) name1258 (
		_w515_,
		_w1436_,
		_w1437_
	);
	LUT2 #(
		.INIT('h8)
	) name1259 (
		_w552_,
		_w1437_,
		_w1438_
	);
	LUT2 #(
		.INIT('h8)
	) name1260 (
		_w628_,
		_w1438_,
		_w1439_
	);
	LUT2 #(
		.INIT('h4)
	) name1261 (
		_w666_,
		_w1439_,
		_w1440_
	);
	LUT2 #(
		.INIT('h1)
	) name1262 (
		_w489_,
		_w533_,
		_w1441_
	);
	LUT2 #(
		.INIT('h1)
	) name1263 (
		_w570_,
		_w608_,
		_w1442_
	);
	LUT2 #(
		.INIT('h1)
	) name1264 (
		_w646_,
		_w984_,
		_w1443_
	);
	LUT2 #(
		.INIT('h1)
	) name1265 (
		_w1018_,
		_w1054_,
		_w1444_
	);
	LUT2 #(
		.INIT('h4)
	) name1266 (
		_w1090_,
		_w1444_,
		_w1445_
	);
	LUT2 #(
		.INIT('h8)
	) name1267 (
		_w1442_,
		_w1443_,
		_w1446_
	);
	LUT2 #(
		.INIT('h8)
	) name1268 (
		_w1441_,
		_w1446_,
		_w1447_
	);
	LUT2 #(
		.INIT('h8)
	) name1269 (
		_w1445_,
		_w1447_,
		_w1448_
	);
	assign \1000(2168)_pad  = _w235_ ;
	assign \1002(1920)_pad  = _w259_ ;
	assign \1004(1977)_pad  = _w286_ ;
	assign \588(1696)_pad  = _w321_ ;
	assign \593(733)_pad  = \889(734)_pad ;
	assign \598(1623)_pad  = _w386_ ;
	assign \599(269)_pad  = \348(126)_pad ;
	assign \600(259)_pad  = \366(130)_pad ;
	assign \601(220)_pad  = _w387_ ;
	assign \604(223)_pad  = \545(150)_pad ;
	assign \606(407)_pad  = \892(408)_pad ;
	assign \611(275)_pad  = \338(124)_pad ;
	assign \612(263)_pad  = \358(128)_pad ;
	assign \615(1750)_pad  = _w438_ ;
	assign \618(1925)_pad  = _w451_ ;
	assign \621(1893)_pad  = _w467_ ;
	assign \626(1752)_pad  = _w438_ ;
	assign \632(1692)_pad  = _w321_ ;
	assign \634(665)_pad  = _w468_ ;
	assign \636(1280)_pad  = _w473_ ;
	assign \639(1275)_pad  = _w478_ ;
	assign \642(2222)_pad  = _w524_ ;
	assign \645(2271)_pad  = _w561_ ;
	assign \648(2295)_pad  = _w599_ ;
	assign \651(2314)_pad  = _w637_ ;
	assign \654(2315)_pad  = _w674_ ;
	assign \656(621)_pad  = _w675_ ;
	assign \658(2483)_pad  = _w964_ ;
	assign \661(2178)_pad  = _w997_ ;
	assign \664(2223)_pad  = _w1033_ ;
	assign \667(2224)_pad  = _w1069_ ;
	assign \670(2225)_pad  = _w1104_ ;
	assign \673(1276)_pad  = _w1109_ ;
	assign \676(2229)_pad  = _w1121_ ;
	assign \679(2272)_pad  = _w1129_ ;
	assign \682(2296)_pad  = _w1137_ ;
	assign \685(2316)_pad  = _w1145_ ;
	assign \688(2317)_pad  = _w1153_ ;
	assign \690(2484)_pad  = _w1161_ ;
	assign \693(2179)_pad  = _w1169_ ;
	assign \696(2226)_pad  = _w1177_ ;
	assign \699(2227)_pad  = _w1185_ ;
	assign \702(2228)_pad  = _w1193_ ;
	assign \704(1281)_pad  = _w1197_ ;
	assign \707(1277)_pad  = _w1202_ ;
	assign \712(2297)_pad  = _w1213_ ;
	assign \715(1278)_pad  = _w1218_ ;
	assign \722(2131)_pad  = _w1229_ ;
	assign \727(2298)_pad  = _w1236_ ;
	assign \732(2300)_pad  = _w1243_ ;
	assign \737(2279)_pad  = _w1250_ ;
	assign \742(2238)_pad  = _w1257_ ;
	assign \747(2187)_pad  = _w1264_ ;
	assign \752(2189)_pad  = _w1271_ ;
	assign \757(2190)_pad  = _w1278_ ;
	assign \762(2184)_pad  = _w1285_ ;
	assign \767(2479)_pad  = _w1292_ ;
	assign \772(2299)_pad  = _w1299_ ;
	assign \777(2278)_pad  = _w1306_ ;
	assign \782(2239)_pad  = _w1313_ ;
	assign \787(2186)_pad  = _w1320_ ;
	assign \792(2188)_pad  = _w1327_ ;
	assign \797(2191)_pad  = _w1334_ ;
	assign \802(2183)_pad  = _w1341_ ;
	assign \807(2480)_pad  = _w1348_ ;
	assign \809(655)_pad  = _w469_ ;
	assign \810(356)_pad  = _w1349_ ;
	assign \813(2260)_pad  = _w1352_ ;
	assign \815(627)_pad  = _w1353_ ;
	assign \820(1283)_pad  = _w1354_ ;
	assign \822(1933)_pad  = _w972_ ;
	assign \824(2274)_pad  = _w669_ ;
	assign \826(2275)_pad  = _w632_ ;
	assign \828(2233)_pad  = _w594_ ;
	assign \830(2182)_pad  = _w556_ ;
	assign \832(2133)_pad  = _w519_ ;
	assign \834(2123)_pad  = _w1078_ ;
	assign \836(2128)_pad  = _w1042_ ;
	assign \838(2064)_pad  = _w1006_ ;
	assign \843(2455)_pad  = _w1359_ ;
	assign \845(845)_pad  = _w1360_ ;
	assign \847(465)_pad  = _w1361_ ;
	assign \848(330)_pad  = \245(98)_pad ;
	assign \849(219)_pad  = \552(152)_pad ;
	assign \850(217)_pad  = \562(155)_pad ;
	assign \851(218)_pad  = \559(154)_pad ;
	assign \854(2268)_pad  = _w1398_ ;
	assign \859(2132)_pad  = _w1405_ ;
	assign \861(2070)_pad  = _w992_ ;
	assign \863(2276)_pad  = _w658_ ;
	assign \865(2277)_pad  = _w619_ ;
	assign \867(2237)_pad  = _w580_ ;
	assign \869(2181)_pad  = _w544_ ;
	assign \871(2127)_pad  = _w502_ ;
	assign \873(2124)_pad  = _w1099_ ;
	assign \875(2125)_pad  = _w1064_ ;
	assign \877(2126)_pad  = _w1028_ ;
	assign \882(2456)_pad  = _w1410_ ;
	assign \998(2163)_pad  = _w1391_ ;
	assign \u2023_syn_3  = _w1424_ ;
	assign \u2095_syn_3  = _w1432_ ;
	assign \u2109_syn_3  = _w1440_ ;
	assign \u2318_syn_3  = _w666_ ;
	assign \u3086_syn_3  = _w1448_ ;
endmodule;