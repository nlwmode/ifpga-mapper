module top( \100(51)_pad  , \103(52)_pad  , \109(54)_pad  , \110(55)_pad  , \111(56)_pad  , \112(57)_pad  , \113(58)_pad  , \114(59)_pad  , \115(60)_pad  , \118(61)_pad  , \1197(165)_pad  , \12(3)_pad  , \121(62)_pad  , \124(63)_pad  , \127(64)_pad  , \130(65)_pad  , \133(66)_pad  , \134(67)_pad  , \135(68)_pad  , \138(69)_pad  , \141(70)_pad  , \144(71)_pad  , \1455(166)_pad  , \147(72)_pad  , \15(4)_pad  , \150(73)_pad  , \151(74)_pad  , \152(75)_pad  , \153(76)_pad  , \154(77)_pad  , \155(78)_pad  , \156(79)_pad  , \157(80)_pad  , \158(81)_pad  , \159(82)_pad  , \160(83)_pad  , \161(84)_pad  , \162(85)_pad  , \163(86)_pad  , \164(87)_pad  , \165(88)_pad  , \166(89)_pad  , \167(90)_pad  , \168(91)_pad  , \169(92)_pad  , \170(93)_pad  , \171(94)_pad  , \172(95)_pad  , \173(96)_pad  , \174(97)_pad  , \175(98)_pad  , \176(99)_pad  , \177(100)_pad  , \178(101)_pad  , \179(102)_pad  , \18(5)_pad  , \180(103)_pad  , \181(104)_pad  , \182(105)_pad  , \183(106)_pad  , \184(107)_pad  , \185(108)_pad  , \186(109)_pad  , \187(110)_pad  , \188(111)_pad  , \189(112)_pad  , \190(113)_pad  , \191(114)_pad  , \192(115)_pad  , \193(116)_pad  , \194(117)_pad  , \195(118)_pad  , \196(119)_pad  , \197(120)_pad  , \198(121)_pad  , \199(122)_pad  , \200(123)_pad  , \201(124)_pad  , \202(125)_pad  , \203(126)_pad  , \204(127)_pad  , \205(128)_pad  , \206(129)_pad  , \207(130)_pad  , \208(131)_pad  , \209(132)_pad  , \210(133)_pad  , \211(134)_pad  , \212(135)_pad  , \213(136)_pad  , \214(137)_pad  , \215(138)_pad  , \216(139)_pad  , \217(140)_pad  , \218(141)_pad  , \219(142)_pad  , \220(143)_pad  , \2204(174)_pad  , \221(144)_pad  , \222(145)_pad  , \223(146)_pad  , \224(147)_pad  , \225(148)_pad  , \226(149)_pad  , \227(150)_pad  , \228(151)_pad  , \229(152)_pad  , \23(6)_pad  , \230(153)_pad  , \231(154)_pad  , \232(155)_pad  , \233(156)_pad  , \234(157)_pad  , \235(158)_pad  , \236(159)_pad  , \237(160)_pad  , \238(161)_pad  , \239(162)_pad  , \240(163)_pad  , \26(7)_pad  , \29(8)_pad  , \32(9)_pad  , \35(10)_pad  , \38(11)_pad  , \41(12)_pad  , \436(286)_pad  , \438(274)_pad  , \44(13)_pad  , \440(277)_pad  , \442(280)_pad  , \444(282)_pad  , \446(393)_pad  , \448(284)_pad  , \450(288)_pad  , \4526(205)_pad  , \4528(206)_pad  , \453(596)_pad  , \47(14)_pad  , \478(269)_pad  , \480(250)_pad  , \482(253)_pad  , \484(256)_pad  , \486(258)_pad  , \488(260)_pad  , \490(263)_pad  , \492(265)_pad  , \494(267)_pad  , \496(271)_pad  , \5(1)_pad  , \50(15)_pad  , \522(226)_pad  , \524(210)_pad  , \526(212)_pad  , \528(214)_pad  , \53(16)_pad  , \530(216)_pad  , \532(218)_pad  , \534(220)_pad  , \536(222)_pad  , \538(224)_pad  , \54(17)_pad  , \540(227)_pad  , \542(246)_pad  , \544(230)_pad  , \546(232)_pad  , \548(234)_pad  , \55(18)_pad  , \550(236)_pad  , \552(238)_pad  , \554(240)_pad  , \556(242)_pad  , \558(244)_pad  , \56(19)_pad  , \560(248)_pad  , \57(20)_pad  , \58(21)_pad  , \59(22)_pad  , \60(23)_pad  , \61(24)_pad  , \62(25)_pad  , \63(26)_pad  , \64(27)_pad  , \65(28)_pad  , \66(29)_pad  , \69(30)_pad  , \70(31)_pad  , \73(32)_pad  , \74(33)_pad  , \75(34)_pad  , \76(35)_pad  , \77(36)_pad  , \78(37)_pad  , \79(38)_pad  , \80(39)_pad  , \81(40)_pad  , \82(41)_pad  , \83(42)_pad  , \84(43)_pad  , \85(44)_pad  , \86(45)_pad  , \87(46)_pad  , \88(47)_pad  , \89(48)_pad  , \9(2)_pad  , \94(49)_pad  , \97(50)_pad  , \252(3450)_pad  , \258(3122)_pad  , \270(3109)_pad  , \278(536)_pad  , \281(547)_pad  , \284(384)_pad  , \286(419)_pad  , \292(392)_pad  , \295(3352)_pad  , \298(3387)_pad  , \301(3388)_pad  , \304(3390)_pad  , \307(3389)_pad  , \310(3393)_pad  , \313(3396)_pad  , \316(3397)_pad  , \319(3398)_pad  , \321(3715)_pad  , \324(3363)_pad  , \327(3408)_pad  , \330(3411)_pad  , \333(3416)_pad  , \336(3412)_pad  , \338(3716)_pad  , \344(3382)_pad  , \347(3420)_pad  , \350(3421)_pad  , \353(3425)_pad  , \356(3424)_pad  , \359(3426)_pad  , \362(3429)_pad  , \365(3430)_pad  , \368(3431)_pad  , \370(3718)_pad  , \373(2994)_pad  , \376(3206)_pad  , \379(3207)_pad  , \382(3148)_pad  , \385(3151)_pad  , \388(3093)_pad  , \391(3094)_pad  , \394(3095)_pad  , \397(3097)_pad  , \399(3717)_pad  , \402(395)_pad  , \404(390)_pad  , \406(388)_pad  , \408(385)_pad  , \410(387)_pad  , \412(3369)_pad  , \414(3338)_pad  , \416(3368)_pad  , \418(3449)_pad  , \419(3444)_pad  , \422(3451)_pad  );
  input \100(51)_pad  ;
  input \103(52)_pad  ;
  input \109(54)_pad  ;
  input \110(55)_pad  ;
  input \111(56)_pad  ;
  input \112(57)_pad  ;
  input \113(58)_pad  ;
  input \114(59)_pad  ;
  input \115(60)_pad  ;
  input \118(61)_pad  ;
  input \1197(165)_pad  ;
  input \12(3)_pad  ;
  input \121(62)_pad  ;
  input \124(63)_pad  ;
  input \127(64)_pad  ;
  input \130(65)_pad  ;
  input \133(66)_pad  ;
  input \134(67)_pad  ;
  input \135(68)_pad  ;
  input \138(69)_pad  ;
  input \141(70)_pad  ;
  input \144(71)_pad  ;
  input \1455(166)_pad  ;
  input \147(72)_pad  ;
  input \15(4)_pad  ;
  input \150(73)_pad  ;
  input \151(74)_pad  ;
  input \152(75)_pad  ;
  input \153(76)_pad  ;
  input \154(77)_pad  ;
  input \155(78)_pad  ;
  input \156(79)_pad  ;
  input \157(80)_pad  ;
  input \158(81)_pad  ;
  input \159(82)_pad  ;
  input \160(83)_pad  ;
  input \161(84)_pad  ;
  input \162(85)_pad  ;
  input \163(86)_pad  ;
  input \164(87)_pad  ;
  input \165(88)_pad  ;
  input \166(89)_pad  ;
  input \167(90)_pad  ;
  input \168(91)_pad  ;
  input \169(92)_pad  ;
  input \170(93)_pad  ;
  input \171(94)_pad  ;
  input \172(95)_pad  ;
  input \173(96)_pad  ;
  input \174(97)_pad  ;
  input \175(98)_pad  ;
  input \176(99)_pad  ;
  input \177(100)_pad  ;
  input \178(101)_pad  ;
  input \179(102)_pad  ;
  input \18(5)_pad  ;
  input \180(103)_pad  ;
  input \181(104)_pad  ;
  input \182(105)_pad  ;
  input \183(106)_pad  ;
  input \184(107)_pad  ;
  input \185(108)_pad  ;
  input \186(109)_pad  ;
  input \187(110)_pad  ;
  input \188(111)_pad  ;
  input \189(112)_pad  ;
  input \190(113)_pad  ;
  input \191(114)_pad  ;
  input \192(115)_pad  ;
  input \193(116)_pad  ;
  input \194(117)_pad  ;
  input \195(118)_pad  ;
  input \196(119)_pad  ;
  input \197(120)_pad  ;
  input \198(121)_pad  ;
  input \199(122)_pad  ;
  input \200(123)_pad  ;
  input \201(124)_pad  ;
  input \202(125)_pad  ;
  input \203(126)_pad  ;
  input \204(127)_pad  ;
  input \205(128)_pad  ;
  input \206(129)_pad  ;
  input \207(130)_pad  ;
  input \208(131)_pad  ;
  input \209(132)_pad  ;
  input \210(133)_pad  ;
  input \211(134)_pad  ;
  input \212(135)_pad  ;
  input \213(136)_pad  ;
  input \214(137)_pad  ;
  input \215(138)_pad  ;
  input \216(139)_pad  ;
  input \217(140)_pad  ;
  input \218(141)_pad  ;
  input \219(142)_pad  ;
  input \220(143)_pad  ;
  input \2204(174)_pad  ;
  input \221(144)_pad  ;
  input \222(145)_pad  ;
  input \223(146)_pad  ;
  input \224(147)_pad  ;
  input \225(148)_pad  ;
  input \226(149)_pad  ;
  input \227(150)_pad  ;
  input \228(151)_pad  ;
  input \229(152)_pad  ;
  input \23(6)_pad  ;
  input \230(153)_pad  ;
  input \231(154)_pad  ;
  input \232(155)_pad  ;
  input \233(156)_pad  ;
  input \234(157)_pad  ;
  input \235(158)_pad  ;
  input \236(159)_pad  ;
  input \237(160)_pad  ;
  input \238(161)_pad  ;
  input \239(162)_pad  ;
  input \240(163)_pad  ;
  input \26(7)_pad  ;
  input \29(8)_pad  ;
  input \32(9)_pad  ;
  input \35(10)_pad  ;
  input \38(11)_pad  ;
  input \41(12)_pad  ;
  input \436(286)_pad  ;
  input \438(274)_pad  ;
  input \44(13)_pad  ;
  input \440(277)_pad  ;
  input \442(280)_pad  ;
  input \444(282)_pad  ;
  input \446(393)_pad  ;
  input \448(284)_pad  ;
  input \450(288)_pad  ;
  input \4526(205)_pad  ;
  input \4528(206)_pad  ;
  input \453(596)_pad  ;
  input \47(14)_pad  ;
  input \478(269)_pad  ;
  input \480(250)_pad  ;
  input \482(253)_pad  ;
  input \484(256)_pad  ;
  input \486(258)_pad  ;
  input \488(260)_pad  ;
  input \490(263)_pad  ;
  input \492(265)_pad  ;
  input \494(267)_pad  ;
  input \496(271)_pad  ;
  input \5(1)_pad  ;
  input \50(15)_pad  ;
  input \522(226)_pad  ;
  input \524(210)_pad  ;
  input \526(212)_pad  ;
  input \528(214)_pad  ;
  input \53(16)_pad  ;
  input \530(216)_pad  ;
  input \532(218)_pad  ;
  input \534(220)_pad  ;
  input \536(222)_pad  ;
  input \538(224)_pad  ;
  input \54(17)_pad  ;
  input \540(227)_pad  ;
  input \542(246)_pad  ;
  input \544(230)_pad  ;
  input \546(232)_pad  ;
  input \548(234)_pad  ;
  input \55(18)_pad  ;
  input \550(236)_pad  ;
  input \552(238)_pad  ;
  input \554(240)_pad  ;
  input \556(242)_pad  ;
  input \558(244)_pad  ;
  input \56(19)_pad  ;
  input \560(248)_pad  ;
  input \57(20)_pad  ;
  input \58(21)_pad  ;
  input \59(22)_pad  ;
  input \60(23)_pad  ;
  input \61(24)_pad  ;
  input \62(25)_pad  ;
  input \63(26)_pad  ;
  input \64(27)_pad  ;
  input \65(28)_pad  ;
  input \66(29)_pad  ;
  input \69(30)_pad  ;
  input \70(31)_pad  ;
  input \73(32)_pad  ;
  input \74(33)_pad  ;
  input \75(34)_pad  ;
  input \76(35)_pad  ;
  input \77(36)_pad  ;
  input \78(37)_pad  ;
  input \79(38)_pad  ;
  input \80(39)_pad  ;
  input \81(40)_pad  ;
  input \82(41)_pad  ;
  input \83(42)_pad  ;
  input \84(43)_pad  ;
  input \85(44)_pad  ;
  input \86(45)_pad  ;
  input \87(46)_pad  ;
  input \88(47)_pad  ;
  input \89(48)_pad  ;
  input \9(2)_pad  ;
  input \94(49)_pad  ;
  input \97(50)_pad  ;
  output \252(3450)_pad  ;
  output \258(3122)_pad  ;
  output \270(3109)_pad  ;
  output \278(536)_pad  ;
  output \281(547)_pad  ;
  output \284(384)_pad  ;
  output \286(419)_pad  ;
  output \292(392)_pad  ;
  output \295(3352)_pad  ;
  output \298(3387)_pad  ;
  output \301(3388)_pad  ;
  output \304(3390)_pad  ;
  output \307(3389)_pad  ;
  output \310(3393)_pad  ;
  output \313(3396)_pad  ;
  output \316(3397)_pad  ;
  output \319(3398)_pad  ;
  output \321(3715)_pad  ;
  output \324(3363)_pad  ;
  output \327(3408)_pad  ;
  output \330(3411)_pad  ;
  output \333(3416)_pad  ;
  output \336(3412)_pad  ;
  output \338(3716)_pad  ;
  output \344(3382)_pad  ;
  output \347(3420)_pad  ;
  output \350(3421)_pad  ;
  output \353(3425)_pad  ;
  output \356(3424)_pad  ;
  output \359(3426)_pad  ;
  output \362(3429)_pad  ;
  output \365(3430)_pad  ;
  output \368(3431)_pad  ;
  output \370(3718)_pad  ;
  output \373(2994)_pad  ;
  output \376(3206)_pad  ;
  output \379(3207)_pad  ;
  output \382(3148)_pad  ;
  output \385(3151)_pad  ;
  output \388(3093)_pad  ;
  output \391(3094)_pad  ;
  output \394(3095)_pad  ;
  output \397(3097)_pad  ;
  output \399(3717)_pad  ;
  output \402(395)_pad  ;
  output \404(390)_pad  ;
  output \406(388)_pad  ;
  output \408(385)_pad  ;
  output \410(387)_pad  ;
  output \412(3369)_pad  ;
  output \414(3338)_pad  ;
  output \416(3368)_pad  ;
  output \418(3449)_pad  ;
  output \419(3444)_pad  ;
  output \422(3451)_pad  ;
  wire n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 ;
  assign n207 = ~\18(5)_pad  & \94(49)_pad  ;
  assign n208 = \18(5)_pad  & \195(118)_pad  ;
  assign n209 = ~n207 & ~n208 ;
  assign n210 = ~\18(5)_pad  & \59(22)_pad  ;
  assign n211 = \18(5)_pad  & ~\536(222)_pad  ;
  assign n212 = ~n210 & ~n211 ;
  assign n213 = n209 & n212 ;
  assign n214 = ~\18(5)_pad  & \97(50)_pad  ;
  assign n215 = \18(5)_pad  & \196(119)_pad  ;
  assign n216 = ~n214 & ~n215 ;
  assign n217 = ~\18(5)_pad  & \78(37)_pad  ;
  assign n218 = \18(5)_pad  & ~\538(224)_pad  ;
  assign n219 = ~n217 & ~n218 ;
  assign n220 = n216 & n219 ;
  assign n221 = ~n213 & ~n220 ;
  assign n222 = ~\18(5)_pad  & \47(14)_pad  ;
  assign n223 = \18(5)_pad  & \193(116)_pad  ;
  assign n224 = ~n222 & ~n223 ;
  assign n225 = ~\18(5)_pad  & \80(39)_pad  ;
  assign n226 = \18(5)_pad  & ~\532(218)_pad  ;
  assign n227 = ~n225 & ~n226 ;
  assign n228 = ~n224 & ~n227 ;
  assign n229 = \121(62)_pad  & ~\18(5)_pad  ;
  assign n230 = \18(5)_pad  & \194(117)_pad  ;
  assign n231 = ~n229 & ~n230 ;
  assign n232 = ~\18(5)_pad  & \81(40)_pad  ;
  assign n233 = \18(5)_pad  & ~\534(220)_pad  ;
  assign n234 = ~n232 & ~n233 ;
  assign n235 = ~n231 & ~n234 ;
  assign n236 = ~n209 & ~n212 ;
  assign n237 = ~n235 & ~n236 ;
  assign n238 = ~n228 & n237 ;
  assign n239 = ~n221 & n238 ;
  assign n240 = ~\18(5)_pad  & \23(6)_pad  ;
  assign n241 = \18(5)_pad  & \205(128)_pad  ;
  assign n242 = ~n240 & ~n241 ;
  assign n243 = ~\18(5)_pad  & \75(34)_pad  ;
  assign n244 = \18(5)_pad  & ~\554(240)_pad  ;
  assign n245 = ~n243 & ~n244 ;
  assign n246 = n242 & n245 ;
  assign n247 = \103(52)_pad  & ~\18(5)_pad  ;
  assign n248 = \18(5)_pad  & \204(127)_pad  ;
  assign n249 = ~n247 & ~n248 ;
  assign n250 = ~\18(5)_pad  & \73(32)_pad  ;
  assign n251 = \18(5)_pad  & ~\552(238)_pad  ;
  assign n252 = ~n250 & ~n251 ;
  assign n253 = n249 & n252 ;
  assign n254 = ~n246 & ~n253 ;
  assign n255 = ~n242 & ~n245 ;
  assign n256 = ~\18(5)_pad  & \26(7)_pad  ;
  assign n257 = \18(5)_pad  & \206(129)_pad  ;
  assign n258 = ~n256 & ~n257 ;
  assign n259 = ~\18(5)_pad  & \76(35)_pad  ;
  assign n260 = \18(5)_pad  & ~\556(242)_pad  ;
  assign n261 = ~n259 & ~n260 ;
  assign n262 = ~n258 & ~n261 ;
  assign n263 = ~n255 & ~n262 ;
  assign n264 = n254 & ~n263 ;
  assign n265 = ~\18(5)_pad  & \41(12)_pad  ;
  assign n266 = \70(31)_pad  & n265 ;
  assign n267 = ~\18(5)_pad  & ~\70(31)_pad  ;
  assign n268 = ~\41(12)_pad  & n267 ;
  assign n269 = \89(48)_pad  & ~n268 ;
  assign n270 = ~\18(5)_pad  & \29(8)_pad  ;
  assign n271 = \18(5)_pad  & \207(130)_pad  ;
  assign n272 = ~n270 & ~n271 ;
  assign n273 = ~\18(5)_pad  & \74(33)_pad  ;
  assign n274 = \18(5)_pad  & ~\558(244)_pad  ;
  assign n275 = ~n273 & ~n274 ;
  assign n276 = ~n272 & ~n275 ;
  assign n277 = ~n269 & ~n276 ;
  assign n278 = ~n266 & n277 ;
  assign n279 = n258 & n261 ;
  assign n280 = n272 & n275 ;
  assign n281 = ~n279 & ~n280 ;
  assign n282 = n254 & n281 ;
  assign n283 = ~n278 & n282 ;
  assign n284 = ~n264 & ~n283 ;
  assign n285 = \124(63)_pad  & ~\18(5)_pad  ;
  assign n286 = \18(5)_pad  & \201(124)_pad  ;
  assign n287 = ~n285 & ~n286 ;
  assign n288 = ~\18(5)_pad  & \55(18)_pad  ;
  assign n289 = \18(5)_pad  & ~\546(232)_pad  ;
  assign n290 = ~n288 & ~n289 ;
  assign n291 = n287 & n290 ;
  assign n292 = \127(64)_pad  & ~\18(5)_pad  ;
  assign n293 = \18(5)_pad  & \202(125)_pad  ;
  assign n294 = ~n292 & ~n293 ;
  assign n295 = ~\18(5)_pad  & \54(17)_pad  ;
  assign n296 = \18(5)_pad  & ~\548(234)_pad  ;
  assign n297 = ~n295 & ~n296 ;
  assign n298 = ~n294 & ~n297 ;
  assign n299 = ~n291 & n298 ;
  assign n300 = \100(51)_pad  & ~\18(5)_pad  ;
  assign n301 = \18(5)_pad  & \200(123)_pad  ;
  assign n302 = ~n300 & ~n301 ;
  assign n303 = ~\18(5)_pad  & \56(19)_pad  ;
  assign n304 = \18(5)_pad  & ~\544(230)_pad  ;
  assign n305 = ~n303 & ~n304 ;
  assign n306 = ~n302 & ~n305 ;
  assign n307 = ~n287 & ~n290 ;
  assign n308 = ~n306 & ~n307 ;
  assign n309 = ~n299 & n308 ;
  assign n310 = ~n249 & ~n252 ;
  assign n311 = \130(65)_pad  & ~\18(5)_pad  ;
  assign n312 = \18(5)_pad  & \203(126)_pad  ;
  assign n313 = ~n311 & ~n312 ;
  assign n314 = ~\18(5)_pad  & \53(16)_pad  ;
  assign n315 = \18(5)_pad  & ~\550(236)_pad  ;
  assign n316 = ~n314 & ~n315 ;
  assign n317 = ~n313 & ~n316 ;
  assign n318 = ~n310 & ~n317 ;
  assign n319 = n309 & n318 ;
  assign n320 = n284 & n319 ;
  assign n321 = n294 & n297 ;
  assign n322 = ~n291 & ~n321 ;
  assign n323 = n313 & n316 ;
  assign n324 = ~n298 & ~n323 ;
  assign n325 = n322 & n324 ;
  assign n326 = n309 & ~n325 ;
  assign n327 = \118(61)_pad  & ~\18(5)_pad  ;
  assign n328 = \18(5)_pad  & \187(110)_pad  ;
  assign n329 = ~n327 & ~n328 ;
  assign n330 = ~\18(5)_pad  & \77(36)_pad  ;
  assign n331 = \18(5)_pad  & ~\522(226)_pad  ;
  assign n332 = ~n330 & ~n331 ;
  assign n333 = n329 & n332 ;
  assign n334 = n302 & n305 ;
  assign n335 = ~n333 & ~n334 ;
  assign n336 = ~n326 & n335 ;
  assign n337 = ~n320 & n336 ;
  assign n338 = ~n216 & ~n219 ;
  assign n339 = ~n329 & ~n332 ;
  assign n340 = ~n338 & ~n339 ;
  assign n341 = n238 & n340 ;
  assign n342 = ~n337 & n341 ;
  assign n343 = ~n239 & ~n342 ;
  assign n344 = n231 & n234 ;
  assign n345 = n224 & n227 ;
  assign n346 = ~n344 & ~n345 ;
  assign n347 = ~n228 & ~n346 ;
  assign n348 = ~\18(5)_pad  & \66(29)_pad  ;
  assign n349 = \18(5)_pad  & \189(112)_pad  ;
  assign n350 = ~n348 & ~n349 ;
  assign n351 = ~\18(5)_pad  & \62(25)_pad  ;
  assign n352 = \18(5)_pad  & ~\524(210)_pad  ;
  assign n353 = ~n351 & ~n352 ;
  assign n354 = n350 & n353 ;
  assign n355 = ~\18(5)_pad  & \32(9)_pad  ;
  assign n356 = \18(5)_pad  & \191(114)_pad  ;
  assign n357 = ~n355 & ~n356 ;
  assign n358 = ~\18(5)_pad  & \60(23)_pad  ;
  assign n359 = \18(5)_pad  & ~\528(214)_pad  ;
  assign n360 = ~n358 & ~n359 ;
  assign n361 = n357 & n360 ;
  assign n362 = ~n354 & ~n361 ;
  assign n363 = ~n357 & ~n360 ;
  assign n364 = ~\18(5)_pad  & \50(15)_pad  ;
  assign n365 = \18(5)_pad  & \190(113)_pad  ;
  assign n366 = ~n364 & ~n365 ;
  assign n367 = ~\18(5)_pad  & \61(24)_pad  ;
  assign n368 = \18(5)_pad  & ~\526(212)_pad  ;
  assign n369 = ~n367 & ~n368 ;
  assign n370 = n366 & n369 ;
  assign n371 = ~n363 & ~n370 ;
  assign n372 = n362 & n371 ;
  assign n373 = ~n366 & ~n369 ;
  assign n374 = ~n350 & ~n353 ;
  assign n375 = ~n373 & ~n374 ;
  assign n376 = ~\18(5)_pad  & \35(10)_pad  ;
  assign n377 = \18(5)_pad  & \192(115)_pad  ;
  assign n378 = ~n376 & ~n377 ;
  assign n379 = ~\18(5)_pad  & \79(38)_pad  ;
  assign n380 = \18(5)_pad  & ~\530(216)_pad  ;
  assign n381 = ~n379 & ~n380 ;
  assign n382 = ~n378 & ~n381 ;
  assign n383 = n378 & n381 ;
  assign n384 = ~n382 & ~n383 ;
  assign n385 = n375 & n384 ;
  assign n386 = n372 & n385 ;
  assign n387 = ~n347 & n386 ;
  assign n388 = n343 & n387 ;
  assign n389 = n375 & n382 ;
  assign n390 = n372 & n389 ;
  assign n391 = n363 & ~n370 ;
  assign n392 = n375 & ~n391 ;
  assign n393 = ~n354 & ~n392 ;
  assign n394 = ~n390 & ~n393 ;
  assign n395 = ~n388 & n394 ;
  assign n396 = \12(3)_pad  & \9(2)_pad  ;
  assign n397 = ~\167(90)_pad  & \18(5)_pad  ;
  assign n398 = ~n396 & ~n397 ;
  assign n399 = \18(5)_pad  & ~\444(282)_pad  ;
  assign n400 = \112(57)_pad  & ~\18(5)_pad  ;
  assign n401 = ~n399 & ~n400 ;
  assign n402 = n398 & ~n401 ;
  assign n403 = ~\168(91)_pad  & \18(5)_pad  ;
  assign n404 = ~n396 & ~n403 ;
  assign n405 = \18(5)_pad  & ~\446(393)_pad  ;
  assign n406 = ~\18(5)_pad  & \87(46)_pad  ;
  assign n407 = ~n405 & ~n406 ;
  assign n408 = n404 & ~n407 ;
  assign n409 = ~n402 & ~n408 ;
  assign n410 = ~n398 & n401 ;
  assign n411 = ~n404 & n407 ;
  assign n412 = ~n410 & ~n411 ;
  assign n413 = n409 & n412 ;
  assign n414 = ~\169(92)_pad  & \18(5)_pad  ;
  assign n415 = ~n396 & ~n414 ;
  assign n416 = \18(5)_pad  & ~\448(284)_pad  ;
  assign n417 = \111(56)_pad  & ~\18(5)_pad  ;
  assign n418 = ~n416 & ~n417 ;
  assign n419 = ~n415 & n418 ;
  assign n420 = n415 & ~n418 ;
  assign n421 = ~n419 & ~n420 ;
  assign n422 = n413 & n421 ;
  assign n423 = \1455(166)_pad  & \2204(174)_pad  ;
  assign n424 = ~\38(11)_pad  & \4528(206)_pad  ;
  assign n425 = ~n423 & n424 ;
  assign n426 = ~\166(89)_pad  & \18(5)_pad  ;
  assign n427 = ~n396 & ~n426 ;
  assign n428 = \18(5)_pad  & ~\442(280)_pad  ;
  assign n429 = ~\18(5)_pad  & \88(47)_pad  ;
  assign n430 = ~n428 & ~n429 ;
  assign n431 = ~n427 & n430 ;
  assign n432 = ~\1455(166)_pad  & ~\2204(174)_pad  ;
  assign n433 = \4528(206)_pad  & n432 ;
  assign n434 = \38(11)_pad  & ~n433 ;
  assign n435 = ~n431 & ~n434 ;
  assign n436 = ~n425 & n435 ;
  assign n437 = n427 & ~n430 ;
  assign n438 = \18(5)_pad  & ~\436(286)_pad  ;
  assign n439 = \113(58)_pad  & ~\18(5)_pad  ;
  assign n440 = ~n438 & ~n439 ;
  assign n441 = ~n396 & ~n440 ;
  assign n442 = n396 & n440 ;
  assign n443 = ~n441 & ~n442 ;
  assign n444 = ~n437 & n443 ;
  assign n445 = n436 & n444 ;
  assign n446 = n422 & n445 ;
  assign n447 = n431 & ~n434 ;
  assign n448 = n425 & ~n434 ;
  assign n449 = ~n447 & ~n448 ;
  assign n450 = n413 & n420 ;
  assign n451 = ~n409 & ~n410 ;
  assign n452 = ~n437 & ~n451 ;
  assign n453 = ~n450 & n452 ;
  assign n454 = n421 & n441 ;
  assign n455 = n413 & n454 ;
  assign n456 = ~n434 & ~n455 ;
  assign n457 = n453 & n456 ;
  assign n458 = n449 & ~n457 ;
  assign n459 = ~n446 & ~n458 ;
  assign n460 = ~\177(100)_pad  & \18(5)_pad  ;
  assign n461 = ~n396 & ~n460 ;
  assign n462 = \18(5)_pad  & ~\488(260)_pad  ;
  assign n463 = ~\18(5)_pad  & \64(27)_pad  ;
  assign n464 = ~n462 & ~n463 ;
  assign n465 = n461 & ~n464 ;
  assign n466 = \178(101)_pad  & \18(5)_pad  ;
  assign n467 = \135(68)_pad  & ~\18(5)_pad  ;
  assign n468 = ~n466 & ~n467 ;
  assign n469 = \18(5)_pad  & ~\490(263)_pad  ;
  assign n470 = ~\18(5)_pad  & \85(44)_pad  ;
  assign n471 = ~n469 & ~n470 ;
  assign n472 = ~n468 & ~n471 ;
  assign n473 = ~n465 & ~n472 ;
  assign n474 = ~\175(98)_pad  & \18(5)_pad  ;
  assign n475 = ~n396 & ~n474 ;
  assign n476 = \18(5)_pad  & ~\484(256)_pad  ;
  assign n477 = ~\18(5)_pad  & \86(45)_pad  ;
  assign n478 = ~n476 & ~n477 ;
  assign n479 = ~n475 & n478 ;
  assign n480 = ~\176(99)_pad  & \18(5)_pad  ;
  assign n481 = ~n396 & ~n480 ;
  assign n482 = \18(5)_pad  & ~\486(258)_pad  ;
  assign n483 = ~\18(5)_pad  & \63(26)_pad  ;
  assign n484 = ~n482 & ~n483 ;
  assign n485 = n481 & ~n484 ;
  assign n486 = ~n479 & ~n485 ;
  assign n487 = \179(102)_pad  & \18(5)_pad  ;
  assign n488 = \144(71)_pad  & ~\18(5)_pad  ;
  assign n489 = ~n487 & ~n488 ;
  assign n490 = \18(5)_pad  & ~\492(265)_pad  ;
  assign n491 = ~\18(5)_pad  & \84(43)_pad  ;
  assign n492 = ~n490 & ~n491 ;
  assign n493 = n489 & n492 ;
  assign n494 = n468 & n471 ;
  assign n495 = ~n493 & ~n494 ;
  assign n496 = n486 & n495 ;
  assign n497 = n473 & n496 ;
  assign n498 = ~\174(97)_pad  & \18(5)_pad  ;
  assign n499 = ~n396 & ~n498 ;
  assign n500 = \18(5)_pad  & ~\482(253)_pad  ;
  assign n501 = \109(54)_pad  & ~\18(5)_pad  ;
  assign n502 = ~n500 & ~n501 ;
  assign n503 = ~n499 & n502 ;
  assign n504 = ~\173(96)_pad  & \18(5)_pad  ;
  assign n505 = ~n396 & ~n504 ;
  assign n506 = \18(5)_pad  & ~\480(250)_pad  ;
  assign n507 = \110(55)_pad  & ~\18(5)_pad  ;
  assign n508 = ~n506 & ~n507 ;
  assign n509 = ~n505 & n508 ;
  assign n510 = ~n503 & ~n509 ;
  assign n511 = n505 & ~n508 ;
  assign n512 = \18(5)_pad  & \180(103)_pad  ;
  assign n513 = \138(69)_pad  & ~\18(5)_pad  ;
  assign n514 = ~n512 & ~n513 ;
  assign n515 = \18(5)_pad  & ~\494(267)_pad  ;
  assign n516 = ~\18(5)_pad  & \83(42)_pad  ;
  assign n517 = ~n515 & ~n516 ;
  assign n518 = n514 & n517 ;
  assign n519 = \171(94)_pad  & \18(5)_pad  ;
  assign n520 = \147(72)_pad  & ~\18(5)_pad  ;
  assign n521 = ~n519 & ~n520 ;
  assign n522 = \18(5)_pad  & ~\478(269)_pad  ;
  assign n523 = ~\18(5)_pad  & \65(28)_pad  ;
  assign n524 = ~n522 & ~n523 ;
  assign n525 = n521 & n524 ;
  assign n526 = ~n518 & ~n525 ;
  assign n527 = ~n511 & n526 ;
  assign n528 = n510 & n527 ;
  assign n529 = n497 & n528 ;
  assign n530 = ~n514 & ~n517 ;
  assign n531 = ~n489 & ~n492 ;
  assign n532 = ~n521 & ~n524 ;
  assign n533 = ~n531 & ~n532 ;
  assign n534 = ~n530 & n533 ;
  assign n535 = n499 & ~n502 ;
  assign n536 = n475 & ~n478 ;
  assign n537 = ~n535 & ~n536 ;
  assign n538 = ~n461 & n464 ;
  assign n539 = ~n481 & n484 ;
  assign n540 = ~n538 & ~n539 ;
  assign n541 = n537 & n540 ;
  assign n542 = n534 & n541 ;
  assign n543 = n386 & n542 ;
  assign n544 = n529 & n543 ;
  assign n545 = ~n347 & n544 ;
  assign n546 = n343 & n545 ;
  assign n547 = n529 & n542 ;
  assign n548 = ~n394 & n547 ;
  assign n549 = ~n510 & ~n511 ;
  assign n550 = n518 & ~n531 ;
  assign n551 = n495 & ~n550 ;
  assign n552 = ~n534 & n551 ;
  assign n553 = n473 & ~n485 ;
  assign n554 = ~n552 & n553 ;
  assign n555 = ~n485 & ~n540 ;
  assign n556 = ~n479 & ~n555 ;
  assign n557 = ~n554 & n556 ;
  assign n558 = ~n511 & n537 ;
  assign n559 = ~n557 & n558 ;
  assign n560 = ~n549 & ~n559 ;
  assign n561 = ~n458 & ~n560 ;
  assign n562 = ~n548 & n561 ;
  assign n563 = ~n546 & n562 ;
  assign n564 = ~n459 & ~n563 ;
  assign n565 = ~\155(78)_pad  & \18(5)_pad  ;
  assign n566 = ~n396 & ~n565 ;
  assign n567 = ~\484(256)_pad  & n566 ;
  assign n568 = \484(256)_pad  & ~n566 ;
  assign n569 = ~n567 & ~n568 ;
  assign n570 = ~\156(79)_pad  & \18(5)_pad  ;
  assign n571 = ~n396 & ~n570 ;
  assign n572 = ~\486(258)_pad  & n571 ;
  assign n573 = \486(258)_pad  & ~n571 ;
  assign n574 = ~n572 & ~n573 ;
  assign n575 = n569 & n574 ;
  assign n576 = \151(74)_pad  & \18(5)_pad  ;
  assign n577 = ~n520 & ~n576 ;
  assign n578 = ~\478(269)_pad  & ~n577 ;
  assign n579 = \478(269)_pad  & n577 ;
  assign n580 = ~n578 & ~n579 ;
  assign n581 = \159(82)_pad  & \18(5)_pad  ;
  assign n582 = ~n488 & ~n581 ;
  assign n583 = ~\492(265)_pad  & ~n582 ;
  assign n584 = \492(265)_pad  & n582 ;
  assign n585 = ~n583 & ~n584 ;
  assign n586 = \160(83)_pad  & \18(5)_pad  ;
  assign n587 = ~n513 & ~n586 ;
  assign n588 = ~\494(267)_pad  & ~n587 ;
  assign n589 = \494(267)_pad  & n587 ;
  assign n590 = ~n588 & ~n589 ;
  assign n591 = n585 & n590 ;
  assign n592 = n580 & n591 ;
  assign n593 = \158(81)_pad  & \18(5)_pad  ;
  assign n594 = ~n467 & ~n593 ;
  assign n595 = ~\490(263)_pad  & ~n594 ;
  assign n596 = \490(263)_pad  & n594 ;
  assign n597 = ~n595 & ~n596 ;
  assign n598 = ~\157(80)_pad  & \18(5)_pad  ;
  assign n599 = ~n396 & ~n598 ;
  assign n600 = ~\488(260)_pad  & n599 ;
  assign n601 = \488(260)_pad  & ~n599 ;
  assign n602 = ~n600 & ~n601 ;
  assign n603 = n597 & n602 ;
  assign n604 = ~\154(77)_pad  & \18(5)_pad  ;
  assign n605 = ~n396 & ~n604 ;
  assign n606 = ~\482(253)_pad  & n605 ;
  assign n607 = \482(253)_pad  & ~n605 ;
  assign n608 = ~n606 & ~n607 ;
  assign n609 = ~\153(76)_pad  & \18(5)_pad  ;
  assign n610 = ~n396 & ~n609 ;
  assign n611 = ~\480(250)_pad  & n610 ;
  assign n612 = \480(250)_pad  & ~n610 ;
  assign n613 = ~n611 & ~n612 ;
  assign n614 = n608 & n613 ;
  assign n615 = n603 & n614 ;
  assign n616 = n592 & n615 ;
  assign n617 = n575 & n616 ;
  assign n618 = n578 & ~n589 ;
  assign n619 = ~n583 & ~n588 ;
  assign n620 = ~n618 & n619 ;
  assign n621 = ~n596 & ~n601 ;
  assign n622 = ~n584 & n621 ;
  assign n623 = ~n620 & n622 ;
  assign n624 = n595 & ~n601 ;
  assign n625 = ~n600 & ~n624 ;
  assign n626 = ~n623 & n625 ;
  assign n627 = n608 & ~n612 ;
  assign n628 = n575 & n627 ;
  assign n629 = ~n626 & n628 ;
  assign n630 = \18(5)_pad  & ~\216(139)_pad  ;
  assign n631 = ~n396 & ~n630 ;
  assign n632 = ~\448(284)_pad  & n631 ;
  assign n633 = \18(5)_pad  & ~\209(132)_pad  ;
  assign n634 = ~n396 & ~n633 ;
  assign n635 = ~\436(286)_pad  & n634 ;
  assign n636 = ~n632 & ~n635 ;
  assign n637 = \18(5)_pad  & ~\215(138)_pad  ;
  assign n638 = ~n396 & ~n637 ;
  assign n639 = \446(393)_pad  & ~n638 ;
  assign n640 = \448(284)_pad  & ~n631 ;
  assign n641 = ~n639 & ~n640 ;
  assign n642 = ~n636 & n641 ;
  assign n643 = ~\446(393)_pad  & n638 ;
  assign n644 = \18(5)_pad  & ~\214(137)_pad  ;
  assign n645 = ~n396 & ~n644 ;
  assign n646 = ~\444(282)_pad  & n645 ;
  assign n647 = ~n643 & ~n646 ;
  assign n648 = ~n642 & n647 ;
  assign n649 = ~n567 & ~n572 ;
  assign n650 = ~n568 & ~n607 ;
  assign n651 = ~n649 & n650 ;
  assign n652 = ~n606 & ~n611 ;
  assign n653 = ~n651 & n652 ;
  assign n654 = ~n612 & ~n653 ;
  assign n655 = n648 & ~n654 ;
  assign n656 = ~n629 & n655 ;
  assign n657 = ~n617 & n656 ;
  assign n658 = \18(5)_pad  & \231(154)_pad  ;
  assign n659 = ~n300 & ~n658 ;
  assign n660 = \544(230)_pad  & n659 ;
  assign n661 = \18(5)_pad  & \233(156)_pad  ;
  assign n662 = ~n292 & ~n661 ;
  assign n663 = ~\548(234)_pad  & ~n662 ;
  assign n664 = \18(5)_pad  & \234(157)_pad  ;
  assign n665 = ~n311 & ~n664 ;
  assign n666 = ~\550(236)_pad  & ~n665 ;
  assign n667 = ~n663 & ~n666 ;
  assign n668 = \18(5)_pad  & \232(155)_pad  ;
  assign n669 = ~n285 & ~n668 ;
  assign n670 = \546(232)_pad  & n669 ;
  assign n671 = \548(234)_pad  & n662 ;
  assign n672 = ~n670 & ~n671 ;
  assign n673 = ~n667 & n672 ;
  assign n674 = ~\546(232)_pad  & ~n669 ;
  assign n675 = ~\544(230)_pad  & ~n659 ;
  assign n676 = ~n674 & ~n675 ;
  assign n677 = ~n673 & n676 ;
  assign n678 = ~n660 & ~n677 ;
  assign n679 = \18(5)_pad  & \220(143)_pad  ;
  assign n680 = ~n364 & ~n679 ;
  assign n681 = ~\526(212)_pad  & ~n680 ;
  assign n682 = \526(212)_pad  & n680 ;
  assign n683 = ~n681 & ~n682 ;
  assign n684 = \18(5)_pad  & \221(144)_pad  ;
  assign n685 = ~n355 & ~n684 ;
  assign n686 = ~\528(214)_pad  & ~n685 ;
  assign n687 = \528(214)_pad  & n685 ;
  assign n688 = ~n686 & ~n687 ;
  assign n689 = \18(5)_pad  & \222(145)_pad  ;
  assign n690 = ~n376 & ~n689 ;
  assign n691 = ~\530(216)_pad  & ~n690 ;
  assign n692 = \530(216)_pad  & n690 ;
  assign n693 = ~n691 & ~n692 ;
  assign n694 = n688 & n693 ;
  assign n695 = n683 & n694 ;
  assign n696 = \18(5)_pad  & \217(140)_pad  ;
  assign n697 = ~n327 & ~n696 ;
  assign n698 = ~\522(226)_pad  & ~n697 ;
  assign n699 = \522(226)_pad  & n697 ;
  assign n700 = ~n698 & ~n699 ;
  assign n701 = \18(5)_pad  & \226(149)_pad  ;
  assign n702 = ~n214 & ~n701 ;
  assign n703 = \538(224)_pad  & n702 ;
  assign n704 = ~\538(224)_pad  & ~n702 ;
  assign n705 = ~n703 & ~n704 ;
  assign n706 = \18(5)_pad  & \225(148)_pad  ;
  assign n707 = ~n207 & ~n706 ;
  assign n708 = ~\536(222)_pad  & ~n707 ;
  assign n709 = \536(222)_pad  & n707 ;
  assign n710 = ~n708 & ~n709 ;
  assign n711 = n705 & n710 ;
  assign n712 = n700 & n711 ;
  assign n713 = \18(5)_pad  & \224(147)_pad  ;
  assign n714 = ~n229 & ~n713 ;
  assign n715 = \534(220)_pad  & n714 ;
  assign n716 = ~\534(220)_pad  & ~n714 ;
  assign n717 = ~n715 & ~n716 ;
  assign n718 = \18(5)_pad  & \223(146)_pad  ;
  assign n719 = ~n222 & ~n718 ;
  assign n720 = ~\532(218)_pad  & ~n719 ;
  assign n721 = \532(218)_pad  & n719 ;
  assign n722 = ~n720 & ~n721 ;
  assign n723 = n717 & n722 ;
  assign n724 = \18(5)_pad  & \219(142)_pad  ;
  assign n725 = ~n348 & ~n724 ;
  assign n726 = \524(210)_pad  & n725 ;
  assign n727 = ~\524(210)_pad  & ~n725 ;
  assign n728 = ~n726 & ~n727 ;
  assign n729 = n723 & n728 ;
  assign n730 = n712 & n729 ;
  assign n731 = n695 & n730 ;
  assign n732 = n678 & n731 ;
  assign n733 = \18(5)_pad  & \236(159)_pad  ;
  assign n734 = ~n240 & ~n733 ;
  assign n735 = ~\554(240)_pad  & ~n734 ;
  assign n736 = \554(240)_pad  & n734 ;
  assign n737 = \18(5)_pad  & \235(158)_pad  ;
  assign n738 = ~n247 & ~n737 ;
  assign n739 = \552(238)_pad  & n738 ;
  assign n740 = ~n736 & ~n739 ;
  assign n741 = n735 & n740 ;
  assign n742 = \18(5)_pad  & \238(161)_pad  ;
  assign n743 = ~n270 & ~n742 ;
  assign n744 = \558(244)_pad  & n743 ;
  assign n745 = ~\542(246)_pad  & n265 ;
  assign n746 = ~n744 & n745 ;
  assign n747 = \18(5)_pad  & \237(160)_pad  ;
  assign n748 = ~n256 & ~n747 ;
  assign n749 = ~\556(242)_pad  & ~n748 ;
  assign n750 = ~\558(244)_pad  & ~n743 ;
  assign n751 = ~n749 & ~n750 ;
  assign n752 = ~n746 & n751 ;
  assign n753 = \556(242)_pad  & n748 ;
  assign n754 = n740 & ~n753 ;
  assign n755 = ~n752 & n754 ;
  assign n756 = ~n741 & ~n755 ;
  assign n757 = ~\552(238)_pad  & ~n738 ;
  assign n758 = ~n749 & ~n753 ;
  assign n759 = ~\18(5)_pad  & \542(246)_pad  ;
  assign n760 = n265 & ~n759 ;
  assign n761 = ~n265 & n759 ;
  assign n762 = ~n760 & ~n761 ;
  assign n763 = ~n744 & ~n750 ;
  assign n764 = n762 & n763 ;
  assign n765 = \4526(205)_pad  & ~n735 ;
  assign n766 = n740 & n765 ;
  assign n767 = n764 & n766 ;
  assign n768 = n758 & n767 ;
  assign n769 = ~n757 & ~n768 ;
  assign n770 = n756 & n769 ;
  assign n771 = ~n663 & ~n671 ;
  assign n772 = \550(236)_pad  & n665 ;
  assign n773 = ~n666 & ~n772 ;
  assign n774 = n771 & n773 ;
  assign n775 = ~n670 & ~n674 ;
  assign n776 = ~n660 & ~n675 ;
  assign n777 = n775 & n776 ;
  assign n778 = n774 & n777 ;
  assign n779 = n695 & n778 ;
  assign n780 = n730 & n779 ;
  assign n781 = ~n770 & n780 ;
  assign n782 = ~n732 & ~n781 ;
  assign n783 = ~n681 & ~n727 ;
  assign n784 = n683 & ~n721 ;
  assign n785 = n694 & n784 ;
  assign n786 = ~n686 & ~n691 ;
  assign n787 = ~n682 & ~n687 ;
  assign n788 = ~n786 & n787 ;
  assign n789 = ~n785 & ~n788 ;
  assign n790 = n698 & ~n703 ;
  assign n791 = ~n704 & ~n708 ;
  assign n792 = ~n790 & n791 ;
  assign n793 = ~n709 & ~n715 ;
  assign n794 = ~n792 & n793 ;
  assign n795 = ~n716 & ~n720 ;
  assign n796 = ~n788 & n795 ;
  assign n797 = ~n794 & n796 ;
  assign n798 = ~n789 & ~n797 ;
  assign n799 = n783 & ~n798 ;
  assign n800 = ~n726 & ~n799 ;
  assign n801 = n656 & ~n800 ;
  assign n802 = n782 & n801 ;
  assign n803 = ~n657 & ~n802 ;
  assign n804 = ~n639 & ~n643 ;
  assign n805 = ~n632 & ~n640 ;
  assign n806 = n804 & n805 ;
  assign n807 = \436(286)_pad  & ~n634 ;
  assign n808 = ~n635 & ~n807 ;
  assign n809 = n806 & n808 ;
  assign n810 = n648 & ~n809 ;
  assign n811 = \18(5)_pad  & ~\213(136)_pad  ;
  assign n812 = ~n396 & ~n811 ;
  assign n813 = ~\442(280)_pad  & n812 ;
  assign n814 = \442(280)_pad  & ~n812 ;
  assign n815 = ~n813 & ~n814 ;
  assign n816 = \444(282)_pad  & ~n645 ;
  assign n817 = n815 & ~n816 ;
  assign n818 = ~n810 & n817 ;
  assign n819 = n803 & n818 ;
  assign n820 = \440(277)_pad  & \4528(206)_pad  ;
  assign n821 = \438(274)_pad  & n820 ;
  assign n822 = \38(11)_pad  & ~n821 ;
  assign n823 = ~n813 & ~n822 ;
  assign n824 = ~n819 & n823 ;
  assign n825 = \438(274)_pad  & \4528(206)_pad  ;
  assign n826 = ~n820 & ~n825 ;
  assign n827 = ~\38(11)_pad  & ~n826 ;
  assign n828 = ~n824 & ~n827 ;
  assign n829 = \163(86)_pad  & \453(596)_pad  ;
  assign n830 = \133(66)_pad  & \134(67)_pad  ;
  assign n831 = ~\5(1)_pad  & n830 ;
  assign n832 = \1197(165)_pad  & ~\5(1)_pad  ;
  assign n833 = n782 & ~n800 ;
  assign n834 = ~n580 & ~n833 ;
  assign n835 = n580 & ~n800 ;
  assign n836 = n782 & n835 ;
  assign n837 = ~n834 & ~n836 ;
  assign n838 = n575 & n608 ;
  assign n839 = n592 & n603 ;
  assign n840 = n626 & ~n839 ;
  assign n841 = n626 & ~n800 ;
  assign n842 = n782 & n841 ;
  assign n843 = ~n840 & ~n842 ;
  assign n844 = n838 & n843 ;
  assign n845 = ~n606 & ~n651 ;
  assign n846 = ~n613 & n845 ;
  assign n847 = ~n844 & n846 ;
  assign n848 = n575 & n614 ;
  assign n849 = n843 & n848 ;
  assign n850 = n613 & ~n845 ;
  assign n851 = ~n849 & ~n850 ;
  assign n852 = ~n847 & n851 ;
  assign n853 = ~n568 & ~n649 ;
  assign n854 = ~n843 & ~n853 ;
  assign n855 = ~n567 & n573 ;
  assign n856 = ~n568 & ~n855 ;
  assign n857 = ~n608 & n856 ;
  assign n858 = ~n854 & n857 ;
  assign n859 = n608 & ~n856 ;
  assign n860 = n608 & ~n853 ;
  assign n861 = ~n843 & n860 ;
  assign n862 = ~n859 & ~n861 ;
  assign n863 = ~n858 & n862 ;
  assign n864 = n574 & ~n843 ;
  assign n865 = ~n569 & ~n573 ;
  assign n866 = n569 & n573 ;
  assign n867 = ~n865 & ~n866 ;
  assign n868 = ~n864 & ~n867 ;
  assign n869 = n575 & ~n843 ;
  assign n870 = ~n868 & ~n869 ;
  assign n871 = ~n574 & n843 ;
  assign n872 = ~n864 & ~n871 ;
  assign n873 = ~n578 & ~n800 ;
  assign n874 = n782 & n873 ;
  assign n875 = n585 & ~n589 ;
  assign n876 = ~n579 & n875 ;
  assign n877 = ~n874 & n876 ;
  assign n878 = n585 & n588 ;
  assign n879 = ~n583 & ~n595 ;
  assign n880 = ~n878 & n879 ;
  assign n881 = ~n877 & n880 ;
  assign n882 = ~n596 & n602 ;
  assign n883 = ~n881 & n882 ;
  assign n884 = ~n596 & ~n881 ;
  assign n885 = ~n602 & ~n884 ;
  assign n886 = ~n883 & ~n885 ;
  assign n887 = ~n583 & ~n878 ;
  assign n888 = ~n877 & n887 ;
  assign n889 = ~n597 & ~n888 ;
  assign n890 = ~n583 & n597 ;
  assign n891 = ~n878 & n890 ;
  assign n892 = ~n877 & n891 ;
  assign n893 = ~n889 & ~n892 ;
  assign n894 = ~n877 & ~n878 ;
  assign n895 = ~n579 & ~n589 ;
  assign n896 = ~n874 & n895 ;
  assign n897 = ~n585 & ~n588 ;
  assign n898 = ~n896 & n897 ;
  assign n899 = n894 & ~n898 ;
  assign n900 = ~n579 & ~n874 ;
  assign n901 = ~n590 & ~n900 ;
  assign n902 = ~n579 & n590 ;
  assign n903 = ~n874 & n902 ;
  assign n904 = ~n901 & ~n903 ;
  assign n905 = ~n585 & ~n590 ;
  assign n906 = ~n591 & ~n905 ;
  assign n907 = ~n578 & ~n588 ;
  assign n908 = ~n618 & ~n907 ;
  assign n909 = ~n584 & ~n596 ;
  assign n910 = ~n620 & n909 ;
  assign n911 = n908 & n910 ;
  assign n912 = ~n584 & ~n620 ;
  assign n913 = ~n595 & n908 ;
  assign n914 = ~n912 & n913 ;
  assign n915 = ~n911 & ~n914 ;
  assign n916 = ~n595 & ~n912 ;
  assign n917 = ~n908 & ~n910 ;
  assign n918 = ~n916 & n917 ;
  assign n919 = n915 & ~n918 ;
  assign n920 = ~n580 & ~n919 ;
  assign n921 = n580 & n919 ;
  assign n922 = ~n920 & ~n921 ;
  assign n923 = n833 & ~n922 ;
  assign n924 = ~n592 & n916 ;
  assign n925 = n580 & ~n596 ;
  assign n926 = n591 & n925 ;
  assign n927 = ~n910 & ~n926 ;
  assign n928 = n579 & ~n588 ;
  assign n929 = ~n895 & ~n928 ;
  assign n930 = n927 & ~n929 ;
  assign n931 = ~n924 & n930 ;
  assign n932 = ~n927 & n929 ;
  assign n933 = ~n592 & n929 ;
  assign n934 = n916 & n933 ;
  assign n935 = ~n932 & ~n934 ;
  assign n936 = ~n931 & n935 ;
  assign n937 = n580 & n936 ;
  assign n938 = ~n920 & ~n937 ;
  assign n939 = ~n833 & n938 ;
  assign n940 = ~n923 & ~n939 ;
  assign n941 = n906 & ~n940 ;
  assign n942 = ~n906 & n940 ;
  assign n943 = ~n941 & ~n942 ;
  assign n944 = ~n597 & ~n602 ;
  assign n945 = ~n603 & ~n944 ;
  assign n946 = ~n608 & ~n613 ;
  assign n947 = ~n614 & ~n946 ;
  assign n948 = n945 & n947 ;
  assign n949 = ~n945 & ~n947 ;
  assign n950 = ~n948 & ~n949 ;
  assign n951 = ~n838 & n856 ;
  assign n952 = n845 & n951 ;
  assign n953 = n569 & n572 ;
  assign n954 = ~n569 & ~n572 ;
  assign n955 = ~n953 & ~n954 ;
  assign n956 = \486(258)_pad  & ~n566 ;
  assign n957 = ~n571 & n956 ;
  assign n958 = \484(256)_pad  & \486(258)_pad  ;
  assign n959 = ~n571 & n958 ;
  assign n960 = ~n568 & ~n959 ;
  assign n961 = ~n957 & n960 ;
  assign n962 = n606 & ~n961 ;
  assign n963 = ~n955 & ~n962 ;
  assign n964 = ~n952 & n963 ;
  assign n965 = n955 & n962 ;
  assign n966 = n845 & n955 ;
  assign n967 = n951 & n966 ;
  assign n968 = ~n965 & ~n967 ;
  assign n969 = ~n964 & n968 ;
  assign n970 = n843 & n969 ;
  assign n971 = ~n606 & ~n853 ;
  assign n972 = ~n651 & ~n971 ;
  assign n973 = ~n867 & n972 ;
  assign n974 = n867 & ~n972 ;
  assign n975 = ~n973 & ~n974 ;
  assign n976 = ~n843 & ~n975 ;
  assign n977 = ~n970 & ~n976 ;
  assign n978 = n950 & ~n977 ;
  assign n979 = ~n943 & n978 ;
  assign n980 = n950 & n977 ;
  assign n981 = n943 & n980 ;
  assign n982 = ~n979 & ~n981 ;
  assign n983 = ~n950 & n977 ;
  assign n984 = ~n943 & n983 ;
  assign n985 = ~n950 & ~n977 ;
  assign n986 = n943 & n985 ;
  assign n987 = ~n984 & ~n986 ;
  assign n988 = n982 & n987 ;
  assign n989 = ~n629 & ~n654 ;
  assign n990 = ~n617 & n989 ;
  assign n991 = ~n800 & n989 ;
  assign n992 = n782 & n991 ;
  assign n993 = ~n990 & ~n992 ;
  assign n994 = ~n808 & n993 ;
  assign n995 = n808 & ~n993 ;
  assign n996 = ~n994 & ~n995 ;
  assign n997 = ~n810 & ~n816 ;
  assign n998 = n803 & n997 ;
  assign n999 = ~n815 & ~n998 ;
  assign n1000 = ~n819 & ~n999 ;
  assign n1001 = ~n646 & ~n816 ;
  assign n1002 = ~n642 & ~n643 ;
  assign n1003 = ~n809 & n1002 ;
  assign n1004 = ~n1001 & n1003 ;
  assign n1005 = ~n1001 & n1002 ;
  assign n1006 = ~n993 & n1005 ;
  assign n1007 = ~n1004 & ~n1006 ;
  assign n1008 = ~n993 & n1002 ;
  assign n1009 = n1001 & ~n1003 ;
  assign n1010 = ~n1008 & n1009 ;
  assign n1011 = n1007 & ~n1010 ;
  assign n1012 = ~n635 & ~n993 ;
  assign n1013 = ~n640 & ~n807 ;
  assign n1014 = ~n1012 & n1013 ;
  assign n1015 = ~n632 & ~n804 ;
  assign n1016 = ~n1014 & n1015 ;
  assign n1017 = n632 & n804 ;
  assign n1018 = n804 & n1013 ;
  assign n1019 = ~n1012 & n1018 ;
  assign n1020 = ~n1017 & ~n1019 ;
  assign n1021 = ~n1016 & n1020 ;
  assign n1022 = ~n805 & ~n807 ;
  assign n1023 = ~n1012 & n1022 ;
  assign n1024 = n805 & n807 ;
  assign n1025 = ~n635 & n805 ;
  assign n1026 = ~n993 & n1025 ;
  assign n1027 = ~n1024 & ~n1026 ;
  assign n1028 = ~n1023 & n1027 ;
  assign n1029 = ~n804 & ~n805 ;
  assign n1030 = ~n806 & ~n1029 ;
  assign n1031 = n815 & n1030 ;
  assign n1032 = ~n815 & ~n1030 ;
  assign n1033 = ~n1031 & ~n1032 ;
  assign n1034 = n635 & ~n640 ;
  assign n1035 = ~n636 & ~n1034 ;
  assign n1036 = n648 & n1035 ;
  assign n1037 = ~n816 & n1035 ;
  assign n1038 = ~n1002 & n1037 ;
  assign n1039 = ~n1036 & ~n1038 ;
  assign n1040 = ~n816 & ~n1002 ;
  assign n1041 = ~n648 & ~n1035 ;
  assign n1042 = ~n1040 & n1041 ;
  assign n1043 = n1039 & ~n1042 ;
  assign n1044 = ~n808 & ~n1001 ;
  assign n1045 = ~n1043 & n1044 ;
  assign n1046 = n808 & ~n1001 ;
  assign n1047 = n1043 & n1046 ;
  assign n1048 = ~n1045 & ~n1047 ;
  assign n1049 = n808 & n1001 ;
  assign n1050 = ~n1043 & n1049 ;
  assign n1051 = ~n808 & n1001 ;
  assign n1052 = n1043 & n1051 ;
  assign n1053 = ~n1050 & ~n1052 ;
  assign n1054 = n1048 & n1053 ;
  assign n1055 = ~n993 & ~n1054 ;
  assign n1056 = ~n1033 & n1055 ;
  assign n1057 = ~n808 & ~n1043 ;
  assign n1058 = ~n816 & ~n1003 ;
  assign n1059 = ~n810 & ~n1058 ;
  assign n1060 = ~n632 & n807 ;
  assign n1061 = ~n1013 & ~n1060 ;
  assign n1062 = ~n1059 & n1061 ;
  assign n1063 = ~n810 & ~n1061 ;
  assign n1064 = ~n1058 & n1063 ;
  assign n1065 = n808 & ~n1064 ;
  assign n1066 = ~n1062 & n1065 ;
  assign n1067 = ~n1057 & ~n1066 ;
  assign n1068 = ~n1001 & ~n1067 ;
  assign n1069 = n1001 & ~n1057 ;
  assign n1070 = ~n1066 & n1069 ;
  assign n1071 = ~n1068 & ~n1070 ;
  assign n1072 = n993 & ~n1033 ;
  assign n1073 = n1071 & n1072 ;
  assign n1074 = ~n1056 & ~n1073 ;
  assign n1075 = n993 & n1071 ;
  assign n1076 = n1033 & ~n1055 ;
  assign n1077 = ~n1075 & n1076 ;
  assign n1078 = n1074 & ~n1077 ;
  assign n1079 = n806 & n1049 ;
  assign n1080 = n815 & n1079 ;
  assign n1081 = n993 & n1080 ;
  assign n1082 = ~n814 & ~n816 ;
  assign n1083 = ~n648 & n1082 ;
  assign n1084 = ~\38(11)_pad  & ~n820 ;
  assign n1085 = ~n825 & ~n1084 ;
  assign n1086 = ~\38(11)_pad  & ~\440(277)_pad  ;
  assign n1087 = n825 & n1086 ;
  assign n1088 = ~n1085 & ~n1087 ;
  assign n1089 = ~n813 & n1088 ;
  assign n1090 = ~n1083 & n1089 ;
  assign n1091 = ~n1081 & n1090 ;
  assign n1092 = ~n813 & ~n1083 ;
  assign n1093 = ~n1081 & n1092 ;
  assign n1094 = \38(11)_pad  & n820 ;
  assign n1095 = ~n825 & ~n1094 ;
  assign n1096 = \38(11)_pad  & \438(274)_pad  ;
  assign n1097 = n820 & n1096 ;
  assign n1098 = ~n1095 & ~n1097 ;
  assign n1099 = ~n1093 & ~n1098 ;
  assign n1100 = ~n1091 & ~n1099 ;
  assign n1101 = ~n1078 & ~n1100 ;
  assign n1102 = n1078 & n1100 ;
  assign n1103 = ~n1101 & ~n1102 ;
  assign n1104 = ~n660 & n700 ;
  assign n1105 = ~n677 & n1104 ;
  assign n1106 = n700 & n778 ;
  assign n1107 = ~n1105 & ~n1106 ;
  assign n1108 = n756 & ~n1105 ;
  assign n1109 = n769 & n1108 ;
  assign n1110 = ~n1107 & ~n1109 ;
  assign n1111 = n660 & ~n700 ;
  assign n1112 = n676 & ~n700 ;
  assign n1113 = ~n673 & n1112 ;
  assign n1114 = ~n1111 & ~n1113 ;
  assign n1115 = ~n778 & ~n1114 ;
  assign n1116 = n756 & ~n1114 ;
  assign n1117 = n769 & n1116 ;
  assign n1118 = ~n1115 & ~n1117 ;
  assign n1119 = ~n1110 & n1118 ;
  assign n1120 = ~n681 & ~n788 ;
  assign n1121 = ~n695 & n1120 ;
  assign n1122 = ~n721 & ~n795 ;
  assign n1123 = ~n721 & n793 ;
  assign n1124 = ~n792 & n1123 ;
  assign n1125 = ~n1122 & ~n1124 ;
  assign n1126 = n1120 & n1125 ;
  assign n1127 = ~n1121 & ~n1126 ;
  assign n1128 = ~n678 & ~n778 ;
  assign n1129 = ~n678 & n756 ;
  assign n1130 = n769 & n1129 ;
  assign n1131 = ~n1128 & ~n1130 ;
  assign n1132 = n712 & n723 ;
  assign n1133 = ~n1121 & n1132 ;
  assign n1134 = n1131 & n1133 ;
  assign n1135 = ~n1127 & ~n1134 ;
  assign n1136 = n728 & ~n1135 ;
  assign n1137 = ~n728 & n1135 ;
  assign n1138 = ~n1136 & ~n1137 ;
  assign n1139 = n1131 & n1132 ;
  assign n1140 = ~n687 & ~n786 ;
  assign n1141 = n1125 & ~n1140 ;
  assign n1142 = ~n1139 & n1141 ;
  assign n1143 = ~n686 & n692 ;
  assign n1144 = ~n687 & ~n1143 ;
  assign n1145 = ~n683 & n1144 ;
  assign n1146 = ~n1142 & n1145 ;
  assign n1147 = ~n1142 & n1144 ;
  assign n1148 = n683 & ~n1147 ;
  assign n1149 = ~n1146 & ~n1148 ;
  assign n1150 = n693 & n1125 ;
  assign n1151 = ~n1139 & n1150 ;
  assign n1152 = ~n688 & ~n692 ;
  assign n1153 = n688 & n692 ;
  assign n1154 = ~n1152 & ~n1153 ;
  assign n1155 = ~n1151 & ~n1154 ;
  assign n1156 = n694 & n1125 ;
  assign n1157 = ~n1139 & n1156 ;
  assign n1158 = ~n1155 & ~n1157 ;
  assign n1159 = ~n693 & ~n1125 ;
  assign n1160 = ~n693 & n1132 ;
  assign n1161 = n1131 & n1160 ;
  assign n1162 = ~n1159 & ~n1161 ;
  assign n1163 = ~n1151 & n1162 ;
  assign n1164 = ~n709 & ~n792 ;
  assign n1165 = ~n716 & ~n1164 ;
  assign n1166 = ~n715 & ~n1165 ;
  assign n1167 = n712 & ~n715 ;
  assign n1168 = n1131 & n1167 ;
  assign n1169 = ~n1166 & ~n1168 ;
  assign n1170 = n722 & ~n1169 ;
  assign n1171 = ~n722 & n1169 ;
  assign n1172 = ~n1170 & ~n1171 ;
  assign n1173 = ~n717 & n1164 ;
  assign n1174 = n712 & ~n717 ;
  assign n1175 = n1131 & n1174 ;
  assign n1176 = ~n1173 & ~n1175 ;
  assign n1177 = n712 & n1131 ;
  assign n1178 = n717 & ~n1164 ;
  assign n1179 = ~n1177 & n1178 ;
  assign n1180 = n1176 & ~n1179 ;
  assign n1181 = ~n698 & ~n704 ;
  assign n1182 = ~n1110 & n1181 ;
  assign n1183 = ~n703 & n710 ;
  assign n1184 = ~n1182 & n1183 ;
  assign n1185 = n703 & ~n710 ;
  assign n1186 = ~n710 & n1181 ;
  assign n1187 = ~n1110 & n1186 ;
  assign n1188 = ~n1185 & ~n1187 ;
  assign n1189 = ~n1184 & n1188 ;
  assign n1190 = ~n698 & ~n1110 ;
  assign n1191 = ~n705 & ~n1190 ;
  assign n1192 = ~n698 & n705 ;
  assign n1193 = ~n1110 & n1192 ;
  assign n1194 = ~n1191 & ~n1193 ;
  assign n1195 = ~n705 & ~n710 ;
  assign n1196 = ~n711 & ~n1195 ;
  assign n1197 = ~n790 & ~n1181 ;
  assign n1198 = n794 & n1197 ;
  assign n1199 = ~n716 & n1197 ;
  assign n1200 = ~n1164 & n1199 ;
  assign n1201 = ~n1198 & ~n1200 ;
  assign n1202 = ~n794 & ~n1197 ;
  assign n1203 = ~n1165 & n1202 ;
  assign n1204 = n1201 & ~n1203 ;
  assign n1205 = n1119 & ~n1204 ;
  assign n1206 = ~n1118 & n1204 ;
  assign n1207 = ~n712 & ~n1164 ;
  assign n1208 = n699 & n704 ;
  assign n1209 = ~n699 & n703 ;
  assign n1210 = ~n1208 & ~n1209 ;
  assign n1211 = n715 & n1210 ;
  assign n1212 = ~n1207 & n1211 ;
  assign n1213 = n716 & n1210 ;
  assign n1214 = n1207 & n1213 ;
  assign n1215 = ~n1212 & ~n1214 ;
  assign n1216 = ~n715 & ~n1210 ;
  assign n1217 = ~n1207 & n1216 ;
  assign n1218 = ~n716 & ~n1210 ;
  assign n1219 = n1207 & n1218 ;
  assign n1220 = ~n1217 & ~n1219 ;
  assign n1221 = n1215 & n1220 ;
  assign n1222 = n1110 & n1221 ;
  assign n1223 = ~n1206 & ~n1222 ;
  assign n1224 = ~n1205 & n1223 ;
  assign n1225 = n1196 & ~n1224 ;
  assign n1226 = ~n1196 & n1223 ;
  assign n1227 = ~n1205 & n1226 ;
  assign n1228 = ~n717 & ~n722 ;
  assign n1229 = ~n723 & ~n1228 ;
  assign n1230 = n683 & ~n728 ;
  assign n1231 = ~n1229 & n1230 ;
  assign n1232 = ~n683 & ~n728 ;
  assign n1233 = n1229 & n1232 ;
  assign n1234 = ~n1231 & ~n1233 ;
  assign n1235 = ~n683 & n728 ;
  assign n1236 = ~n1229 & n1235 ;
  assign n1237 = n683 & n728 ;
  assign n1238 = n1229 & n1237 ;
  assign n1239 = ~n1236 & ~n1238 ;
  assign n1240 = n1234 & n1239 ;
  assign n1241 = ~n1227 & ~n1240 ;
  assign n1242 = ~n1225 & n1241 ;
  assign n1243 = ~n681 & ~n1140 ;
  assign n1244 = ~n788 & ~n1243 ;
  assign n1245 = ~n1154 & n1244 ;
  assign n1246 = n1154 & ~n1244 ;
  assign n1247 = ~n1245 & ~n1246 ;
  assign n1248 = n1125 & n1247 ;
  assign n1249 = ~n1139 & n1248 ;
  assign n1250 = n1121 & n1144 ;
  assign n1251 = n688 & n691 ;
  assign n1252 = ~n688 & ~n691 ;
  assign n1253 = ~n1251 & ~n1252 ;
  assign n1254 = \530(216)_pad  & n685 ;
  assign n1255 = n690 & n1254 ;
  assign n1256 = \528(214)_pad  & \530(216)_pad  ;
  assign n1257 = n690 & n1256 ;
  assign n1258 = ~n687 & ~n1257 ;
  assign n1259 = ~n1255 & n1258 ;
  assign n1260 = n681 & ~n1259 ;
  assign n1261 = n1253 & ~n1260 ;
  assign n1262 = ~n1250 & n1261 ;
  assign n1263 = ~n1253 & n1260 ;
  assign n1264 = n1144 & ~n1253 ;
  assign n1265 = n1121 & n1264 ;
  assign n1266 = ~n1263 & ~n1265 ;
  assign n1267 = ~n1125 & n1266 ;
  assign n1268 = n1132 & n1266 ;
  assign n1269 = n1131 & n1268 ;
  assign n1270 = ~n1267 & ~n1269 ;
  assign n1271 = ~n1262 & ~n1270 ;
  assign n1272 = ~n1249 & ~n1271 ;
  assign n1273 = n1196 & n1240 ;
  assign n1274 = ~n1224 & n1273 ;
  assign n1275 = ~n1196 & n1240 ;
  assign n1276 = n1224 & n1275 ;
  assign n1277 = ~n1274 & ~n1276 ;
  assign n1278 = n1272 & n1277 ;
  assign n1279 = ~n1242 & n1278 ;
  assign n1280 = ~n1272 & ~n1277 ;
  assign n1281 = ~n1225 & ~n1272 ;
  assign n1282 = n1241 & n1281 ;
  assign n1283 = ~n1280 & ~n1282 ;
  assign n1284 = ~n1279 & n1283 ;
  assign n1285 = \4526(205)_pad  & n762 ;
  assign n1286 = ~\18(5)_pad  & ~\4526(205)_pad  ;
  assign n1287 = \41(12)_pad  & ~\542(246)_pad  ;
  assign n1288 = n1286 & n1287 ;
  assign n1289 = ~\41(12)_pad  & ~\4526(205)_pad  ;
  assign n1290 = n759 & n1289 ;
  assign n1291 = ~n1288 & ~n1290 ;
  assign n1292 = ~n1285 & n1291 ;
  assign n1293 = ~n673 & ~n674 ;
  assign n1294 = n756 & n1293 ;
  assign n1295 = n769 & n1294 ;
  assign n1296 = n774 & n775 ;
  assign n1297 = n1293 & ~n1296 ;
  assign n1298 = ~n776 & ~n1297 ;
  assign n1299 = ~n1295 & n1298 ;
  assign n1300 = n776 & n1293 ;
  assign n1301 = n756 & n1300 ;
  assign n1302 = n769 & n1301 ;
  assign n1303 = ~n674 & n776 ;
  assign n1304 = ~n673 & n1303 ;
  assign n1305 = ~n1296 & n1304 ;
  assign n1306 = ~n1302 & ~n1305 ;
  assign n1307 = ~n1299 & n1306 ;
  assign n1308 = ~n667 & ~n671 ;
  assign n1309 = n756 & ~n1308 ;
  assign n1310 = n769 & n1309 ;
  assign n1311 = ~n663 & n772 ;
  assign n1312 = ~n671 & ~n1311 ;
  assign n1313 = ~n775 & n1312 ;
  assign n1314 = ~n1310 & n1313 ;
  assign n1315 = n775 & ~n1312 ;
  assign n1316 = n775 & ~n1308 ;
  assign n1317 = n756 & n1316 ;
  assign n1318 = n769 & n1317 ;
  assign n1319 = ~n1315 & ~n1318 ;
  assign n1320 = ~n1314 & n1319 ;
  assign n1321 = ~n757 & n773 ;
  assign n1322 = ~n768 & n1321 ;
  assign n1323 = n756 & n1322 ;
  assign n1324 = n771 & ~n772 ;
  assign n1325 = ~n771 & n772 ;
  assign n1326 = ~n1324 & ~n1325 ;
  assign n1327 = ~n1323 & n1326 ;
  assign n1328 = n756 & n774 ;
  assign n1329 = n769 & n1328 ;
  assign n1330 = ~n1327 & ~n1329 ;
  assign n1331 = ~n770 & ~n773 ;
  assign n1332 = ~n1323 & ~n1331 ;
  assign n1333 = ~n739 & ~n757 ;
  assign n1334 = ~n746 & ~n750 ;
  assign n1335 = n763 & n1285 ;
  assign n1336 = n1334 & ~n1335 ;
  assign n1337 = ~n735 & ~n736 ;
  assign n1338 = n758 & n1337 ;
  assign n1339 = ~n1336 & n1338 ;
  assign n1340 = n749 & n1337 ;
  assign n1341 = ~n735 & ~n1340 ;
  assign n1342 = ~n1339 & n1341 ;
  assign n1343 = ~n1333 & ~n1342 ;
  assign n1344 = ~n735 & n1333 ;
  assign n1345 = ~n1340 & n1344 ;
  assign n1346 = ~n1339 & n1345 ;
  assign n1347 = ~n1343 & ~n1346 ;
  assign n1348 = ~n1339 & ~n1340 ;
  assign n1349 = n758 & ~n1336 ;
  assign n1350 = ~n749 & ~n1337 ;
  assign n1351 = ~n1349 & n1350 ;
  assign n1352 = n1348 & ~n1351 ;
  assign n1353 = ~n758 & n1336 ;
  assign n1354 = ~n1349 & ~n1353 ;
  assign n1355 = ~\4526(205)_pad  & \542(246)_pad  ;
  assign n1356 = ~n1289 & ~n1355 ;
  assign n1357 = \18(5)_pad  & ~\4526(205)_pad  ;
  assign n1358 = ~\18(5)_pad  & ~\41(12)_pad  ;
  assign n1359 = \542(246)_pad  & n1358 ;
  assign n1360 = ~n1357 & ~n1359 ;
  assign n1361 = n1356 & n1360 ;
  assign n1362 = n763 & n1361 ;
  assign n1363 = ~n763 & ~n1361 ;
  assign n1364 = ~n1362 & ~n1363 ;
  assign n1365 = ~n674 & ~n1308 ;
  assign n1366 = ~n673 & ~n1365 ;
  assign n1367 = ~n1326 & ~n1366 ;
  assign n1368 = n1326 & n1366 ;
  assign n1369 = ~n1367 & ~n1368 ;
  assign n1370 = n770 & n1369 ;
  assign n1371 = n666 & n771 ;
  assign n1372 = ~n666 & ~n771 ;
  assign n1373 = ~n1371 & ~n1372 ;
  assign n1374 = n674 & ~n774 ;
  assign n1375 = ~n1308 & n1374 ;
  assign n1376 = ~n1373 & n1375 ;
  assign n1377 = n1312 & ~n1373 ;
  assign n1378 = n1297 & n1377 ;
  assign n1379 = ~n1376 & ~n1378 ;
  assign n1380 = n1297 & n1312 ;
  assign n1381 = n1373 & ~n1375 ;
  assign n1382 = ~n1380 & n1381 ;
  assign n1383 = ~n770 & ~n1382 ;
  assign n1384 = n1379 & n1383 ;
  assign n1385 = ~n1370 & ~n1384 ;
  assign n1386 = ~n752 & ~n753 ;
  assign n1387 = n758 & n764 ;
  assign n1388 = ~n1386 & ~n1387 ;
  assign n1389 = ~n736 & ~n1388 ;
  assign n1390 = ~n735 & ~n1386 ;
  assign n1391 = ~n1387 & n1390 ;
  assign n1392 = ~n1389 & ~n1391 ;
  assign n1393 = n750 & ~n761 ;
  assign n1394 = n745 & ~n761 ;
  assign n1395 = ~n744 & n1394 ;
  assign n1396 = ~n1393 & ~n1395 ;
  assign n1397 = ~n761 & ~n764 ;
  assign n1398 = n1334 & ~n1397 ;
  assign n1399 = n1396 & ~n1398 ;
  assign n1400 = n1285 & ~n1399 ;
  assign n1401 = ~n1392 & n1400 ;
  assign n1402 = n1285 & n1399 ;
  assign n1403 = n1392 & n1402 ;
  assign n1404 = ~n1401 & ~n1403 ;
  assign n1405 = ~n745 & ~n750 ;
  assign n1406 = ~n746 & ~n1405 ;
  assign n1407 = n736 & ~n1406 ;
  assign n1408 = n1386 & n1407 ;
  assign n1409 = n735 & ~n1406 ;
  assign n1410 = ~n1386 & n1409 ;
  assign n1411 = ~n1408 & ~n1410 ;
  assign n1412 = ~n735 & n1406 ;
  assign n1413 = ~n1386 & n1412 ;
  assign n1414 = ~n736 & n1406 ;
  assign n1415 = n1386 & n1414 ;
  assign n1416 = ~n1413 & ~n1415 ;
  assign n1417 = n1411 & n1416 ;
  assign n1418 = ~n1291 & n1417 ;
  assign n1419 = n1292 & ~n1417 ;
  assign n1420 = ~n1418 & ~n1419 ;
  assign n1421 = n1404 & n1420 ;
  assign n1422 = n1385 & n1421 ;
  assign n1423 = ~n1385 & ~n1421 ;
  assign n1424 = ~n1422 & ~n1423 ;
  assign n1425 = n758 & ~n1337 ;
  assign n1426 = ~n758 & n1337 ;
  assign n1427 = ~n1425 & ~n1426 ;
  assign n1428 = ~n776 & n1333 ;
  assign n1429 = ~n1427 & n1428 ;
  assign n1430 = n776 & n1333 ;
  assign n1431 = n1427 & n1430 ;
  assign n1432 = ~n1429 & ~n1431 ;
  assign n1433 = n776 & ~n1333 ;
  assign n1434 = ~n1427 & n1433 ;
  assign n1435 = ~n776 & ~n1333 ;
  assign n1436 = n1427 & n1435 ;
  assign n1437 = ~n1434 & ~n1436 ;
  assign n1438 = n1432 & n1437 ;
  assign n1439 = n763 & ~n775 ;
  assign n1440 = ~n763 & n775 ;
  assign n1441 = ~n1439 & ~n1440 ;
  assign n1442 = ~n1438 & ~n1441 ;
  assign n1443 = ~n1424 & n1442 ;
  assign n1444 = ~n1438 & n1441 ;
  assign n1445 = n1424 & n1444 ;
  assign n1446 = ~n1443 & ~n1445 ;
  assign n1447 = n1438 & ~n1441 ;
  assign n1448 = n1424 & n1447 ;
  assign n1449 = n1438 & n1441 ;
  assign n1450 = ~n1424 & n1449 ;
  assign n1451 = ~n1448 & ~n1450 ;
  assign n1452 = n1446 & n1451 ;
  assign n1453 = ~\5(1)_pad  & ~\57(20)_pad  ;
  assign n1454 = \228(151)_pad  & \240(163)_pad  ;
  assign n1455 = \150(73)_pad  & \184(107)_pad  ;
  assign n1456 = n1454 & n1455 ;
  assign n1457 = \218(141)_pad  & \230(153)_pad  ;
  assign n1458 = \152(75)_pad  & \210(133)_pad  ;
  assign n1459 = n1457 & n1458 ;
  assign n1460 = \185(108)_pad  & \186(109)_pad  ;
  assign n1461 = \182(105)_pad  & \183(106)_pad  ;
  assign n1462 = n1460 & n1461 ;
  assign n1463 = \188(111)_pad  & \199(122)_pad  ;
  assign n1464 = \162(85)_pad  & \172(95)_pad  ;
  assign n1465 = n1463 & n1464 ;
  assign n1466 = n685 & ~n702 ;
  assign n1467 = ~n685 & n702 ;
  assign n1468 = ~n1466 & ~n1467 ;
  assign n1469 = n680 & ~n707 ;
  assign n1470 = ~n680 & n707 ;
  assign n1471 = ~n1469 & ~n1470 ;
  assign n1472 = n1468 & ~n1471 ;
  assign n1473 = ~n1468 & n1471 ;
  assign n1474 = ~n1472 & ~n1473 ;
  assign n1475 = ~n714 & ~n1474 ;
  assign n1476 = n714 & n1474 ;
  assign n1477 = ~n1475 & ~n1476 ;
  assign n1478 = \115(60)_pad  & ~\18(5)_pad  ;
  assign n1479 = \18(5)_pad  & \227(150)_pad  ;
  assign n1480 = ~n1478 & ~n1479 ;
  assign n1481 = n719 & n1480 ;
  assign n1482 = ~n719 & ~n1480 ;
  assign n1483 = ~n1481 & ~n1482 ;
  assign n1484 = ~n697 & ~n725 ;
  assign n1485 = n690 & n1484 ;
  assign n1486 = n1483 & n1485 ;
  assign n1487 = ~n697 & n725 ;
  assign n1488 = n690 & n1487 ;
  assign n1489 = ~n1483 & n1488 ;
  assign n1490 = ~n1486 & ~n1489 ;
  assign n1491 = n697 & ~n725 ;
  assign n1492 = n690 & n1491 ;
  assign n1493 = ~n1483 & n1492 ;
  assign n1494 = n697 & n725 ;
  assign n1495 = n690 & n1494 ;
  assign n1496 = n1483 & n1495 ;
  assign n1497 = ~n1493 & ~n1496 ;
  assign n1498 = n1490 & n1497 ;
  assign n1499 = ~n690 & n1487 ;
  assign n1500 = n1483 & n1499 ;
  assign n1501 = ~n690 & n1484 ;
  assign n1502 = ~n1483 & n1501 ;
  assign n1503 = ~n1500 & ~n1502 ;
  assign n1504 = ~n690 & n1491 ;
  assign n1505 = n1483 & n1504 ;
  assign n1506 = ~n690 & n1494 ;
  assign n1507 = ~n1483 & n1506 ;
  assign n1508 = ~n1505 & ~n1507 ;
  assign n1509 = n1503 & n1508 ;
  assign n1510 = n1498 & n1509 ;
  assign n1511 = n1477 & ~n1510 ;
  assign n1512 = ~n1477 & n1510 ;
  assign n1513 = \211(134)_pad  & ~\212(135)_pad  ;
  assign n1514 = ~\211(134)_pad  & \212(135)_pad  ;
  assign n1515 = ~n1513 & ~n1514 ;
  assign n1516 = \209(132)_pad  & n1515 ;
  assign n1517 = \18(5)_pad  & ~n396 ;
  assign n1518 = ~\209(132)_pad  & ~n1515 ;
  assign n1519 = n1517 & ~n1518 ;
  assign n1520 = ~n1516 & n1519 ;
  assign n1521 = \215(138)_pad  & \216(139)_pad  ;
  assign n1522 = ~\215(138)_pad  & ~\216(139)_pad  ;
  assign n1523 = ~n1521 & ~n1522 ;
  assign n1524 = n1517 & n1523 ;
  assign n1525 = \213(136)_pad  & \214(137)_pad  ;
  assign n1526 = ~\213(136)_pad  & ~\214(137)_pad  ;
  assign n1527 = ~n1525 & ~n1526 ;
  assign n1528 = n1517 & n1527 ;
  assign n1529 = ~n1524 & ~n1528 ;
  assign n1530 = ~n1520 & n1529 ;
  assign n1531 = ~n1524 & n1528 ;
  assign n1532 = n1520 & n1531 ;
  assign n1533 = ~n1530 & ~n1532 ;
  assign n1534 = ~n1520 & ~n1528 ;
  assign n1535 = ~n1516 & n1528 ;
  assign n1536 = n1519 & n1535 ;
  assign n1537 = n1524 & ~n1536 ;
  assign n1538 = ~n1534 & n1537 ;
  assign n1539 = n1533 & ~n1538 ;
  assign n1540 = ~n1512 & ~n1539 ;
  assign n1541 = ~n1511 & n1540 ;
  assign n1542 = n665 & n738 ;
  assign n1543 = ~n665 & ~n738 ;
  assign n1544 = ~n1542 & ~n1543 ;
  assign n1545 = ~n659 & ~n669 ;
  assign n1546 = ~n1544 & n1545 ;
  assign n1547 = ~n659 & n669 ;
  assign n1548 = n1544 & n1547 ;
  assign n1549 = ~n1546 & ~n1548 ;
  assign n1550 = n659 & n669 ;
  assign n1551 = ~n1544 & n1550 ;
  assign n1552 = n659 & ~n669 ;
  assign n1553 = n1544 & n1552 ;
  assign n1554 = ~n1551 & ~n1553 ;
  assign n1555 = n1549 & n1554 ;
  assign n1556 = n734 & n748 ;
  assign n1557 = ~n734 & ~n748 ;
  assign n1558 = ~n1556 & ~n1557 ;
  assign n1559 = n662 & ~n1558 ;
  assign n1560 = ~n662 & n1558 ;
  assign n1561 = ~n1559 & ~n1560 ;
  assign n1562 = ~\18(5)_pad  & \44(13)_pad  ;
  assign n1563 = \18(5)_pad  & \239(162)_pad  ;
  assign n1564 = ~n1562 & ~n1563 ;
  assign n1565 = \18(5)_pad  & \229(152)_pad  ;
  assign n1566 = ~n265 & ~n1565 ;
  assign n1567 = n743 & n1566 ;
  assign n1568 = ~n743 & ~n1566 ;
  assign n1569 = ~n1567 & ~n1568 ;
  assign n1570 = ~n1564 & ~n1569 ;
  assign n1571 = ~n1561 & n1570 ;
  assign n1572 = ~n1555 & n1571 ;
  assign n1573 = ~n1564 & n1569 ;
  assign n1574 = ~n1561 & n1573 ;
  assign n1575 = n1555 & n1574 ;
  assign n1576 = ~n1572 & ~n1575 ;
  assign n1577 = n1564 & ~n1569 ;
  assign n1578 = ~n1561 & n1577 ;
  assign n1579 = n1555 & n1578 ;
  assign n1580 = n1564 & n1569 ;
  assign n1581 = ~n1561 & n1580 ;
  assign n1582 = ~n1555 & n1581 ;
  assign n1583 = ~n1579 & ~n1582 ;
  assign n1584 = n1576 & n1583 ;
  assign n1585 = n1561 & n1570 ;
  assign n1586 = n1555 & n1585 ;
  assign n1587 = n1561 & n1573 ;
  assign n1588 = ~n1555 & n1587 ;
  assign n1589 = ~n1586 & ~n1588 ;
  assign n1590 = n1561 & n1577 ;
  assign n1591 = ~n1555 & n1590 ;
  assign n1592 = n1561 & n1580 ;
  assign n1593 = n1555 & n1592 ;
  assign n1594 = ~n1591 & ~n1593 ;
  assign n1595 = n1589 & n1594 ;
  assign n1596 = n1584 & n1595 ;
  assign n1597 = n582 & n587 ;
  assign n1598 = ~n582 & ~n587 ;
  assign n1599 = ~n1597 & ~n1598 ;
  assign n1600 = n594 & ~n1599 ;
  assign n1601 = ~n594 & n1599 ;
  assign n1602 = ~n1600 & ~n1601 ;
  assign n1603 = ~\153(76)_pad  & ~\154(77)_pad  ;
  assign n1604 = \18(5)_pad  & ~n1603 ;
  assign n1605 = \153(76)_pad  & \154(77)_pad  ;
  assign n1606 = ~n396 & ~n1605 ;
  assign n1607 = n1604 & n1606 ;
  assign n1608 = n577 & n1607 ;
  assign n1609 = ~n577 & ~n1607 ;
  assign n1610 = ~n1608 & ~n1609 ;
  assign n1611 = \161(84)_pad  & \18(5)_pad  ;
  assign n1612 = \141(70)_pad  & ~\18(5)_pad  ;
  assign n1613 = ~n1611 & ~n1612 ;
  assign n1614 = ~n599 & ~n1613 ;
  assign n1615 = n599 & n1613 ;
  assign n1616 = ~n1614 & ~n1615 ;
  assign n1617 = ~\155(78)_pad  & ~\156(79)_pad  ;
  assign n1618 = \18(5)_pad  & ~n1617 ;
  assign n1619 = \155(78)_pad  & \156(79)_pad  ;
  assign n1620 = ~n396 & ~n1619 ;
  assign n1621 = n1618 & n1620 ;
  assign n1622 = ~n1616 & n1621 ;
  assign n1623 = ~n1610 & n1622 ;
  assign n1624 = ~n1616 & ~n1621 ;
  assign n1625 = n1610 & n1624 ;
  assign n1626 = ~n1623 & ~n1625 ;
  assign n1627 = n1616 & ~n1621 ;
  assign n1628 = ~n1610 & n1627 ;
  assign n1629 = n1616 & n1621 ;
  assign n1630 = n1610 & n1629 ;
  assign n1631 = ~n1628 & ~n1630 ;
  assign n1632 = n1626 & n1631 ;
  assign n1633 = ~n1602 & n1632 ;
  assign n1634 = n1602 & ~n1632 ;
  assign n1635 = ~n1633 & ~n1634 ;
  assign n1636 = ~n1596 & n1635 ;
  assign n1637 = n1541 & n1636 ;
  assign n1638 = n401 & ~n407 ;
  assign n1639 = ~n401 & n407 ;
  assign n1640 = ~n1638 & ~n1639 ;
  assign n1641 = n418 & n1640 ;
  assign n1642 = ~n418 & ~n1640 ;
  assign n1643 = ~n1641 & ~n1642 ;
  assign n1644 = ~\438(274)_pad  & ~\440(277)_pad  ;
  assign n1645 = \438(274)_pad  & \440(277)_pad  ;
  assign n1646 = ~n1644 & ~n1645 ;
  assign n1647 = \18(5)_pad  & ~n1646 ;
  assign n1648 = ~n423 & ~n432 ;
  assign n1649 = ~\18(5)_pad  & ~n1648 ;
  assign n1650 = ~n1647 & ~n1649 ;
  assign n1651 = \18(5)_pad  & ~\450(288)_pad  ;
  assign n1652 = \114(59)_pad  & ~\18(5)_pad  ;
  assign n1653 = ~n1651 & ~n1652 ;
  assign n1654 = n430 & n440 ;
  assign n1655 = ~n430 & ~n440 ;
  assign n1656 = ~n1654 & ~n1655 ;
  assign n1657 = n1653 & ~n1656 ;
  assign n1658 = ~n1653 & n1656 ;
  assign n1659 = ~n1657 & ~n1658 ;
  assign n1660 = ~n1650 & n1659 ;
  assign n1661 = n1650 & ~n1659 ;
  assign n1662 = ~n1660 & ~n1661 ;
  assign n1663 = ~n1643 & ~n1662 ;
  assign n1664 = n1643 & n1662 ;
  assign n1665 = ~n1663 & ~n1664 ;
  assign n1666 = n261 & n316 ;
  assign n1667 = ~n261 & ~n316 ;
  assign n1668 = ~n1666 & ~n1667 ;
  assign n1669 = ~n252 & n290 ;
  assign n1670 = ~n275 & n1669 ;
  assign n1671 = n1668 & n1670 ;
  assign n1672 = n252 & n290 ;
  assign n1673 = ~n275 & n1672 ;
  assign n1674 = ~n1668 & n1673 ;
  assign n1675 = ~n1671 & ~n1674 ;
  assign n1676 = n275 & n1669 ;
  assign n1677 = ~n1668 & n1676 ;
  assign n1678 = n275 & n1672 ;
  assign n1679 = n1668 & n1678 ;
  assign n1680 = ~n1677 & ~n1679 ;
  assign n1681 = n1675 & n1680 ;
  assign n1682 = n252 & ~n290 ;
  assign n1683 = ~n275 & n1682 ;
  assign n1684 = n1668 & n1683 ;
  assign n1685 = ~n252 & ~n290 ;
  assign n1686 = ~n275 & n1685 ;
  assign n1687 = ~n1668 & n1686 ;
  assign n1688 = ~n1684 & ~n1687 ;
  assign n1689 = n275 & n1685 ;
  assign n1690 = n1668 & n1689 ;
  assign n1691 = n275 & n1682 ;
  assign n1692 = ~n1668 & n1691 ;
  assign n1693 = ~n1690 & ~n1692 ;
  assign n1694 = n1688 & n1693 ;
  assign n1695 = n1681 & n1694 ;
  assign n1696 = ~\18(5)_pad  & ~\69(30)_pad  ;
  assign n1697 = \18(5)_pad  & \560(248)_pad  ;
  assign n1698 = ~n1696 & ~n1697 ;
  assign n1699 = n245 & n1698 ;
  assign n1700 = ~n245 & ~n1698 ;
  assign n1701 = ~n1699 & ~n1700 ;
  assign n1702 = \18(5)_pad  & \542(246)_pad  ;
  assign n1703 = ~n267 & ~n1702 ;
  assign n1704 = n297 & ~n1703 ;
  assign n1705 = ~n305 & n1704 ;
  assign n1706 = n1701 & n1705 ;
  assign n1707 = ~n297 & ~n1703 ;
  assign n1708 = ~n305 & n1707 ;
  assign n1709 = ~n1701 & n1708 ;
  assign n1710 = ~n1706 & ~n1709 ;
  assign n1711 = n297 & n1703 ;
  assign n1712 = ~n305 & n1711 ;
  assign n1713 = ~n1701 & n1712 ;
  assign n1714 = ~n297 & n1703 ;
  assign n1715 = ~n305 & n1714 ;
  assign n1716 = n1701 & n1715 ;
  assign n1717 = ~n1713 & ~n1716 ;
  assign n1718 = n1710 & n1717 ;
  assign n1719 = n305 & n1707 ;
  assign n1720 = n1701 & n1719 ;
  assign n1721 = n305 & n1704 ;
  assign n1722 = ~n1701 & n1721 ;
  assign n1723 = ~n1720 & ~n1722 ;
  assign n1724 = n305 & n1714 ;
  assign n1725 = ~n1701 & n1724 ;
  assign n1726 = n305 & n1711 ;
  assign n1727 = n1701 & n1726 ;
  assign n1728 = ~n1725 & ~n1727 ;
  assign n1729 = n1723 & n1728 ;
  assign n1730 = n1718 & n1729 ;
  assign n1731 = ~n1695 & ~n1730 ;
  assign n1732 = n1695 & n1730 ;
  assign n1733 = ~n1731 & ~n1732 ;
  assign n1734 = ~n1665 & n1733 ;
  assign n1735 = n464 & n484 ;
  assign n1736 = ~n464 & ~n484 ;
  assign n1737 = ~n1735 & ~n1736 ;
  assign n1738 = n508 & n524 ;
  assign n1739 = ~n1737 & n1738 ;
  assign n1740 = ~n508 & n524 ;
  assign n1741 = n1737 & n1740 ;
  assign n1742 = ~n1739 & ~n1741 ;
  assign n1743 = ~n508 & ~n524 ;
  assign n1744 = ~n1737 & n1743 ;
  assign n1745 = n508 & ~n524 ;
  assign n1746 = n1737 & n1745 ;
  assign n1747 = ~n1744 & ~n1746 ;
  assign n1748 = n1742 & n1747 ;
  assign n1749 = n492 & n502 ;
  assign n1750 = ~n492 & ~n502 ;
  assign n1751 = ~n1749 & ~n1750 ;
  assign n1752 = n517 & ~n1751 ;
  assign n1753 = ~n517 & n1751 ;
  assign n1754 = ~n1752 & ~n1753 ;
  assign n1755 = ~\18(5)_pad  & ~\82(41)_pad  ;
  assign n1756 = \18(5)_pad  & \496(271)_pad  ;
  assign n1757 = ~n1755 & ~n1756 ;
  assign n1758 = n478 & n1757 ;
  assign n1759 = ~n478 & ~n1757 ;
  assign n1760 = ~n1758 & ~n1759 ;
  assign n1761 = ~n471 & ~n1760 ;
  assign n1762 = n1754 & n1761 ;
  assign n1763 = ~n1748 & n1762 ;
  assign n1764 = n471 & ~n1760 ;
  assign n1765 = n1754 & n1764 ;
  assign n1766 = n1748 & n1765 ;
  assign n1767 = ~n1763 & ~n1766 ;
  assign n1768 = ~n1754 & n1764 ;
  assign n1769 = ~n1748 & n1768 ;
  assign n1770 = ~n1754 & n1761 ;
  assign n1771 = n1748 & n1770 ;
  assign n1772 = ~n1769 & ~n1771 ;
  assign n1773 = n1767 & n1772 ;
  assign n1774 = n471 & n1760 ;
  assign n1775 = n1754 & n1774 ;
  assign n1776 = ~n1748 & n1775 ;
  assign n1777 = ~n471 & n1760 ;
  assign n1778 = n1754 & n1777 ;
  assign n1779 = n1748 & n1778 ;
  assign n1780 = ~n1776 & ~n1779 ;
  assign n1781 = ~n1754 & n1777 ;
  assign n1782 = ~n1748 & n1781 ;
  assign n1783 = ~n1754 & n1774 ;
  assign n1784 = n1748 & n1783 ;
  assign n1785 = ~n1782 & ~n1784 ;
  assign n1786 = n1780 & n1785 ;
  assign n1787 = n1773 & n1786 ;
  assign n1788 = \18(5)_pad  & ~\540(227)_pad  ;
  assign n1789 = ~\18(5)_pad  & \58(21)_pad  ;
  assign n1790 = ~n1788 & ~n1789 ;
  assign n1791 = n369 & n1790 ;
  assign n1792 = ~n369 & ~n1790 ;
  assign n1793 = ~n1791 & ~n1792 ;
  assign n1794 = ~n234 & ~n353 ;
  assign n1795 = n332 & n1794 ;
  assign n1796 = ~n1793 & n1795 ;
  assign n1797 = ~n332 & n1794 ;
  assign n1798 = n1793 & n1797 ;
  assign n1799 = ~n1796 & ~n1798 ;
  assign n1800 = n234 & ~n353 ;
  assign n1801 = ~n332 & n1800 ;
  assign n1802 = ~n1793 & n1801 ;
  assign n1803 = n332 & n1800 ;
  assign n1804 = n1793 & n1803 ;
  assign n1805 = ~n1802 & ~n1804 ;
  assign n1806 = n1799 & n1805 ;
  assign n1807 = n234 & n353 ;
  assign n1808 = n332 & n1807 ;
  assign n1809 = ~n1793 & n1808 ;
  assign n1810 = ~n332 & n1807 ;
  assign n1811 = n1793 & n1810 ;
  assign n1812 = ~n1809 & ~n1811 ;
  assign n1813 = ~n234 & n353 ;
  assign n1814 = ~n332 & n1813 ;
  assign n1815 = ~n1793 & n1814 ;
  assign n1816 = n332 & n1813 ;
  assign n1817 = n1793 & n1816 ;
  assign n1818 = ~n1815 & ~n1817 ;
  assign n1819 = n1812 & n1818 ;
  assign n1820 = n1806 & n1819 ;
  assign n1821 = ~n212 & n227 ;
  assign n1822 = n212 & ~n227 ;
  assign n1823 = ~n1821 & ~n1822 ;
  assign n1824 = n219 & ~n381 ;
  assign n1825 = ~n219 & n381 ;
  assign n1826 = ~n1824 & ~n1825 ;
  assign n1827 = n360 & n1826 ;
  assign n1828 = ~n360 & ~n1826 ;
  assign n1829 = ~n1827 & ~n1828 ;
  assign n1830 = ~n1823 & n1829 ;
  assign n1831 = ~n1820 & n1830 ;
  assign n1832 = ~n1823 & ~n1829 ;
  assign n1833 = n1820 & n1832 ;
  assign n1834 = ~n1831 & ~n1833 ;
  assign n1835 = n1823 & ~n1829 ;
  assign n1836 = ~n1820 & n1835 ;
  assign n1837 = n1823 & n1829 ;
  assign n1838 = n1820 & n1837 ;
  assign n1839 = ~n1836 & ~n1838 ;
  assign n1840 = n1834 & n1839 ;
  assign n1841 = ~n1787 & n1840 ;
  assign n1842 = n1734 & n1841 ;
  assign n1843 = n249 & ~n294 ;
  assign n1844 = ~n249 & n294 ;
  assign n1845 = ~n1843 & ~n1844 ;
  assign n1846 = ~n287 & n313 ;
  assign n1847 = ~n1845 & n1846 ;
  assign n1848 = ~n287 & ~n313 ;
  assign n1849 = n1845 & n1848 ;
  assign n1850 = ~n1847 & ~n1849 ;
  assign n1851 = n287 & ~n313 ;
  assign n1852 = ~n1845 & n1851 ;
  assign n1853 = n287 & n313 ;
  assign n1854 = n1845 & n1853 ;
  assign n1855 = ~n1852 & ~n1854 ;
  assign n1856 = n1850 & n1855 ;
  assign n1857 = n242 & n272 ;
  assign n1858 = ~n242 & ~n272 ;
  assign n1859 = ~n1857 & ~n1858 ;
  assign n1860 = n258 & ~n1859 ;
  assign n1861 = ~n258 & n1859 ;
  assign n1862 = ~n1860 & ~n1861 ;
  assign n1863 = \18(5)_pad  & \208(131)_pad  ;
  assign n1864 = ~n1562 & ~n1863 ;
  assign n1865 = \18(5)_pad  & \198(121)_pad  ;
  assign n1866 = ~n265 & ~n1865 ;
  assign n1867 = n302 & n1866 ;
  assign n1868 = ~n302 & ~n1866 ;
  assign n1869 = ~n1867 & ~n1868 ;
  assign n1870 = ~n1864 & ~n1869 ;
  assign n1871 = ~n1862 & n1870 ;
  assign n1872 = ~n1856 & n1871 ;
  assign n1873 = ~n1864 & n1869 ;
  assign n1874 = ~n1862 & n1873 ;
  assign n1875 = n1856 & n1874 ;
  assign n1876 = ~n1872 & ~n1875 ;
  assign n1877 = n1864 & ~n1869 ;
  assign n1878 = ~n1862 & n1877 ;
  assign n1879 = n1856 & n1878 ;
  assign n1880 = n1864 & n1869 ;
  assign n1881 = ~n1862 & n1880 ;
  assign n1882 = ~n1856 & n1881 ;
  assign n1883 = ~n1879 & ~n1882 ;
  assign n1884 = n1876 & n1883 ;
  assign n1885 = n1862 & n1870 ;
  assign n1886 = n1856 & n1885 ;
  assign n1887 = n1862 & n1873 ;
  assign n1888 = ~n1856 & n1887 ;
  assign n1889 = ~n1886 & ~n1888 ;
  assign n1890 = n1862 & n1877 ;
  assign n1891 = ~n1856 & n1890 ;
  assign n1892 = n1862 & n1880 ;
  assign n1893 = n1856 & n1892 ;
  assign n1894 = ~n1891 & ~n1893 ;
  assign n1895 = n1889 & n1894 ;
  assign n1896 = n1884 & n1895 ;
  assign n1897 = n350 & n357 ;
  assign n1898 = ~n350 & ~n357 ;
  assign n1899 = ~n1897 & ~n1898 ;
  assign n1900 = n209 & n231 ;
  assign n1901 = ~n209 & ~n231 ;
  assign n1902 = ~n1900 & ~n1901 ;
  assign n1903 = ~n1899 & n1902 ;
  assign n1904 = n1899 & ~n1902 ;
  assign n1905 = ~n1903 & ~n1904 ;
  assign n1906 = ~n366 & ~n1905 ;
  assign n1907 = n366 & n1905 ;
  assign n1908 = ~n1906 & ~n1907 ;
  assign n1909 = \18(5)_pad  & \197(120)_pad  ;
  assign n1910 = ~n1478 & ~n1909 ;
  assign n1911 = n329 & n1910 ;
  assign n1912 = ~n329 & ~n1910 ;
  assign n1913 = ~n1911 & ~n1912 ;
  assign n1914 = ~n224 & ~n378 ;
  assign n1915 = ~n216 & n1914 ;
  assign n1916 = ~n1913 & n1915 ;
  assign n1917 = n224 & ~n378 ;
  assign n1918 = ~n216 & n1917 ;
  assign n1919 = n1913 & n1918 ;
  assign n1920 = ~n1916 & ~n1919 ;
  assign n1921 = n216 & n1917 ;
  assign n1922 = ~n1913 & n1921 ;
  assign n1923 = n216 & n1914 ;
  assign n1924 = n1913 & n1923 ;
  assign n1925 = ~n1922 & ~n1924 ;
  assign n1926 = n1920 & n1925 ;
  assign n1927 = ~n224 & n378 ;
  assign n1928 = n216 & n1927 ;
  assign n1929 = ~n1913 & n1928 ;
  assign n1930 = n224 & n378 ;
  assign n1931 = n216 & n1930 ;
  assign n1932 = n1913 & n1931 ;
  assign n1933 = ~n1929 & ~n1932 ;
  assign n1934 = ~n216 & n1930 ;
  assign n1935 = ~n1913 & n1934 ;
  assign n1936 = ~n216 & n1927 ;
  assign n1937 = n1913 & n1936 ;
  assign n1938 = ~n1935 & ~n1937 ;
  assign n1939 = n1933 & n1938 ;
  assign n1940 = n1926 & n1939 ;
  assign n1941 = n1908 & ~n1940 ;
  assign n1942 = ~n1908 & n1940 ;
  assign n1943 = \164(87)_pad  & ~\165(88)_pad  ;
  assign n1944 = ~\164(87)_pad  & \165(88)_pad  ;
  assign n1945 = ~n1943 & ~n1944 ;
  assign n1946 = \170(93)_pad  & n1945 ;
  assign n1947 = ~\170(93)_pad  & ~n1945 ;
  assign n1948 = n1517 & ~n1947 ;
  assign n1949 = ~n1946 & n1948 ;
  assign n1950 = ~\166(89)_pad  & ~\167(90)_pad  ;
  assign n1951 = \18(5)_pad  & ~n1950 ;
  assign n1952 = \166(89)_pad  & \167(90)_pad  ;
  assign n1953 = ~n396 & ~n1952 ;
  assign n1954 = n1951 & n1953 ;
  assign n1955 = ~\168(91)_pad  & ~\169(92)_pad  ;
  assign n1956 = \18(5)_pad  & ~n1955 ;
  assign n1957 = \168(91)_pad  & \169(92)_pad  ;
  assign n1958 = ~n396 & ~n1957 ;
  assign n1959 = n1956 & n1958 ;
  assign n1960 = ~n1954 & ~n1959 ;
  assign n1961 = ~n1949 & n1960 ;
  assign n1962 = ~n1954 & n1959 ;
  assign n1963 = n1949 & n1962 ;
  assign n1964 = ~n1961 & ~n1963 ;
  assign n1965 = ~n1949 & ~n1959 ;
  assign n1966 = ~n1946 & n1959 ;
  assign n1967 = n1948 & n1966 ;
  assign n1968 = n1954 & ~n1967 ;
  assign n1969 = ~n1965 & n1968 ;
  assign n1970 = n1964 & ~n1969 ;
  assign n1971 = ~n1942 & ~n1970 ;
  assign n1972 = ~n1941 & n1971 ;
  assign n1973 = n468 & n514 ;
  assign n1974 = ~n468 & ~n514 ;
  assign n1975 = ~n1973 & ~n1974 ;
  assign n1976 = n489 & ~n1975 ;
  assign n1977 = ~n489 & n1975 ;
  assign n1978 = ~n1976 & ~n1977 ;
  assign n1979 = ~\173(96)_pad  & ~\174(97)_pad  ;
  assign n1980 = \18(5)_pad  & ~n1979 ;
  assign n1981 = \173(96)_pad  & \174(97)_pad  ;
  assign n1982 = ~n396 & ~n1981 ;
  assign n1983 = n1980 & n1982 ;
  assign n1984 = n461 & n1983 ;
  assign n1985 = ~n461 & ~n1983 ;
  assign n1986 = ~n1984 & ~n1985 ;
  assign n1987 = \18(5)_pad  & \181(104)_pad  ;
  assign n1988 = ~n1612 & ~n1987 ;
  assign n1989 = n521 & n1988 ;
  assign n1990 = ~n521 & ~n1988 ;
  assign n1991 = ~n1989 & ~n1990 ;
  assign n1992 = ~\175(98)_pad  & ~\176(99)_pad  ;
  assign n1993 = \18(5)_pad  & ~n1992 ;
  assign n1994 = \175(98)_pad  & \176(99)_pad  ;
  assign n1995 = ~n396 & ~n1994 ;
  assign n1996 = n1993 & n1995 ;
  assign n1997 = ~n1991 & ~n1996 ;
  assign n1998 = n1986 & n1997 ;
  assign n1999 = ~n1991 & n1996 ;
  assign n2000 = ~n1986 & n1999 ;
  assign n2001 = ~n1998 & ~n2000 ;
  assign n2002 = n1991 & n1996 ;
  assign n2003 = n1986 & n2002 ;
  assign n2004 = n1991 & ~n1996 ;
  assign n2005 = ~n1986 & n2004 ;
  assign n2006 = ~n2003 & ~n2005 ;
  assign n2007 = n2001 & n2006 ;
  assign n2008 = ~n1978 & n2007 ;
  assign n2009 = n1978 & ~n2007 ;
  assign n2010 = ~n2008 & ~n2009 ;
  assign n2011 = n1972 & n2010 ;
  assign n2012 = ~n1896 & n2011 ;
  assign n2013 = ~n1896 & n2010 ;
  assign n2014 = n1462 & n1465 ;
  assign n2015 = n1456 & n2014 ;
  assign n2016 = n1459 & n2015 ;
  assign n2017 = ~n1511 & n2016 ;
  assign n2018 = n1540 & n2017 ;
  assign n2019 = n1636 & n2018 ;
  assign n2020 = n2013 & n2019 ;
  assign n2021 = n1842 & n1972 ;
  assign n2022 = n2020 & n2021 ;
  assign n2023 = ~n1084 & ~n1094 ;
  assign n2024 = ~n813 & ~n2023 ;
  assign n2025 = ~n819 & n2024 ;
  assign n2026 = ~n813 & ~n819 ;
  assign n2027 = n2023 & ~n2026 ;
  assign n2028 = ~n2025 & ~n2027 ;
  assign n2029 = ~n813 & ~n1098 ;
  assign n2030 = ~n819 & n2029 ;
  assign n2031 = ~n1088 & ~n2026 ;
  assign n2032 = ~n2030 & ~n2031 ;
  assign \252(3450)_pad  = ~n395 ;
  assign \258(3122)_pad  = n564 ;
  assign \270(3109)_pad  = n828 ;
  assign \278(536)_pad  = n829 ;
  assign \281(547)_pad  = ~n831 ;
  assign \284(384)_pad  = ~n832 ;
  assign \286(419)_pad  = ~\15(4)_pad  ;
  assign \292(392)_pad  = ~n831 ;
  assign \295(3352)_pad  = ~n837 ;
  assign \298(3387)_pad  = n852 ;
  assign \301(3388)_pad  = ~n863 ;
  assign \304(3390)_pad  = ~n870 ;
  assign \307(3389)_pad  = ~n872 ;
  assign \310(3393)_pad  = n886 ;
  assign \313(3396)_pad  = ~n893 ;
  assign \316(3397)_pad  = n899 ;
  assign \319(3398)_pad  = n904 ;
  assign \321(3715)_pad  = n988 ;
  assign \324(3363)_pad  = ~n996 ;
  assign \327(3408)_pad  = n1000 ;
  assign \330(3411)_pad  = n1011 ;
  assign \333(3416)_pad  = n1021 ;
  assign \336(3412)_pad  = ~n1028 ;
  assign \338(3716)_pad  = n1103 ;
  assign \344(3382)_pad  = n1119 ;
  assign \347(3420)_pad  = n1138 ;
  assign \350(3421)_pad  = ~n1149 ;
  assign \353(3425)_pad  = ~n1158 ;
  assign \356(3424)_pad  = ~n1163 ;
  assign \359(3426)_pad  = n1172 ;
  assign \362(3429)_pad  = ~n1180 ;
  assign \365(3430)_pad  = n1189 ;
  assign \368(3431)_pad  = ~n1194 ;
  assign \370(3718)_pad  = ~n1284 ;
  assign \373(2994)_pad  = n1292 ;
  assign \376(3206)_pad  = ~n1307 ;
  assign \379(3207)_pad  = ~n1320 ;
  assign \382(3148)_pad  = ~n1330 ;
  assign \385(3151)_pad  = ~n1332 ;
  assign \388(3093)_pad  = ~n1347 ;
  assign \391(3094)_pad  = n1352 ;
  assign \394(3095)_pad  = n1354 ;
  assign \397(3097)_pad  = n1364 ;
  assign \399(3717)_pad  = ~n1452 ;
  assign \402(395)_pad  = ~n1453 ;
  assign \404(390)_pad  = ~n1456 ;
  assign \406(388)_pad  = ~n1459 ;
  assign \408(385)_pad  = ~n1462 ;
  assign \410(387)_pad  = ~n1465 ;
  assign \412(3369)_pad  = ~n1637 ;
  assign \414(3338)_pad  = ~n1842 ;
  assign \416(3368)_pad  = ~n2012 ;
  assign \418(3449)_pad  = ~n2022 ;
  assign \419(3444)_pad  = ~n2028 ;
  assign \422(3451)_pad  = ~n2032 ;
endmodule
