module top (\pi000 , \pi001 , \pi002 , \pi003 , \pi004 , \pi005 , \pi006 , \pi007 , \pi008 , \pi009 , \pi010 , \pi011 , \pi012 , \pi013 , \pi014 , \pi015 , \pi016 , \pi017 , \pi018 , \pi019 , \pi020 , \pi021 , \pi022 , \pi023 , \pi024 , \pi025 , \pi026 , \pi027 , \pi028 , \pi029 , \pi030 , \pi031 , \pi032 , \pi033 , \pi034 , \pi035 , \pi036 , \pi037 , \pi038 , \pi039 , \pi040 , \pi041 , \pi042 , \pi043 , \pi044 , \pi045 , \pi046 , \pi047 , \pi048 , \pi049 , \pi050 , \pi051 , \pi052 , \pi053 , \pi054 , \pi055 , \pi056 , \pi057 , \pi058 , \pi059 , \pi060 , \pi061 , \pi062 , \pi063 , \pi064 , \pi065 , \pi066 , \pi067 , \pi068 , \pi069 , \pi070 , \pi071 , \pi072 , \pi073 , \pi074 , \pi075 , \pi076 , \pi077 , \pi078 , \pi079 , \pi080 , \pi081 , \pi082 , \pi083 , \pi084 , \pi085 , \pi086 , \pi087 , \pi088 , \pi089 , \pi090 , \pi091 , \pi092 , \pi093 , \pi094 , \pi095 , \pi096 , \pi097 , \pi098 , \pi099 , \pi100 , \pi101 , \pi102 , \pi103 , \pi104 , \pi105 , \pi106 , \pi107 , \pi108 , \pi109 , \pi110 , \pi111 , \pi112 , \pi113 , \pi114 , \pi115 , \pi116 , \pi117 , \pi118 , \pi119 , \pi120 , \pi121 , \pi122 , \pi123 , \pi124 , \pi125 , \pi126 , \pi127 , \pi128 , \pi129 , \pi130 , \pi131 , \pi132 , \pi133 , \pi134 , \pi135 , \pi136 , \pi137 , \pi138 , \pi139 , \pi140 , \pi141 , \pi142 , \pi143 , \pi144 , \pi145 , \pi146 , \po000 , \po001 , \po002 , \po003 , \po004 , \po005 , \po006 , \po007 , \po008 , \po009 , \po010 , \po011 , \po012 , \po013 , \po014 , \po015 , \po016 , \po017 , \po018 , \po019 , \po020 , \po021 , \po022 , \po023 , \po024 , \po025 , \po026 , \po027 , \po028 , \po029 , \po030 , \po031 , \po032 , \po033 , \po034 , \po035 , \po036 , \po037 , \po038 , \po039 , \po040 , \po041 , \po042 , \po043 , \po044 , \po045 , \po046 , \po047 , \po048 , \po049 , \po050 , \po051 , \po052 , \po053 , \po054 , \po055 , \po056 , \po057 , \po058 , \po059 , \po060 , \po061 , \po062 , \po063 , \po064 , \po065 , \po066 , \po067 , \po068 , \po069 , \po070 , \po071 , \po072 , \po073 , \po074 , \po075 , \po076 , \po077 , \po078 , \po079 , \po080 , \po081 , \po082 , \po083 , \po084 , \po085 , \po086 , \po087 , \po088 , \po089 , \po090 , \po091 , \po092 , \po093 , \po094 , \po095 , \po096 , \po097 , \po098 , \po099 , \po100 , \po101 , \po102 , \po103 , \po104 , \po105 , \po106 , \po107 , \po108 , \po109 , \po110 , \po111 , \po112 , \po113 , \po114 , \po115 , \po116 , \po117 , \po118 , \po119 , \po120 , \po121 , \po122 , \po123 , \po124 , \po125 , \po126 , \po127 , \po128 , \po129 , \po130 , \po131 , \po132 , \po133 , \po134 , \po135 , \po136 , \po137 , \po138 , \po139 , \po140 , \po141 );
	input \pi000  ;
	input \pi001  ;
	input \pi002  ;
	input \pi003  ;
	input \pi004  ;
	input \pi005  ;
	input \pi006  ;
	input \pi007  ;
	input \pi008  ;
	input \pi009  ;
	input \pi010  ;
	input \pi011  ;
	input \pi012  ;
	input \pi013  ;
	input \pi014  ;
	input \pi015  ;
	input \pi016  ;
	input \pi017  ;
	input \pi018  ;
	input \pi019  ;
	input \pi020  ;
	input \pi021  ;
	input \pi022  ;
	input \pi023  ;
	input \pi024  ;
	input \pi025  ;
	input \pi026  ;
	input \pi027  ;
	input \pi028  ;
	input \pi029  ;
	input \pi030  ;
	input \pi031  ;
	input \pi032  ;
	input \pi033  ;
	input \pi034  ;
	input \pi035  ;
	input \pi036  ;
	input \pi037  ;
	input \pi038  ;
	input \pi039  ;
	input \pi040  ;
	input \pi041  ;
	input \pi042  ;
	input \pi043  ;
	input \pi044  ;
	input \pi045  ;
	input \pi046  ;
	input \pi047  ;
	input \pi048  ;
	input \pi049  ;
	input \pi050  ;
	input \pi051  ;
	input \pi052  ;
	input \pi053  ;
	input \pi054  ;
	input \pi055  ;
	input \pi056  ;
	input \pi057  ;
	input \pi058  ;
	input \pi059  ;
	input \pi060  ;
	input \pi061  ;
	input \pi062  ;
	input \pi063  ;
	input \pi064  ;
	input \pi065  ;
	input \pi066  ;
	input \pi067  ;
	input \pi068  ;
	input \pi069  ;
	input \pi070  ;
	input \pi071  ;
	input \pi072  ;
	input \pi073  ;
	input \pi074  ;
	input \pi075  ;
	input \pi076  ;
	input \pi077  ;
	input \pi078  ;
	input \pi079  ;
	input \pi080  ;
	input \pi081  ;
	input \pi082  ;
	input \pi083  ;
	input \pi084  ;
	input \pi085  ;
	input \pi086  ;
	input \pi087  ;
	input \pi088  ;
	input \pi089  ;
	input \pi090  ;
	input \pi091  ;
	input \pi092  ;
	input \pi093  ;
	input \pi094  ;
	input \pi095  ;
	input \pi096  ;
	input \pi097  ;
	input \pi098  ;
	input \pi099  ;
	input \pi100  ;
	input \pi101  ;
	input \pi102  ;
	input \pi103  ;
	input \pi104  ;
	input \pi105  ;
	input \pi106  ;
	input \pi107  ;
	input \pi108  ;
	input \pi109  ;
	input \pi110  ;
	input \pi111  ;
	input \pi112  ;
	input \pi113  ;
	input \pi114  ;
	input \pi115  ;
	input \pi116  ;
	input \pi117  ;
	input \pi118  ;
	input \pi119  ;
	input \pi120  ;
	input \pi121  ;
	input \pi122  ;
	input \pi123  ;
	input \pi124  ;
	input \pi125  ;
	input \pi126  ;
	input \pi127  ;
	input \pi128  ;
	input \pi129  ;
	input \pi130  ;
	input \pi131  ;
	input \pi132  ;
	input \pi133  ;
	input \pi134  ;
	input \pi135  ;
	input \pi136  ;
	input \pi137  ;
	input \pi138  ;
	input \pi139  ;
	input \pi140  ;
	input \pi141  ;
	input \pi142  ;
	input \pi143  ;
	input \pi144  ;
	input \pi145  ;
	input \pi146  ;
	output \po000  ;
	output \po001  ;
	output \po002  ;
	output \po003  ;
	output \po004  ;
	output \po005  ;
	output \po006  ;
	output \po007  ;
	output \po008  ;
	output \po009  ;
	output \po010  ;
	output \po011  ;
	output \po012  ;
	output \po013  ;
	output \po014  ;
	output \po015  ;
	output \po016  ;
	output \po017  ;
	output \po018  ;
	output \po019  ;
	output \po020  ;
	output \po021  ;
	output \po022  ;
	output \po023  ;
	output \po024  ;
	output \po025  ;
	output \po026  ;
	output \po027  ;
	output \po028  ;
	output \po029  ;
	output \po030  ;
	output \po031  ;
	output \po032  ;
	output \po033  ;
	output \po034  ;
	output \po035  ;
	output \po036  ;
	output \po037  ;
	output \po038  ;
	output \po039  ;
	output \po040  ;
	output \po041  ;
	output \po042  ;
	output \po043  ;
	output \po044  ;
	output \po045  ;
	output \po046  ;
	output \po047  ;
	output \po048  ;
	output \po049  ;
	output \po050  ;
	output \po051  ;
	output \po052  ;
	output \po053  ;
	output \po054  ;
	output \po055  ;
	output \po056  ;
	output \po057  ;
	output \po058  ;
	output \po059  ;
	output \po060  ;
	output \po061  ;
	output \po062  ;
	output \po063  ;
	output \po064  ;
	output \po065  ;
	output \po066  ;
	output \po067  ;
	output \po068  ;
	output \po069  ;
	output \po070  ;
	output \po071  ;
	output \po072  ;
	output \po073  ;
	output \po074  ;
	output \po075  ;
	output \po076  ;
	output \po077  ;
	output \po078  ;
	output \po079  ;
	output \po080  ;
	output \po081  ;
	output \po082  ;
	output \po083  ;
	output \po084  ;
	output \po085  ;
	output \po086  ;
	output \po087  ;
	output \po088  ;
	output \po089  ;
	output \po090  ;
	output \po091  ;
	output \po092  ;
	output \po093  ;
	output \po094  ;
	output \po095  ;
	output \po096  ;
	output \po097  ;
	output \po098  ;
	output \po099  ;
	output \po100  ;
	output \po101  ;
	output \po102  ;
	output \po103  ;
	output \po104  ;
	output \po105  ;
	output \po106  ;
	output \po107  ;
	output \po108  ;
	output \po109  ;
	output \po110  ;
	output \po111  ;
	output \po112  ;
	output \po113  ;
	output \po114  ;
	output \po115  ;
	output \po116  ;
	output \po117  ;
	output \po118  ;
	output \po119  ;
	output \po120  ;
	output \po121  ;
	output \po122  ;
	output \po123  ;
	output \po124  ;
	output \po125  ;
	output \po126  ;
	output \po127  ;
	output \po128  ;
	output \po129  ;
	output \po130  ;
	output \po131  ;
	output \po132  ;
	output \po133  ;
	output \po134  ;
	output \po135  ;
	output \po136  ;
	output \po137  ;
	output \po138  ;
	output \po139  ;
	output \po140  ;
	output \po141  ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\pi003 ,
		\pi129 ,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\pi008 ,
		\pi021 ,
		_w149_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\pi011 ,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\pi007 ,
		\pi013 ,
		_w151_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		\pi014 ,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\pi006 ,
		\pi012 ,
		_w153_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\pi004 ,
		\pi019 ,
		_w154_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		\pi016 ,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\pi017 ,
		\pi018 ,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		_w155_,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\pi005 ,
		\pi022 ,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w153_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		_w157_,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		\pi009 ,
		_w150_,
		_w161_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w152_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		_w160_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\pi054 ,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		\pi000 ,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\pi009 ,
		\pi011 ,
		_w166_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		\pi056 ,
		_w158_,
		_w167_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w166_,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\pi056 ,
		_w158_,
		_w169_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		\pi007 ,
		_w149_,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w149_,
		_w151_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w170_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\pi014 ,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		\pi007 ,
		_w149_,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		\pi008 ,
		\pi021 ,
		_w175_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\pi013 ,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		_w174_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		\pi014 ,
		_w171_,
		_w178_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		\pi010 ,
		_w177_,
		_w179_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		_w178_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		_w173_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		\pi010 ,
		\pi014 ,
		_w182_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w171_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w181_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		_w160_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		_w166_,
		_w169_,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name39 (
		_w185_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		\pi054 ,
		_w168_,
		_w188_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		_w187_,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w165_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		_w148_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\pi010 ,
		\pi022 ,
		_w192_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		\pi013 ,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		\pi005 ,
		\pi006 ,
		_w194_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		\pi007 ,
		\pi012 ,
		_w195_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		_w194_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w155_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\pi014 ,
		\pi018 ,
		_w198_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w150_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w193_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w197_,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		\pi017 ,
		\pi054 ,
		_w202_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		_w201_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\pi001 ,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w150_,
		_w157_,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		\pi013 ,
		_w196_,
		_w206_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		\pi009 ,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		_w194_,
		_w195_,
		_w208_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		\pi005 ,
		\pi007 ,
		_w209_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		_w153_,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		\pi009 ,
		_w208_,
		_w211_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		_w210_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		_w206_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		\pi013 ,
		_w196_,
		_w214_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		\pi022 ,
		\pi054 ,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		\pi010 ,
		\pi014 ,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		_w215_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		_w214_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		_w205_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w207_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		_w213_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w204_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h2)
	) name75 (
		_w148_,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		\pi122 ,
		\pi127 ,
		_w224_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		\pi082 ,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		\pi042 ,
		\pi044 ,
		_w226_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		\pi038 ,
		\pi040 ,
		_w227_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		_w226_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		\pi046 ,
		\pi050 ,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		_w228_,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		\pi041 ,
		\pi043 ,
		_w231_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		\pi047 ,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		_w230_,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		\pi048 ,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		\pi002 ,
		\pi020 ,
		_w235_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		\pi015 ,
		\pi049 ,
		_w236_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		_w235_,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		\pi024 ,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		\pi045 ,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		_w224_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		_w234_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w225_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		\pi065 ,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		\pi082 ,
		_w224_,
		_w244_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		\pi045 ,
		_w234_,
		_w245_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		\pi024 ,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w236_,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h4)
	) name100 (
		\pi020 ,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h2)
	) name101 (
		\pi082 ,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w244_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h2)
	) name103 (
		\pi002 ,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		_w243_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		\pi129 ,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h2)
	) name106 (
		\pi000 ,
		\pi113 ,
		_w254_
	);
	LUT2 #(
		.INIT('h4)
	) name107 (
		\pi123 ,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		\pi009 ,
		\pi014 ,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		_w193_,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		_w195_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		_w194_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		_w205_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		\pi061 ,
		\pi118 ,
		_w261_
	);
	LUT2 #(
		.INIT('h4)
	) name114 (
		_w260_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		_w255_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		\pi129 ,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		\pi004 ,
		\pi054 ,
		_w265_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		\pi054 ,
		_w205_,
		_w266_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		\pi022 ,
		_w182_,
		_w267_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		_w207_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		_w266_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w265_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h2)
	) name123 (
		_w148_,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h2)
	) name124 (
		\pi005 ,
		\pi054 ,
		_w272_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		\pi054 ,
		_w196_,
		_w273_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		\pi016 ,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		\pi017 ,
		_w150_,
		_w275_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		_w257_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		\pi059 ,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		\pi018 ,
		_w154_,
		_w278_
	);
	LUT2 #(
		.INIT('h4)
	) name131 (
		\pi029 ,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		\pi025 ,
		\pi028 ,
		_w280_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		_w279_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		_w274_,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		_w277_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		_w272_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h2)
	) name137 (
		_w148_,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h2)
	) name138 (
		\pi006 ,
		\pi054 ,
		_w286_
	);
	LUT2 #(
		.INIT('h2)
	) name139 (
		\pi025 ,
		\pi028 ,
		_w287_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		_w279_,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		_w274_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		_w277_,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		_w286_,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h2)
	) name144 (
		_w148_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h2)
	) name145 (
		\pi007 ,
		\pi054 ,
		_w293_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		\pi054 ,
		_w155_,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w259_,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h4)
	) name148 (
		\pi011 ,
		_w156_,
		_w296_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		_w295_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		\pi008 ,
		\pi021 ,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		_w297_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		_w293_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h2)
	) name153 (
		_w148_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h2)
	) name154 (
		\pi008 ,
		\pi054 ,
		_w302_
	);
	LUT2 #(
		.INIT('h4)
	) name155 (
		\pi008 ,
		\pi021 ,
		_w303_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		_w297_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w302_,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		_w148_,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h2)
	) name159 (
		\pi009 ,
		\pi054 ,
		_w307_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		_w192_,
		_w294_,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		_w149_,
		_w156_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		_w206_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		\pi011 ,
		_w256_,
		_w311_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		_w308_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		_w310_,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w307_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h2)
	) name167 (
		_w148_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h2)
	) name168 (
		\pi010 ,
		\pi054 ,
		_w316_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		\pi009 ,
		_w309_,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		_w308_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h4)
	) name171 (
		\pi011 ,
		\pi014 ,
		_w319_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		_w206_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		_w318_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		_w316_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h2)
	) name175 (
		_w148_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		\pi011 ,
		\pi054 ,
		_w324_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		\pi022 ,
		_w166_,
		_w325_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		_w216_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		_w294_,
		_w326_,
		_w327_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		_w310_,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		_w324_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h2)
	) name182 (
		_w148_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h2)
	) name183 (
		\pi012 ,
		\pi054 ,
		_w331_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		\pi018 ,
		_w275_,
		_w332_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		_w295_,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		_w331_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h2)
	) name187 (
		_w148_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h2)
	) name188 (
		\pi013 ,
		\pi054 ,
		_w336_
	);
	LUT2 #(
		.INIT('h4)
	) name189 (
		\pi018 ,
		_w295_,
		_w337_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		\pi025 ,
		\pi028 ,
		_w338_
	);
	LUT2 #(
		.INIT('h2)
	) name191 (
		\pi029 ,
		\pi059 ,
		_w339_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		_w338_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		_w275_,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		_w337_,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		_w336_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h2)
	) name196 (
		_w148_,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h2)
	) name197 (
		\pi014 ,
		\pi054 ,
		_w345_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		\pi011 ,
		\pi013 ,
		_w346_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w217_,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		_w197_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		_w317_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		_w345_,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h2)
	) name203 (
		_w148_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		\pi015 ,
		_w244_,
		_w352_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		_w235_,
		_w247_,
		_w353_
	);
	LUT2 #(
		.INIT('h4)
	) name206 (
		\pi049 ,
		_w246_,
		_w354_
	);
	LUT2 #(
		.INIT('h2)
	) name207 (
		\pi015 ,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		_w353_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h2)
	) name209 (
		\pi082 ,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h2)
	) name210 (
		\pi082 ,
		_w247_,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		\pi070 ,
		_w224_,
		_w359_
	);
	LUT2 #(
		.INIT('h4)
	) name212 (
		_w358_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w352_,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h4)
	) name214 (
		_w357_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		\pi129 ,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h2)
	) name216 (
		\pi016 ,
		\pi054 ,
		_w364_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		\pi005 ,
		\pi006 ,
		_w365_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		_w258_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		_w266_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		_w364_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		_w148_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		\pi017 ,
		\pi054 ,
		_w370_
	);
	LUT2 #(
		.INIT('h4)
	) name223 (
		\pi029 ,
		\pi054 ,
		_w371_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		\pi059 ,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		_w338_,
		_w372_,
		_w373_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		_w260_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		_w370_,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h2)
	) name228 (
		_w148_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h2)
	) name229 (
		\pi018 ,
		\pi054 ,
		_w377_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w273_,
		_w276_,
		_w378_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		\pi016 ,
		_w278_,
		_w379_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		_w378_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		_w377_,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h2)
	) name234 (
		_w148_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h2)
	) name235 (
		\pi019 ,
		\pi054 ,
		_w383_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		\pi017 ,
		_w150_,
		_w384_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		_w337_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		_w383_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h2)
	) name239 (
		_w148_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		\pi002 ,
		_w248_,
		_w388_
	);
	LUT2 #(
		.INIT('h2)
	) name241 (
		\pi020 ,
		_w247_,
		_w389_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w388_,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h2)
	) name243 (
		\pi082 ,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		\pi020 ,
		_w244_,
		_w392_
	);
	LUT2 #(
		.INIT('h1)
	) name245 (
		\pi071 ,
		_w224_,
		_w393_
	);
	LUT2 #(
		.INIT('h4)
	) name246 (
		_w249_,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		_w392_,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h4)
	) name248 (
		_w391_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name249 (
		\pi129 ,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		\pi021 ,
		\pi054 ,
		_w398_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		\pi004 ,
		\pi016 ,
		_w399_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		\pi018 ,
		\pi019 ,
		_w400_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		_w399_,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		_w378_,
		_w401_,
		_w402_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w398_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h2)
	) name256 (
		_w148_,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h2)
	) name257 (
		\pi022 ,
		\pi054 ,
		_w405_
	);
	LUT2 #(
		.INIT('h2)
	) name258 (
		\pi005 ,
		\pi011 ,
		_w406_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		_w153_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		_w152_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		_w318_,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w405_,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		_w148_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h4)
	) name264 (
		\pi023 ,
		\pi055 ,
		_w412_
	);
	LUT2 #(
		.INIT('h2)
	) name265 (
		\pi061 ,
		\pi129 ,
		_w413_
	);
	LUT2 #(
		.INIT('h4)
	) name266 (
		_w412_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		\pi082 ,
		_w230_,
		_w415_
	);
	LUT2 #(
		.INIT('h2)
	) name268 (
		\pi024 ,
		\pi045 ,
		_w416_
	);
	LUT2 #(
		.INIT('h4)
	) name269 (
		\pi048 ,
		_w416_,
		_w417_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		_w232_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		_w415_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h2)
	) name272 (
		\pi082 ,
		_w245_,
		_w420_
	);
	LUT2 #(
		.INIT('h2)
	) name273 (
		\pi082 ,
		_w237_,
		_w421_
	);
	LUT2 #(
		.INIT('h2)
	) name274 (
		_w224_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h1)
	) name275 (
		_w420_,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		\pi024 ,
		_w423_,
		_w424_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		_w237_,
		_w245_,
		_w425_
	);
	LUT2 #(
		.INIT('h2)
	) name278 (
		\pi082 ,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h2)
	) name279 (
		\pi063 ,
		_w224_,
		_w427_
	);
	LUT2 #(
		.INIT('h4)
	) name280 (
		_w426_,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		\pi129 ,
		_w419_,
		_w429_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		_w424_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		_w428_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		\pi053 ,
		\pi058 ,
		_w432_
	);
	LUT2 #(
		.INIT('h2)
	) name285 (
		\pi025 ,
		\pi116 ,
		_w433_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		\pi026 ,
		\pi027 ,
		_w434_
	);
	LUT2 #(
		.INIT('h4)
	) name287 (
		\pi085 ,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		_w433_,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w432_,
		_w436_,
		_w437_
	);
	LUT2 #(
		.INIT('h4)
	) name290 (
		\pi053 ,
		\pi058 ,
		_w438_
	);
	LUT2 #(
		.INIT('h2)
	) name291 (
		\pi053 ,
		\pi058 ,
		_w439_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w438_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		\pi039 ,
		\pi052 ,
		_w441_
	);
	LUT2 #(
		.INIT('h4)
	) name294 (
		\pi051 ,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h8)
	) name295 (
		\pi116 ,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		_w433_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h2)
	) name297 (
		\pi027 ,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		\pi095 ,
		\pi100 ,
		_w446_
	);
	LUT2 #(
		.INIT('h4)
	) name299 (
		\pi097 ,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		\pi110 ,
		_w447_,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		\pi051 ,
		\pi052 ,
		_w449_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		\pi039 ,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h2)
	) name303 (
		\pi027 ,
		_w450_,
		_w451_
	);
	LUT2 #(
		.INIT('h2)
	) name304 (
		\pi025 ,
		_w448_,
		_w452_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		_w451_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		_w445_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		\pi085 ,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		\pi096 ,
		\pi110 ,
		_w456_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		\pi085 ,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h2)
	) name310 (
		\pi085 ,
		\pi116 ,
		_w458_
	);
	LUT2 #(
		.INIT('h2)
	) name311 (
		\pi100 ,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h4)
	) name312 (
		_w457_,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('h8)
	) name313 (
		\pi025 ,
		_w458_,
		_w461_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		_w460_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		\pi027 ,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		_w455_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		\pi026 ,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h2)
	) name318 (
		\pi026 ,
		\pi085 ,
		_w466_
	);
	LUT2 #(
		.INIT('h4)
	) name319 (
		_w443_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h1)
	) name320 (
		\pi025 ,
		\pi116 ,
		_w468_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		\pi027 ,
		_w468_,
		_w469_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		_w467_,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		_w465_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		\pi053 ,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h2)
	) name325 (
		_w440_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h2)
	) name326 (
		_w148_,
		_w437_,
		_w474_
	);
	LUT2 #(
		.INIT('h4)
	) name327 (
		_w473_,
		_w474_,
		_w475_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		\pi027 ,
		_w432_,
		_w476_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		\pi026 ,
		\pi116 ,
		_w477_
	);
	LUT2 #(
		.INIT('h2)
	) name330 (
		_w460_,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h1)
	) name331 (
		_w467_,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		_w148_,
		_w476_,
		_w480_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		_w479_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h4)
	) name334 (
		\pi026 ,
		_w148_,
		_w482_
	);
	LUT2 #(
		.INIT('h2)
	) name335 (
		\pi027 ,
		\pi085 ,
		_w483_
	);
	LUT2 #(
		.INIT('h4)
	) name336 (
		_w443_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		\pi085 ,
		\pi116 ,
		_w485_
	);
	LUT2 #(
		.INIT('h4)
	) name338 (
		\pi085 ,
		\pi095 ,
		_w486_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		_w456_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		_w485_,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		\pi027 ,
		\pi116 ,
		_w489_
	);
	LUT2 #(
		.INIT('h1)
	) name342 (
		\pi100 ,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('h4)
	) name343 (
		_w488_,
		_w490_,
		_w491_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		_w484_,
		_w491_,
		_w492_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		_w432_,
		_w482_,
		_w493_
	);
	LUT2 #(
		.INIT('h4)
	) name346 (
		_w492_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		\pi028 ,
		\pi116 ,
		_w495_
	);
	LUT2 #(
		.INIT('h8)
	) name348 (
		\pi100 ,
		\pi116 ,
		_w496_
	);
	LUT2 #(
		.INIT('h2)
	) name349 (
		_w434_,
		_w495_,
		_w497_
	);
	LUT2 #(
		.INIT('h4)
	) name350 (
		_w496_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		\pi085 ,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h1)
	) name352 (
		\pi026 ,
		_w450_,
		_w500_
	);
	LUT2 #(
		.INIT('h8)
	) name353 (
		_w489_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h4)
	) name354 (
		\pi027 ,
		_w442_,
		_w502_
	);
	LUT2 #(
		.INIT('h1)
	) name355 (
		_w500_,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w448_,
		_w503_,
		_w504_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		\pi026 ,
		\pi027 ,
		_w505_
	);
	LUT2 #(
		.INIT('h1)
	) name358 (
		_w434_,
		_w505_,
		_w506_
	);
	LUT2 #(
		.INIT('h4)
	) name359 (
		\pi116 ,
		_w506_,
		_w507_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		_w504_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h2)
	) name361 (
		\pi028 ,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h4)
	) name362 (
		\pi026 ,
		\pi095 ,
		_w510_
	);
	LUT2 #(
		.INIT('h4)
	) name363 (
		\pi100 ,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		_w456_,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h8)
	) name365 (
		\pi026 ,
		_w443_,
		_w513_
	);
	LUT2 #(
		.INIT('h1)
	) name366 (
		_w512_,
		_w513_,
		_w514_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		\pi027 ,
		_w514_,
		_w515_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		\pi085 ,
		_w501_,
		_w516_
	);
	LUT2 #(
		.INIT('h4)
	) name369 (
		_w515_,
		_w516_,
		_w517_
	);
	LUT2 #(
		.INIT('h4)
	) name370 (
		_w509_,
		_w517_,
		_w518_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		\pi053 ,
		_w499_,
		_w519_
	);
	LUT2 #(
		.INIT('h4)
	) name372 (
		_w518_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h2)
	) name373 (
		\pi053 ,
		\pi116 ,
		_w521_
	);
	LUT2 #(
		.INIT('h8)
	) name374 (
		\pi028 ,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		_w435_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h1)
	) name376 (
		_w520_,
		_w523_,
		_w524_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		\pi058 ,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h2)
	) name378 (
		\pi058 ,
		\pi116 ,
		_w526_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		\pi026 ,
		\pi053 ,
		_w527_
	);
	LUT2 #(
		.INIT('h4)
	) name380 (
		\pi085 ,
		_w527_,
		_w528_
	);
	LUT2 #(
		.INIT('h4)
	) name381 (
		\pi027 ,
		\pi028 ,
		_w529_
	);
	LUT2 #(
		.INIT('h8)
	) name382 (
		_w526_,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h8)
	) name383 (
		_w528_,
		_w530_,
		_w531_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		_w525_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h2)
	) name385 (
		_w148_,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h2)
	) name386 (
		\pi029 ,
		_w448_,
		_w534_
	);
	LUT2 #(
		.INIT('h8)
	) name387 (
		_w446_,
		_w456_,
		_w535_
	);
	LUT2 #(
		.INIT('h8)
	) name388 (
		\pi097 ,
		_w535_,
		_w536_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		\pi058 ,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h4)
	) name390 (
		_w534_,
		_w537_,
		_w538_
	);
	LUT2 #(
		.INIT('h2)
	) name391 (
		\pi029 ,
		\pi116 ,
		_w539_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		\pi097 ,
		\pi116 ,
		_w540_
	);
	LUT2 #(
		.INIT('h2)
	) name393 (
		\pi058 ,
		_w539_,
		_w541_
	);
	LUT2 #(
		.INIT('h4)
	) name394 (
		_w540_,
		_w541_,
		_w542_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		\pi053 ,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h4)
	) name396 (
		_w538_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h8)
	) name397 (
		_w439_,
		_w539_,
		_w545_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		_w544_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		\pi027 ,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		\pi027 ,
		_w432_,
		_w548_
	);
	LUT2 #(
		.INIT('h8)
	) name401 (
		_w539_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		_w547_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		\pi085 ,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h8)
	) name404 (
		\pi085 ,
		_w539_,
		_w552_
	);
	LUT2 #(
		.INIT('h8)
	) name405 (
		_w476_,
		_w552_,
		_w553_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		_w551_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		\pi026 ,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h8)
	) name408 (
		_w466_,
		_w476_,
		_w556_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		_w539_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		_w555_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h2)
	) name411 (
		_w148_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h4)
	) name412 (
		\pi088 ,
		\pi106 ,
		_w560_
	);
	LUT2 #(
		.INIT('h1)
	) name413 (
		\pi030 ,
		\pi109 ,
		_w561_
	);
	LUT2 #(
		.INIT('h4)
	) name414 (
		\pi060 ,
		\pi109 ,
		_w562_
	);
	LUT2 #(
		.INIT('h1)
	) name415 (
		_w561_,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		\pi106 ,
		_w563_,
		_w564_
	);
	LUT2 #(
		.INIT('h1)
	) name417 (
		\pi129 ,
		_w560_,
		_w565_
	);
	LUT2 #(
		.INIT('h4)
	) name418 (
		_w564_,
		_w565_,
		_w566_
	);
	LUT2 #(
		.INIT('h4)
	) name419 (
		\pi089 ,
		\pi106 ,
		_w567_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		\pi031 ,
		\pi109 ,
		_w568_
	);
	LUT2 #(
		.INIT('h4)
	) name421 (
		\pi030 ,
		\pi109 ,
		_w569_
	);
	LUT2 #(
		.INIT('h1)
	) name422 (
		_w568_,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		\pi106 ,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name424 (
		\pi129 ,
		_w567_,
		_w572_
	);
	LUT2 #(
		.INIT('h4)
	) name425 (
		_w571_,
		_w572_,
		_w573_
	);
	LUT2 #(
		.INIT('h4)
	) name426 (
		\pi099 ,
		\pi106 ,
		_w574_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		\pi032 ,
		\pi109 ,
		_w575_
	);
	LUT2 #(
		.INIT('h4)
	) name428 (
		\pi031 ,
		\pi109 ,
		_w576_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		_w575_,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('h1)
	) name430 (
		\pi106 ,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		\pi129 ,
		_w574_,
		_w579_
	);
	LUT2 #(
		.INIT('h4)
	) name432 (
		_w578_,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h4)
	) name433 (
		\pi090 ,
		\pi106 ,
		_w581_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		\pi033 ,
		\pi109 ,
		_w582_
	);
	LUT2 #(
		.INIT('h4)
	) name435 (
		\pi032 ,
		\pi109 ,
		_w583_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		_w582_,
		_w583_,
		_w584_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		\pi106 ,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h1)
	) name438 (
		\pi129 ,
		_w581_,
		_w586_
	);
	LUT2 #(
		.INIT('h4)
	) name439 (
		_w585_,
		_w586_,
		_w587_
	);
	LUT2 #(
		.INIT('h4)
	) name440 (
		\pi091 ,
		\pi106 ,
		_w588_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		\pi034 ,
		\pi109 ,
		_w589_
	);
	LUT2 #(
		.INIT('h4)
	) name442 (
		\pi033 ,
		\pi109 ,
		_w590_
	);
	LUT2 #(
		.INIT('h1)
	) name443 (
		_w589_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		\pi106 ,
		_w591_,
		_w592_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		\pi129 ,
		_w588_,
		_w593_
	);
	LUT2 #(
		.INIT('h4)
	) name446 (
		_w592_,
		_w593_,
		_w594_
	);
	LUT2 #(
		.INIT('h4)
	) name447 (
		\pi092 ,
		\pi106 ,
		_w595_
	);
	LUT2 #(
		.INIT('h1)
	) name448 (
		\pi035 ,
		\pi109 ,
		_w596_
	);
	LUT2 #(
		.INIT('h4)
	) name449 (
		\pi034 ,
		\pi109 ,
		_w597_
	);
	LUT2 #(
		.INIT('h1)
	) name450 (
		_w596_,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h1)
	) name451 (
		\pi106 ,
		_w598_,
		_w599_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		\pi129 ,
		_w595_,
		_w600_
	);
	LUT2 #(
		.INIT('h4)
	) name453 (
		_w599_,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h4)
	) name454 (
		\pi098 ,
		\pi106 ,
		_w602_
	);
	LUT2 #(
		.INIT('h1)
	) name455 (
		\pi036 ,
		\pi109 ,
		_w603_
	);
	LUT2 #(
		.INIT('h4)
	) name456 (
		\pi035 ,
		\pi109 ,
		_w604_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		_w603_,
		_w604_,
		_w605_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		\pi106 ,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		\pi129 ,
		_w602_,
		_w607_
	);
	LUT2 #(
		.INIT('h4)
	) name460 (
		_w606_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h4)
	) name461 (
		\pi093 ,
		\pi106 ,
		_w609_
	);
	LUT2 #(
		.INIT('h1)
	) name462 (
		\pi037 ,
		\pi109 ,
		_w610_
	);
	LUT2 #(
		.INIT('h4)
	) name463 (
		\pi036 ,
		\pi109 ,
		_w611_
	);
	LUT2 #(
		.INIT('h1)
	) name464 (
		_w610_,
		_w611_,
		_w612_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		\pi106 ,
		_w612_,
		_w613_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		\pi129 ,
		_w609_,
		_w614_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		_w613_,
		_w614_,
		_w615_
	);
	LUT2 #(
		.INIT('h4)
	) name468 (
		\pi044 ,
		\pi082 ,
		_w616_
	);
	LUT2 #(
		.INIT('h4)
	) name469 (
		\pi042 ,
		_w616_,
		_w617_
	);
	LUT2 #(
		.INIT('h4)
	) name470 (
		\pi040 ,
		_w617_,
		_w618_
	);
	LUT2 #(
		.INIT('h2)
	) name471 (
		\pi038 ,
		_w225_,
		_w619_
	);
	LUT2 #(
		.INIT('h4)
	) name472 (
		_w618_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h4)
	) name473 (
		\pi048 ,
		_w239_,
		_w621_
	);
	LUT2 #(
		.INIT('h8)
	) name474 (
		_w232_,
		_w621_,
		_w622_
	);
	LUT2 #(
		.INIT('h8)
	) name475 (
		_w229_,
		_w622_,
		_w623_
	);
	LUT2 #(
		.INIT('h8)
	) name476 (
		\pi082 ,
		_w228_,
		_w624_
	);
	LUT2 #(
		.INIT('h4)
	) name477 (
		_w623_,
		_w624_,
		_w625_
	);
	LUT2 #(
		.INIT('h2)
	) name478 (
		\pi082 ,
		_w228_,
		_w626_
	);
	LUT2 #(
		.INIT('h1)
	) name479 (
		\pi074 ,
		_w224_,
		_w627_
	);
	LUT2 #(
		.INIT('h4)
	) name480 (
		_w626_,
		_w627_,
		_w628_
	);
	LUT2 #(
		.INIT('h1)
	) name481 (
		_w620_,
		_w628_,
		_w629_
	);
	LUT2 #(
		.INIT('h4)
	) name482 (
		_w625_,
		_w629_,
		_w630_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		\pi129 ,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h8)
	) name484 (
		\pi109 ,
		_w449_,
		_w632_
	);
	LUT2 #(
		.INIT('h2)
	) name485 (
		\pi039 ,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h4)
	) name486 (
		\pi051 ,
		\pi109 ,
		_w634_
	);
	LUT2 #(
		.INIT('h8)
	) name487 (
		_w441_,
		_w634_,
		_w635_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		\pi106 ,
		_w635_,
		_w636_
	);
	LUT2 #(
		.INIT('h4)
	) name489 (
		_w633_,
		_w636_,
		_w637_
	);
	LUT2 #(
		.INIT('h1)
	) name490 (
		\pi129 ,
		_w637_,
		_w638_
	);
	LUT2 #(
		.INIT('h2)
	) name491 (
		\pi082 ,
		_w226_,
		_w639_
	);
	LUT2 #(
		.INIT('h4)
	) name492 (
		\pi038 ,
		_w623_,
		_w640_
	);
	LUT2 #(
		.INIT('h2)
	) name493 (
		\pi082 ,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h2)
	) name494 (
		_w224_,
		_w641_,
		_w642_
	);
	LUT2 #(
		.INIT('h1)
	) name495 (
		_w639_,
		_w642_,
		_w643_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		\pi040 ,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h8)
	) name497 (
		\pi040 ,
		_w617_,
		_w645_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		_w226_,
		_w640_,
		_w646_
	);
	LUT2 #(
		.INIT('h2)
	) name499 (
		\pi082 ,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h2)
	) name500 (
		\pi073 ,
		_w224_,
		_w648_
	);
	LUT2 #(
		.INIT('h4)
	) name501 (
		_w647_,
		_w648_,
		_w649_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		\pi129 ,
		_w645_,
		_w650_
	);
	LUT2 #(
		.INIT('h4)
	) name503 (
		_w649_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h4)
	) name504 (
		_w644_,
		_w651_,
		_w652_
	);
	LUT2 #(
		.INIT('h4)
	) name505 (
		\pi047 ,
		_w621_,
		_w653_
	);
	LUT2 #(
		.INIT('h4)
	) name506 (
		\pi043 ,
		_w653_,
		_w654_
	);
	LUT2 #(
		.INIT('h4)
	) name507 (
		\pi041 ,
		_w230_,
		_w655_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		\pi082 ,
		_w655_,
		_w656_
	);
	LUT2 #(
		.INIT('h4)
	) name509 (
		_w654_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h2)
	) name510 (
		\pi041 ,
		_w225_,
		_w658_
	);
	LUT2 #(
		.INIT('h4)
	) name511 (
		_w415_,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h2)
	) name512 (
		\pi082 ,
		_w655_,
		_w660_
	);
	LUT2 #(
		.INIT('h1)
	) name513 (
		\pi076 ,
		_w224_,
		_w661_
	);
	LUT2 #(
		.INIT('h4)
	) name514 (
		_w660_,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h1)
	) name515 (
		_w659_,
		_w662_,
		_w663_
	);
	LUT2 #(
		.INIT('h4)
	) name516 (
		_w657_,
		_w663_,
		_w664_
	);
	LUT2 #(
		.INIT('h1)
	) name517 (
		\pi129 ,
		_w664_,
		_w665_
	);
	LUT2 #(
		.INIT('h8)
	) name518 (
		_w227_,
		_w623_,
		_w666_
	);
	LUT2 #(
		.INIT('h2)
	) name519 (
		\pi082 ,
		_w666_,
		_w667_
	);
	LUT2 #(
		.INIT('h1)
	) name520 (
		\pi072 ,
		_w224_,
		_w668_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		_w667_,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h1)
	) name522 (
		_w639_,
		_w669_,
		_w670_
	);
	LUT2 #(
		.INIT('h2)
	) name523 (
		\pi042 ,
		_w616_,
		_w671_
	);
	LUT2 #(
		.INIT('h4)
	) name524 (
		_w225_,
		_w671_,
		_w672_
	);
	LUT2 #(
		.INIT('h1)
	) name525 (
		_w670_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		\pi129 ,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h2)
	) name527 (
		\pi043 ,
		_w225_,
		_w675_
	);
	LUT2 #(
		.INIT('h4)
	) name528 (
		_w656_,
		_w675_,
		_w676_
	);
	LUT2 #(
		.INIT('h8)
	) name529 (
		_w230_,
		_w231_,
		_w677_
	);
	LUT2 #(
		.INIT('h2)
	) name530 (
		\pi082 ,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		\pi077 ,
		_w224_,
		_w679_
	);
	LUT2 #(
		.INIT('h4)
	) name532 (
		_w678_,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h8)
	) name533 (
		\pi082 ,
		_w677_,
		_w681_
	);
	LUT2 #(
		.INIT('h4)
	) name534 (
		_w653_,
		_w681_,
		_w682_
	);
	LUT2 #(
		.INIT('h1)
	) name535 (
		_w676_,
		_w680_,
		_w683_
	);
	LUT2 #(
		.INIT('h4)
	) name536 (
		_w682_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		\pi129 ,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h8)
	) name538 (
		\pi044 ,
		\pi082 ,
		_w686_
	);
	LUT2 #(
		.INIT('h4)
	) name539 (
		\pi042 ,
		_w666_,
		_w687_
	);
	LUT2 #(
		.INIT('h2)
	) name540 (
		\pi082 ,
		_w687_,
		_w688_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		\pi067 ,
		_w224_,
		_w689_
	);
	LUT2 #(
		.INIT('h8)
	) name542 (
		\pi044 ,
		_w224_,
		_w690_
	);
	LUT2 #(
		.INIT('h1)
	) name543 (
		_w689_,
		_w690_,
		_w691_
	);
	LUT2 #(
		.INIT('h4)
	) name544 (
		_w688_,
		_w691_,
		_w692_
	);
	LUT2 #(
		.INIT('h1)
	) name545 (
		\pi129 ,
		_w686_,
		_w693_
	);
	LUT2 #(
		.INIT('h4)
	) name546 (
		_w692_,
		_w693_,
		_w694_
	);
	LUT2 #(
		.INIT('h2)
	) name547 (
		\pi082 ,
		_w234_,
		_w695_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		_w244_,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h2)
	) name549 (
		\pi045 ,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h2)
	) name550 (
		\pi082 ,
		_w238_,
		_w698_
	);
	LUT2 #(
		.INIT('h1)
	) name551 (
		\pi068 ,
		_w224_,
		_w699_
	);
	LUT2 #(
		.INIT('h1)
	) name552 (
		_w698_,
		_w699_,
		_w700_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		_w420_,
		_w700_,
		_w701_
	);
	LUT2 #(
		.INIT('h1)
	) name554 (
		_w697_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		\pi129 ,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h4)
	) name556 (
		\pi075 ,
		_w225_,
		_w704_
	);
	LUT2 #(
		.INIT('h1)
	) name557 (
		\pi075 ,
		_w224_,
		_w705_
	);
	LUT2 #(
		.INIT('h2)
	) name558 (
		\pi082 ,
		_w622_,
		_w706_
	);
	LUT2 #(
		.INIT('h1)
	) name559 (
		_w705_,
		_w706_,
		_w707_
	);
	LUT2 #(
		.INIT('h2)
	) name560 (
		_w230_,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h4)
	) name561 (
		\pi050 ,
		_w624_,
		_w709_
	);
	LUT2 #(
		.INIT('h2)
	) name562 (
		\pi046 ,
		_w225_,
		_w710_
	);
	LUT2 #(
		.INIT('h4)
	) name563 (
		_w709_,
		_w710_,
		_w711_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w704_,
		_w711_,
		_w712_
	);
	LUT2 #(
		.INIT('h4)
	) name565 (
		_w708_,
		_w712_,
		_w713_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		\pi129 ,
		_w713_,
		_w714_
	);
	LUT2 #(
		.INIT('h2)
	) name567 (
		\pi082 ,
		_w621_,
		_w715_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		\pi064 ,
		_w224_,
		_w716_
	);
	LUT2 #(
		.INIT('h1)
	) name569 (
		_w715_,
		_w716_,
		_w717_
	);
	LUT2 #(
		.INIT('h2)
	) name570 (
		\pi082 ,
		_w233_,
		_w718_
	);
	LUT2 #(
		.INIT('h1)
	) name571 (
		_w717_,
		_w718_,
		_w719_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		_w244_,
		_w678_,
		_w720_
	);
	LUT2 #(
		.INIT('h2)
	) name573 (
		\pi047 ,
		_w720_,
		_w721_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		_w719_,
		_w721_,
		_w722_
	);
	LUT2 #(
		.INIT('h1)
	) name575 (
		\pi129 ,
		_w722_,
		_w723_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		_w244_,
		_w718_,
		_w724_
	);
	LUT2 #(
		.INIT('h2)
	) name577 (
		\pi048 ,
		_w724_,
		_w725_
	);
	LUT2 #(
		.INIT('h2)
	) name578 (
		\pi082 ,
		_w239_,
		_w726_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		\pi062 ,
		_w224_,
		_w727_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		_w726_,
		_w727_,
		_w728_
	);
	LUT2 #(
		.INIT('h1)
	) name581 (
		_w695_,
		_w728_,
		_w729_
	);
	LUT2 #(
		.INIT('h1)
	) name582 (
		_w725_,
		_w729_,
		_w730_
	);
	LUT2 #(
		.INIT('h1)
	) name583 (
		\pi129 ,
		_w730_,
		_w731_
	);
	LUT2 #(
		.INIT('h4)
	) name584 (
		_w246_,
		_w421_,
		_w732_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		_w244_,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h2)
	) name586 (
		\pi049 ,
		_w733_,
		_w734_
	);
	LUT2 #(
		.INIT('h2)
	) name587 (
		\pi069 ,
		_w421_,
		_w735_
	);
	LUT2 #(
		.INIT('h2)
	) name588 (
		\pi082 ,
		_w354_,
		_w736_
	);
	LUT2 #(
		.INIT('h1)
	) name589 (
		_w422_,
		_w735_,
		_w737_
	);
	LUT2 #(
		.INIT('h4)
	) name590 (
		_w736_,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h1)
	) name591 (
		_w734_,
		_w738_,
		_w739_
	);
	LUT2 #(
		.INIT('h1)
	) name592 (
		\pi129 ,
		_w739_,
		_w740_
	);
	LUT2 #(
		.INIT('h4)
	) name593 (
		\pi046 ,
		_w622_,
		_w741_
	);
	LUT2 #(
		.INIT('h2)
	) name594 (
		\pi082 ,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h2)
	) name595 (
		_w224_,
		_w742_,
		_w743_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		_w626_,
		_w743_,
		_w744_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		\pi050 ,
		_w744_,
		_w745_
	);
	LUT2 #(
		.INIT('h8)
	) name598 (
		\pi050 ,
		_w624_,
		_w746_
	);
	LUT2 #(
		.INIT('h8)
	) name599 (
		_w228_,
		_w741_,
		_w747_
	);
	LUT2 #(
		.INIT('h2)
	) name600 (
		\pi082 ,
		_w747_,
		_w748_
	);
	LUT2 #(
		.INIT('h2)
	) name601 (
		\pi066 ,
		_w224_,
		_w749_
	);
	LUT2 #(
		.INIT('h4)
	) name602 (
		_w748_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		\pi129 ,
		_w746_,
		_w751_
	);
	LUT2 #(
		.INIT('h4)
	) name604 (
		_w750_,
		_w751_,
		_w752_
	);
	LUT2 #(
		.INIT('h4)
	) name605 (
		_w745_,
		_w752_,
		_w753_
	);
	LUT2 #(
		.INIT('h2)
	) name606 (
		\pi051 ,
		\pi109 ,
		_w754_
	);
	LUT2 #(
		.INIT('h1)
	) name607 (
		\pi106 ,
		_w634_,
		_w755_
	);
	LUT2 #(
		.INIT('h4)
	) name608 (
		_w754_,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h1)
	) name609 (
		\pi129 ,
		_w756_,
		_w757_
	);
	LUT2 #(
		.INIT('h2)
	) name610 (
		\pi052 ,
		_w634_,
		_w758_
	);
	LUT2 #(
		.INIT('h1)
	) name611 (
		\pi106 ,
		_w632_,
		_w759_
	);
	LUT2 #(
		.INIT('h4)
	) name612 (
		_w758_,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h1)
	) name613 (
		\pi129 ,
		_w760_,
		_w761_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		\pi058 ,
		_w535_,
		_w762_
	);
	LUT2 #(
		.INIT('h4)
	) name615 (
		\pi053 ,
		\pi097 ,
		_w763_
	);
	LUT2 #(
		.INIT('h4)
	) name616 (
		_w762_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('h1)
	) name617 (
		_w521_,
		_w764_,
		_w765_
	);
	LUT2 #(
		.INIT('h2)
	) name618 (
		_w148_,
		_w526_,
		_w766_
	);
	LUT2 #(
		.INIT('h8)
	) name619 (
		_w435_,
		_w766_,
		_w767_
	);
	LUT2 #(
		.INIT('h4)
	) name620 (
		_w765_,
		_w767_,
		_w768_
	);
	LUT2 #(
		.INIT('h4)
	) name621 (
		\pi129 ,
		_w242_,
		_w769_
	);
	LUT2 #(
		.INIT('h1)
	) name622 (
		\pi123 ,
		\pi129 ,
		_w770_
	);
	LUT2 #(
		.INIT('h2)
	) name623 (
		\pi114 ,
		\pi122 ,
		_w771_
	);
	LUT2 #(
		.INIT('h8)
	) name624 (
		_w770_,
		_w771_,
		_w772_
	);
	LUT2 #(
		.INIT('h4)
	) name625 (
		\pi026 ,
		\pi037 ,
		_w773_
	);
	LUT2 #(
		.INIT('h4)
	) name626 (
		\pi058 ,
		_w773_,
		_w774_
	);
	LUT2 #(
		.INIT('h4)
	) name627 (
		\pi026 ,
		\pi058 ,
		_w775_
	);
	LUT2 #(
		.INIT('h4)
	) name628 (
		\pi058 ,
		_w477_,
		_w776_
	);
	LUT2 #(
		.INIT('h1)
	) name629 (
		_w775_,
		_w776_,
		_w777_
	);
	LUT2 #(
		.INIT('h2)
	) name630 (
		\pi094 ,
		_w777_,
		_w778_
	);
	LUT2 #(
		.INIT('h2)
	) name631 (
		\pi037 ,
		\pi116 ,
		_w779_
	);
	LUT2 #(
		.INIT('h1)
	) name632 (
		_w775_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h1)
	) name633 (
		_w526_,
		_w780_,
		_w781_
	);
	LUT2 #(
		.INIT('h1)
	) name634 (
		_w778_,
		_w781_,
		_w782_
	);
	LUT2 #(
		.INIT('h1)
	) name635 (
		\pi053 ,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		_w774_,
		_w783_,
		_w784_
	);
	LUT2 #(
		.INIT('h1)
	) name637 (
		\pi053 ,
		\pi085 ,
		_w785_
	);
	LUT2 #(
		.INIT('h8)
	) name638 (
		_w774_,
		_w785_,
		_w786_
	);
	LUT2 #(
		.INIT('h2)
	) name639 (
		\pi027 ,
		_w786_,
		_w787_
	);
	LUT2 #(
		.INIT('h4)
	) name640 (
		\pi053 ,
		_w774_,
		_w788_
	);
	LUT2 #(
		.INIT('h2)
	) name641 (
		\pi085 ,
		_w788_,
		_w789_
	);
	LUT2 #(
		.INIT('h2)
	) name642 (
		_w148_,
		_w787_,
		_w790_
	);
	LUT2 #(
		.INIT('h4)
	) name643 (
		_w789_,
		_w790_,
		_w791_
	);
	LUT2 #(
		.INIT('h4)
	) name644 (
		_w784_,
		_w791_,
		_w792_
	);
	LUT2 #(
		.INIT('h4)
	) name645 (
		\pi116 ,
		_w528_,
		_w793_
	);
	LUT2 #(
		.INIT('h2)
	) name646 (
		\pi085 ,
		_w527_,
		_w794_
	);
	LUT2 #(
		.INIT('h8)
	) name647 (
		\pi026 ,
		\pi053 ,
		_w795_
	);
	LUT2 #(
		.INIT('h1)
	) name648 (
		\pi058 ,
		_w795_,
		_w796_
	);
	LUT2 #(
		.INIT('h4)
	) name649 (
		_w794_,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('h1)
	) name650 (
		_w793_,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('h2)
	) name651 (
		\pi057 ,
		_w798_,
		_w799_
	);
	LUT2 #(
		.INIT('h8)
	) name652 (
		\pi058 ,
		\pi060 ,
		_w800_
	);
	LUT2 #(
		.INIT('h8)
	) name653 (
		\pi116 ,
		_w800_,
		_w801_
	);
	LUT2 #(
		.INIT('h8)
	) name654 (
		_w528_,
		_w801_,
		_w802_
	);
	LUT2 #(
		.INIT('h1)
	) name655 (
		_w799_,
		_w802_,
		_w803_
	);
	LUT2 #(
		.INIT('h1)
	) name656 (
		\pi027 ,
		_w803_,
		_w804_
	);
	LUT2 #(
		.INIT('h2)
	) name657 (
		\pi057 ,
		\pi058 ,
		_w805_
	);
	LUT2 #(
		.INIT('h8)
	) name658 (
		_w528_,
		_w805_,
		_w806_
	);
	LUT2 #(
		.INIT('h1)
	) name659 (
		_w804_,
		_w806_,
		_w807_
	);
	LUT2 #(
		.INIT('h2)
	) name660 (
		_w148_,
		_w807_,
		_w808_
	);
	LUT2 #(
		.INIT('h8)
	) name661 (
		_w434_,
		_w526_,
		_w809_
	);
	LUT2 #(
		.INIT('h4)
	) name662 (
		\pi058 ,
		_w506_,
		_w810_
	);
	LUT2 #(
		.INIT('h8)
	) name663 (
		_w443_,
		_w810_,
		_w811_
	);
	LUT2 #(
		.INIT('h1)
	) name664 (
		_w809_,
		_w811_,
		_w812_
	);
	LUT2 #(
		.INIT('h8)
	) name665 (
		_w148_,
		_w785_,
		_w813_
	);
	LUT2 #(
		.INIT('h4)
	) name666 (
		_w812_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h2)
	) name667 (
		\pi059 ,
		\pi116 ,
		_w815_
	);
	LUT2 #(
		.INIT('h4)
	) name668 (
		_w440_,
		_w815_,
		_w816_
	);
	LUT2 #(
		.INIT('h1)
	) name669 (
		\pi059 ,
		_w448_,
		_w817_
	);
	LUT2 #(
		.INIT('h4)
	) name670 (
		\pi096 ,
		_w448_,
		_w818_
	);
	LUT2 #(
		.INIT('h2)
	) name671 (
		_w432_,
		_w817_,
		_w819_
	);
	LUT2 #(
		.INIT('h4)
	) name672 (
		_w818_,
		_w819_,
		_w820_
	);
	LUT2 #(
		.INIT('h1)
	) name673 (
		_w816_,
		_w820_,
		_w821_
	);
	LUT2 #(
		.INIT('h1)
	) name674 (
		\pi085 ,
		_w821_,
		_w822_
	);
	LUT2 #(
		.INIT('h8)
	) name675 (
		\pi085 ,
		_w432_,
		_w823_
	);
	LUT2 #(
		.INIT('h8)
	) name676 (
		_w815_,
		_w823_,
		_w824_
	);
	LUT2 #(
		.INIT('h1)
	) name677 (
		_w822_,
		_w824_,
		_w825_
	);
	LUT2 #(
		.INIT('h1)
	) name678 (
		\pi027 ,
		_w825_,
		_w826_
	);
	LUT2 #(
		.INIT('h4)
	) name679 (
		\pi085 ,
		_w815_,
		_w827_
	);
	LUT2 #(
		.INIT('h8)
	) name680 (
		_w548_,
		_w827_,
		_w828_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		_w826_,
		_w828_,
		_w829_
	);
	LUT2 #(
		.INIT('h1)
	) name682 (
		\pi026 ,
		_w829_,
		_w830_
	);
	LUT2 #(
		.INIT('h8)
	) name683 (
		_w556_,
		_w815_,
		_w831_
	);
	LUT2 #(
		.INIT('h1)
	) name684 (
		_w830_,
		_w831_,
		_w832_
	);
	LUT2 #(
		.INIT('h2)
	) name685 (
		_w148_,
		_w832_,
		_w833_
	);
	LUT2 #(
		.INIT('h1)
	) name686 (
		\pi117 ,
		\pi122 ,
		_w834_
	);
	LUT2 #(
		.INIT('h2)
	) name687 (
		\pi060 ,
		_w834_,
		_w835_
	);
	LUT2 #(
		.INIT('h8)
	) name688 (
		\pi123 ,
		_w834_,
		_w836_
	);
	LUT2 #(
		.INIT('h1)
	) name689 (
		_w835_,
		_w836_,
		_w837_
	);
	LUT2 #(
		.INIT('h1)
	) name690 (
		\pi114 ,
		\pi122 ,
		_w838_
	);
	LUT2 #(
		.INIT('h2)
	) name691 (
		\pi123 ,
		\pi129 ,
		_w839_
	);
	LUT2 #(
		.INIT('h8)
	) name692 (
		_w838_,
		_w839_,
		_w840_
	);
	LUT2 #(
		.INIT('h2)
	) name693 (
		\pi136 ,
		\pi137 ,
		_w841_
	);
	LUT2 #(
		.INIT('h8)
	) name694 (
		\pi131 ,
		\pi132 ,
		_w842_
	);
	LUT2 #(
		.INIT('h8)
	) name695 (
		\pi133 ,
		_w842_,
		_w843_
	);
	LUT2 #(
		.INIT('h4)
	) name696 (
		\pi138 ,
		_w843_,
		_w844_
	);
	LUT2 #(
		.INIT('h8)
	) name697 (
		_w841_,
		_w844_,
		_w845_
	);
	LUT2 #(
		.INIT('h1)
	) name698 (
		\pi062 ,
		_w845_,
		_w846_
	);
	LUT2 #(
		.INIT('h8)
	) name699 (
		\pi140 ,
		_w845_,
		_w847_
	);
	LUT2 #(
		.INIT('h1)
	) name700 (
		\pi129 ,
		_w846_,
		_w848_
	);
	LUT2 #(
		.INIT('h4)
	) name701 (
		_w847_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h1)
	) name702 (
		\pi063 ,
		_w845_,
		_w850_
	);
	LUT2 #(
		.INIT('h8)
	) name703 (
		\pi142 ,
		_w845_,
		_w851_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		\pi129 ,
		_w850_,
		_w852_
	);
	LUT2 #(
		.INIT('h4)
	) name705 (
		_w851_,
		_w852_,
		_w853_
	);
	LUT2 #(
		.INIT('h1)
	) name706 (
		\pi064 ,
		_w845_,
		_w854_
	);
	LUT2 #(
		.INIT('h8)
	) name707 (
		\pi139 ,
		_w845_,
		_w855_
	);
	LUT2 #(
		.INIT('h1)
	) name708 (
		\pi129 ,
		_w854_,
		_w856_
	);
	LUT2 #(
		.INIT('h4)
	) name709 (
		_w855_,
		_w856_,
		_w857_
	);
	LUT2 #(
		.INIT('h1)
	) name710 (
		\pi065 ,
		_w845_,
		_w858_
	);
	LUT2 #(
		.INIT('h8)
	) name711 (
		\pi146 ,
		_w845_,
		_w859_
	);
	LUT2 #(
		.INIT('h1)
	) name712 (
		\pi129 ,
		_w858_,
		_w860_
	);
	LUT2 #(
		.INIT('h4)
	) name713 (
		_w859_,
		_w860_,
		_w861_
	);
	LUT2 #(
		.INIT('h1)
	) name714 (
		\pi136 ,
		\pi137 ,
		_w862_
	);
	LUT2 #(
		.INIT('h8)
	) name715 (
		_w844_,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h1)
	) name716 (
		\pi066 ,
		_w863_,
		_w864_
	);
	LUT2 #(
		.INIT('h8)
	) name717 (
		\pi143 ,
		_w863_,
		_w865_
	);
	LUT2 #(
		.INIT('h1)
	) name718 (
		\pi129 ,
		_w864_,
		_w866_
	);
	LUT2 #(
		.INIT('h4)
	) name719 (
		_w865_,
		_w866_,
		_w867_
	);
	LUT2 #(
		.INIT('h1)
	) name720 (
		\pi067 ,
		_w863_,
		_w868_
	);
	LUT2 #(
		.INIT('h8)
	) name721 (
		\pi139 ,
		_w863_,
		_w869_
	);
	LUT2 #(
		.INIT('h1)
	) name722 (
		\pi129 ,
		_w868_,
		_w870_
	);
	LUT2 #(
		.INIT('h4)
	) name723 (
		_w869_,
		_w870_,
		_w871_
	);
	LUT2 #(
		.INIT('h1)
	) name724 (
		\pi068 ,
		_w845_,
		_w872_
	);
	LUT2 #(
		.INIT('h8)
	) name725 (
		\pi141 ,
		_w845_,
		_w873_
	);
	LUT2 #(
		.INIT('h1)
	) name726 (
		\pi129 ,
		_w872_,
		_w874_
	);
	LUT2 #(
		.INIT('h4)
	) name727 (
		_w873_,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h1)
	) name728 (
		\pi069 ,
		_w845_,
		_w876_
	);
	LUT2 #(
		.INIT('h8)
	) name729 (
		\pi143 ,
		_w845_,
		_w877_
	);
	LUT2 #(
		.INIT('h1)
	) name730 (
		\pi129 ,
		_w876_,
		_w878_
	);
	LUT2 #(
		.INIT('h4)
	) name731 (
		_w877_,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('h1)
	) name732 (
		\pi070 ,
		_w845_,
		_w880_
	);
	LUT2 #(
		.INIT('h8)
	) name733 (
		\pi144 ,
		_w845_,
		_w881_
	);
	LUT2 #(
		.INIT('h1)
	) name734 (
		\pi129 ,
		_w880_,
		_w882_
	);
	LUT2 #(
		.INIT('h4)
	) name735 (
		_w881_,
		_w882_,
		_w883_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		\pi071 ,
		_w845_,
		_w884_
	);
	LUT2 #(
		.INIT('h8)
	) name737 (
		\pi145 ,
		_w845_,
		_w885_
	);
	LUT2 #(
		.INIT('h1)
	) name738 (
		\pi129 ,
		_w884_,
		_w886_
	);
	LUT2 #(
		.INIT('h4)
	) name739 (
		_w885_,
		_w886_,
		_w887_
	);
	LUT2 #(
		.INIT('h1)
	) name740 (
		\pi072 ,
		_w863_,
		_w888_
	);
	LUT2 #(
		.INIT('h8)
	) name741 (
		\pi140 ,
		_w863_,
		_w889_
	);
	LUT2 #(
		.INIT('h1)
	) name742 (
		\pi129 ,
		_w888_,
		_w890_
	);
	LUT2 #(
		.INIT('h4)
	) name743 (
		_w889_,
		_w890_,
		_w891_
	);
	LUT2 #(
		.INIT('h1)
	) name744 (
		\pi073 ,
		_w863_,
		_w892_
	);
	LUT2 #(
		.INIT('h8)
	) name745 (
		\pi141 ,
		_w863_,
		_w893_
	);
	LUT2 #(
		.INIT('h1)
	) name746 (
		\pi129 ,
		_w892_,
		_w894_
	);
	LUT2 #(
		.INIT('h4)
	) name747 (
		_w893_,
		_w894_,
		_w895_
	);
	LUT2 #(
		.INIT('h1)
	) name748 (
		\pi074 ,
		_w863_,
		_w896_
	);
	LUT2 #(
		.INIT('h8)
	) name749 (
		\pi142 ,
		_w863_,
		_w897_
	);
	LUT2 #(
		.INIT('h1)
	) name750 (
		\pi129 ,
		_w896_,
		_w898_
	);
	LUT2 #(
		.INIT('h4)
	) name751 (
		_w897_,
		_w898_,
		_w899_
	);
	LUT2 #(
		.INIT('h1)
	) name752 (
		\pi075 ,
		_w863_,
		_w900_
	);
	LUT2 #(
		.INIT('h8)
	) name753 (
		\pi144 ,
		_w863_,
		_w901_
	);
	LUT2 #(
		.INIT('h1)
	) name754 (
		\pi129 ,
		_w900_,
		_w902_
	);
	LUT2 #(
		.INIT('h4)
	) name755 (
		_w901_,
		_w902_,
		_w903_
	);
	LUT2 #(
		.INIT('h1)
	) name756 (
		\pi076 ,
		_w863_,
		_w904_
	);
	LUT2 #(
		.INIT('h8)
	) name757 (
		\pi145 ,
		_w863_,
		_w905_
	);
	LUT2 #(
		.INIT('h1)
	) name758 (
		\pi129 ,
		_w904_,
		_w906_
	);
	LUT2 #(
		.INIT('h4)
	) name759 (
		_w905_,
		_w906_,
		_w907_
	);
	LUT2 #(
		.INIT('h1)
	) name760 (
		\pi077 ,
		_w863_,
		_w908_
	);
	LUT2 #(
		.INIT('h8)
	) name761 (
		\pi146 ,
		_w863_,
		_w909_
	);
	LUT2 #(
		.INIT('h1)
	) name762 (
		\pi129 ,
		_w908_,
		_w910_
	);
	LUT2 #(
		.INIT('h4)
	) name763 (
		_w909_,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h4)
	) name764 (
		\pi136 ,
		\pi137 ,
		_w912_
	);
	LUT2 #(
		.INIT('h8)
	) name765 (
		_w844_,
		_w912_,
		_w913_
	);
	LUT2 #(
		.INIT('h1)
	) name766 (
		\pi078 ,
		_w913_,
		_w914_
	);
	LUT2 #(
		.INIT('h4)
	) name767 (
		\pi142 ,
		_w913_,
		_w915_
	);
	LUT2 #(
		.INIT('h1)
	) name768 (
		\pi129 ,
		_w914_,
		_w916_
	);
	LUT2 #(
		.INIT('h4)
	) name769 (
		_w915_,
		_w916_,
		_w917_
	);
	LUT2 #(
		.INIT('h1)
	) name770 (
		\pi079 ,
		_w913_,
		_w918_
	);
	LUT2 #(
		.INIT('h4)
	) name771 (
		\pi143 ,
		_w913_,
		_w919_
	);
	LUT2 #(
		.INIT('h1)
	) name772 (
		\pi129 ,
		_w918_,
		_w920_
	);
	LUT2 #(
		.INIT('h4)
	) name773 (
		_w919_,
		_w920_,
		_w921_
	);
	LUT2 #(
		.INIT('h1)
	) name774 (
		\pi080 ,
		_w913_,
		_w922_
	);
	LUT2 #(
		.INIT('h4)
	) name775 (
		\pi144 ,
		_w913_,
		_w923_
	);
	LUT2 #(
		.INIT('h1)
	) name776 (
		\pi129 ,
		_w922_,
		_w924_
	);
	LUT2 #(
		.INIT('h4)
	) name777 (
		_w923_,
		_w924_,
		_w925_
	);
	LUT2 #(
		.INIT('h1)
	) name778 (
		\pi081 ,
		_w913_,
		_w926_
	);
	LUT2 #(
		.INIT('h4)
	) name779 (
		\pi145 ,
		_w913_,
		_w927_
	);
	LUT2 #(
		.INIT('h1)
	) name780 (
		\pi129 ,
		_w926_,
		_w928_
	);
	LUT2 #(
		.INIT('h4)
	) name781 (
		_w927_,
		_w928_,
		_w929_
	);
	LUT2 #(
		.INIT('h1)
	) name782 (
		\pi082 ,
		_w913_,
		_w930_
	);
	LUT2 #(
		.INIT('h4)
	) name783 (
		\pi146 ,
		_w913_,
		_w931_
	);
	LUT2 #(
		.INIT('h1)
	) name784 (
		\pi129 ,
		_w930_,
		_w932_
	);
	LUT2 #(
		.INIT('h4)
	) name785 (
		_w931_,
		_w932_,
		_w933_
	);
	LUT2 #(
		.INIT('h2)
	) name786 (
		\pi136 ,
		\pi138 ,
		_w934_
	);
	LUT2 #(
		.INIT('h8)
	) name787 (
		\pi031 ,
		_w934_,
		_w935_
	);
	LUT2 #(
		.INIT('h1)
	) name788 (
		\pi087 ,
		\pi138 ,
		_w936_
	);
	LUT2 #(
		.INIT('h8)
	) name789 (
		\pi115 ,
		\pi138 ,
		_w937_
	);
	LUT2 #(
		.INIT('h1)
	) name790 (
		\pi136 ,
		_w936_,
		_w938_
	);
	LUT2 #(
		.INIT('h4)
	) name791 (
		_w937_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h1)
	) name792 (
		_w935_,
		_w939_,
		_w940_
	);
	LUT2 #(
		.INIT('h2)
	) name793 (
		\pi137 ,
		_w940_,
		_w941_
	);
	LUT2 #(
		.INIT('h4)
	) name794 (
		\pi089 ,
		\pi138 ,
		_w942_
	);
	LUT2 #(
		.INIT('h2)
	) name795 (
		\pi062 ,
		\pi138 ,
		_w943_
	);
	LUT2 #(
		.INIT('h2)
	) name796 (
		\pi136 ,
		_w942_,
		_w944_
	);
	LUT2 #(
		.INIT('h4)
	) name797 (
		_w943_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h4)
	) name798 (
		\pi119 ,
		\pi138 ,
		_w946_
	);
	LUT2 #(
		.INIT('h2)
	) name799 (
		\pi072 ,
		\pi138 ,
		_w947_
	);
	LUT2 #(
		.INIT('h1)
	) name800 (
		\pi136 ,
		_w946_,
		_w948_
	);
	LUT2 #(
		.INIT('h4)
	) name801 (
		_w947_,
		_w948_,
		_w949_
	);
	LUT2 #(
		.INIT('h1)
	) name802 (
		_w945_,
		_w949_,
		_w950_
	);
	LUT2 #(
		.INIT('h1)
	) name803 (
		\pi137 ,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h1)
	) name804 (
		_w941_,
		_w951_,
		_w952_
	);
	LUT2 #(
		.INIT('h1)
	) name805 (
		\pi084 ,
		_w913_,
		_w953_
	);
	LUT2 #(
		.INIT('h4)
	) name806 (
		\pi141 ,
		_w913_,
		_w954_
	);
	LUT2 #(
		.INIT('h1)
	) name807 (
		\pi129 ,
		_w953_,
		_w955_
	);
	LUT2 #(
		.INIT('h4)
	) name808 (
		_w954_,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h4)
	) name809 (
		\pi085 ,
		_w448_,
		_w957_
	);
	LUT2 #(
		.INIT('h8)
	) name810 (
		\pi096 ,
		_w957_,
		_w958_
	);
	LUT2 #(
		.INIT('h1)
	) name811 (
		_w458_,
		_w958_,
		_w959_
	);
	LUT2 #(
		.INIT('h8)
	) name812 (
		_w476_,
		_w482_,
		_w960_
	);
	LUT2 #(
		.INIT('h4)
	) name813 (
		_w959_,
		_w960_,
		_w961_
	);
	LUT2 #(
		.INIT('h1)
	) name814 (
		\pi086 ,
		_w913_,
		_w962_
	);
	LUT2 #(
		.INIT('h4)
	) name815 (
		\pi139 ,
		_w913_,
		_w963_
	);
	LUT2 #(
		.INIT('h1)
	) name816 (
		\pi129 ,
		_w962_,
		_w964_
	);
	LUT2 #(
		.INIT('h4)
	) name817 (
		_w963_,
		_w964_,
		_w965_
	);
	LUT2 #(
		.INIT('h1)
	) name818 (
		\pi087 ,
		_w913_,
		_w966_
	);
	LUT2 #(
		.INIT('h4)
	) name819 (
		\pi140 ,
		_w913_,
		_w967_
	);
	LUT2 #(
		.INIT('h1)
	) name820 (
		\pi129 ,
		_w966_,
		_w968_
	);
	LUT2 #(
		.INIT('h4)
	) name821 (
		_w967_,
		_w968_,
		_w969_
	);
	LUT2 #(
		.INIT('h8)
	) name822 (
		\pi137 ,
		_w934_,
		_w970_
	);
	LUT2 #(
		.INIT('h8)
	) name823 (
		_w843_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h1)
	) name824 (
		\pi088 ,
		_w971_,
		_w972_
	);
	LUT2 #(
		.INIT('h4)
	) name825 (
		\pi139 ,
		_w971_,
		_w973_
	);
	LUT2 #(
		.INIT('h1)
	) name826 (
		\pi129 ,
		_w972_,
		_w974_
	);
	LUT2 #(
		.INIT('h4)
	) name827 (
		_w973_,
		_w974_,
		_w975_
	);
	LUT2 #(
		.INIT('h1)
	) name828 (
		\pi089 ,
		_w971_,
		_w976_
	);
	LUT2 #(
		.INIT('h4)
	) name829 (
		\pi140 ,
		_w971_,
		_w977_
	);
	LUT2 #(
		.INIT('h1)
	) name830 (
		\pi129 ,
		_w976_,
		_w978_
	);
	LUT2 #(
		.INIT('h4)
	) name831 (
		_w977_,
		_w978_,
		_w979_
	);
	LUT2 #(
		.INIT('h1)
	) name832 (
		\pi090 ,
		_w971_,
		_w980_
	);
	LUT2 #(
		.INIT('h4)
	) name833 (
		\pi142 ,
		_w971_,
		_w981_
	);
	LUT2 #(
		.INIT('h1)
	) name834 (
		\pi129 ,
		_w980_,
		_w982_
	);
	LUT2 #(
		.INIT('h4)
	) name835 (
		_w981_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h1)
	) name836 (
		\pi091 ,
		_w971_,
		_w984_
	);
	LUT2 #(
		.INIT('h4)
	) name837 (
		\pi143 ,
		_w971_,
		_w985_
	);
	LUT2 #(
		.INIT('h1)
	) name838 (
		\pi129 ,
		_w984_,
		_w986_
	);
	LUT2 #(
		.INIT('h4)
	) name839 (
		_w985_,
		_w986_,
		_w987_
	);
	LUT2 #(
		.INIT('h1)
	) name840 (
		\pi092 ,
		_w971_,
		_w988_
	);
	LUT2 #(
		.INIT('h4)
	) name841 (
		\pi144 ,
		_w971_,
		_w989_
	);
	LUT2 #(
		.INIT('h1)
	) name842 (
		\pi129 ,
		_w988_,
		_w990_
	);
	LUT2 #(
		.INIT('h4)
	) name843 (
		_w989_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h1)
	) name844 (
		\pi093 ,
		_w971_,
		_w992_
	);
	LUT2 #(
		.INIT('h4)
	) name845 (
		\pi146 ,
		_w971_,
		_w993_
	);
	LUT2 #(
		.INIT('h1)
	) name846 (
		\pi129 ,
		_w992_,
		_w994_
	);
	LUT2 #(
		.INIT('h4)
	) name847 (
		_w993_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h8)
	) name848 (
		\pi082 ,
		\pi138 ,
		_w996_
	);
	LUT2 #(
		.INIT('h8)
	) name849 (
		_w862_,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h8)
	) name850 (
		_w843_,
		_w997_,
		_w998_
	);
	LUT2 #(
		.INIT('h1)
	) name851 (
		\pi094 ,
		_w998_,
		_w999_
	);
	LUT2 #(
		.INIT('h4)
	) name852 (
		\pi142 ,
		_w998_,
		_w1000_
	);
	LUT2 #(
		.INIT('h1)
	) name853 (
		\pi129 ,
		_w999_,
		_w1001_
	);
	LUT2 #(
		.INIT('h4)
	) name854 (
		_w1000_,
		_w1001_,
		_w1002_
	);
	LUT2 #(
		.INIT('h1)
	) name855 (
		\pi003 ,
		\pi110 ,
		_w1003_
	);
	LUT2 #(
		.INIT('h1)
	) name856 (
		_w843_,
		_w1003_,
		_w1004_
	);
	LUT2 #(
		.INIT('h1)
	) name857 (
		_w998_,
		_w1004_,
		_w1005_
	);
	LUT2 #(
		.INIT('h8)
	) name858 (
		\pi095 ,
		_w1005_,
		_w1006_
	);
	LUT2 #(
		.INIT('h8)
	) name859 (
		\pi143 ,
		_w998_,
		_w1007_
	);
	LUT2 #(
		.INIT('h1)
	) name860 (
		_w1006_,
		_w1007_,
		_w1008_
	);
	LUT2 #(
		.INIT('h1)
	) name861 (
		\pi129 ,
		_w1008_,
		_w1009_
	);
	LUT2 #(
		.INIT('h8)
	) name862 (
		\pi096 ,
		_w1005_,
		_w1010_
	);
	LUT2 #(
		.INIT('h8)
	) name863 (
		\pi146 ,
		_w998_,
		_w1011_
	);
	LUT2 #(
		.INIT('h1)
	) name864 (
		_w1010_,
		_w1011_,
		_w1012_
	);
	LUT2 #(
		.INIT('h1)
	) name865 (
		\pi129 ,
		_w1012_,
		_w1013_
	);
	LUT2 #(
		.INIT('h8)
	) name866 (
		\pi097 ,
		_w1005_,
		_w1014_
	);
	LUT2 #(
		.INIT('h8)
	) name867 (
		\pi145 ,
		_w998_,
		_w1015_
	);
	LUT2 #(
		.INIT('h1)
	) name868 (
		_w1014_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('h1)
	) name869 (
		\pi129 ,
		_w1016_,
		_w1017_
	);
	LUT2 #(
		.INIT('h1)
	) name870 (
		\pi098 ,
		_w971_,
		_w1018_
	);
	LUT2 #(
		.INIT('h4)
	) name871 (
		\pi145 ,
		_w971_,
		_w1019_
	);
	LUT2 #(
		.INIT('h1)
	) name872 (
		\pi129 ,
		_w1018_,
		_w1020_
	);
	LUT2 #(
		.INIT('h4)
	) name873 (
		_w1019_,
		_w1020_,
		_w1021_
	);
	LUT2 #(
		.INIT('h1)
	) name874 (
		\pi099 ,
		_w971_,
		_w1022_
	);
	LUT2 #(
		.INIT('h4)
	) name875 (
		\pi141 ,
		_w971_,
		_w1023_
	);
	LUT2 #(
		.INIT('h1)
	) name876 (
		\pi129 ,
		_w1022_,
		_w1024_
	);
	LUT2 #(
		.INIT('h4)
	) name877 (
		_w1023_,
		_w1024_,
		_w1025_
	);
	LUT2 #(
		.INIT('h8)
	) name878 (
		\pi100 ,
		_w1005_,
		_w1026_
	);
	LUT2 #(
		.INIT('h8)
	) name879 (
		\pi144 ,
		_w998_,
		_w1027_
	);
	LUT2 #(
		.INIT('h1)
	) name880 (
		_w1026_,
		_w1027_,
		_w1028_
	);
	LUT2 #(
		.INIT('h1)
	) name881 (
		\pi129 ,
		_w1028_,
		_w1029_
	);
	LUT2 #(
		.INIT('h8)
	) name882 (
		\pi037 ,
		_w934_,
		_w1030_
	);
	LUT2 #(
		.INIT('h1)
	) name883 (
		\pi082 ,
		\pi138 ,
		_w1031_
	);
	LUT2 #(
		.INIT('h4)
	) name884 (
		\pi096 ,
		\pi138 ,
		_w1032_
	);
	LUT2 #(
		.INIT('h1)
	) name885 (
		\pi136 ,
		_w1031_,
		_w1033_
	);
	LUT2 #(
		.INIT('h4)
	) name886 (
		_w1032_,
		_w1033_,
		_w1034_
	);
	LUT2 #(
		.INIT('h1)
	) name887 (
		_w1030_,
		_w1034_,
		_w1035_
	);
	LUT2 #(
		.INIT('h2)
	) name888 (
		\pi137 ,
		_w1035_,
		_w1036_
	);
	LUT2 #(
		.INIT('h4)
	) name889 (
		\pi093 ,
		\pi138 ,
		_w1037_
	);
	LUT2 #(
		.INIT('h2)
	) name890 (
		\pi065 ,
		\pi138 ,
		_w1038_
	);
	LUT2 #(
		.INIT('h2)
	) name891 (
		\pi136 ,
		_w1037_,
		_w1039_
	);
	LUT2 #(
		.INIT('h4)
	) name892 (
		_w1038_,
		_w1039_,
		_w1040_
	);
	LUT2 #(
		.INIT('h4)
	) name893 (
		\pi124 ,
		\pi138 ,
		_w1041_
	);
	LUT2 #(
		.INIT('h2)
	) name894 (
		\pi077 ,
		\pi138 ,
		_w1042_
	);
	LUT2 #(
		.INIT('h1)
	) name895 (
		\pi136 ,
		_w1041_,
		_w1043_
	);
	LUT2 #(
		.INIT('h4)
	) name896 (
		_w1042_,
		_w1043_,
		_w1044_
	);
	LUT2 #(
		.INIT('h1)
	) name897 (
		_w1040_,
		_w1044_,
		_w1045_
	);
	LUT2 #(
		.INIT('h1)
	) name898 (
		\pi137 ,
		_w1045_,
		_w1046_
	);
	LUT2 #(
		.INIT('h1)
	) name899 (
		_w1036_,
		_w1046_,
		_w1047_
	);
	LUT2 #(
		.INIT('h8)
	) name900 (
		\pi091 ,
		_w841_,
		_w1048_
	);
	LUT2 #(
		.INIT('h8)
	) name901 (
		\pi095 ,
		_w912_,
		_w1049_
	);
	LUT2 #(
		.INIT('h1)
	) name902 (
		_w1048_,
		_w1049_,
		_w1050_
	);
	LUT2 #(
		.INIT('h2)
	) name903 (
		\pi138 ,
		_w1050_,
		_w1051_
	);
	LUT2 #(
		.INIT('h1)
	) name904 (
		\pi079 ,
		\pi136 ,
		_w1052_
	);
	LUT2 #(
		.INIT('h4)
	) name905 (
		\pi034 ,
		\pi136 ,
		_w1053_
	);
	LUT2 #(
		.INIT('h2)
	) name906 (
		\pi137 ,
		_w1052_,
		_w1054_
	);
	LUT2 #(
		.INIT('h4)
	) name907 (
		_w1053_,
		_w1054_,
		_w1055_
	);
	LUT2 #(
		.INIT('h2)
	) name908 (
		\pi066 ,
		\pi136 ,
		_w1056_
	);
	LUT2 #(
		.INIT('h8)
	) name909 (
		\pi069 ,
		\pi136 ,
		_w1057_
	);
	LUT2 #(
		.INIT('h1)
	) name910 (
		\pi137 ,
		_w1056_,
		_w1058_
	);
	LUT2 #(
		.INIT('h4)
	) name911 (
		_w1057_,
		_w1058_,
		_w1059_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		_w1055_,
		_w1059_,
		_w1060_
	);
	LUT2 #(
		.INIT('h1)
	) name913 (
		\pi138 ,
		_w1060_,
		_w1061_
	);
	LUT2 #(
		.INIT('h1)
	) name914 (
		_w1051_,
		_w1061_,
		_w1062_
	);
	LUT2 #(
		.INIT('h8)
	) name915 (
		\pi090 ,
		_w841_,
		_w1063_
	);
	LUT2 #(
		.INIT('h8)
	) name916 (
		\pi094 ,
		_w912_,
		_w1064_
	);
	LUT2 #(
		.INIT('h1)
	) name917 (
		_w1063_,
		_w1064_,
		_w1065_
	);
	LUT2 #(
		.INIT('h2)
	) name918 (
		\pi138 ,
		_w1065_,
		_w1066_
	);
	LUT2 #(
		.INIT('h1)
	) name919 (
		\pi078 ,
		\pi136 ,
		_w1067_
	);
	LUT2 #(
		.INIT('h4)
	) name920 (
		\pi033 ,
		\pi136 ,
		_w1068_
	);
	LUT2 #(
		.INIT('h2)
	) name921 (
		\pi137 ,
		_w1067_,
		_w1069_
	);
	LUT2 #(
		.INIT('h4)
	) name922 (
		_w1068_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h2)
	) name923 (
		\pi074 ,
		\pi136 ,
		_w1071_
	);
	LUT2 #(
		.INIT('h8)
	) name924 (
		\pi063 ,
		\pi136 ,
		_w1072_
	);
	LUT2 #(
		.INIT('h1)
	) name925 (
		\pi137 ,
		_w1071_,
		_w1073_
	);
	LUT2 #(
		.INIT('h4)
	) name926 (
		_w1072_,
		_w1073_,
		_w1074_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		_w1070_,
		_w1074_,
		_w1075_
	);
	LUT2 #(
		.INIT('h1)
	) name928 (
		\pi138 ,
		_w1075_,
		_w1076_
	);
	LUT2 #(
		.INIT('h1)
	) name929 (
		_w1066_,
		_w1076_,
		_w1077_
	);
	LUT2 #(
		.INIT('h8)
	) name930 (
		\pi099 ,
		_w841_,
		_w1078_
	);
	LUT2 #(
		.INIT('h4)
	) name931 (
		\pi112 ,
		_w912_,
		_w1079_
	);
	LUT2 #(
		.INIT('h1)
	) name932 (
		_w1078_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h2)
	) name933 (
		\pi138 ,
		_w1080_,
		_w1081_
	);
	LUT2 #(
		.INIT('h1)
	) name934 (
		\pi084 ,
		\pi136 ,
		_w1082_
	);
	LUT2 #(
		.INIT('h4)
	) name935 (
		\pi032 ,
		\pi136 ,
		_w1083_
	);
	LUT2 #(
		.INIT('h2)
	) name936 (
		\pi137 ,
		_w1082_,
		_w1084_
	);
	LUT2 #(
		.INIT('h4)
	) name937 (
		_w1083_,
		_w1084_,
		_w1085_
	);
	LUT2 #(
		.INIT('h2)
	) name938 (
		\pi073 ,
		\pi136 ,
		_w1086_
	);
	LUT2 #(
		.INIT('h8)
	) name939 (
		\pi068 ,
		\pi136 ,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name940 (
		\pi137 ,
		_w1086_,
		_w1088_
	);
	LUT2 #(
		.INIT('h4)
	) name941 (
		_w1087_,
		_w1088_,
		_w1089_
	);
	LUT2 #(
		.INIT('h1)
	) name942 (
		_w1085_,
		_w1089_,
		_w1090_
	);
	LUT2 #(
		.INIT('h1)
	) name943 (
		\pi138 ,
		_w1090_,
		_w1091_
	);
	LUT2 #(
		.INIT('h1)
	) name944 (
		_w1081_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h8)
	) name945 (
		\pi035 ,
		_w934_,
		_w1093_
	);
	LUT2 #(
		.INIT('h1)
	) name946 (
		\pi080 ,
		\pi138 ,
		_w1094_
	);
	LUT2 #(
		.INIT('h4)
	) name947 (
		\pi100 ,
		\pi138 ,
		_w1095_
	);
	LUT2 #(
		.INIT('h1)
	) name948 (
		\pi136 ,
		_w1094_,
		_w1096_
	);
	LUT2 #(
		.INIT('h4)
	) name949 (
		_w1095_,
		_w1096_,
		_w1097_
	);
	LUT2 #(
		.INIT('h1)
	) name950 (
		_w1093_,
		_w1097_,
		_w1098_
	);
	LUT2 #(
		.INIT('h2)
	) name951 (
		\pi137 ,
		_w1098_,
		_w1099_
	);
	LUT2 #(
		.INIT('h4)
	) name952 (
		\pi092 ,
		\pi138 ,
		_w1100_
	);
	LUT2 #(
		.INIT('h2)
	) name953 (
		\pi070 ,
		\pi138 ,
		_w1101_
	);
	LUT2 #(
		.INIT('h2)
	) name954 (
		\pi136 ,
		_w1100_,
		_w1102_
	);
	LUT2 #(
		.INIT('h4)
	) name955 (
		_w1101_,
		_w1102_,
		_w1103_
	);
	LUT2 #(
		.INIT('h4)
	) name956 (
		\pi125 ,
		\pi138 ,
		_w1104_
	);
	LUT2 #(
		.INIT('h2)
	) name957 (
		\pi075 ,
		\pi138 ,
		_w1105_
	);
	LUT2 #(
		.INIT('h1)
	) name958 (
		\pi136 ,
		_w1104_,
		_w1106_
	);
	LUT2 #(
		.INIT('h4)
	) name959 (
		_w1105_,
		_w1106_,
		_w1107_
	);
	LUT2 #(
		.INIT('h1)
	) name960 (
		_w1103_,
		_w1107_,
		_w1108_
	);
	LUT2 #(
		.INIT('h1)
	) name961 (
		\pi137 ,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h1)
	) name962 (
		_w1099_,
		_w1109_,
		_w1110_
	);
	LUT2 #(
		.INIT('h4)
	) name963 (
		\pi026 ,
		_w476_,
		_w1111_
	);
	LUT2 #(
		.INIT('h8)
	) name964 (
		_w957_,
		_w1111_,
		_w1112_
	);
	LUT2 #(
		.INIT('h1)
	) name965 (
		_w485_,
		_w1112_,
		_w1113_
	);
	LUT2 #(
		.INIT('h2)
	) name966 (
		_w148_,
		_w1113_,
		_w1114_
	);
	LUT2 #(
		.INIT('h8)
	) name967 (
		\pi036 ,
		_w934_,
		_w1115_
	);
	LUT2 #(
		.INIT('h1)
	) name968 (
		\pi081 ,
		\pi138 ,
		_w1116_
	);
	LUT2 #(
		.INIT('h4)
	) name969 (
		\pi097 ,
		\pi138 ,
		_w1117_
	);
	LUT2 #(
		.INIT('h1)
	) name970 (
		\pi136 ,
		_w1116_,
		_w1118_
	);
	LUT2 #(
		.INIT('h4)
	) name971 (
		_w1117_,
		_w1118_,
		_w1119_
	);
	LUT2 #(
		.INIT('h1)
	) name972 (
		_w1115_,
		_w1119_,
		_w1120_
	);
	LUT2 #(
		.INIT('h2)
	) name973 (
		\pi137 ,
		_w1120_,
		_w1121_
	);
	LUT2 #(
		.INIT('h4)
	) name974 (
		\pi098 ,
		\pi138 ,
		_w1122_
	);
	LUT2 #(
		.INIT('h2)
	) name975 (
		\pi071 ,
		\pi138 ,
		_w1123_
	);
	LUT2 #(
		.INIT('h2)
	) name976 (
		\pi136 ,
		_w1122_,
		_w1124_
	);
	LUT2 #(
		.INIT('h4)
	) name977 (
		_w1123_,
		_w1124_,
		_w1125_
	);
	LUT2 #(
		.INIT('h4)
	) name978 (
		\pi023 ,
		\pi138 ,
		_w1126_
	);
	LUT2 #(
		.INIT('h2)
	) name979 (
		\pi076 ,
		\pi138 ,
		_w1127_
	);
	LUT2 #(
		.INIT('h1)
	) name980 (
		\pi136 ,
		_w1126_,
		_w1128_
	);
	LUT2 #(
		.INIT('h4)
	) name981 (
		_w1127_,
		_w1128_,
		_w1129_
	);
	LUT2 #(
		.INIT('h1)
	) name982 (
		_w1125_,
		_w1129_,
		_w1130_
	);
	LUT2 #(
		.INIT('h1)
	) name983 (
		\pi137 ,
		_w1130_,
		_w1131_
	);
	LUT2 #(
		.INIT('h1)
	) name984 (
		_w1121_,
		_w1131_,
		_w1132_
	);
	LUT2 #(
		.INIT('h8)
	) name985 (
		\pi030 ,
		_w934_,
		_w1133_
	);
	LUT2 #(
		.INIT('h1)
	) name986 (
		\pi086 ,
		\pi138 ,
		_w1134_
	);
	LUT2 #(
		.INIT('h4)
	) name987 (
		\pi111 ,
		\pi138 ,
		_w1135_
	);
	LUT2 #(
		.INIT('h1)
	) name988 (
		\pi136 ,
		_w1134_,
		_w1136_
	);
	LUT2 #(
		.INIT('h4)
	) name989 (
		_w1135_,
		_w1136_,
		_w1137_
	);
	LUT2 #(
		.INIT('h1)
	) name990 (
		_w1133_,
		_w1137_,
		_w1138_
	);
	LUT2 #(
		.INIT('h2)
	) name991 (
		\pi137 ,
		_w1138_,
		_w1139_
	);
	LUT2 #(
		.INIT('h4)
	) name992 (
		\pi088 ,
		\pi138 ,
		_w1140_
	);
	LUT2 #(
		.INIT('h2)
	) name993 (
		\pi064 ,
		\pi138 ,
		_w1141_
	);
	LUT2 #(
		.INIT('h2)
	) name994 (
		\pi136 ,
		_w1140_,
		_w1142_
	);
	LUT2 #(
		.INIT('h4)
	) name995 (
		_w1141_,
		_w1142_,
		_w1143_
	);
	LUT2 #(
		.INIT('h4)
	) name996 (
		\pi120 ,
		\pi138 ,
		_w1144_
	);
	LUT2 #(
		.INIT('h2)
	) name997 (
		\pi067 ,
		\pi138 ,
		_w1145_
	);
	LUT2 #(
		.INIT('h1)
	) name998 (
		\pi136 ,
		_w1144_,
		_w1146_
	);
	LUT2 #(
		.INIT('h4)
	) name999 (
		_w1145_,
		_w1146_,
		_w1147_
	);
	LUT2 #(
		.INIT('h1)
	) name1000 (
		_w1143_,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h1)
	) name1001 (
		\pi137 ,
		_w1148_,
		_w1149_
	);
	LUT2 #(
		.INIT('h1)
	) name1002 (
		_w1139_,
		_w1149_,
		_w1150_
	);
	LUT2 #(
		.INIT('h8)
	) name1003 (
		\pi116 ,
		_w148_,
		_w1151_
	);
	LUT2 #(
		.INIT('h4)
	) name1004 (
		\pi026 ,
		_w450_,
		_w1152_
	);
	LUT2 #(
		.INIT('h8)
	) name1005 (
		_w506_,
		_w1151_,
		_w1153_
	);
	LUT2 #(
		.INIT('h4)
	) name1006 (
		_w1152_,
		_w1153_,
		_w1154_
	);
	LUT2 #(
		.INIT('h4)
	) name1007 (
		\pi097 ,
		_w438_,
		_w1155_
	);
	LUT2 #(
		.INIT('h1)
	) name1008 (
		_w439_,
		_w1155_,
		_w1156_
	);
	LUT2 #(
		.INIT('h2)
	) name1009 (
		_w1151_,
		_w1156_,
		_w1157_
	);
	LUT2 #(
		.INIT('h4)
	) name1010 (
		\pi129 ,
		_w843_,
		_w1158_
	);
	LUT2 #(
		.INIT('h1)
	) name1011 (
		\pi111 ,
		_w997_,
		_w1159_
	);
	LUT2 #(
		.INIT('h4)
	) name1012 (
		\pi139 ,
		_w997_,
		_w1160_
	);
	LUT2 #(
		.INIT('h2)
	) name1013 (
		_w1158_,
		_w1159_,
		_w1161_
	);
	LUT2 #(
		.INIT('h4)
	) name1014 (
		_w1160_,
		_w1161_,
		_w1162_
	);
	LUT2 #(
		.INIT('h4)
	) name1015 (
		\pi141 ,
		_w997_,
		_w1163_
	);
	LUT2 #(
		.INIT('h2)
	) name1016 (
		\pi112 ,
		_w997_,
		_w1164_
	);
	LUT2 #(
		.INIT('h2)
	) name1017 (
		_w1158_,
		_w1163_,
		_w1165_
	);
	LUT2 #(
		.INIT('h4)
	) name1018 (
		_w1164_,
		_w1165_,
		_w1166_
	);
	LUT2 #(
		.INIT('h4)
	) name1019 (
		\pi011 ,
		_w215_,
		_w1167_
	);
	LUT2 #(
		.INIT('h4)
	) name1020 (
		\pi054 ,
		\pi113 ,
		_w1168_
	);
	LUT2 #(
		.INIT('h2)
	) name1021 (
		_w148_,
		_w1168_,
		_w1169_
	);
	LUT2 #(
		.INIT('h4)
	) name1022 (
		_w1167_,
		_w1169_,
		_w1170_
	);
	LUT2 #(
		.INIT('h4)
	) name1023 (
		\pi140 ,
		_w997_,
		_w1171_
	);
	LUT2 #(
		.INIT('h2)
	) name1024 (
		\pi115 ,
		_w997_,
		_w1172_
	);
	LUT2 #(
		.INIT('h2)
	) name1025 (
		_w1158_,
		_w1171_,
		_w1173_
	);
	LUT2 #(
		.INIT('h4)
	) name1026 (
		_w1172_,
		_w1173_,
		_w1174_
	);
	LUT2 #(
		.INIT('h1)
	) name1027 (
		\pi004 ,
		\pi009 ,
		_w1175_
	);
	LUT2 #(
		.INIT('h8)
	) name1028 (
		_w195_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h8)
	) name1029 (
		\pi054 ,
		_w148_,
		_w1177_
	);
	LUT2 #(
		.INIT('h4)
	) name1030 (
		_w1176_,
		_w1177_,
		_w1178_
	);
	LUT2 #(
		.INIT('h2)
	) name1031 (
		\pi122 ,
		\pi129 ,
		_w1179_
	);
	LUT2 #(
		.INIT('h1)
	) name1032 (
		\pi054 ,
		\pi118 ,
		_w1180_
	);
	LUT2 #(
		.INIT('h2)
	) name1033 (
		\pi054 ,
		_w340_,
		_w1181_
	);
	LUT2 #(
		.INIT('h1)
	) name1034 (
		\pi129 ,
		_w1180_,
		_w1182_
	);
	LUT2 #(
		.INIT('h4)
	) name1035 (
		_w1181_,
		_w1182_,
		_w1183_
	);
	LUT2 #(
		.INIT('h1)
	) name1036 (
		\pi129 ,
		_w446_,
		_w1184_
	);
	LUT2 #(
		.INIT('h4)
	) name1037 (
		\pi120 ,
		_w1003_,
		_w1185_
	);
	LUT2 #(
		.INIT('h1)
	) name1038 (
		\pi111 ,
		\pi129 ,
		_w1186_
	);
	LUT2 #(
		.INIT('h4)
	) name1039 (
		_w1185_,
		_w1186_,
		_w1187_
	);
	LUT2 #(
		.INIT('h8)
	) name1040 (
		\pi081 ,
		\pi120 ,
		_w1188_
	);
	LUT2 #(
		.INIT('h4)
	) name1041 (
		\pi129 ,
		_w1188_,
		_w1189_
	);
	LUT2 #(
		.INIT('h1)
	) name1042 (
		\pi129 ,
		\pi134 ,
		_w1190_
	);
	LUT2 #(
		.INIT('h1)
	) name1043 (
		\pi129 ,
		\pi135 ,
		_w1191_
	);
	LUT2 #(
		.INIT('h2)
	) name1044 (
		\pi057 ,
		\pi129 ,
		_w1192_
	);
	LUT2 #(
		.INIT('h4)
	) name1045 (
		\pi096 ,
		\pi125 ,
		_w1193_
	);
	LUT2 #(
		.INIT('h1)
	) name1046 (
		\pi003 ,
		_w1193_,
		_w1194_
	);
	LUT2 #(
		.INIT('h1)
	) name1047 (
		\pi129 ,
		_w1194_,
		_w1195_
	);
	LUT2 #(
		.INIT('h4)
	) name1048 (
		\pi126 ,
		\pi132 ,
		_w1196_
	);
	LUT2 #(
		.INIT('h8)
	) name1049 (
		\pi133 ,
		_w1196_,
		_w1197_
	);
	assign \po000  = \pi108 ;
	assign \po001  = \pi083 ;
	assign \po002  = \pi104 ;
	assign \po003  = \pi103 ;
	assign \po004  = \pi102 ;
	assign \po005  = \pi105 ;
	assign \po006  = \pi107 ;
	assign \po007  = \pi101 ;
	assign \po008  = \pi126 ;
	assign \po009  = \pi121 ;
	assign \po010  = \pi001 ;
	assign \po011  = \pi000 ;
	assign \po012  = 1'b0;
	assign \po013  = \pi130 ;
	assign \po014  = \pi128 ;
	assign \po015  = _w191_ ;
	assign \po016  = _w223_ ;
	assign \po017  = _w253_ ;
	assign \po018  = _w264_ ;
	assign \po019  = _w271_ ;
	assign \po020  = _w285_ ;
	assign \po021  = _w292_ ;
	assign \po022  = _w301_ ;
	assign \po023  = _w306_ ;
	assign \po024  = _w315_ ;
	assign \po025  = _w323_ ;
	assign \po026  = _w330_ ;
	assign \po027  = _w335_ ;
	assign \po028  = _w344_ ;
	assign \po029  = _w351_ ;
	assign \po030  = _w363_ ;
	assign \po031  = _w369_ ;
	assign \po032  = _w376_ ;
	assign \po033  = _w382_ ;
	assign \po034  = _w387_ ;
	assign \po035  = _w397_ ;
	assign \po036  = _w404_ ;
	assign \po037  = _w411_ ;
	assign \po038  = _w414_ ;
	assign \po039  = _w431_ ;
	assign \po040  = _w475_ ;
	assign \po041  = _w481_ ;
	assign \po042  = _w494_ ;
	assign \po043  = _w533_ ;
	assign \po044  = _w559_ ;
	assign \po045  = _w566_ ;
	assign \po046  = _w573_ ;
	assign \po047  = _w580_ ;
	assign \po048  = _w587_ ;
	assign \po049  = _w594_ ;
	assign \po050  = _w601_ ;
	assign \po051  = _w608_ ;
	assign \po052  = _w615_ ;
	assign \po053  = _w631_ ;
	assign \po054  = _w638_ ;
	assign \po055  = _w652_ ;
	assign \po056  = _w665_ ;
	assign \po057  = _w674_ ;
	assign \po058  = _w685_ ;
	assign \po059  = _w694_ ;
	assign \po060  = _w703_ ;
	assign \po061  = _w714_ ;
	assign \po062  = _w723_ ;
	assign \po063  = _w731_ ;
	assign \po064  = _w740_ ;
	assign \po065  = _w753_ ;
	assign \po066  = _w757_ ;
	assign \po067  = _w761_ ;
	assign \po068  = _w768_ ;
	assign \po069  = _w769_ ;
	assign \po070  = _w772_ ;
	assign \po071  = _w792_ ;
	assign \po072  = _w808_ ;
	assign \po073  = _w814_ ;
	assign \po074  = _w833_ ;
	assign \po075  = _w837_ ;
	assign \po076  = _w840_ ;
	assign \po077  = _w849_ ;
	assign \po078  = _w853_ ;
	assign \po079  = _w857_ ;
	assign \po080  = _w861_ ;
	assign \po081  = _w867_ ;
	assign \po082  = _w871_ ;
	assign \po083  = _w875_ ;
	assign \po084  = _w879_ ;
	assign \po085  = _w883_ ;
	assign \po086  = _w887_ ;
	assign \po087  = _w891_ ;
	assign \po088  = _w895_ ;
	assign \po089  = _w899_ ;
	assign \po090  = _w903_ ;
	assign \po091  = _w907_ ;
	assign \po092  = _w911_ ;
	assign \po093  = _w917_ ;
	assign \po094  = _w921_ ;
	assign \po095  = _w925_ ;
	assign \po096  = _w929_ ;
	assign \po097  = _w933_ ;
	assign \po098  = _w952_ ;
	assign \po099  = _w956_ ;
	assign \po100  = _w961_ ;
	assign \po101  = _w965_ ;
	assign \po102  = _w969_ ;
	assign \po103  = _w975_ ;
	assign \po104  = _w979_ ;
	assign \po105  = _w983_ ;
	assign \po106  = _w987_ ;
	assign \po107  = _w991_ ;
	assign \po108  = _w995_ ;
	assign \po109  = _w1002_ ;
	assign \po110  = _w1009_ ;
	assign \po111  = _w1013_ ;
	assign \po112  = _w1017_ ;
	assign \po113  = _w1021_ ;
	assign \po114  = _w1025_ ;
	assign \po115  = _w1029_ ;
	assign \po116  = _w1047_ ;
	assign \po117  = _w1062_ ;
	assign \po118  = _w1077_ ;
	assign \po119  = _w1092_ ;
	assign \po120  = _w1110_ ;
	assign \po121  = _w1114_ ;
	assign \po122  = _w1132_ ;
	assign \po123  = _w1150_ ;
	assign \po124  = _w1154_ ;
	assign \po125  = _w1157_ ;
	assign \po126  = _w1162_ ;
	assign \po127  = _w1166_ ;
	assign \po128  = _w1170_ ;
	assign \po129  = _w770_ ;
	assign \po130  = _w1174_ ;
	assign \po131  = _w1178_ ;
	assign \po132  = _w1179_ ;
	assign \po133  = _w1183_ ;
	assign \po134  = _w1184_ ;
	assign \po135  = _w1187_ ;
	assign \po136  = _w1189_ ;
	assign \po137  = _w1190_ ;
	assign \po138  = _w1191_ ;
	assign \po139  = _w1192_ ;
	assign \po140  = _w1195_ ;
	assign \po141  = _w1197_ ;
endmodule;