module top( \A[0]_pad  , \A[10]_pad  , \A[11]_pad  , \A[12]_pad  , \A[13]_pad  , \A[14]_pad  , \A[15]_pad  , \A[1]_pad  , \A[2]_pad  , \A[3]_pad  , \A[4]_pad  , \A[5]_pad  , \A[6]_pad  , \A[7]_pad  , \A[8]_pad  , \A[9]_pad  , busrq_n_pad , \di[0]_pad  , \di[1]_pad  , \di[2]_pad  , \di[3]_pad  , \di[4]_pad  , \di[5]_pad  , \di[6]_pad  , \di[7]_pad  , \di_reg_reg[0]/P0001  , \di_reg_reg[1]/P0001  , \di_reg_reg[2]/P0001  , \di_reg_reg[3]/P0001  , \di_reg_reg[4]/P0001  , \di_reg_reg[5]/P0001  , \di_reg_reg[6]/P0001  , \di_reg_reg[7]/P0001  , \do[0]_pad  , \do[1]_pad  , \do[2]_pad  , \do[3]_pad  , \do[4]_pad  , \do[5]_pad  , \do[6]_pad  , \do[7]_pad  , \i_tv80_core_ACC_reg[0]/P0001  , \i_tv80_core_ACC_reg[1]/P0001  , \i_tv80_core_ACC_reg[2]/P0001  , \i_tv80_core_ACC_reg[3]/P0001  , \i_tv80_core_ACC_reg[4]/P0001  , \i_tv80_core_ACC_reg[5]/P0001  , \i_tv80_core_ACC_reg[6]/P0001  , \i_tv80_core_ACC_reg[7]/P0001  , \i_tv80_core_ALU_Op_r_reg[0]/P0001  , \i_tv80_core_ALU_Op_r_reg[1]/P0001  , \i_tv80_core_ALU_Op_r_reg[2]/NET0131  , \i_tv80_core_ALU_Op_r_reg[3]/P0001  , \i_tv80_core_Alternate_reg/P0001  , \i_tv80_core_Ap_reg[0]/P0001  , \i_tv80_core_Ap_reg[1]/P0001  , \i_tv80_core_Ap_reg[2]/P0001  , \i_tv80_core_Ap_reg[3]/P0001  , \i_tv80_core_Ap_reg[4]/P0001  , \i_tv80_core_Ap_reg[5]/P0001  , \i_tv80_core_Ap_reg[6]/P0001  , \i_tv80_core_Ap_reg[7]/P0001  , \i_tv80_core_Arith16_r_reg/P0001  , \i_tv80_core_Auto_Wait_t1_reg/P0001  , \i_tv80_core_Auto_Wait_t2_reg/P0001  , \i_tv80_core_BTR_r_reg/P0001  , \i_tv80_core_BusA_reg[0]/P0001  , \i_tv80_core_BusA_reg[1]/P0001  , \i_tv80_core_BusA_reg[2]/P0001  , \i_tv80_core_BusA_reg[3]/P0001  , \i_tv80_core_BusA_reg[4]/P0001  , \i_tv80_core_BusA_reg[5]/P0001  , \i_tv80_core_BusA_reg[6]/P0001  , \i_tv80_core_BusA_reg[7]/P0001  , \i_tv80_core_BusAck_reg/P0001  , \i_tv80_core_BusB_reg[0]/P0001  , \i_tv80_core_BusB_reg[1]/P0001  , \i_tv80_core_BusB_reg[2]/P0001  , \i_tv80_core_BusB_reg[3]/P0001  , \i_tv80_core_BusB_reg[4]/P0001  , \i_tv80_core_BusB_reg[5]/P0001  , \i_tv80_core_BusB_reg[6]/P0001  , \i_tv80_core_BusB_reg[7]/P0001  , \i_tv80_core_BusReq_s_reg/P0001  , \i_tv80_core_F_reg[0]/P0001  , \i_tv80_core_F_reg[1]/P0001  , \i_tv80_core_F_reg[2]/P0001  , \i_tv80_core_F_reg[3]/P0001  , \i_tv80_core_F_reg[4]/P0001  , \i_tv80_core_F_reg[5]/P0001  , \i_tv80_core_F_reg[6]/P0001  , \i_tv80_core_F_reg[7]/P0001  , \i_tv80_core_Fp_reg[0]/P0001  , \i_tv80_core_Fp_reg[1]/P0001  , \i_tv80_core_Fp_reg[2]/P0001  , \i_tv80_core_Fp_reg[3]/P0001  , \i_tv80_core_Fp_reg[4]/P0001  , \i_tv80_core_Fp_reg[5]/P0001  , \i_tv80_core_Fp_reg[6]/P0001  , \i_tv80_core_Fp_reg[7]/P0001  , \i_tv80_core_Halt_FF_reg/P0001  , \i_tv80_core_INT_s_reg/P0001  , \i_tv80_core_IR_reg[0]/P0001  , \i_tv80_core_IR_reg[1]/P0001  , \i_tv80_core_IR_reg[2]/P0001  , \i_tv80_core_IR_reg[3]/P0001  , \i_tv80_core_IR_reg[4]/P0001  , \i_tv80_core_IR_reg[5]/P0001  , \i_tv80_core_IR_reg[6]/P0001  , \i_tv80_core_IR_reg[7]/P0001  , \i_tv80_core_ISet_reg[0]/NET0131  , \i_tv80_core_ISet_reg[1]/P0001  , \i_tv80_core_IStatus_reg[0]/P0001  , \i_tv80_core_IStatus_reg[1]/P0001  , \i_tv80_core_I_reg[0]/P0001  , \i_tv80_core_I_reg[1]/P0001  , \i_tv80_core_I_reg[2]/P0001  , \i_tv80_core_I_reg[3]/P0001  , \i_tv80_core_I_reg[4]/P0001  , \i_tv80_core_I_reg[5]/P0001  , \i_tv80_core_I_reg[6]/P0001  , \i_tv80_core_I_reg[7]/P0001  , \i_tv80_core_IncDecZ_reg/P0002  , \i_tv80_core_IntCycle_reg/P0001  , \i_tv80_core_IntE_FF1_reg/P0001  , \i_tv80_core_IntE_FF2_reg/P0001  , \i_tv80_core_NMICycle_reg/P0001  , \i_tv80_core_NMI_s_reg/P0001  , \i_tv80_core_No_BTR_reg/P0001  , \i_tv80_core_Oldnmi_n_reg/P0001  , \i_tv80_core_PC_reg[0]/P0001  , \i_tv80_core_PC_reg[10]/P0001  , \i_tv80_core_PC_reg[11]/P0001  , \i_tv80_core_PC_reg[12]/P0001  , \i_tv80_core_PC_reg[13]/P0001  , \i_tv80_core_PC_reg[14]/P0001  , \i_tv80_core_PC_reg[15]/P0001  , \i_tv80_core_PC_reg[1]/P0001  , \i_tv80_core_PC_reg[2]/P0001  , \i_tv80_core_PC_reg[3]/P0001  , \i_tv80_core_PC_reg[4]/P0001  , \i_tv80_core_PC_reg[5]/P0001  , \i_tv80_core_PC_reg[6]/P0001  , \i_tv80_core_PC_reg[7]/P0001  , \i_tv80_core_PC_reg[8]/P0001  , \i_tv80_core_PC_reg[9]/P0001  , \i_tv80_core_Pre_XY_F_M_reg[0]/P0001  , \i_tv80_core_Pre_XY_F_M_reg[1]/P0001  , \i_tv80_core_Pre_XY_F_M_reg[2]/P0001  , \i_tv80_core_PreserveC_r_reg/P0001  , \i_tv80_core_R_reg[0]/P0001  , \i_tv80_core_R_reg[1]/P0001  , \i_tv80_core_R_reg[2]/P0001  , \i_tv80_core_R_reg[3]/P0001  , \i_tv80_core_R_reg[4]/P0001  , \i_tv80_core_R_reg[5]/P0001  , \i_tv80_core_R_reg[6]/P0001  , \i_tv80_core_R_reg[7]/P0001  , \i_tv80_core_Read_To_Reg_r_reg[0]/P0001  , \i_tv80_core_Read_To_Reg_r_reg[1]/P0001  , \i_tv80_core_Read_To_Reg_r_reg[2]/P0001  , \i_tv80_core_Read_To_Reg_r_reg[3]/P0001  , \i_tv80_core_Read_To_Reg_r_reg[4]/P0001  , \i_tv80_core_RegAddrA_r_reg[0]/NET0131  , \i_tv80_core_RegAddrA_r_reg[1]/NET0131  , \i_tv80_core_RegAddrA_r_reg[2]/NET0131  , \i_tv80_core_RegAddrB_r_reg[0]/P0001  , \i_tv80_core_RegAddrB_r_reg[1]/P0001  , \i_tv80_core_RegAddrB_r_reg[2]/P0001  , \i_tv80_core_RegAddrC_reg[0]/P0001  , \i_tv80_core_RegAddrC_reg[1]/NET0131  , \i_tv80_core_RegAddrC_reg[2]/NET0131  , \i_tv80_core_RegBusA_r_reg[0]/P0001  , \i_tv80_core_RegBusA_r_reg[10]/P0001  , \i_tv80_core_RegBusA_r_reg[11]/P0001  , \i_tv80_core_RegBusA_r_reg[12]/P0001  , \i_tv80_core_RegBusA_r_reg[13]/P0001  , \i_tv80_core_RegBusA_r_reg[14]/P0001  , \i_tv80_core_RegBusA_r_reg[15]/P0001  , \i_tv80_core_RegBusA_r_reg[1]/P0001  , \i_tv80_core_RegBusA_r_reg[2]/P0001  , \i_tv80_core_RegBusA_r_reg[3]/P0001  , \i_tv80_core_RegBusA_r_reg[4]/P0001  , \i_tv80_core_RegBusA_r_reg[5]/P0001  , \i_tv80_core_RegBusA_r_reg[6]/P0001  , \i_tv80_core_RegBusA_r_reg[7]/P0001  , \i_tv80_core_RegBusA_r_reg[8]/P0001  , \i_tv80_core_RegBusA_r_reg[9]/P0001  , \i_tv80_core_SP_reg[0]/P0001  , \i_tv80_core_SP_reg[10]/P0001  , \i_tv80_core_SP_reg[11]/P0001  , \i_tv80_core_SP_reg[12]/P0001  , \i_tv80_core_SP_reg[13]/P0001  , \i_tv80_core_SP_reg[14]/P0001  , \i_tv80_core_SP_reg[15]/P0001  , \i_tv80_core_SP_reg[1]/P0001  , \i_tv80_core_SP_reg[2]/P0001  , \i_tv80_core_SP_reg[3]/P0001  , \i_tv80_core_SP_reg[4]/P0001  , \i_tv80_core_SP_reg[5]/P0001  , \i_tv80_core_SP_reg[6]/P0001  , \i_tv80_core_SP_reg[7]/P0001  , \i_tv80_core_SP_reg[8]/P0001  , \i_tv80_core_SP_reg[9]/P0001  , \i_tv80_core_Save_ALU_r_reg/P0001  , \i_tv80_core_TmpAddr_reg[0]/P0001  , \i_tv80_core_TmpAddr_reg[10]/P0001  , \i_tv80_core_TmpAddr_reg[11]/P0001  , \i_tv80_core_TmpAddr_reg[12]/P0001  , \i_tv80_core_TmpAddr_reg[13]/P0001  , \i_tv80_core_TmpAddr_reg[14]/P0001  , \i_tv80_core_TmpAddr_reg[15]/P0001  , \i_tv80_core_TmpAddr_reg[1]/P0001  , \i_tv80_core_TmpAddr_reg[2]/P0001  , \i_tv80_core_TmpAddr_reg[3]/P0001  , \i_tv80_core_TmpAddr_reg[4]/P0001  , \i_tv80_core_TmpAddr_reg[5]/P0001  , \i_tv80_core_TmpAddr_reg[6]/P0001  , \i_tv80_core_TmpAddr_reg[7]/P0001  , \i_tv80_core_TmpAddr_reg[8]/P0001  , \i_tv80_core_TmpAddr_reg[9]/P0001  , \i_tv80_core_XY_Ind_reg/P0001  , \i_tv80_core_XY_State_reg[0]/NET0131  , \i_tv80_core_XY_State_reg[1]/P0001  , \i_tv80_core_Z16_r_reg/P0001  , \i_tv80_core_i_reg_RegsH_reg[0][0]/P0001  , \i_tv80_core_i_reg_RegsH_reg[0][1]/P0001  , \i_tv80_core_i_reg_RegsH_reg[0][2]/P0001  , \i_tv80_core_i_reg_RegsH_reg[0][3]/P0001  , \i_tv80_core_i_reg_RegsH_reg[0][4]/P0001  , \i_tv80_core_i_reg_RegsH_reg[0][5]/P0001  , \i_tv80_core_i_reg_RegsH_reg[0][6]/P0001  , \i_tv80_core_i_reg_RegsH_reg[0][7]/P0002  , \i_tv80_core_i_reg_RegsH_reg[1][0]/P0001  , \i_tv80_core_i_reg_RegsH_reg[1][1]/P0001  , \i_tv80_core_i_reg_RegsH_reg[1][2]/P0001  , \i_tv80_core_i_reg_RegsH_reg[1][3]/P0001  , \i_tv80_core_i_reg_RegsH_reg[1][4]/P0001  , \i_tv80_core_i_reg_RegsH_reg[1][5]/P0001  , \i_tv80_core_i_reg_RegsH_reg[1][6]/P0001  , \i_tv80_core_i_reg_RegsH_reg[1][7]/P0002  , \i_tv80_core_i_reg_RegsH_reg[2][0]/P0001  , \i_tv80_core_i_reg_RegsH_reg[2][1]/P0001  , \i_tv80_core_i_reg_RegsH_reg[2][2]/P0001  , \i_tv80_core_i_reg_RegsH_reg[2][3]/P0001  , \i_tv80_core_i_reg_RegsH_reg[2][4]/P0001  , \i_tv80_core_i_reg_RegsH_reg[2][5]/P0001  , \i_tv80_core_i_reg_RegsH_reg[2][6]/P0001  , \i_tv80_core_i_reg_RegsH_reg[2][7]/P0002  , \i_tv80_core_i_reg_RegsH_reg[3][0]/P0001  , \i_tv80_core_i_reg_RegsH_reg[3][1]/P0001  , \i_tv80_core_i_reg_RegsH_reg[3][2]/P0001  , \i_tv80_core_i_reg_RegsH_reg[3][3]/P0001  , \i_tv80_core_i_reg_RegsH_reg[3][4]/P0001  , \i_tv80_core_i_reg_RegsH_reg[3][5]/P0001  , \i_tv80_core_i_reg_RegsH_reg[3][6]/P0001  , \i_tv80_core_i_reg_RegsH_reg[3][7]/P0002  , \i_tv80_core_i_reg_RegsH_reg[4][0]/P0001  , \i_tv80_core_i_reg_RegsH_reg[4][1]/P0001  , \i_tv80_core_i_reg_RegsH_reg[4][2]/P0001  , \i_tv80_core_i_reg_RegsH_reg[4][3]/P0001  , \i_tv80_core_i_reg_RegsH_reg[4][4]/P0001  , \i_tv80_core_i_reg_RegsH_reg[4][5]/P0001  , \i_tv80_core_i_reg_RegsH_reg[4][6]/P0001  , \i_tv80_core_i_reg_RegsH_reg[4][7]/P0002  , \i_tv80_core_i_reg_RegsH_reg[5][0]/P0001  , \i_tv80_core_i_reg_RegsH_reg[5][1]/P0001  , \i_tv80_core_i_reg_RegsH_reg[5][2]/P0001  , \i_tv80_core_i_reg_RegsH_reg[5][3]/P0001  , \i_tv80_core_i_reg_RegsH_reg[5][4]/P0001  , \i_tv80_core_i_reg_RegsH_reg[5][5]/P0001  , \i_tv80_core_i_reg_RegsH_reg[5][6]/P0001  , \i_tv80_core_i_reg_RegsH_reg[5][7]/P0002  , \i_tv80_core_i_reg_RegsH_reg[6][0]/P0001  , \i_tv80_core_i_reg_RegsH_reg[6][1]/P0001  , \i_tv80_core_i_reg_RegsH_reg[6][2]/P0001  , \i_tv80_core_i_reg_RegsH_reg[6][3]/P0001  , \i_tv80_core_i_reg_RegsH_reg[6][4]/P0001  , \i_tv80_core_i_reg_RegsH_reg[6][5]/P0001  , \i_tv80_core_i_reg_RegsH_reg[6][6]/P0001  , \i_tv80_core_i_reg_RegsH_reg[6][7]/P0002  , \i_tv80_core_i_reg_RegsH_reg[7][0]/P0001  , \i_tv80_core_i_reg_RegsH_reg[7][1]/P0001  , \i_tv80_core_i_reg_RegsH_reg[7][2]/P0001  , \i_tv80_core_i_reg_RegsH_reg[7][3]/P0001  , \i_tv80_core_i_reg_RegsH_reg[7][4]/P0001  , \i_tv80_core_i_reg_RegsH_reg[7][5]/P0001  , \i_tv80_core_i_reg_RegsH_reg[7][6]/P0001  , \i_tv80_core_i_reg_RegsH_reg[7][7]/P0002  , \i_tv80_core_i_reg_RegsL_reg[0][0]/P0001  , \i_tv80_core_i_reg_RegsL_reg[0][1]/P0001  , \i_tv80_core_i_reg_RegsL_reg[0][2]/P0001  , \i_tv80_core_i_reg_RegsL_reg[0][3]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[0][4]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[0][5]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[0][6]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[0][7]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[1][0]/P0001  , \i_tv80_core_i_reg_RegsL_reg[1][1]/P0001  , \i_tv80_core_i_reg_RegsL_reg[1][2]/P0001  , \i_tv80_core_i_reg_RegsL_reg[1][3]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[1][4]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[1][5]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[1][6]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[1][7]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[2][0]/P0001  , \i_tv80_core_i_reg_RegsL_reg[2][1]/P0001  , \i_tv80_core_i_reg_RegsL_reg[2][2]/P0001  , \i_tv80_core_i_reg_RegsL_reg[2][3]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[2][4]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[2][5]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[2][6]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[2][7]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[3][0]/P0001  , \i_tv80_core_i_reg_RegsL_reg[3][1]/P0001  , \i_tv80_core_i_reg_RegsL_reg[3][2]/P0001  , \i_tv80_core_i_reg_RegsL_reg[3][3]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[3][4]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[3][5]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[3][6]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[3][7]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[4][0]/P0001  , \i_tv80_core_i_reg_RegsL_reg[4][1]/P0001  , \i_tv80_core_i_reg_RegsL_reg[4][2]/P0001  , \i_tv80_core_i_reg_RegsL_reg[4][3]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[4][4]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[4][5]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[4][6]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[4][7]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[5][0]/P0001  , \i_tv80_core_i_reg_RegsL_reg[5][1]/P0001  , \i_tv80_core_i_reg_RegsL_reg[5][2]/P0001  , \i_tv80_core_i_reg_RegsL_reg[5][3]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[5][4]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[5][5]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[5][6]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[5][7]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[6][0]/P0001  , \i_tv80_core_i_reg_RegsL_reg[6][1]/P0001  , \i_tv80_core_i_reg_RegsL_reg[6][2]/P0001  , \i_tv80_core_i_reg_RegsL_reg[6][3]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[6][4]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[6][5]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[6][6]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[6][7]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[7][0]/P0001  , \i_tv80_core_i_reg_RegsL_reg[7][1]/P0001  , \i_tv80_core_i_reg_RegsL_reg[7][2]/P0001  , \i_tv80_core_i_reg_RegsL_reg[7][3]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[7][4]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[7][5]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[7][6]/NET0131  , \i_tv80_core_i_reg_RegsL_reg[7][7]/NET0131  , \i_tv80_core_mcycle_reg[0]/P0001  , \i_tv80_core_mcycle_reg[1]/P0001  , \i_tv80_core_mcycle_reg[2]/P0001  , \i_tv80_core_mcycles_reg[0]/P0001  , \i_tv80_core_mcycles_reg[1]/P0001  , \i_tv80_core_mcycles_reg[2]/P0001  , \i_tv80_core_tstate_reg[0]/P0001  , \i_tv80_core_tstate_reg[1]/NET0131  , \i_tv80_core_tstate_reg[2]/NET0131  , int_n_pad , \m1_n_pad  , nmi_n_pad , reset_n_pad , wait_n_pad , \_al_n0  , \_al_n1  , \g28227/_0_  , \g28233/_0_  , \g28274/_0_  , \g28275/_0_  , \g28276/_0_  , \g28277/_0_  , \g28278/_0_  , \g28279/_0_  , \g28280/_0_  , \g28281/_0_  , \g28282/_0_  , \g28283/_0_  , \g28284/_0_  , \g28285/_0_  , \g28286/_0_  , \g28287/_0_  , \g28288/_0_  , \g28289/_0_  , \g28290/_0_  , \g28294/_0_  , \g28295/_0_  , \g28296/_0_  , \g28297/_0_  , \g28298/_0_  , \g28299/_0_  , \g28300/_0_  , \g28301/_0_  , \g28349/_0_  , \g28350/_0_  , \g28351/_0_  , \g28352/_0_  , \g28353/_0_  , \g28354/_0_  , \g28355/_0_  , \g28356/_0_  , \g28357/_0_  , \g28358/_0_  , \g28359/_0_  , \g28360/_0_  , \g28414/_0_  , \g28417/_0_  , \g28418/_0_  , \g28421/_0_  , \g28422/_0_  , \g28423/_0_  , \g28424/_0_  , \g28425/_0_  , \g28426/_0_  , \g28427/_0_  , \g28428/_0_  , \g28429/_0_  , \g28464/_0_  , \g28466/_0_  , \g28470/_0_  , \g28471/_0_  , \g28472/_0_  , \g28473/_0_  , \g28478/_0_  , \g28479/_0_  , \g28500/_0_  , \g28501/_0_  , \g28502/_0_  , \g28503/_0_  , \g28507/_0_  , \g28509/_0_  , \g28536/_0_  , \g28539/_0_  , \g28540/_0_  , \g28543/_0_  , \g28555/_0_  , \g28561/_0_  , \g28562/_0_  , \g28563/_0_  , \g28604/_0_  , \g28606/_0_  , \g28607/_0_  , \g28608/_0_  , \g28609/_0_  , \g28610/_0_  , \g28611/_0_  , \g28612/_0_  , \g28613/_0_  , \g28614/_0_  , \g28616/_0_  , \g28617/_0_  , \g28618/_0_  , \g28660/_0_  , \g28661/_0_  , \g28662/_0_  , \g28663/_0_  , \g28664/_0_  , \g28665/_0_  , \g28666/_0_  , \g28691/_0_  , \g28693/_0_  , \g28694/_0_  , \g28727/_0_  , \g28728/_0_  , \g28729/_0_  , \g28730/_0_  , \g28731/_0_  , \g28732/_0_  , \g28733/_0_  , \g28734/_0_  , \g28750/_0_  , \g28759/_0_  , \g28787/_0_  , \g28788/_0_  , \g28789/_0_  , \g28790/_0_  , \g28791/_0_  , \g28792/_0_  , \g28793/_0_  , \g28794/_0_  , \g28810/_0_  , \g28811/_0_  , \g28812/_0_  , \g28813/_0_  , \g28814/_0_  , \g28835/_0_  , \g28836/_0_  , \g28856/_0_  , \g28857/_0_  , \g28858/_0_  , \g28859/_0_  , \g28860/_0_  , \g28861/_0_  , \g28862/_0_  , \g28863/_0_  , \g28894/_0_  , \g28898/_0_  , \g28914/_0_  , \g28917/_0_  , \g28922/_0_  , \g28923/_0_  , \g28953/_0_  , \g28954/_0_  , \g28955/_0_  , \g28956/_0_  , \g28957/_0_  , \g28958/_0_  , \g28959/_0_  , \g28960/_0_  , \g28970/_0_  , \g28971/_0_  , \g28972/_0_  , \g28973/_0_  , \g28974/_0_  , \g28975/_0_  , \g28976/_0_  , \g28977/_0_  , \g28978/_0_  , \g28979/_0_  , \g28980/_0_  , \g28981/_0_  , \g28982/_0_  , \g28983/_0_  , \g28984/_0_  , \g28985/_0_  , \g28986/_0_  , \g28987/_0_  , \g28988/_0_  , \g28993/_0_  , \g28994/_0_  , \g29029/_0_  , \g29081/_0_  , \g29082/_0_  , \g29083/_0_  , \g29084/_0_  , \g29085/_0_  , \g29086/_0_  , \g29093/_0_  , \g29188/_0_  , \g29189/_0_  , \g29190/_0_  , \g29191/_0_  , \g29192/_0_  , \g29193/_0_  , \g29221/_0_  , \g29222/_0_  , \g29223/_0_  , \g29224/_0_  , \g29225/_0_  , \g29227/_0_  , \g29228/_0_  , \g29229/_0_  , \g29366/_0_  , \g29385/_0_  , \g29387/_0_  , \g29388/_0_  , \g29405/_0_  , \g29450/_0_  , \g29451/_0_  , \g29472/_0_  , \g29552/_0_  , \g29553/_0_  , \g29559/_0_  , \g29561/_0_  , \g29562/_0_  , \g29563/_0_  , \g29564/_0_  , \g29565/_0_  , \g29566/_0_  , \g29577/_0_  , \g29623/_0_  , \g29624/_0_  , \g29625/_0_  , \g29626/_0_  , \g29627/_0_  , \g29628/_0_  , \g29629/_0_  , \g29630/_0_  , \g29657/_0_  , \g29658/_0_  , \g29679/_0_  , \g29689/_3_  , \g29728/_0_  , \g29828/_0_  , \g29909/_3_  , \g29966/_0_  , \g30036/_3_  , \g30038/_3_  , \g30040/_3_  , \g30080/_0_  , \g30081/_0_  , \g30107/_0_  , \g30176/_0_  , \g30189/_3_  , \g30192/_3_  , \g30194/_3_  , \g30354/_0_  , \g30377/_0_  , \g30454/_2_  , \g30479/_2_  , \g30490/_0_  , \g30492/_1_  , \g30495/_0_  , \g30497/_1_  , \g30501/_1_  , \g30503/_1_  , \g30509/_1_  , \g30513/_0_  , \g30514/_0_  , \g30517/_0_  , \g30523/_0_  , \g30678/_0_  , \g30982/_0_  , \g30983/_0_  , \g30984/_0_  , \g30985/_0_  , \g30986/_0_  , \g30987/_0_  , \g30988/_0_  , \g30998/_0_  , \g31212/_0_  , \g31235/_0_  , \g31236/_0_  , \g31296/_3_  , \g31303/_0_  , \g31306/_0_  , \g31312/_0_  , \g31356/_0_  , \g31397/_0_  , \g31430/_0_  , \g31440/_3_  , \g31455/_3_  , \g31459/_0_  , \g31511/_0_  , \g31512/_0_  , \g31561/_0_  , \g31603/_0_  , \g31604/_0_  , \g31666/_0_  , \g31794/_0_  , \g31795/_0_  , \g31796/_0_  , \g31854/_0_  , \g31855/_0_  , \g31856/_0_  , \g31871/_0_  , \g31920/_0_  , \g31934/_0_  , \g31935/_0_  , \g31943/_0_  , \g32128/_0_  , \g32129/_0_  , \g32130/_0_  , \g32131/_0_  , \g32132/_0_  , \g32133/_0_  , \g32134/_0_  , \g32135/_0_  , \g32136/_0_  , \g32137/_0_  , \g32140/_0_  , \g32141/_0_  , \g32142/_0_  , \g32143/_0_  , \g32144/_0_  , \g32145/_0_  , \g32146/_0_  , \g32147/_0_  , \g32475/_0_  , \g32639/_0_  , \g32640/_0_  , \g32641/_0_  , \g32642/_0_  , \g32643/_0_  , \g32644/_0_  , \g32645/_0_  , \g32646/_0_  , \g32647/_0_  , \g32648/_0_  , \g32649/_0_  , \g32650/_0_  , \g32651/_0_  , \g32652/_0_  , \g32653/_0_  , \g32654/_0_  , \g32798/_3_  , \g33177/_0_  , \g33187/_0_  , \g33306/_0_  , \g33307/_0_  , \g33308/_0_  , \g33309/_0_  , \g33310/_0_  , \g33311/_0_  , \g33312/_0_  , \g33313/_0_  , \g34088/_0_  , \g35570/_0_  , \g35594/_0_  , \g35838/_0_  , \g37467/_0_  , \g37492/_0_  , \g37503/_0_  , \g37513/_0_  , \g37524/_0_  , \g37727/_0_  , \g37748/_0_  , \g37758/_0_  , \g37767/_0_  , \g37777/_0_  , \g37790/_0_  , \g37809/_0_  , \g37840/_0_  , \g37852/_0_  , \g38312_dup/_0_  , \g38324/_0_  , \g38354/_0_  , \g38781/_1_  , \g38840/_0_  , \g38851/_0_  , \g38866/_0_  , \g38892/_1_  , \g38932/_0_  , \g38943/_0_  , \g39103/_0_  , \g39113/_2__syn_2  , \g39127/_0_  , \g44/_0_  , halt_n_pad );
  input \A[0]_pad  ;
  input \A[10]_pad  ;
  input \A[11]_pad  ;
  input \A[12]_pad  ;
  input \A[13]_pad  ;
  input \A[14]_pad  ;
  input \A[15]_pad  ;
  input \A[1]_pad  ;
  input \A[2]_pad  ;
  input \A[3]_pad  ;
  input \A[4]_pad  ;
  input \A[5]_pad  ;
  input \A[6]_pad  ;
  input \A[7]_pad  ;
  input \A[8]_pad  ;
  input \A[9]_pad  ;
  input busrq_n_pad ;
  input \di[0]_pad  ;
  input \di[1]_pad  ;
  input \di[2]_pad  ;
  input \di[3]_pad  ;
  input \di[4]_pad  ;
  input \di[5]_pad  ;
  input \di[6]_pad  ;
  input \di[7]_pad  ;
  input \di_reg_reg[0]/P0001  ;
  input \di_reg_reg[1]/P0001  ;
  input \di_reg_reg[2]/P0001  ;
  input \di_reg_reg[3]/P0001  ;
  input \di_reg_reg[4]/P0001  ;
  input \di_reg_reg[5]/P0001  ;
  input \di_reg_reg[6]/P0001  ;
  input \di_reg_reg[7]/P0001  ;
  input \do[0]_pad  ;
  input \do[1]_pad  ;
  input \do[2]_pad  ;
  input \do[3]_pad  ;
  input \do[4]_pad  ;
  input \do[5]_pad  ;
  input \do[6]_pad  ;
  input \do[7]_pad  ;
  input \i_tv80_core_ACC_reg[0]/P0001  ;
  input \i_tv80_core_ACC_reg[1]/P0001  ;
  input \i_tv80_core_ACC_reg[2]/P0001  ;
  input \i_tv80_core_ACC_reg[3]/P0001  ;
  input \i_tv80_core_ACC_reg[4]/P0001  ;
  input \i_tv80_core_ACC_reg[5]/P0001  ;
  input \i_tv80_core_ACC_reg[6]/P0001  ;
  input \i_tv80_core_ACC_reg[7]/P0001  ;
  input \i_tv80_core_ALU_Op_r_reg[0]/P0001  ;
  input \i_tv80_core_ALU_Op_r_reg[1]/P0001  ;
  input \i_tv80_core_ALU_Op_r_reg[2]/NET0131  ;
  input \i_tv80_core_ALU_Op_r_reg[3]/P0001  ;
  input \i_tv80_core_Alternate_reg/P0001  ;
  input \i_tv80_core_Ap_reg[0]/P0001  ;
  input \i_tv80_core_Ap_reg[1]/P0001  ;
  input \i_tv80_core_Ap_reg[2]/P0001  ;
  input \i_tv80_core_Ap_reg[3]/P0001  ;
  input \i_tv80_core_Ap_reg[4]/P0001  ;
  input \i_tv80_core_Ap_reg[5]/P0001  ;
  input \i_tv80_core_Ap_reg[6]/P0001  ;
  input \i_tv80_core_Ap_reg[7]/P0001  ;
  input \i_tv80_core_Arith16_r_reg/P0001  ;
  input \i_tv80_core_Auto_Wait_t1_reg/P0001  ;
  input \i_tv80_core_Auto_Wait_t2_reg/P0001  ;
  input \i_tv80_core_BTR_r_reg/P0001  ;
  input \i_tv80_core_BusA_reg[0]/P0001  ;
  input \i_tv80_core_BusA_reg[1]/P0001  ;
  input \i_tv80_core_BusA_reg[2]/P0001  ;
  input \i_tv80_core_BusA_reg[3]/P0001  ;
  input \i_tv80_core_BusA_reg[4]/P0001  ;
  input \i_tv80_core_BusA_reg[5]/P0001  ;
  input \i_tv80_core_BusA_reg[6]/P0001  ;
  input \i_tv80_core_BusA_reg[7]/P0001  ;
  input \i_tv80_core_BusAck_reg/P0001  ;
  input \i_tv80_core_BusB_reg[0]/P0001  ;
  input \i_tv80_core_BusB_reg[1]/P0001  ;
  input \i_tv80_core_BusB_reg[2]/P0001  ;
  input \i_tv80_core_BusB_reg[3]/P0001  ;
  input \i_tv80_core_BusB_reg[4]/P0001  ;
  input \i_tv80_core_BusB_reg[5]/P0001  ;
  input \i_tv80_core_BusB_reg[6]/P0001  ;
  input \i_tv80_core_BusB_reg[7]/P0001  ;
  input \i_tv80_core_BusReq_s_reg/P0001  ;
  input \i_tv80_core_F_reg[0]/P0001  ;
  input \i_tv80_core_F_reg[1]/P0001  ;
  input \i_tv80_core_F_reg[2]/P0001  ;
  input \i_tv80_core_F_reg[3]/P0001  ;
  input \i_tv80_core_F_reg[4]/P0001  ;
  input \i_tv80_core_F_reg[5]/P0001  ;
  input \i_tv80_core_F_reg[6]/P0001  ;
  input \i_tv80_core_F_reg[7]/P0001  ;
  input \i_tv80_core_Fp_reg[0]/P0001  ;
  input \i_tv80_core_Fp_reg[1]/P0001  ;
  input \i_tv80_core_Fp_reg[2]/P0001  ;
  input \i_tv80_core_Fp_reg[3]/P0001  ;
  input \i_tv80_core_Fp_reg[4]/P0001  ;
  input \i_tv80_core_Fp_reg[5]/P0001  ;
  input \i_tv80_core_Fp_reg[6]/P0001  ;
  input \i_tv80_core_Fp_reg[7]/P0001  ;
  input \i_tv80_core_Halt_FF_reg/P0001  ;
  input \i_tv80_core_INT_s_reg/P0001  ;
  input \i_tv80_core_IR_reg[0]/P0001  ;
  input \i_tv80_core_IR_reg[1]/P0001  ;
  input \i_tv80_core_IR_reg[2]/P0001  ;
  input \i_tv80_core_IR_reg[3]/P0001  ;
  input \i_tv80_core_IR_reg[4]/P0001  ;
  input \i_tv80_core_IR_reg[5]/P0001  ;
  input \i_tv80_core_IR_reg[6]/P0001  ;
  input \i_tv80_core_IR_reg[7]/P0001  ;
  input \i_tv80_core_ISet_reg[0]/NET0131  ;
  input \i_tv80_core_ISet_reg[1]/P0001  ;
  input \i_tv80_core_IStatus_reg[0]/P0001  ;
  input \i_tv80_core_IStatus_reg[1]/P0001  ;
  input \i_tv80_core_I_reg[0]/P0001  ;
  input \i_tv80_core_I_reg[1]/P0001  ;
  input \i_tv80_core_I_reg[2]/P0001  ;
  input \i_tv80_core_I_reg[3]/P0001  ;
  input \i_tv80_core_I_reg[4]/P0001  ;
  input \i_tv80_core_I_reg[5]/P0001  ;
  input \i_tv80_core_I_reg[6]/P0001  ;
  input \i_tv80_core_I_reg[7]/P0001  ;
  input \i_tv80_core_IncDecZ_reg/P0002  ;
  input \i_tv80_core_IntCycle_reg/P0001  ;
  input \i_tv80_core_IntE_FF1_reg/P0001  ;
  input \i_tv80_core_IntE_FF2_reg/P0001  ;
  input \i_tv80_core_NMICycle_reg/P0001  ;
  input \i_tv80_core_NMI_s_reg/P0001  ;
  input \i_tv80_core_No_BTR_reg/P0001  ;
  input \i_tv80_core_Oldnmi_n_reg/P0001  ;
  input \i_tv80_core_PC_reg[0]/P0001  ;
  input \i_tv80_core_PC_reg[10]/P0001  ;
  input \i_tv80_core_PC_reg[11]/P0001  ;
  input \i_tv80_core_PC_reg[12]/P0001  ;
  input \i_tv80_core_PC_reg[13]/P0001  ;
  input \i_tv80_core_PC_reg[14]/P0001  ;
  input \i_tv80_core_PC_reg[15]/P0001  ;
  input \i_tv80_core_PC_reg[1]/P0001  ;
  input \i_tv80_core_PC_reg[2]/P0001  ;
  input \i_tv80_core_PC_reg[3]/P0001  ;
  input \i_tv80_core_PC_reg[4]/P0001  ;
  input \i_tv80_core_PC_reg[5]/P0001  ;
  input \i_tv80_core_PC_reg[6]/P0001  ;
  input \i_tv80_core_PC_reg[7]/P0001  ;
  input \i_tv80_core_PC_reg[8]/P0001  ;
  input \i_tv80_core_PC_reg[9]/P0001  ;
  input \i_tv80_core_Pre_XY_F_M_reg[0]/P0001  ;
  input \i_tv80_core_Pre_XY_F_M_reg[1]/P0001  ;
  input \i_tv80_core_Pre_XY_F_M_reg[2]/P0001  ;
  input \i_tv80_core_PreserveC_r_reg/P0001  ;
  input \i_tv80_core_R_reg[0]/P0001  ;
  input \i_tv80_core_R_reg[1]/P0001  ;
  input \i_tv80_core_R_reg[2]/P0001  ;
  input \i_tv80_core_R_reg[3]/P0001  ;
  input \i_tv80_core_R_reg[4]/P0001  ;
  input \i_tv80_core_R_reg[5]/P0001  ;
  input \i_tv80_core_R_reg[6]/P0001  ;
  input \i_tv80_core_R_reg[7]/P0001  ;
  input \i_tv80_core_Read_To_Reg_r_reg[0]/P0001  ;
  input \i_tv80_core_Read_To_Reg_r_reg[1]/P0001  ;
  input \i_tv80_core_Read_To_Reg_r_reg[2]/P0001  ;
  input \i_tv80_core_Read_To_Reg_r_reg[3]/P0001  ;
  input \i_tv80_core_Read_To_Reg_r_reg[4]/P0001  ;
  input \i_tv80_core_RegAddrA_r_reg[0]/NET0131  ;
  input \i_tv80_core_RegAddrA_r_reg[1]/NET0131  ;
  input \i_tv80_core_RegAddrA_r_reg[2]/NET0131  ;
  input \i_tv80_core_RegAddrB_r_reg[0]/P0001  ;
  input \i_tv80_core_RegAddrB_r_reg[1]/P0001  ;
  input \i_tv80_core_RegAddrB_r_reg[2]/P0001  ;
  input \i_tv80_core_RegAddrC_reg[0]/P0001  ;
  input \i_tv80_core_RegAddrC_reg[1]/NET0131  ;
  input \i_tv80_core_RegAddrC_reg[2]/NET0131  ;
  input \i_tv80_core_RegBusA_r_reg[0]/P0001  ;
  input \i_tv80_core_RegBusA_r_reg[10]/P0001  ;
  input \i_tv80_core_RegBusA_r_reg[11]/P0001  ;
  input \i_tv80_core_RegBusA_r_reg[12]/P0001  ;
  input \i_tv80_core_RegBusA_r_reg[13]/P0001  ;
  input \i_tv80_core_RegBusA_r_reg[14]/P0001  ;
  input \i_tv80_core_RegBusA_r_reg[15]/P0001  ;
  input \i_tv80_core_RegBusA_r_reg[1]/P0001  ;
  input \i_tv80_core_RegBusA_r_reg[2]/P0001  ;
  input \i_tv80_core_RegBusA_r_reg[3]/P0001  ;
  input \i_tv80_core_RegBusA_r_reg[4]/P0001  ;
  input \i_tv80_core_RegBusA_r_reg[5]/P0001  ;
  input \i_tv80_core_RegBusA_r_reg[6]/P0001  ;
  input \i_tv80_core_RegBusA_r_reg[7]/P0001  ;
  input \i_tv80_core_RegBusA_r_reg[8]/P0001  ;
  input \i_tv80_core_RegBusA_r_reg[9]/P0001  ;
  input \i_tv80_core_SP_reg[0]/P0001  ;
  input \i_tv80_core_SP_reg[10]/P0001  ;
  input \i_tv80_core_SP_reg[11]/P0001  ;
  input \i_tv80_core_SP_reg[12]/P0001  ;
  input \i_tv80_core_SP_reg[13]/P0001  ;
  input \i_tv80_core_SP_reg[14]/P0001  ;
  input \i_tv80_core_SP_reg[15]/P0001  ;
  input \i_tv80_core_SP_reg[1]/P0001  ;
  input \i_tv80_core_SP_reg[2]/P0001  ;
  input \i_tv80_core_SP_reg[3]/P0001  ;
  input \i_tv80_core_SP_reg[4]/P0001  ;
  input \i_tv80_core_SP_reg[5]/P0001  ;
  input \i_tv80_core_SP_reg[6]/P0001  ;
  input \i_tv80_core_SP_reg[7]/P0001  ;
  input \i_tv80_core_SP_reg[8]/P0001  ;
  input \i_tv80_core_SP_reg[9]/P0001  ;
  input \i_tv80_core_Save_ALU_r_reg/P0001  ;
  input \i_tv80_core_TmpAddr_reg[0]/P0001  ;
  input \i_tv80_core_TmpAddr_reg[10]/P0001  ;
  input \i_tv80_core_TmpAddr_reg[11]/P0001  ;
  input \i_tv80_core_TmpAddr_reg[12]/P0001  ;
  input \i_tv80_core_TmpAddr_reg[13]/P0001  ;
  input \i_tv80_core_TmpAddr_reg[14]/P0001  ;
  input \i_tv80_core_TmpAddr_reg[15]/P0001  ;
  input \i_tv80_core_TmpAddr_reg[1]/P0001  ;
  input \i_tv80_core_TmpAddr_reg[2]/P0001  ;
  input \i_tv80_core_TmpAddr_reg[3]/P0001  ;
  input \i_tv80_core_TmpAddr_reg[4]/P0001  ;
  input \i_tv80_core_TmpAddr_reg[5]/P0001  ;
  input \i_tv80_core_TmpAddr_reg[6]/P0001  ;
  input \i_tv80_core_TmpAddr_reg[7]/P0001  ;
  input \i_tv80_core_TmpAddr_reg[8]/P0001  ;
  input \i_tv80_core_TmpAddr_reg[9]/P0001  ;
  input \i_tv80_core_XY_Ind_reg/P0001  ;
  input \i_tv80_core_XY_State_reg[0]/NET0131  ;
  input \i_tv80_core_XY_State_reg[1]/P0001  ;
  input \i_tv80_core_Z16_r_reg/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[0][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[0][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[0][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[0][3]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[0][4]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[0][5]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[0][6]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[0][7]/P0002  ;
  input \i_tv80_core_i_reg_RegsH_reg[1][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[1][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[1][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[1][3]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[1][4]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[1][5]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[1][6]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[1][7]/P0002  ;
  input \i_tv80_core_i_reg_RegsH_reg[2][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[2][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[2][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[2][3]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[2][4]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[2][5]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[2][6]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[2][7]/P0002  ;
  input \i_tv80_core_i_reg_RegsH_reg[3][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[3][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[3][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[3][3]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[3][4]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[3][5]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[3][6]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[3][7]/P0002  ;
  input \i_tv80_core_i_reg_RegsH_reg[4][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[4][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[4][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[4][3]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[4][4]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[4][5]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[4][6]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[4][7]/P0002  ;
  input \i_tv80_core_i_reg_RegsH_reg[5][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[5][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[5][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[5][3]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[5][4]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[5][5]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[5][6]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[5][7]/P0002  ;
  input \i_tv80_core_i_reg_RegsH_reg[6][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[6][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[6][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[6][3]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[6][4]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[6][5]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[6][6]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[6][7]/P0002  ;
  input \i_tv80_core_i_reg_RegsH_reg[7][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[7][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[7][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[7][3]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[7][4]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[7][5]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[7][6]/P0001  ;
  input \i_tv80_core_i_reg_RegsH_reg[7][7]/P0002  ;
  input \i_tv80_core_i_reg_RegsL_reg[0][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[0][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[0][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[0][3]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[0][4]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[0][5]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[0][6]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[0][7]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[1][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[1][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[1][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[1][3]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[1][4]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[1][5]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[1][6]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[1][7]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[2][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[2][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[2][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[2][3]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[2][4]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[2][5]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[2][6]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[2][7]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[3][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[3][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[3][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[3][3]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[3][4]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[3][5]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[3][6]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[3][7]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[4][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[4][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[4][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[4][3]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[4][4]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[4][5]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[4][6]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[4][7]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[5][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[5][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[5][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[5][3]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[5][4]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[5][5]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[5][6]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[5][7]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[6][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[6][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[6][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[6][3]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[6][4]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[6][5]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[6][6]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[6][7]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[7][0]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[7][1]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[7][2]/P0001  ;
  input \i_tv80_core_i_reg_RegsL_reg[7][3]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[7][4]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[7][5]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[7][6]/NET0131  ;
  input \i_tv80_core_i_reg_RegsL_reg[7][7]/NET0131  ;
  input \i_tv80_core_mcycle_reg[0]/P0001  ;
  input \i_tv80_core_mcycle_reg[1]/P0001  ;
  input \i_tv80_core_mcycle_reg[2]/P0001  ;
  input \i_tv80_core_mcycles_reg[0]/P0001  ;
  input \i_tv80_core_mcycles_reg[1]/P0001  ;
  input \i_tv80_core_mcycles_reg[2]/P0001  ;
  input \i_tv80_core_tstate_reg[0]/P0001  ;
  input \i_tv80_core_tstate_reg[1]/NET0131  ;
  input \i_tv80_core_tstate_reg[2]/NET0131  ;
  input int_n_pad ;
  input \m1_n_pad  ;
  input nmi_n_pad ;
  input reset_n_pad ;
  input wait_n_pad ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g28227/_0_  ;
  output \g28233/_0_  ;
  output \g28274/_0_  ;
  output \g28275/_0_  ;
  output \g28276/_0_  ;
  output \g28277/_0_  ;
  output \g28278/_0_  ;
  output \g28279/_0_  ;
  output \g28280/_0_  ;
  output \g28281/_0_  ;
  output \g28282/_0_  ;
  output \g28283/_0_  ;
  output \g28284/_0_  ;
  output \g28285/_0_  ;
  output \g28286/_0_  ;
  output \g28287/_0_  ;
  output \g28288/_0_  ;
  output \g28289/_0_  ;
  output \g28290/_0_  ;
  output \g28294/_0_  ;
  output \g28295/_0_  ;
  output \g28296/_0_  ;
  output \g28297/_0_  ;
  output \g28298/_0_  ;
  output \g28299/_0_  ;
  output \g28300/_0_  ;
  output \g28301/_0_  ;
  output \g28349/_0_  ;
  output \g28350/_0_  ;
  output \g28351/_0_  ;
  output \g28352/_0_  ;
  output \g28353/_0_  ;
  output \g28354/_0_  ;
  output \g28355/_0_  ;
  output \g28356/_0_  ;
  output \g28357/_0_  ;
  output \g28358/_0_  ;
  output \g28359/_0_  ;
  output \g28360/_0_  ;
  output \g28414/_0_  ;
  output \g28417/_0_  ;
  output \g28418/_0_  ;
  output \g28421/_0_  ;
  output \g28422/_0_  ;
  output \g28423/_0_  ;
  output \g28424/_0_  ;
  output \g28425/_0_  ;
  output \g28426/_0_  ;
  output \g28427/_0_  ;
  output \g28428/_0_  ;
  output \g28429/_0_  ;
  output \g28464/_0_  ;
  output \g28466/_0_  ;
  output \g28470/_0_  ;
  output \g28471/_0_  ;
  output \g28472/_0_  ;
  output \g28473/_0_  ;
  output \g28478/_0_  ;
  output \g28479/_0_  ;
  output \g28500/_0_  ;
  output \g28501/_0_  ;
  output \g28502/_0_  ;
  output \g28503/_0_  ;
  output \g28507/_0_  ;
  output \g28509/_0_  ;
  output \g28536/_0_  ;
  output \g28539/_0_  ;
  output \g28540/_0_  ;
  output \g28543/_0_  ;
  output \g28555/_0_  ;
  output \g28561/_0_  ;
  output \g28562/_0_  ;
  output \g28563/_0_  ;
  output \g28604/_0_  ;
  output \g28606/_0_  ;
  output \g28607/_0_  ;
  output \g28608/_0_  ;
  output \g28609/_0_  ;
  output \g28610/_0_  ;
  output \g28611/_0_  ;
  output \g28612/_0_  ;
  output \g28613/_0_  ;
  output \g28614/_0_  ;
  output \g28616/_0_  ;
  output \g28617/_0_  ;
  output \g28618/_0_  ;
  output \g28660/_0_  ;
  output \g28661/_0_  ;
  output \g28662/_0_  ;
  output \g28663/_0_  ;
  output \g28664/_0_  ;
  output \g28665/_0_  ;
  output \g28666/_0_  ;
  output \g28691/_0_  ;
  output \g28693/_0_  ;
  output \g28694/_0_  ;
  output \g28727/_0_  ;
  output \g28728/_0_  ;
  output \g28729/_0_  ;
  output \g28730/_0_  ;
  output \g28731/_0_  ;
  output \g28732/_0_  ;
  output \g28733/_0_  ;
  output \g28734/_0_  ;
  output \g28750/_0_  ;
  output \g28759/_0_  ;
  output \g28787/_0_  ;
  output \g28788/_0_  ;
  output \g28789/_0_  ;
  output \g28790/_0_  ;
  output \g28791/_0_  ;
  output \g28792/_0_  ;
  output \g28793/_0_  ;
  output \g28794/_0_  ;
  output \g28810/_0_  ;
  output \g28811/_0_  ;
  output \g28812/_0_  ;
  output \g28813/_0_  ;
  output \g28814/_0_  ;
  output \g28835/_0_  ;
  output \g28836/_0_  ;
  output \g28856/_0_  ;
  output \g28857/_0_  ;
  output \g28858/_0_  ;
  output \g28859/_0_  ;
  output \g28860/_0_  ;
  output \g28861/_0_  ;
  output \g28862/_0_  ;
  output \g28863/_0_  ;
  output \g28894/_0_  ;
  output \g28898/_0_  ;
  output \g28914/_0_  ;
  output \g28917/_0_  ;
  output \g28922/_0_  ;
  output \g28923/_0_  ;
  output \g28953/_0_  ;
  output \g28954/_0_  ;
  output \g28955/_0_  ;
  output \g28956/_0_  ;
  output \g28957/_0_  ;
  output \g28958/_0_  ;
  output \g28959/_0_  ;
  output \g28960/_0_  ;
  output \g28970/_0_  ;
  output \g28971/_0_  ;
  output \g28972/_0_  ;
  output \g28973/_0_  ;
  output \g28974/_0_  ;
  output \g28975/_0_  ;
  output \g28976/_0_  ;
  output \g28977/_0_  ;
  output \g28978/_0_  ;
  output \g28979/_0_  ;
  output \g28980/_0_  ;
  output \g28981/_0_  ;
  output \g28982/_0_  ;
  output \g28983/_0_  ;
  output \g28984/_0_  ;
  output \g28985/_0_  ;
  output \g28986/_0_  ;
  output \g28987/_0_  ;
  output \g28988/_0_  ;
  output \g28993/_0_  ;
  output \g28994/_0_  ;
  output \g29029/_0_  ;
  output \g29081/_0_  ;
  output \g29082/_0_  ;
  output \g29083/_0_  ;
  output \g29084/_0_  ;
  output \g29085/_0_  ;
  output \g29086/_0_  ;
  output \g29093/_0_  ;
  output \g29188/_0_  ;
  output \g29189/_0_  ;
  output \g29190/_0_  ;
  output \g29191/_0_  ;
  output \g29192/_0_  ;
  output \g29193/_0_  ;
  output \g29221/_0_  ;
  output \g29222/_0_  ;
  output \g29223/_0_  ;
  output \g29224/_0_  ;
  output \g29225/_0_  ;
  output \g29227/_0_  ;
  output \g29228/_0_  ;
  output \g29229/_0_  ;
  output \g29366/_0_  ;
  output \g29385/_0_  ;
  output \g29387/_0_  ;
  output \g29388/_0_  ;
  output \g29405/_0_  ;
  output \g29450/_0_  ;
  output \g29451/_0_  ;
  output \g29472/_0_  ;
  output \g29552/_0_  ;
  output \g29553/_0_  ;
  output \g29559/_0_  ;
  output \g29561/_0_  ;
  output \g29562/_0_  ;
  output \g29563/_0_  ;
  output \g29564/_0_  ;
  output \g29565/_0_  ;
  output \g29566/_0_  ;
  output \g29577/_0_  ;
  output \g29623/_0_  ;
  output \g29624/_0_  ;
  output \g29625/_0_  ;
  output \g29626/_0_  ;
  output \g29627/_0_  ;
  output \g29628/_0_  ;
  output \g29629/_0_  ;
  output \g29630/_0_  ;
  output \g29657/_0_  ;
  output \g29658/_0_  ;
  output \g29679/_0_  ;
  output \g29689/_3_  ;
  output \g29728/_0_  ;
  output \g29828/_0_  ;
  output \g29909/_3_  ;
  output \g29966/_0_  ;
  output \g30036/_3_  ;
  output \g30038/_3_  ;
  output \g30040/_3_  ;
  output \g30080/_0_  ;
  output \g30081/_0_  ;
  output \g30107/_0_  ;
  output \g30176/_0_  ;
  output \g30189/_3_  ;
  output \g30192/_3_  ;
  output \g30194/_3_  ;
  output \g30354/_0_  ;
  output \g30377/_0_  ;
  output \g30454/_2_  ;
  output \g30479/_2_  ;
  output \g30490/_0_  ;
  output \g30492/_1_  ;
  output \g30495/_0_  ;
  output \g30497/_1_  ;
  output \g30501/_1_  ;
  output \g30503/_1_  ;
  output \g30509/_1_  ;
  output \g30513/_0_  ;
  output \g30514/_0_  ;
  output \g30517/_0_  ;
  output \g30523/_0_  ;
  output \g30678/_0_  ;
  output \g30982/_0_  ;
  output \g30983/_0_  ;
  output \g30984/_0_  ;
  output \g30985/_0_  ;
  output \g30986/_0_  ;
  output \g30987/_0_  ;
  output \g30988/_0_  ;
  output \g30998/_0_  ;
  output \g31212/_0_  ;
  output \g31235/_0_  ;
  output \g31236/_0_  ;
  output \g31296/_3_  ;
  output \g31303/_0_  ;
  output \g31306/_0_  ;
  output \g31312/_0_  ;
  output \g31356/_0_  ;
  output \g31397/_0_  ;
  output \g31430/_0_  ;
  output \g31440/_3_  ;
  output \g31455/_3_  ;
  output \g31459/_0_  ;
  output \g31511/_0_  ;
  output \g31512/_0_  ;
  output \g31561/_0_  ;
  output \g31603/_0_  ;
  output \g31604/_0_  ;
  output \g31666/_0_  ;
  output \g31794/_0_  ;
  output \g31795/_0_  ;
  output \g31796/_0_  ;
  output \g31854/_0_  ;
  output \g31855/_0_  ;
  output \g31856/_0_  ;
  output \g31871/_0_  ;
  output \g31920/_0_  ;
  output \g31934/_0_  ;
  output \g31935/_0_  ;
  output \g31943/_0_  ;
  output \g32128/_0_  ;
  output \g32129/_0_  ;
  output \g32130/_0_  ;
  output \g32131/_0_  ;
  output \g32132/_0_  ;
  output \g32133/_0_  ;
  output \g32134/_0_  ;
  output \g32135/_0_  ;
  output \g32136/_0_  ;
  output \g32137/_0_  ;
  output \g32140/_0_  ;
  output \g32141/_0_  ;
  output \g32142/_0_  ;
  output \g32143/_0_  ;
  output \g32144/_0_  ;
  output \g32145/_0_  ;
  output \g32146/_0_  ;
  output \g32147/_0_  ;
  output \g32475/_0_  ;
  output \g32639/_0_  ;
  output \g32640/_0_  ;
  output \g32641/_0_  ;
  output \g32642/_0_  ;
  output \g32643/_0_  ;
  output \g32644/_0_  ;
  output \g32645/_0_  ;
  output \g32646/_0_  ;
  output \g32647/_0_  ;
  output \g32648/_0_  ;
  output \g32649/_0_  ;
  output \g32650/_0_  ;
  output \g32651/_0_  ;
  output \g32652/_0_  ;
  output \g32653/_0_  ;
  output \g32654/_0_  ;
  output \g32798/_3_  ;
  output \g33177/_0_  ;
  output \g33187/_0_  ;
  output \g33306/_0_  ;
  output \g33307/_0_  ;
  output \g33308/_0_  ;
  output \g33309/_0_  ;
  output \g33310/_0_  ;
  output \g33311/_0_  ;
  output \g33312/_0_  ;
  output \g33313/_0_  ;
  output \g34088/_0_  ;
  output \g35570/_0_  ;
  output \g35594/_0_  ;
  output \g35838/_0_  ;
  output \g37467/_0_  ;
  output \g37492/_0_  ;
  output \g37503/_0_  ;
  output \g37513/_0_  ;
  output \g37524/_0_  ;
  output \g37727/_0_  ;
  output \g37748/_0_  ;
  output \g37758/_0_  ;
  output \g37767/_0_  ;
  output \g37777/_0_  ;
  output \g37790/_0_  ;
  output \g37809/_0_  ;
  output \g37840/_0_  ;
  output \g37852/_0_  ;
  output \g38312_dup/_0_  ;
  output \g38324/_0_  ;
  output \g38354/_0_  ;
  output \g38781/_1_  ;
  output \g38840/_0_  ;
  output \g38851/_0_  ;
  output \g38866/_0_  ;
  output \g38892/_1_  ;
  output \g38932/_0_  ;
  output \g38943/_0_  ;
  output \g39103/_0_  ;
  output \g39113/_2__syn_2  ;
  output \g39127/_0_  ;
  output \g44/_0_  ;
  output halt_n_pad ;
  wire n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 ;
  assign n368 = \i_tv80_core_ALU_Op_r_reg[0]/P0001  & ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  ;
  assign n369 = ~\i_tv80_core_ALU_Op_r_reg[2]/NET0131  & \i_tv80_core_ALU_Op_r_reg[3]/P0001  ;
  assign n370 = n368 & n369 ;
  assign n378 = \i_tv80_core_mcycle_reg[0]/P0001  & \i_tv80_core_mcycle_reg[1]/P0001  ;
  assign n379 = ~\i_tv80_core_mcycle_reg[0]/P0001  & ~\i_tv80_core_mcycle_reg[1]/P0001  ;
  assign n380 = ~n378 & ~n379 ;
  assign n381 = ~\i_tv80_core_mcycle_reg[2]/P0001  & n380 ;
  assign n371 = ~\i_tv80_core_IR_reg[5]/P0001  & ~\i_tv80_core_IR_reg[6]/P0001  ;
  assign n372 = ~\i_tv80_core_IR_reg[2]/P0001  & ~\i_tv80_core_IR_reg[3]/P0001  ;
  assign n373 = n371 & n372 ;
  assign n374 = ~\i_tv80_core_IR_reg[0]/P0001  & ~\i_tv80_core_IR_reg[1]/P0001  ;
  assign n375 = \i_tv80_core_IR_reg[4]/P0001  & ~\i_tv80_core_IR_reg[7]/P0001  ;
  assign n376 = n374 & n375 ;
  assign n377 = n373 & n376 ;
  assign n382 = ~\i_tv80_core_ISet_reg[0]/NET0131  & ~\i_tv80_core_ISet_reg[1]/P0001  ;
  assign n383 = n377 & n382 ;
  assign n384 = n381 & n383 ;
  assign n385 = \i_tv80_core_Save_ALU_r_reg/P0001  & ~n384 ;
  assign n386 = ~n370 & ~n385 ;
  assign n389 = ~\i_tv80_core_BusA_reg[6]/P0001  & ~\i_tv80_core_BusB_reg[6]/P0001  ;
  assign n390 = \i_tv80_core_ALU_Op_r_reg[2]/NET0131  & n368 ;
  assign n391 = \i_tv80_core_BusA_reg[6]/P0001  & \i_tv80_core_BusB_reg[6]/P0001  ;
  assign n392 = n390 & ~n391 ;
  assign n393 = ~\i_tv80_core_ALU_Op_r_reg[0]/P0001  & \i_tv80_core_ALU_Op_r_reg[2]/NET0131  ;
  assign n394 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~n391 ;
  assign n395 = n393 & ~n394 ;
  assign n396 = ~n392 & ~n395 ;
  assign n397 = ~n389 & ~n396 ;
  assign n398 = \i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~\i_tv80_core_BusB_reg[5]/P0001  ;
  assign n399 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & \i_tv80_core_BusB_reg[5]/P0001  ;
  assign n400 = ~n398 & ~n399 ;
  assign n401 = ~\i_tv80_core_BusA_reg[5]/P0001  & n400 ;
  assign n402 = \i_tv80_core_BusA_reg[5]/P0001  & ~n400 ;
  assign n403 = ~n401 & ~n402 ;
  assign n404 = \i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~\i_tv80_core_BusB_reg[4]/P0001  ;
  assign n405 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & \i_tv80_core_BusB_reg[4]/P0001  ;
  assign n406 = ~n404 & ~n405 ;
  assign n407 = \i_tv80_core_BusA_reg[4]/P0001  & ~n406 ;
  assign n408 = ~\i_tv80_core_BusA_reg[4]/P0001  & n406 ;
  assign n409 = ~n407 & ~n408 ;
  assign n410 = \i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~\i_tv80_core_BusB_reg[1]/P0001  ;
  assign n411 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & \i_tv80_core_BusB_reg[1]/P0001  ;
  assign n412 = ~n410 & ~n411 ;
  assign n413 = ~\i_tv80_core_BusA_reg[1]/P0001  & n412 ;
  assign n414 = \i_tv80_core_BusA_reg[1]/P0001  & ~n412 ;
  assign n415 = ~n413 & ~n414 ;
  assign n416 = \i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~\i_tv80_core_BusB_reg[0]/P0001  ;
  assign n417 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & \i_tv80_core_BusB_reg[0]/P0001  ;
  assign n418 = ~n416 & ~n417 ;
  assign n419 = \i_tv80_core_BusA_reg[0]/P0001  & ~n418 ;
  assign n420 = ~\i_tv80_core_BusA_reg[0]/P0001  & n418 ;
  assign n421 = ~n419 & ~n420 ;
  assign n422 = ~\i_tv80_core_ALU_Op_r_reg[2]/NET0131  & \i_tv80_core_F_reg[0]/P0001  ;
  assign n423 = \i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~n422 ;
  assign n424 = ~\i_tv80_core_ALU_Op_r_reg[0]/P0001  & ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  ;
  assign n387 = \i_tv80_core_ALU_Op_r_reg[0]/P0001  & \i_tv80_core_ALU_Op_r_reg[1]/P0001  ;
  assign n425 = ~n387 & n422 ;
  assign n426 = ~n424 & n425 ;
  assign n427 = ~n423 & ~n426 ;
  assign n428 = n421 & ~n427 ;
  assign n429 = n415 & n428 ;
  assign n430 = \i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~\i_tv80_core_BusB_reg[2]/P0001  ;
  assign n431 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & \i_tv80_core_BusB_reg[2]/P0001  ;
  assign n432 = ~n430 & ~n431 ;
  assign n433 = \i_tv80_core_BusA_reg[2]/P0001  & ~n432 ;
  assign n434 = ~\i_tv80_core_BusA_reg[2]/P0001  & n432 ;
  assign n435 = ~n433 & ~n434 ;
  assign n436 = ~n413 & n419 ;
  assign n437 = ~n414 & ~n436 ;
  assign n438 = n435 & ~n437 ;
  assign n439 = ~n435 & n437 ;
  assign n440 = ~n438 & ~n439 ;
  assign n441 = n429 & n440 ;
  assign n442 = \i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~\i_tv80_core_BusB_reg[3]/P0001  ;
  assign n443 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & \i_tv80_core_BusB_reg[3]/P0001  ;
  assign n444 = ~n442 & ~n443 ;
  assign n445 = \i_tv80_core_BusA_reg[3]/P0001  & ~n444 ;
  assign n446 = ~\i_tv80_core_BusA_reg[3]/P0001  & n444 ;
  assign n447 = ~n445 & ~n446 ;
  assign n448 = ~n434 & ~n437 ;
  assign n449 = ~n433 & ~n448 ;
  assign n450 = n447 & ~n449 ;
  assign n451 = ~n447 & n449 ;
  assign n452 = ~n450 & ~n451 ;
  assign n453 = n441 & n452 ;
  assign n454 = ~n446 & ~n449 ;
  assign n455 = ~n445 & ~n454 ;
  assign n456 = n453 & ~n455 ;
  assign n457 = ~n453 & n455 ;
  assign n458 = ~n456 & ~n457 ;
  assign n459 = n409 & n458 ;
  assign n460 = n403 & n459 ;
  assign n461 = \i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~\i_tv80_core_BusB_reg[6]/P0001  ;
  assign n462 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & \i_tv80_core_BusB_reg[6]/P0001  ;
  assign n463 = ~n461 & ~n462 ;
  assign n464 = \i_tv80_core_BusA_reg[6]/P0001  & ~n463 ;
  assign n465 = ~\i_tv80_core_BusA_reg[6]/P0001  & n463 ;
  assign n466 = ~n464 & ~n465 ;
  assign n467 = ~n401 & n407 ;
  assign n468 = ~n402 & ~n467 ;
  assign n469 = n466 & ~n468 ;
  assign n470 = ~n466 & n468 ;
  assign n471 = ~n469 & ~n470 ;
  assign n473 = n460 & n471 ;
  assign n388 = \i_tv80_core_ALU_Op_r_reg[2]/NET0131  & ~n387 ;
  assign n472 = ~n460 & ~n471 ;
  assign n474 = ~n388 & ~n472 ;
  assign n475 = ~n473 & n474 ;
  assign n476 = ~n397 & ~n475 ;
  assign n477 = ~\i_tv80_core_BusA_reg[4]/P0001  & ~\i_tv80_core_BusB_reg[4]/P0001  ;
  assign n478 = \i_tv80_core_BusA_reg[4]/P0001  & \i_tv80_core_BusB_reg[4]/P0001  ;
  assign n479 = n390 & ~n478 ;
  assign n480 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~n478 ;
  assign n481 = n393 & ~n480 ;
  assign n482 = ~n479 & ~n481 ;
  assign n483 = ~n477 & ~n482 ;
  assign n484 = ~n409 & ~n458 ;
  assign n485 = ~n388 & ~n459 ;
  assign n486 = ~n484 & n485 ;
  assign n487 = ~n483 & ~n486 ;
  assign n488 = ~n476 & ~n487 ;
  assign n489 = n476 & n487 ;
  assign n490 = ~n488 & ~n489 ;
  assign n491 = ~\i_tv80_core_BusA_reg[1]/P0001  & ~\i_tv80_core_BusB_reg[1]/P0001  ;
  assign n492 = \i_tv80_core_BusA_reg[1]/P0001  & \i_tv80_core_BusB_reg[1]/P0001  ;
  assign n493 = n390 & ~n492 ;
  assign n494 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~n492 ;
  assign n495 = n393 & ~n494 ;
  assign n496 = ~n493 & ~n495 ;
  assign n497 = ~n491 & ~n496 ;
  assign n498 = ~n419 & ~n428 ;
  assign n500 = ~n415 & n498 ;
  assign n499 = n415 & ~n498 ;
  assign n501 = ~n388 & ~n499 ;
  assign n502 = ~n500 & n501 ;
  assign n503 = ~n497 & ~n502 ;
  assign n504 = ~\i_tv80_core_BusA_reg[0]/P0001  & ~\i_tv80_core_BusB_reg[0]/P0001  ;
  assign n505 = \i_tv80_core_BusA_reg[0]/P0001  & \i_tv80_core_BusB_reg[0]/P0001  ;
  assign n506 = n390 & ~n505 ;
  assign n507 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~n505 ;
  assign n508 = n393 & ~n507 ;
  assign n509 = ~n506 & ~n508 ;
  assign n510 = ~n504 & ~n509 ;
  assign n511 = ~n421 & n427 ;
  assign n512 = ~n388 & ~n428 ;
  assign n513 = ~n511 & n512 ;
  assign n514 = ~n510 & ~n513 ;
  assign n515 = n503 & ~n514 ;
  assign n516 = ~n503 & n514 ;
  assign n517 = ~n515 & ~n516 ;
  assign n526 = ~n407 & ~n459 ;
  assign n528 = ~n403 & n526 ;
  assign n527 = n403 & ~n526 ;
  assign n529 = ~n388 & ~n527 ;
  assign n530 = ~n528 & n529 ;
  assign n518 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & n393 ;
  assign n519 = \i_tv80_core_BusA_reg[5]/P0001  & \i_tv80_core_BusB_reg[5]/P0001  ;
  assign n520 = n518 & n519 ;
  assign n521 = ~\i_tv80_core_BusA_reg[5]/P0001  & ~\i_tv80_core_BusB_reg[5]/P0001  ;
  assign n522 = \i_tv80_core_ALU_Op_r_reg[1]/P0001  & n393 ;
  assign n523 = n390 & ~n519 ;
  assign n524 = ~n522 & ~n523 ;
  assign n525 = ~n521 & ~n524 ;
  assign n531 = ~n520 & ~n525 ;
  assign n532 = ~n530 & n531 ;
  assign n533 = ~\i_tv80_core_BusA_reg[7]/P0001  & ~\i_tv80_core_BusB_reg[7]/P0001  ;
  assign n534 = \i_tv80_core_BusA_reg[7]/P0001  & \i_tv80_core_BusB_reg[7]/P0001  ;
  assign n535 = n390 & ~n534 ;
  assign n536 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~n534 ;
  assign n537 = n393 & ~n536 ;
  assign n538 = ~n535 & ~n537 ;
  assign n539 = ~n533 & ~n538 ;
  assign n540 = \i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~\i_tv80_core_BusB_reg[7]/P0001  ;
  assign n541 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & \i_tv80_core_BusB_reg[7]/P0001  ;
  assign n542 = ~n540 & ~n541 ;
  assign n543 = ~\i_tv80_core_BusA_reg[7]/P0001  & n542 ;
  assign n544 = \i_tv80_core_BusA_reg[7]/P0001  & ~n542 ;
  assign n545 = ~n543 & ~n544 ;
  assign n546 = ~n465 & ~n468 ;
  assign n547 = ~n464 & ~n546 ;
  assign n548 = ~n473 & n547 ;
  assign n549 = n473 & ~n547 ;
  assign n550 = ~n548 & ~n549 ;
  assign n552 = n545 & n550 ;
  assign n551 = ~n545 & ~n550 ;
  assign n553 = ~n388 & ~n551 ;
  assign n554 = ~n552 & n553 ;
  assign n555 = ~n539 & ~n554 ;
  assign n556 = ~\i_tv80_core_BusA_reg[3]/P0001  & ~\i_tv80_core_BusB_reg[3]/P0001  ;
  assign n557 = \i_tv80_core_BusA_reg[3]/P0001  & \i_tv80_core_BusB_reg[3]/P0001  ;
  assign n558 = n390 & ~n557 ;
  assign n559 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~n557 ;
  assign n560 = n393 & ~n559 ;
  assign n561 = ~n558 & ~n560 ;
  assign n562 = ~n556 & ~n561 ;
  assign n563 = ~n441 & ~n452 ;
  assign n564 = ~n388 & ~n453 ;
  assign n565 = ~n563 & n564 ;
  assign n566 = ~n562 & ~n565 ;
  assign n567 = n555 & ~n566 ;
  assign n568 = ~n555 & n566 ;
  assign n569 = ~n567 & ~n568 ;
  assign n570 = n532 & n569 ;
  assign n571 = ~n532 & ~n569 ;
  assign n572 = ~n570 & ~n571 ;
  assign n579 = ~n429 & ~n440 ;
  assign n580 = ~n388 & ~n441 ;
  assign n581 = ~n579 & n580 ;
  assign n573 = \i_tv80_core_BusA_reg[2]/P0001  & \i_tv80_core_BusB_reg[2]/P0001  ;
  assign n574 = n518 & n573 ;
  assign n575 = ~\i_tv80_core_BusA_reg[2]/P0001  & ~\i_tv80_core_BusB_reg[2]/P0001  ;
  assign n576 = n390 & ~n573 ;
  assign n577 = ~n522 & ~n576 ;
  assign n578 = ~n575 & ~n577 ;
  assign n582 = ~n574 & ~n578 ;
  assign n583 = ~n581 & n582 ;
  assign n584 = n572 & ~n583 ;
  assign n585 = ~n572 & n583 ;
  assign n586 = ~n584 & ~n585 ;
  assign n587 = n517 & n586 ;
  assign n588 = ~n517 & ~n586 ;
  assign n589 = ~n587 & ~n588 ;
  assign n591 = n490 & n589 ;
  assign n590 = ~n490 & ~n589 ;
  assign n592 = n388 & ~n590 ;
  assign n593 = ~n591 & n592 ;
  assign n595 = ~n543 & ~n548 ;
  assign n594 = ~n544 & n548 ;
  assign n596 = ~n388 & ~n594 ;
  assign n597 = ~n595 & n596 ;
  assign n598 = ~\i_tv80_core_Arith16_r_reg/P0001  & ~n597 ;
  assign n599 = ~n593 & n598 ;
  assign n600 = \i_tv80_core_Arith16_r_reg/P0001  & ~\i_tv80_core_F_reg[2]/P0001  ;
  assign n601 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n600 ;
  assign n602 = ~n599 & n601 ;
  assign n736 = ~\i_tv80_core_BusA_reg[1]/P0001  & ~\i_tv80_core_BusA_reg[2]/P0001  ;
  assign n737 = \i_tv80_core_BusA_reg[3]/P0001  & ~n736 ;
  assign n738 = ~\i_tv80_core_F_reg[4]/P0001  & ~n737 ;
  assign n739 = ~\i_tv80_core_BusA_reg[1]/P0001  & n738 ;
  assign n740 = \i_tv80_core_BusA_reg[1]/P0001  & ~n738 ;
  assign n741 = ~n739 & ~n740 ;
  assign n719 = ~\i_tv80_core_BusA_reg[5]/P0001  & ~\i_tv80_core_BusA_reg[6]/P0001  ;
  assign n742 = \i_tv80_core_BusA_reg[1]/P0001  & \i_tv80_core_BusA_reg[2]/P0001  ;
  assign n743 = ~\i_tv80_core_BusA_reg[3]/P0001  & ~n742 ;
  assign n744 = ~\i_tv80_core_BusA_reg[4]/P0001  & n743 ;
  assign n745 = ~n738 & n744 ;
  assign n746 = n719 & n745 ;
  assign n747 = \i_tv80_core_BusA_reg[7]/P0001  & n746 ;
  assign n748 = ~\i_tv80_core_BusA_reg[7]/P0001  & ~n746 ;
  assign n749 = ~n747 & ~n748 ;
  assign n720 = \i_tv80_core_BusA_reg[5]/P0001  & \i_tv80_core_BusA_reg[6]/P0001  ;
  assign n721 = ~n719 & ~n720 ;
  assign n750 = \i_tv80_core_BusA_reg[5]/P0001  & n745 ;
  assign n751 = ~\i_tv80_core_BusA_reg[5]/P0001  & ~n745 ;
  assign n752 = ~n750 & ~n751 ;
  assign n753 = ~n721 & n752 ;
  assign n754 = \i_tv80_core_BusA_reg[4]/P0001  & n737 ;
  assign n755 = n719 & ~n754 ;
  assign n756 = \i_tv80_core_BusA_reg[7]/P0001  & ~n755 ;
  assign n757 = ~\i_tv80_core_F_reg[0]/P0001  & ~n756 ;
  assign n758 = ~n753 & ~n757 ;
  assign n760 = n749 & n758 ;
  assign n759 = ~n749 & ~n758 ;
  assign n761 = \i_tv80_core_F_reg[1]/P0001  & ~n759 ;
  assign n762 = ~n760 & n761 ;
  assign n763 = ~\i_tv80_core_F_reg[1]/P0001  & ~n756 ;
  assign n765 = \i_tv80_core_BusA_reg[5]/P0001  & n754 ;
  assign n766 = \i_tv80_core_BusA_reg[6]/P0001  & n765 ;
  assign n764 = \i_tv80_core_F_reg[0]/P0001  & ~n755 ;
  assign n767 = ~\i_tv80_core_BusA_reg[7]/P0001  & ~n764 ;
  assign n768 = ~n766 & n767 ;
  assign n769 = n763 & ~n768 ;
  assign n770 = ~n762 & ~n769 ;
  assign n771 = n741 & ~n770 ;
  assign n772 = ~n741 & n770 ;
  assign n773 = ~n771 & ~n772 ;
  assign n774 = ~\i_tv80_core_BusA_reg[7]/P0001  & \i_tv80_core_F_reg[1]/P0001  ;
  assign n775 = ~n753 & n774 ;
  assign n776 = ~n757 & ~n763 ;
  assign n777 = ~n775 & n776 ;
  assign n778 = n773 & n777 ;
  assign n779 = ~n773 & ~n777 ;
  assign n780 = ~n778 & ~n779 ;
  assign n781 = \i_tv80_core_F_reg[4]/P0001  & n743 ;
  assign n782 = \i_tv80_core_BusA_reg[4]/P0001  & ~n781 ;
  assign n783 = ~n745 & ~n782 ;
  assign n784 = \i_tv80_core_F_reg[1]/P0001  & ~n783 ;
  assign n785 = ~\i_tv80_core_BusA_reg[4]/P0001  & ~n737 ;
  assign n786 = ~\i_tv80_core_F_reg[1]/P0001  & ~n754 ;
  assign n787 = ~n785 & n786 ;
  assign n788 = ~n784 & ~n787 ;
  assign n789 = \i_tv80_core_F_reg[1]/P0001  & ~n752 ;
  assign n790 = ~\i_tv80_core_BusA_reg[5]/P0001  & ~n754 ;
  assign n791 = ~n765 & ~n790 ;
  assign n792 = ~\i_tv80_core_F_reg[1]/P0001  & ~n791 ;
  assign n793 = ~n789 & ~n792 ;
  assign n794 = n757 & ~n793 ;
  assign n795 = ~n757 & n793 ;
  assign n796 = ~n794 & ~n795 ;
  assign n797 = n788 & ~n796 ;
  assign n798 = ~n788 & n796 ;
  assign n799 = ~n797 & ~n798 ;
  assign n800 = ~n750 & ~n757 ;
  assign n801 = ~n751 & ~n800 ;
  assign n803 = ~n721 & ~n801 ;
  assign n802 = n721 & n801 ;
  assign n804 = \i_tv80_core_F_reg[1]/P0001  & ~n802 ;
  assign n805 = ~n803 & n804 ;
  assign n806 = ~n757 & ~n791 ;
  assign n808 = ~\i_tv80_core_BusA_reg[6]/P0001  & ~n765 ;
  assign n809 = ~n766 & ~n808 ;
  assign n810 = ~n806 & ~n809 ;
  assign n807 = n721 & n806 ;
  assign n811 = ~\i_tv80_core_F_reg[1]/P0001  & ~n807 ;
  assign n812 = ~n810 & n811 ;
  assign n813 = ~n805 & ~n812 ;
  assign n814 = \i_tv80_core_F_reg[4]/P0001  & ~n736 ;
  assign n815 = ~\i_tv80_core_BusA_reg[3]/P0001  & ~n814 ;
  assign n816 = ~\i_tv80_core_F_reg[1]/P0001  & ~n737 ;
  assign n817 = ~n815 & n816 ;
  assign n818 = ~n738 & ~n742 ;
  assign n820 = \i_tv80_core_BusA_reg[3]/P0001  & n818 ;
  assign n819 = ~\i_tv80_core_BusA_reg[3]/P0001  & ~n818 ;
  assign n821 = \i_tv80_core_F_reg[1]/P0001  & ~n819 ;
  assign n822 = ~n820 & n821 ;
  assign n823 = ~n817 & ~n822 ;
  assign n824 = \i_tv80_core_BusA_reg[0]/P0001  & ~n823 ;
  assign n825 = ~\i_tv80_core_BusA_reg[0]/P0001  & n823 ;
  assign n826 = ~n824 & ~n825 ;
  assign n827 = \i_tv80_core_F_reg[1]/P0001  & ~n738 ;
  assign n828 = ~n739 & ~n827 ;
  assign n829 = ~n736 & ~n742 ;
  assign n830 = ~n828 & ~n829 ;
  assign n831 = n828 & n829 ;
  assign n832 = ~n830 & ~n831 ;
  assign n833 = n826 & n832 ;
  assign n834 = ~n826 & ~n832 ;
  assign n835 = ~n833 & ~n834 ;
  assign n836 = n813 & ~n835 ;
  assign n837 = ~n813 & n835 ;
  assign n838 = ~n836 & ~n837 ;
  assign n839 = n799 & n838 ;
  assign n840 = ~n799 & ~n838 ;
  assign n841 = ~n839 & ~n840 ;
  assign n843 = ~n780 & n841 ;
  assign n735 = \i_tv80_core_ALU_Op_r_reg[3]/P0001  & n518 ;
  assign n842 = n780 & ~n841 ;
  assign n844 = n735 & ~n842 ;
  assign n845 = ~n843 & n844 ;
  assign n605 = \i_tv80_core_BusA_reg[2]/P0001  & \i_tv80_core_IR_reg[3]/P0001  ;
  assign n606 = \i_tv80_core_BusA_reg[0]/P0001  & ~\i_tv80_core_IR_reg[3]/P0001  ;
  assign n607 = ~n605 & ~n606 ;
  assign n608 = \i_tv80_core_BusA_reg[4]/P0001  & \i_tv80_core_IR_reg[3]/P0001  ;
  assign n609 = \i_tv80_core_BusA_reg[2]/P0001  & ~\i_tv80_core_IR_reg[3]/P0001  ;
  assign n610 = ~n608 & ~n609 ;
  assign n611 = n607 & n610 ;
  assign n612 = ~n607 & ~n610 ;
  assign n613 = ~n611 & ~n612 ;
  assign n614 = ~\i_tv80_core_BusA_reg[5]/P0001  & ~\i_tv80_core_IR_reg[3]/P0001  ;
  assign n615 = ~\i_tv80_core_BusA_reg[7]/P0001  & \i_tv80_core_IR_reg[3]/P0001  ;
  assign n616 = ~n614 & ~n615 ;
  assign n617 = n613 & ~n616 ;
  assign n618 = ~n613 & n616 ;
  assign n619 = ~n617 & ~n618 ;
  assign n624 = \i_tv80_core_IR_reg[3]/P0001  & ~\i_tv80_core_IR_reg[4]/P0001  ;
  assign n625 = \i_tv80_core_IR_reg[5]/P0001  & n624 ;
  assign n626 = \i_tv80_core_BusA_reg[7]/P0001  & n625 ;
  assign n627 = \i_tv80_core_BusA_reg[0]/P0001  & \i_tv80_core_IR_reg[3]/P0001  ;
  assign n628 = ~\i_tv80_core_IR_reg[4]/P0001  & ~\i_tv80_core_IR_reg[5]/P0001  ;
  assign n629 = n627 & n628 ;
  assign n620 = \i_tv80_core_IR_reg[4]/P0001  & ~\i_tv80_core_IR_reg[5]/P0001  ;
  assign n621 = \i_tv80_core_F_reg[0]/P0001  & \i_tv80_core_IR_reg[3]/P0001  ;
  assign n622 = n620 & n621 ;
  assign n623 = \i_tv80_core_BusA_reg[6]/P0001  & ~\i_tv80_core_IR_reg[3]/P0001  ;
  assign n630 = ~n622 & ~n623 ;
  assign n631 = ~n629 & n630 ;
  assign n632 = ~n626 & n631 ;
  assign n633 = \i_tv80_core_BusA_reg[5]/P0001  & \i_tv80_core_IR_reg[3]/P0001  ;
  assign n634 = \i_tv80_core_BusA_reg[3]/P0001  & ~\i_tv80_core_IR_reg[3]/P0001  ;
  assign n635 = ~n633 & ~n634 ;
  assign n636 = \i_tv80_core_BusA_reg[6]/P0001  & \i_tv80_core_IR_reg[3]/P0001  ;
  assign n637 = \i_tv80_core_BusA_reg[4]/P0001  & ~\i_tv80_core_IR_reg[3]/P0001  ;
  assign n638 = ~n636 & ~n637 ;
  assign n639 = n635 & n638 ;
  assign n640 = ~n635 & ~n638 ;
  assign n641 = ~n639 & ~n640 ;
  assign n642 = \i_tv80_core_BusA_reg[3]/P0001  & \i_tv80_core_IR_reg[3]/P0001  ;
  assign n643 = \i_tv80_core_BusA_reg[1]/P0001  & ~\i_tv80_core_IR_reg[3]/P0001  ;
  assign n644 = ~n642 & ~n643 ;
  assign n649 = \i_tv80_core_BusA_reg[7]/P0001  & ~\i_tv80_core_IR_reg[3]/P0001  ;
  assign n650 = n628 & n649 ;
  assign n645 = ~\i_tv80_core_IR_reg[3]/P0001  & \i_tv80_core_IR_reg[4]/P0001  ;
  assign n646 = ~\i_tv80_core_F_reg[0]/P0001  & ~\i_tv80_core_IR_reg[5]/P0001  ;
  assign n647 = n645 & ~n646 ;
  assign n648 = \i_tv80_core_BusA_reg[1]/P0001  & \i_tv80_core_IR_reg[3]/P0001  ;
  assign n651 = ~n647 & ~n648 ;
  assign n652 = ~n650 & n651 ;
  assign n653 = ~n644 & ~n652 ;
  assign n654 = n644 & n652 ;
  assign n655 = ~n653 & ~n654 ;
  assign n656 = n641 & ~n655 ;
  assign n657 = ~n641 & n655 ;
  assign n658 = ~n656 & ~n657 ;
  assign n659 = n632 & n658 ;
  assign n660 = ~n632 & ~n658 ;
  assign n661 = ~n659 & ~n660 ;
  assign n663 = ~n619 & n661 ;
  assign n662 = n619 & ~n661 ;
  assign n664 = ~n382 & ~n662 ;
  assign n665 = ~n663 & n664 ;
  assign n603 = ~\i_tv80_core_F_reg[2]/P0001  & n382 ;
  assign n604 = n369 & n424 ;
  assign n666 = ~n603 & n604 ;
  assign n667 = ~n665 & n666 ;
  assign n701 = \i_tv80_core_ALU_Op_r_reg[0]/P0001  & \i_tv80_core_BusB_reg[4]/P0001  ;
  assign n702 = ~\i_tv80_core_ALU_Op_r_reg[0]/P0001  & \i_tv80_core_BusB_reg[0]/P0001  ;
  assign n703 = ~n701 & ~n702 ;
  assign n704 = ~\i_tv80_core_BusA_reg[4]/P0001  & ~\i_tv80_core_BusA_reg[7]/P0001  ;
  assign n705 = \i_tv80_core_BusA_reg[4]/P0001  & \i_tv80_core_BusA_reg[7]/P0001  ;
  assign n706 = ~n704 & ~n705 ;
  assign n707 = \i_tv80_core_ALU_Op_r_reg[0]/P0001  & \i_tv80_core_BusB_reg[6]/P0001  ;
  assign n708 = ~\i_tv80_core_ALU_Op_r_reg[0]/P0001  & \i_tv80_core_BusB_reg[2]/P0001  ;
  assign n709 = ~n707 & ~n708 ;
  assign n710 = n706 & ~n709 ;
  assign n711 = ~n706 & n709 ;
  assign n712 = ~n710 & ~n711 ;
  assign n713 = n703 & n712 ;
  assign n714 = ~n703 & ~n712 ;
  assign n715 = ~n713 & ~n714 ;
  assign n716 = \i_tv80_core_ALU_Op_r_reg[0]/P0001  & \i_tv80_core_BusB_reg[5]/P0001  ;
  assign n717 = ~\i_tv80_core_ALU_Op_r_reg[0]/P0001  & \i_tv80_core_BusB_reg[1]/P0001  ;
  assign n718 = ~n716 & ~n717 ;
  assign n722 = \i_tv80_core_ALU_Op_r_reg[0]/P0001  & \i_tv80_core_BusB_reg[7]/P0001  ;
  assign n723 = ~\i_tv80_core_ALU_Op_r_reg[0]/P0001  & \i_tv80_core_BusB_reg[3]/P0001  ;
  assign n724 = ~n722 & ~n723 ;
  assign n725 = n721 & ~n724 ;
  assign n726 = ~n721 & n724 ;
  assign n727 = ~n725 & ~n726 ;
  assign n728 = n718 & n727 ;
  assign n729 = ~n718 & ~n727 ;
  assign n730 = ~n728 & ~n729 ;
  assign n732 = n715 & ~n730 ;
  assign n699 = \i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n424 ;
  assign n700 = n388 & n699 ;
  assign n731 = ~n715 & n730 ;
  assign n733 = n700 & ~n731 ;
  assign n734 = ~n732 & n733 ;
  assign n686 = ~\i_tv80_core_IR_reg[5]/P0001  & n624 ;
  assign n687 = \i_tv80_core_BusB_reg[1]/P0001  & n686 ;
  assign n681 = ~\i_tv80_core_IR_reg[4]/P0001  & \i_tv80_core_IR_reg[5]/P0001  ;
  assign n682 = \i_tv80_core_IR_reg[3]/P0001  & n681 ;
  assign n683 = \i_tv80_core_BusB_reg[5]/P0001  & n682 ;
  assign n668 = ~\i_tv80_core_IR_reg[3]/P0001  & ~\i_tv80_core_IR_reg[4]/P0001  ;
  assign n684 = ~\i_tv80_core_IR_reg[5]/P0001  & n668 ;
  assign n685 = \i_tv80_core_BusB_reg[0]/P0001  & n684 ;
  assign n691 = ~n683 & ~n685 ;
  assign n692 = ~n687 & n691 ;
  assign n669 = \i_tv80_core_IR_reg[5]/P0001  & n668 ;
  assign n670 = \i_tv80_core_BusB_reg[4]/P0001  & n669 ;
  assign n688 = n370 & ~n670 ;
  assign n671 = ~\i_tv80_core_IR_reg[5]/P0001  & n645 ;
  assign n672 = \i_tv80_core_BusB_reg[2]/P0001  & n671 ;
  assign n673 = \i_tv80_core_IR_reg[5]/P0001  & n645 ;
  assign n674 = \i_tv80_core_BusB_reg[6]/P0001  & n673 ;
  assign n689 = ~n672 & ~n674 ;
  assign n675 = \i_tv80_core_IR_reg[4]/P0001  & \i_tv80_core_IR_reg[5]/P0001  ;
  assign n676 = \i_tv80_core_IR_reg[3]/P0001  & n675 ;
  assign n677 = \i_tv80_core_BusB_reg[7]/P0001  & n676 ;
  assign n678 = \i_tv80_core_IR_reg[3]/P0001  & \i_tv80_core_IR_reg[4]/P0001  ;
  assign n679 = ~\i_tv80_core_IR_reg[5]/P0001  & n678 ;
  assign n680 = \i_tv80_core_BusB_reg[3]/P0001  & n679 ;
  assign n690 = ~n677 & ~n680 ;
  assign n693 = n689 & n690 ;
  assign n694 = n688 & n693 ;
  assign n695 = n692 & n694 ;
  assign n696 = \i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~n393 ;
  assign n697 = \i_tv80_core_ALU_Op_r_reg[3]/P0001  & n696 ;
  assign n698 = \i_tv80_core_F_reg[2]/P0001  & n697 ;
  assign n846 = ~n695 & ~n698 ;
  assign n847 = ~n734 & n846 ;
  assign n848 = ~n667 & n847 ;
  assign n849 = ~n845 & n848 ;
  assign n850 = ~n602 & n849 ;
  assign n851 = ~n386 & ~n850 ;
  assign n859 = \i_tv80_core_mcycle_reg[0]/P0001  & ~\i_tv80_core_mcycle_reg[2]/P0001  ;
  assign n860 = ~\i_tv80_core_mcycle_reg[1]/P0001  & n859 ;
  assign n861 = ~\i_tv80_core_mcycle_reg[0]/P0001  & \i_tv80_core_mcycle_reg[1]/P0001  ;
  assign n862 = \i_tv80_core_mcycle_reg[2]/P0001  & n861 ;
  assign n863 = ~n860 & ~n862 ;
  assign n856 = \i_tv80_core_mcycle_reg[1]/P0001  & ~\i_tv80_core_mcycle_reg[2]/P0001  ;
  assign n956 = \i_tv80_core_mcycle_reg[0]/P0001  & n856 ;
  assign n960 = ~\i_tv80_core_F_reg[0]/P0001  & n671 ;
  assign n961 = \i_tv80_core_F_reg[7]/P0001  & n676 ;
  assign n966 = ~n960 & ~n961 ;
  assign n962 = \i_tv80_core_F_reg[6]/P0001  & n686 ;
  assign n963 = ~\i_tv80_core_F_reg[6]/P0001  & n684 ;
  assign n967 = ~n962 & ~n963 ;
  assign n968 = n966 & n967 ;
  assign n957 = ~\i_tv80_core_F_reg[2]/P0001  & n669 ;
  assign n964 = ~n622 & ~n957 ;
  assign n958 = ~\i_tv80_core_F_reg[7]/P0001  & n673 ;
  assign n959 = \i_tv80_core_F_reg[2]/P0001  & n625 ;
  assign n965 = ~n958 & ~n959 ;
  assign n969 = n964 & n965 ;
  assign n970 = n968 & n969 ;
  assign n971 = n956 & n970 ;
  assign n972 = n859 & ~n971 ;
  assign n885 = ~\i_tv80_core_IR_reg[0]/P0001  & \i_tv80_core_IR_reg[2]/P0001  ;
  assign n867 = \i_tv80_core_IR_reg[6]/P0001  & \i_tv80_core_IR_reg[7]/P0001  ;
  assign n973 = ~\i_tv80_core_IR_reg[1]/P0001  & n867 ;
  assign n974 = n885 & n973 ;
  assign n975 = ~n972 & n974 ;
  assign n912 = \i_tv80_core_IR_reg[0]/P0001  & \i_tv80_core_IR_reg[3]/P0001  ;
  assign n853 = ~\i_tv80_core_IR_reg[1]/P0001  & ~\i_tv80_core_IR_reg[2]/P0001  ;
  assign n913 = ~\i_tv80_core_IR_reg[6]/P0001  & ~\i_tv80_core_IR_reg[7]/P0001  ;
  assign n914 = n853 & n913 ;
  assign n915 = n912 & n914 ;
  assign n916 = \i_tv80_core_IR_reg[2]/P0001  & ~\i_tv80_core_IR_reg[3]/P0001  ;
  assign n917 = ~\i_tv80_core_IR_reg[7]/P0001  & n675 ;
  assign n918 = ~\i_tv80_core_IR_reg[6]/P0001  & n917 ;
  assign n919 = n916 & n918 ;
  assign n920 = ~\i_tv80_core_IR_reg[1]/P0001  & n919 ;
  assign n921 = \i_tv80_core_IR_reg[0]/P0001  & n920 ;
  assign n922 = ~n915 & ~n921 ;
  assign n923 = ~n381 & ~n922 ;
  assign n891 = ~\i_tv80_core_IR_reg[2]/P0001  & \i_tv80_core_IR_reg[5]/P0001  ;
  assign n892 = ~\i_tv80_core_IR_reg[6]/P0001  & n891 ;
  assign n893 = ~\i_tv80_core_IR_reg[3]/P0001  & n892 ;
  assign n889 = ~\i_tv80_core_IR_reg[0]/P0001  & \i_tv80_core_IR_reg[1]/P0001  ;
  assign n895 = ~\i_tv80_core_IR_reg[4]/P0001  & ~\i_tv80_core_IR_reg[7]/P0001  ;
  assign n896 = n889 & n895 ;
  assign n910 = n893 & n896 ;
  assign n911 = ~n860 & n910 ;
  assign n924 = ~\i_tv80_core_IR_reg[0]/P0001  & ~n381 ;
  assign n925 = n920 & n924 ;
  assign n926 = ~n911 & ~n925 ;
  assign n927 = ~n923 & n926 ;
  assign n874 = ~\i_tv80_core_IR_reg[2]/P0001  & \i_tv80_core_IR_reg[3]/P0001  ;
  assign n1075 = n371 & n874 ;
  assign n1076 = n896 & n1075 ;
  assign n1077 = ~n860 & n1076 ;
  assign n904 = \i_tv80_core_IR_reg[1]/P0001  & ~\i_tv80_core_IR_reg[6]/P0001  ;
  assign n1013 = \i_tv80_core_IR_reg[0]/P0001  & ~\i_tv80_core_IR_reg[7]/P0001  ;
  assign n1063 = ~\i_tv80_core_IR_reg[2]/P0001  & n1013 ;
  assign n1064 = n904 & n1063 ;
  assign n1078 = ~\i_tv80_core_IR_reg[3]/P0001  & n1064 ;
  assign n1079 = ~n1077 & ~n1078 ;
  assign n886 = \i_tv80_core_IR_reg[1]/P0001  & n885 ;
  assign n952 = ~\i_tv80_core_IR_reg[3]/P0001  & n917 ;
  assign n953 = \i_tv80_core_IR_reg[6]/P0001  & n952 ;
  assign n1080 = ~n886 & n953 ;
  assign n1081 = ~n860 & n1080 ;
  assign n1082 = n1079 & ~n1081 ;
  assign n876 = \i_tv80_core_IR_reg[0]/P0001  & \i_tv80_core_IR_reg[1]/P0001  ;
  assign n943 = ~\i_tv80_core_IR_reg[2]/P0001  & n867 ;
  assign n1066 = n876 & n943 ;
  assign n1067 = n673 & n1066 ;
  assign n852 = ~\i_tv80_core_IR_reg[0]/P0001  & ~\i_tv80_core_IR_reg[7]/P0001  ;
  assign n1028 = \i_tv80_core_IR_reg[1]/P0001  & \i_tv80_core_IR_reg[2]/P0001  ;
  assign n1068 = n852 & n1028 ;
  assign n1069 = ~n673 & n1068 ;
  assign n882 = ~\i_tv80_core_IR_reg[4]/P0001  & \i_tv80_core_IR_reg[7]/P0001  ;
  assign n883 = n876 & n882 ;
  assign n873 = ~\i_tv80_core_IR_reg[5]/P0001  & \i_tv80_core_IR_reg[6]/P0001  ;
  assign n1070 = n372 & n873 ;
  assign n1071 = n883 & n1070 ;
  assign n1072 = ~n1069 & ~n1071 ;
  assign n1073 = ~n1067 & n1072 ;
  assign n1074 = ~n860 & ~n1073 ;
  assign n928 = n374 & n895 ;
  assign n929 = n373 & n928 ;
  assign n930 = ~\i_tv80_core_IntCycle_reg/P0001  & ~\i_tv80_core_NMICycle_reg/P0001  ;
  assign n931 = \i_tv80_core_mcycle_reg[1]/P0001  & n930 ;
  assign n1083 = ~\i_tv80_core_mcycle_reg[2]/P0001  & ~n379 ;
  assign n1084 = ~n931 & n1083 ;
  assign n1085 = n929 & ~n1084 ;
  assign n1065 = \i_tv80_core_IR_reg[3]/P0001  & n1064 ;
  assign n880 = \i_tv80_core_IR_reg[5]/P0001  & \i_tv80_core_IR_reg[6]/P0001  ;
  assign n881 = n874 & n880 ;
  assign n877 = \i_tv80_core_IR_reg[4]/P0001  & \i_tv80_core_IR_reg[7]/P0001  ;
  assign n940 = \i_tv80_core_IR_reg[0]/P0001  & ~\i_tv80_core_IR_reg[1]/P0001  ;
  assign n1086 = n877 & n940 ;
  assign n1087 = n881 & n1086 ;
  assign n1088 = ~n1065 & ~n1087 ;
  assign n1089 = ~n1085 & n1088 ;
  assign n1090 = ~n1074 & n1089 ;
  assign n1091 = n1082 & n1090 ;
  assign n1092 = n927 & n1091 ;
  assign n1093 = ~n975 & n1092 ;
  assign n1094 = ~\i_tv80_core_ISet_reg[0]/NET0131  & ~n1093 ;
  assign n1095 = ~\i_tv80_core_ISet_reg[1]/P0001  & ~n1094 ;
  assign n936 = \i_tv80_core_IR_reg[2]/P0001  & \i_tv80_core_IR_reg[6]/P0001  ;
  assign n997 = n876 & n895 ;
  assign n998 = n936 & n997 ;
  assign n1034 = \i_tv80_core_IR_reg[5]/P0001  & n998 ;
  assign n1035 = ~n859 & n1034 ;
  assign n946 = ~\i_tv80_core_IR_reg[1]/P0001  & n936 ;
  assign n1042 = n852 & n946 ;
  assign n989 = \i_tv80_core_IR_reg[6]/P0001  & ~\i_tv80_core_IR_reg[7]/P0001  ;
  assign n1036 = n853 & n989 ;
  assign n1037 = n896 & n936 ;
  assign n1043 = ~n1036 & ~n1037 ;
  assign n1044 = ~n1042 & n1043 ;
  assign n1026 = ~\i_tv80_core_IR_reg[3]/P0001  & \i_tv80_core_IR_reg[5]/P0001  ;
  assign n1027 = \i_tv80_core_IR_reg[0]/P0001  & ~n1026 ;
  assign n1031 = ~n1027 & n1028 ;
  assign n1029 = \i_tv80_core_IR_reg[6]/P0001  & n375 ;
  assign n999 = \i_tv80_core_IR_reg[3]/P0001  & ~\i_tv80_core_IR_reg[5]/P0001  ;
  assign n1030 = ~\i_tv80_core_IR_reg[0]/P0001  & ~n999 ;
  assign n1032 = n1029 & ~n1030 ;
  assign n1033 = n1031 & n1032 ;
  assign n1038 = n889 & n916 ;
  assign n1039 = n1029 & n1038 ;
  assign n990 = n876 & n989 ;
  assign n1040 = n874 & n990 ;
  assign n1041 = ~n1039 & ~n1040 ;
  assign n1045 = ~n1033 & n1041 ;
  assign n1046 = n1044 & n1045 ;
  assign n1047 = ~n1035 & n1046 ;
  assign n1048 = ~n860 & ~n1047 ;
  assign n993 = \i_tv80_core_IR_reg[1]/P0001  & \i_tv80_core_IR_reg[6]/P0001  ;
  assign n1049 = ~\i_tv80_core_IR_reg[2]/P0001  & n993 ;
  assign n1050 = n852 & n1049 ;
  assign n1051 = ~n381 & n1050 ;
  assign n1052 = \i_tv80_core_ISet_reg[1]/P0001  & ~n1051 ;
  assign n1053 = ~n1048 & n1052 ;
  assign n1096 = ~n862 & ~n1053 ;
  assign n1097 = ~n1095 & n1096 ;
  assign n1098 = ~n863 & ~n1097 ;
  assign n1099 = \i_tv80_core_tstate_reg[1]/NET0131  & ~n1098 ;
  assign n1100 = ~\i_tv80_core_tstate_reg[1]/NET0131  & n1098 ;
  assign n1101 = ~n1099 & ~n1100 ;
  assign n864 = \i_tv80_core_tstate_reg[2]/NET0131  & ~n863 ;
  assign n865 = ~\i_tv80_core_tstate_reg[2]/NET0131  & n863 ;
  assign n866 = ~n864 & ~n865 ;
  assign n884 = n881 & n883 ;
  assign n887 = n867 & n886 ;
  assign n888 = ~n884 & ~n887 ;
  assign n890 = n375 & n889 ;
  assign n894 = n890 & n893 ;
  assign n897 = \i_tv80_core_IR_reg[3]/P0001  & n892 ;
  assign n898 = n896 & n897 ;
  assign n899 = ~n894 & ~n898 ;
  assign n900 = n888 & n899 ;
  assign n868 = ~\i_tv80_core_IR_reg[1]/P0001  & \i_tv80_core_IR_reg[2]/P0001  ;
  assign n869 = n867 & n868 ;
  assign n870 = n686 & n869 ;
  assign n871 = \i_tv80_core_IR_reg[0]/P0001  & n870 ;
  assign n872 = ~n859 & n871 ;
  assign n875 = n873 & n874 ;
  assign n878 = n876 & n877 ;
  assign n879 = n875 & n878 ;
  assign n901 = \i_tv80_core_IR_reg[2]/P0001  & ~\i_tv80_core_IR_reg[7]/P0001  ;
  assign n902 = \i_tv80_core_IR_reg[0]/P0001  & ~\i_tv80_core_IR_reg[5]/P0001  ;
  assign n903 = n901 & n902 ;
  assign n905 = n903 & n904 ;
  assign n906 = ~n879 & ~n905 ;
  assign n907 = ~n872 & n906 ;
  assign n908 = n900 & n907 ;
  assign n909 = ~n860 & ~n908 ;
  assign n950 = ~n860 & ~n886 ;
  assign n951 = ~\i_tv80_core_IR_reg[6]/P0001  & \i_tv80_core_IR_reg[7]/P0001  ;
  assign n954 = ~n951 & ~n953 ;
  assign n955 = n950 & ~n954 ;
  assign n932 = n859 & n930 ;
  assign n933 = ~n856 & ~n932 ;
  assign n934 = ~n931 & ~n933 ;
  assign n935 = n929 & ~n934 ;
  assign n937 = \i_tv80_core_IR_reg[1]/P0001  & n936 ;
  assign n938 = \i_tv80_core_IR_reg[0]/P0001  & \i_tv80_core_IR_reg[7]/P0001  ;
  assign n939 = n937 & n938 ;
  assign n979 = ~n377 & ~n939 ;
  assign n980 = ~n935 & n979 ;
  assign n941 = n882 & n940 ;
  assign n942 = n875 & n941 ;
  assign n944 = n374 & n943 ;
  assign n945 = ~n942 & ~n944 ;
  assign n947 = ~\i_tv80_core_IR_reg[3]/P0001  & n938 ;
  assign n948 = n946 & n947 ;
  assign n949 = n945 & ~n948 ;
  assign n976 = n372 & n883 ;
  assign n977 = n880 & n976 ;
  assign n978 = ~n859 & n977 ;
  assign n981 = n949 & ~n978 ;
  assign n982 = n980 & n981 ;
  assign n983 = ~n955 & n982 ;
  assign n984 = ~n909 & n983 ;
  assign n985 = n927 & n984 ;
  assign n986 = ~n975 & n985 ;
  assign n987 = ~\i_tv80_core_ISet_reg[0]/NET0131  & ~n986 ;
  assign n988 = ~\i_tv80_core_ISet_reg[1]/P0001  & ~n987 ;
  assign n1005 = \i_tv80_core_IR_reg[7]/P0001  & n892 ;
  assign n1006 = \i_tv80_core_IR_reg[1]/P0001  & n1005 ;
  assign n1020 = ~\i_tv80_core_IR_reg[0]/P0001  & n1006 ;
  assign n1021 = ~n859 & n1020 ;
  assign n1008 = n372 & n990 ;
  assign n1009 = ~\i_tv80_core_IR_reg[7]/P0001  & n676 ;
  assign n1010 = n937 & n1009 ;
  assign n1011 = ~n1008 & ~n1010 ;
  assign n1012 = ~\i_tv80_core_IR_reg[1]/P0001  & n1005 ;
  assign n1014 = n946 & n1013 ;
  assign n1015 = ~n951 & ~n989 ;
  assign n1016 = \i_tv80_core_IR_reg[2]/P0001  & ~\i_tv80_core_IR_reg[6]/P0001  ;
  assign n1017 = ~n371 & ~n1016 ;
  assign n1018 = ~n1015 & n1017 ;
  assign n1019 = ~n1014 & n1018 ;
  assign n1022 = ~n1012 & n1019 ;
  assign n1023 = n1011 & n1022 ;
  assign n1024 = ~n1021 & n1023 ;
  assign n1025 = ~n860 & ~n1024 ;
  assign n991 = \i_tv80_core_IR_reg[2]/P0001  & n671 ;
  assign n992 = n990 & n991 ;
  assign n994 = n678 & n993 ;
  assign n995 = n903 & n994 ;
  assign n996 = ~n992 & ~n995 ;
  assign n1000 = n998 & n999 ;
  assign n1001 = n873 & n916 ;
  assign n1002 = n997 & n1001 ;
  assign n1003 = ~n1000 & ~n1002 ;
  assign n1004 = n996 & n1003 ;
  assign n1007 = \i_tv80_core_IR_reg[0]/P0001  & n1006 ;
  assign n1054 = n1004 & ~n1007 ;
  assign n1055 = ~n1025 & n1054 ;
  assign n1056 = n1053 & n1055 ;
  assign n1057 = ~n862 & ~n1056 ;
  assign n1058 = ~n988 & n1057 ;
  assign n1059 = ~n863 & ~n1058 ;
  assign n1060 = \i_tv80_core_tstate_reg[0]/P0001  & ~n1059 ;
  assign n1061 = ~\i_tv80_core_tstate_reg[0]/P0001  & n1059 ;
  assign n1062 = ~n1060 & ~n1061 ;
  assign n1102 = ~n866 & ~n1062 ;
  assign n1103 = ~n1101 & n1102 ;
  assign n854 = \i_tv80_core_IR_reg[6]/P0001  & n853 ;
  assign n855 = n852 & n854 ;
  assign n857 = ~\i_tv80_core_mcycle_reg[0]/P0001  & n856 ;
  assign n858 = \i_tv80_core_ISet_reg[1]/P0001  & n857 ;
  assign n1104 = n855 & n858 ;
  assign n1105 = n1103 & n1104 ;
  assign n1106 = \i_tv80_core_tstate_reg[0]/P0001  & \i_tv80_core_tstate_reg[1]/NET0131  ;
  assign n1107 = ~\i_tv80_core_tstate_reg[2]/NET0131  & n1106 ;
  assign n1108 = \i_tv80_core_ISet_reg[1]/P0001  & n989 ;
  assign n1109 = n902 & n1028 ;
  assign n1110 = n1108 & n1109 ;
  assign n1111 = n1107 & n1110 ;
  assign n1112 = \i_tv80_core_IR_reg[4]/P0001  & n1111 ;
  assign n1113 = ~\i_tv80_core_tstate_reg[2]/NET0131  & n860 ;
  assign n1114 = ~\i_tv80_core_IR_reg[6]/P0001  & n853 ;
  assign n1115 = n382 & n852 ;
  assign n1116 = n686 & n1115 ;
  assign n1117 = n1114 & n1116 ;
  assign n1118 = ~n1113 & n1117 ;
  assign n1119 = ~\i_tv80_core_F_reg[2]/P0001  & ~n1118 ;
  assign n1120 = ~\i_tv80_core_Fp_reg[2]/P0001  & n1118 ;
  assign n1121 = ~n1119 & ~n1120 ;
  assign n1122 = ~n1112 & ~n1121 ;
  assign n1123 = ~\i_tv80_core_IntE_FF2_reg/P0001  & n1112 ;
  assign n1124 = n386 & ~n1123 ;
  assign n1125 = ~n1122 & n1124 ;
  assign n1126 = ~n1105 & ~n1125 ;
  assign n1127 = ~n851 & n1126 ;
  assign n1128 = \i_tv80_core_ISet_reg[1]/P0001  & n956 ;
  assign n1129 = n1012 & n1128 ;
  assign n1130 = ~\di_reg_reg[0]/P0001  & ~\di_reg_reg[7]/P0001  ;
  assign n1131 = \di_reg_reg[0]/P0001  & \di_reg_reg[7]/P0001  ;
  assign n1132 = ~n1130 & ~n1131 ;
  assign n1133 = ~\di_reg_reg[3]/P0001  & ~\di_reg_reg[5]/P0001  ;
  assign n1134 = \di_reg_reg[3]/P0001  & \di_reg_reg[5]/P0001  ;
  assign n1135 = ~n1133 & ~n1134 ;
  assign n1136 = n1132 & ~n1135 ;
  assign n1137 = ~n1132 & n1135 ;
  assign n1138 = ~n1136 & ~n1137 ;
  assign n1139 = ~\di_reg_reg[1]/P0001  & ~\di_reg_reg[6]/P0001  ;
  assign n1140 = \di_reg_reg[1]/P0001  & \di_reg_reg[6]/P0001  ;
  assign n1141 = ~n1139 & ~n1140 ;
  assign n1142 = ~\di_reg_reg[2]/P0001  & ~\di_reg_reg[4]/P0001  ;
  assign n1143 = \di_reg_reg[2]/P0001  & \di_reg_reg[4]/P0001  ;
  assign n1144 = ~n1142 & ~n1143 ;
  assign n1145 = n1141 & ~n1144 ;
  assign n1146 = ~n1141 & n1144 ;
  assign n1147 = ~n1145 & ~n1146 ;
  assign n1148 = n1138 & n1147 ;
  assign n1149 = ~n1138 & ~n1147 ;
  assign n1150 = ~n1148 & ~n1149 ;
  assign n1151 = n1105 & n1150 ;
  assign n1152 = ~n1129 & ~n1151 ;
  assign n1153 = ~n1127 & n1152 ;
  assign n1154 = \i_tv80_core_IncDecZ_reg/P0002  & n1129 ;
  assign n1155 = \i_tv80_core_tstate_reg[0]/P0001  & ~\i_tv80_core_tstate_reg[1]/NET0131  ;
  assign n1156 = ~\i_tv80_core_tstate_reg[2]/NET0131  & n1155 ;
  assign n1157 = ~\i_tv80_core_Auto_Wait_t1_reg/P0001  & n1156 ;
  assign n1158 = ~\i_tv80_core_Save_ALU_r_reg/P0001  & ~n1157 ;
  assign n1159 = \i_tv80_core_ALU_Op_r_reg[2]/NET0131  & n387 ;
  assign n1160 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & \i_tv80_core_Save_ALU_r_reg/P0001  ;
  assign n1161 = n1159 & n1160 ;
  assign n1162 = ~n1158 & ~n1161 ;
  assign n1163 = \i_tv80_core_Read_To_Reg_r_reg[3]/P0001  & \i_tv80_core_Read_To_Reg_r_reg[4]/P0001  ;
  assign n1164 = n1162 & n1163 ;
  assign n1165 = \i_tv80_core_Read_To_Reg_r_reg[0]/P0001  & \i_tv80_core_Read_To_Reg_r_reg[1]/P0001  ;
  assign n1166 = ~\i_tv80_core_Read_To_Reg_r_reg[2]/P0001  & n1165 ;
  assign n1167 = n1164 & n1166 ;
  assign n1168 = ~n1154 & ~n1167 ;
  assign n1169 = ~n1153 & n1168 ;
  assign n1183 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n583 ;
  assign n1174 = n735 & n832 ;
  assign n1177 = \i_tv80_core_ALU_Op_r_reg[0]/P0001  & n671 ;
  assign n1175 = \i_tv80_core_ALU_Op_r_reg[1]/P0001  & n369 ;
  assign n1176 = ~\i_tv80_core_BusB_reg[2]/P0001  & ~n671 ;
  assign n1178 = n1175 & ~n1176 ;
  assign n1179 = ~n1177 & n1178 ;
  assign n1181 = n700 & ~n709 ;
  assign n1180 = n370 & n672 ;
  assign n1182 = n604 & ~n644 ;
  assign n1184 = \i_tv80_core_Save_ALU_r_reg/P0001  & ~n1182 ;
  assign n1185 = ~n1180 & n1184 ;
  assign n1186 = ~n1181 & n1185 ;
  assign n1187 = ~n1179 & n1186 ;
  assign n1188 = ~n1174 & n1187 ;
  assign n1189 = ~n1183 & n1188 ;
  assign n1170 = ~n886 & n989 ;
  assign n1171 = ~n673 & n1170 ;
  assign n1172 = n382 & n1171 ;
  assign n1173 = ~\di_reg_reg[2]/P0001  & ~\i_tv80_core_Save_ALU_r_reg/P0001  ;
  assign n1190 = ~n1172 & ~n1173 ;
  assign n1191 = ~n1189 & n1190 ;
  assign n1192 = \i_tv80_core_BusB_reg[2]/P0001  & n1172 ;
  assign n1193 = ~n1191 & ~n1192 ;
  assign n1194 = n1167 & n1193 ;
  assign n1195 = ~\i_tv80_core_BusAck_reg/P0001  & ~n1194 ;
  assign n1196 = ~n1169 & n1195 ;
  assign n1197 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_F_reg[2]/P0001  ;
  assign n1198 = reset_n_pad & ~n1197 ;
  assign n1199 = ~n1196 & n1198 ;
  assign n1222 = \i_tv80_core_Arith16_r_reg/P0001  & \i_tv80_core_F_reg[6]/P0001  ;
  assign n1223 = ~\i_tv80_core_F_reg[6]/P0001  & \i_tv80_core_Z16_r_reg/P0001  ;
  assign n1224 = ~\i_tv80_core_Arith16_r_reg/P0001  & ~n1223 ;
  assign n1225 = n514 & n1224 ;
  assign n1226 = n503 & n1225 ;
  assign n1227 = n583 & n1226 ;
  assign n1228 = n566 & n1227 ;
  assign n1229 = n532 & n1228 ;
  assign n1230 = n489 & n1229 ;
  assign n1231 = n555 & n1230 ;
  assign n1232 = ~n1222 & ~n1231 ;
  assign n1233 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n1232 ;
  assign n1249 = n735 & ~n832 ;
  assign n1250 = n825 & n1249 ;
  assign n1251 = n797 & n1250 ;
  assign n1252 = n813 & n1251 ;
  assign n1253 = n772 & n1252 ;
  assign n1234 = \i_tv80_core_F_reg[6]/P0001  & n382 ;
  assign n1235 = ~n382 & n632 ;
  assign n1236 = n611 & ~n616 ;
  assign n1237 = n639 & n1236 ;
  assign n1238 = n654 & n1237 ;
  assign n1239 = n1235 & n1238 ;
  assign n1240 = ~n1234 & ~n1239 ;
  assign n1241 = n604 & ~n1240 ;
  assign n1244 = n709 & n718 ;
  assign n1245 = n724 & n1244 ;
  assign n1242 = n704 & n719 ;
  assign n1243 = n703 & n1242 ;
  assign n1246 = n700 & n1243 ;
  assign n1247 = n1245 & n1246 ;
  assign n1248 = \i_tv80_core_F_reg[6]/P0001  & n697 ;
  assign n1254 = ~n1247 & ~n1248 ;
  assign n1255 = ~n695 & n1254 ;
  assign n1256 = ~n1241 & n1255 ;
  assign n1257 = ~n1253 & n1256 ;
  assign n1258 = ~n1233 & n1257 ;
  assign n1259 = ~n386 & ~n1258 ;
  assign n1260 = \i_tv80_core_Fp_reg[6]/P0001  & n1118 ;
  assign n1261 = \i_tv80_core_F_reg[6]/P0001  & ~n1118 ;
  assign n1262 = ~n1260 & ~n1261 ;
  assign n1263 = n386 & ~n1262 ;
  assign n1264 = ~n1105 & ~n1263 ;
  assign n1265 = ~n1259 & n1264 ;
  assign n1266 = n1130 & n1133 ;
  assign n1267 = n1139 & n1142 ;
  assign n1268 = n1266 & n1267 ;
  assign n1269 = n1105 & ~n1268 ;
  assign n1270 = ~n1265 & ~n1269 ;
  assign n1271 = ~n1167 & ~n1270 ;
  assign n1210 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n476 ;
  assign n1202 = n735 & ~n813 ;
  assign n1204 = \i_tv80_core_ALU_Op_r_reg[0]/P0001  & n673 ;
  assign n1203 = ~\i_tv80_core_BusB_reg[6]/P0001  & ~n673 ;
  assign n1205 = n1175 & ~n1203 ;
  assign n1206 = ~n1204 & n1205 ;
  assign n1208 = n370 & n674 ;
  assign n1207 = \i_tv80_core_BusA_reg[6]/P0001  & n700 ;
  assign n1209 = n604 & n616 ;
  assign n1211 = \i_tv80_core_Save_ALU_r_reg/P0001  & ~n1209 ;
  assign n1212 = ~n1207 & n1211 ;
  assign n1213 = ~n1208 & n1212 ;
  assign n1214 = ~n1206 & n1213 ;
  assign n1215 = ~n1202 & n1214 ;
  assign n1216 = ~n1210 & n1215 ;
  assign n1201 = ~\di_reg_reg[6]/P0001  & ~\i_tv80_core_Save_ALU_r_reg/P0001  ;
  assign n1217 = ~n1172 & ~n1201 ;
  assign n1218 = ~n1216 & n1217 ;
  assign n1219 = \i_tv80_core_BusB_reg[6]/P0001  & n1172 ;
  assign n1220 = ~n1218 & ~n1219 ;
  assign n1221 = n1167 & n1220 ;
  assign n1272 = ~\i_tv80_core_BusAck_reg/P0001  & ~n1221 ;
  assign n1273 = ~n1271 & n1272 ;
  assign n1200 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_F_reg[6]/P0001  ;
  assign n1274 = reset_n_pad & ~n1200 ;
  assign n1275 = ~n1273 & n1274 ;
  assign n1276 = n881 & n941 ;
  assign n1277 = n382 & n1276 ;
  assign n1289 = \i_tv80_core_RegAddrC_reg[1]/NET0131  & ~\i_tv80_core_RegAddrC_reg[2]/NET0131  ;
  assign n1290 = ~\i_tv80_core_RegAddrC_reg[0]/P0001  & n1289 ;
  assign n1291 = \i_tv80_core_i_reg_RegsL_reg[2][2]/P0001  & n1290 ;
  assign n1278 = ~\i_tv80_core_RegAddrC_reg[1]/NET0131  & ~\i_tv80_core_RegAddrC_reg[2]/NET0131  ;
  assign n1292 = \i_tv80_core_RegAddrC_reg[0]/P0001  & n1278 ;
  assign n1293 = \i_tv80_core_i_reg_RegsL_reg[1][2]/P0001  & n1292 ;
  assign n1300 = ~n1291 & ~n1293 ;
  assign n1284 = \i_tv80_core_RegAddrC_reg[1]/NET0131  & \i_tv80_core_RegAddrC_reg[2]/NET0131  ;
  assign n1294 = \i_tv80_core_RegAddrC_reg[0]/P0001  & n1284 ;
  assign n1295 = \i_tv80_core_i_reg_RegsL_reg[7][2]/P0001  & n1294 ;
  assign n1296 = \i_tv80_core_RegAddrC_reg[0]/P0001  & n1289 ;
  assign n1297 = \i_tv80_core_i_reg_RegsL_reg[3][2]/P0001  & n1296 ;
  assign n1301 = ~n1295 & ~n1297 ;
  assign n1302 = n1300 & n1301 ;
  assign n1279 = ~\i_tv80_core_RegAddrC_reg[0]/P0001  & n1278 ;
  assign n1280 = \i_tv80_core_i_reg_RegsL_reg[0][2]/P0001  & n1279 ;
  assign n1281 = ~\i_tv80_core_RegAddrC_reg[1]/NET0131  & \i_tv80_core_RegAddrC_reg[2]/NET0131  ;
  assign n1282 = ~\i_tv80_core_RegAddrC_reg[0]/P0001  & n1281 ;
  assign n1283 = \i_tv80_core_i_reg_RegsL_reg[4][2]/P0001  & n1282 ;
  assign n1298 = ~n1280 & ~n1283 ;
  assign n1285 = ~\i_tv80_core_RegAddrC_reg[0]/P0001  & n1284 ;
  assign n1286 = \i_tv80_core_i_reg_RegsL_reg[6][2]/P0001  & n1285 ;
  assign n1287 = \i_tv80_core_RegAddrC_reg[0]/P0001  & n1281 ;
  assign n1288 = \i_tv80_core_i_reg_RegsL_reg[5][2]/P0001  & n1287 ;
  assign n1299 = ~n1286 & ~n1288 ;
  assign n1303 = n1298 & n1299 ;
  assign n1304 = n1302 & n1303 ;
  assign n1305 = n1277 & ~n1304 ;
  assign n1306 = ~\i_tv80_core_ISet_reg[0]/NET0131  & n956 ;
  assign n1307 = ~\i_tv80_core_ISet_reg[1]/P0001  & n1306 ;
  assign n1308 = n939 & n1307 ;
  assign n1311 = ~n871 & ~n974 ;
  assign n1309 = ~\i_tv80_core_mcycle_reg[1]/P0001  & \i_tv80_core_mcycle_reg[2]/P0001  ;
  assign n1310 = \i_tv80_core_mcycle_reg[0]/P0001  & n1309 ;
  assign n1312 = n382 & n1310 ;
  assign n1313 = ~n1311 & n1312 ;
  assign n1314 = ~n1308 & ~n1313 ;
  assign n1315 = ~\i_tv80_core_IStatus_reg[0]/P0001  & \i_tv80_core_IStatus_reg[1]/P0001  ;
  assign n1316 = \i_tv80_core_IntCycle_reg/P0001  & n1315 ;
  assign n1317 = n956 & n1316 ;
  assign n1318 = n1314 & ~n1317 ;
  assign n1319 = \i_tv80_core_TmpAddr_reg[2]/P0001  & ~n1318 ;
  assign n1320 = ~\i_tv80_core_mcycle_reg[2]/P0001  & \i_tv80_core_mcycles_reg[2]/P0001  ;
  assign n1321 = \i_tv80_core_mcycle_reg[0]/P0001  & ~\i_tv80_core_mcycles_reg[0]/P0001  ;
  assign n1326 = ~n1320 & ~n1321 ;
  assign n1322 = \i_tv80_core_mcycle_reg[1]/P0001  & ~\i_tv80_core_mcycles_reg[1]/P0001  ;
  assign n1323 = ~\i_tv80_core_mcycle_reg[1]/P0001  & \i_tv80_core_mcycles_reg[1]/P0001  ;
  assign n1327 = ~n1322 & ~n1323 ;
  assign n1324 = ~\i_tv80_core_mcycle_reg[0]/P0001  & \i_tv80_core_mcycles_reg[0]/P0001  ;
  assign n1325 = \i_tv80_core_mcycle_reg[2]/P0001  & ~\i_tv80_core_mcycles_reg[2]/P0001  ;
  assign n1328 = ~n1324 & ~n1325 ;
  assign n1329 = n1327 & n1328 ;
  assign n1330 = n1326 & n1329 ;
  assign n1331 = \i_tv80_core_NMICycle_reg/P0001  & n1330 ;
  assign n1332 = n1314 & n1331 ;
  assign n1333 = ~n1319 & ~n1332 ;
  assign n1334 = n686 & n1066 ;
  assign n1335 = n889 & n919 ;
  assign n1336 = ~n1334 & ~n1335 ;
  assign n1337 = n862 & ~n1336 ;
  assign n1364 = \i_tv80_core_IR_reg[6]/P0001  & n1069 ;
  assign n1365 = ~n860 & n1364 ;
  assign n1394 = n1311 & ~n1365 ;
  assign n1366 = n875 & n883 ;
  assign n1367 = \i_tv80_core_IR_reg[3]/P0001  & n936 ;
  assign n1368 = \i_tv80_core_IR_reg[5]/P0001  & n941 ;
  assign n1369 = n1367 & n1368 ;
  assign n1370 = ~n1366 & ~n1369 ;
  assign n1371 = n376 & n1075 ;
  assign n1372 = \i_tv80_core_IR_reg[6]/P0001  & n976 ;
  assign n1373 = ~n1371 & ~n1372 ;
  assign n1395 = n1370 & n1373 ;
  assign n1396 = n1394 & n1395 ;
  assign n1362 = ~n857 & n1335 ;
  assign n1361 = ~\i_tv80_core_IR_reg[6]/P0001  & n1069 ;
  assign n1392 = n945 & ~n1065 ;
  assign n1393 = ~n1361 & n1392 ;
  assign n1397 = ~n1362 & n1393 ;
  assign n1398 = n1396 & n1397 ;
  assign n1363 = ~n381 & n921 ;
  assign n1384 = n875 & n1086 ;
  assign n1377 = n928 & n1075 ;
  assign n1378 = n878 & n881 ;
  assign n1385 = ~n1377 & ~n1378 ;
  assign n1386 = ~n1384 & n1385 ;
  assign n1379 = \i_tv80_core_IR_reg[0]/P0001  & n1028 ;
  assign n1380 = n918 & n1379 ;
  assign n1381 = n681 & n901 ;
  assign n1382 = n904 & n1381 ;
  assign n1383 = \i_tv80_core_IR_reg[0]/P0001  & n1382 ;
  assign n1387 = ~n1380 & ~n1383 ;
  assign n1388 = n1386 & n1387 ;
  assign n1375 = n1086 & n1367 ;
  assign n1376 = ~n1276 & ~n1375 ;
  assign n1374 = n376 & n893 ;
  assign n1389 = ~n1171 & ~n1374 ;
  assign n1390 = n1376 & n1389 ;
  assign n1391 = n1388 & n1390 ;
  assign n1399 = ~n1363 & n1391 ;
  assign n1400 = n1398 & n1399 ;
  assign n1407 = n376 & n897 ;
  assign n1408 = ~n377 & ~n1407 ;
  assign n1409 = ~n905 & n1408 ;
  assign n1401 = n890 & n1075 ;
  assign n1402 = n373 & n890 ;
  assign n1403 = n373 & n896 ;
  assign n1404 = ~n1402 & ~n1403 ;
  assign n1405 = ~n1401 & n1404 ;
  assign n1406 = ~n860 & ~n1405 ;
  assign n1410 = \i_tv80_core_IR_reg[5]/P0001  & n1039 ;
  assign n1411 = ~n1067 & ~n1410 ;
  assign n1412 = ~n886 & n951 ;
  assign n1413 = n1411 & ~n1412 ;
  assign n1414 = ~n1406 & n1413 ;
  assign n1415 = n1409 & n1414 ;
  assign n1338 = n897 & n928 ;
  assign n1339 = n893 & n928 ;
  assign n1340 = ~n1087 & ~n1339 ;
  assign n1341 = ~n1338 & n1340 ;
  assign n1342 = ~n925 & n1341 ;
  assign n1343 = n1082 & n1342 ;
  assign n1416 = ~n884 & ~n898 ;
  assign n1350 = n878 & n1070 ;
  assign n1351 = ~n939 & ~n1350 ;
  assign n1352 = ~n910 & n1351 ;
  assign n1353 = \i_tv80_core_IR_reg[7]/P0001  & n886 ;
  assign n1354 = ~\i_tv80_core_IR_reg[6]/P0001  & n1353 ;
  assign n1355 = ~n860 & n1354 ;
  assign n1422 = n1352 & ~n1355 ;
  assign n1423 = n1416 & n1422 ;
  assign n1417 = ~n879 & ~n887 ;
  assign n1418 = ~n915 & n1417 ;
  assign n1356 = n889 & n943 ;
  assign n1357 = n868 & n913 ;
  assign n1358 = ~n673 & n1357 ;
  assign n1359 = ~n1356 & ~n1358 ;
  assign n1360 = n890 & n897 ;
  assign n1419 = n1359 & ~n1360 ;
  assign n1420 = n1418 & n1419 ;
  assign n1344 = n854 & n947 ;
  assign n1345 = ~n929 & ~n948 ;
  assign n1346 = ~n1344 & n1345 ;
  assign n1347 = ~\i_tv80_core_IR_reg[3]/P0001  & n1013 ;
  assign n1348 = n1114 & n1347 ;
  assign n1349 = ~n894 & ~n1348 ;
  assign n1421 = n1346 & n1349 ;
  assign n1424 = n1420 & n1421 ;
  assign n1425 = n1423 & n1424 ;
  assign n1426 = n1343 & n1425 ;
  assign n1427 = n1415 & n1426 ;
  assign n1428 = n1400 & n1427 ;
  assign n1429 = n382 & ~n1428 ;
  assign n1430 = \i_tv80_core_ISet_reg[0]/NET0131  & ~\i_tv80_core_ISet_reg[1]/P0001  ;
  assign n1431 = n856 & ~n989 ;
  assign n1432 = ~\i_tv80_core_mcycle_reg[0]/P0001  & ~n1431 ;
  assign n1433 = n886 & ~n1309 ;
  assign n1434 = ~n956 & n1433 ;
  assign n1435 = ~n1432 & n1434 ;
  assign n1436 = n1430 & ~n1435 ;
  assign n1440 = \i_tv80_core_IR_reg[0]/P0001  & n1012 ;
  assign n1441 = ~n1036 & ~n1440 ;
  assign n1442 = ~n860 & ~n1441 ;
  assign n1437 = ~n381 & n1007 ;
  assign n1439 = ~n1033 & ~n1050 ;
  assign n1438 = ~n856 & n1034 ;
  assign n1443 = n996 & ~n1438 ;
  assign n1444 = n1439 & n1443 ;
  assign n1445 = ~n1437 & n1444 ;
  assign n1446 = ~n1442 & n1445 ;
  assign n1447 = ~n1037 & ~n1039 ;
  assign n1448 = ~n1010 & n1447 ;
  assign n1449 = n1003 & n1019 ;
  assign n1450 = n1448 & n1449 ;
  assign n1451 = n1013 & n1049 ;
  assign n1452 = ~n1042 & ~n1451 ;
  assign n1453 = n924 & n1005 ;
  assign n1454 = n1452 & ~n1453 ;
  assign n1455 = n1450 & n1454 ;
  assign n1456 = n1446 & n1455 ;
  assign n1457 = \i_tv80_core_ISet_reg[1]/P0001  & ~n1456 ;
  assign n1458 = ~n1436 & ~n1457 ;
  assign n1459 = ~n1429 & n1458 ;
  assign n1460 = ~n862 & ~n1459 ;
  assign n1461 = ~n1337 & ~n1460 ;
  assign n1462 = \i_tv80_core_mcycle_reg[2]/P0001  & n378 ;
  assign n1463 = ~n1430 & n1462 ;
  assign n1582 = ~n1461 & ~n1463 ;
  assign n1469 = ~n381 & n1014 ;
  assign n1471 = \i_tv80_core_ISet_reg[1]/P0001  & n1018 ;
  assign n1472 = n1452 & n1471 ;
  assign n1473 = ~n1469 & n1472 ;
  assign n1476 = n1004 & n1473 ;
  assign n1468 = ~n1034 & ~n1440 ;
  assign n1470 = ~n857 & n1007 ;
  assign n1477 = n1468 & ~n1470 ;
  assign n1478 = n1476 & n1477 ;
  assign n1464 = ~n1020 & ~n1036 ;
  assign n1465 = ~n860 & ~n1464 ;
  assign n1466 = n374 & n1005 ;
  assign n1467 = ~n857 & n1466 ;
  assign n1474 = n1439 & n1448 ;
  assign n1475 = ~n1467 & n1474 ;
  assign n1479 = ~n1465 & n1475 ;
  assign n1480 = n1478 & n1479 ;
  assign n1505 = ~n1338 & ~n1354 ;
  assign n1491 = ~n857 & n1350 ;
  assign n1492 = n929 & n930 ;
  assign n1506 = ~n1491 & ~n1492 ;
  assign n1507 = n1505 & n1506 ;
  assign n1516 = n900 & n1507 ;
  assign n1498 = ~n857 & n879 ;
  assign n1499 = ~n1348 & n1359 ;
  assign n1500 = ~n1498 & n1499 ;
  assign n1501 = ~n381 & ~n1346 ;
  assign n1517 = n1500 & ~n1501 ;
  assign n1518 = n1516 & n1517 ;
  assign n1510 = n1340 & n1370 ;
  assign n1481 = ~\i_tv80_core_mcycle_reg[0]/P0001  & n1309 ;
  assign n1482 = ~n956 & ~n1481 ;
  assign n1483 = n871 & n1482 ;
  assign n1484 = ~n1071 & ~n1360 ;
  assign n1511 = ~n1483 & n1484 ;
  assign n1514 = n1510 & n1511 ;
  assign n1502 = n382 & ~n1069 ;
  assign n1503 = ~n1371 & n1502 ;
  assign n1504 = ~n910 & ~n1065 ;
  assign n1508 = n1503 & n1504 ;
  assign n1509 = n1079 & ~n1080 ;
  assign n1515 = n1508 & n1509 ;
  assign n1519 = n1514 & n1515 ;
  assign n1522 = n1518 & n1519 ;
  assign n1523 = n1415 & n1522 ;
  assign n1496 = ~n971 & ~n1482 ;
  assign n1497 = n974 & ~n1496 ;
  assign n1493 = n860 & n970 ;
  assign n1494 = n381 & ~n1493 ;
  assign n1495 = n944 & ~n1494 ;
  assign n1490 = ~\i_tv80_core_IR_reg[0]/P0001  & n919 ;
  assign n1485 = ~n939 & ~n942 ;
  assign n1486 = ~n381 & ~n1485 ;
  assign n1487 = \i_tv80_core_mcycle_reg[2]/P0001  & n379 ;
  assign n1488 = ~n1083 & ~n1487 ;
  assign n1489 = n977 & n1488 ;
  assign n1512 = ~n1486 & ~n1489 ;
  assign n1513 = ~n1490 & n1512 ;
  assign n1520 = n922 & n1513 ;
  assign n1521 = n1391 & n1520 ;
  assign n1524 = ~n1495 & n1521 ;
  assign n1525 = ~n1497 & n1524 ;
  assign n1526 = n1523 & n1525 ;
  assign n1527 = ~n1480 & ~n1526 ;
  assign n1528 = ~n862 & ~n1527 ;
  assign n1529 = ~n1463 & n1528 ;
  assign n1539 = ~n860 & n1403 ;
  assign n1538 = ~n929 & ~n1412 ;
  assign n1544 = ~n1491 & n1538 ;
  assign n1545 = ~n1539 & n1544 ;
  assign n1549 = n1409 & n1545 ;
  assign n1532 = ~n1344 & n1411 ;
  assign n1550 = n1500 & n1532 ;
  assign n1551 = n1549 & n1550 ;
  assign n1533 = n890 & n892 ;
  assign n1534 = n898 & ~n1487 ;
  assign n1535 = ~n1533 & ~n1534 ;
  assign n1536 = ~n956 & ~n1535 ;
  assign n1541 = ~n948 & ~n1401 ;
  assign n1542 = ~n1402 & n1541 ;
  assign n1540 = ~n915 & ~n939 ;
  assign n1543 = n888 & n1540 ;
  assign n1546 = n1542 & n1543 ;
  assign n1537 = n910 & n1482 ;
  assign n1547 = ~n1355 & ~n1537 ;
  assign n1548 = n1546 & n1547 ;
  assign n1552 = ~n1536 & n1548 ;
  assign n1553 = n1551 & n1552 ;
  assign n1554 = n1343 & n1553 ;
  assign n1555 = n1400 & n1554 ;
  assign n1556 = n382 & ~n1555 ;
  assign n1559 = n924 & n1006 ;
  assign n1558 = ~n860 & n1466 ;
  assign n1557 = n1451 & n1482 ;
  assign n1560 = ~n1042 & ~n1557 ;
  assign n1561 = ~n1558 & n1560 ;
  assign n1562 = ~n1559 & n1561 ;
  assign n1563 = n1450 & n1562 ;
  assign n1564 = n1446 & n1563 ;
  assign n1565 = \i_tv80_core_ISet_reg[1]/P0001  & ~n1564 ;
  assign n1566 = ~n1436 & ~n1565 ;
  assign n1567 = ~n1556 & n1566 ;
  assign n1568 = ~n862 & ~n1567 ;
  assign n1569 = ~n1337 & ~n1568 ;
  assign n1570 = ~n1463 & ~n1569 ;
  assign n1583 = ~n1529 & ~n1570 ;
  assign n1595 = ~n1582 & n1583 ;
  assign n1596 = n860 & ~n1336 ;
  assign n1597 = ~n1595 & ~n1596 ;
  assign n1593 = ~\i_tv80_core_XY_State_reg[0]/NET0131  & ~\i_tv80_core_XY_State_reg[1]/P0001  ;
  assign n1598 = ~\i_tv80_core_XY_Ind_reg/P0001  & ~n1593 ;
  assign n1599 = ~n1597 & n1598 ;
  assign n1601 = \i_tv80_core_PC_reg[2]/P0001  & n1599 ;
  assign n1600 = \i_tv80_core_TmpAddr_reg[2]/P0001  & ~n1599 ;
  assign n1602 = ~n1593 & ~n1600 ;
  assign n1603 = ~n1601 & n1602 ;
  assign n1594 = n1304 & n1593 ;
  assign n1604 = ~n1594 & n1595 ;
  assign n1605 = ~n1603 & n1604 ;
  assign n1584 = n1582 & n1583 ;
  assign n1573 = n892 & n896 ;
  assign n1574 = n382 & n1573 ;
  assign n1575 = \i_tv80_core_ISet_reg[1]/P0001  & n993 ;
  assign n1576 = n1063 & n1575 ;
  assign n1577 = ~n1574 & ~n1576 ;
  assign n1578 = n1481 & ~n1577 ;
  assign n1579 = \i_tv80_core_TmpAddr_reg[0]/P0001  & n1578 ;
  assign n1580 = \i_tv80_core_TmpAddr_reg[1]/P0001  & n1579 ;
  assign n1581 = ~\i_tv80_core_TmpAddr_reg[2]/P0001  & ~n1580 ;
  assign n1585 = \i_tv80_core_TmpAddr_reg[2]/P0001  & n1580 ;
  assign n1586 = ~n1581 & ~n1585 ;
  assign n1587 = n1584 & n1586 ;
  assign n1530 = n1461 & n1529 ;
  assign n1531 = ~n1304 & n1530 ;
  assign n1571 = n1527 & n1570 ;
  assign n1572 = \i_tv80_core_PC_reg[2]/P0001  & n1571 ;
  assign n1606 = ~n1531 & ~n1572 ;
  assign n1607 = ~n1587 & n1606 ;
  assign n1588 = n1528 & n1582 ;
  assign n1589 = n1569 & n1588 ;
  assign n1590 = \di_reg_reg[2]/P0001  & n1589 ;
  assign n1591 = ~n1569 & n1588 ;
  assign n1592 = \i_tv80_core_SP_reg[2]/P0001  & n1591 ;
  assign n1608 = ~n1590 & ~n1592 ;
  assign n1609 = n1607 & n1608 ;
  assign n1610 = ~n1605 & n1609 ;
  assign n1611 = n1318 & ~n1610 ;
  assign n1612 = n1333 & ~n1611 ;
  assign n1613 = ~n1277 & ~n1612 ;
  assign n1614 = ~n1305 & ~n1613 ;
  assign n1615 = n1014 & n1128 ;
  assign n1616 = \i_tv80_core_IntCycle_reg/P0001  & ~\i_tv80_core_NMICycle_reg/P0001  ;
  assign n1617 = n929 & n1616 ;
  assign n1618 = n1310 & n1617 ;
  assign n1619 = ~n970 & n1356 ;
  assign n1620 = n945 & ~n1071 ;
  assign n1621 = ~n1619 & n1620 ;
  assign n1622 = n956 & ~n1621 ;
  assign n1623 = ~n1618 & ~n1622 ;
  assign n1624 = n382 & ~n1623 ;
  assign n1625 = ~n1615 & ~n1624 ;
  assign n1626 = ~n1614 & n1625 ;
  assign n1627 = \i_tv80_core_TmpAddr_reg[2]/P0001  & ~n1625 ;
  assign n1628 = n1103 & ~n1627 ;
  assign n1629 = ~n1626 & n1628 ;
  assign n1630 = ~\A[2]_pad  & ~n1103 ;
  assign n1631 = ~n1113 & ~n1630 ;
  assign n1632 = ~n1629 & n1631 ;
  assign n1633 = ~\i_tv80_core_tstate_reg[0]/P0001  & \i_tv80_core_tstate_reg[1]/NET0131  ;
  assign n1634 = ~\i_tv80_core_tstate_reg[2]/NET0131  & n1633 ;
  assign n1635 = wait_n_pad & n1634 ;
  assign n1637 = ~\i_tv80_core_R_reg[2]/P0001  & n1635 ;
  assign n1636 = ~\A[2]_pad  & ~n1635 ;
  assign n1638 = n1113 & ~n1636 ;
  assign n1639 = ~n1637 & n1638 ;
  assign n1640 = ~\i_tv80_core_BusAck_reg/P0001  & ~n1639 ;
  assign n1641 = ~n1632 & n1640 ;
  assign n1642 = ~\A[2]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n1643 = reset_n_pad & ~n1642 ;
  assign n1644 = ~n1641 & n1643 ;
  assign n1649 = \i_tv80_core_i_reg_RegsL_reg[2][1]/P0001  & n1290 ;
  assign n1650 = \i_tv80_core_i_reg_RegsL_reg[1][1]/P0001  & n1292 ;
  assign n1655 = ~n1649 & ~n1650 ;
  assign n1651 = \i_tv80_core_i_reg_RegsL_reg[7][1]/P0001  & n1294 ;
  assign n1652 = \i_tv80_core_i_reg_RegsL_reg[3][1]/P0001  & n1296 ;
  assign n1656 = ~n1651 & ~n1652 ;
  assign n1657 = n1655 & n1656 ;
  assign n1645 = \i_tv80_core_i_reg_RegsL_reg[0][1]/P0001  & n1279 ;
  assign n1646 = \i_tv80_core_i_reg_RegsL_reg[4][1]/P0001  & n1282 ;
  assign n1653 = ~n1645 & ~n1646 ;
  assign n1647 = \i_tv80_core_i_reg_RegsL_reg[6][1]/P0001  & n1285 ;
  assign n1648 = \i_tv80_core_i_reg_RegsL_reg[5][1]/P0001  & n1287 ;
  assign n1654 = ~n1647 & ~n1648 ;
  assign n1658 = n1653 & n1654 ;
  assign n1659 = n1657 & n1658 ;
  assign n1660 = n1277 & ~n1659 ;
  assign n1661 = \i_tv80_core_TmpAddr_reg[1]/P0001  & ~n1318 ;
  assign n1662 = ~n1332 & ~n1661 ;
  assign n1672 = \i_tv80_core_PC_reg[1]/P0001  & n1599 ;
  assign n1671 = \i_tv80_core_TmpAddr_reg[1]/P0001  & ~n1599 ;
  assign n1673 = ~n1593 & ~n1671 ;
  assign n1674 = ~n1672 & n1673 ;
  assign n1670 = n1593 & n1659 ;
  assign n1675 = n1595 & ~n1670 ;
  assign n1676 = ~n1674 & n1675 ;
  assign n1665 = ~\i_tv80_core_TmpAddr_reg[1]/P0001  & ~n1579 ;
  assign n1666 = ~n1580 & ~n1665 ;
  assign n1667 = n1584 & n1666 ;
  assign n1663 = n1530 & ~n1659 ;
  assign n1664 = \i_tv80_core_PC_reg[1]/P0001  & n1571 ;
  assign n1677 = ~n1663 & ~n1664 ;
  assign n1678 = ~n1667 & n1677 ;
  assign n1668 = \di_reg_reg[1]/P0001  & n1589 ;
  assign n1669 = \i_tv80_core_SP_reg[1]/P0001  & n1591 ;
  assign n1679 = ~n1668 & ~n1669 ;
  assign n1680 = n1678 & n1679 ;
  assign n1681 = ~n1676 & n1680 ;
  assign n1682 = n1318 & ~n1681 ;
  assign n1683 = n1662 & ~n1682 ;
  assign n1684 = ~n1277 & ~n1683 ;
  assign n1685 = ~n1660 & ~n1684 ;
  assign n1686 = n1625 & ~n1685 ;
  assign n1687 = \i_tv80_core_TmpAddr_reg[1]/P0001  & ~n1625 ;
  assign n1688 = n1103 & ~n1687 ;
  assign n1689 = ~n1686 & n1688 ;
  assign n1690 = ~\A[1]_pad  & ~n1103 ;
  assign n1691 = ~n1113 & ~n1690 ;
  assign n1692 = ~n1689 & n1691 ;
  assign n1694 = ~\i_tv80_core_R_reg[1]/P0001  & n1635 ;
  assign n1693 = ~\A[1]_pad  & ~n1635 ;
  assign n1695 = n1113 & ~n1693 ;
  assign n1696 = ~n1694 & n1695 ;
  assign n1697 = ~\i_tv80_core_BusAck_reg/P0001  & ~n1696 ;
  assign n1698 = ~n1692 & n1697 ;
  assign n1699 = ~\A[1]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n1700 = reset_n_pad & ~n1699 ;
  assign n1701 = ~n1698 & n1700 ;
  assign n1706 = \i_tv80_core_i_reg_RegsL_reg[2][5]/NET0131  & n1290 ;
  assign n1707 = \i_tv80_core_i_reg_RegsL_reg[1][5]/NET0131  & n1292 ;
  assign n1712 = ~n1706 & ~n1707 ;
  assign n1708 = \i_tv80_core_i_reg_RegsL_reg[7][5]/NET0131  & n1294 ;
  assign n1709 = \i_tv80_core_i_reg_RegsL_reg[3][5]/NET0131  & n1296 ;
  assign n1713 = ~n1708 & ~n1709 ;
  assign n1714 = n1712 & n1713 ;
  assign n1702 = \i_tv80_core_i_reg_RegsL_reg[0][5]/NET0131  & n1279 ;
  assign n1703 = \i_tv80_core_i_reg_RegsL_reg[4][5]/NET0131  & n1282 ;
  assign n1710 = ~n1702 & ~n1703 ;
  assign n1704 = \i_tv80_core_i_reg_RegsL_reg[6][5]/NET0131  & n1285 ;
  assign n1705 = \i_tv80_core_i_reg_RegsL_reg[5][5]/NET0131  & n1287 ;
  assign n1711 = ~n1704 & ~n1705 ;
  assign n1715 = n1710 & n1711 ;
  assign n1716 = n1714 & n1715 ;
  assign n1717 = n1277 & ~n1716 ;
  assign n1718 = \i_tv80_core_TmpAddr_reg[5]/P0001  & ~n1318 ;
  assign n1719 = ~n1332 & ~n1718 ;
  assign n1733 = \i_tv80_core_PC_reg[5]/P0001  & n1599 ;
  assign n1732 = \i_tv80_core_TmpAddr_reg[5]/P0001  & ~n1599 ;
  assign n1734 = ~n1593 & ~n1732 ;
  assign n1735 = ~n1733 & n1734 ;
  assign n1731 = n1593 & n1716 ;
  assign n1736 = n1595 & ~n1731 ;
  assign n1737 = ~n1735 & n1736 ;
  assign n1722 = \i_tv80_core_TmpAddr_reg[2]/P0001  & \i_tv80_core_TmpAddr_reg[3]/P0001  ;
  assign n1723 = n1580 & n1722 ;
  assign n1724 = \i_tv80_core_TmpAddr_reg[4]/P0001  & n1723 ;
  assign n1725 = \i_tv80_core_TmpAddr_reg[5]/P0001  & n1724 ;
  assign n1726 = ~\i_tv80_core_TmpAddr_reg[5]/P0001  & ~n1724 ;
  assign n1727 = ~n1725 & ~n1726 ;
  assign n1728 = n1584 & n1727 ;
  assign n1720 = n1530 & ~n1716 ;
  assign n1721 = \i_tv80_core_PC_reg[5]/P0001  & n1571 ;
  assign n1738 = ~n1720 & ~n1721 ;
  assign n1739 = ~n1728 & n1738 ;
  assign n1729 = \di_reg_reg[5]/P0001  & n1589 ;
  assign n1730 = \i_tv80_core_SP_reg[5]/P0001  & n1591 ;
  assign n1740 = ~n1729 & ~n1730 ;
  assign n1741 = n1739 & n1740 ;
  assign n1742 = ~n1737 & n1741 ;
  assign n1743 = n1318 & ~n1742 ;
  assign n1744 = n1719 & ~n1743 ;
  assign n1745 = ~n1277 & ~n1744 ;
  assign n1746 = ~n1717 & ~n1745 ;
  assign n1747 = n1625 & ~n1746 ;
  assign n1748 = \i_tv80_core_TmpAddr_reg[5]/P0001  & ~n1625 ;
  assign n1749 = n1103 & ~n1748 ;
  assign n1750 = ~n1747 & n1749 ;
  assign n1751 = ~\A[5]_pad  & ~n1103 ;
  assign n1752 = ~n1113 & ~n1751 ;
  assign n1753 = ~n1750 & n1752 ;
  assign n1755 = ~\i_tv80_core_R_reg[5]/P0001  & n1635 ;
  assign n1754 = ~\A[5]_pad  & ~n1635 ;
  assign n1756 = n1113 & ~n1754 ;
  assign n1757 = ~n1755 & n1756 ;
  assign n1758 = ~\i_tv80_core_BusAck_reg/P0001  & ~n1757 ;
  assign n1759 = ~n1753 & n1758 ;
  assign n1760 = ~\A[5]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n1761 = reset_n_pad & ~n1760 ;
  assign n1762 = ~n1759 & n1761 ;
  assign n1767 = \i_tv80_core_i_reg_RegsL_reg[2][6]/NET0131  & n1290 ;
  assign n1768 = \i_tv80_core_i_reg_RegsL_reg[1][6]/NET0131  & n1292 ;
  assign n1773 = ~n1767 & ~n1768 ;
  assign n1769 = \i_tv80_core_i_reg_RegsL_reg[7][6]/NET0131  & n1294 ;
  assign n1770 = \i_tv80_core_i_reg_RegsL_reg[5][6]/NET0131  & n1287 ;
  assign n1774 = ~n1769 & ~n1770 ;
  assign n1775 = n1773 & n1774 ;
  assign n1763 = \i_tv80_core_i_reg_RegsL_reg[0][6]/NET0131  & n1279 ;
  assign n1764 = \i_tv80_core_i_reg_RegsL_reg[6][6]/NET0131  & n1285 ;
  assign n1771 = ~n1763 & ~n1764 ;
  assign n1765 = \i_tv80_core_i_reg_RegsL_reg[4][6]/NET0131  & n1282 ;
  assign n1766 = \i_tv80_core_i_reg_RegsL_reg[3][6]/NET0131  & n1296 ;
  assign n1772 = ~n1765 & ~n1766 ;
  assign n1776 = n1771 & n1772 ;
  assign n1777 = n1775 & n1776 ;
  assign n1778 = n1277 & ~n1777 ;
  assign n1779 = \i_tv80_core_TmpAddr_reg[6]/P0001  & ~n1318 ;
  assign n1780 = ~n1332 & ~n1779 ;
  assign n1791 = \i_tv80_core_PC_reg[6]/P0001  & n1599 ;
  assign n1790 = \i_tv80_core_TmpAddr_reg[6]/P0001  & ~n1599 ;
  assign n1792 = ~n1593 & ~n1790 ;
  assign n1793 = ~n1791 & n1792 ;
  assign n1789 = n1593 & n1777 ;
  assign n1794 = n1595 & ~n1789 ;
  assign n1795 = ~n1793 & n1794 ;
  assign n1783 = ~\i_tv80_core_TmpAddr_reg[6]/P0001  & ~n1725 ;
  assign n1784 = \i_tv80_core_TmpAddr_reg[6]/P0001  & n1725 ;
  assign n1785 = ~n1783 & ~n1784 ;
  assign n1786 = n1584 & n1785 ;
  assign n1781 = n1530 & ~n1777 ;
  assign n1782 = \i_tv80_core_PC_reg[6]/P0001  & n1571 ;
  assign n1796 = ~n1781 & ~n1782 ;
  assign n1797 = ~n1786 & n1796 ;
  assign n1787 = \i_tv80_core_SP_reg[6]/P0001  & n1591 ;
  assign n1788 = \di_reg_reg[6]/P0001  & n1589 ;
  assign n1798 = ~n1787 & ~n1788 ;
  assign n1799 = n1797 & n1798 ;
  assign n1800 = ~n1795 & n1799 ;
  assign n1801 = n1318 & ~n1800 ;
  assign n1802 = n1780 & ~n1801 ;
  assign n1803 = ~n1277 & ~n1802 ;
  assign n1804 = ~n1778 & ~n1803 ;
  assign n1805 = n1625 & ~n1804 ;
  assign n1806 = \i_tv80_core_TmpAddr_reg[6]/P0001  & ~n1625 ;
  assign n1807 = n1103 & ~n1806 ;
  assign n1808 = ~n1805 & n1807 ;
  assign n1809 = ~\A[6]_pad  & ~n1103 ;
  assign n1810 = ~n1113 & ~n1809 ;
  assign n1811 = ~n1808 & n1810 ;
  assign n1813 = ~\i_tv80_core_R_reg[6]/P0001  & n1635 ;
  assign n1812 = ~\A[6]_pad  & ~n1635 ;
  assign n1814 = n1113 & ~n1812 ;
  assign n1815 = ~n1813 & n1814 ;
  assign n1816 = ~\i_tv80_core_BusAck_reg/P0001  & ~n1815 ;
  assign n1817 = ~n1811 & n1816 ;
  assign n1818 = ~\A[6]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n1819 = reset_n_pad & ~n1818 ;
  assign n1820 = ~n1817 & n1819 ;
  assign n1832 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n555 ;
  assign n1826 = n735 & ~n770 ;
  assign n1831 = n604 & ~n632 ;
  assign n1828 = \i_tv80_core_ALU_Op_r_reg[0]/P0001  & n676 ;
  assign n1827 = ~\i_tv80_core_BusB_reg[7]/P0001  & ~n676 ;
  assign n1829 = n1175 & ~n1827 ;
  assign n1830 = ~n1828 & n1829 ;
  assign n1823 = \i_tv80_core_BusA_reg[7]/P0001  & n700 ;
  assign n1824 = n370 & n677 ;
  assign n1825 = ~n1823 & ~n1824 ;
  assign n1833 = \i_tv80_core_Save_ALU_r_reg/P0001  & n1825 ;
  assign n1834 = ~n1830 & n1833 ;
  assign n1835 = ~n1831 & n1834 ;
  assign n1836 = ~n1826 & n1835 ;
  assign n1837 = ~n1832 & n1836 ;
  assign n1822 = ~\di_reg_reg[7]/P0001  & ~\i_tv80_core_Save_ALU_r_reg/P0001  ;
  assign n1838 = ~n1172 & ~n1822 ;
  assign n1839 = ~n1837 & n1838 ;
  assign n1840 = \i_tv80_core_BusB_reg[7]/P0001  & n1172 ;
  assign n1841 = ~n1839 & ~n1840 ;
  assign n1842 = n1167 & ~n1841 ;
  assign n1844 = \i_tv80_core_Fp_reg[7]/P0001  & n1118 ;
  assign n1845 = \i_tv80_core_F_reg[7]/P0001  & ~n1118 ;
  assign n1846 = ~n1844 & ~n1845 ;
  assign n1847 = n386 & n1846 ;
  assign n1848 = ~\i_tv80_core_Arith16_r_reg/P0001  & n555 ;
  assign n1849 = \i_tv80_core_Arith16_r_reg/P0001  & ~\i_tv80_core_F_reg[7]/P0001  ;
  assign n1850 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n1849 ;
  assign n1851 = ~n1848 & n1850 ;
  assign n1853 = ~\i_tv80_core_F_reg[7]/P0001  & n382 ;
  assign n1854 = n604 & ~n1853 ;
  assign n1855 = ~n1235 & n1854 ;
  assign n1852 = \i_tv80_core_F_reg[7]/P0001  & n697 ;
  assign n1856 = n1825 & ~n1852 ;
  assign n1857 = ~n386 & n1856 ;
  assign n1858 = ~n1855 & n1857 ;
  assign n1859 = ~n1826 & n1858 ;
  assign n1860 = ~n1851 & n1859 ;
  assign n1861 = ~n1847 & ~n1860 ;
  assign n1862 = ~n1105 & ~n1861 ;
  assign n1843 = ~\di_reg_reg[7]/P0001  & n1105 ;
  assign n1863 = ~n1167 & ~n1843 ;
  assign n1864 = ~n1862 & n1863 ;
  assign n1865 = ~n1842 & ~n1864 ;
  assign n1866 = ~\i_tv80_core_BusAck_reg/P0001  & ~n1865 ;
  assign n1821 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_F_reg[7]/P0001  ;
  assign n1867 = reset_n_pad & ~n1821 ;
  assign n1868 = ~n1866 & n1867 ;
  assign n1873 = \i_tv80_core_i_reg_RegsL_reg[2][0]/P0001  & n1290 ;
  assign n1874 = \i_tv80_core_i_reg_RegsL_reg[1][0]/P0001  & n1292 ;
  assign n1879 = ~n1873 & ~n1874 ;
  assign n1875 = \i_tv80_core_i_reg_RegsL_reg[7][0]/P0001  & n1294 ;
  assign n1876 = \i_tv80_core_i_reg_RegsL_reg[3][0]/P0001  & n1296 ;
  assign n1880 = ~n1875 & ~n1876 ;
  assign n1881 = n1879 & n1880 ;
  assign n1869 = \i_tv80_core_i_reg_RegsL_reg[0][0]/P0001  & n1279 ;
  assign n1870 = \i_tv80_core_i_reg_RegsL_reg[4][0]/P0001  & n1282 ;
  assign n1877 = ~n1869 & ~n1870 ;
  assign n1871 = \i_tv80_core_i_reg_RegsL_reg[6][0]/P0001  & n1285 ;
  assign n1872 = \i_tv80_core_i_reg_RegsL_reg[5][0]/P0001  & n1287 ;
  assign n1878 = ~n1871 & ~n1872 ;
  assign n1882 = n1877 & n1878 ;
  assign n1883 = n1881 & n1882 ;
  assign n1884 = n1277 & ~n1883 ;
  assign n1885 = \i_tv80_core_TmpAddr_reg[0]/P0001  & ~n1314 ;
  assign n1886 = n1314 & ~n1331 ;
  assign n1887 = \i_tv80_core_TmpAddr_reg[0]/P0001  & n1317 ;
  assign n1890 = ~\i_tv80_core_TmpAddr_reg[0]/P0001  & ~n1599 ;
  assign n1891 = ~\i_tv80_core_PC_reg[0]/P0001  & n1599 ;
  assign n1892 = ~n1890 & ~n1891 ;
  assign n1893 = ~n1593 & ~n1892 ;
  assign n1889 = n1593 & n1883 ;
  assign n1894 = n1595 & ~n1889 ;
  assign n1895 = ~n1893 & n1894 ;
  assign n1897 = ~\i_tv80_core_TmpAddr_reg[0]/P0001  & ~n1578 ;
  assign n1898 = ~n1579 & ~n1897 ;
  assign n1899 = n1584 & n1898 ;
  assign n1888 = n1530 & ~n1883 ;
  assign n1896 = \i_tv80_core_PC_reg[0]/P0001  & n1571 ;
  assign n1902 = ~n1888 & ~n1896 ;
  assign n1903 = ~n1899 & n1902 ;
  assign n1900 = \di_reg_reg[0]/P0001  & n1589 ;
  assign n1901 = \i_tv80_core_SP_reg[0]/P0001  & n1591 ;
  assign n1904 = ~n1900 & ~n1901 ;
  assign n1905 = n1903 & n1904 ;
  assign n1906 = ~n1895 & n1905 ;
  assign n1907 = ~n1317 & ~n1906 ;
  assign n1908 = ~n1887 & ~n1907 ;
  assign n1909 = n1886 & ~n1908 ;
  assign n1910 = ~n1885 & ~n1909 ;
  assign n1911 = ~n1277 & ~n1910 ;
  assign n1912 = ~n1884 & ~n1911 ;
  assign n1913 = n1625 & ~n1912 ;
  assign n1914 = \i_tv80_core_TmpAddr_reg[0]/P0001  & ~n1625 ;
  assign n1915 = n1103 & ~n1914 ;
  assign n1916 = ~n1913 & n1915 ;
  assign n1917 = ~\A[0]_pad  & ~n1103 ;
  assign n1918 = ~n1113 & ~n1917 ;
  assign n1919 = ~n1916 & n1918 ;
  assign n1921 = ~\i_tv80_core_R_reg[0]/P0001  & n1635 ;
  assign n1920 = ~\A[0]_pad  & ~n1635 ;
  assign n1922 = n1113 & ~n1920 ;
  assign n1923 = ~n1921 & n1922 ;
  assign n1924 = ~\i_tv80_core_BusAck_reg/P0001  & ~n1923 ;
  assign n1925 = ~n1919 & n1924 ;
  assign n1926 = ~\A[0]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n1927 = reset_n_pad & ~n1926 ;
  assign n1928 = ~n1925 & n1927 ;
  assign n1929 = \i_tv80_core_I_reg[2]/P0001  & n1317 ;
  assign n1935 = \i_tv80_core_i_reg_RegsH_reg[6][2]/P0001  & n1285 ;
  assign n1936 = \i_tv80_core_i_reg_RegsH_reg[5][2]/P0001  & n1287 ;
  assign n1941 = ~n1935 & ~n1936 ;
  assign n1937 = \i_tv80_core_i_reg_RegsH_reg[7][2]/P0001  & n1294 ;
  assign n1938 = \i_tv80_core_i_reg_RegsH_reg[3][2]/P0001  & n1296 ;
  assign n1942 = ~n1937 & ~n1938 ;
  assign n1943 = n1941 & n1942 ;
  assign n1931 = \i_tv80_core_i_reg_RegsH_reg[0][2]/P0001  & n1279 ;
  assign n1932 = \i_tv80_core_i_reg_RegsH_reg[4][2]/P0001  & n1282 ;
  assign n1939 = ~n1931 & ~n1932 ;
  assign n1933 = \i_tv80_core_i_reg_RegsH_reg[2][2]/P0001  & n1290 ;
  assign n1934 = \i_tv80_core_i_reg_RegsH_reg[1][2]/P0001  & n1292 ;
  assign n1940 = ~n1933 & ~n1934 ;
  assign n1944 = n1939 & n1940 ;
  assign n1945 = n1943 & n1944 ;
  assign n1946 = n1593 & ~n1945 ;
  assign n1948 = ~\i_tv80_core_PC_reg[10]/P0001  & n1599 ;
  assign n1947 = ~\i_tv80_core_TmpAddr_reg[10]/P0001  & ~n1599 ;
  assign n1949 = ~n1593 & ~n1947 ;
  assign n1950 = ~n1948 & n1949 ;
  assign n1951 = ~n1946 & ~n1950 ;
  assign n1952 = n1595 & ~n1951 ;
  assign n1930 = \i_tv80_core_SP_reg[10]/P0001  & n1591 ;
  assign n1953 = \i_tv80_core_PC_reg[10]/P0001  & n1571 ;
  assign n1970 = n1530 & ~n1945 ;
  assign n1971 = ~n1953 & ~n1970 ;
  assign n1972 = ~n1930 & n1971 ;
  assign n1954 = ~\di_reg_reg[2]/P0001  & ~n1578 ;
  assign n1956 = \i_tv80_core_TmpAddr_reg[4]/P0001  & \i_tv80_core_TmpAddr_reg[5]/P0001  ;
  assign n1957 = \i_tv80_core_TmpAddr_reg[6]/P0001  & \i_tv80_core_TmpAddr_reg[7]/P0001  ;
  assign n1958 = n1956 & n1957 ;
  assign n1955 = \i_tv80_core_TmpAddr_reg[0]/P0001  & \i_tv80_core_TmpAddr_reg[1]/P0001  ;
  assign n1959 = n1722 & n1955 ;
  assign n1960 = n1958 & n1959 ;
  assign n1961 = \i_tv80_core_TmpAddr_reg[8]/P0001  & n1960 ;
  assign n1962 = \i_tv80_core_TmpAddr_reg[9]/P0001  & n1961 ;
  assign n1963 = ~\i_tv80_core_TmpAddr_reg[10]/P0001  & ~n1962 ;
  assign n1964 = \i_tv80_core_TmpAddr_reg[10]/P0001  & n1962 ;
  assign n1965 = ~n1963 & ~n1964 ;
  assign n1966 = n1578 & ~n1965 ;
  assign n1967 = ~n1954 & ~n1966 ;
  assign n1968 = n1584 & n1967 ;
  assign n1969 = \i_tv80_core_ACC_reg[2]/P0001  & n1589 ;
  assign n1973 = ~n1968 & ~n1969 ;
  assign n1974 = n1972 & n1973 ;
  assign n1975 = ~n1952 & n1974 ;
  assign n1976 = ~n1317 & ~n1975 ;
  assign n1977 = ~n1929 & ~n1976 ;
  assign n1978 = n1886 & ~n1977 ;
  assign n1979 = \i_tv80_core_TmpAddr_reg[10]/P0001  & ~n1314 ;
  assign n1980 = ~n1978 & ~n1979 ;
  assign n1981 = ~n1277 & ~n1980 ;
  assign n1982 = n1277 & ~n1945 ;
  assign n1983 = ~n1981 & ~n1982 ;
  assign n1984 = n1625 & ~n1983 ;
  assign n1985 = \di_reg_reg[2]/P0001  & ~n1625 ;
  assign n1986 = n1103 & ~n1985 ;
  assign n1987 = ~n1984 & n1986 ;
  assign n1988 = ~\A[10]_pad  & ~n1103 ;
  assign n1989 = ~n1113 & ~n1988 ;
  assign n1990 = ~n1987 & n1989 ;
  assign n1992 = ~\i_tv80_core_I_reg[2]/P0001  & n1635 ;
  assign n1991 = ~\A[10]_pad  & ~n1635 ;
  assign n1993 = n1113 & ~n1991 ;
  assign n1994 = ~n1992 & n1993 ;
  assign n1995 = ~\i_tv80_core_BusAck_reg/P0001  & ~n1994 ;
  assign n1996 = ~n1990 & n1995 ;
  assign n1997 = ~\A[10]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n1998 = reset_n_pad & ~n1997 ;
  assign n1999 = ~n1996 & n1998 ;
  assign n2000 = \i_tv80_core_I_reg[3]/P0001  & n1317 ;
  assign n2006 = \i_tv80_core_i_reg_RegsH_reg[6][3]/P0001  & n1285 ;
  assign n2007 = \i_tv80_core_i_reg_RegsH_reg[5][3]/P0001  & n1287 ;
  assign n2012 = ~n2006 & ~n2007 ;
  assign n2008 = \i_tv80_core_i_reg_RegsH_reg[7][3]/P0001  & n1294 ;
  assign n2009 = \i_tv80_core_i_reg_RegsH_reg[3][3]/P0001  & n1296 ;
  assign n2013 = ~n2008 & ~n2009 ;
  assign n2014 = n2012 & n2013 ;
  assign n2002 = \i_tv80_core_i_reg_RegsH_reg[0][3]/P0001  & n1279 ;
  assign n2003 = \i_tv80_core_i_reg_RegsH_reg[4][3]/P0001  & n1282 ;
  assign n2010 = ~n2002 & ~n2003 ;
  assign n2004 = \i_tv80_core_i_reg_RegsH_reg[2][3]/P0001  & n1290 ;
  assign n2005 = \i_tv80_core_i_reg_RegsH_reg[1][3]/P0001  & n1292 ;
  assign n2011 = ~n2004 & ~n2005 ;
  assign n2015 = n2010 & n2011 ;
  assign n2016 = n2014 & n2015 ;
  assign n2017 = n1593 & ~n2016 ;
  assign n2019 = ~\i_tv80_core_PC_reg[11]/P0001  & n1599 ;
  assign n2018 = ~\i_tv80_core_TmpAddr_reg[11]/P0001  & ~n1599 ;
  assign n2020 = ~n1593 & ~n2018 ;
  assign n2021 = ~n2019 & n2020 ;
  assign n2022 = ~n2017 & ~n2021 ;
  assign n2023 = n1595 & ~n2022 ;
  assign n2001 = \i_tv80_core_SP_reg[11]/P0001  & n1591 ;
  assign n2024 = \i_tv80_core_PC_reg[11]/P0001  & n1571 ;
  assign n2033 = n1530 & ~n2016 ;
  assign n2034 = ~n2024 & ~n2033 ;
  assign n2035 = ~n2001 & n2034 ;
  assign n2025 = ~\di_reg_reg[3]/P0001  & ~n1578 ;
  assign n2026 = ~\i_tv80_core_TmpAddr_reg[11]/P0001  & ~n1964 ;
  assign n2027 = \i_tv80_core_TmpAddr_reg[11]/P0001  & n1964 ;
  assign n2028 = ~n2026 & ~n2027 ;
  assign n2029 = n1578 & ~n2028 ;
  assign n2030 = ~n2025 & ~n2029 ;
  assign n2031 = n1584 & n2030 ;
  assign n2032 = \i_tv80_core_ACC_reg[3]/P0001  & n1589 ;
  assign n2036 = ~n2031 & ~n2032 ;
  assign n2037 = n2035 & n2036 ;
  assign n2038 = ~n2023 & n2037 ;
  assign n2039 = ~n1317 & ~n2038 ;
  assign n2040 = ~n2000 & ~n2039 ;
  assign n2041 = n1886 & ~n2040 ;
  assign n2042 = \i_tv80_core_TmpAddr_reg[11]/P0001  & ~n1314 ;
  assign n2043 = ~n2041 & ~n2042 ;
  assign n2044 = ~n1277 & ~n2043 ;
  assign n2045 = n1277 & ~n2016 ;
  assign n2046 = ~n2044 & ~n2045 ;
  assign n2047 = n1625 & ~n2046 ;
  assign n2048 = \di_reg_reg[3]/P0001  & ~n1625 ;
  assign n2049 = n1103 & ~n2048 ;
  assign n2050 = ~n2047 & n2049 ;
  assign n2051 = ~\A[11]_pad  & ~n1103 ;
  assign n2052 = ~n1113 & ~n2051 ;
  assign n2053 = ~n2050 & n2052 ;
  assign n2055 = ~\i_tv80_core_I_reg[3]/P0001  & n1635 ;
  assign n2054 = ~\A[11]_pad  & ~n1635 ;
  assign n2056 = n1113 & ~n2054 ;
  assign n2057 = ~n2055 & n2056 ;
  assign n2058 = ~\i_tv80_core_BusAck_reg/P0001  & ~n2057 ;
  assign n2059 = ~n2053 & n2058 ;
  assign n2060 = ~\A[11]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n2061 = reset_n_pad & ~n2060 ;
  assign n2062 = ~n2059 & n2061 ;
  assign n2063 = \i_tv80_core_I_reg[4]/P0001  & n1317 ;
  assign n2069 = \i_tv80_core_i_reg_RegsH_reg[2][4]/P0001  & n1290 ;
  assign n2070 = \i_tv80_core_i_reg_RegsH_reg[1][4]/P0001  & n1292 ;
  assign n2075 = ~n2069 & ~n2070 ;
  assign n2071 = \i_tv80_core_i_reg_RegsH_reg[7][4]/P0001  & n1294 ;
  assign n2072 = \i_tv80_core_i_reg_RegsH_reg[3][4]/P0001  & n1296 ;
  assign n2076 = ~n2071 & ~n2072 ;
  assign n2077 = n2075 & n2076 ;
  assign n2065 = \i_tv80_core_i_reg_RegsH_reg[0][4]/P0001  & n1279 ;
  assign n2066 = \i_tv80_core_i_reg_RegsH_reg[4][4]/P0001  & n1282 ;
  assign n2073 = ~n2065 & ~n2066 ;
  assign n2067 = \i_tv80_core_i_reg_RegsH_reg[6][4]/P0001  & n1285 ;
  assign n2068 = \i_tv80_core_i_reg_RegsH_reg[5][4]/P0001  & n1287 ;
  assign n2074 = ~n2067 & ~n2068 ;
  assign n2078 = n2073 & n2074 ;
  assign n2079 = n2077 & n2078 ;
  assign n2080 = n1593 & ~n2079 ;
  assign n2082 = ~\i_tv80_core_PC_reg[12]/P0001  & n1599 ;
  assign n2081 = ~\i_tv80_core_TmpAddr_reg[12]/P0001  & ~n1599 ;
  assign n2083 = ~n1593 & ~n2081 ;
  assign n2084 = ~n2082 & n2083 ;
  assign n2085 = ~n2080 & ~n2084 ;
  assign n2086 = n1595 & ~n2085 ;
  assign n2064 = \i_tv80_core_SP_reg[12]/P0001  & n1591 ;
  assign n2087 = \i_tv80_core_PC_reg[12]/P0001  & n1571 ;
  assign n2096 = n1530 & ~n2079 ;
  assign n2097 = ~n2087 & ~n2096 ;
  assign n2098 = ~n2064 & n2097 ;
  assign n2088 = ~\di_reg_reg[4]/P0001  & ~n1578 ;
  assign n2089 = ~\i_tv80_core_TmpAddr_reg[12]/P0001  & ~n2027 ;
  assign n2090 = \i_tv80_core_TmpAddr_reg[12]/P0001  & n2027 ;
  assign n2091 = ~n2089 & ~n2090 ;
  assign n2092 = n1578 & ~n2091 ;
  assign n2093 = ~n2088 & ~n2092 ;
  assign n2094 = n1584 & n2093 ;
  assign n2095 = \i_tv80_core_ACC_reg[4]/P0001  & n1589 ;
  assign n2099 = ~n2094 & ~n2095 ;
  assign n2100 = n2098 & n2099 ;
  assign n2101 = ~n2086 & n2100 ;
  assign n2102 = ~n1317 & ~n2101 ;
  assign n2103 = ~n2063 & ~n2102 ;
  assign n2104 = n1886 & ~n2103 ;
  assign n2105 = \i_tv80_core_TmpAddr_reg[12]/P0001  & ~n1314 ;
  assign n2106 = ~n2104 & ~n2105 ;
  assign n2107 = ~n1277 & ~n2106 ;
  assign n2108 = n1277 & ~n2079 ;
  assign n2109 = ~n2107 & ~n2108 ;
  assign n2110 = n1625 & ~n2109 ;
  assign n2111 = \di_reg_reg[4]/P0001  & ~n1625 ;
  assign n2112 = n1103 & ~n2111 ;
  assign n2113 = ~n2110 & n2112 ;
  assign n2114 = ~\A[12]_pad  & ~n1103 ;
  assign n2115 = ~n1113 & ~n2114 ;
  assign n2116 = ~n2113 & n2115 ;
  assign n2118 = ~\i_tv80_core_I_reg[4]/P0001  & n1635 ;
  assign n2117 = ~\A[12]_pad  & ~n1635 ;
  assign n2119 = n1113 & ~n2117 ;
  assign n2120 = ~n2118 & n2119 ;
  assign n2121 = ~\i_tv80_core_BusAck_reg/P0001  & ~n2120 ;
  assign n2122 = ~n2116 & n2121 ;
  assign n2123 = ~\A[12]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n2124 = reset_n_pad & ~n2123 ;
  assign n2125 = ~n2122 & n2124 ;
  assign n2126 = \i_tv80_core_I_reg[5]/P0001  & n1317 ;
  assign n2132 = \i_tv80_core_i_reg_RegsH_reg[6][5]/P0001  & n1285 ;
  assign n2133 = \i_tv80_core_i_reg_RegsH_reg[5][5]/P0001  & n1287 ;
  assign n2138 = ~n2132 & ~n2133 ;
  assign n2134 = \i_tv80_core_i_reg_RegsH_reg[7][5]/P0001  & n1294 ;
  assign n2135 = \i_tv80_core_i_reg_RegsH_reg[3][5]/P0001  & n1296 ;
  assign n2139 = ~n2134 & ~n2135 ;
  assign n2140 = n2138 & n2139 ;
  assign n2128 = \i_tv80_core_i_reg_RegsH_reg[0][5]/P0001  & n1279 ;
  assign n2129 = \i_tv80_core_i_reg_RegsH_reg[4][5]/P0001  & n1282 ;
  assign n2136 = ~n2128 & ~n2129 ;
  assign n2130 = \i_tv80_core_i_reg_RegsH_reg[2][5]/P0001  & n1290 ;
  assign n2131 = \i_tv80_core_i_reg_RegsH_reg[1][5]/P0001  & n1292 ;
  assign n2137 = ~n2130 & ~n2131 ;
  assign n2141 = n2136 & n2137 ;
  assign n2142 = n2140 & n2141 ;
  assign n2143 = n1593 & ~n2142 ;
  assign n2145 = ~\i_tv80_core_PC_reg[13]/P0001  & n1599 ;
  assign n2144 = ~\i_tv80_core_TmpAddr_reg[13]/P0001  & ~n1599 ;
  assign n2146 = ~n1593 & ~n2144 ;
  assign n2147 = ~n2145 & n2146 ;
  assign n2148 = ~n2143 & ~n2147 ;
  assign n2149 = n1595 & ~n2148 ;
  assign n2127 = \i_tv80_core_SP_reg[13]/P0001  & n1591 ;
  assign n2150 = \i_tv80_core_PC_reg[13]/P0001  & n1571 ;
  assign n2159 = n1530 & ~n2142 ;
  assign n2160 = ~n2150 & ~n2159 ;
  assign n2161 = ~n2127 & n2160 ;
  assign n2151 = ~\di_reg_reg[5]/P0001  & ~n1578 ;
  assign n2152 = ~\i_tv80_core_TmpAddr_reg[13]/P0001  & ~n2090 ;
  assign n2153 = \i_tv80_core_TmpAddr_reg[13]/P0001  & n2090 ;
  assign n2154 = ~n2152 & ~n2153 ;
  assign n2155 = n1578 & ~n2154 ;
  assign n2156 = ~n2151 & ~n2155 ;
  assign n2157 = n1584 & n2156 ;
  assign n2158 = \i_tv80_core_ACC_reg[5]/P0001  & n1589 ;
  assign n2162 = ~n2157 & ~n2158 ;
  assign n2163 = n2161 & n2162 ;
  assign n2164 = ~n2149 & n2163 ;
  assign n2165 = ~n1317 & ~n2164 ;
  assign n2166 = ~n2126 & ~n2165 ;
  assign n2167 = n1886 & ~n2166 ;
  assign n2168 = \i_tv80_core_TmpAddr_reg[13]/P0001  & ~n1314 ;
  assign n2169 = ~n2167 & ~n2168 ;
  assign n2170 = ~n1277 & ~n2169 ;
  assign n2171 = n1277 & ~n2142 ;
  assign n2172 = ~n2170 & ~n2171 ;
  assign n2173 = n1625 & ~n2172 ;
  assign n2174 = \di_reg_reg[5]/P0001  & ~n1625 ;
  assign n2175 = n1103 & ~n2174 ;
  assign n2176 = ~n2173 & n2175 ;
  assign n2177 = ~\A[13]_pad  & ~n1103 ;
  assign n2178 = ~n1113 & ~n2177 ;
  assign n2179 = ~n2176 & n2178 ;
  assign n2181 = ~\i_tv80_core_I_reg[5]/P0001  & n1635 ;
  assign n2180 = ~\A[13]_pad  & ~n1635 ;
  assign n2182 = n1113 & ~n2180 ;
  assign n2183 = ~n2181 & n2182 ;
  assign n2184 = ~\i_tv80_core_BusAck_reg/P0001  & ~n2183 ;
  assign n2185 = ~n2179 & n2184 ;
  assign n2186 = ~\A[13]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n2187 = reset_n_pad & ~n2186 ;
  assign n2188 = ~n2185 & n2187 ;
  assign n2189 = \i_tv80_core_I_reg[6]/P0001  & n1317 ;
  assign n2195 = \i_tv80_core_i_reg_RegsH_reg[6][6]/P0001  & n1285 ;
  assign n2196 = \i_tv80_core_i_reg_RegsH_reg[5][6]/P0001  & n1287 ;
  assign n2201 = ~n2195 & ~n2196 ;
  assign n2197 = \i_tv80_core_i_reg_RegsH_reg[7][6]/P0001  & n1294 ;
  assign n2198 = \i_tv80_core_i_reg_RegsH_reg[3][6]/P0001  & n1296 ;
  assign n2202 = ~n2197 & ~n2198 ;
  assign n2203 = n2201 & n2202 ;
  assign n2191 = \i_tv80_core_i_reg_RegsH_reg[0][6]/P0001  & n1279 ;
  assign n2192 = \i_tv80_core_i_reg_RegsH_reg[4][6]/P0001  & n1282 ;
  assign n2199 = ~n2191 & ~n2192 ;
  assign n2193 = \i_tv80_core_i_reg_RegsH_reg[2][6]/P0001  & n1290 ;
  assign n2194 = \i_tv80_core_i_reg_RegsH_reg[1][6]/P0001  & n1292 ;
  assign n2200 = ~n2193 & ~n2194 ;
  assign n2204 = n2199 & n2200 ;
  assign n2205 = n2203 & n2204 ;
  assign n2206 = n1593 & ~n2205 ;
  assign n2208 = ~\i_tv80_core_PC_reg[14]/P0001  & n1599 ;
  assign n2207 = ~\i_tv80_core_TmpAddr_reg[14]/P0001  & ~n1599 ;
  assign n2209 = ~n1593 & ~n2207 ;
  assign n2210 = ~n2208 & n2209 ;
  assign n2211 = ~n2206 & ~n2210 ;
  assign n2212 = n1595 & ~n2211 ;
  assign n2190 = \i_tv80_core_SP_reg[14]/P0001  & n1591 ;
  assign n2213 = \i_tv80_core_PC_reg[14]/P0001  & n1571 ;
  assign n2222 = n1530 & ~n2205 ;
  assign n2223 = ~n2213 & ~n2222 ;
  assign n2224 = ~n2190 & n2223 ;
  assign n2214 = ~\di_reg_reg[6]/P0001  & ~n1578 ;
  assign n2215 = ~\i_tv80_core_TmpAddr_reg[14]/P0001  & ~n2153 ;
  assign n2216 = \i_tv80_core_TmpAddr_reg[14]/P0001  & n2153 ;
  assign n2217 = ~n2215 & ~n2216 ;
  assign n2218 = n1578 & ~n2217 ;
  assign n2219 = ~n2214 & ~n2218 ;
  assign n2220 = n1584 & n2219 ;
  assign n2221 = \i_tv80_core_ACC_reg[6]/P0001  & n1589 ;
  assign n2225 = ~n2220 & ~n2221 ;
  assign n2226 = n2224 & n2225 ;
  assign n2227 = ~n2212 & n2226 ;
  assign n2228 = ~n1317 & ~n2227 ;
  assign n2229 = ~n2189 & ~n2228 ;
  assign n2230 = n1886 & ~n2229 ;
  assign n2231 = \i_tv80_core_TmpAddr_reg[14]/P0001  & ~n1314 ;
  assign n2232 = ~n2230 & ~n2231 ;
  assign n2233 = ~n1277 & ~n2232 ;
  assign n2234 = n1277 & ~n2205 ;
  assign n2235 = ~n2233 & ~n2234 ;
  assign n2236 = n1625 & ~n2235 ;
  assign n2237 = \di_reg_reg[6]/P0001  & ~n1625 ;
  assign n2238 = n1103 & ~n2237 ;
  assign n2239 = ~n2236 & n2238 ;
  assign n2240 = ~\A[14]_pad  & ~n1103 ;
  assign n2241 = ~n1113 & ~n2240 ;
  assign n2242 = ~n2239 & n2241 ;
  assign n2244 = ~\i_tv80_core_I_reg[6]/P0001  & n1635 ;
  assign n2243 = ~\A[14]_pad  & ~n1635 ;
  assign n2245 = n1113 & ~n2243 ;
  assign n2246 = ~n2244 & n2245 ;
  assign n2247 = ~\i_tv80_core_BusAck_reg/P0001  & ~n2246 ;
  assign n2248 = ~n2242 & n2247 ;
  assign n2249 = ~\A[14]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n2250 = reset_n_pad & ~n2249 ;
  assign n2251 = ~n2248 & n2250 ;
  assign n2252 = \i_tv80_core_I_reg[7]/P0001  & n1317 ;
  assign n2258 = \i_tv80_core_i_reg_RegsH_reg[6][7]/P0002  & n1285 ;
  assign n2259 = \i_tv80_core_i_reg_RegsH_reg[5][7]/P0002  & n1287 ;
  assign n2264 = ~n2258 & ~n2259 ;
  assign n2260 = \i_tv80_core_i_reg_RegsH_reg[2][7]/P0002  & n1290 ;
  assign n2261 = \i_tv80_core_i_reg_RegsH_reg[3][7]/P0002  & n1296 ;
  assign n2265 = ~n2260 & ~n2261 ;
  assign n2266 = n2264 & n2265 ;
  assign n2254 = \i_tv80_core_i_reg_RegsH_reg[1][7]/P0002  & n1292 ;
  assign n2255 = \i_tv80_core_i_reg_RegsH_reg[4][7]/P0002  & n1282 ;
  assign n2262 = ~n2254 & ~n2255 ;
  assign n2256 = \i_tv80_core_i_reg_RegsH_reg[7][7]/P0002  & n1294 ;
  assign n2257 = \i_tv80_core_i_reg_RegsH_reg[0][7]/P0002  & n1279 ;
  assign n2263 = ~n2256 & ~n2257 ;
  assign n2267 = n2262 & n2263 ;
  assign n2268 = n2266 & n2267 ;
  assign n2269 = n1593 & ~n2268 ;
  assign n2271 = ~\i_tv80_core_PC_reg[15]/P0001  & n1599 ;
  assign n2270 = ~\i_tv80_core_TmpAddr_reg[15]/P0001  & ~n1599 ;
  assign n2272 = ~n1593 & ~n2270 ;
  assign n2273 = ~n2271 & n2272 ;
  assign n2274 = ~n2269 & ~n2273 ;
  assign n2275 = n1595 & ~n2274 ;
  assign n2253 = \i_tv80_core_SP_reg[15]/P0001  & n1591 ;
  assign n2276 = \i_tv80_core_PC_reg[15]/P0001  & n1571 ;
  assign n2285 = n1530 & ~n2268 ;
  assign n2286 = ~n2276 & ~n2285 ;
  assign n2287 = ~n2253 & n2286 ;
  assign n2277 = ~\di_reg_reg[7]/P0001  & ~n1578 ;
  assign n2278 = ~\i_tv80_core_TmpAddr_reg[15]/P0001  & ~n2216 ;
  assign n2279 = \i_tv80_core_TmpAddr_reg[15]/P0001  & n2216 ;
  assign n2280 = ~n2278 & ~n2279 ;
  assign n2281 = n1578 & ~n2280 ;
  assign n2282 = ~n2277 & ~n2281 ;
  assign n2283 = n1584 & n2282 ;
  assign n2284 = \i_tv80_core_ACC_reg[7]/P0001  & n1589 ;
  assign n2288 = ~n2283 & ~n2284 ;
  assign n2289 = n2287 & n2288 ;
  assign n2290 = ~n2275 & n2289 ;
  assign n2291 = ~n1317 & ~n2290 ;
  assign n2292 = ~n2252 & ~n2291 ;
  assign n2293 = n1886 & ~n2292 ;
  assign n2294 = \i_tv80_core_TmpAddr_reg[15]/P0001  & ~n1314 ;
  assign n2295 = ~n2293 & ~n2294 ;
  assign n2296 = ~n1277 & ~n2295 ;
  assign n2297 = n1277 & ~n2268 ;
  assign n2298 = ~n2296 & ~n2297 ;
  assign n2299 = n1625 & ~n2298 ;
  assign n2300 = \di_reg_reg[7]/P0001  & ~n1625 ;
  assign n2301 = n1103 & ~n2300 ;
  assign n2302 = ~n2299 & n2301 ;
  assign n2303 = ~\A[15]_pad  & ~n1103 ;
  assign n2304 = ~n1113 & ~n2303 ;
  assign n2305 = ~n2302 & n2304 ;
  assign n2307 = ~\i_tv80_core_I_reg[7]/P0001  & n1635 ;
  assign n2306 = ~\A[15]_pad  & ~n1635 ;
  assign n2308 = n1113 & ~n2306 ;
  assign n2309 = ~n2307 & n2308 ;
  assign n2310 = ~\i_tv80_core_BusAck_reg/P0001  & ~n2309 ;
  assign n2311 = ~n2305 & n2310 ;
  assign n2312 = ~\A[15]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n2313 = reset_n_pad & ~n2312 ;
  assign n2314 = ~n2311 & n2313 ;
  assign n2315 = \i_tv80_core_TmpAddr_reg[3]/P0001  & n1317 ;
  assign n2320 = \i_tv80_core_i_reg_RegsL_reg[6][3]/NET0131  & n1285 ;
  assign n2321 = \i_tv80_core_i_reg_RegsL_reg[5][3]/NET0131  & n1287 ;
  assign n2326 = ~n2320 & ~n2321 ;
  assign n2322 = \i_tv80_core_i_reg_RegsL_reg[2][3]/NET0131  & n1290 ;
  assign n2323 = \i_tv80_core_i_reg_RegsL_reg[0][3]/NET0131  & n1279 ;
  assign n2327 = ~n2322 & ~n2323 ;
  assign n2328 = n2326 & n2327 ;
  assign n2316 = \i_tv80_core_i_reg_RegsL_reg[1][3]/NET0131  & n1292 ;
  assign n2317 = \i_tv80_core_i_reg_RegsL_reg[7][3]/NET0131  & n1294 ;
  assign n2324 = ~n2316 & ~n2317 ;
  assign n2318 = \i_tv80_core_i_reg_RegsL_reg[4][3]/NET0131  & n1282 ;
  assign n2319 = \i_tv80_core_i_reg_RegsL_reg[3][3]/NET0131  & n1296 ;
  assign n2325 = ~n2318 & ~n2319 ;
  assign n2329 = n2324 & n2325 ;
  assign n2330 = n2328 & n2329 ;
  assign n2332 = n1593 & ~n2330 ;
  assign n2334 = ~\i_tv80_core_PC_reg[3]/P0001  & n1599 ;
  assign n2333 = ~\i_tv80_core_TmpAddr_reg[3]/P0001  & ~n1599 ;
  assign n2335 = ~n1593 & ~n2333 ;
  assign n2336 = ~n2334 & n2335 ;
  assign n2337 = ~n2332 & ~n2336 ;
  assign n2338 = n1595 & ~n2337 ;
  assign n2340 = ~\i_tv80_core_TmpAddr_reg[3]/P0001  & ~n1585 ;
  assign n2341 = ~n1723 & ~n2340 ;
  assign n2342 = n1584 & n2341 ;
  assign n2331 = n1530 & ~n2330 ;
  assign n2339 = \i_tv80_core_PC_reg[3]/P0001  & n1571 ;
  assign n2345 = ~n2331 & ~n2339 ;
  assign n2346 = ~n2342 & n2345 ;
  assign n2343 = \di_reg_reg[3]/P0001  & n1589 ;
  assign n2344 = \i_tv80_core_SP_reg[3]/P0001  & n1591 ;
  assign n2347 = ~n2343 & ~n2344 ;
  assign n2348 = n2346 & n2347 ;
  assign n2349 = ~n2338 & n2348 ;
  assign n2350 = ~n1317 & ~n2349 ;
  assign n2351 = ~n2315 & ~n2350 ;
  assign n2352 = n1886 & ~n2351 ;
  assign n2353 = \i_tv80_core_TmpAddr_reg[3]/P0001  & ~n1314 ;
  assign n2354 = ~n2352 & ~n2353 ;
  assign n2355 = ~n1277 & ~n2354 ;
  assign n2356 = n1277 & ~n2330 ;
  assign n2357 = ~n2355 & ~n2356 ;
  assign n2358 = n1625 & ~n2357 ;
  assign n2359 = \i_tv80_core_TmpAddr_reg[3]/P0001  & ~n1625 ;
  assign n2360 = n1103 & ~n2359 ;
  assign n2361 = ~n2358 & n2360 ;
  assign n2362 = ~\A[3]_pad  & ~n1103 ;
  assign n2363 = ~n1113 & ~n2362 ;
  assign n2364 = ~n2361 & n2363 ;
  assign n2366 = ~\i_tv80_core_R_reg[3]/P0001  & n1635 ;
  assign n2365 = ~\A[3]_pad  & ~n1635 ;
  assign n2367 = n1113 & ~n2365 ;
  assign n2368 = ~n2366 & n2367 ;
  assign n2369 = ~\i_tv80_core_BusAck_reg/P0001  & ~n2368 ;
  assign n2370 = ~n2364 & n2369 ;
  assign n2371 = ~\A[3]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n2372 = reset_n_pad & ~n2371 ;
  assign n2373 = ~n2370 & n2372 ;
  assign n2374 = \i_tv80_core_TmpAddr_reg[4]/P0001  & n1317 ;
  assign n2379 = \i_tv80_core_i_reg_RegsL_reg[2][4]/NET0131  & n1290 ;
  assign n2380 = \i_tv80_core_i_reg_RegsL_reg[1][4]/NET0131  & n1292 ;
  assign n2385 = ~n2379 & ~n2380 ;
  assign n2381 = \i_tv80_core_i_reg_RegsL_reg[7][4]/NET0131  & n1294 ;
  assign n2382 = \i_tv80_core_i_reg_RegsL_reg[3][4]/NET0131  & n1296 ;
  assign n2386 = ~n2381 & ~n2382 ;
  assign n2387 = n2385 & n2386 ;
  assign n2375 = \i_tv80_core_i_reg_RegsL_reg[0][4]/NET0131  & n1279 ;
  assign n2376 = \i_tv80_core_i_reg_RegsL_reg[4][4]/NET0131  & n1282 ;
  assign n2383 = ~n2375 & ~n2376 ;
  assign n2377 = \i_tv80_core_i_reg_RegsL_reg[6][4]/NET0131  & n1285 ;
  assign n2378 = \i_tv80_core_i_reg_RegsL_reg[5][4]/NET0131  & n1287 ;
  assign n2384 = ~n2377 & ~n2378 ;
  assign n2388 = n2383 & n2384 ;
  assign n2389 = n2387 & n2388 ;
  assign n2391 = n1593 & ~n2389 ;
  assign n2393 = ~\i_tv80_core_PC_reg[4]/P0001  & n1599 ;
  assign n2392 = ~\i_tv80_core_TmpAddr_reg[4]/P0001  & ~n1599 ;
  assign n2394 = ~n1593 & ~n2392 ;
  assign n2395 = ~n2393 & n2394 ;
  assign n2396 = ~n2391 & ~n2395 ;
  assign n2397 = n1595 & ~n2396 ;
  assign n2399 = ~\i_tv80_core_TmpAddr_reg[4]/P0001  & ~n1723 ;
  assign n2400 = ~n1724 & ~n2399 ;
  assign n2401 = n1584 & n2400 ;
  assign n2390 = n1530 & ~n2389 ;
  assign n2398 = \i_tv80_core_PC_reg[4]/P0001  & n1571 ;
  assign n2404 = ~n2390 & ~n2398 ;
  assign n2405 = ~n2401 & n2404 ;
  assign n2402 = \di_reg_reg[4]/P0001  & n1589 ;
  assign n2403 = \i_tv80_core_SP_reg[4]/P0001  & n1591 ;
  assign n2406 = ~n2402 & ~n2403 ;
  assign n2407 = n2405 & n2406 ;
  assign n2408 = ~n2397 & n2407 ;
  assign n2409 = ~n1317 & ~n2408 ;
  assign n2410 = ~n2374 & ~n2409 ;
  assign n2411 = n1886 & ~n2410 ;
  assign n2412 = \i_tv80_core_TmpAddr_reg[4]/P0001  & ~n1314 ;
  assign n2413 = ~n2411 & ~n2412 ;
  assign n2414 = ~n1277 & ~n2413 ;
  assign n2415 = n1277 & ~n2389 ;
  assign n2416 = ~n2414 & ~n2415 ;
  assign n2417 = n1625 & ~n2416 ;
  assign n2418 = \i_tv80_core_TmpAddr_reg[4]/P0001  & ~n1625 ;
  assign n2419 = n1103 & ~n2418 ;
  assign n2420 = ~n2417 & n2419 ;
  assign n2421 = ~\A[4]_pad  & ~n1103 ;
  assign n2422 = ~n1113 & ~n2421 ;
  assign n2423 = ~n2420 & n2422 ;
  assign n2425 = ~\i_tv80_core_R_reg[4]/P0001  & n1635 ;
  assign n2424 = ~\A[4]_pad  & ~n1635 ;
  assign n2426 = n1113 & ~n2424 ;
  assign n2427 = ~n2425 & n2426 ;
  assign n2428 = ~\i_tv80_core_BusAck_reg/P0001  & ~n2427 ;
  assign n2429 = ~n2423 & n2428 ;
  assign n2430 = ~\A[4]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n2431 = reset_n_pad & ~n2430 ;
  assign n2432 = ~n2429 & n2431 ;
  assign n2433 = \i_tv80_core_TmpAddr_reg[7]/P0001  & n1317 ;
  assign n2455 = \i_tv80_core_TmpAddr_reg[7]/P0001  & ~n1599 ;
  assign n2454 = \i_tv80_core_PC_reg[7]/P0001  & n1599 ;
  assign n2456 = ~n1593 & ~n2454 ;
  assign n2457 = ~n2455 & n2456 ;
  assign n2438 = \i_tv80_core_i_reg_RegsL_reg[2][7]/NET0131  & n1290 ;
  assign n2439 = \i_tv80_core_i_reg_RegsL_reg[1][7]/NET0131  & n1292 ;
  assign n2444 = ~n2438 & ~n2439 ;
  assign n2440 = \i_tv80_core_i_reg_RegsL_reg[7][7]/NET0131  & n1294 ;
  assign n2441 = \i_tv80_core_i_reg_RegsL_reg[3][7]/NET0131  & n1296 ;
  assign n2445 = ~n2440 & ~n2441 ;
  assign n2446 = n2444 & n2445 ;
  assign n2434 = \i_tv80_core_i_reg_RegsL_reg[0][7]/NET0131  & n1279 ;
  assign n2435 = \i_tv80_core_i_reg_RegsL_reg[4][7]/NET0131  & n1282 ;
  assign n2442 = ~n2434 & ~n2435 ;
  assign n2436 = \i_tv80_core_i_reg_RegsL_reg[6][7]/NET0131  & n1285 ;
  assign n2437 = \i_tv80_core_i_reg_RegsL_reg[5][7]/NET0131  & n1287 ;
  assign n2443 = ~n2436 & ~n2437 ;
  assign n2447 = n2442 & n2443 ;
  assign n2448 = n2446 & n2447 ;
  assign n2453 = n1593 & n2448 ;
  assign n2458 = n1595 & ~n2453 ;
  assign n2459 = ~n2457 & n2458 ;
  assign n2451 = \di_reg_reg[7]/P0001  & n1589 ;
  assign n2449 = n1530 & ~n2448 ;
  assign n2450 = \i_tv80_core_PC_reg[7]/P0001  & n1571 ;
  assign n2464 = ~n2449 & ~n2450 ;
  assign n2465 = ~n2451 & n2464 ;
  assign n2452 = \i_tv80_core_SP_reg[7]/P0001  & n1591 ;
  assign n2460 = n1578 & n1960 ;
  assign n2461 = ~\i_tv80_core_TmpAddr_reg[7]/P0001  & ~n1784 ;
  assign n2462 = ~n2460 & ~n2461 ;
  assign n2463 = n1584 & n2462 ;
  assign n2466 = ~n2452 & ~n2463 ;
  assign n2467 = n2465 & n2466 ;
  assign n2468 = ~n2459 & n2467 ;
  assign n2469 = ~n1317 & ~n2468 ;
  assign n2470 = ~n2433 & ~n2469 ;
  assign n2471 = n1886 & ~n2470 ;
  assign n2472 = \i_tv80_core_TmpAddr_reg[7]/P0001  & ~n1314 ;
  assign n2473 = ~n2471 & ~n2472 ;
  assign n2474 = ~n1277 & ~n2473 ;
  assign n2475 = n1277 & ~n2448 ;
  assign n2476 = ~n2474 & ~n2475 ;
  assign n2477 = n1625 & ~n2476 ;
  assign n2478 = \i_tv80_core_TmpAddr_reg[7]/P0001  & ~n1625 ;
  assign n2479 = n1103 & ~n2478 ;
  assign n2480 = ~n2477 & n2479 ;
  assign n2481 = ~\A[7]_pad  & ~n1103 ;
  assign n2482 = ~n1113 & ~n2481 ;
  assign n2483 = ~n2480 & n2482 ;
  assign n2485 = ~\i_tv80_core_R_reg[7]/P0001  & n1635 ;
  assign n2484 = ~\A[7]_pad  & ~n1635 ;
  assign n2486 = n1113 & ~n2484 ;
  assign n2487 = ~n2485 & n2486 ;
  assign n2488 = ~\i_tv80_core_BusAck_reg/P0001  & ~n2487 ;
  assign n2489 = ~n2483 & n2488 ;
  assign n2490 = ~\A[7]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n2491 = reset_n_pad & ~n2490 ;
  assign n2492 = ~n2489 & n2491 ;
  assign n2493 = \i_tv80_core_I_reg[0]/P0001  & n1317 ;
  assign n2499 = \i_tv80_core_i_reg_RegsH_reg[2][0]/P0001  & n1290 ;
  assign n2500 = \i_tv80_core_i_reg_RegsH_reg[1][0]/P0001  & n1292 ;
  assign n2505 = ~n2499 & ~n2500 ;
  assign n2501 = \i_tv80_core_i_reg_RegsH_reg[7][0]/P0001  & n1294 ;
  assign n2502 = \i_tv80_core_i_reg_RegsH_reg[3][0]/P0001  & n1296 ;
  assign n2506 = ~n2501 & ~n2502 ;
  assign n2507 = n2505 & n2506 ;
  assign n2495 = \i_tv80_core_i_reg_RegsH_reg[0][0]/P0001  & n1279 ;
  assign n2496 = \i_tv80_core_i_reg_RegsH_reg[4][0]/P0001  & n1282 ;
  assign n2503 = ~n2495 & ~n2496 ;
  assign n2497 = \i_tv80_core_i_reg_RegsH_reg[6][0]/P0001  & n1285 ;
  assign n2498 = \i_tv80_core_i_reg_RegsH_reg[5][0]/P0001  & n1287 ;
  assign n2504 = ~n2497 & ~n2498 ;
  assign n2508 = n2503 & n2504 ;
  assign n2509 = n2507 & n2508 ;
  assign n2510 = n1593 & ~n2509 ;
  assign n2512 = ~\i_tv80_core_PC_reg[8]/P0001  & n1599 ;
  assign n2511 = ~\i_tv80_core_TmpAddr_reg[8]/P0001  & ~n1599 ;
  assign n2513 = ~n1593 & ~n2511 ;
  assign n2514 = ~n2512 & n2513 ;
  assign n2515 = ~n2510 & ~n2514 ;
  assign n2516 = n1595 & ~n2515 ;
  assign n2494 = \i_tv80_core_SP_reg[8]/P0001  & n1591 ;
  assign n2517 = \i_tv80_core_PC_reg[8]/P0001  & n1571 ;
  assign n2525 = n1530 & ~n2509 ;
  assign n2526 = ~n2517 & ~n2525 ;
  assign n2527 = ~n2494 & n2526 ;
  assign n2518 = ~\di_reg_reg[0]/P0001  & ~n1578 ;
  assign n2519 = ~\i_tv80_core_TmpAddr_reg[8]/P0001  & ~n1960 ;
  assign n2520 = ~n1961 & ~n2519 ;
  assign n2521 = n1578 & ~n2520 ;
  assign n2522 = ~n2518 & ~n2521 ;
  assign n2523 = n1584 & n2522 ;
  assign n2524 = \i_tv80_core_ACC_reg[0]/P0001  & n1589 ;
  assign n2528 = ~n2523 & ~n2524 ;
  assign n2529 = n2527 & n2528 ;
  assign n2530 = ~n2516 & n2529 ;
  assign n2531 = ~n1317 & ~n2530 ;
  assign n2532 = ~n2493 & ~n2531 ;
  assign n2533 = n1886 & ~n2532 ;
  assign n2534 = \i_tv80_core_TmpAddr_reg[8]/P0001  & ~n1314 ;
  assign n2535 = ~n2533 & ~n2534 ;
  assign n2536 = ~n1277 & ~n2535 ;
  assign n2537 = n1277 & ~n2509 ;
  assign n2538 = ~n2536 & ~n2537 ;
  assign n2539 = n1625 & ~n2538 ;
  assign n2540 = \di_reg_reg[0]/P0001  & ~n1625 ;
  assign n2541 = n1103 & ~n2540 ;
  assign n2542 = ~n2539 & n2541 ;
  assign n2543 = ~\A[8]_pad  & ~n1103 ;
  assign n2544 = ~n1113 & ~n2543 ;
  assign n2545 = ~n2542 & n2544 ;
  assign n2547 = ~\i_tv80_core_I_reg[0]/P0001  & n1635 ;
  assign n2546 = ~\A[8]_pad  & ~n1635 ;
  assign n2548 = n1113 & ~n2546 ;
  assign n2549 = ~n2547 & n2548 ;
  assign n2550 = ~\i_tv80_core_BusAck_reg/P0001  & ~n2549 ;
  assign n2551 = ~n2545 & n2550 ;
  assign n2552 = ~\A[8]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n2553 = reset_n_pad & ~n2552 ;
  assign n2554 = ~n2551 & n2553 ;
  assign n2555 = \i_tv80_core_I_reg[1]/P0001  & n1317 ;
  assign n2561 = \i_tv80_core_i_reg_RegsH_reg[2][1]/P0001  & n1290 ;
  assign n2562 = \i_tv80_core_i_reg_RegsH_reg[1][1]/P0001  & n1292 ;
  assign n2567 = ~n2561 & ~n2562 ;
  assign n2563 = \i_tv80_core_i_reg_RegsH_reg[7][1]/P0001  & n1294 ;
  assign n2564 = \i_tv80_core_i_reg_RegsH_reg[3][1]/P0001  & n1296 ;
  assign n2568 = ~n2563 & ~n2564 ;
  assign n2569 = n2567 & n2568 ;
  assign n2557 = \i_tv80_core_i_reg_RegsH_reg[0][1]/P0001  & n1279 ;
  assign n2558 = \i_tv80_core_i_reg_RegsH_reg[4][1]/P0001  & n1282 ;
  assign n2565 = ~n2557 & ~n2558 ;
  assign n2559 = \i_tv80_core_i_reg_RegsH_reg[6][1]/P0001  & n1285 ;
  assign n2560 = \i_tv80_core_i_reg_RegsH_reg[5][1]/P0001  & n1287 ;
  assign n2566 = ~n2559 & ~n2560 ;
  assign n2570 = n2565 & n2566 ;
  assign n2571 = n2569 & n2570 ;
  assign n2572 = n1593 & ~n2571 ;
  assign n2574 = ~\i_tv80_core_PC_reg[9]/P0001  & n1599 ;
  assign n2573 = ~\i_tv80_core_TmpAddr_reg[9]/P0001  & ~n1599 ;
  assign n2575 = ~n1593 & ~n2573 ;
  assign n2576 = ~n2574 & n2575 ;
  assign n2577 = ~n2572 & ~n2576 ;
  assign n2578 = n1595 & ~n2577 ;
  assign n2556 = \i_tv80_core_SP_reg[9]/P0001  & n1591 ;
  assign n2579 = \i_tv80_core_PC_reg[9]/P0001  & n1571 ;
  assign n2587 = n1530 & ~n2571 ;
  assign n2588 = ~n2579 & ~n2587 ;
  assign n2589 = ~n2556 & n2588 ;
  assign n2580 = ~\di_reg_reg[1]/P0001  & ~n1578 ;
  assign n2581 = ~\i_tv80_core_TmpAddr_reg[9]/P0001  & ~n1961 ;
  assign n2582 = ~n1962 & ~n2581 ;
  assign n2583 = n1578 & ~n2582 ;
  assign n2584 = ~n2580 & ~n2583 ;
  assign n2585 = n1584 & n2584 ;
  assign n2586 = \i_tv80_core_ACC_reg[1]/P0001  & n1589 ;
  assign n2590 = ~n2585 & ~n2586 ;
  assign n2591 = n2589 & n2590 ;
  assign n2592 = ~n2578 & n2591 ;
  assign n2593 = ~n1317 & ~n2592 ;
  assign n2594 = ~n2555 & ~n2593 ;
  assign n2595 = n1886 & ~n2594 ;
  assign n2596 = \i_tv80_core_TmpAddr_reg[9]/P0001  & ~n1314 ;
  assign n2597 = ~n2595 & ~n2596 ;
  assign n2598 = ~n1277 & ~n2597 ;
  assign n2599 = n1277 & ~n2571 ;
  assign n2600 = ~n2598 & ~n2599 ;
  assign n2601 = n1625 & ~n2600 ;
  assign n2602 = \di_reg_reg[1]/P0001  & ~n1625 ;
  assign n2603 = n1103 & ~n2602 ;
  assign n2604 = ~n2601 & n2603 ;
  assign n2605 = ~\A[9]_pad  & ~n1103 ;
  assign n2606 = ~n1113 & ~n2605 ;
  assign n2607 = ~n2604 & n2606 ;
  assign n2609 = ~\i_tv80_core_I_reg[1]/P0001  & n1635 ;
  assign n2608 = ~\A[9]_pad  & ~n1635 ;
  assign n2610 = n1113 & ~n2608 ;
  assign n2611 = ~n2609 & n2610 ;
  assign n2612 = ~\i_tv80_core_BusAck_reg/P0001  & ~n2611 ;
  assign n2613 = ~n2607 & n2612 ;
  assign n2614 = ~\A[9]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n2615 = reset_n_pad & ~n2614 ;
  assign n2616 = ~n2613 & n2615 ;
  assign n2617 = n860 & n1107 ;
  assign n2618 = ~n1634 & ~n2617 ;
  assign n2624 = n970 & ~n1487 ;
  assign n2625 = n974 & ~n1482 ;
  assign n2626 = ~n2624 & n2625 ;
  assign n2631 = n929 & ~n930 ;
  assign n2632 = ~n939 & ~n2631 ;
  assign n2633 = n381 & ~n2632 ;
  assign n2627 = ~n856 & ~n1309 ;
  assign n2628 = \i_tv80_core_mcycle_reg[0]/P0001  & ~n2627 ;
  assign n2629 = n977 & n2628 ;
  assign n2630 = n856 & n1344 ;
  assign n2634 = ~n2629 & ~n2630 ;
  assign n2635 = ~n2633 & n2634 ;
  assign n2636 = ~n2626 & n2635 ;
  assign n2619 = n871 & ~n1482 ;
  assign n2620 = n381 & n948 ;
  assign n2621 = ~n2619 & ~n2620 ;
  assign n2622 = n856 & ~n945 ;
  assign n2623 = n2621 & ~n2622 ;
  assign n2637 = ~n1064 & n2623 ;
  assign n2638 = n2636 & n2637 ;
  assign n2639 = n382 & ~n2638 ;
  assign n2640 = n381 & n1012 ;
  assign n2641 = n856 & n1014 ;
  assign n2642 = n956 & n1466 ;
  assign n2643 = ~n2641 & ~n2642 ;
  assign n2644 = ~n2640 & n2643 ;
  assign n2645 = \i_tv80_core_ISet_reg[1]/P0001  & ~n2644 ;
  assign n2646 = ~n2639 & ~n2645 ;
  assign n2647 = ~n1634 & n2646 ;
  assign n2648 = ~n2618 & ~n2647 ;
  assign n2649 = n1593 & n2648 ;
  assign n2661 = ~\i_tv80_core_tstate_reg[0]/P0001  & ~\i_tv80_core_tstate_reg[1]/NET0131  ;
  assign n2662 = \i_tv80_core_tstate_reg[2]/NET0131  & n2661 ;
  assign n2663 = n382 & n2662 ;
  assign n2664 = n884 & n2663 ;
  assign n2665 = \i_tv80_core_RegAddrA_r_reg[1]/NET0131  & ~n2664 ;
  assign n2666 = n382 & n1107 ;
  assign n2667 = n884 & n2666 ;
  assign n2668 = ~n2665 & ~n2667 ;
  assign n2669 = ~n2649 & ~n2668 ;
  assign n2650 = \i_tv80_core_IR_reg[5]/P0001  & n1064 ;
  assign n2651 = n2623 & n2636 ;
  assign n2652 = ~n2650 & n2651 ;
  assign n2653 = n382 & ~n2652 ;
  assign n2655 = n857 & n1012 ;
  assign n2654 = n956 & n1006 ;
  assign n2656 = ~n2641 & ~n2654 ;
  assign n2657 = ~n2655 & n2656 ;
  assign n2658 = \i_tv80_core_ISet_reg[1]/P0001  & ~n2657 ;
  assign n2659 = ~n2653 & ~n2658 ;
  assign n2660 = n2649 & ~n2659 ;
  assign n2670 = \i_tv80_core_ISet_reg[1]/P0001  & ~n2643 ;
  assign n2671 = \i_tv80_core_IR_reg[4]/P0001  & n1064 ;
  assign n2672 = n2651 & ~n2671 ;
  assign n2673 = n382 & ~n2672 ;
  assign n2674 = ~n2670 & ~n2673 ;
  assign n2675 = ~n2659 & n2674 ;
  assign n2676 = n2648 & n2675 ;
  assign n2677 = ~n2660 & ~n2676 ;
  assign n2678 = ~n2669 & n2677 ;
  assign n2679 = n2649 & n2674 ;
  assign n2680 = ~\i_tv80_core_RegAddrA_r_reg[0]/NET0131  & ~n2664 ;
  assign n2681 = ~n2667 & ~n2680 ;
  assign n2682 = ~n2649 & ~n2681 ;
  assign n2683 = ~n2676 & n2682 ;
  assign n2684 = ~n2679 & ~n2683 ;
  assign n2685 = n2678 & ~n2684 ;
  assign n2686 = ~n2664 & ~n2667 ;
  assign n2687 = \i_tv80_core_Alternate_reg/P0001  & ~n2686 ;
  assign n2688 = \i_tv80_core_RegAddrA_r_reg[2]/NET0131  & n2686 ;
  assign n2689 = ~n2649 & n2688 ;
  assign n2690 = ~n2687 & ~n2689 ;
  assign n2691 = ~n2676 & ~n2690 ;
  assign n2692 = \i_tv80_core_Alternate_reg/P0001  & n2649 ;
  assign n2693 = \i_tv80_core_XY_State_reg[1]/P0001  & n2676 ;
  assign n2694 = ~n2692 & ~n2693 ;
  assign n2695 = ~n2691 & n2694 ;
  assign n2696 = n2685 & n2695 ;
  assign n2699 = ~n2659 & ~n2674 ;
  assign n2697 = n860 & ~n1107 ;
  assign n2698 = ~n2646 & ~n2697 ;
  assign n2700 = ~n860 & ~n1635 ;
  assign n2701 = n2698 & ~n2700 ;
  assign n2702 = ~n2699 & n2701 ;
  assign n2703 = \i_tv80_core_Read_To_Reg_r_reg[1]/P0001  & \i_tv80_core_Read_To_Reg_r_reg[2]/P0001  ;
  assign n2704 = ~\i_tv80_core_Read_To_Reg_r_reg[3]/P0001  & \i_tv80_core_Read_To_Reg_r_reg[4]/P0001  ;
  assign n2705 = ~n2703 & n2704 ;
  assign n2706 = \i_tv80_core_Read_To_Reg_r_reg[0]/P0001  & n2705 ;
  assign n2707 = n1162 & n2706 ;
  assign n2708 = n2686 & ~n2707 ;
  assign n2709 = ~n2702 & n2708 ;
  assign n2710 = ~\i_tv80_core_BusAck_reg/P0001  & ~n2709 ;
  assign n2711 = n2696 & n2710 ;
  assign n2712 = \i_tv80_core_IR_reg[0]/P0001  & n2655 ;
  assign n2713 = ~n2654 & ~n2712 ;
  assign n2714 = \i_tv80_core_IR_reg[3]/P0001  & ~n2713 ;
  assign n2715 = \i_tv80_core_IR_reg[0]/P0001  & n860 ;
  assign n2716 = ~\i_tv80_core_IR_reg[3]/P0001  & \i_tv80_core_mcycle_reg[1]/P0001  ;
  assign n2717 = ~\i_tv80_core_IR_reg[0]/P0001  & ~n2716 ;
  assign n2718 = n1083 & n2717 ;
  assign n2719 = ~n2715 & ~n2718 ;
  assign n2720 = n1012 & ~n2719 ;
  assign n2721 = ~n2714 & ~n2720 ;
  assign n2722 = \i_tv80_core_ISet_reg[1]/P0001  & ~n2721 ;
  assign n2723 = n977 & n1310 ;
  assign n2724 = ~n1065 & ~n2723 ;
  assign n2725 = n2621 & n2724 ;
  assign n2726 = ~n2633 & n2725 ;
  assign n2727 = ~n2626 & n2726 ;
  assign n2728 = n382 & ~n2727 ;
  assign n2729 = ~n2722 & ~n2728 ;
  assign n2738 = n2678 & n2684 ;
  assign n2741 = n2695 & n2738 ;
  assign n2742 = \i_tv80_core_i_reg_RegsL_reg[1][1]/P0001  & n2741 ;
  assign n2730 = ~n2678 & n2684 ;
  assign n2743 = n2695 & n2730 ;
  assign n2744 = \i_tv80_core_i_reg_RegsL_reg[3][1]/P0001  & n2743 ;
  assign n2750 = ~n2742 & ~n2744 ;
  assign n2735 = ~n2678 & ~n2684 ;
  assign n2745 = n2695 & n2735 ;
  assign n2746 = \i_tv80_core_i_reg_RegsL_reg[2][1]/P0001  & n2745 ;
  assign n2747 = \i_tv80_core_i_reg_RegsL_reg[0][1]/P0001  & n2696 ;
  assign n2751 = ~n2746 & ~n2747 ;
  assign n2752 = n2750 & n2751 ;
  assign n2731 = ~n2695 & n2730 ;
  assign n2732 = \i_tv80_core_i_reg_RegsL_reg[7][1]/P0001  & n2731 ;
  assign n2733 = n2685 & ~n2695 ;
  assign n2734 = \i_tv80_core_i_reg_RegsL_reg[4][1]/P0001  & n2733 ;
  assign n2748 = ~n2732 & ~n2734 ;
  assign n2736 = ~n2695 & n2735 ;
  assign n2737 = \i_tv80_core_i_reg_RegsL_reg[6][1]/P0001  & n2736 ;
  assign n2739 = ~n2695 & n2738 ;
  assign n2740 = \i_tv80_core_i_reg_RegsL_reg[5][1]/P0001  & n2739 ;
  assign n2749 = ~n2737 & ~n2740 ;
  assign n2753 = n2748 & n2749 ;
  assign n2754 = n2752 & n2753 ;
  assign n2755 = ~n2729 & ~n2754 ;
  assign n2760 = \i_tv80_core_i_reg_RegsL_reg[2][2]/P0001  & n2745 ;
  assign n2761 = \i_tv80_core_i_reg_RegsL_reg[7][2]/P0001  & n2731 ;
  assign n2766 = ~n2760 & ~n2761 ;
  assign n2762 = \i_tv80_core_i_reg_RegsL_reg[4][2]/P0001  & n2733 ;
  assign n2763 = \i_tv80_core_i_reg_RegsL_reg[3][2]/P0001  & n2743 ;
  assign n2767 = ~n2762 & ~n2763 ;
  assign n2768 = n2766 & n2767 ;
  assign n2756 = \i_tv80_core_i_reg_RegsL_reg[0][2]/P0001  & n2696 ;
  assign n2757 = \i_tv80_core_i_reg_RegsL_reg[5][2]/P0001  & n2739 ;
  assign n2764 = ~n2756 & ~n2757 ;
  assign n2758 = \i_tv80_core_i_reg_RegsL_reg[6][2]/P0001  & n2736 ;
  assign n2759 = \i_tv80_core_i_reg_RegsL_reg[1][2]/P0001  & n2741 ;
  assign n2765 = ~n2758 & ~n2759 ;
  assign n2769 = n2764 & n2765 ;
  assign n2770 = n2768 & n2769 ;
  assign n2771 = ~n2729 & ~n2770 ;
  assign n2772 = ~n2755 & ~n2771 ;
  assign n2773 = n2729 & n2770 ;
  assign n2778 = \i_tv80_core_i_reg_RegsL_reg[0][0]/P0001  & n2696 ;
  assign n2779 = \i_tv80_core_i_reg_RegsL_reg[1][0]/P0001  & n2741 ;
  assign n2784 = ~n2778 & ~n2779 ;
  assign n2780 = \i_tv80_core_i_reg_RegsL_reg[2][0]/P0001  & n2745 ;
  assign n2781 = \i_tv80_core_i_reg_RegsL_reg[3][0]/P0001  & n2743 ;
  assign n2785 = ~n2780 & ~n2781 ;
  assign n2786 = n2784 & n2785 ;
  assign n2774 = \i_tv80_core_i_reg_RegsL_reg[4][0]/P0001  & n2733 ;
  assign n2775 = \i_tv80_core_i_reg_RegsL_reg[5][0]/P0001  & n2739 ;
  assign n2782 = ~n2774 & ~n2775 ;
  assign n2776 = \i_tv80_core_i_reg_RegsL_reg[7][0]/P0001  & n2731 ;
  assign n2777 = \i_tv80_core_i_reg_RegsL_reg[6][0]/P0001  & n2736 ;
  assign n2783 = ~n2776 & ~n2777 ;
  assign n2787 = n2782 & n2783 ;
  assign n2788 = n2786 & n2787 ;
  assign n2789 = n2729 & n2754 ;
  assign n2790 = ~n2788 & ~n2789 ;
  assign n2791 = ~n2773 & n2790 ;
  assign n2792 = n2772 & ~n2791 ;
  assign n2797 = \i_tv80_core_i_reg_RegsL_reg[2][4]/NET0131  & n2745 ;
  assign n2798 = \i_tv80_core_i_reg_RegsL_reg[7][4]/NET0131  & n2731 ;
  assign n2803 = ~n2797 & ~n2798 ;
  assign n2799 = \i_tv80_core_i_reg_RegsL_reg[3][4]/NET0131  & n2743 ;
  assign n2800 = \i_tv80_core_i_reg_RegsL_reg[4][4]/NET0131  & n2733 ;
  assign n2804 = ~n2799 & ~n2800 ;
  assign n2805 = n2803 & n2804 ;
  assign n2793 = \i_tv80_core_i_reg_RegsL_reg[0][4]/NET0131  & n2696 ;
  assign n2794 = \i_tv80_core_i_reg_RegsL_reg[5][4]/NET0131  & n2739 ;
  assign n2801 = ~n2793 & ~n2794 ;
  assign n2795 = \i_tv80_core_i_reg_RegsL_reg[1][4]/NET0131  & n2741 ;
  assign n2796 = \i_tv80_core_i_reg_RegsL_reg[6][4]/NET0131  & n2736 ;
  assign n2802 = ~n2795 & ~n2796 ;
  assign n2806 = n2801 & n2802 ;
  assign n2807 = n2805 & n2806 ;
  assign n2808 = n2729 & n2807 ;
  assign n2813 = \i_tv80_core_i_reg_RegsL_reg[5][5]/NET0131  & n2739 ;
  assign n2814 = \i_tv80_core_i_reg_RegsL_reg[4][5]/NET0131  & n2733 ;
  assign n2819 = ~n2813 & ~n2814 ;
  assign n2815 = \i_tv80_core_i_reg_RegsL_reg[6][5]/NET0131  & n2736 ;
  assign n2816 = \i_tv80_core_i_reg_RegsL_reg[7][5]/NET0131  & n2731 ;
  assign n2820 = ~n2815 & ~n2816 ;
  assign n2821 = n2819 & n2820 ;
  assign n2809 = \i_tv80_core_i_reg_RegsL_reg[0][5]/NET0131  & n2696 ;
  assign n2810 = \i_tv80_core_i_reg_RegsL_reg[2][5]/NET0131  & n2745 ;
  assign n2817 = ~n2809 & ~n2810 ;
  assign n2811 = \i_tv80_core_i_reg_RegsL_reg[1][5]/NET0131  & n2741 ;
  assign n2812 = \i_tv80_core_i_reg_RegsL_reg[3][5]/NET0131  & n2743 ;
  assign n2818 = ~n2811 & ~n2812 ;
  assign n2822 = n2817 & n2818 ;
  assign n2823 = n2821 & n2822 ;
  assign n2824 = n2729 & n2823 ;
  assign n2825 = ~n2808 & ~n2824 ;
  assign n2830 = \i_tv80_core_i_reg_RegsL_reg[4][3]/NET0131  & n2733 ;
  assign n2831 = \i_tv80_core_i_reg_RegsL_reg[5][3]/NET0131  & n2739 ;
  assign n2836 = ~n2830 & ~n2831 ;
  assign n2832 = \i_tv80_core_i_reg_RegsL_reg[7][3]/NET0131  & n2731 ;
  assign n2833 = \i_tv80_core_i_reg_RegsL_reg[6][3]/NET0131  & n2736 ;
  assign n2837 = ~n2832 & ~n2833 ;
  assign n2838 = n2836 & n2837 ;
  assign n2826 = \i_tv80_core_i_reg_RegsL_reg[1][3]/NET0131  & n2741 ;
  assign n2827 = \i_tv80_core_i_reg_RegsL_reg[3][3]/NET0131  & n2743 ;
  assign n2834 = ~n2826 & ~n2827 ;
  assign n2828 = \i_tv80_core_i_reg_RegsL_reg[0][3]/NET0131  & n2696 ;
  assign n2829 = \i_tv80_core_i_reg_RegsL_reg[2][3]/NET0131  & n2745 ;
  assign n2835 = ~n2828 & ~n2829 ;
  assign n2839 = n2834 & n2835 ;
  assign n2840 = n2838 & n2839 ;
  assign n2841 = n2729 & n2840 ;
  assign n2846 = \i_tv80_core_i_reg_RegsL_reg[0][6]/NET0131  & n2696 ;
  assign n2847 = \i_tv80_core_i_reg_RegsL_reg[6][6]/NET0131  & n2736 ;
  assign n2852 = ~n2846 & ~n2847 ;
  assign n2848 = \i_tv80_core_i_reg_RegsL_reg[7][6]/NET0131  & n2731 ;
  assign n2849 = \i_tv80_core_i_reg_RegsL_reg[2][6]/NET0131  & n2745 ;
  assign n2853 = ~n2848 & ~n2849 ;
  assign n2854 = n2852 & n2853 ;
  assign n2842 = \i_tv80_core_i_reg_RegsL_reg[3][6]/NET0131  & n2743 ;
  assign n2843 = \i_tv80_core_i_reg_RegsL_reg[1][6]/NET0131  & n2741 ;
  assign n2850 = ~n2842 & ~n2843 ;
  assign n2844 = \i_tv80_core_i_reg_RegsL_reg[5][6]/NET0131  & n2739 ;
  assign n2845 = \i_tv80_core_i_reg_RegsL_reg[4][6]/NET0131  & n2733 ;
  assign n2851 = ~n2844 & ~n2845 ;
  assign n2855 = n2850 & n2851 ;
  assign n2856 = n2854 & n2855 ;
  assign n2857 = n2729 & n2856 ;
  assign n2858 = ~n2841 & ~n2857 ;
  assign n2859 = n2825 & n2858 ;
  assign n2860 = ~n2792 & n2859 ;
  assign n2861 = ~n2729 & ~n2807 ;
  assign n2862 = ~n2729 & ~n2840 ;
  assign n2863 = ~n2861 & ~n2862 ;
  assign n2864 = ~n2729 & ~n2823 ;
  assign n2865 = ~n2729 & ~n2856 ;
  assign n2866 = ~n2864 & ~n2865 ;
  assign n2867 = n2863 & n2866 ;
  assign n2868 = ~n2860 & n2867 ;
  assign n2873 = \i_tv80_core_i_reg_RegsL_reg[4][7]/NET0131  & n2733 ;
  assign n2874 = \i_tv80_core_i_reg_RegsL_reg[5][7]/NET0131  & n2739 ;
  assign n2879 = ~n2873 & ~n2874 ;
  assign n2875 = \i_tv80_core_i_reg_RegsL_reg[3][7]/NET0131  & n2743 ;
  assign n2876 = \i_tv80_core_i_reg_RegsL_reg[0][7]/NET0131  & n2696 ;
  assign n2880 = ~n2875 & ~n2876 ;
  assign n2881 = n2879 & n2880 ;
  assign n2869 = \i_tv80_core_i_reg_RegsL_reg[1][7]/NET0131  & n2741 ;
  assign n2870 = \i_tv80_core_i_reg_RegsL_reg[6][7]/NET0131  & n2736 ;
  assign n2877 = ~n2869 & ~n2870 ;
  assign n2871 = \i_tv80_core_i_reg_RegsL_reg[7][7]/NET0131  & n2731 ;
  assign n2872 = \i_tv80_core_i_reg_RegsL_reg[2][7]/NET0131  & n2745 ;
  assign n2878 = ~n2871 & ~n2872 ;
  assign n2882 = n2877 & n2878 ;
  assign n2883 = n2881 & n2882 ;
  assign n2884 = n2729 & n2883 ;
  assign n2885 = ~n2729 & ~n2883 ;
  assign n2886 = ~n2884 & ~n2885 ;
  assign n2887 = ~n2868 & n2886 ;
  assign n2888 = n2868 & ~n2886 ;
  assign n2889 = ~n2887 & ~n2888 ;
  assign n2890 = ~n2618 & n2698 ;
  assign n2891 = ~n2664 & n2890 ;
  assign n2892 = ~n2667 & n2891 ;
  assign n2893 = n2889 & n2892 ;
  assign n2894 = \i_tv80_core_RegBusA_r_reg[7]/P0001  & n2664 ;
  assign n2895 = ~n2664 & ~n2890 ;
  assign n2896 = ~n1841 & n2895 ;
  assign n2897 = ~n2894 & ~n2896 ;
  assign n2898 = ~n2667 & ~n2897 ;
  assign n2901 = \i_tv80_core_RegAddrB_r_reg[2]/P0001  & ~n2667 ;
  assign n2902 = \i_tv80_core_Alternate_reg/P0001  & n2667 ;
  assign n2903 = ~n2901 & ~n2902 ;
  assign n2899 = \i_tv80_core_RegAddrB_r_reg[1]/P0001  & ~n2667 ;
  assign n2906 = ~\i_tv80_core_RegAddrB_r_reg[0]/P0001  & ~n2667 ;
  assign n2913 = ~n2899 & ~n2906 ;
  assign n2916 = ~n2903 & n2913 ;
  assign n2917 = \i_tv80_core_i_reg_RegsL_reg[5][7]/NET0131  & n2916 ;
  assign n2910 = ~\i_tv80_core_RegAddrB_r_reg[1]/P0001  & n2906 ;
  assign n2918 = ~n2903 & n2910 ;
  assign n2919 = \i_tv80_core_i_reg_RegsL_reg[4][7]/NET0131  & n2918 ;
  assign n2926 = ~n2917 & ~n2919 ;
  assign n2907 = \i_tv80_core_RegAddrB_r_reg[1]/P0001  & n2906 ;
  assign n2920 = ~n2903 & n2907 ;
  assign n2921 = \i_tv80_core_i_reg_RegsL_reg[6][7]/NET0131  & n2920 ;
  assign n2900 = \i_tv80_core_RegAddrB_r_reg[0]/P0001  & n2899 ;
  assign n2922 = n2900 & n2903 ;
  assign n2923 = \i_tv80_core_i_reg_RegsL_reg[3][7]/NET0131  & n2922 ;
  assign n2927 = ~n2921 & ~n2923 ;
  assign n2928 = n2926 & n2927 ;
  assign n2904 = n2900 & ~n2903 ;
  assign n2905 = \i_tv80_core_i_reg_RegsL_reg[7][7]/NET0131  & n2904 ;
  assign n2908 = n2903 & n2907 ;
  assign n2909 = \i_tv80_core_i_reg_RegsL_reg[2][7]/NET0131  & n2908 ;
  assign n2924 = ~n2905 & ~n2909 ;
  assign n2911 = n2903 & n2910 ;
  assign n2912 = \i_tv80_core_i_reg_RegsL_reg[0][7]/NET0131  & n2911 ;
  assign n2914 = n2903 & n2913 ;
  assign n2915 = \i_tv80_core_i_reg_RegsL_reg[1][7]/NET0131  & n2914 ;
  assign n2925 = ~n2912 & ~n2915 ;
  assign n2929 = n2924 & n2925 ;
  assign n2930 = n2928 & n2929 ;
  assign n2931 = n2667 & ~n2930 ;
  assign n2932 = ~n2898 & ~n2931 ;
  assign n2933 = ~n2893 & n2932 ;
  assign n2934 = n2711 & ~n2933 ;
  assign n2935 = \i_tv80_core_i_reg_RegsL_reg[0][7]/NET0131  & ~n2711 ;
  assign n2936 = ~n2934 & ~n2935 ;
  assign n2937 = n2710 & n2741 ;
  assign n2938 = ~n2933 & n2937 ;
  assign n2939 = \i_tv80_core_i_reg_RegsL_reg[1][7]/NET0131  & ~n2937 ;
  assign n2940 = ~n2938 & ~n2939 ;
  assign n2941 = n2710 & n2745 ;
  assign n2942 = ~n2933 & n2941 ;
  assign n2943 = \i_tv80_core_i_reg_RegsL_reg[2][7]/NET0131  & ~n2941 ;
  assign n2944 = ~n2942 & ~n2943 ;
  assign n2945 = n2710 & n2743 ;
  assign n2946 = ~n2933 & n2945 ;
  assign n2947 = \i_tv80_core_i_reg_RegsL_reg[3][7]/NET0131  & ~n2945 ;
  assign n2948 = ~n2946 & ~n2947 ;
  assign n2949 = n2710 & n2733 ;
  assign n2950 = ~n2933 & n2949 ;
  assign n2951 = \i_tv80_core_i_reg_RegsL_reg[4][7]/NET0131  & ~n2949 ;
  assign n2952 = ~n2950 & ~n2951 ;
  assign n2953 = n2710 & n2739 ;
  assign n2954 = ~n2933 & n2953 ;
  assign n2955 = \i_tv80_core_i_reg_RegsL_reg[5][7]/NET0131  & ~n2953 ;
  assign n2956 = ~n2954 & ~n2955 ;
  assign n2957 = n2710 & n2736 ;
  assign n2958 = ~n2933 & n2957 ;
  assign n2959 = \i_tv80_core_i_reg_RegsL_reg[6][7]/NET0131  & ~n2957 ;
  assign n2960 = ~n2958 & ~n2959 ;
  assign n2961 = n2710 & n2731 ;
  assign n2962 = ~n2933 & n2961 ;
  assign n2963 = \i_tv80_core_i_reg_RegsL_reg[7][7]/NET0131  & ~n2961 ;
  assign n2964 = ~n2962 & ~n2963 ;
  assign n2966 = n2703 & n2704 ;
  assign n2967 = n1162 & n2966 ;
  assign n2968 = ~\i_tv80_core_Read_To_Reg_r_reg[0]/P0001  & n2967 ;
  assign n2969 = ~n1841 & n2968 ;
  assign n2971 = \i_tv80_core_ISet_reg[1]/P0001  & n1481 ;
  assign n2972 = ~\i_tv80_core_IR_reg[3]/P0001  & n2971 ;
  assign n2973 = n1034 & n2972 ;
  assign n2974 = \i_tv80_core_IR_reg[3]/P0001  & n1034 ;
  assign n2975 = n2971 & n2974 ;
  assign n2976 = ~\i_tv80_core_BusB_reg[7]/P0001  & ~n2975 ;
  assign n2977 = ~\i_tv80_core_BusB_reg[3]/P0001  & n2975 ;
  assign n2978 = ~n2976 & ~n2977 ;
  assign n2979 = ~n2973 & ~n2978 ;
  assign n2980 = ~\i_tv80_core_BusA_reg[3]/P0001  & n2973 ;
  assign n2981 = ~n2979 & ~n2980 ;
  assign n2982 = n1157 & ~n2981 ;
  assign n2970 = ~\do[7]_pad  & ~n1157 ;
  assign n2983 = ~n2968 & ~n2970 ;
  assign n2984 = ~n2982 & n2983 ;
  assign n2985 = ~\i_tv80_core_BusAck_reg/P0001  & ~n2984 ;
  assign n2986 = ~n2969 & n2985 ;
  assign n2965 = ~\do[7]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n2987 = reset_n_pad & ~n2965 ;
  assign n2988 = ~n2986 & n2987 ;
  assign n2990 = ~\i_tv80_core_Read_To_Reg_r_reg[1]/P0001  & ~\i_tv80_core_Read_To_Reg_r_reg[2]/P0001  ;
  assign n2991 = n1164 & n2990 ;
  assign n2992 = ~\i_tv80_core_Read_To_Reg_r_reg[0]/P0001  & n2991 ;
  assign n2994 = n382 & n675 ;
  assign n2995 = ~\i_tv80_core_IR_reg[2]/P0001  & n912 ;
  assign n2996 = n973 & n2995 ;
  assign n2997 = n2994 & n2996 ;
  assign n2998 = n2448 & n2997 ;
  assign n2999 = n860 & n2662 ;
  assign n3000 = ~n1635 & ~n2999 ;
  assign n3001 = n2699 & ~n3000 ;
  assign n3004 = \di_reg_reg[7]/P0001  & n1107 ;
  assign n3005 = ~n1107 & ~n2729 ;
  assign n3006 = ~n3004 & ~n3005 ;
  assign n3007 = n1107 & ~n2448 ;
  assign n3008 = \i_tv80_core_SP_reg[7]/P0001  & ~n1107 ;
  assign n3009 = ~n3007 & ~n3008 ;
  assign n3010 = ~n3006 & ~n3009 ;
  assign n3011 = n3006 & n3009 ;
  assign n3012 = ~n3010 & ~n3011 ;
  assign n3013 = \di_reg_reg[4]/P0001  & n1107 ;
  assign n3014 = ~n3005 & ~n3013 ;
  assign n3015 = n1107 & ~n2389 ;
  assign n3016 = \i_tv80_core_SP_reg[4]/P0001  & ~n1107 ;
  assign n3017 = ~n3015 & ~n3016 ;
  assign n3018 = ~n3014 & ~n3017 ;
  assign n3019 = n3014 & n3017 ;
  assign n3020 = \di_reg_reg[3]/P0001  & n1107 ;
  assign n3021 = ~n3005 & ~n3020 ;
  assign n3022 = n1107 & ~n2330 ;
  assign n3023 = \i_tv80_core_SP_reg[3]/P0001  & ~n1107 ;
  assign n3024 = ~n3022 & ~n3023 ;
  assign n3025 = n3021 & n3024 ;
  assign n3026 = \di_reg_reg[2]/P0001  & n1107 ;
  assign n3027 = ~n3005 & ~n3026 ;
  assign n3028 = n1107 & ~n1304 ;
  assign n3029 = \i_tv80_core_SP_reg[2]/P0001  & ~n1107 ;
  assign n3030 = ~n3028 & ~n3029 ;
  assign n3031 = ~n3027 & ~n3030 ;
  assign n3032 = n3027 & n3030 ;
  assign n3033 = \di_reg_reg[1]/P0001  & n1107 ;
  assign n3034 = ~n3005 & ~n3033 ;
  assign n3035 = n1107 & ~n1659 ;
  assign n3036 = \i_tv80_core_SP_reg[1]/P0001  & ~n1107 ;
  assign n3037 = ~n3035 & ~n3036 ;
  assign n3038 = n3034 & n3037 ;
  assign n3039 = \i_tv80_core_SP_reg[0]/P0001  & ~n1107 ;
  assign n3040 = \di_reg_reg[0]/P0001  & n1107 ;
  assign n3041 = ~n1883 & n3040 ;
  assign n3042 = ~n3039 & ~n3041 ;
  assign n3043 = ~n3038 & ~n3042 ;
  assign n3044 = ~n3034 & ~n3037 ;
  assign n3045 = ~n3043 & ~n3044 ;
  assign n3046 = ~n3032 & ~n3045 ;
  assign n3047 = ~n3031 & ~n3046 ;
  assign n3048 = ~n3025 & ~n3047 ;
  assign n3049 = ~n3021 & ~n3024 ;
  assign n3050 = ~n3048 & ~n3049 ;
  assign n3051 = ~n3019 & ~n3050 ;
  assign n3052 = ~n3018 & ~n3051 ;
  assign n3053 = \di_reg_reg[6]/P0001  & n1107 ;
  assign n3054 = ~n3005 & ~n3053 ;
  assign n3055 = n1107 & ~n1777 ;
  assign n3056 = \i_tv80_core_SP_reg[6]/P0001  & ~n1107 ;
  assign n3057 = ~n3055 & ~n3056 ;
  assign n3058 = n3054 & n3057 ;
  assign n3059 = \di_reg_reg[5]/P0001  & n1107 ;
  assign n3060 = ~n3005 & ~n3059 ;
  assign n3061 = n1107 & ~n1716 ;
  assign n3062 = \i_tv80_core_SP_reg[5]/P0001  & ~n1107 ;
  assign n3063 = ~n3061 & ~n3062 ;
  assign n3064 = n3060 & n3063 ;
  assign n3065 = ~n3058 & ~n3064 ;
  assign n3066 = ~n3052 & n3065 ;
  assign n3067 = ~n3060 & ~n3063 ;
  assign n3068 = ~n3054 & ~n3057 ;
  assign n3069 = ~n3067 & ~n3068 ;
  assign n3070 = ~n3058 & ~n3069 ;
  assign n3071 = ~n3066 & ~n3070 ;
  assign n3072 = n3012 & ~n3071 ;
  assign n3073 = ~n3012 & n3071 ;
  assign n3074 = ~n3072 & ~n3073 ;
  assign n3075 = n3001 & n3074 ;
  assign n3002 = ~n2646 & n3001 ;
  assign n3003 = \i_tv80_core_SP_reg[7]/P0001  & ~n3002 ;
  assign n3076 = ~n2997 & ~n3003 ;
  assign n3077 = ~n3075 & n3076 ;
  assign n3078 = ~n2998 & ~n3077 ;
  assign n3079 = ~n1113 & ~n3078 ;
  assign n3080 = ~\i_tv80_core_SP_reg[7]/P0001  & n1113 ;
  assign n3081 = ~n3079 & ~n3080 ;
  assign n3082 = ~n2992 & ~n3081 ;
  assign n2993 = n1841 & n2992 ;
  assign n3083 = ~\i_tv80_core_BusAck_reg/P0001  & ~n2993 ;
  assign n3084 = ~n3082 & n3083 ;
  assign n2989 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[7]/P0001  ;
  assign n3085 = reset_n_pad & ~n2989 ;
  assign n3086 = ~n3084 & n3085 ;
  assign n3109 = ~n544 & ~n595 ;
  assign n3111 = ~\i_tv80_core_ALU_Op_r_reg[1]/P0001  & ~\i_tv80_core_ALU_Op_r_reg[2]/NET0131  ;
  assign n3112 = ~n3109 & ~n3111 ;
  assign n3110 = ~n696 & n3109 ;
  assign n3113 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n3110 ;
  assign n3114 = ~n3112 & n3113 ;
  assign n3118 = ~\i_tv80_core_PreserveC_r_reg/P0001  & ~n386 ;
  assign n3117 = n735 & ~n757 ;
  assign n3115 = ~n627 & ~n649 ;
  assign n3116 = n604 & ~n3115 ;
  assign n3119 = \i_tv80_core_F_reg[0]/P0001  & n699 ;
  assign n3120 = ~n3116 & ~n3119 ;
  assign n3121 = ~n3117 & n3120 ;
  assign n3122 = n3118 & n3121 ;
  assign n3123 = ~n3114 & n3122 ;
  assign n3126 = n382 & n1380 ;
  assign n3127 = n1103 & n3126 ;
  assign n3129 = \i_tv80_core_F_reg[0]/P0001  & ~n3127 ;
  assign n3128 = ~n621 & n3127 ;
  assign n3130 = ~n1117 & ~n3128 ;
  assign n3131 = ~n3129 & n3130 ;
  assign n3125 = ~\i_tv80_core_Fp_reg[0]/P0001  & n1117 ;
  assign n3132 = ~n1113 & ~n3125 ;
  assign n3133 = ~n3131 & n3132 ;
  assign n3124 = \i_tv80_core_F_reg[0]/P0001  & n1113 ;
  assign n3134 = ~n3118 & ~n3124 ;
  assign n3135 = ~n3133 & n3134 ;
  assign n3136 = ~n3123 & ~n3135 ;
  assign n3137 = ~n1167 & ~n3136 ;
  assign n3095 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n514 ;
  assign n3089 = \i_tv80_core_BusA_reg[0]/P0001  & n735 ;
  assign n3098 = \i_tv80_core_Save_ALU_r_reg/P0001  & ~n3089 ;
  assign n3090 = n700 & ~n703 ;
  assign n3097 = n370 & n685 ;
  assign n3099 = ~n3090 & ~n3097 ;
  assign n3100 = n3098 & n3099 ;
  assign n3092 = \i_tv80_core_ALU_Op_r_reg[0]/P0001  & n684 ;
  assign n3091 = ~\i_tv80_core_BusB_reg[0]/P0001  & ~n684 ;
  assign n3093 = n1175 & ~n3091 ;
  assign n3094 = ~n3092 & n3093 ;
  assign n3096 = n604 & ~n652 ;
  assign n3101 = ~n3094 & ~n3096 ;
  assign n3102 = n3100 & n3101 ;
  assign n3103 = ~n3095 & n3102 ;
  assign n3088 = ~\di_reg_reg[0]/P0001  & ~\i_tv80_core_Save_ALU_r_reg/P0001  ;
  assign n3104 = ~n1172 & ~n3088 ;
  assign n3105 = ~n3103 & n3104 ;
  assign n3106 = \i_tv80_core_BusB_reg[0]/P0001  & n1172 ;
  assign n3107 = ~n3105 & ~n3106 ;
  assign n3108 = n1167 & n3107 ;
  assign n3138 = ~\i_tv80_core_BusAck_reg/P0001  & ~n3108 ;
  assign n3139 = ~n3137 & n3138 ;
  assign n3087 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_F_reg[0]/P0001  ;
  assign n3140 = reset_n_pad & ~n3087 ;
  assign n3141 = ~n3139 & n3140 ;
  assign n3151 = \i_tv80_core_Ap_reg[7]/P0001  & n1117 ;
  assign n3152 = n382 & n912 ;
  assign n3153 = n1382 & n3152 ;
  assign n3154 = n1103 & n3153 ;
  assign n3155 = ~n1117 & n3154 ;
  assign n3156 = ~\i_tv80_core_ACC_reg[7]/P0001  & n3155 ;
  assign n3157 = ~n3151 & ~n3156 ;
  assign n3158 = ~n1113 & ~n3157 ;
  assign n3159 = ~n1113 & n3154 ;
  assign n3160 = ~n1118 & ~n3159 ;
  assign n3161 = \i_tv80_core_ACC_reg[7]/P0001  & n3160 ;
  assign n3162 = ~n3158 & ~n3161 ;
  assign n3163 = ~n1112 & ~n3162 ;
  assign n3143 = \i_tv80_core_Read_To_Reg_r_reg[0]/P0001  & n2967 ;
  assign n3145 = n678 & n1110 ;
  assign n3146 = \i_tv80_core_R_reg[7]/P0001  & n3145 ;
  assign n3147 = ~n645 & n1110 ;
  assign n3148 = \i_tv80_core_I_reg[7]/P0001  & ~n3147 ;
  assign n3149 = ~n3146 & ~n3148 ;
  assign n3150 = n1111 & ~n3149 ;
  assign n3164 = ~n3143 & ~n3150 ;
  assign n3165 = ~n3163 & n3164 ;
  assign n3144 = n1841 & n3143 ;
  assign n3166 = ~\i_tv80_core_BusAck_reg/P0001  & ~n3144 ;
  assign n3167 = ~n3165 & n3166 ;
  assign n3142 = \i_tv80_core_ACC_reg[7]/P0001  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n3168 = reset_n_pad & ~n3142 ;
  assign n3169 = ~n3167 & n3168 ;
  assign n3170 = ~n2646 & n2699 ;
  assign n3171 = \i_tv80_core_SP_reg[15]/P0001  & ~n3170 ;
  assign n3172 = n1107 & ~n2268 ;
  assign n3173 = \i_tv80_core_SP_reg[15]/P0001  & ~n1107 ;
  assign n3174 = ~n3172 & ~n3173 ;
  assign n3175 = n3006 & ~n3174 ;
  assign n3176 = ~n3006 & n3174 ;
  assign n3177 = ~n3175 & ~n3176 ;
  assign n3178 = n1107 & ~n2142 ;
  assign n3179 = \i_tv80_core_SP_reg[13]/P0001  & ~n1107 ;
  assign n3180 = ~n3178 & ~n3179 ;
  assign n3181 = n3006 & n3180 ;
  assign n3182 = n1107 & ~n2205 ;
  assign n3183 = \i_tv80_core_SP_reg[14]/P0001  & ~n1107 ;
  assign n3184 = ~n3182 & ~n3183 ;
  assign n3185 = n3006 & n3184 ;
  assign n3186 = ~n3181 & ~n3185 ;
  assign n3187 = n1107 & ~n2509 ;
  assign n3188 = \i_tv80_core_SP_reg[8]/P0001  & ~n1107 ;
  assign n3189 = ~n3187 & ~n3188 ;
  assign n3190 = n3006 & n3189 ;
  assign n3191 = ~n3011 & ~n3190 ;
  assign n3192 = ~n3071 & n3191 ;
  assign n3193 = ~n3006 & ~n3189 ;
  assign n3194 = ~n3010 & ~n3193 ;
  assign n3195 = ~n3192 & n3194 ;
  assign n3196 = n1107 & ~n1945 ;
  assign n3197 = \i_tv80_core_SP_reg[10]/P0001  & ~n1107 ;
  assign n3198 = ~n3196 & ~n3197 ;
  assign n3199 = n3006 & n3198 ;
  assign n3200 = n1107 & ~n2571 ;
  assign n3201 = \i_tv80_core_SP_reg[9]/P0001  & ~n1107 ;
  assign n3202 = ~n3200 & ~n3201 ;
  assign n3203 = n3006 & n3202 ;
  assign n3204 = ~n3199 & ~n3203 ;
  assign n3205 = ~n3195 & n3204 ;
  assign n3206 = ~n3006 & ~n3202 ;
  assign n3207 = ~n3006 & ~n3198 ;
  assign n3208 = ~n3206 & ~n3207 ;
  assign n3209 = ~n3205 & n3208 ;
  assign n3210 = n1107 & ~n2016 ;
  assign n3211 = \i_tv80_core_SP_reg[11]/P0001  & ~n1107 ;
  assign n3212 = ~n3210 & ~n3211 ;
  assign n3213 = n3006 & n3212 ;
  assign n3214 = n1107 & ~n2079 ;
  assign n3215 = \i_tv80_core_SP_reg[12]/P0001  & ~n1107 ;
  assign n3216 = ~n3214 & ~n3215 ;
  assign n3217 = n3006 & n3216 ;
  assign n3218 = ~n3213 & ~n3217 ;
  assign n3219 = ~n3209 & n3218 ;
  assign n3220 = n3186 & n3219 ;
  assign n3222 = ~n3006 & ~n3212 ;
  assign n3223 = ~n3006 & ~n3216 ;
  assign n3224 = ~n3222 & ~n3223 ;
  assign n3225 = n3186 & ~n3224 ;
  assign n3221 = ~n3006 & ~n3180 ;
  assign n3226 = ~n3006 & ~n3184 ;
  assign n3227 = ~n3221 & ~n3226 ;
  assign n3228 = ~n3225 & n3227 ;
  assign n3229 = ~n3220 & n3228 ;
  assign n3230 = n3177 & n3229 ;
  assign n3231 = ~n3177 & ~n3229 ;
  assign n3232 = ~n3230 & ~n3231 ;
  assign n3233 = n2699 & n3232 ;
  assign n3234 = ~n3171 & ~n3233 ;
  assign n3235 = ~n3000 & ~n3234 ;
  assign n3236 = \i_tv80_core_SP_reg[15]/P0001  & n3000 ;
  assign n3237 = ~n2997 & ~n3236 ;
  assign n3238 = ~n3235 & n3237 ;
  assign n3239 = n2268 & n2997 ;
  assign n3240 = ~n1113 & ~n3239 ;
  assign n3241 = ~n3238 & n3240 ;
  assign n3242 = \i_tv80_core_Read_To_Reg_r_reg[0]/P0001  & n2991 ;
  assign n3243 = \i_tv80_core_SP_reg[15]/P0001  & n1113 ;
  assign n3244 = ~n3242 & ~n3243 ;
  assign n3245 = ~n3241 & n3244 ;
  assign n3246 = n1841 & n3242 ;
  assign n3247 = ~\i_tv80_core_BusAck_reg/P0001  & ~n3246 ;
  assign n3248 = ~n3245 & n3247 ;
  assign n3249 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[15]/P0001  ;
  assign n3250 = reset_n_pad & ~n3249 ;
  assign n3251 = ~n3248 & n3250 ;
  assign n3256 = \i_tv80_core_i_reg_RegsH_reg[6][2]/P0001  & n2736 ;
  assign n3257 = \i_tv80_core_i_reg_RegsH_reg[0][2]/P0001  & n2696 ;
  assign n3262 = ~n3256 & ~n3257 ;
  assign n3258 = \i_tv80_core_i_reg_RegsH_reg[3][2]/P0001  & n2743 ;
  assign n3259 = \i_tv80_core_i_reg_RegsH_reg[7][2]/P0001  & n2731 ;
  assign n3263 = ~n3258 & ~n3259 ;
  assign n3264 = n3262 & n3263 ;
  assign n3252 = \i_tv80_core_i_reg_RegsH_reg[5][2]/P0001  & n2739 ;
  assign n3253 = \i_tv80_core_i_reg_RegsH_reg[2][2]/P0001  & n2745 ;
  assign n3260 = ~n3252 & ~n3253 ;
  assign n3254 = \i_tv80_core_i_reg_RegsH_reg[1][2]/P0001  & n2741 ;
  assign n3255 = \i_tv80_core_i_reg_RegsH_reg[4][2]/P0001  & n2733 ;
  assign n3261 = ~n3254 & ~n3255 ;
  assign n3265 = n3260 & n3261 ;
  assign n3266 = n3264 & n3265 ;
  assign n3267 = n2729 & n3266 ;
  assign n3272 = \i_tv80_core_i_reg_RegsH_reg[5][1]/P0001  & n2739 ;
  assign n3273 = \i_tv80_core_i_reg_RegsH_reg[1][1]/P0001  & n2741 ;
  assign n3278 = ~n3272 & ~n3273 ;
  assign n3274 = \i_tv80_core_i_reg_RegsH_reg[0][1]/P0001  & n2696 ;
  assign n3275 = \i_tv80_core_i_reg_RegsH_reg[2][1]/P0001  & n2745 ;
  assign n3279 = ~n3274 & ~n3275 ;
  assign n3280 = n3278 & n3279 ;
  assign n3268 = \i_tv80_core_i_reg_RegsH_reg[6][1]/P0001  & n2736 ;
  assign n3269 = \i_tv80_core_i_reg_RegsH_reg[7][1]/P0001  & n2731 ;
  assign n3276 = ~n3268 & ~n3269 ;
  assign n3270 = \i_tv80_core_i_reg_RegsH_reg[4][1]/P0001  & n2733 ;
  assign n3271 = \i_tv80_core_i_reg_RegsH_reg[3][1]/P0001  & n2743 ;
  assign n3277 = ~n3270 & ~n3271 ;
  assign n3281 = n3276 & n3277 ;
  assign n3282 = n3280 & n3281 ;
  assign n3283 = n2729 & n3282 ;
  assign n3284 = ~n3267 & ~n3283 ;
  assign n3289 = \i_tv80_core_i_reg_RegsH_reg[6][0]/P0001  & n2736 ;
  assign n3290 = \i_tv80_core_i_reg_RegsH_reg[2][0]/P0001  & n2745 ;
  assign n3295 = ~n3289 & ~n3290 ;
  assign n3291 = \i_tv80_core_i_reg_RegsH_reg[1][0]/P0001  & n2741 ;
  assign n3292 = \i_tv80_core_i_reg_RegsH_reg[7][0]/P0001  & n2731 ;
  assign n3296 = ~n3291 & ~n3292 ;
  assign n3297 = n3295 & n3296 ;
  assign n3285 = \i_tv80_core_i_reg_RegsH_reg[4][0]/P0001  & n2733 ;
  assign n3286 = \i_tv80_core_i_reg_RegsH_reg[3][0]/P0001  & n2743 ;
  assign n3293 = ~n3285 & ~n3286 ;
  assign n3287 = \i_tv80_core_i_reg_RegsH_reg[5][0]/P0001  & n2739 ;
  assign n3288 = \i_tv80_core_i_reg_RegsH_reg[0][0]/P0001  & n2696 ;
  assign n3294 = ~n3287 & ~n3288 ;
  assign n3298 = n3293 & n3294 ;
  assign n3299 = n3297 & n3298 ;
  assign n3300 = n2729 & n3299 ;
  assign n3301 = n3284 & ~n3300 ;
  assign n3302 = ~n2884 & n3301 ;
  assign n3303 = ~n2868 & n3302 ;
  assign n3304 = ~n2729 & ~n3299 ;
  assign n3305 = ~n2885 & ~n3304 ;
  assign n3306 = ~n2729 & ~n3266 ;
  assign n3307 = ~n2729 & ~n3282 ;
  assign n3308 = ~n3306 & ~n3307 ;
  assign n3309 = n3305 & n3308 ;
  assign n3310 = ~n3303 & n3309 ;
  assign n3315 = \i_tv80_core_i_reg_RegsH_reg[3][6]/P0001  & n2743 ;
  assign n3316 = \i_tv80_core_i_reg_RegsH_reg[2][6]/P0001  & n2745 ;
  assign n3321 = ~n3315 & ~n3316 ;
  assign n3317 = \i_tv80_core_i_reg_RegsH_reg[7][6]/P0001  & n2731 ;
  assign n3318 = \i_tv80_core_i_reg_RegsH_reg[1][6]/P0001  & n2741 ;
  assign n3322 = ~n3317 & ~n3318 ;
  assign n3323 = n3321 & n3322 ;
  assign n3311 = \i_tv80_core_i_reg_RegsH_reg[4][6]/P0001  & n2733 ;
  assign n3312 = \i_tv80_core_i_reg_RegsH_reg[6][6]/P0001  & n2736 ;
  assign n3319 = ~n3311 & ~n3312 ;
  assign n3313 = \i_tv80_core_i_reg_RegsH_reg[5][6]/P0001  & n2739 ;
  assign n3314 = \i_tv80_core_i_reg_RegsH_reg[0][6]/P0001  & n2696 ;
  assign n3320 = ~n3313 & ~n3314 ;
  assign n3324 = n3319 & n3320 ;
  assign n3325 = n3323 & n3324 ;
  assign n3326 = n2729 & n3325 ;
  assign n3331 = \i_tv80_core_i_reg_RegsH_reg[2][3]/P0001  & n2745 ;
  assign n3332 = \i_tv80_core_i_reg_RegsH_reg[3][3]/P0001  & n2743 ;
  assign n3337 = ~n3331 & ~n3332 ;
  assign n3333 = \i_tv80_core_i_reg_RegsH_reg[0][3]/P0001  & n2696 ;
  assign n3334 = \i_tv80_core_i_reg_RegsH_reg[4][3]/P0001  & n2733 ;
  assign n3338 = ~n3333 & ~n3334 ;
  assign n3339 = n3337 & n3338 ;
  assign n3327 = \i_tv80_core_i_reg_RegsH_reg[1][3]/P0001  & n2741 ;
  assign n3328 = \i_tv80_core_i_reg_RegsH_reg[7][3]/P0001  & n2731 ;
  assign n3335 = ~n3327 & ~n3328 ;
  assign n3329 = \i_tv80_core_i_reg_RegsH_reg[5][3]/P0001  & n2739 ;
  assign n3330 = \i_tv80_core_i_reg_RegsH_reg[6][3]/P0001  & n2736 ;
  assign n3336 = ~n3329 & ~n3330 ;
  assign n3340 = n3335 & n3336 ;
  assign n3341 = n3339 & n3340 ;
  assign n3342 = n2729 & n3341 ;
  assign n3347 = \i_tv80_core_i_reg_RegsH_reg[0][4]/P0001  & n2696 ;
  assign n3348 = \i_tv80_core_i_reg_RegsH_reg[5][4]/P0001  & n2739 ;
  assign n3353 = ~n3347 & ~n3348 ;
  assign n3349 = \i_tv80_core_i_reg_RegsH_reg[6][4]/P0001  & n2736 ;
  assign n3350 = \i_tv80_core_i_reg_RegsH_reg[2][4]/P0001  & n2745 ;
  assign n3354 = ~n3349 & ~n3350 ;
  assign n3355 = n3353 & n3354 ;
  assign n3343 = \i_tv80_core_i_reg_RegsH_reg[1][4]/P0001  & n2741 ;
  assign n3344 = \i_tv80_core_i_reg_RegsH_reg[3][4]/P0001  & n2743 ;
  assign n3351 = ~n3343 & ~n3344 ;
  assign n3345 = \i_tv80_core_i_reg_RegsH_reg[7][4]/P0001  & n2731 ;
  assign n3346 = \i_tv80_core_i_reg_RegsH_reg[4][4]/P0001  & n2733 ;
  assign n3352 = ~n3345 & ~n3346 ;
  assign n3356 = n3351 & n3352 ;
  assign n3357 = n3355 & n3356 ;
  assign n3358 = n2729 & n3357 ;
  assign n3359 = ~n3342 & ~n3358 ;
  assign n3364 = \i_tv80_core_i_reg_RegsH_reg[6][5]/P0001  & n2736 ;
  assign n3365 = \i_tv80_core_i_reg_RegsH_reg[3][5]/P0001  & n2743 ;
  assign n3370 = ~n3364 & ~n3365 ;
  assign n3366 = \i_tv80_core_i_reg_RegsH_reg[5][5]/P0001  & n2739 ;
  assign n3367 = \i_tv80_core_i_reg_RegsH_reg[4][5]/P0001  & n2733 ;
  assign n3371 = ~n3366 & ~n3367 ;
  assign n3372 = n3370 & n3371 ;
  assign n3360 = \i_tv80_core_i_reg_RegsH_reg[2][5]/P0001  & n2745 ;
  assign n3361 = \i_tv80_core_i_reg_RegsH_reg[7][5]/P0001  & n2731 ;
  assign n3368 = ~n3360 & ~n3361 ;
  assign n3362 = \i_tv80_core_i_reg_RegsH_reg[0][5]/P0001  & n2696 ;
  assign n3363 = \i_tv80_core_i_reg_RegsH_reg[1][5]/P0001  & n2741 ;
  assign n3369 = ~n3362 & ~n3363 ;
  assign n3373 = n3368 & n3369 ;
  assign n3374 = n3372 & n3373 ;
  assign n3375 = n2729 & n3374 ;
  assign n3376 = n3359 & ~n3375 ;
  assign n3377 = ~n3326 & n3376 ;
  assign n3378 = ~n3310 & n3377 ;
  assign n3379 = ~n2729 & ~n3325 ;
  assign n3380 = ~n2729 & ~n3341 ;
  assign n3381 = ~n2729 & ~n3357 ;
  assign n3382 = ~n3380 & ~n3381 ;
  assign n3383 = ~n2729 & ~n3374 ;
  assign n3384 = n3382 & ~n3383 ;
  assign n3385 = ~n3379 & n3384 ;
  assign n3386 = ~n3378 & n3385 ;
  assign n3391 = \i_tv80_core_i_reg_RegsH_reg[2][7]/P0002  & n2745 ;
  assign n3392 = \i_tv80_core_i_reg_RegsH_reg[3][7]/P0002  & n2743 ;
  assign n3397 = ~n3391 & ~n3392 ;
  assign n3393 = \i_tv80_core_i_reg_RegsH_reg[7][7]/P0002  & n2731 ;
  assign n3394 = \i_tv80_core_i_reg_RegsH_reg[6][7]/P0002  & n2736 ;
  assign n3398 = ~n3393 & ~n3394 ;
  assign n3399 = n3397 & n3398 ;
  assign n3387 = \i_tv80_core_i_reg_RegsH_reg[4][7]/P0002  & n2733 ;
  assign n3388 = \i_tv80_core_i_reg_RegsH_reg[5][7]/P0002  & n2739 ;
  assign n3395 = ~n3387 & ~n3388 ;
  assign n3389 = \i_tv80_core_i_reg_RegsH_reg[0][7]/P0002  & n2696 ;
  assign n3390 = \i_tv80_core_i_reg_RegsH_reg[1][7]/P0002  & n2741 ;
  assign n3396 = ~n3389 & ~n3390 ;
  assign n3400 = n3395 & n3396 ;
  assign n3401 = n3399 & n3400 ;
  assign n3402 = n2729 & ~n3401 ;
  assign n3403 = ~n2729 & n3401 ;
  assign n3404 = ~n3402 & ~n3403 ;
  assign n3405 = n3386 & n3404 ;
  assign n3406 = ~n3386 & ~n3404 ;
  assign n3407 = ~n3405 & ~n3406 ;
  assign n3408 = n2891 & n3407 ;
  assign n3409 = \i_tv80_core_RegBusA_r_reg[15]/P0001  & n2664 ;
  assign n3410 = ~n2896 & ~n3409 ;
  assign n3411 = ~n2667 & n3410 ;
  assign n3412 = ~n3408 & n3411 ;
  assign n3417 = \i_tv80_core_i_reg_RegsH_reg[7][7]/P0002  & n2904 ;
  assign n3418 = \i_tv80_core_i_reg_RegsH_reg[6][7]/P0002  & n2920 ;
  assign n3423 = ~n3417 & ~n3418 ;
  assign n3419 = \i_tv80_core_i_reg_RegsH_reg[5][7]/P0002  & n2916 ;
  assign n3420 = \i_tv80_core_i_reg_RegsH_reg[1][7]/P0002  & n2914 ;
  assign n3424 = ~n3419 & ~n3420 ;
  assign n3425 = n3423 & n3424 ;
  assign n3413 = \i_tv80_core_i_reg_RegsH_reg[4][7]/P0002  & n2918 ;
  assign n3414 = \i_tv80_core_i_reg_RegsH_reg[0][7]/P0002  & n2911 ;
  assign n3421 = ~n3413 & ~n3414 ;
  assign n3415 = \i_tv80_core_i_reg_RegsH_reg[2][7]/P0002  & n2908 ;
  assign n3416 = \i_tv80_core_i_reg_RegsH_reg[3][7]/P0002  & n2922 ;
  assign n3422 = ~n3415 & ~n3416 ;
  assign n3426 = n3421 & n3422 ;
  assign n3427 = n3425 & n3426 ;
  assign n3428 = n2667 & n3427 ;
  assign n3429 = ~n3412 & ~n3428 ;
  assign n3430 = n2696 & ~n3429 ;
  assign n3431 = ~\i_tv80_core_i_reg_RegsH_reg[0][7]/P0002  & ~n2696 ;
  assign n3432 = ~n3430 & ~n3431 ;
  assign n3433 = n2741 & ~n3429 ;
  assign n3434 = ~\i_tv80_core_i_reg_RegsH_reg[1][7]/P0002  & ~n2741 ;
  assign n3435 = ~n3433 & ~n3434 ;
  assign n3436 = n2745 & ~n3429 ;
  assign n3437 = ~\i_tv80_core_i_reg_RegsH_reg[2][7]/P0002  & ~n2745 ;
  assign n3438 = ~n3436 & ~n3437 ;
  assign n3439 = n2743 & ~n3429 ;
  assign n3440 = ~\i_tv80_core_i_reg_RegsH_reg[3][7]/P0002  & ~n2743 ;
  assign n3441 = ~n3439 & ~n3440 ;
  assign n3442 = n2733 & ~n3429 ;
  assign n3443 = ~\i_tv80_core_i_reg_RegsH_reg[4][7]/P0002  & ~n2733 ;
  assign n3444 = ~n3442 & ~n3443 ;
  assign n3445 = n2739 & ~n3429 ;
  assign n3446 = ~\i_tv80_core_i_reg_RegsH_reg[5][7]/P0002  & ~n2739 ;
  assign n3447 = ~n3445 & ~n3446 ;
  assign n3448 = n2736 & ~n3429 ;
  assign n3449 = ~\i_tv80_core_i_reg_RegsH_reg[6][7]/P0002  & ~n2736 ;
  assign n3450 = ~n3448 & ~n3449 ;
  assign n3451 = ~\i_tv80_core_Read_To_Reg_r_reg[0]/P0001  & n2705 ;
  assign n3452 = n1162 & n3451 ;
  assign n3453 = n2686 & ~n3452 ;
  assign n3454 = ~n2702 & n3453 ;
  assign n3455 = ~\i_tv80_core_BusAck_reg/P0001  & ~n3454 ;
  assign n3456 = n2696 & n3455 ;
  assign n3457 = ~n3326 & ~n3379 ;
  assign n3458 = ~n2861 & ~n2864 ;
  assign n3459 = ~n2755 & ~n2790 ;
  assign n3460 = ~n2773 & ~n2841 ;
  assign n3461 = ~n3459 & n3460 ;
  assign n3462 = ~n2771 & ~n2862 ;
  assign n3463 = ~n3461 & n3462 ;
  assign n3464 = n2825 & ~n3463 ;
  assign n3465 = n3458 & ~n3464 ;
  assign n3466 = ~n2857 & ~n2884 ;
  assign n3467 = ~n3300 & n3466 ;
  assign n3468 = ~n3283 & n3467 ;
  assign n3469 = ~n3465 & n3468 ;
  assign n3470 = ~n2865 & ~n2885 ;
  assign n3471 = ~n3304 & ~n3307 ;
  assign n3472 = n3470 & n3471 ;
  assign n3473 = ~n3469 & n3472 ;
  assign n3474 = ~n3267 & n3376 ;
  assign n3475 = ~n3473 & n3474 ;
  assign n3476 = ~n3306 & n3384 ;
  assign n3477 = ~n3475 & n3476 ;
  assign n3478 = n3457 & ~n3477 ;
  assign n3479 = ~n3457 & n3477 ;
  assign n3480 = ~n3478 & ~n3479 ;
  assign n3481 = n2891 & n3480 ;
  assign n3486 = \i_tv80_core_i_reg_RegsH_reg[4][6]/P0001  & n2918 ;
  assign n3487 = \i_tv80_core_i_reg_RegsH_reg[5][6]/P0001  & n2916 ;
  assign n3492 = ~n3486 & ~n3487 ;
  assign n3488 = \i_tv80_core_i_reg_RegsH_reg[3][6]/P0001  & n2922 ;
  assign n3489 = \i_tv80_core_i_reg_RegsH_reg[0][6]/P0001  & n2911 ;
  assign n3493 = ~n3488 & ~n3489 ;
  assign n3494 = n3492 & n3493 ;
  assign n3482 = \i_tv80_core_i_reg_RegsH_reg[2][6]/P0001  & n2908 ;
  assign n3483 = \i_tv80_core_i_reg_RegsH_reg[1][6]/P0001  & n2914 ;
  assign n3490 = ~n3482 & ~n3483 ;
  assign n3484 = \i_tv80_core_i_reg_RegsH_reg[7][6]/P0001  & n2904 ;
  assign n3485 = \i_tv80_core_i_reg_RegsH_reg[6][6]/P0001  & n2920 ;
  assign n3491 = ~n3484 & ~n3485 ;
  assign n3495 = n3490 & n3491 ;
  assign n3496 = n3494 & n3495 ;
  assign n3497 = n2667 & ~n3496 ;
  assign n3498 = ~n1220 & n2895 ;
  assign n3499 = \i_tv80_core_RegBusA_r_reg[14]/P0001  & n2664 ;
  assign n3500 = ~n3498 & ~n3499 ;
  assign n3501 = ~n2667 & ~n3500 ;
  assign n3502 = ~n3497 & ~n3501 ;
  assign n3503 = ~n3481 & n3502 ;
  assign n3504 = n3456 & ~n3503 ;
  assign n3505 = \i_tv80_core_i_reg_RegsH_reg[0][6]/P0001  & ~n3456 ;
  assign n3506 = ~n3504 & ~n3505 ;
  assign n3507 = n2743 & n3455 ;
  assign n3508 = ~n3503 & n3507 ;
  assign n3509 = \i_tv80_core_i_reg_RegsH_reg[3][6]/P0001  & ~n3507 ;
  assign n3510 = ~n3508 & ~n3509 ;
  assign n3511 = n2733 & n3455 ;
  assign n3512 = ~n3503 & n3511 ;
  assign n3513 = \i_tv80_core_i_reg_RegsH_reg[4][6]/P0001  & ~n3511 ;
  assign n3514 = ~n3512 & ~n3513 ;
  assign n3515 = n2731 & n3455 ;
  assign n3516 = ~n3503 & n3515 ;
  assign n3517 = \i_tv80_core_i_reg_RegsH_reg[7][6]/P0001  & ~n3515 ;
  assign n3518 = ~n3516 & ~n3517 ;
  assign n3519 = \i_tv80_core_i_reg_RegsL_reg[0][6]/NET0131  & ~n2711 ;
  assign n3520 = ~n2857 & ~n2865 ;
  assign n3521 = ~n3465 & n3520 ;
  assign n3522 = n3465 & ~n3520 ;
  assign n3523 = ~n3521 & ~n3522 ;
  assign n3524 = n2891 & n3523 ;
  assign n3525 = \i_tv80_core_RegBusA_r_reg[6]/P0001  & n2664 ;
  assign n3526 = ~n3498 & ~n3525 ;
  assign n3527 = ~n3524 & n3526 ;
  assign n3528 = ~n2667 & ~n3527 ;
  assign n3533 = \i_tv80_core_i_reg_RegsL_reg[7][6]/NET0131  & n2904 ;
  assign n3534 = \i_tv80_core_i_reg_RegsL_reg[6][6]/NET0131  & n2920 ;
  assign n3539 = ~n3533 & ~n3534 ;
  assign n3535 = \i_tv80_core_i_reg_RegsL_reg[1][6]/NET0131  & n2914 ;
  assign n3536 = \i_tv80_core_i_reg_RegsL_reg[2][6]/NET0131  & n2908 ;
  assign n3540 = ~n3535 & ~n3536 ;
  assign n3541 = n3539 & n3540 ;
  assign n3529 = \i_tv80_core_i_reg_RegsL_reg[0][6]/NET0131  & n2911 ;
  assign n3530 = \i_tv80_core_i_reg_RegsL_reg[3][6]/NET0131  & n2922 ;
  assign n3537 = ~n3529 & ~n3530 ;
  assign n3531 = \i_tv80_core_i_reg_RegsL_reg[4][6]/NET0131  & n2918 ;
  assign n3532 = \i_tv80_core_i_reg_RegsL_reg[5][6]/NET0131  & n2916 ;
  assign n3538 = ~n3531 & ~n3532 ;
  assign n3542 = n3537 & n3538 ;
  assign n3543 = n3541 & n3542 ;
  assign n3544 = n2667 & ~n3543 ;
  assign n3545 = ~n3528 & ~n3544 ;
  assign n3546 = n2711 & ~n3545 ;
  assign n3547 = ~n3519 & ~n3546 ;
  assign n3548 = \i_tv80_core_i_reg_RegsL_reg[1][6]/NET0131  & ~n2937 ;
  assign n3549 = n2937 & ~n3545 ;
  assign n3550 = ~n3548 & ~n3549 ;
  assign n3551 = \i_tv80_core_i_reg_RegsL_reg[2][6]/NET0131  & ~n2941 ;
  assign n3552 = n2941 & ~n3545 ;
  assign n3553 = ~n3551 & ~n3552 ;
  assign n3554 = \i_tv80_core_i_reg_RegsL_reg[3][6]/NET0131  & ~n2945 ;
  assign n3555 = n2945 & ~n3545 ;
  assign n3556 = ~n3554 & ~n3555 ;
  assign n3557 = \i_tv80_core_i_reg_RegsL_reg[4][6]/NET0131  & ~n2949 ;
  assign n3558 = n2949 & ~n3545 ;
  assign n3559 = ~n3557 & ~n3558 ;
  assign n3560 = \i_tv80_core_i_reg_RegsL_reg[5][6]/NET0131  & ~n2953 ;
  assign n3561 = n2953 & ~n3545 ;
  assign n3562 = ~n3560 & ~n3561 ;
  assign n3563 = \i_tv80_core_i_reg_RegsL_reg[6][6]/NET0131  & ~n2957 ;
  assign n3564 = n2957 & ~n3545 ;
  assign n3565 = ~n3563 & ~n3564 ;
  assign n3566 = \i_tv80_core_i_reg_RegsL_reg[7][6]/NET0131  & ~n2961 ;
  assign n3567 = n2961 & ~n3545 ;
  assign n3568 = ~n3566 & ~n3567 ;
  assign n3574 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n532 ;
  assign n3570 = n735 & n796 ;
  assign n3575 = n370 & n682 ;
  assign n3576 = \i_tv80_core_ALU_Op_r_reg[0]/P0001  & ~n625 ;
  assign n3577 = n1175 & n3576 ;
  assign n3578 = ~n3575 & ~n3577 ;
  assign n3579 = \i_tv80_core_BusB_reg[5]/P0001  & ~n3578 ;
  assign n3580 = \i_tv80_core_BusA_reg[5]/P0001  & n700 ;
  assign n3581 = n604 & ~n638 ;
  assign n3582 = ~n3580 & ~n3581 ;
  assign n3571 = ~\i_tv80_core_ALU_Op_r_reg[0]/P0001  & n1175 ;
  assign n3572 = ~\i_tv80_core_BusB_reg[5]/P0001  & ~n682 ;
  assign n3573 = n3571 & ~n3572 ;
  assign n3583 = \i_tv80_core_Save_ALU_r_reg/P0001  & ~n3573 ;
  assign n3584 = n3582 & n3583 ;
  assign n3585 = ~n3579 & n3584 ;
  assign n3586 = ~n3570 & n3585 ;
  assign n3587 = ~n3574 & n3586 ;
  assign n3569 = ~\di_reg_reg[5]/P0001  & ~\i_tv80_core_Save_ALU_r_reg/P0001  ;
  assign n3588 = ~n1172 & ~n3569 ;
  assign n3589 = ~n3587 & n3588 ;
  assign n3590 = \i_tv80_core_BusB_reg[5]/P0001  & n1172 ;
  assign n3591 = ~n3589 & ~n3590 ;
  assign n3592 = n2895 & ~n3591 ;
  assign n3593 = \i_tv80_core_RegBusA_r_reg[13]/P0001  & n2664 ;
  assign n3594 = ~n3592 & ~n3593 ;
  assign n3595 = ~n2667 & ~n3594 ;
  assign n3596 = ~n3375 & ~n3383 ;
  assign n3601 = n2790 & ~n2808 ;
  assign n3602 = n3460 & n3601 ;
  assign n3603 = n2772 & n2863 ;
  assign n3604 = ~n3602 & n3603 ;
  assign n3605 = ~n2824 & n3467 ;
  assign n3606 = ~n3604 & n3605 ;
  assign n3607 = n3284 & n3359 ;
  assign n3608 = n3606 & n3607 ;
  assign n3597 = n2866 & n3305 ;
  assign n3598 = n3284 & ~n3597 ;
  assign n3599 = n3308 & ~n3598 ;
  assign n3600 = n3359 & ~n3599 ;
  assign n3609 = n3382 & ~n3600 ;
  assign n3610 = ~n3608 & n3609 ;
  assign n3611 = n3596 & ~n3610 ;
  assign n3612 = ~n3596 & n3610 ;
  assign n3613 = ~n3611 & ~n3612 ;
  assign n3614 = n2890 & n3613 ;
  assign n3615 = ~n3595 & ~n3614 ;
  assign n3620 = \i_tv80_core_i_reg_RegsH_reg[4][5]/P0001  & n2918 ;
  assign n3621 = \i_tv80_core_i_reg_RegsH_reg[5][5]/P0001  & n2916 ;
  assign n3626 = ~n3620 & ~n3621 ;
  assign n3622 = \i_tv80_core_i_reg_RegsH_reg[7][5]/P0001  & n2904 ;
  assign n3623 = \i_tv80_core_i_reg_RegsH_reg[2][5]/P0001  & n2908 ;
  assign n3627 = ~n3622 & ~n3623 ;
  assign n3628 = n3626 & n3627 ;
  assign n3616 = \i_tv80_core_i_reg_RegsH_reg[6][5]/P0001  & n2920 ;
  assign n3617 = \i_tv80_core_i_reg_RegsH_reg[3][5]/P0001  & n2922 ;
  assign n3624 = ~n3616 & ~n3617 ;
  assign n3618 = \i_tv80_core_i_reg_RegsH_reg[1][5]/P0001  & n2914 ;
  assign n3619 = \i_tv80_core_i_reg_RegsH_reg[0][5]/P0001  & n2911 ;
  assign n3625 = ~n3618 & ~n3619 ;
  assign n3629 = n3624 & n3625 ;
  assign n3630 = n3628 & n3629 ;
  assign n3631 = n2667 & ~n3630 ;
  assign n3632 = n3615 & ~n3631 ;
  assign n3633 = n3456 & ~n3632 ;
  assign n3634 = \i_tv80_core_i_reg_RegsH_reg[0][5]/P0001  & ~n3456 ;
  assign n3635 = ~n3633 & ~n3634 ;
  assign n3636 = n2741 & n3455 ;
  assign n3637 = ~n3358 & ~n3381 ;
  assign n3638 = n3464 & n3466 ;
  assign n3639 = n3301 & ~n3342 ;
  assign n3640 = n3638 & n3639 ;
  assign n3641 = n3458 & n3470 ;
  assign n3642 = ~n3306 & ~n3380 ;
  assign n3643 = n3471 & n3642 ;
  assign n3644 = n3641 & n3643 ;
  assign n3645 = ~n3640 & n3644 ;
  assign n3646 = n3637 & ~n3645 ;
  assign n3647 = ~n3637 & n3645 ;
  assign n3648 = ~n3646 & ~n3647 ;
  assign n3649 = n2892 & n3648 ;
  assign n3659 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n487 ;
  assign n3651 = n735 & ~n788 ;
  assign n3653 = \i_tv80_core_ALU_Op_r_reg[0]/P0001  & n669 ;
  assign n3652 = ~\i_tv80_core_BusB_reg[4]/P0001  & ~n669 ;
  assign n3654 = n1175 & ~n3652 ;
  assign n3655 = ~n3653 & n3654 ;
  assign n3657 = \i_tv80_core_BusA_reg[4]/P0001  & n700 ;
  assign n3656 = n370 & n670 ;
  assign n3658 = n604 & ~n635 ;
  assign n3660 = \i_tv80_core_Save_ALU_r_reg/P0001  & ~n3658 ;
  assign n3661 = ~n3656 & n3660 ;
  assign n3662 = ~n3657 & n3661 ;
  assign n3663 = ~n3655 & n3662 ;
  assign n3664 = ~n3651 & n3663 ;
  assign n3665 = ~n3659 & n3664 ;
  assign n3650 = ~\di_reg_reg[4]/P0001  & ~\i_tv80_core_Save_ALU_r_reg/P0001  ;
  assign n3666 = ~n1172 & ~n3650 ;
  assign n3667 = ~n3665 & n3666 ;
  assign n3668 = \i_tv80_core_BusB_reg[4]/P0001  & n1172 ;
  assign n3669 = ~n3667 & ~n3668 ;
  assign n3670 = n2895 & ~n3669 ;
  assign n3671 = \i_tv80_core_RegBusA_r_reg[12]/P0001  & n2664 ;
  assign n3672 = ~n3670 & ~n3671 ;
  assign n3673 = ~n2667 & ~n3672 ;
  assign n3678 = \i_tv80_core_i_reg_RegsH_reg[4][4]/P0001  & n2918 ;
  assign n3679 = \i_tv80_core_i_reg_RegsH_reg[5][4]/P0001  & n2916 ;
  assign n3684 = ~n3678 & ~n3679 ;
  assign n3680 = \i_tv80_core_i_reg_RegsH_reg[7][4]/P0001  & n2904 ;
  assign n3681 = \i_tv80_core_i_reg_RegsH_reg[2][4]/P0001  & n2908 ;
  assign n3685 = ~n3680 & ~n3681 ;
  assign n3686 = n3684 & n3685 ;
  assign n3674 = \i_tv80_core_i_reg_RegsH_reg[6][4]/P0001  & n2920 ;
  assign n3675 = \i_tv80_core_i_reg_RegsH_reg[3][4]/P0001  & n2922 ;
  assign n3682 = ~n3674 & ~n3675 ;
  assign n3676 = \i_tv80_core_i_reg_RegsH_reg[1][4]/P0001  & n2914 ;
  assign n3677 = \i_tv80_core_i_reg_RegsH_reg[0][4]/P0001  & n2911 ;
  assign n3683 = ~n3676 & ~n3677 ;
  assign n3687 = n3682 & n3683 ;
  assign n3688 = n3686 & n3687 ;
  assign n3689 = n2667 & ~n3688 ;
  assign n3690 = ~n3673 & ~n3689 ;
  assign n3691 = ~n3649 & n3690 ;
  assign n3692 = n3636 & ~n3691 ;
  assign n3693 = \i_tv80_core_i_reg_RegsH_reg[1][4]/P0001  & ~n3636 ;
  assign n3694 = ~n3692 & ~n3693 ;
  assign n3695 = n3507 & ~n3691 ;
  assign n3696 = \i_tv80_core_i_reg_RegsH_reg[3][4]/P0001  & ~n3507 ;
  assign n3697 = ~n3695 & ~n3696 ;
  assign n3698 = n3507 & ~n3632 ;
  assign n3699 = \i_tv80_core_i_reg_RegsH_reg[3][5]/P0001  & ~n3507 ;
  assign n3700 = ~n3698 & ~n3699 ;
  assign n3701 = n3511 & ~n3691 ;
  assign n3702 = \i_tv80_core_i_reg_RegsH_reg[4][4]/P0001  & ~n3511 ;
  assign n3703 = ~n3701 & ~n3702 ;
  assign n3704 = n3511 & ~n3632 ;
  assign n3705 = \i_tv80_core_i_reg_RegsH_reg[4][5]/P0001  & ~n3511 ;
  assign n3706 = ~n3704 & ~n3705 ;
  assign n3707 = n3515 & ~n3691 ;
  assign n3708 = \i_tv80_core_i_reg_RegsH_reg[7][4]/P0001  & ~n3515 ;
  assign n3709 = ~n3707 & ~n3708 ;
  assign n3710 = n3515 & ~n3632 ;
  assign n3711 = \i_tv80_core_i_reg_RegsH_reg[7][5]/P0001  & ~n3515 ;
  assign n3712 = ~n3710 & ~n3711 ;
  assign n3714 = ~n1220 & n2968 ;
  assign n3716 = ~\i_tv80_core_BusB_reg[6]/P0001  & ~n2975 ;
  assign n3717 = ~\i_tv80_core_BusB_reg[2]/P0001  & n2975 ;
  assign n3718 = ~n3716 & ~n3717 ;
  assign n3719 = ~n2973 & ~n3718 ;
  assign n3720 = ~\i_tv80_core_BusA_reg[2]/P0001  & n2973 ;
  assign n3721 = ~n3719 & ~n3720 ;
  assign n3722 = n1157 & ~n3721 ;
  assign n3715 = ~\do[6]_pad  & ~n1157 ;
  assign n3723 = ~n2968 & ~n3715 ;
  assign n3724 = ~n3722 & n3723 ;
  assign n3725 = ~\i_tv80_core_BusAck_reg/P0001  & ~n3724 ;
  assign n3726 = ~n3714 & n3725 ;
  assign n3713 = ~\do[6]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n3727 = reset_n_pad & ~n3713 ;
  assign n3728 = ~n3726 & n3727 ;
  assign n3733 = ~n3058 & ~n3068 ;
  assign n3734 = n3052 & ~n3067 ;
  assign n3735 = ~n3064 & ~n3734 ;
  assign n3736 = n3733 & ~n3735 ;
  assign n3737 = ~n3733 & n3735 ;
  assign n3738 = ~n3736 & ~n3737 ;
  assign n3739 = n3001 & ~n3738 ;
  assign n3732 = \i_tv80_core_SP_reg[6]/P0001  & ~n3002 ;
  assign n3740 = ~n2997 & ~n3732 ;
  assign n3741 = ~n3739 & n3740 ;
  assign n3731 = n1777 & n2997 ;
  assign n3742 = ~n1113 & ~n3731 ;
  assign n3743 = ~n3741 & n3742 ;
  assign n3744 = \i_tv80_core_SP_reg[6]/P0001  & n1113 ;
  assign n3745 = ~n2992 & ~n3744 ;
  assign n3746 = ~n3743 & n3745 ;
  assign n3730 = n1220 & n2992 ;
  assign n3747 = ~\i_tv80_core_BusAck_reg/P0001  & ~n3730 ;
  assign n3748 = ~n3746 & n3747 ;
  assign n3729 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[6]/P0001  ;
  assign n3749 = reset_n_pad & ~n3729 ;
  assign n3750 = ~n3748 & n3749 ;
  assign n3777 = \i_tv80_core_Ap_reg[3]/P0001  & n1117 ;
  assign n3778 = ~\i_tv80_core_ACC_reg[3]/P0001  & n3155 ;
  assign n3779 = ~n3777 & ~n3778 ;
  assign n3780 = ~n1113 & ~n3779 ;
  assign n3781 = \i_tv80_core_ACC_reg[3]/P0001  & n3160 ;
  assign n3782 = ~n3780 & ~n3781 ;
  assign n3783 = ~n1112 & ~n3782 ;
  assign n3773 = \i_tv80_core_I_reg[3]/P0001  & ~n3147 ;
  assign n3774 = \i_tv80_core_R_reg[3]/P0001  & n3145 ;
  assign n3775 = ~n3773 & ~n3774 ;
  assign n3776 = n1111 & ~n3775 ;
  assign n3784 = ~n3143 & ~n3776 ;
  assign n3785 = ~n3783 & n3784 ;
  assign n3753 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n566 ;
  assign n3760 = n735 & ~n823 ;
  assign n3758 = n700 & ~n724 ;
  assign n3759 = n604 & ~n610 ;
  assign n3761 = ~n3758 & ~n3759 ;
  assign n3762 = ~n3760 & n3761 ;
  assign n3752 = n679 & n3571 ;
  assign n3755 = ~n679 & ~n1175 ;
  assign n3754 = ~n370 & n679 ;
  assign n3756 = \i_tv80_core_BusB_reg[3]/P0001  & ~n3754 ;
  assign n3757 = ~n3755 & n3756 ;
  assign n3763 = ~n3752 & ~n3757 ;
  assign n3764 = n3762 & n3763 ;
  assign n3765 = ~n3753 & n3764 ;
  assign n3766 = \i_tv80_core_Save_ALU_r_reg/P0001  & ~n3765 ;
  assign n3767 = \di_reg_reg[3]/P0001  & ~\i_tv80_core_Save_ALU_r_reg/P0001  ;
  assign n3768 = ~n3766 & ~n3767 ;
  assign n3769 = ~n1172 & ~n3768 ;
  assign n3770 = \i_tv80_core_BusB_reg[3]/P0001  & n1172 ;
  assign n3771 = ~n3769 & ~n3770 ;
  assign n3772 = n3143 & n3771 ;
  assign n3786 = ~\i_tv80_core_BusAck_reg/P0001  & ~n3772 ;
  assign n3787 = ~n3785 & n3786 ;
  assign n3751 = \i_tv80_core_ACC_reg[3]/P0001  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n3788 = reset_n_pad & ~n3751 ;
  assign n3789 = ~n3787 & n3788 ;
  assign n3796 = \i_tv80_core_Ap_reg[5]/P0001  & n1117 ;
  assign n3797 = ~\i_tv80_core_ACC_reg[5]/P0001  & n3155 ;
  assign n3798 = ~n3796 & ~n3797 ;
  assign n3799 = ~n1113 & ~n3798 ;
  assign n3800 = \i_tv80_core_ACC_reg[5]/P0001  & n3160 ;
  assign n3801 = ~n3799 & ~n3800 ;
  assign n3802 = ~n1112 & ~n3801 ;
  assign n3792 = \i_tv80_core_I_reg[5]/P0001  & ~n3147 ;
  assign n3793 = \i_tv80_core_R_reg[5]/P0001  & n3145 ;
  assign n3794 = ~n3792 & ~n3793 ;
  assign n3795 = n1111 & ~n3794 ;
  assign n3803 = ~n3143 & ~n3795 ;
  assign n3804 = ~n3802 & n3803 ;
  assign n3791 = n3143 & n3591 ;
  assign n3805 = ~\i_tv80_core_BusAck_reg/P0001  & ~n3791 ;
  assign n3806 = ~n3804 & n3805 ;
  assign n3790 = \i_tv80_core_ACC_reg[5]/P0001  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n3807 = reset_n_pad & ~n3790 ;
  assign n3808 = ~n3806 & n3807 ;
  assign n3815 = \i_tv80_core_Ap_reg[6]/P0001  & n1117 ;
  assign n3816 = ~\i_tv80_core_ACC_reg[6]/P0001  & n3155 ;
  assign n3817 = ~n3815 & ~n3816 ;
  assign n3818 = ~n1113 & ~n3817 ;
  assign n3819 = \i_tv80_core_ACC_reg[6]/P0001  & n3160 ;
  assign n3820 = ~n3818 & ~n3819 ;
  assign n3821 = ~n1112 & ~n3820 ;
  assign n3811 = \i_tv80_core_R_reg[6]/P0001  & n3145 ;
  assign n3812 = \i_tv80_core_I_reg[6]/P0001  & ~n3147 ;
  assign n3813 = ~n3811 & ~n3812 ;
  assign n3814 = n1111 & ~n3813 ;
  assign n3822 = ~n3143 & ~n3814 ;
  assign n3823 = ~n3821 & n3822 ;
  assign n3810 = n1220 & n3143 ;
  assign n3824 = ~\i_tv80_core_BusAck_reg/P0001  & ~n3810 ;
  assign n3825 = ~n3823 & n3824 ;
  assign n3809 = \i_tv80_core_ACC_reg[6]/P0001  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n3826 = reset_n_pad & ~n3809 ;
  assign n3827 = ~n3825 & n3826 ;
  assign n3828 = ~n2205 & n2997 ;
  assign n3829 = \i_tv80_core_SP_reg[14]/P0001  & ~n3002 ;
  assign n3830 = ~n3185 & ~n3226 ;
  assign n3831 = n3065 & ~n3734 ;
  assign n3832 = ~n3068 & ~n3831 ;
  assign n3833 = ~n3011 & ~n3832 ;
  assign n3834 = ~n3010 & ~n3833 ;
  assign n3835 = ~n3190 & ~n3203 ;
  assign n3836 = ~n3834 & n3835 ;
  assign n3837 = ~n3193 & ~n3206 ;
  assign n3838 = ~n3836 & n3837 ;
  assign n3839 = ~n3199 & ~n3213 ;
  assign n3840 = ~n3181 & ~n3217 ;
  assign n3841 = n3839 & n3840 ;
  assign n3842 = ~n3838 & n3841 ;
  assign n3843 = ~n3207 & ~n3222 ;
  assign n3844 = ~n3221 & ~n3223 ;
  assign n3845 = n3843 & n3844 ;
  assign n3846 = ~n3842 & n3845 ;
  assign n3847 = n3830 & ~n3846 ;
  assign n3848 = ~n3830 & n3846 ;
  assign n3849 = ~n3847 & ~n3848 ;
  assign n3850 = n2699 & n3849 ;
  assign n3851 = ~n3829 & ~n3850 ;
  assign n3852 = ~\i_tv80_core_SP_reg[14]/P0001  & n3000 ;
  assign n3853 = ~n2997 & ~n3852 ;
  assign n3854 = ~n3851 & n3853 ;
  assign n3855 = ~n3828 & ~n3854 ;
  assign n3856 = ~n1113 & ~n3855 ;
  assign n3857 = \i_tv80_core_SP_reg[14]/P0001  & n1113 ;
  assign n3858 = ~n3242 & ~n3857 ;
  assign n3859 = ~n3856 & n3858 ;
  assign n3860 = n1220 & n3242 ;
  assign n3861 = ~\i_tv80_core_BusAck_reg/P0001  & ~n3860 ;
  assign n3862 = ~n3859 & n3861 ;
  assign n3863 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[14]/P0001  ;
  assign n3864 = reset_n_pad & ~n3863 ;
  assign n3865 = ~n3862 & n3864 ;
  assign n3866 = ~n3267 & ~n3306 ;
  assign n3867 = ~n3473 & n3866 ;
  assign n3868 = n3473 & ~n3866 ;
  assign n3869 = ~n3867 & ~n3868 ;
  assign n3870 = n2890 & n3869 ;
  assign n3871 = \i_tv80_core_RegBusA_r_reg[10]/P0001  & n2664 ;
  assign n3872 = ~n1193 & n2895 ;
  assign n3873 = ~n3871 & ~n3872 ;
  assign n3874 = ~n2667 & ~n3873 ;
  assign n3879 = \i_tv80_core_i_reg_RegsH_reg[4][2]/P0001  & n2918 ;
  assign n3880 = \i_tv80_core_i_reg_RegsH_reg[5][2]/P0001  & n2916 ;
  assign n3885 = ~n3879 & ~n3880 ;
  assign n3881 = \i_tv80_core_i_reg_RegsH_reg[7][2]/P0001  & n2904 ;
  assign n3882 = \i_tv80_core_i_reg_RegsH_reg[2][2]/P0001  & n2908 ;
  assign n3886 = ~n3881 & ~n3882 ;
  assign n3887 = n3885 & n3886 ;
  assign n3875 = \i_tv80_core_i_reg_RegsH_reg[6][2]/P0001  & n2920 ;
  assign n3876 = \i_tv80_core_i_reg_RegsH_reg[3][2]/P0001  & n2922 ;
  assign n3883 = ~n3875 & ~n3876 ;
  assign n3877 = \i_tv80_core_i_reg_RegsH_reg[1][2]/P0001  & n2914 ;
  assign n3878 = \i_tv80_core_i_reg_RegsH_reg[0][2]/P0001  & n2911 ;
  assign n3884 = ~n3877 & ~n3878 ;
  assign n3888 = n3883 & n3884 ;
  assign n3889 = n3887 & n3888 ;
  assign n3890 = n2667 & ~n3889 ;
  assign n3891 = ~n3874 & ~n3890 ;
  assign n3892 = ~n3870 & n3891 ;
  assign n3893 = n3456 & ~n3892 ;
  assign n3894 = \i_tv80_core_i_reg_RegsH_reg[0][2]/P0001  & ~n3456 ;
  assign n3895 = ~n3893 & ~n3894 ;
  assign n3896 = n3507 & ~n3892 ;
  assign n3897 = \i_tv80_core_i_reg_RegsH_reg[3][2]/P0001  & ~n3507 ;
  assign n3898 = ~n3896 & ~n3897 ;
  assign n3899 = n3511 & ~n3892 ;
  assign n3900 = \i_tv80_core_i_reg_RegsH_reg[4][2]/P0001  & ~n3511 ;
  assign n3901 = ~n3899 & ~n3900 ;
  assign n3902 = n3515 & ~n3892 ;
  assign n3903 = \i_tv80_core_i_reg_RegsH_reg[7][2]/P0001  & ~n3515 ;
  assign n3904 = ~n3902 & ~n3903 ;
  assign n3911 = \i_tv80_core_Ap_reg[2]/P0001  & n1117 ;
  assign n3912 = ~\i_tv80_core_ACC_reg[2]/P0001  & n3155 ;
  assign n3913 = ~n3911 & ~n3912 ;
  assign n3914 = ~n1113 & ~n3913 ;
  assign n3915 = \i_tv80_core_ACC_reg[2]/P0001  & n3160 ;
  assign n3916 = ~n3914 & ~n3915 ;
  assign n3917 = ~n1112 & ~n3916 ;
  assign n3907 = \i_tv80_core_I_reg[2]/P0001  & ~n3147 ;
  assign n3908 = \i_tv80_core_R_reg[2]/P0001  & n3145 ;
  assign n3909 = ~n3907 & ~n3908 ;
  assign n3910 = n1111 & ~n3909 ;
  assign n3918 = ~n3143 & ~n3910 ;
  assign n3919 = ~n3917 & n3918 ;
  assign n3906 = n1193 & n3143 ;
  assign n3920 = ~\i_tv80_core_BusAck_reg/P0001  & ~n3906 ;
  assign n3921 = ~n3919 & n3920 ;
  assign n3905 = \i_tv80_core_ACC_reg[2]/P0001  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n3922 = reset_n_pad & ~n3905 ;
  assign n3923 = ~n3921 & n3922 ;
  assign n3930 = \i_tv80_core_Ap_reg[4]/P0001  & n1117 ;
  assign n3931 = ~\i_tv80_core_ACC_reg[4]/P0001  & n3155 ;
  assign n3932 = ~n3930 & ~n3931 ;
  assign n3933 = ~n1113 & ~n3932 ;
  assign n3934 = \i_tv80_core_ACC_reg[4]/P0001  & n3160 ;
  assign n3935 = ~n3933 & ~n3934 ;
  assign n3936 = ~n1112 & ~n3935 ;
  assign n3926 = \i_tv80_core_R_reg[4]/P0001  & n3145 ;
  assign n3927 = \i_tv80_core_I_reg[4]/P0001  & ~n3147 ;
  assign n3928 = ~n3926 & ~n3927 ;
  assign n3929 = n1111 & ~n3928 ;
  assign n3937 = ~n3143 & ~n3929 ;
  assign n3938 = ~n3936 & n3937 ;
  assign n3925 = n3143 & n3669 ;
  assign n3939 = ~\i_tv80_core_BusAck_reg/P0001  & ~n3925 ;
  assign n3940 = ~n3938 & n3939 ;
  assign n3924 = \i_tv80_core_ACC_reg[4]/P0001  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n3941 = reset_n_pad & ~n3924 ;
  assign n3942 = ~n3940 & n3941 ;
  assign n3949 = \i_tv80_core_Ap_reg[0]/P0001  & n1117 ;
  assign n3950 = ~\i_tv80_core_ACC_reg[0]/P0001  & n3155 ;
  assign n3951 = ~n3949 & ~n3950 ;
  assign n3952 = ~n1113 & ~n3951 ;
  assign n3953 = \i_tv80_core_ACC_reg[0]/P0001  & n3160 ;
  assign n3954 = ~n3952 & ~n3953 ;
  assign n3955 = ~n1112 & ~n3954 ;
  assign n3945 = \i_tv80_core_I_reg[0]/P0001  & ~n3147 ;
  assign n3946 = \i_tv80_core_R_reg[0]/P0001  & n3145 ;
  assign n3947 = ~n3945 & ~n3946 ;
  assign n3948 = n1111 & ~n3947 ;
  assign n3956 = ~n3143 & ~n3948 ;
  assign n3957 = ~n3955 & n3956 ;
  assign n3944 = n3107 & n3143 ;
  assign n3958 = ~\i_tv80_core_BusAck_reg/P0001  & ~n3944 ;
  assign n3959 = ~n3957 & n3958 ;
  assign n3943 = \i_tv80_core_ACC_reg[0]/P0001  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n3960 = reset_n_pad & ~n3943 ;
  assign n3961 = ~n3959 & n3960 ;
  assign n3988 = \i_tv80_core_Ap_reg[1]/P0001  & n1117 ;
  assign n3989 = ~\i_tv80_core_ACC_reg[1]/P0001  & n3155 ;
  assign n3990 = ~n3988 & ~n3989 ;
  assign n3991 = ~n1113 & ~n3990 ;
  assign n3992 = \i_tv80_core_ACC_reg[1]/P0001  & n3160 ;
  assign n3993 = ~n3991 & ~n3992 ;
  assign n3994 = ~n1112 & ~n3993 ;
  assign n3984 = \i_tv80_core_R_reg[1]/P0001  & n3145 ;
  assign n3985 = \i_tv80_core_I_reg[1]/P0001  & ~n3147 ;
  assign n3986 = ~n3984 & ~n3985 ;
  assign n3987 = n1111 & ~n3986 ;
  assign n3995 = ~n3143 & ~n3987 ;
  assign n3996 = ~n3994 & n3995 ;
  assign n3964 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n503 ;
  assign n3963 = n735 & n741 ;
  assign n3966 = \i_tv80_core_ALU_Op_r_reg[0]/P0001  & n686 ;
  assign n3965 = ~\i_tv80_core_BusB_reg[1]/P0001  & ~n686 ;
  assign n3967 = n1175 & ~n3965 ;
  assign n3968 = ~n3966 & n3967 ;
  assign n3970 = n370 & n687 ;
  assign n3969 = n700 & ~n718 ;
  assign n3971 = n604 & ~n607 ;
  assign n3972 = ~n3969 & ~n3971 ;
  assign n3973 = ~n3970 & n3972 ;
  assign n3974 = ~n3968 & n3973 ;
  assign n3975 = ~n3963 & n3974 ;
  assign n3976 = ~n3964 & n3975 ;
  assign n3977 = \i_tv80_core_Save_ALU_r_reg/P0001  & ~n3976 ;
  assign n3978 = \di_reg_reg[1]/P0001  & ~\i_tv80_core_Save_ALU_r_reg/P0001  ;
  assign n3979 = ~n3977 & ~n3978 ;
  assign n3980 = ~n1172 & ~n3979 ;
  assign n3981 = \i_tv80_core_BusB_reg[1]/P0001  & n1172 ;
  assign n3982 = ~n3980 & ~n3981 ;
  assign n3983 = n3143 & n3982 ;
  assign n3997 = ~\i_tv80_core_BusAck_reg/P0001  & ~n3983 ;
  assign n3998 = ~n3996 & n3997 ;
  assign n3962 = \i_tv80_core_ACC_reg[1]/P0001  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n3999 = reset_n_pad & ~n3962 ;
  assign n4000 = ~n3998 & n3999 ;
  assign n4005 = \i_tv80_core_i_reg_RegsH_reg[3][3]/P0001  & n2922 ;
  assign n4006 = \i_tv80_core_i_reg_RegsH_reg[2][3]/P0001  & n2908 ;
  assign n4011 = ~n4005 & ~n4006 ;
  assign n4007 = \i_tv80_core_i_reg_RegsH_reg[7][3]/P0001  & n2904 ;
  assign n4008 = \i_tv80_core_i_reg_RegsH_reg[0][3]/P0001  & n2911 ;
  assign n4012 = ~n4007 & ~n4008 ;
  assign n4013 = n4011 & n4012 ;
  assign n4001 = \i_tv80_core_i_reg_RegsH_reg[6][3]/P0001  & n2920 ;
  assign n4002 = \i_tv80_core_i_reg_RegsH_reg[1][3]/P0001  & n2914 ;
  assign n4009 = ~n4001 & ~n4002 ;
  assign n4003 = \i_tv80_core_i_reg_RegsH_reg[4][3]/P0001  & n2918 ;
  assign n4004 = \i_tv80_core_i_reg_RegsH_reg[5][3]/P0001  & n2916 ;
  assign n4010 = ~n4003 & ~n4004 ;
  assign n4014 = n4009 & n4010 ;
  assign n4015 = n4013 & n4014 ;
  assign n4016 = n2667 & n4015 ;
  assign n4018 = ~n3342 & ~n3380 ;
  assign n4019 = ~n3310 & n4018 ;
  assign n4020 = n3310 & ~n4018 ;
  assign n4021 = ~n4019 & ~n4020 ;
  assign n4022 = n2891 & n4021 ;
  assign n4017 = n2895 & ~n3771 ;
  assign n4023 = \i_tv80_core_RegBusA_r_reg[11]/P0001  & n2664 ;
  assign n4024 = ~n2667 & ~n4023 ;
  assign n4025 = ~n4017 & n4024 ;
  assign n4026 = ~n4022 & n4025 ;
  assign n4027 = ~n4016 & ~n4026 ;
  assign n4028 = n3456 & ~n4027 ;
  assign n4029 = ~\i_tv80_core_i_reg_RegsH_reg[0][3]/P0001  & ~n3456 ;
  assign n4030 = ~n4028 & ~n4029 ;
  assign n4031 = n3636 & ~n4027 ;
  assign n4032 = ~\i_tv80_core_i_reg_RegsH_reg[1][3]/P0001  & ~n3636 ;
  assign n4033 = ~n4031 & ~n4032 ;
  assign n4034 = n2745 & n3455 ;
  assign n4035 = n3597 & ~n3606 ;
  assign n4036 = ~n3283 & ~n3307 ;
  assign n4037 = ~n4035 & n4036 ;
  assign n4038 = n4035 & ~n4036 ;
  assign n4039 = ~n4037 & ~n4038 ;
  assign n4040 = n2892 & n4039 ;
  assign n4041 = \i_tv80_core_RegBusA_r_reg[9]/P0001  & n2664 ;
  assign n4042 = n2895 & ~n3982 ;
  assign n4043 = ~n4041 & ~n4042 ;
  assign n4044 = ~n2667 & ~n4043 ;
  assign n4049 = \i_tv80_core_i_reg_RegsH_reg[4][1]/P0001  & n2918 ;
  assign n4050 = \i_tv80_core_i_reg_RegsH_reg[5][1]/P0001  & n2916 ;
  assign n4055 = ~n4049 & ~n4050 ;
  assign n4051 = \i_tv80_core_i_reg_RegsH_reg[7][1]/P0001  & n2904 ;
  assign n4052 = \i_tv80_core_i_reg_RegsH_reg[2][1]/P0001  & n2908 ;
  assign n4056 = ~n4051 & ~n4052 ;
  assign n4057 = n4055 & n4056 ;
  assign n4045 = \i_tv80_core_i_reg_RegsH_reg[6][1]/P0001  & n2920 ;
  assign n4046 = \i_tv80_core_i_reg_RegsH_reg[3][1]/P0001  & n2922 ;
  assign n4053 = ~n4045 & ~n4046 ;
  assign n4047 = \i_tv80_core_i_reg_RegsH_reg[1][1]/P0001  & n2914 ;
  assign n4048 = \i_tv80_core_i_reg_RegsH_reg[0][1]/P0001  & n2911 ;
  assign n4054 = ~n4047 & ~n4048 ;
  assign n4058 = n4053 & n4054 ;
  assign n4059 = n4057 & n4058 ;
  assign n4060 = n2667 & ~n4059 ;
  assign n4061 = ~n4044 & ~n4060 ;
  assign n4062 = ~n4040 & n4061 ;
  assign n4063 = n4034 & ~n4062 ;
  assign n4064 = \i_tv80_core_i_reg_RegsH_reg[2][1]/P0001  & ~n4034 ;
  assign n4065 = ~n4063 & ~n4064 ;
  assign n4066 = ~n4027 & n4034 ;
  assign n4067 = ~\i_tv80_core_i_reg_RegsH_reg[2][3]/P0001  & ~n4034 ;
  assign n4068 = ~n4066 & ~n4067 ;
  assign n4069 = n3507 & ~n4062 ;
  assign n4070 = \i_tv80_core_i_reg_RegsH_reg[3][1]/P0001  & ~n3507 ;
  assign n4071 = ~n4069 & ~n4070 ;
  assign n4072 = n3507 & ~n4027 ;
  assign n4073 = ~\i_tv80_core_i_reg_RegsH_reg[3][3]/P0001  & ~n3507 ;
  assign n4074 = ~n4072 & ~n4073 ;
  assign n4075 = n3511 & ~n4062 ;
  assign n4076 = \i_tv80_core_i_reg_RegsH_reg[4][1]/P0001  & ~n3511 ;
  assign n4077 = ~n4075 & ~n4076 ;
  assign n4078 = n3511 & ~n4027 ;
  assign n4079 = ~\i_tv80_core_i_reg_RegsH_reg[4][3]/P0001  & ~n3511 ;
  assign n4080 = ~n4078 & ~n4079 ;
  assign n4081 = n2739 & n3455 ;
  assign n4082 = ~n4062 & n4081 ;
  assign n4083 = \i_tv80_core_i_reg_RegsH_reg[5][1]/P0001  & ~n4081 ;
  assign n4084 = ~n4082 & ~n4083 ;
  assign n4085 = ~n4027 & n4081 ;
  assign n4086 = ~\i_tv80_core_i_reg_RegsH_reg[5][3]/P0001  & ~n4081 ;
  assign n4087 = ~n4085 & ~n4086 ;
  assign n4088 = n2736 & n3455 ;
  assign n4089 = ~n4027 & n4088 ;
  assign n4090 = ~\i_tv80_core_i_reg_RegsH_reg[6][3]/P0001  & ~n4088 ;
  assign n4091 = ~n4089 & ~n4090 ;
  assign n4092 = n3515 & ~n4062 ;
  assign n4093 = \i_tv80_core_i_reg_RegsH_reg[7][1]/P0001  & ~n3515 ;
  assign n4094 = ~n4092 & ~n4093 ;
  assign n4095 = n3515 & ~n4027 ;
  assign n4096 = ~\i_tv80_core_i_reg_RegsH_reg[7][3]/P0001  & ~n3515 ;
  assign n4097 = ~n4095 & ~n4096 ;
  assign n4102 = \i_tv80_core_i_reg_RegsH_reg[7][0]/P0001  & n2904 ;
  assign n4103 = \i_tv80_core_i_reg_RegsH_reg[6][0]/P0001  & n2920 ;
  assign n4108 = ~n4102 & ~n4103 ;
  assign n4104 = \i_tv80_core_i_reg_RegsH_reg[3][0]/P0001  & n2922 ;
  assign n4105 = \i_tv80_core_i_reg_RegsH_reg[5][0]/P0001  & n2916 ;
  assign n4109 = ~n4104 & ~n4105 ;
  assign n4110 = n4108 & n4109 ;
  assign n4098 = \i_tv80_core_i_reg_RegsH_reg[2][0]/P0001  & n2908 ;
  assign n4099 = \i_tv80_core_i_reg_RegsH_reg[4][0]/P0001  & n2918 ;
  assign n4106 = ~n4098 & ~n4099 ;
  assign n4100 = \i_tv80_core_i_reg_RegsH_reg[1][0]/P0001  & n2914 ;
  assign n4101 = \i_tv80_core_i_reg_RegsH_reg[0][0]/P0001  & n2911 ;
  assign n4107 = ~n4100 & ~n4101 ;
  assign n4111 = n4106 & n4107 ;
  assign n4112 = n4110 & n4111 ;
  assign n4113 = n2667 & ~n4112 ;
  assign n4115 = ~n3638 & n3641 ;
  assign n4116 = ~n3300 & ~n3304 ;
  assign n4117 = ~n4115 & n4116 ;
  assign n4118 = n4115 & ~n4116 ;
  assign n4119 = ~n4117 & ~n4118 ;
  assign n4120 = n2891 & n4119 ;
  assign n4114 = \i_tv80_core_RegBusA_r_reg[8]/P0001  & n2664 ;
  assign n4121 = n2895 & ~n3107 ;
  assign n4122 = ~n4114 & ~n4121 ;
  assign n4123 = ~n4120 & n4122 ;
  assign n4124 = ~n2667 & ~n4123 ;
  assign n4125 = ~n4113 & ~n4124 ;
  assign n4126 = n3636 & ~n4125 ;
  assign n4127 = \i_tv80_core_i_reg_RegsH_reg[1][0]/P0001  & ~n3636 ;
  assign n4128 = ~n4126 & ~n4127 ;
  assign n4129 = n4034 & ~n4125 ;
  assign n4130 = \i_tv80_core_i_reg_RegsH_reg[2][0]/P0001  & ~n4034 ;
  assign n4131 = ~n4129 & ~n4130 ;
  assign n4132 = n3507 & ~n4125 ;
  assign n4133 = \i_tv80_core_i_reg_RegsH_reg[3][0]/P0001  & ~n3507 ;
  assign n4134 = ~n4132 & ~n4133 ;
  assign n4135 = n3511 & ~n4125 ;
  assign n4136 = \i_tv80_core_i_reg_RegsH_reg[4][0]/P0001  & ~n3511 ;
  assign n4137 = ~n4135 & ~n4136 ;
  assign n4138 = n4081 & ~n4125 ;
  assign n4139 = \i_tv80_core_i_reg_RegsH_reg[5][0]/P0001  & ~n4081 ;
  assign n4140 = ~n4138 & ~n4139 ;
  assign n4141 = n4088 & ~n4125 ;
  assign n4142 = \i_tv80_core_i_reg_RegsH_reg[6][0]/P0001  & ~n4088 ;
  assign n4143 = ~n4141 & ~n4142 ;
  assign n4144 = n3515 & ~n4125 ;
  assign n4145 = \i_tv80_core_i_reg_RegsH_reg[7][0]/P0001  & ~n3515 ;
  assign n4146 = ~n4144 & ~n4145 ;
  assign n4148 = n1167 & ~n3982 ;
  assign n4150 = ~\i_tv80_core_F_reg[1]/P0001  & ~n3154 ;
  assign n4151 = ~n3127 & ~n4150 ;
  assign n4152 = ~n1117 & ~n4151 ;
  assign n4149 = n386 & ~n1113 ;
  assign n4153 = ~\i_tv80_core_Fp_reg[1]/P0001  & n1117 ;
  assign n4154 = n4149 & ~n4153 ;
  assign n4155 = ~n4152 & n4154 ;
  assign n4156 = \i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~\i_tv80_core_F_reg[1]/P0001  ;
  assign n4157 = ~n696 & ~n735 ;
  assign n4158 = ~n4156 & ~n4157 ;
  assign n4159 = ~n386 & n4158 ;
  assign n4160 = \i_tv80_core_F_reg[1]/P0001  & n1113 ;
  assign n4161 = n386 & n4160 ;
  assign n4162 = ~n4159 & ~n4161 ;
  assign n4163 = ~n4155 & n4162 ;
  assign n4164 = ~\i_tv80_core_IR_reg[0]/P0001  & n1156 ;
  assign n4165 = n1129 & n4164 ;
  assign n4166 = ~n1167 & ~n4165 ;
  assign n4167 = ~n1105 & n4166 ;
  assign n4168 = ~n4163 & n4167 ;
  assign n4169 = ~n4148 & ~n4168 ;
  assign n4170 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4169 ;
  assign n4147 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_F_reg[1]/P0001  ;
  assign n4171 = reset_n_pad & ~n4147 ;
  assign n4172 = ~n4170 & n4171 ;
  assign n4187 = ~n3126 & ~n3153 ;
  assign n4188 = n1103 & ~n4187 ;
  assign n4189 = ~n1113 & n4188 ;
  assign n4190 = ~n1118 & ~n4189 ;
  assign n4191 = ~\i_tv80_core_F_reg[3]/P0001  & n4190 ;
  assign n4193 = ~\i_tv80_core_ACC_reg[3]/P0001  & ~n3126 ;
  assign n4194 = \i_tv80_core_ACC_reg[3]/P0001  & n3126 ;
  assign n4195 = ~n4193 & ~n4194 ;
  assign n4196 = n4188 & n4195 ;
  assign n4197 = ~n1117 & ~n4196 ;
  assign n4192 = \i_tv80_core_Fp_reg[3]/P0001  & n1117 ;
  assign n4198 = ~n1113 & ~n4192 ;
  assign n4199 = ~n4197 & n4198 ;
  assign n4200 = ~n4191 & ~n4199 ;
  assign n4201 = n386 & ~n4200 ;
  assign n4180 = n566 & ~n1159 ;
  assign n4179 = ~\i_tv80_core_BusB_reg[3]/P0001  & n1159 ;
  assign n4181 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n4179 ;
  assign n4182 = ~n4180 & n4181 ;
  assign n4176 = n370 & ~n886 ;
  assign n4177 = \i_tv80_core_BusB_reg[3]/P0001  & n4176 ;
  assign n4178 = \i_tv80_core_F_reg[3]/P0001  & n697 ;
  assign n4183 = ~n4177 & ~n4178 ;
  assign n4184 = ~n386 & n4183 ;
  assign n4185 = n3762 & n4184 ;
  assign n4186 = ~n4182 & n4185 ;
  assign n4202 = ~n4165 & ~n4186 ;
  assign n4203 = ~n4201 & n4202 ;
  assign n4175 = ~n3765 & n4165 ;
  assign n4204 = ~n1167 & ~n4175 ;
  assign n4205 = ~n4203 & n4204 ;
  assign n4174 = n1167 & n3771 ;
  assign n4206 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4174 ;
  assign n4207 = ~n4205 & n4206 ;
  assign n4173 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_F_reg[3]/P0001  ;
  assign n4208 = reset_n_pad & ~n4173 ;
  assign n4209 = ~n4207 & n4208 ;
  assign n4213 = ~\i_tv80_core_F_reg[5]/P0001  & n4190 ;
  assign n4215 = ~\i_tv80_core_ACC_reg[5]/P0001  & ~n3126 ;
  assign n4216 = \i_tv80_core_ACC_reg[5]/P0001  & n3126 ;
  assign n4217 = ~n4215 & ~n4216 ;
  assign n4218 = n4188 & n4217 ;
  assign n4219 = ~n1117 & ~n4218 ;
  assign n4214 = \i_tv80_core_Fp_reg[5]/P0001  & n1117 ;
  assign n4220 = ~n1113 & ~n4214 ;
  assign n4221 = ~n4219 & n4220 ;
  assign n4222 = ~n4213 & ~n4221 ;
  assign n4223 = n386 & ~n4222 ;
  assign n4227 = n532 & ~n1159 ;
  assign n4226 = ~\i_tv80_core_BusB_reg[5]/P0001  & n1159 ;
  assign n4228 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n4226 ;
  assign n4229 = ~n4227 & n4228 ;
  assign n4224 = \i_tv80_core_F_reg[5]/P0001  & n697 ;
  assign n4225 = \i_tv80_core_BusB_reg[5]/P0001  & n4176 ;
  assign n4230 = ~n4224 & ~n4225 ;
  assign n4231 = n3582 & n4230 ;
  assign n4232 = ~n386 & n4231 ;
  assign n4233 = ~n3570 & n4232 ;
  assign n4234 = ~n4229 & n4233 ;
  assign n4235 = ~n4165 & ~n4234 ;
  assign n4236 = ~n4223 & n4235 ;
  assign n4212 = ~n3976 & n4165 ;
  assign n4237 = ~n1167 & ~n4212 ;
  assign n4238 = ~n4236 & n4237 ;
  assign n4211 = n1167 & n3591 ;
  assign n4239 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4211 ;
  assign n4240 = ~n4238 & n4239 ;
  assign n4210 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_F_reg[5]/P0001  ;
  assign n4241 = reset_n_pad & ~n4210 ;
  assign n4242 = ~n4240 & n4241 ;
  assign n4243 = \i_tv80_core_i_reg_RegsL_reg[0][5]/NET0131  & ~n2711 ;
  assign n4244 = ~n2824 & ~n2864 ;
  assign n4245 = n3604 & ~n4244 ;
  assign n4246 = ~n3604 & n4244 ;
  assign n4247 = ~n4245 & ~n4246 ;
  assign n4248 = n2891 & n4247 ;
  assign n4249 = \i_tv80_core_RegBusA_r_reg[5]/P0001  & n2664 ;
  assign n4250 = ~n3592 & ~n4249 ;
  assign n4251 = ~n4248 & n4250 ;
  assign n4252 = ~n2667 & ~n4251 ;
  assign n4257 = \i_tv80_core_i_reg_RegsL_reg[1][5]/NET0131  & n2914 ;
  assign n4258 = \i_tv80_core_i_reg_RegsL_reg[0][5]/NET0131  & n2911 ;
  assign n4263 = ~n4257 & ~n4258 ;
  assign n4259 = \i_tv80_core_i_reg_RegsL_reg[3][5]/NET0131  & n2922 ;
  assign n4260 = \i_tv80_core_i_reg_RegsL_reg[5][5]/NET0131  & n2916 ;
  assign n4264 = ~n4259 & ~n4260 ;
  assign n4265 = n4263 & n4264 ;
  assign n4253 = \i_tv80_core_i_reg_RegsL_reg[2][5]/NET0131  & n2908 ;
  assign n4254 = \i_tv80_core_i_reg_RegsL_reg[4][5]/NET0131  & n2918 ;
  assign n4261 = ~n4253 & ~n4254 ;
  assign n4255 = \i_tv80_core_i_reg_RegsL_reg[7][5]/NET0131  & n2904 ;
  assign n4256 = \i_tv80_core_i_reg_RegsL_reg[6][5]/NET0131  & n2920 ;
  assign n4262 = ~n4255 & ~n4256 ;
  assign n4266 = n4261 & n4262 ;
  assign n4267 = n4265 & n4266 ;
  assign n4268 = n2667 & ~n4267 ;
  assign n4269 = ~n4252 & ~n4268 ;
  assign n4270 = n2711 & ~n4269 ;
  assign n4271 = ~n4243 & ~n4270 ;
  assign n4272 = \i_tv80_core_i_reg_RegsL_reg[1][5]/NET0131  & ~n2937 ;
  assign n4273 = n2937 & ~n4269 ;
  assign n4274 = ~n4272 & ~n4273 ;
  assign n4275 = \i_tv80_core_i_reg_RegsL_reg[2][5]/NET0131  & ~n2941 ;
  assign n4276 = n2941 & ~n4269 ;
  assign n4277 = ~n4275 & ~n4276 ;
  assign n4278 = \i_tv80_core_i_reg_RegsL_reg[3][5]/NET0131  & ~n2945 ;
  assign n4279 = n2945 & ~n4269 ;
  assign n4280 = ~n4278 & ~n4279 ;
  assign n4281 = \i_tv80_core_i_reg_RegsL_reg[4][5]/NET0131  & ~n2949 ;
  assign n4282 = n2949 & ~n4269 ;
  assign n4283 = ~n4281 & ~n4282 ;
  assign n4284 = \i_tv80_core_i_reg_RegsL_reg[5][5]/NET0131  & ~n2953 ;
  assign n4285 = n2953 & ~n4269 ;
  assign n4286 = ~n4284 & ~n4285 ;
  assign n4287 = \i_tv80_core_i_reg_RegsL_reg[6][5]/NET0131  & ~n2957 ;
  assign n4288 = n2957 & ~n4269 ;
  assign n4289 = ~n4287 & ~n4288 ;
  assign n4290 = \i_tv80_core_i_reg_RegsL_reg[7][5]/NET0131  & ~n2961 ;
  assign n4291 = n2961 & ~n4269 ;
  assign n4292 = ~n4290 & ~n4291 ;
  assign n4294 = n1311 & ~n1573 ;
  assign n4295 = n1307 & ~n4294 ;
  assign n4296 = n1128 & n1451 ;
  assign n4297 = ~n4295 & ~n4296 ;
  assign n4298 = n1107 & ~n4297 ;
  assign n4300 = n862 & n1107 ;
  assign n4301 = n3849 & n4300 ;
  assign n4302 = n1308 & n1635 ;
  assign n4303 = ~n4300 & ~n4302 ;
  assign n4304 = \i_tv80_core_TmpAddr_reg[14]/P0001  & n4303 ;
  assign n4305 = ~n4301 & ~n4304 ;
  assign n4306 = ~n4298 & ~n4305 ;
  assign n4299 = \di_reg_reg[6]/P0001  & n4298 ;
  assign n4307 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4299 ;
  assign n4308 = ~n4306 & n4307 ;
  assign n4293 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[14]/P0001  ;
  assign n4309 = reset_n_pad & ~n4293 ;
  assign n4310 = ~n4308 & n4309 ;
  assign n4314 = \i_tv80_core_SP_reg[10]/P0001  & ~n3170 ;
  assign n4315 = ~n3199 & ~n3207 ;
  assign n4316 = ~n3838 & n4315 ;
  assign n4317 = n3838 & ~n4315 ;
  assign n4318 = ~n4316 & ~n4317 ;
  assign n4319 = n2699 & n4318 ;
  assign n4320 = ~n4314 & ~n4319 ;
  assign n4321 = ~n3000 & ~n4320 ;
  assign n4313 = \i_tv80_core_SP_reg[10]/P0001  & n3000 ;
  assign n4322 = ~n2997 & ~n4313 ;
  assign n4323 = ~n4321 & n4322 ;
  assign n4312 = n1945 & n2997 ;
  assign n4324 = ~n1113 & ~n4312 ;
  assign n4325 = ~n4323 & n4324 ;
  assign n4311 = \i_tv80_core_SP_reg[10]/P0001  & n1113 ;
  assign n4326 = ~n3242 & ~n4311 ;
  assign n4327 = ~n4325 & n4326 ;
  assign n4328 = n1193 & n3242 ;
  assign n4329 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4328 ;
  assign n4330 = ~n4327 & n4329 ;
  assign n4331 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[10]/P0001  ;
  assign n4332 = reset_n_pad & ~n4331 ;
  assign n4333 = ~n4330 & n4332 ;
  assign n4334 = \i_tv80_core_i_reg_RegsL_reg[0][4]/NET0131  & ~n2711 ;
  assign n4335 = ~n2808 & ~n2861 ;
  assign n4336 = ~n3463 & n4335 ;
  assign n4337 = n3463 & ~n4335 ;
  assign n4338 = ~n4336 & ~n4337 ;
  assign n4339 = n2891 & n4338 ;
  assign n4340 = \i_tv80_core_RegBusA_r_reg[4]/P0001  & n2664 ;
  assign n4341 = ~n3670 & ~n4340 ;
  assign n4342 = ~n4339 & n4341 ;
  assign n4343 = ~n2667 & ~n4342 ;
  assign n4348 = \i_tv80_core_i_reg_RegsL_reg[7][4]/NET0131  & n2904 ;
  assign n4349 = \i_tv80_core_i_reg_RegsL_reg[6][4]/NET0131  & n2920 ;
  assign n4354 = ~n4348 & ~n4349 ;
  assign n4350 = \i_tv80_core_i_reg_RegsL_reg[4][4]/NET0131  & n2918 ;
  assign n4351 = \i_tv80_core_i_reg_RegsL_reg[2][4]/NET0131  & n2908 ;
  assign n4355 = ~n4350 & ~n4351 ;
  assign n4356 = n4354 & n4355 ;
  assign n4344 = \i_tv80_core_i_reg_RegsL_reg[5][4]/NET0131  & n2916 ;
  assign n4345 = \i_tv80_core_i_reg_RegsL_reg[3][4]/NET0131  & n2922 ;
  assign n4352 = ~n4344 & ~n4345 ;
  assign n4346 = \i_tv80_core_i_reg_RegsL_reg[1][4]/NET0131  & n2914 ;
  assign n4347 = \i_tv80_core_i_reg_RegsL_reg[0][4]/NET0131  & n2911 ;
  assign n4353 = ~n4346 & ~n4347 ;
  assign n4357 = n4352 & n4353 ;
  assign n4358 = n4356 & n4357 ;
  assign n4359 = n2667 & ~n4358 ;
  assign n4360 = ~n4343 & ~n4359 ;
  assign n4361 = n2711 & ~n4360 ;
  assign n4362 = ~n4334 & ~n4361 ;
  assign n4363 = \i_tv80_core_i_reg_RegsL_reg[1][4]/NET0131  & ~n2937 ;
  assign n4364 = n2937 & ~n4360 ;
  assign n4365 = ~n4363 & ~n4364 ;
  assign n4366 = \i_tv80_core_i_reg_RegsL_reg[2][4]/NET0131  & ~n2941 ;
  assign n4367 = n2941 & ~n4360 ;
  assign n4368 = ~n4366 & ~n4367 ;
  assign n4369 = \i_tv80_core_i_reg_RegsL_reg[3][4]/NET0131  & ~n2945 ;
  assign n4370 = n2945 & ~n4360 ;
  assign n4371 = ~n4369 & ~n4370 ;
  assign n4372 = \i_tv80_core_i_reg_RegsL_reg[4][4]/NET0131  & ~n2949 ;
  assign n4373 = n2949 & ~n4360 ;
  assign n4374 = ~n4372 & ~n4373 ;
  assign n4375 = \i_tv80_core_i_reg_RegsL_reg[5][4]/NET0131  & ~n2953 ;
  assign n4376 = n2953 & ~n4360 ;
  assign n4377 = ~n4375 & ~n4376 ;
  assign n4378 = \i_tv80_core_i_reg_RegsL_reg[6][4]/NET0131  & ~n2957 ;
  assign n4379 = n2957 & ~n4360 ;
  assign n4380 = ~n4378 & ~n4379 ;
  assign n4381 = \i_tv80_core_i_reg_RegsL_reg[7][4]/NET0131  & ~n2961 ;
  assign n4382 = n2961 & ~n4360 ;
  assign n4383 = ~n4381 & ~n4382 ;
  assign n4384 = ~n879 & ~n1350 ;
  assign n4385 = n1307 & ~n4384 ;
  assign n4386 = n857 & ~n1464 ;
  assign n4387 = \i_tv80_core_IR_reg[0]/P0001  & n2654 ;
  assign n4388 = ~n4386 & ~n4387 ;
  assign n4389 = \i_tv80_core_ISet_reg[1]/P0001  & ~n4388 ;
  assign n4390 = ~n4385 & ~n4389 ;
  assign n4391 = ~\i_tv80_core_Auto_Wait_t1_reg/P0001  & ~n4390 ;
  assign n4392 = n860 & ~n930 ;
  assign n4393 = ~\i_tv80_core_Auto_Wait_t2_reg/P0001  & n4392 ;
  assign n4394 = ~n4391 & ~n4393 ;
  assign n4395 = ~wait_n_pad & n1634 ;
  assign n4396 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_BusReq_s_reg/P0001  ;
  assign n4397 = ~n4395 & ~n4396 ;
  assign n4398 = n4394 & n4397 ;
  assign n4399 = ~n1103 & n4398 ;
  assign n4403 = ~\i_tv80_core_tstate_reg[0]/P0001  & n4399 ;
  assign n4400 = \i_tv80_core_tstate_reg[0]/P0001  & ~n4399 ;
  assign n4401 = ~\i_tv80_core_BusReq_s_reg/P0001  & n1103 ;
  assign n4402 = ~n4395 & n4401 ;
  assign n4404 = ~n4400 & ~n4402 ;
  assign n4405 = ~n4403 & n4404 ;
  assign n4406 = reset_n_pad & ~n4405 ;
  assign n4407 = \i_tv80_core_BusReq_s_reg/P0001  & n1103 ;
  assign n4408 = n4397 & ~n4407 ;
  assign n4409 = \i_tv80_core_tstate_reg[1]/NET0131  & ~n4408 ;
  assign n4412 = n1106 & n4394 ;
  assign n4413 = ~n1103 & ~n4412 ;
  assign n4410 = \i_tv80_core_tstate_reg[0]/P0001  & n4394 ;
  assign n4411 = ~\i_tv80_core_tstate_reg[1]/NET0131  & ~n4410 ;
  assign n4414 = n4397 & ~n4411 ;
  assign n4415 = n4413 & n4414 ;
  assign n4416 = ~n4409 & ~n4415 ;
  assign n4417 = reset_n_pad & ~n4416 ;
  assign n4418 = ~n4407 & ~n4413 ;
  assign n4419 = ~n4395 & ~n4418 ;
  assign n4420 = ~n4396 & ~n4419 ;
  assign n4421 = \i_tv80_core_tstate_reg[2]/NET0131  & ~n4420 ;
  assign n4422 = n1107 & n4399 ;
  assign n4423 = ~n4421 & ~n4422 ;
  assign n4424 = reset_n_pad & ~n4423 ;
  assign n4426 = n2968 & ~n3591 ;
  assign n4428 = ~\i_tv80_core_BusB_reg[5]/P0001  & ~n2975 ;
  assign n4429 = ~\i_tv80_core_BusB_reg[1]/P0001  & n2975 ;
  assign n4430 = ~n4428 & ~n4429 ;
  assign n4431 = ~n2973 & ~n4430 ;
  assign n4432 = ~\i_tv80_core_BusA_reg[1]/P0001  & n2973 ;
  assign n4433 = ~n4431 & ~n4432 ;
  assign n4434 = n1157 & ~n4433 ;
  assign n4427 = ~\do[5]_pad  & ~n1157 ;
  assign n4435 = ~n2968 & ~n4427 ;
  assign n4436 = ~n4434 & n4435 ;
  assign n4437 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4436 ;
  assign n4438 = ~n4426 & n4437 ;
  assign n4425 = ~\do[5]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n4439 = reset_n_pad & ~n4425 ;
  assign n4440 = ~n4438 & n4439 ;
  assign n4443 = n1716 & n2997 ;
  assign n4445 = ~n3064 & ~n3067 ;
  assign n4446 = ~n3052 & n4445 ;
  assign n4447 = n3052 & ~n4445 ;
  assign n4448 = ~n4446 & ~n4447 ;
  assign n4449 = n3001 & n4448 ;
  assign n4444 = \i_tv80_core_SP_reg[5]/P0001  & ~n3002 ;
  assign n4450 = ~n2997 & ~n4444 ;
  assign n4451 = ~n4449 & n4450 ;
  assign n4452 = ~n4443 & ~n4451 ;
  assign n4453 = ~n1113 & ~n4452 ;
  assign n4454 = ~\i_tv80_core_SP_reg[5]/P0001  & n1113 ;
  assign n4455 = ~n4453 & ~n4454 ;
  assign n4456 = ~n2992 & ~n4455 ;
  assign n4442 = n2992 & n3591 ;
  assign n4457 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4442 ;
  assign n4458 = ~n4456 & n4457 ;
  assign n4441 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[5]/P0001  ;
  assign n4459 = reset_n_pad & ~n4441 ;
  assign n4460 = ~n4458 & n4459 ;
  assign n4464 = ~n3217 & ~n3223 ;
  assign n4465 = ~n3838 & n3839 ;
  assign n4466 = n3843 & ~n4465 ;
  assign n4467 = n4464 & ~n4466 ;
  assign n4468 = ~n4464 & n4466 ;
  assign n4469 = ~n4467 & ~n4468 ;
  assign n4470 = n3001 & n4469 ;
  assign n4463 = \i_tv80_core_SP_reg[12]/P0001  & ~n3002 ;
  assign n4471 = ~n2997 & ~n4463 ;
  assign n4472 = ~n4470 & n4471 ;
  assign n4462 = n2079 & n2997 ;
  assign n4473 = ~n1113 & ~n4462 ;
  assign n4474 = ~n4472 & n4473 ;
  assign n4461 = \i_tv80_core_SP_reg[12]/P0001  & n1113 ;
  assign n4475 = ~n3242 & ~n4461 ;
  assign n4476 = ~n4474 & n4475 ;
  assign n4477 = n3242 & n3669 ;
  assign n4478 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4477 ;
  assign n4479 = ~n4476 & n4478 ;
  assign n4480 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[12]/P0001  ;
  assign n4481 = reset_n_pad & ~n4480 ;
  assign n4482 = ~n4479 & n4481 ;
  assign n4485 = \i_tv80_core_SP_reg[13]/P0001  & ~n3170 ;
  assign n4486 = ~n3181 & ~n3221 ;
  assign n4487 = ~n3219 & n3224 ;
  assign n4488 = n4486 & ~n4487 ;
  assign n4489 = ~n4486 & n4487 ;
  assign n4490 = ~n4488 & ~n4489 ;
  assign n4491 = n2699 & n4490 ;
  assign n4492 = ~n4485 & ~n4491 ;
  assign n4493 = ~n3000 & ~n4492 ;
  assign n4484 = \i_tv80_core_SP_reg[13]/P0001  & n3000 ;
  assign n4494 = ~n2997 & ~n4484 ;
  assign n4495 = ~n4493 & n4494 ;
  assign n4483 = n2142 & n2997 ;
  assign n4496 = ~n1113 & ~n4483 ;
  assign n4497 = ~n4495 & n4496 ;
  assign n4498 = \i_tv80_core_SP_reg[13]/P0001  & n1113 ;
  assign n4499 = ~n3242 & ~n4498 ;
  assign n4500 = ~n4497 & n4499 ;
  assign n4501 = n3242 & n3591 ;
  assign n4502 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4501 ;
  assign n4503 = ~n4500 & n4502 ;
  assign n4504 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[13]/P0001  ;
  assign n4505 = reset_n_pad & ~n4504 ;
  assign n4506 = ~n4503 & n4505 ;
  assign n4507 = \i_tv80_core_i_reg_RegsL_reg[0][3]/NET0131  & ~n2711 ;
  assign n4508 = ~n2841 & ~n2862 ;
  assign n4509 = ~n2792 & n4508 ;
  assign n4510 = n2792 & ~n4508 ;
  assign n4511 = ~n4509 & ~n4510 ;
  assign n4512 = n2891 & n4511 ;
  assign n4513 = \i_tv80_core_RegBusA_r_reg[3]/P0001  & n2664 ;
  assign n4514 = ~n4017 & ~n4513 ;
  assign n4515 = ~n4512 & n4514 ;
  assign n4516 = ~n2667 & ~n4515 ;
  assign n4521 = \i_tv80_core_i_reg_RegsL_reg[3][3]/NET0131  & n2922 ;
  assign n4522 = \i_tv80_core_i_reg_RegsL_reg[2][3]/NET0131  & n2908 ;
  assign n4527 = ~n4521 & ~n4522 ;
  assign n4523 = \i_tv80_core_i_reg_RegsL_reg[4][3]/NET0131  & n2918 ;
  assign n4524 = \i_tv80_core_i_reg_RegsL_reg[0][3]/NET0131  & n2911 ;
  assign n4528 = ~n4523 & ~n4524 ;
  assign n4529 = n4527 & n4528 ;
  assign n4517 = \i_tv80_core_i_reg_RegsL_reg[5][3]/NET0131  & n2916 ;
  assign n4518 = \i_tv80_core_i_reg_RegsL_reg[1][3]/NET0131  & n2914 ;
  assign n4525 = ~n4517 & ~n4518 ;
  assign n4519 = \i_tv80_core_i_reg_RegsL_reg[7][3]/NET0131  & n2904 ;
  assign n4520 = \i_tv80_core_i_reg_RegsL_reg[6][3]/NET0131  & n2920 ;
  assign n4526 = ~n4519 & ~n4520 ;
  assign n4530 = n4525 & n4526 ;
  assign n4531 = n4529 & n4530 ;
  assign n4532 = n2667 & ~n4531 ;
  assign n4533 = ~n4516 & ~n4532 ;
  assign n4534 = n2711 & ~n4533 ;
  assign n4535 = ~n4507 & ~n4534 ;
  assign n4536 = \i_tv80_core_i_reg_RegsL_reg[1][3]/NET0131  & ~n2937 ;
  assign n4537 = n2937 & ~n4533 ;
  assign n4538 = ~n4536 & ~n4537 ;
  assign n4539 = \i_tv80_core_i_reg_RegsL_reg[2][3]/NET0131  & ~n2941 ;
  assign n4540 = n2941 & ~n4533 ;
  assign n4541 = ~n4539 & ~n4540 ;
  assign n4542 = \i_tv80_core_i_reg_RegsL_reg[3][3]/NET0131  & ~n2945 ;
  assign n4543 = n2945 & ~n4533 ;
  assign n4544 = ~n4542 & ~n4543 ;
  assign n4545 = \i_tv80_core_i_reg_RegsL_reg[4][3]/NET0131  & ~n2949 ;
  assign n4546 = n2949 & ~n4533 ;
  assign n4547 = ~n4545 & ~n4546 ;
  assign n4548 = \i_tv80_core_i_reg_RegsL_reg[5][3]/NET0131  & ~n2953 ;
  assign n4549 = n2953 & ~n4533 ;
  assign n4550 = ~n4548 & ~n4549 ;
  assign n4551 = \i_tv80_core_i_reg_RegsL_reg[6][3]/NET0131  & ~n2957 ;
  assign n4552 = n2957 & ~n4533 ;
  assign n4553 = ~n4551 & ~n4552 ;
  assign n4554 = \i_tv80_core_i_reg_RegsL_reg[7][3]/NET0131  & ~n2961 ;
  assign n4555 = n2961 & ~n4533 ;
  assign n4556 = ~n4554 & ~n4555 ;
  assign n4558 = n2968 & ~n3669 ;
  assign n4560 = ~\i_tv80_core_BusB_reg[4]/P0001  & ~n2975 ;
  assign n4561 = ~\i_tv80_core_BusB_reg[0]/P0001  & n2975 ;
  assign n4562 = ~n4560 & ~n4561 ;
  assign n4563 = ~n2973 & ~n4562 ;
  assign n4564 = ~\i_tv80_core_BusA_reg[0]/P0001  & n2973 ;
  assign n4565 = ~n4563 & ~n4564 ;
  assign n4566 = n1157 & ~n4565 ;
  assign n4559 = ~\do[4]_pad  & ~n1157 ;
  assign n4567 = ~n2968 & ~n4559 ;
  assign n4568 = ~n4566 & n4567 ;
  assign n4569 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4568 ;
  assign n4570 = ~n4558 & n4569 ;
  assign n4557 = ~\do[4]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n4571 = reset_n_pad & ~n4557 ;
  assign n4572 = ~n4570 & n4571 ;
  assign n4575 = n2389 & n2997 ;
  assign n4577 = ~n3018 & ~n3019 ;
  assign n4578 = n3050 & ~n4577 ;
  assign n4579 = ~n3050 & n4577 ;
  assign n4580 = ~n4578 & ~n4579 ;
  assign n4581 = n3001 & n4580 ;
  assign n4576 = \i_tv80_core_SP_reg[4]/P0001  & ~n3002 ;
  assign n4582 = ~n2997 & ~n4576 ;
  assign n4583 = ~n4581 & n4582 ;
  assign n4584 = ~n4575 & ~n4583 ;
  assign n4585 = ~n1113 & ~n4584 ;
  assign n4586 = ~\i_tv80_core_SP_reg[4]/P0001  & n1113 ;
  assign n4587 = ~n4585 & ~n4586 ;
  assign n4588 = ~n2992 & ~n4587 ;
  assign n4574 = n2992 & n3669 ;
  assign n4589 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4574 ;
  assign n4590 = ~n4588 & n4589 ;
  assign n4573 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[4]/P0001  ;
  assign n4591 = reset_n_pad & ~n4573 ;
  assign n4592 = ~n4590 & n4591 ;
  assign n4594 = ~n862 & ~n1462 ;
  assign n4595 = n1430 & ~n1462 ;
  assign n4596 = ~n4594 & ~n4595 ;
  assign n4597 = \i_tv80_core_IncDecZ_reg/P0002  & \i_tv80_core_mcycle_reg[1]/P0001  ;
  assign n4598 = n384 & n4597 ;
  assign n4599 = ~\i_tv80_core_No_BTR_reg/P0001  & ~n1330 ;
  assign n4600 = ~n4598 & n4599 ;
  assign n4601 = ~n4596 & n4600 ;
  assign n4602 = \i_tv80_core_mcycle_reg[0]/P0001  & n4601 ;
  assign n4603 = \i_tv80_core_Pre_XY_F_M_reg[0]/P0001  & n4596 ;
  assign n4604 = ~n4602 & ~n4603 ;
  assign n4605 = ~n1599 & n4604 ;
  assign n4606 = n4402 & n4605 ;
  assign n4593 = \i_tv80_core_mcycle_reg[0]/P0001  & ~n4402 ;
  assign n4607 = reset_n_pad & ~n4593 ;
  assign n4608 = ~n4606 & n4607 ;
  assign n4610 = n1167 & ~n3669 ;
  assign n4612 = ~\i_tv80_core_F_reg[4]/P0001  & ~n4188 ;
  assign n4613 = ~n3128 & ~n4612 ;
  assign n4614 = ~n1117 & ~n4613 ;
  assign n4611 = ~\i_tv80_core_Fp_reg[4]/P0001  & n1117 ;
  assign n4615 = n4149 & ~n4611 ;
  assign n4616 = ~n4614 & n4615 ;
  assign n4624 = n458 & n3111 ;
  assign n4623 = ~n458 & n696 ;
  assign n4625 = ~n518 & ~n4623 ;
  assign n4626 = ~n4624 & n4625 ;
  assign n4627 = ~\i_tv80_core_ALU_Op_r_reg[3]/P0001  & ~n4626 ;
  assign n4619 = \i_tv80_core_F_reg[1]/P0001  & ~n781 ;
  assign n4620 = n735 & ~n816 ;
  assign n4621 = ~n4619 & n4620 ;
  assign n4622 = \i_tv80_core_F_reg[4]/P0001  & n697 ;
  assign n4628 = ~n4621 & ~n4622 ;
  assign n4629 = ~n4627 & n4628 ;
  assign n4630 = n385 & ~n4629 ;
  assign n4617 = \i_tv80_core_F_reg[4]/P0001  & n1113 ;
  assign n4618 = ~n385 & n4617 ;
  assign n4631 = ~n370 & ~n4618 ;
  assign n4632 = ~n4630 & n4631 ;
  assign n4633 = ~n4616 & n4632 ;
  assign n4634 = n4167 & ~n4633 ;
  assign n4635 = ~n4610 & ~n4634 ;
  assign n4636 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4635 ;
  assign n4609 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_F_reg[4]/P0001  ;
  assign n4637 = reset_n_pad & ~n4609 ;
  assign n4638 = ~n4636 & n4637 ;
  assign n4639 = \i_tv80_core_mcycle_reg[1]/P0001  & reset_n_pad ;
  assign n4640 = ~n4402 & n4639 ;
  assign n4641 = \i_tv80_core_Pre_XY_F_M_reg[0]/P0001  & \i_tv80_core_Pre_XY_F_M_reg[1]/P0001  ;
  assign n4642 = ~\i_tv80_core_Pre_XY_F_M_reg[0]/P0001  & ~\i_tv80_core_Pre_XY_F_M_reg[1]/P0001  ;
  assign n4643 = ~n4641 & ~n4642 ;
  assign n4644 = n4596 & n4643 ;
  assign n4645 = n380 & n4601 ;
  assign n4646 = ~n4644 & ~n4645 ;
  assign n4647 = ~n1599 & n4646 ;
  assign n4648 = reset_n_pad & ~n4396 ;
  assign n4649 = n4402 & n4648 ;
  assign n4650 = ~n4647 & n4649 ;
  assign n4651 = ~n4640 & ~n4650 ;
  assign n4659 = ~n378 & ~n1599 ;
  assign n4660 = n4402 & ~n4659 ;
  assign n4661 = ~\i_tv80_core_mcycle_reg[2]/P0001  & ~n4660 ;
  assign n4652 = \i_tv80_core_Pre_XY_F_M_reg[2]/P0001  & ~n4641 ;
  assign n4653 = ~\i_tv80_core_Pre_XY_F_M_reg[2]/P0001  & n4641 ;
  assign n4654 = ~n4652 & ~n4653 ;
  assign n4655 = n4596 & ~n4654 ;
  assign n4656 = ~n4601 & ~n4655 ;
  assign n4657 = ~n1599 & n4656 ;
  assign n4658 = n4402 & n4657 ;
  assign n4662 = reset_n_pad & ~n4658 ;
  assign n4663 = ~n4661 & n4662 ;
  assign n4664 = \i_tv80_core_i_reg_RegsL_reg[0][2]/P0001  & ~n2711 ;
  assign n4665 = ~n2771 & ~n2773 ;
  assign n4666 = ~n3459 & ~n4665 ;
  assign n4667 = n3459 & n4665 ;
  assign n4668 = ~n4666 & ~n4667 ;
  assign n4669 = n2891 & ~n4668 ;
  assign n4670 = \i_tv80_core_RegBusA_r_reg[2]/P0001  & n2664 ;
  assign n4671 = ~n3872 & ~n4670 ;
  assign n4672 = ~n4669 & n4671 ;
  assign n4673 = ~n2667 & ~n4672 ;
  assign n4678 = \i_tv80_core_i_reg_RegsL_reg[4][2]/P0001  & n2918 ;
  assign n4679 = \i_tv80_core_i_reg_RegsL_reg[5][2]/P0001  & n2916 ;
  assign n4684 = ~n4678 & ~n4679 ;
  assign n4680 = \i_tv80_core_i_reg_RegsL_reg[7][2]/P0001  & n2904 ;
  assign n4681 = \i_tv80_core_i_reg_RegsL_reg[2][2]/P0001  & n2908 ;
  assign n4685 = ~n4680 & ~n4681 ;
  assign n4686 = n4684 & n4685 ;
  assign n4674 = \i_tv80_core_i_reg_RegsL_reg[6][2]/P0001  & n2920 ;
  assign n4675 = \i_tv80_core_i_reg_RegsL_reg[3][2]/P0001  & n2922 ;
  assign n4682 = ~n4674 & ~n4675 ;
  assign n4676 = \i_tv80_core_i_reg_RegsL_reg[1][2]/P0001  & n2914 ;
  assign n4677 = \i_tv80_core_i_reg_RegsL_reg[0][2]/P0001  & n2911 ;
  assign n4683 = ~n4676 & ~n4677 ;
  assign n4687 = n4682 & n4683 ;
  assign n4688 = n4686 & n4687 ;
  assign n4689 = n2667 & ~n4688 ;
  assign n4690 = ~n4673 & ~n4689 ;
  assign n4691 = n2711 & ~n4690 ;
  assign n4692 = ~n4664 & ~n4691 ;
  assign n4693 = \i_tv80_core_i_reg_RegsL_reg[1][2]/P0001  & ~n2937 ;
  assign n4694 = n2937 & ~n4690 ;
  assign n4695 = ~n4693 & ~n4694 ;
  assign n4696 = \i_tv80_core_i_reg_RegsL_reg[2][2]/P0001  & ~n2941 ;
  assign n4697 = n2941 & ~n4690 ;
  assign n4698 = ~n4696 & ~n4697 ;
  assign n4699 = \i_tv80_core_i_reg_RegsL_reg[3][2]/P0001  & ~n2945 ;
  assign n4700 = n2945 & ~n4690 ;
  assign n4701 = ~n4699 & ~n4700 ;
  assign n4702 = \i_tv80_core_i_reg_RegsL_reg[4][2]/P0001  & ~n2949 ;
  assign n4703 = n2949 & ~n4690 ;
  assign n4704 = ~n4702 & ~n4703 ;
  assign n4705 = \i_tv80_core_i_reg_RegsL_reg[5][2]/P0001  & ~n2953 ;
  assign n4706 = n2953 & ~n4690 ;
  assign n4707 = ~n4705 & ~n4706 ;
  assign n4708 = \i_tv80_core_i_reg_RegsL_reg[6][2]/P0001  & ~n2957 ;
  assign n4709 = n2957 & ~n4690 ;
  assign n4710 = ~n4708 & ~n4709 ;
  assign n4711 = \i_tv80_core_i_reg_RegsL_reg[7][2]/P0001  & ~n2961 ;
  assign n4712 = n2961 & ~n4690 ;
  assign n4713 = ~n4711 & ~n4712 ;
  assign n4714 = ~n4596 & ~n4600 ;
  assign n4715 = ~n1599 & n4714 ;
  assign n4716 = n4401 & n4715 ;
  assign n4717 = \i_tv80_core_IntCycle_reg/P0001  & ~n4716 ;
  assign n4722 = n382 & n1334 ;
  assign n4723 = n869 & n3152 ;
  assign n4724 = ~n628 & n4723 ;
  assign n4725 = ~n4722 & ~n4724 ;
  assign n4726 = n4716 & n4725 ;
  assign n4718 = \i_tv80_core_IR_reg[3]/P0001  & n2994 ;
  assign n4719 = n1066 & n4718 ;
  assign n4720 = \i_tv80_core_INT_s_reg/P0001  & \i_tv80_core_IntE_FF1_reg/P0001  ;
  assign n4721 = ~n4719 & n4720 ;
  assign n4727 = ~\i_tv80_core_NMI_s_reg/P0001  & n4721 ;
  assign n4728 = n4726 & n4727 ;
  assign n4729 = ~n4717 & ~n4728 ;
  assign n4730 = reset_n_pad & ~n4729 ;
  assign n4731 = n1634 & n4719 ;
  assign n4732 = ~\i_tv80_core_IntE_FF2_reg/P0001  & ~n4731 ;
  assign n4733 = n1067 & n2666 ;
  assign n4734 = reset_n_pad & ~n4733 ;
  assign n4735 = ~n4732 & n4734 ;
  assign n4736 = ~n4728 & n4735 ;
  assign n4738 = n886 & n989 ;
  assign n4739 = n382 & n673 ;
  assign n4740 = n4738 & n4739 ;
  assign n4741 = ~\i_tv80_core_Halt_FF_reg/P0001  & n930 ;
  assign n4742 = ~n4740 & n4741 ;
  assign n4743 = ~n1313 & n4742 ;
  assign n4744 = n1625 & n4743 ;
  assign n4745 = n1635 & n4744 ;
  assign n4747 = ~n1338 & ~n1339 ;
  assign n4748 = ~n1374 & n4747 ;
  assign n4749 = ~n1371 & n1408 ;
  assign n4750 = n4748 & n4749 ;
  assign n4751 = n956 & ~n4750 ;
  assign n4752 = n382 & n4751 ;
  assign n4753 = \i_tv80_core_BTR_r_reg/P0001  & ~n4752 ;
  assign n4754 = ~\di_reg_reg[0]/P0001  & n4752 ;
  assign n4755 = ~n4753 & ~n4754 ;
  assign n4756 = ~\i_tv80_core_PC_reg[0]/P0001  & ~n4755 ;
  assign n4757 = \i_tv80_core_PC_reg[0]/P0001  & n4755 ;
  assign n4758 = ~n4756 & ~n4757 ;
  assign n4759 = n4745 & n4758 ;
  assign n4746 = \i_tv80_core_PC_reg[0]/P0001  & ~n4745 ;
  assign n4760 = n1113 & ~n4746 ;
  assign n4761 = ~n4759 & n4760 ;
  assign n4795 = \i_tv80_core_PC_reg[0]/P0001  & ~n1317 ;
  assign n4796 = ~n1887 & ~n4795 ;
  assign n4797 = n1886 & ~n4796 ;
  assign n4798 = ~n1885 & ~n4797 ;
  assign n4799 = ~n1277 & ~n4798 ;
  assign n4800 = ~n1884 & ~n4799 ;
  assign n4801 = n1625 & ~n4800 ;
  assign n4802 = n1915 & ~n4801 ;
  assign n4762 = ~n879 & ~n1335 ;
  assign n4763 = n4750 & n4762 ;
  assign n4764 = ~\i_tv80_core_mcycle_reg[0]/P0001  & ~n4763 ;
  assign n4766 = ~n910 & ~n974 ;
  assign n4767 = n899 & n4766 ;
  assign n4765 = ~n871 & ~n1356 ;
  assign n4768 = n1484 & n4765 ;
  assign n4769 = n4767 & n4768 ;
  assign n4770 = ~n4764 & n4769 ;
  assign n4771 = n856 & ~n4770 ;
  assign n4775 = n856 & n1348 ;
  assign n4776 = n857 & n1353 ;
  assign n4777 = \i_tv80_core_IR_reg[6]/P0001  & n4776 ;
  assign n4778 = ~n4775 & ~n4777 ;
  assign n4779 = n1481 & n1617 ;
  assign n4772 = n857 & n1350 ;
  assign n4773 = n857 & n1069 ;
  assign n4774 = ~\i_tv80_core_IR_reg[6]/P0001  & n4773 ;
  assign n4780 = ~n4772 & ~n4774 ;
  assign n4781 = ~n4779 & n4780 ;
  assign n4782 = n4778 & n4781 ;
  assign n4783 = ~n4751 & n4782 ;
  assign n4784 = ~n4771 & n4783 ;
  assign n4785 = n382 & ~n4784 ;
  assign n4787 = ~n1335 & ~n1430 ;
  assign n4788 = n1462 & ~n4787 ;
  assign n4786 = n856 & n1576 ;
  assign n4789 = ~\i_tv80_core_BTR_r_reg/P0001  & ~n862 ;
  assign n4790 = ~n4786 & n4789 ;
  assign n4791 = ~n4788 & n4790 ;
  assign n4792 = ~n4785 & n4791 ;
  assign n4793 = n1635 & ~n4792 ;
  assign n4803 = ~\i_tv80_core_PC_reg[0]/P0001  & ~n1103 ;
  assign n4804 = ~n4793 & ~n4803 ;
  assign n4805 = ~n4802 & n4804 ;
  assign n4794 = n4758 & n4793 ;
  assign n4806 = ~n1113 & ~n4794 ;
  assign n4807 = ~n4805 & n4806 ;
  assign n4808 = ~n4761 & ~n4807 ;
  assign n4809 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4808 ;
  assign n4737 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PC_reg[0]/P0001  ;
  assign n4810 = reset_n_pad & ~n4737 ;
  assign n4811 = ~n4809 & n4810 ;
  assign n4813 = \di_reg_reg[7]/P0001  & n4752 ;
  assign n4814 = ~n4753 & ~n4813 ;
  assign n4815 = \i_tv80_core_PC_reg[10]/P0001  & ~n4814 ;
  assign n4816 = ~\i_tv80_core_PC_reg[10]/P0001  & n4814 ;
  assign n4817 = ~n4815 & ~n4816 ;
  assign n4823 = \i_tv80_core_PC_reg[7]/P0001  & ~n4814 ;
  assign n4824 = \di_reg_reg[6]/P0001  & n4752 ;
  assign n4825 = ~n4753 & ~n4824 ;
  assign n4826 = ~\i_tv80_core_PC_reg[6]/P0001  & n4825 ;
  assign n4827 = \i_tv80_core_PC_reg[6]/P0001  & ~n4825 ;
  assign n4828 = \di_reg_reg[5]/P0001  & n4752 ;
  assign n4829 = ~n4753 & ~n4828 ;
  assign n4830 = ~\i_tv80_core_PC_reg[5]/P0001  & n4829 ;
  assign n4831 = \i_tv80_core_PC_reg[5]/P0001  & ~n4829 ;
  assign n4832 = \di_reg_reg[4]/P0001  & n4752 ;
  assign n4833 = ~n4753 & ~n4832 ;
  assign n4834 = ~\i_tv80_core_PC_reg[4]/P0001  & n4833 ;
  assign n4835 = \i_tv80_core_PC_reg[4]/P0001  & ~n4833 ;
  assign n4836 = \di_reg_reg[3]/P0001  & n4752 ;
  assign n4837 = ~n4753 & ~n4836 ;
  assign n4838 = ~\i_tv80_core_PC_reg[3]/P0001  & n4837 ;
  assign n4839 = \i_tv80_core_PC_reg[3]/P0001  & ~n4837 ;
  assign n4840 = \di_reg_reg[2]/P0001  & n4752 ;
  assign n4841 = ~n4753 & ~n4840 ;
  assign n4842 = ~\i_tv80_core_PC_reg[2]/P0001  & n4841 ;
  assign n4843 = \i_tv80_core_PC_reg[2]/P0001  & ~n4841 ;
  assign n4844 = \di_reg_reg[1]/P0001  & n4752 ;
  assign n4845 = ~n4753 & ~n4844 ;
  assign n4846 = ~\i_tv80_core_PC_reg[1]/P0001  & n4845 ;
  assign n4847 = \i_tv80_core_PC_reg[1]/P0001  & ~n4845 ;
  assign n4848 = ~n4757 & ~n4847 ;
  assign n4849 = ~n4846 & ~n4848 ;
  assign n4850 = ~n4843 & ~n4849 ;
  assign n4851 = ~n4842 & ~n4850 ;
  assign n4852 = ~n4839 & ~n4851 ;
  assign n4853 = ~n4838 & ~n4852 ;
  assign n4854 = ~n4835 & ~n4853 ;
  assign n4855 = ~n4834 & ~n4854 ;
  assign n4856 = ~n4831 & ~n4855 ;
  assign n4857 = ~n4830 & ~n4856 ;
  assign n4858 = ~n4827 & ~n4857 ;
  assign n4859 = ~n4826 & ~n4858 ;
  assign n4860 = ~n4823 & ~n4859 ;
  assign n4820 = ~\i_tv80_core_PC_reg[8]/P0001  & n4814 ;
  assign n4821 = ~\i_tv80_core_PC_reg[7]/P0001  & n4814 ;
  assign n4822 = ~n4820 & ~n4821 ;
  assign n4861 = ~\i_tv80_core_PC_reg[9]/P0001  & n4814 ;
  assign n4862 = n4822 & ~n4861 ;
  assign n4863 = ~n4860 & n4862 ;
  assign n4818 = \i_tv80_core_PC_reg[8]/P0001  & ~n4814 ;
  assign n4819 = \i_tv80_core_PC_reg[9]/P0001  & ~n4814 ;
  assign n4864 = ~n4818 & ~n4819 ;
  assign n4865 = ~n4863 & n4864 ;
  assign n4866 = n4817 & n4865 ;
  assign n4867 = ~n4817 & ~n4865 ;
  assign n4868 = ~n4866 & ~n4867 ;
  assign n4873 = n4793 & n4868 ;
  assign n4883 = \i_tv80_core_PC_reg[10]/P0001  & ~n1103 ;
  assign n4874 = \i_tv80_core_PC_reg[10]/P0001  & ~n1317 ;
  assign n4875 = ~n1929 & ~n4874 ;
  assign n4876 = n1886 & ~n4875 ;
  assign n4877 = ~n1979 & ~n4876 ;
  assign n4878 = ~n1277 & ~n4877 ;
  assign n4879 = ~n1982 & ~n4878 ;
  assign n4880 = n1625 & ~n4879 ;
  assign n4881 = ~n1985 & ~n4880 ;
  assign n4882 = n1103 & ~n4881 ;
  assign n4884 = ~n4793 & ~n4882 ;
  assign n4885 = ~n4883 & n4884 ;
  assign n4886 = ~n1113 & ~n4885 ;
  assign n4887 = ~n4873 & n4886 ;
  assign n4869 = n4745 & n4868 ;
  assign n4870 = ~\i_tv80_core_PC_reg[10]/P0001  & ~n4745 ;
  assign n4871 = n1113 & ~n4870 ;
  assign n4872 = ~n4869 & n4871 ;
  assign n4888 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4872 ;
  assign n4889 = ~n4887 & n4888 ;
  assign n4812 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PC_reg[10]/P0001  ;
  assign n4890 = reset_n_pad & ~n4812 ;
  assign n4891 = ~n4889 & n4890 ;
  assign n4893 = ~\i_tv80_core_PC_reg[11]/P0001  & n4814 ;
  assign n4894 = \i_tv80_core_PC_reg[11]/P0001  & ~n4814 ;
  assign n4895 = ~n4893 & ~n4894 ;
  assign n4896 = n4822 & n4859 ;
  assign n4897 = ~n4818 & ~n4823 ;
  assign n4898 = ~n4896 & n4897 ;
  assign n4899 = ~n4816 & ~n4861 ;
  assign n4900 = ~n4898 & n4899 ;
  assign n4901 = ~n4815 & ~n4819 ;
  assign n4902 = ~n4900 & n4901 ;
  assign n4903 = n4895 & ~n4902 ;
  assign n4904 = ~n4895 & n4902 ;
  assign n4905 = ~n4903 & ~n4904 ;
  assign n4910 = n4793 & ~n4905 ;
  assign n4920 = \i_tv80_core_PC_reg[11]/P0001  & ~n1103 ;
  assign n4911 = \i_tv80_core_PC_reg[11]/P0001  & ~n1317 ;
  assign n4912 = ~n2000 & ~n4911 ;
  assign n4913 = n1886 & ~n4912 ;
  assign n4914 = ~n2042 & ~n4913 ;
  assign n4915 = ~n1277 & ~n4914 ;
  assign n4916 = ~n2045 & ~n4915 ;
  assign n4917 = n1625 & ~n4916 ;
  assign n4918 = ~n2048 & ~n4917 ;
  assign n4919 = n1103 & ~n4918 ;
  assign n4921 = ~n4793 & ~n4919 ;
  assign n4922 = ~n4920 & n4921 ;
  assign n4923 = ~n1113 & ~n4922 ;
  assign n4924 = ~n4910 & n4923 ;
  assign n4906 = n4745 & ~n4905 ;
  assign n4907 = ~\i_tv80_core_PC_reg[11]/P0001  & ~n4745 ;
  assign n4908 = n1113 & ~n4907 ;
  assign n4909 = ~n4906 & n4908 ;
  assign n4925 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4909 ;
  assign n4926 = ~n4924 & n4925 ;
  assign n4892 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PC_reg[11]/P0001  ;
  assign n4927 = reset_n_pad & ~n4892 ;
  assign n4928 = ~n4926 & n4927 ;
  assign n4930 = \i_tv80_core_PC_reg[12]/P0001  & ~n4814 ;
  assign n4931 = ~\i_tv80_core_PC_reg[12]/P0001  & n4814 ;
  assign n4932 = ~n4930 & ~n4931 ;
  assign n4933 = ~n4815 & ~n4894 ;
  assign n4934 = ~n4816 & ~n4893 ;
  assign n4935 = ~n4865 & n4934 ;
  assign n4936 = n4933 & ~n4935 ;
  assign n4937 = n4932 & ~n4936 ;
  assign n4938 = ~n4932 & n4936 ;
  assign n4939 = ~n4937 & ~n4938 ;
  assign n4944 = n4793 & ~n4939 ;
  assign n4954 = \i_tv80_core_PC_reg[12]/P0001  & ~n1103 ;
  assign n4945 = \i_tv80_core_PC_reg[12]/P0001  & ~n1317 ;
  assign n4946 = ~n2063 & ~n4945 ;
  assign n4947 = n1886 & ~n4946 ;
  assign n4948 = ~n2105 & ~n4947 ;
  assign n4949 = ~n1277 & ~n4948 ;
  assign n4950 = ~n2108 & ~n4949 ;
  assign n4951 = n1625 & ~n4950 ;
  assign n4952 = ~n2111 & ~n4951 ;
  assign n4953 = n1103 & ~n4952 ;
  assign n4955 = ~n4793 & ~n4953 ;
  assign n4956 = ~n4954 & n4955 ;
  assign n4957 = ~n1113 & ~n4956 ;
  assign n4958 = ~n4944 & n4957 ;
  assign n4940 = n4745 & ~n4939 ;
  assign n4941 = ~\i_tv80_core_PC_reg[12]/P0001  & ~n4745 ;
  assign n4942 = n1113 & ~n4941 ;
  assign n4943 = ~n4940 & n4942 ;
  assign n4959 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4943 ;
  assign n4960 = ~n4958 & n4959 ;
  assign n4929 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PC_reg[12]/P0001  ;
  assign n4961 = reset_n_pad & ~n4929 ;
  assign n4962 = ~n4960 & n4961 ;
  assign n4966 = \i_tv80_core_PC_reg[13]/P0001  & ~n4814 ;
  assign n4967 = ~\i_tv80_core_PC_reg[13]/P0001  & n4814 ;
  assign n4968 = ~n4966 & ~n4967 ;
  assign n4969 = ~n4893 & ~n4931 ;
  assign n4970 = ~n4902 & n4969 ;
  assign n4971 = ~n4894 & ~n4930 ;
  assign n4972 = ~n4970 & n4971 ;
  assign n4973 = n4968 & ~n4972 ;
  assign n4974 = ~n4968 & n4972 ;
  assign n4975 = ~n4973 & ~n4974 ;
  assign n4976 = n4745 & ~n4975 ;
  assign n4965 = ~\i_tv80_core_PC_reg[13]/P0001  & ~n4745 ;
  assign n4977 = ~\i_tv80_core_BusAck_reg/P0001  & ~n4965 ;
  assign n4978 = ~n4976 & n4977 ;
  assign n4963 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_PC_reg[13]/P0001  ;
  assign n4964 = ~\i_tv80_core_BusAck_reg/P0001  & ~n1113 ;
  assign n4979 = ~n4963 & ~n4964 ;
  assign n4980 = ~n4978 & n4979 ;
  assign n4981 = n4793 & n4975 ;
  assign n4982 = \i_tv80_core_PC_reg[13]/P0001  & ~n1317 ;
  assign n4983 = ~n2126 & ~n4982 ;
  assign n4984 = n1886 & ~n4983 ;
  assign n4985 = ~n2168 & ~n4984 ;
  assign n4986 = ~n1277 & ~n4985 ;
  assign n4987 = ~n2171 & ~n4986 ;
  assign n4988 = n1625 & ~n4987 ;
  assign n4989 = n2175 & ~n4988 ;
  assign n4990 = ~\i_tv80_core_PC_reg[13]/P0001  & ~n1103 ;
  assign n4991 = ~n4793 & ~n4990 ;
  assign n4992 = ~n4989 & n4991 ;
  assign n4993 = n4964 & ~n4992 ;
  assign n4994 = ~n4981 & n4993 ;
  assign n4995 = reset_n_pad & ~n4994 ;
  assign n4996 = ~n4980 & n4995 ;
  assign n4997 = \i_tv80_core_PC_reg[14]/P0001  & ~n4814 ;
  assign n4998 = ~\i_tv80_core_PC_reg[14]/P0001  & n4814 ;
  assign n4999 = ~n4997 & ~n4998 ;
  assign n5000 = n4935 & ~n4967 ;
  assign n5001 = n4933 & ~n4966 ;
  assign n5002 = ~n5000 & n5001 ;
  assign n5003 = ~n4931 & ~n5002 ;
  assign n5004 = ~n4930 & ~n5003 ;
  assign n5005 = n4999 & n5004 ;
  assign n5006 = ~n4999 & ~n5004 ;
  assign n5007 = ~n5005 & ~n5006 ;
  assign n5024 = n4745 & n5007 ;
  assign n5023 = ~\i_tv80_core_PC_reg[14]/P0001  & ~n4745 ;
  assign n5025 = n1113 & ~n5023 ;
  assign n5026 = ~n5024 & n5025 ;
  assign n5008 = n4793 & n5007 ;
  assign n5018 = \i_tv80_core_PC_reg[14]/P0001  & ~n1103 ;
  assign n5009 = \i_tv80_core_PC_reg[14]/P0001  & ~n1317 ;
  assign n5010 = ~n2189 & ~n5009 ;
  assign n5011 = n1886 & ~n5010 ;
  assign n5012 = ~n2231 & ~n5011 ;
  assign n5013 = ~n1277 & ~n5012 ;
  assign n5014 = ~n2234 & ~n5013 ;
  assign n5015 = n1625 & ~n5014 ;
  assign n5016 = ~n2237 & ~n5015 ;
  assign n5017 = n1103 & ~n5016 ;
  assign n5019 = ~n4793 & ~n5017 ;
  assign n5020 = ~n5018 & n5019 ;
  assign n5021 = ~n1113 & ~n5020 ;
  assign n5022 = ~n5008 & n5021 ;
  assign n5027 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5022 ;
  assign n5028 = ~n5026 & n5027 ;
  assign n5029 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PC_reg[14]/P0001  ;
  assign n5030 = reset_n_pad & ~n5029 ;
  assign n5031 = ~n5028 & n5030 ;
  assign n5032 = ~n4967 & ~n4998 ;
  assign n5033 = ~n4972 & n5032 ;
  assign n5034 = ~n4966 & ~n4997 ;
  assign n5035 = ~n5033 & n5034 ;
  assign n5036 = \i_tv80_core_PC_reg[15]/P0001  & ~n4814 ;
  assign n5037 = ~\i_tv80_core_PC_reg[15]/P0001  & n4814 ;
  assign n5038 = ~n5036 & ~n5037 ;
  assign n5039 = n5035 & n5038 ;
  assign n5040 = ~n5035 & ~n5038 ;
  assign n5041 = ~n5039 & ~n5040 ;
  assign n5042 = ~n4792 & n5041 ;
  assign n5043 = \i_tv80_core_PC_reg[15]/P0001  & ~n1103 ;
  assign n5044 = \i_tv80_core_PC_reg[15]/P0001  & ~n1317 ;
  assign n5045 = ~n2252 & ~n5044 ;
  assign n5046 = n1886 & ~n5045 ;
  assign n5047 = ~n2294 & ~n5046 ;
  assign n5048 = ~n1277 & ~n5047 ;
  assign n5049 = ~n2297 & ~n5048 ;
  assign n5050 = n1625 & ~n5049 ;
  assign n5051 = ~n2300 & ~n5050 ;
  assign n5052 = n1103 & ~n5051 ;
  assign n5053 = ~n5043 & ~n5052 ;
  assign n5054 = n4792 & n5053 ;
  assign n5055 = n1635 & ~n5054 ;
  assign n5056 = ~n5042 & n5055 ;
  assign n5057 = ~n1635 & ~n5053 ;
  assign n5058 = ~n1113 & ~n5057 ;
  assign n5059 = ~n5056 & n5058 ;
  assign n5060 = n4744 & n5041 ;
  assign n5061 = ~\i_tv80_core_PC_reg[15]/P0001  & ~n4744 ;
  assign n5062 = n1635 & ~n5061 ;
  assign n5063 = ~n5060 & n5062 ;
  assign n5064 = \i_tv80_core_PC_reg[15]/P0001  & ~n1635 ;
  assign n5065 = n1113 & ~n5064 ;
  assign n5066 = ~n5063 & n5065 ;
  assign n5067 = ~n5059 & ~n5066 ;
  assign n5068 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5067 ;
  assign n5069 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PC_reg[15]/P0001  ;
  assign n5070 = reset_n_pad & ~n5069 ;
  assign n5071 = ~n5068 & n5070 ;
  assign n5074 = ~n4846 & ~n4847 ;
  assign n5075 = n4757 & ~n5074 ;
  assign n5076 = ~n4757 & n5074 ;
  assign n5077 = ~n5075 & ~n5076 ;
  assign n5078 = n4745 & ~n5077 ;
  assign n5073 = \i_tv80_core_PC_reg[1]/P0001  & ~n4745 ;
  assign n5079 = n1113 & ~n5073 ;
  assign n5080 = ~n5078 & n5079 ;
  assign n5082 = \i_tv80_core_PC_reg[1]/P0001  & n1318 ;
  assign n5083 = n1662 & ~n5082 ;
  assign n5084 = ~n1277 & ~n5083 ;
  assign n5085 = ~n1660 & ~n5084 ;
  assign n5086 = n1625 & ~n5085 ;
  assign n5087 = n1688 & ~n5086 ;
  assign n5088 = ~\i_tv80_core_PC_reg[1]/P0001  & ~n1103 ;
  assign n5089 = ~n4793 & ~n5088 ;
  assign n5090 = ~n5087 & n5089 ;
  assign n5081 = n4793 & ~n5077 ;
  assign n5091 = ~n1113 & ~n5081 ;
  assign n5092 = ~n5090 & n5091 ;
  assign n5093 = ~n5080 & ~n5092 ;
  assign n5094 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5093 ;
  assign n5072 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PC_reg[1]/P0001  ;
  assign n5095 = reset_n_pad & ~n5072 ;
  assign n5096 = ~n5094 & n5095 ;
  assign n5099 = ~n4842 & ~n4843 ;
  assign n5100 = ~n4849 & n5099 ;
  assign n5101 = n4849 & ~n5099 ;
  assign n5102 = ~n5100 & ~n5101 ;
  assign n5103 = n4745 & ~n5102 ;
  assign n5098 = \i_tv80_core_PC_reg[2]/P0001  & ~n4745 ;
  assign n5104 = n1113 & ~n5098 ;
  assign n5105 = ~n5103 & n5104 ;
  assign n5107 = \i_tv80_core_PC_reg[2]/P0001  & n1318 ;
  assign n5108 = n1333 & ~n5107 ;
  assign n5109 = ~n1277 & ~n5108 ;
  assign n5110 = ~n1305 & ~n5109 ;
  assign n5111 = n1625 & ~n5110 ;
  assign n5112 = n1628 & ~n5111 ;
  assign n5113 = ~\i_tv80_core_PC_reg[2]/P0001  & ~n1103 ;
  assign n5114 = ~n4793 & ~n5113 ;
  assign n5115 = ~n5112 & n5114 ;
  assign n5106 = n4793 & ~n5102 ;
  assign n5116 = ~n1113 & ~n5106 ;
  assign n5117 = ~n5115 & n5116 ;
  assign n5118 = ~n5105 & ~n5117 ;
  assign n5119 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5118 ;
  assign n5097 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PC_reg[2]/P0001  ;
  assign n5120 = reset_n_pad & ~n5097 ;
  assign n5121 = ~n5119 & n5120 ;
  assign n5132 = ~\i_tv80_core_PC_reg[3]/P0001  & ~n1103 ;
  assign n5133 = \i_tv80_core_PC_reg[3]/P0001  & ~n1317 ;
  assign n5134 = ~n2315 & ~n5133 ;
  assign n5135 = n1886 & ~n5134 ;
  assign n5136 = ~n2353 & ~n5135 ;
  assign n5137 = ~n1277 & ~n5136 ;
  assign n5138 = ~n2356 & ~n5137 ;
  assign n5139 = n1625 & ~n5138 ;
  assign n5140 = n2360 & ~n5139 ;
  assign n5141 = ~n5132 & ~n5140 ;
  assign n5142 = ~n4793 & ~n5141 ;
  assign n5124 = ~n4838 & ~n4839 ;
  assign n5125 = ~n4851 & n5124 ;
  assign n5126 = n4851 & ~n5124 ;
  assign n5127 = ~n5125 & ~n5126 ;
  assign n5131 = n4793 & n5127 ;
  assign n5143 = ~n1113 & ~n5131 ;
  assign n5144 = ~n5142 & n5143 ;
  assign n5128 = n4745 & n5127 ;
  assign n5123 = ~\i_tv80_core_PC_reg[3]/P0001  & ~n4745 ;
  assign n5129 = n1113 & ~n5123 ;
  assign n5130 = ~n5128 & n5129 ;
  assign n5145 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5130 ;
  assign n5146 = ~n5144 & n5145 ;
  assign n5122 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PC_reg[3]/P0001  ;
  assign n5147 = reset_n_pad & ~n5122 ;
  assign n5148 = ~n5146 & n5147 ;
  assign n5159 = ~\i_tv80_core_PC_reg[4]/P0001  & ~n1103 ;
  assign n5160 = \i_tv80_core_PC_reg[4]/P0001  & ~n1317 ;
  assign n5161 = ~n2374 & ~n5160 ;
  assign n5162 = n1886 & ~n5161 ;
  assign n5163 = ~n2412 & ~n5162 ;
  assign n5164 = ~n1277 & ~n5163 ;
  assign n5165 = ~n2415 & ~n5164 ;
  assign n5166 = n1625 & ~n5165 ;
  assign n5167 = n2419 & ~n5166 ;
  assign n5168 = ~n5159 & ~n5167 ;
  assign n5169 = ~n4793 & ~n5168 ;
  assign n5151 = ~n4834 & ~n4835 ;
  assign n5152 = ~n4853 & n5151 ;
  assign n5153 = n4853 & ~n5151 ;
  assign n5154 = ~n5152 & ~n5153 ;
  assign n5158 = n4793 & n5154 ;
  assign n5170 = ~n1113 & ~n5158 ;
  assign n5171 = ~n5169 & n5170 ;
  assign n5155 = n4745 & n5154 ;
  assign n5150 = ~\i_tv80_core_PC_reg[4]/P0001  & ~n4745 ;
  assign n5156 = n1113 & ~n5150 ;
  assign n5157 = ~n5155 & n5156 ;
  assign n5172 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5157 ;
  assign n5173 = ~n5171 & n5172 ;
  assign n5149 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PC_reg[4]/P0001  ;
  assign n5174 = reset_n_pad & ~n5149 ;
  assign n5175 = ~n5173 & n5174 ;
  assign n5186 = ~\i_tv80_core_PC_reg[5]/P0001  & ~n1103 ;
  assign n5187 = \i_tv80_core_PC_reg[5]/P0001  & n1318 ;
  assign n5188 = n1719 & ~n5187 ;
  assign n5189 = ~n1277 & ~n5188 ;
  assign n5190 = ~n1717 & ~n5189 ;
  assign n5191 = n1625 & ~n5190 ;
  assign n5192 = n1749 & ~n5191 ;
  assign n5193 = ~n5186 & ~n5192 ;
  assign n5194 = ~n4793 & ~n5193 ;
  assign n5177 = ~n4830 & ~n4831 ;
  assign n5178 = ~n4855 & n5177 ;
  assign n5179 = n4855 & ~n5177 ;
  assign n5180 = ~n5178 & ~n5179 ;
  assign n5185 = n4793 & n5180 ;
  assign n5195 = ~n1113 & ~n5185 ;
  assign n5196 = ~n5194 & n5195 ;
  assign n5181 = n4745 & n5180 ;
  assign n5182 = ~\i_tv80_core_PC_reg[5]/P0001  & ~n4745 ;
  assign n5183 = n1113 & ~n5182 ;
  assign n5184 = ~n5181 & n5183 ;
  assign n5197 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5184 ;
  assign n5198 = ~n5196 & n5197 ;
  assign n5176 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PC_reg[5]/P0001  ;
  assign n5199 = reset_n_pad & ~n5176 ;
  assign n5200 = ~n5198 & n5199 ;
  assign n5202 = ~n4826 & ~n4827 ;
  assign n5203 = ~n4857 & n5202 ;
  assign n5204 = n4857 & ~n5202 ;
  assign n5205 = ~n5203 & ~n5204 ;
  assign n5219 = n4793 & n5205 ;
  assign n5210 = ~\i_tv80_core_PC_reg[6]/P0001  & ~n1103 ;
  assign n5211 = \i_tv80_core_PC_reg[6]/P0001  & n1318 ;
  assign n5212 = n1780 & ~n5211 ;
  assign n5213 = ~n1277 & ~n5212 ;
  assign n5214 = ~n1778 & ~n5213 ;
  assign n5215 = n1625 & ~n5214 ;
  assign n5216 = n1807 & ~n5215 ;
  assign n5217 = ~n5210 & ~n5216 ;
  assign n5218 = ~n4793 & ~n5217 ;
  assign n5220 = ~n1113 & ~n5218 ;
  assign n5221 = ~n5219 & n5220 ;
  assign n5206 = n4745 & n5205 ;
  assign n5207 = ~\i_tv80_core_PC_reg[6]/P0001  & ~n4745 ;
  assign n5208 = n1113 & ~n5207 ;
  assign n5209 = ~n5206 & n5208 ;
  assign n5222 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5209 ;
  assign n5223 = ~n5221 & n5222 ;
  assign n5201 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PC_reg[6]/P0001  ;
  assign n5224 = reset_n_pad & ~n5201 ;
  assign n5225 = ~n5223 & n5224 ;
  assign n5227 = ~n4821 & ~n4823 ;
  assign n5228 = ~n4859 & n5227 ;
  assign n5229 = n4859 & ~n5227 ;
  assign n5230 = ~n5228 & ~n5229 ;
  assign n5246 = n4793 & n5230 ;
  assign n5235 = ~\i_tv80_core_PC_reg[7]/P0001  & ~n1103 ;
  assign n5236 = \i_tv80_core_PC_reg[7]/P0001  & ~n1317 ;
  assign n5237 = ~n2433 & ~n5236 ;
  assign n5238 = n1886 & ~n5237 ;
  assign n5239 = ~n2472 & ~n5238 ;
  assign n5240 = ~n1277 & ~n5239 ;
  assign n5241 = ~n2475 & ~n5240 ;
  assign n5242 = n1625 & ~n5241 ;
  assign n5243 = n2479 & ~n5242 ;
  assign n5244 = ~n5235 & ~n5243 ;
  assign n5245 = ~n4793 & ~n5244 ;
  assign n5247 = ~n1113 & ~n5245 ;
  assign n5248 = ~n5246 & n5247 ;
  assign n5231 = n4745 & n5230 ;
  assign n5232 = ~\i_tv80_core_PC_reg[7]/P0001  & ~n4745 ;
  assign n5233 = n1113 & ~n5232 ;
  assign n5234 = ~n5231 & n5233 ;
  assign n5249 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5234 ;
  assign n5250 = ~n5248 & n5249 ;
  assign n5226 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PC_reg[7]/P0001  ;
  assign n5251 = reset_n_pad & ~n5226 ;
  assign n5252 = ~n5250 & n5251 ;
  assign n5254 = ~n4818 & ~n4820 ;
  assign n5255 = ~n4821 & ~n4860 ;
  assign n5256 = n5254 & n5255 ;
  assign n5257 = ~n5254 & ~n5255 ;
  assign n5258 = ~n5256 & ~n5257 ;
  assign n5274 = n4793 & ~n5258 ;
  assign n5263 = ~\i_tv80_core_PC_reg[8]/P0001  & ~n1103 ;
  assign n5264 = \i_tv80_core_PC_reg[8]/P0001  & ~n1317 ;
  assign n5265 = ~n2493 & ~n5264 ;
  assign n5266 = n1886 & ~n5265 ;
  assign n5267 = ~n2534 & ~n5266 ;
  assign n5268 = ~n1277 & ~n5267 ;
  assign n5269 = ~n2537 & ~n5268 ;
  assign n5270 = n1625 & ~n5269 ;
  assign n5271 = n2541 & ~n5270 ;
  assign n5272 = ~n5263 & ~n5271 ;
  assign n5273 = ~n4793 & ~n5272 ;
  assign n5275 = ~n1113 & ~n5273 ;
  assign n5276 = ~n5274 & n5275 ;
  assign n5259 = n4745 & ~n5258 ;
  assign n5260 = ~\i_tv80_core_PC_reg[8]/P0001  & ~n4745 ;
  assign n5261 = n1113 & ~n5260 ;
  assign n5262 = ~n5259 & n5261 ;
  assign n5277 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5262 ;
  assign n5278 = ~n5276 & n5277 ;
  assign n5253 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PC_reg[8]/P0001  ;
  assign n5279 = reset_n_pad & ~n5253 ;
  assign n5280 = ~n5278 & n5279 ;
  assign n5282 = ~n4819 & ~n4861 ;
  assign n5283 = ~n4898 & n5282 ;
  assign n5284 = n4898 & ~n5282 ;
  assign n5285 = ~n5283 & ~n5284 ;
  assign n5290 = n4793 & ~n5285 ;
  assign n5300 = \i_tv80_core_PC_reg[9]/P0001  & ~n1103 ;
  assign n5291 = \i_tv80_core_PC_reg[9]/P0001  & ~n1317 ;
  assign n5292 = ~n2555 & ~n5291 ;
  assign n5293 = n1886 & ~n5292 ;
  assign n5294 = ~n2596 & ~n5293 ;
  assign n5295 = ~n1277 & ~n5294 ;
  assign n5296 = ~n2599 & ~n5295 ;
  assign n5297 = n1625 & ~n5296 ;
  assign n5298 = ~n2602 & ~n5297 ;
  assign n5299 = n1103 & ~n5298 ;
  assign n5301 = ~n4793 & ~n5299 ;
  assign n5302 = ~n5300 & n5301 ;
  assign n5303 = ~n1113 & ~n5302 ;
  assign n5304 = ~n5290 & n5303 ;
  assign n5286 = n4745 & ~n5285 ;
  assign n5287 = ~\i_tv80_core_PC_reg[9]/P0001  & ~n4745 ;
  assign n5288 = n1113 & ~n5287 ;
  assign n5289 = ~n5286 & n5288 ;
  assign n5305 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5289 ;
  assign n5306 = ~n5304 & n5305 ;
  assign n5281 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PC_reg[9]/P0001  ;
  assign n5307 = reset_n_pad & ~n5281 ;
  assign n5308 = ~n5306 & n5307 ;
  assign n5309 = ~\i_tv80_core_tstate_reg[2]/NET0131  & n2661 ;
  assign n5310 = n860 & n1635 ;
  assign n5311 = ~\m1_n_pad  & ~n5310 ;
  assign n5312 = ~n5309 & ~n5311 ;
  assign n5313 = ~n4716 & n5312 ;
  assign n5314 = reset_n_pad & ~n5313 ;
  assign n5315 = ~\i_tv80_core_NMI_s_reg/P0001  & ~n4721 ;
  assign n5316 = n4726 & ~n5315 ;
  assign n5319 = ~n1615 & ~n4719 ;
  assign n5320 = n1634 & ~n5319 ;
  assign n5321 = ~\i_tv80_core_IntE_FF1_reg/P0001  & ~n5320 ;
  assign n5317 = ~\i_tv80_core_IntE_FF2_reg/P0001  & n1634 ;
  assign n5318 = n1615 & n5317 ;
  assign n5322 = n4734 & ~n5318 ;
  assign n5323 = ~n5321 & n5322 ;
  assign n5324 = ~n5316 & n5323 ;
  assign n5330 = ~n3203 & ~n3206 ;
  assign n5331 = ~n3195 & n5330 ;
  assign n5332 = n3195 & ~n5330 ;
  assign n5333 = ~n5331 & ~n5332 ;
  assign n5334 = n3001 & n5333 ;
  assign n5329 = \i_tv80_core_SP_reg[9]/P0001  & ~n3002 ;
  assign n5335 = ~n2997 & ~n5329 ;
  assign n5336 = ~n5334 & n5335 ;
  assign n5328 = n2571 & n2997 ;
  assign n5337 = ~n1113 & ~n5328 ;
  assign n5338 = ~n5336 & n5337 ;
  assign n5327 = \i_tv80_core_SP_reg[9]/P0001  & n1113 ;
  assign n5339 = ~n3242 & ~n5327 ;
  assign n5340 = ~n5338 & n5339 ;
  assign n5326 = n3242 & n3982 ;
  assign n5341 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5326 ;
  assign n5342 = ~n5340 & n5341 ;
  assign n5325 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[9]/P0001  ;
  assign n5343 = reset_n_pad & ~n5325 ;
  assign n5344 = ~n5342 & n5343 ;
  assign n5349 = \i_tv80_core_SP_reg[11]/P0001  & ~n3170 ;
  assign n5350 = ~n3213 & ~n3222 ;
  assign n5351 = ~n3209 & n5350 ;
  assign n5352 = n3209 & ~n5350 ;
  assign n5353 = ~n5351 & ~n5352 ;
  assign n5354 = n2699 & n5353 ;
  assign n5355 = ~n5349 & ~n5354 ;
  assign n5356 = ~n3000 & ~n5355 ;
  assign n5348 = \i_tv80_core_SP_reg[11]/P0001  & n3000 ;
  assign n5357 = ~n2997 & ~n5348 ;
  assign n5358 = ~n5356 & n5357 ;
  assign n5347 = n2016 & n2997 ;
  assign n5359 = ~n1113 & ~n5347 ;
  assign n5360 = ~n5358 & n5359 ;
  assign n5346 = \i_tv80_core_SP_reg[11]/P0001  & n1113 ;
  assign n5361 = ~n3242 & ~n5346 ;
  assign n5362 = ~n5360 & n5361 ;
  assign n5345 = n3242 & n3771 ;
  assign n5363 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5345 ;
  assign n5364 = ~n5362 & n5363 ;
  assign n5365 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[11]/P0001  ;
  assign n5366 = reset_n_pad & ~n5365 ;
  assign n5367 = ~n5364 & n5366 ;
  assign n5368 = \i_tv80_core_NMICycle_reg/P0001  & ~n4716 ;
  assign n5369 = \i_tv80_core_NMI_s_reg/P0001  & n4726 ;
  assign n5370 = ~n5368 & ~n5369 ;
  assign n5371 = reset_n_pad & ~n5370 ;
  assign n5374 = n4300 & n4318 ;
  assign n5375 = \i_tv80_core_TmpAddr_reg[10]/P0001  & n4303 ;
  assign n5376 = ~n5374 & ~n5375 ;
  assign n5377 = ~n4298 & ~n5376 ;
  assign n5373 = \di_reg_reg[2]/P0001  & n4298 ;
  assign n5378 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5373 ;
  assign n5379 = ~n5377 & n5378 ;
  assign n5372 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[10]/P0001  ;
  assign n5380 = reset_n_pad & ~n5372 ;
  assign n5381 = ~n5379 & n5380 ;
  assign n5383 = n2968 & ~n3107 ;
  assign n5385 = ~\i_tv80_core_BusB_reg[0]/P0001  & ~n2975 ;
  assign n5386 = ~\i_tv80_core_BusA_reg[0]/P0001  & n2975 ;
  assign n5387 = ~n5385 & ~n5386 ;
  assign n5388 = ~n2973 & ~n5387 ;
  assign n5389 = ~\i_tv80_core_BusB_reg[4]/P0001  & n2973 ;
  assign n5390 = ~n5388 & ~n5389 ;
  assign n5391 = n1157 & ~n5390 ;
  assign n5384 = ~\do[0]_pad  & ~n1157 ;
  assign n5392 = ~n2968 & ~n5384 ;
  assign n5393 = ~n5391 & n5392 ;
  assign n5394 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5393 ;
  assign n5395 = ~n5383 & n5394 ;
  assign n5382 = ~\do[0]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n5396 = reset_n_pad & ~n5382 ;
  assign n5397 = ~n5395 & n5396 ;
  assign n5399 = n2968 & ~n3982 ;
  assign n5401 = ~\i_tv80_core_BusB_reg[1]/P0001  & ~n2975 ;
  assign n5402 = ~\i_tv80_core_BusA_reg[1]/P0001  & n2975 ;
  assign n5403 = ~n5401 & ~n5402 ;
  assign n5404 = ~n2973 & ~n5403 ;
  assign n5405 = ~\i_tv80_core_BusB_reg[5]/P0001  & n2973 ;
  assign n5406 = ~n5404 & ~n5405 ;
  assign n5407 = n1157 & ~n5406 ;
  assign n5400 = ~\do[1]_pad  & ~n1157 ;
  assign n5408 = ~n2968 & ~n5400 ;
  assign n5409 = ~n5407 & n5408 ;
  assign n5410 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5409 ;
  assign n5411 = ~n5399 & n5410 ;
  assign n5398 = ~\do[1]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n5412 = reset_n_pad & ~n5398 ;
  assign n5413 = ~n5411 & n5412 ;
  assign n5415 = ~n1193 & n2968 ;
  assign n5417 = ~\i_tv80_core_BusB_reg[2]/P0001  & ~n2975 ;
  assign n5418 = ~\i_tv80_core_BusA_reg[2]/P0001  & n2975 ;
  assign n5419 = ~n5417 & ~n5418 ;
  assign n5420 = ~n2973 & ~n5419 ;
  assign n5421 = ~\i_tv80_core_BusB_reg[6]/P0001  & n2973 ;
  assign n5422 = ~n5420 & ~n5421 ;
  assign n5423 = n1157 & ~n5422 ;
  assign n5416 = ~\do[2]_pad  & ~n1157 ;
  assign n5424 = ~n2968 & ~n5416 ;
  assign n5425 = ~n5423 & n5424 ;
  assign n5426 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5425 ;
  assign n5427 = ~n5415 & n5426 ;
  assign n5414 = ~\do[2]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n5428 = reset_n_pad & ~n5414 ;
  assign n5429 = ~n5427 & n5428 ;
  assign n5431 = n2968 & ~n3771 ;
  assign n5433 = ~\i_tv80_core_BusB_reg[3]/P0001  & ~n2975 ;
  assign n5434 = ~\i_tv80_core_BusA_reg[3]/P0001  & n2975 ;
  assign n5435 = ~n5433 & ~n5434 ;
  assign n5436 = ~n2973 & ~n5435 ;
  assign n5437 = ~\i_tv80_core_BusB_reg[7]/P0001  & n2973 ;
  assign n5438 = ~n5436 & ~n5437 ;
  assign n5439 = n1157 & ~n5438 ;
  assign n5432 = ~\do[3]_pad  & ~n1157 ;
  assign n5440 = ~n2968 & ~n5432 ;
  assign n5441 = ~n5439 & n5440 ;
  assign n5442 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5441 ;
  assign n5443 = ~n5431 & n5442 ;
  assign n5430 = ~\do[3]_pad  & \i_tv80_core_BusAck_reg/P0001  ;
  assign n5444 = reset_n_pad & ~n5430 ;
  assign n5445 = ~n5443 & n5444 ;
  assign n5450 = ~n3190 & ~n3193 ;
  assign n5451 = ~n3834 & n5450 ;
  assign n5452 = n3834 & ~n5450 ;
  assign n5453 = ~n5451 & ~n5452 ;
  assign n5454 = n3001 & n5453 ;
  assign n5449 = \i_tv80_core_SP_reg[8]/P0001  & ~n3002 ;
  assign n5455 = ~n2997 & ~n5449 ;
  assign n5456 = ~n5454 & n5455 ;
  assign n5448 = n2509 & n2997 ;
  assign n5457 = ~n1113 & ~n5448 ;
  assign n5458 = ~n5456 & n5457 ;
  assign n5447 = \i_tv80_core_SP_reg[8]/P0001  & n1113 ;
  assign n5459 = ~n3242 & ~n5447 ;
  assign n5460 = ~n5458 & n5459 ;
  assign n5461 = n3107 & n3242 ;
  assign n5462 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5461 ;
  assign n5463 = ~n5460 & n5462 ;
  assign n5446 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[8]/P0001  ;
  assign n5464 = reset_n_pad & ~n5446 ;
  assign n5465 = ~n5463 & n5464 ;
  assign n5466 = n1599 & n4401 ;
  assign n5468 = ~\i_tv80_core_mcycle_reg[0]/P0001  & n5466 ;
  assign n5467 = ~\i_tv80_core_Pre_XY_F_M_reg[0]/P0001  & ~n5466 ;
  assign n5469 = reset_n_pad & ~n5467 ;
  assign n5470 = ~n5468 & n5469 ;
  assign n5472 = ~\i_tv80_core_mcycle_reg[1]/P0001  & n5466 ;
  assign n5471 = ~\i_tv80_core_Pre_XY_F_M_reg[1]/P0001  & ~n5466 ;
  assign n5473 = reset_n_pad & ~n5471 ;
  assign n5474 = ~n5472 & n5473 ;
  assign n5476 = ~\i_tv80_core_mcycle_reg[2]/P0001  & n5466 ;
  assign n5475 = ~\i_tv80_core_Pre_XY_F_M_reg[2]/P0001  & ~n5466 ;
  assign n5477 = reset_n_pad & ~n5475 ;
  assign n5478 = ~n5476 & n5477 ;
  assign n5481 = n4300 & n4469 ;
  assign n5482 = \i_tv80_core_TmpAddr_reg[12]/P0001  & n4303 ;
  assign n5483 = ~n5481 & ~n5482 ;
  assign n5484 = ~n4298 & ~n5483 ;
  assign n5480 = \di_reg_reg[4]/P0001  & n4298 ;
  assign n5485 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5480 ;
  assign n5486 = ~n5484 & n5485 ;
  assign n5479 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[12]/P0001  ;
  assign n5487 = reset_n_pad & ~n5479 ;
  assign n5488 = ~n5486 & n5487 ;
  assign n5491 = n4300 & n4490 ;
  assign n5492 = \i_tv80_core_TmpAddr_reg[13]/P0001  & n4303 ;
  assign n5493 = ~n5491 & ~n5492 ;
  assign n5494 = ~n4298 & ~n5493 ;
  assign n5490 = \di_reg_reg[5]/P0001  & n4298 ;
  assign n5495 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5490 ;
  assign n5496 = ~n5494 & n5495 ;
  assign n5489 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[13]/P0001  ;
  assign n5497 = reset_n_pad & ~n5489 ;
  assign n5498 = ~n5496 & n5497 ;
  assign n5501 = n3232 & n4300 ;
  assign n5502 = \i_tv80_core_TmpAddr_reg[15]/P0001  & n4303 ;
  assign n5503 = ~n5501 & ~n5502 ;
  assign n5504 = ~n4298 & ~n5503 ;
  assign n5500 = \di_reg_reg[7]/P0001  & n4298 ;
  assign n5505 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5500 ;
  assign n5506 = ~n5504 & n5505 ;
  assign n5499 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[15]/P0001  ;
  assign n5507 = reset_n_pad & ~n5499 ;
  assign n5508 = ~n5506 & n5507 ;
  assign n5509 = \i_tv80_core_i_reg_RegsL_reg[0][1]/P0001  & ~n2696 ;
  assign n5512 = ~n2755 & n2790 ;
  assign n5510 = ~n2755 & ~n2789 ;
  assign n5511 = n2788 & ~n5510 ;
  assign n5513 = n2891 & ~n5511 ;
  assign n5514 = ~n5512 & n5513 ;
  assign n5515 = \i_tv80_core_RegBusA_r_reg[1]/P0001  & n2664 ;
  assign n5516 = ~n4042 & ~n5515 ;
  assign n5517 = ~n5514 & n5516 ;
  assign n5518 = ~n2667 & ~n5517 ;
  assign n5523 = \i_tv80_core_i_reg_RegsL_reg[4][1]/P0001  & n2918 ;
  assign n5524 = \i_tv80_core_i_reg_RegsL_reg[5][1]/P0001  & n2916 ;
  assign n5529 = ~n5523 & ~n5524 ;
  assign n5525 = \i_tv80_core_i_reg_RegsL_reg[7][1]/P0001  & n2904 ;
  assign n5526 = \i_tv80_core_i_reg_RegsL_reg[2][1]/P0001  & n2908 ;
  assign n5530 = ~n5525 & ~n5526 ;
  assign n5531 = n5529 & n5530 ;
  assign n5519 = \i_tv80_core_i_reg_RegsL_reg[6][1]/P0001  & n2920 ;
  assign n5520 = \i_tv80_core_i_reg_RegsL_reg[3][1]/P0001  & n2922 ;
  assign n5527 = ~n5519 & ~n5520 ;
  assign n5521 = \i_tv80_core_i_reg_RegsL_reg[1][1]/P0001  & n2914 ;
  assign n5522 = \i_tv80_core_i_reg_RegsL_reg[0][1]/P0001  & n2911 ;
  assign n5528 = ~n5521 & ~n5522 ;
  assign n5532 = n5527 & n5528 ;
  assign n5533 = n5531 & n5532 ;
  assign n5534 = n2667 & ~n5533 ;
  assign n5535 = ~n5518 & ~n5534 ;
  assign n5536 = n2696 & ~n5535 ;
  assign n5537 = ~n5509 & ~n5536 ;
  assign n5538 = \i_tv80_core_i_reg_RegsL_reg[1][1]/P0001  & ~n2741 ;
  assign n5539 = n2741 & ~n5535 ;
  assign n5540 = ~n5538 & ~n5539 ;
  assign n5541 = \i_tv80_core_i_reg_RegsL_reg[2][1]/P0001  & ~n2745 ;
  assign n5542 = n2745 & ~n5535 ;
  assign n5543 = ~n5541 & ~n5542 ;
  assign n5544 = \i_tv80_core_i_reg_RegsL_reg[3][1]/P0001  & ~n2743 ;
  assign n5545 = n2743 & ~n5535 ;
  assign n5546 = ~n5544 & ~n5545 ;
  assign n5547 = \i_tv80_core_i_reg_RegsL_reg[4][1]/P0001  & ~n2733 ;
  assign n5548 = n2733 & ~n5535 ;
  assign n5549 = ~n5547 & ~n5548 ;
  assign n5550 = \i_tv80_core_i_reg_RegsL_reg[5][1]/P0001  & ~n2739 ;
  assign n5551 = n2739 & ~n5535 ;
  assign n5552 = ~n5550 & ~n5551 ;
  assign n5553 = \i_tv80_core_i_reg_RegsL_reg[6][1]/P0001  & ~n2736 ;
  assign n5554 = n2736 & ~n5535 ;
  assign n5555 = ~n5553 & ~n5554 ;
  assign n5556 = \i_tv80_core_i_reg_RegsL_reg[7][1]/P0001  & ~n2731 ;
  assign n5557 = n2731 & ~n5535 ;
  assign n5558 = ~n5556 & ~n5557 ;
  assign n5561 = n2330 & n2997 ;
  assign n5563 = ~n3025 & ~n3049 ;
  assign n5564 = n3047 & ~n5563 ;
  assign n5565 = n3048 & ~n3049 ;
  assign n5566 = ~n5564 & ~n5565 ;
  assign n5567 = n3001 & n5566 ;
  assign n5562 = \i_tv80_core_SP_reg[3]/P0001  & ~n3002 ;
  assign n5568 = ~n2997 & ~n5562 ;
  assign n5569 = ~n5567 & n5568 ;
  assign n5570 = ~n5561 & ~n5569 ;
  assign n5571 = ~n1113 & ~n5570 ;
  assign n5572 = ~\i_tv80_core_SP_reg[3]/P0001  & n1113 ;
  assign n5573 = ~n5571 & ~n5572 ;
  assign n5574 = ~n2992 & ~n5573 ;
  assign n5560 = n2992 & n3771 ;
  assign n5575 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5560 ;
  assign n5576 = ~n5574 & n5575 ;
  assign n5559 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[3]/P0001  ;
  assign n5577 = reset_n_pad & ~n5559 ;
  assign n5578 = ~n5576 & n5577 ;
  assign n5581 = ~n2997 & ~n3002 ;
  assign n5582 = ~n1113 & ~n5581 ;
  assign n5583 = \i_tv80_core_SP_reg[0]/P0001  & ~n5582 ;
  assign n5584 = ~n1883 & n2997 ;
  assign n5585 = ~\di_reg_reg[0]/P0001  & n1107 ;
  assign n5586 = n1883 & n5585 ;
  assign n5587 = n3042 & ~n5586 ;
  assign n5588 = ~n2997 & n5587 ;
  assign n5589 = n3001 & n5588 ;
  assign n5590 = ~n5584 & ~n5589 ;
  assign n5591 = ~n1113 & ~n5590 ;
  assign n5592 = ~n2992 & ~n5591 ;
  assign n5593 = ~n5583 & n5592 ;
  assign n5580 = n2992 & n3107 ;
  assign n5594 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5580 ;
  assign n5595 = ~n5593 & n5594 ;
  assign n5579 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[0]/P0001  ;
  assign n5596 = reset_n_pad & ~n5579 ;
  assign n5597 = ~n5595 & n5596 ;
  assign n5601 = ~n3038 & ~n3044 ;
  assign n5602 = n3042 & ~n5601 ;
  assign n5603 = ~n3042 & n5601 ;
  assign n5604 = ~n5602 & ~n5603 ;
  assign n5605 = n3001 & n5604 ;
  assign n5606 = \i_tv80_core_SP_reg[1]/P0001  & ~n3002 ;
  assign n5607 = ~n2997 & ~n5606 ;
  assign n5608 = ~n5605 & n5607 ;
  assign n5600 = n1659 & n2997 ;
  assign n5609 = ~n1113 & ~n5600 ;
  assign n5610 = ~n5608 & n5609 ;
  assign n5611 = \i_tv80_core_SP_reg[1]/P0001  & n1113 ;
  assign n5612 = ~n2992 & ~n5611 ;
  assign n5613 = ~n5610 & n5612 ;
  assign n5599 = n2992 & n3982 ;
  assign n5614 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5599 ;
  assign n5615 = ~n5613 & n5614 ;
  assign n5598 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[1]/P0001  ;
  assign n5616 = reset_n_pad & ~n5598 ;
  assign n5617 = ~n5615 & n5616 ;
  assign n5621 = ~n3031 & ~n3032 ;
  assign n5622 = n3045 & ~n5621 ;
  assign n5623 = ~n3045 & n5621 ;
  assign n5624 = ~n5622 & ~n5623 ;
  assign n5625 = n3001 & n5624 ;
  assign n5626 = \i_tv80_core_SP_reg[2]/P0001  & ~n3002 ;
  assign n5627 = ~n2997 & ~n5626 ;
  assign n5628 = ~n5625 & n5627 ;
  assign n5620 = n1304 & n2997 ;
  assign n5629 = ~n1113 & ~n5620 ;
  assign n5630 = ~n5628 & n5629 ;
  assign n5631 = \i_tv80_core_SP_reg[2]/P0001  & n1113 ;
  assign n5632 = ~n2992 & ~n5631 ;
  assign n5633 = ~n5630 & n5632 ;
  assign n5619 = n1193 & n2992 ;
  assign n5634 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5619 ;
  assign n5635 = ~n5633 & n5634 ;
  assign n5618 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_SP_reg[2]/P0001  ;
  assign n5636 = reset_n_pad & ~n5618 ;
  assign n5637 = ~n5635 & n5636 ;
  assign n5640 = n4300 & n5353 ;
  assign n5641 = \i_tv80_core_TmpAddr_reg[11]/P0001  & n4303 ;
  assign n5642 = ~n5640 & ~n5641 ;
  assign n5643 = ~n4298 & ~n5642 ;
  assign n5639 = \di_reg_reg[3]/P0001  & n4298 ;
  assign n5644 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5639 ;
  assign n5645 = ~n5643 & n5644 ;
  assign n5638 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[11]/P0001  ;
  assign n5646 = reset_n_pad & ~n5638 ;
  assign n5647 = ~n5645 & n5646 ;
  assign n5652 = ~\i_tv80_core_TmpAddr_reg[9]/P0001  & n1113 ;
  assign n5653 = n4300 & n5333 ;
  assign n5649 = \i_tv80_core_TmpAddr_reg[9]/P0001  & n4303 ;
  assign n5654 = ~n1113 & ~n5649 ;
  assign n5655 = ~n5653 & n5654 ;
  assign n5656 = ~n5652 & ~n5655 ;
  assign n5657 = n4297 & ~n5656 ;
  assign n5651 = ~\di_reg_reg[1]/P0001  & ~n4297 ;
  assign n5658 = n1107 & ~n5651 ;
  assign n5659 = ~n5657 & n5658 ;
  assign n5650 = ~n1107 & n5649 ;
  assign n5660 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5650 ;
  assign n5661 = ~n5659 & n5660 ;
  assign n5648 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[9]/P0001  ;
  assign n5662 = reset_n_pad & ~n5648 ;
  assign n5663 = ~n5661 & n5662 ;
  assign n5665 = ~n1014 & ~n1451 ;
  assign n5666 = n858 & ~n5665 ;
  assign n5667 = ~n860 & ~n1481 ;
  assign n5668 = n1617 & ~n5667 ;
  assign n5669 = n945 & n4769 ;
  assign n5670 = n857 & ~n5669 ;
  assign n5671 = ~n5668 & ~n5670 ;
  assign n5672 = n382 & ~n5671 ;
  assign n5673 = ~n5666 & ~n5672 ;
  assign n5674 = n1107 & ~n5673 ;
  assign n5676 = ~n3738 & n4300 ;
  assign n5677 = \i_tv80_core_TmpAddr_reg[6]/P0001  & n4303 ;
  assign n5678 = ~n5676 & ~n5677 ;
  assign n5679 = ~n5674 & ~n5678 ;
  assign n5675 = \di_reg_reg[6]/P0001  & n5674 ;
  assign n5680 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5675 ;
  assign n5681 = ~n5679 & n5680 ;
  assign n5664 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[6]/P0001  ;
  assign n5682 = reset_n_pad & ~n5664 ;
  assign n5683 = ~n5681 & n5682 ;
  assign n5686 = n4300 & n5453 ;
  assign n5685 = \i_tv80_core_TmpAddr_reg[8]/P0001  & n4303 ;
  assign n5687 = ~n4298 & ~n5685 ;
  assign n5688 = ~n5686 & n5687 ;
  assign n5689 = ~\di_reg_reg[0]/P0001  & n4298 ;
  assign n5690 = ~n5688 & ~n5689 ;
  assign n5691 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5690 ;
  assign n5684 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[8]/P0001  ;
  assign n5692 = reset_n_pad & ~n5684 ;
  assign n5693 = ~n5691 & n5692 ;
  assign n5753 = ~n915 & ~n1353 ;
  assign n5754 = ~n977 & n5753 ;
  assign n5755 = n857 & ~n5754 ;
  assign n5713 = ~\i_tv80_core_IR_reg[3]/P0001  & n1383 ;
  assign n5714 = ~n905 & ~n5713 ;
  assign n5756 = ~n1412 & n5714 ;
  assign n5757 = ~n5755 & n5756 ;
  assign n5745 = n1487 & n1573 ;
  assign n5746 = ~n1170 & ~n1358 ;
  assign n5747 = ~n4773 & n5746 ;
  assign n5748 = ~n5745 & n5747 ;
  assign n5749 = \i_tv80_core_IR_reg[3]/P0001  & ~n5748 ;
  assign n5736 = \i_tv80_core_mcycle_reg[0]/P0001  & ~n675 ;
  assign n5735 = ~\i_tv80_core_mcycle_reg[0]/P0001  & n675 ;
  assign n5750 = n4775 & ~n5735 ;
  assign n5751 = ~n2630 & ~n5750 ;
  assign n5752 = ~n5736 & ~n5751 ;
  assign n5758 = ~n5749 & ~n5752 ;
  assign n5759 = n5757 & n5758 ;
  assign n5760 = n382 & ~n5759 ;
  assign n5734 = \i_tv80_core_IR_reg[0]/P0001  & n1430 ;
  assign n5702 = ~n673 & n857 ;
  assign n5703 = n855 & n5702 ;
  assign n5697 = n1309 & n1451 ;
  assign n5737 = ~n5735 & ~n5736 ;
  assign n5738 = n5697 & n5737 ;
  assign n5739 = ~n5703 & ~n5738 ;
  assign n5740 = \i_tv80_core_IR_reg[3]/P0001  & ~n5739 ;
  assign n5707 = n956 & n1034 ;
  assign n5708 = ~n2655 & ~n5707 ;
  assign n5741 = n857 & n1050 ;
  assign n5742 = n5708 & ~n5741 ;
  assign n5743 = ~n5740 & n5742 ;
  assign n5744 = \i_tv80_core_ISet_reg[1]/P0001  & ~n5743 ;
  assign n5761 = ~n5734 & ~n5744 ;
  assign n5762 = ~n5760 & n5761 ;
  assign n5812 = n2754 & ~n5762 ;
  assign n5811 = n3282 & n5762 ;
  assign n5694 = ~\i_tv80_core_mcycle_reg[0]/P0001  & n2630 ;
  assign n5695 = ~n4775 & ~n5694 ;
  assign n5696 = n2994 & ~n5695 ;
  assign n5698 = n676 & n5697 ;
  assign n5699 = ~n1042 & ~n5698 ;
  assign n5700 = \i_tv80_core_ISet_reg[1]/P0001  & ~n5699 ;
  assign n5701 = ~n5696 & ~n5700 ;
  assign n5715 = ~n1171 & ~n1358 ;
  assign n5716 = n4738 & n5702 ;
  assign n5717 = ~n2630 & ~n5716 ;
  assign n5718 = ~n4774 & n5717 ;
  assign n5719 = n5715 & n5718 ;
  assign n5720 = \i_tv80_core_IR_reg[4]/P0001  & ~n5719 ;
  assign n5721 = n620 & n4775 ;
  assign n5723 = ~n857 & n886 ;
  assign n5724 = n951 & ~n5723 ;
  assign n5725 = ~n4777 & ~n5724 ;
  assign n5726 = ~n5721 & n5725 ;
  assign n5722 = n857 & n920 ;
  assign n5727 = n5714 & ~n5722 ;
  assign n5728 = n5726 & n5727 ;
  assign n5729 = ~n5720 & n5728 ;
  assign n5730 = n382 & ~n5729 ;
  assign n5704 = n999 & n5697 ;
  assign n5705 = ~n5703 & ~n5704 ;
  assign n5706 = \i_tv80_core_IR_reg[4]/P0001  & ~n5705 ;
  assign n5709 = ~n1042 & n5708 ;
  assign n5710 = ~n5706 & n5709 ;
  assign n5711 = \i_tv80_core_ISet_reg[1]/P0001  & ~n5710 ;
  assign n5712 = \i_tv80_core_IR_reg[1]/P0001  & n1430 ;
  assign n5731 = ~n5711 & ~n5712 ;
  assign n5732 = ~n5730 & n5731 ;
  assign n5783 = n898 & n1309 ;
  assign n5784 = ~n5722 & ~n5783 ;
  assign n5780 = ~\i_tv80_core_mcycle_reg[0]/P0001  & n977 ;
  assign n5781 = ~n2627 & n5780 ;
  assign n5782 = ~n1412 & ~n5713 ;
  assign n5785 = ~n5781 & n5782 ;
  assign n5786 = n5784 & n5785 ;
  assign n5776 = n2630 & ~n5735 ;
  assign n5777 = ~n4773 & n5715 ;
  assign n5778 = ~n5776 & n5777 ;
  assign n5779 = \i_tv80_core_IR_reg[5]/P0001  & ~n5778 ;
  assign n5775 = n681 & n4775 ;
  assign n5773 = n856 & n915 ;
  assign n5774 = ~n905 & ~n5773 ;
  assign n5787 = ~n4776 & n5774 ;
  assign n5788 = ~n5775 & n5787 ;
  assign n5789 = ~n5779 & n5788 ;
  assign n5790 = n5786 & n5789 ;
  assign n5791 = n382 & ~n5790 ;
  assign n5764 = n624 & n5697 ;
  assign n5765 = ~n5703 & ~n5764 ;
  assign n5766 = \i_tv80_core_IR_reg[5]/P0001  & ~n5765 ;
  assign n5767 = n856 & n1050 ;
  assign n5768 = ~n5707 & ~n5767 ;
  assign n5769 = ~n2655 & n5768 ;
  assign n5770 = ~n5766 & n5769 ;
  assign n5771 = \i_tv80_core_ISet_reg[1]/P0001  & ~n5770 ;
  assign n5772 = \i_tv80_core_IR_reg[2]/P0001  & n1430 ;
  assign n5792 = ~n5771 & ~n5772 ;
  assign n5793 = ~n5791 & n5792 ;
  assign n5794 = ~n5732 & ~n5793 ;
  assign n5813 = n5701 & ~n5794 ;
  assign n5814 = ~n5811 & n5813 ;
  assign n5815 = ~n5812 & n5814 ;
  assign n5733 = ~n5701 & n5732 ;
  assign n5796 = n5733 & n5762 ;
  assign n5797 = n5793 & n5796 ;
  assign n5795 = ~n5762 & n5794 ;
  assign n5763 = n5733 & ~n5762 ;
  assign n5798 = ~\i_tv80_core_IR_reg[0]/P0001  & n868 ;
  assign n5799 = n1108 & n5798 ;
  assign n5800 = ~n5701 & ~n5799 ;
  assign n5801 = ~n5763 & n5800 ;
  assign n5802 = ~n5795 & n5801 ;
  assign n5803 = ~n5797 & n5802 ;
  assign n5804 = \i_tv80_core_BusA_reg[1]/P0001  & n5803 ;
  assign n5805 = \i_tv80_core_SP_reg[9]/P0001  & n5763 ;
  assign n5806 = n5701 & n5762 ;
  assign n5807 = n5794 & n5806 ;
  assign n5808 = \di_reg_reg[1]/P0001  & n5807 ;
  assign n5816 = ~n5805 & ~n5808 ;
  assign n5809 = \i_tv80_core_ACC_reg[1]/P0001  & n5795 ;
  assign n5810 = \i_tv80_core_SP_reg[1]/P0001  & n5797 ;
  assign n5817 = ~n5809 & ~n5810 ;
  assign n5818 = n5816 & n5817 ;
  assign n5819 = ~n5804 & n5818 ;
  assign n5820 = ~n5815 & n5819 ;
  assign n5827 = n3266 & n5762 ;
  assign n5826 = n2770 & ~n5762 ;
  assign n5828 = n5813 & ~n5826 ;
  assign n5829 = ~n5827 & n5828 ;
  assign n5821 = \i_tv80_core_BusA_reg[2]/P0001  & n5803 ;
  assign n5822 = \i_tv80_core_SP_reg[10]/P0001  & n5763 ;
  assign n5823 = \di_reg_reg[2]/P0001  & n5807 ;
  assign n5830 = ~n5822 & ~n5823 ;
  assign n5824 = \i_tv80_core_ACC_reg[2]/P0001  & n5795 ;
  assign n5825 = \i_tv80_core_SP_reg[2]/P0001  & n5797 ;
  assign n5831 = ~n5824 & ~n5825 ;
  assign n5832 = n5830 & n5831 ;
  assign n5833 = ~n5821 & n5832 ;
  assign n5834 = ~n5829 & n5833 ;
  assign n5841 = n2840 & ~n5762 ;
  assign n5840 = n3341 & n5762 ;
  assign n5842 = n5813 & ~n5840 ;
  assign n5843 = ~n5841 & n5842 ;
  assign n5835 = \i_tv80_core_BusA_reg[3]/P0001  & n5803 ;
  assign n5836 = \i_tv80_core_SP_reg[11]/P0001  & n5763 ;
  assign n5837 = \di_reg_reg[3]/P0001  & n5807 ;
  assign n5844 = ~n5836 & ~n5837 ;
  assign n5838 = \i_tv80_core_ACC_reg[3]/P0001  & n5795 ;
  assign n5839 = \i_tv80_core_SP_reg[3]/P0001  & n5797 ;
  assign n5845 = ~n5838 & ~n5839 ;
  assign n5846 = n5844 & n5845 ;
  assign n5847 = ~n5835 & n5846 ;
  assign n5848 = ~n5843 & n5847 ;
  assign n5855 = n2807 & ~n5762 ;
  assign n5854 = n3357 & n5762 ;
  assign n5856 = n5813 & ~n5854 ;
  assign n5857 = ~n5855 & n5856 ;
  assign n5849 = \i_tv80_core_BusA_reg[4]/P0001  & n5803 ;
  assign n5850 = \i_tv80_core_SP_reg[12]/P0001  & n5763 ;
  assign n5851 = \di_reg_reg[4]/P0001  & n5807 ;
  assign n5858 = ~n5850 & ~n5851 ;
  assign n5852 = \i_tv80_core_ACC_reg[4]/P0001  & n5795 ;
  assign n5853 = \i_tv80_core_SP_reg[4]/P0001  & n5797 ;
  assign n5859 = ~n5852 & ~n5853 ;
  assign n5860 = n5858 & n5859 ;
  assign n5861 = ~n5849 & n5860 ;
  assign n5862 = ~n5857 & n5861 ;
  assign n5869 = n2823 & ~n5762 ;
  assign n5868 = n3374 & n5762 ;
  assign n5870 = n5813 & ~n5868 ;
  assign n5871 = ~n5869 & n5870 ;
  assign n5863 = \i_tv80_core_BusA_reg[5]/P0001  & n5803 ;
  assign n5864 = \i_tv80_core_SP_reg[13]/P0001  & n5763 ;
  assign n5865 = \di_reg_reg[5]/P0001  & n5807 ;
  assign n5872 = ~n5864 & ~n5865 ;
  assign n5866 = \i_tv80_core_ACC_reg[5]/P0001  & n5795 ;
  assign n5867 = \i_tv80_core_SP_reg[5]/P0001  & n5797 ;
  assign n5873 = ~n5866 & ~n5867 ;
  assign n5874 = n5872 & n5873 ;
  assign n5875 = ~n5863 & n5874 ;
  assign n5876 = ~n5871 & n5875 ;
  assign n5883 = n2856 & ~n5762 ;
  assign n5882 = n3325 & n5762 ;
  assign n5884 = n5813 & ~n5882 ;
  assign n5885 = ~n5883 & n5884 ;
  assign n5877 = \i_tv80_core_BusA_reg[6]/P0001  & n5803 ;
  assign n5878 = \i_tv80_core_SP_reg[14]/P0001  & n5763 ;
  assign n5879 = \di_reg_reg[6]/P0001  & n5807 ;
  assign n5886 = ~n5878 & ~n5879 ;
  assign n5880 = \i_tv80_core_ACC_reg[6]/P0001  & n5795 ;
  assign n5881 = \i_tv80_core_SP_reg[6]/P0001  & n5797 ;
  assign n5887 = ~n5880 & ~n5881 ;
  assign n5888 = n5886 & n5887 ;
  assign n5889 = ~n5877 & n5888 ;
  assign n5890 = ~n5885 & n5889 ;
  assign n5897 = n2883 & ~n5762 ;
  assign n5896 = n3401 & n5762 ;
  assign n5898 = n5813 & ~n5896 ;
  assign n5899 = ~n5897 & n5898 ;
  assign n5891 = \i_tv80_core_BusA_reg[7]/P0001  & n5803 ;
  assign n5892 = \i_tv80_core_SP_reg[15]/P0001  & n5763 ;
  assign n5893 = \di_reg_reg[7]/P0001  & n5807 ;
  assign n5900 = ~n5892 & ~n5893 ;
  assign n5894 = \i_tv80_core_ACC_reg[7]/P0001  & n5795 ;
  assign n5895 = \i_tv80_core_SP_reg[7]/P0001  & n5797 ;
  assign n5901 = ~n5894 & ~n5895 ;
  assign n5902 = n5900 & n5901 ;
  assign n5903 = ~n5891 & n5902 ;
  assign n5904 = ~n5899 & n5903 ;
  assign n5911 = n3299 & n5762 ;
  assign n5910 = n2788 & ~n5762 ;
  assign n5912 = n5813 & ~n5910 ;
  assign n5913 = ~n5911 & n5912 ;
  assign n5905 = \i_tv80_core_BusA_reg[0]/P0001  & n5803 ;
  assign n5906 = \i_tv80_core_SP_reg[8]/P0001  & n5763 ;
  assign n5907 = \di_reg_reg[0]/P0001  & n5807 ;
  assign n5914 = ~n5906 & ~n5907 ;
  assign n5908 = \i_tv80_core_ACC_reg[0]/P0001  & n5795 ;
  assign n5909 = \i_tv80_core_SP_reg[0]/P0001  & n5797 ;
  assign n5915 = ~n5908 & ~n5909 ;
  assign n5916 = n5914 & n5915 ;
  assign n5917 = ~n5905 & n5916 ;
  assign n5918 = ~n5913 & n5917 ;
  assign n5919 = \i_tv80_core_i_reg_RegsL_reg[0][0]/P0001  & ~n2696 ;
  assign n5920 = n2788 & n2891 ;
  assign n5921 = \i_tv80_core_RegBusA_r_reg[0]/P0001  & n2664 ;
  assign n5922 = ~n4121 & ~n5921 ;
  assign n5923 = ~n5920 & n5922 ;
  assign n5924 = ~n2667 & ~n5923 ;
  assign n5929 = \i_tv80_core_i_reg_RegsL_reg[4][0]/P0001  & n2918 ;
  assign n5930 = \i_tv80_core_i_reg_RegsL_reg[5][0]/P0001  & n2916 ;
  assign n5935 = ~n5929 & ~n5930 ;
  assign n5931 = \i_tv80_core_i_reg_RegsL_reg[7][0]/P0001  & n2904 ;
  assign n5932 = \i_tv80_core_i_reg_RegsL_reg[2][0]/P0001  & n2908 ;
  assign n5936 = ~n5931 & ~n5932 ;
  assign n5937 = n5935 & n5936 ;
  assign n5925 = \i_tv80_core_i_reg_RegsL_reg[6][0]/P0001  & n2920 ;
  assign n5926 = \i_tv80_core_i_reg_RegsL_reg[3][0]/P0001  & n2922 ;
  assign n5933 = ~n5925 & ~n5926 ;
  assign n5927 = \i_tv80_core_i_reg_RegsL_reg[1][0]/P0001  & n2914 ;
  assign n5928 = \i_tv80_core_i_reg_RegsL_reg[0][0]/P0001  & n2911 ;
  assign n5934 = ~n5927 & ~n5928 ;
  assign n5938 = n5933 & n5934 ;
  assign n5939 = n5937 & n5938 ;
  assign n5940 = n2667 & ~n5939 ;
  assign n5941 = ~n5924 & ~n5940 ;
  assign n5942 = n2696 & ~n5941 ;
  assign n5943 = ~n5919 & ~n5942 ;
  assign n5944 = \i_tv80_core_i_reg_RegsL_reg[7][0]/P0001  & ~n2731 ;
  assign n5945 = n2731 & ~n5941 ;
  assign n5946 = ~n5944 & ~n5945 ;
  assign n5947 = \i_tv80_core_i_reg_RegsL_reg[1][0]/P0001  & ~n2741 ;
  assign n5948 = n2741 & ~n5941 ;
  assign n5949 = ~n5947 & ~n5948 ;
  assign n5950 = \i_tv80_core_i_reg_RegsL_reg[2][0]/P0001  & ~n2745 ;
  assign n5951 = n2745 & ~n5941 ;
  assign n5952 = ~n5950 & ~n5951 ;
  assign n5953 = \i_tv80_core_i_reg_RegsL_reg[3][0]/P0001  & ~n2743 ;
  assign n5954 = n2743 & ~n5941 ;
  assign n5955 = ~n5953 & ~n5954 ;
  assign n5956 = \i_tv80_core_i_reg_RegsL_reg[4][0]/P0001  & ~n2733 ;
  assign n5957 = n2733 & ~n5941 ;
  assign n5958 = ~n5956 & ~n5957 ;
  assign n5959 = \i_tv80_core_i_reg_RegsL_reg[5][0]/P0001  & ~n2739 ;
  assign n5960 = n2739 & ~n5941 ;
  assign n5961 = ~n5959 & ~n5960 ;
  assign n5962 = \i_tv80_core_i_reg_RegsL_reg[6][0]/P0001  & ~n2736 ;
  assign n5963 = n2736 & ~n5941 ;
  assign n5964 = ~n5962 & ~n5963 ;
  assign n5967 = \i_tv80_core_TmpAddr_reg[5]/P0001  & ~n4302 ;
  assign n5968 = \i_tv80_core_IR_reg[5]/P0001  & n4302 ;
  assign n5969 = ~n5967 & ~n5968 ;
  assign n5970 = ~n4300 & ~n5969 ;
  assign n5971 = n4300 & n4448 ;
  assign n5972 = ~n5970 & ~n5971 ;
  assign n5973 = ~n5674 & ~n5972 ;
  assign n5966 = \di_reg_reg[5]/P0001  & n5674 ;
  assign n5974 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5966 ;
  assign n5975 = ~n5973 & n5974 ;
  assign n5965 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[5]/P0001  ;
  assign n5976 = reset_n_pad & ~n5965 ;
  assign n5977 = ~n5975 & n5976 ;
  assign n5980 = n3074 & n4300 ;
  assign n5981 = \i_tv80_core_TmpAddr_reg[7]/P0001  & n4303 ;
  assign n5982 = ~n5980 & ~n5981 ;
  assign n5983 = ~n5674 & ~n5982 ;
  assign n5979 = \di_reg_reg[7]/P0001  & n5674 ;
  assign n5984 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5979 ;
  assign n5985 = ~n5983 & n5984 ;
  assign n5978 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[7]/P0001  ;
  assign n5986 = reset_n_pad & ~n5978 ;
  assign n5987 = ~n5985 & n5986 ;
  assign n5988 = \i_tv80_core_Halt_FF_reg/P0001  & n930 ;
  assign n5989 = ~n4396 & n4740 ;
  assign n5990 = n1103 & n5989 ;
  assign n5991 = ~n5988 & ~n5990 ;
  assign n5992 = reset_n_pad & ~n5991 ;
  assign n5993 = ~\i_tv80_core_BusAck_reg/P0001  & n1103 ;
  assign n5994 = ~n1113 & n5993 ;
  assign n5995 = \i_tv80_core_BTR_r_reg/P0001  & reset_n_pad ;
  assign n5996 = ~n5994 & n5995 ;
  assign n5997 = reset_n_pad & n5994 ;
  assign n5998 = ~\i_tv80_core_No_BTR_reg/P0001  & n1005 ;
  assign n5999 = n1128 & n5998 ;
  assign n6000 = n5997 & n5999 ;
  assign n6001 = ~n5996 & ~n6000 ;
  assign n6008 = n4300 & ~n4580 ;
  assign n6005 = \i_tv80_core_IR_reg[4]/P0001  & n4302 ;
  assign n6004 = \i_tv80_core_TmpAddr_reg[4]/P0001  & ~n4302 ;
  assign n6006 = ~n4300 & ~n6004 ;
  assign n6007 = ~n6005 & n6006 ;
  assign n6009 = ~n5674 & ~n6007 ;
  assign n6010 = ~n6008 & n6009 ;
  assign n6003 = \di_reg_reg[4]/P0001  & n5674 ;
  assign n6011 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6003 ;
  assign n6012 = ~n6010 & n6011 ;
  assign n6002 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[4]/P0001  ;
  assign n6013 = reset_n_pad & ~n6002 ;
  assign n6014 = ~n6012 & n6013 ;
  assign n6021 = n4300 & ~n5566 ;
  assign n6018 = \i_tv80_core_IR_reg[3]/P0001  & n4302 ;
  assign n6017 = \i_tv80_core_TmpAddr_reg[3]/P0001  & ~n4302 ;
  assign n6019 = ~n4300 & ~n6017 ;
  assign n6020 = ~n6018 & n6019 ;
  assign n6022 = ~n5674 & ~n6020 ;
  assign n6023 = ~n6021 & n6022 ;
  assign n6016 = \di_reg_reg[3]/P0001  & n5674 ;
  assign n6024 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6016 ;
  assign n6025 = ~n6023 & n6024 ;
  assign n6015 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[3]/P0001  ;
  assign n6026 = reset_n_pad & ~n6015 ;
  assign n6027 = ~n6025 & n6026 ;
  assign n6028 = \i_tv80_core_BusAck_reg/P0001  & reset_n_pad ;
  assign n6029 = \i_tv80_core_Read_To_Reg_r_reg[4]/P0001  & n6028 ;
  assign n6030 = n857 & n1354 ;
  assign n6037 = n377 & n860 ;
  assign n6038 = n5774 & ~n6037 ;
  assign n6039 = ~n6030 & n6038 ;
  assign n6040 = n4778 & n5719 ;
  assign n6041 = n6039 & n6040 ;
  assign n6042 = n5786 & n6041 ;
  assign n6043 = n382 & ~n6042 ;
  assign n6052 = n860 & n1006 ;
  assign n6053 = n5768 & ~n6052 ;
  assign n6054 = \i_tv80_core_IR_reg[3]/P0001  & n5697 ;
  assign n6055 = ~n5703 & ~n6054 ;
  assign n6056 = n6053 & n6055 ;
  assign n6057 = \i_tv80_core_ISet_reg[1]/P0001  & ~n6056 ;
  assign n6031 = ~n860 & ~n6030 ;
  assign n6032 = n5724 & ~n6031 ;
  assign n6033 = ~n950 & ~n5723 ;
  assign n6034 = n1015 & n6033 ;
  assign n6035 = ~n6032 & ~n6034 ;
  assign n6036 = n1430 & ~n6035 ;
  assign n6045 = ~n1076 & ~n1401 ;
  assign n6046 = n857 & ~n6045 ;
  assign n6044 = n1360 & n1481 ;
  assign n6047 = n879 & n956 ;
  assign n6048 = ~n6044 & ~n6047 ;
  assign n6049 = ~n6046 & n6048 ;
  assign n6050 = n382 & ~n6049 ;
  assign n6051 = ~n5799 & ~n6050 ;
  assign n6058 = ~n6036 & n6051 ;
  assign n6059 = ~n6057 & n6058 ;
  assign n6060 = ~n6043 & n6059 ;
  assign n6061 = reset_n_pad & ~n6060 ;
  assign n6062 = n5993 & n6061 ;
  assign n6063 = ~n6029 & ~n6062 ;
  assign n6066 = n4300 & n5624 ;
  assign n6067 = \i_tv80_core_TmpAddr_reg[2]/P0001  & n4303 ;
  assign n6068 = ~n6066 & ~n6067 ;
  assign n6069 = ~n5674 & ~n6068 ;
  assign n6065 = \di_reg_reg[2]/P0001  & n5674 ;
  assign n6070 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6065 ;
  assign n6071 = ~n6069 & n6070 ;
  assign n6064 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[2]/P0001  ;
  assign n6072 = reset_n_pad & ~n6064 ;
  assign n6073 = ~n6071 & n6072 ;
  assign n6074 = \i_tv80_core_Read_To_Reg_r_reg[0]/P0001  & n6028 ;
  assign n6075 = n5762 & n6051 ;
  assign n6076 = reset_n_pad & ~n6075 ;
  assign n6077 = n5993 & n6076 ;
  assign n6078 = ~n6074 & ~n6077 ;
  assign n6080 = n5993 & ~n6051 ;
  assign n6079 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_Read_To_Reg_r_reg[2]/P0001  ;
  assign n6081 = ~\i_tv80_core_BusAck_reg/P0001  & ~n5793 ;
  assign n6082 = n1103 & n6081 ;
  assign n6083 = ~n6079 & ~n6082 ;
  assign n6084 = ~n6080 & n6083 ;
  assign n6085 = reset_n_pad & ~n6084 ;
  assign n6086 = ~n5732 & n5993 ;
  assign n6087 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_Read_To_Reg_r_reg[1]/P0001  ;
  assign n6088 = ~n6080 & ~n6087 ;
  assign n6089 = ~n6086 & n6088 ;
  assign n6090 = reset_n_pad & ~n6089 ;
  assign n6093 = n4300 & n5604 ;
  assign n6094 = \i_tv80_core_TmpAddr_reg[1]/P0001  & n4303 ;
  assign n6095 = ~n6093 & ~n6094 ;
  assign n6096 = ~n5674 & ~n6095 ;
  assign n6092 = \di_reg_reg[1]/P0001  & n5674 ;
  assign n6097 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6092 ;
  assign n6098 = ~n6096 & n6097 ;
  assign n6091 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[1]/P0001  ;
  assign n6099 = reset_n_pad & ~n6091 ;
  assign n6100 = ~n6098 & n6099 ;
  assign n6101 = ~n4396 & ~n4407 ;
  assign n6102 = reset_n_pad & ~n6101 ;
  assign n6103 = \i_tv80_core_Auto_Wait_t1_reg/P0001  & reset_n_pad ;
  assign n6104 = \i_tv80_core_Read_To_Reg_r_reg[3]/P0001  & n6028 ;
  assign n6105 = ~\i_tv80_core_BusAck_reg/P0001  & reset_n_pad ;
  assign n6106 = ~n5701 & n6105 ;
  assign n6107 = n6051 & n6106 ;
  assign n6108 = n1103 & n6107 ;
  assign n6109 = ~n6104 & ~n6108 ;
  assign n6110 = \i_tv80_core_Save_ALU_r_reg/P0001  & n6028 ;
  assign n6114 = ~n1358 & ~n5722 ;
  assign n6115 = ~n4777 & n5782 ;
  assign n6116 = n6039 & n6115 ;
  assign n6117 = n6114 & n6116 ;
  assign n6118 = n382 & ~n6117 ;
  assign n6111 = ~n1042 & ~n2712 ;
  assign n6112 = n6053 & n6111 ;
  assign n6113 = \i_tv80_core_ISet_reg[1]/P0001  & ~n6112 ;
  assign n6119 = ~n6036 & ~n6113 ;
  assign n6120 = ~n6118 & n6119 ;
  assign n6121 = n5997 & ~n6120 ;
  assign n6122 = ~n6110 & ~n6121 ;
  assign n6123 = \i_tv80_core_ALU_Op_r_reg[3]/P0001  & n6028 ;
  assign n6125 = ~n951 & n6033 ;
  assign n6126 = ~n6032 & ~n6125 ;
  assign n6127 = n1430 & ~n6126 ;
  assign n6124 = \i_tv80_core_ISet_reg[1]/P0001  & n5707 ;
  assign n6128 = n382 & ~n5714 ;
  assign n6129 = ~n6124 & ~n6128 ;
  assign n6130 = ~n6127 & n6129 ;
  assign n6131 = n5997 & ~n6130 ;
  assign n6132 = ~n6123 & ~n6131 ;
  assign n6133 = \i_tv80_core_ALU_Op_r_reg[1]/P0001  & n6028 ;
  assign n6138 = ~\i_tv80_core_IR_reg[4]/P0001  & ~n857 ;
  assign n6139 = ~\i_tv80_core_IR_reg[7]/P0001  & n857 ;
  assign n6140 = ~n6138 & ~n6139 ;
  assign n6141 = n886 & ~n6140 ;
  assign n6134 = ~\i_tv80_core_IR_reg[4]/P0001  & ~n860 ;
  assign n6135 = ~\i_tv80_core_IR_reg[7]/P0001  & n860 ;
  assign n6136 = ~n6134 & ~n6135 ;
  assign n6137 = ~n886 & ~n6136 ;
  assign n6142 = n1430 & ~n6137 ;
  assign n6143 = ~n6141 & n6142 ;
  assign n6151 = ~n1080 & n1349 ;
  assign n6152 = n1373 & n4765 ;
  assign n6153 = n6151 & n6152 ;
  assign n6148 = ~n1078 & ~n1360 ;
  assign n6149 = n1538 & n6148 ;
  assign n6146 = ~n887 & ~n1076 ;
  assign n6147 = ~n1402 & n6146 ;
  assign n6150 = n949 & n6147 ;
  assign n6154 = n6149 & n6150 ;
  assign n6155 = n1341 & n1532 ;
  assign n6156 = n6154 & n6155 ;
  assign n6157 = n6153 & n6156 ;
  assign n6144 = ~n1401 & ~n1403 ;
  assign n6145 = n1370 & n6144 ;
  assign n6165 = ~n1374 & ~n1378 ;
  assign n6164 = ~n1065 & ~n1407 ;
  assign n6166 = ~n1069 & ~n1375 ;
  assign n6167 = n6164 & n6166 ;
  assign n6168 = n6165 & n6167 ;
  assign n6169 = n6145 & n6168 ;
  assign n6158 = ~n974 & n1416 ;
  assign n6159 = n4762 & n6158 ;
  assign n6161 = n1352 & ~n1354 ;
  assign n6160 = ~n856 & n915 ;
  assign n6162 = ~n1171 & ~n6160 ;
  assign n6163 = n6161 & n6162 ;
  assign n6170 = n6159 & n6163 ;
  assign n6171 = n6169 & n6170 ;
  assign n6172 = n6157 & n6171 ;
  assign n6173 = \i_tv80_core_IR_reg[4]/P0001  & ~n6172 ;
  assign n6177 = n921 & ~n6138 ;
  assign n6175 = ~\i_tv80_core_IR_reg[1]/P0001  & ~n857 ;
  assign n6176 = n1490 & n6175 ;
  assign n6174 = \i_tv80_core_IR_reg[0]/P0001  & n1358 ;
  assign n6178 = ~n377 & ~n1384 ;
  assign n6179 = ~n1380 & n6178 ;
  assign n6180 = ~n6174 & n6179 ;
  assign n6181 = ~n6176 & n6180 ;
  assign n6182 = ~n6177 & n6181 ;
  assign n6183 = ~n6173 & n6182 ;
  assign n6184 = ~\i_tv80_core_ISet_reg[0]/NET0131  & ~n6183 ;
  assign n6185 = ~\i_tv80_core_ISet_reg[1]/P0001  & ~n6184 ;
  assign n6190 = n1018 & ~n1033 ;
  assign n6191 = ~n995 & ~n1440 ;
  assign n6192 = n6190 & n6191 ;
  assign n6195 = ~n1014 & ~n1036 ;
  assign n6196 = ~n992 & n6195 ;
  assign n6197 = n1041 & n6196 ;
  assign n6193 = ~n856 & n1050 ;
  assign n6194 = \i_tv80_core_IR_reg[3]/P0001  & n6193 ;
  assign n6198 = ~n1467 & ~n6194 ;
  assign n6199 = n6197 & n6198 ;
  assign n6200 = n6192 & n6199 ;
  assign n6201 = \i_tv80_core_IR_reg[4]/P0001  & ~n6200 ;
  assign n6187 = n375 & n1049 ;
  assign n6188 = n5768 & ~n6187 ;
  assign n6189 = ~\i_tv80_core_IR_reg[3]/P0001  & ~n6188 ;
  assign n6186 = n1006 & ~n6134 ;
  assign n6202 = \i_tv80_core_ISet_reg[1]/P0001  & ~n1010 ;
  assign n6203 = ~n6186 & n6202 ;
  assign n6204 = n6111 & n6203 ;
  assign n6205 = ~n6189 & n6204 ;
  assign n6206 = ~n6201 & n6205 ;
  assign n6207 = ~n6185 & ~n6206 ;
  assign n6208 = ~n6143 & ~n6207 ;
  assign n6209 = n5997 & ~n6208 ;
  assign n6210 = ~n6133 & ~n6209 ;
  assign n6211 = \i_tv80_core_ALU_Op_r_reg[2]/NET0131  & n6028 ;
  assign n6212 = ~n1361 & n6164 ;
  assign n6213 = n6145 & n6212 ;
  assign n6214 = n6157 & n6213 ;
  assign n6215 = ~n1364 & n6159 ;
  assign n6216 = n997 & n1016 ;
  assign n6217 = n1376 & ~n6216 ;
  assign n6218 = ~n1380 & n6217 ;
  assign n6219 = n6165 & n6218 ;
  assign n6220 = n6163 & n6219 ;
  assign n6221 = n6215 & n6220 ;
  assign n6222 = n6214 & n6221 ;
  assign n6223 = \i_tv80_core_IR_reg[5]/P0001  & ~n6222 ;
  assign n6224 = ~n857 & ~n902 ;
  assign n6225 = n920 & n6224 ;
  assign n6226 = ~n6223 & ~n6225 ;
  assign n6227 = n382 & ~n6226 ;
  assign n6229 = ~n855 & ~n1467 ;
  assign n6233 = n1041 & ~n6193 ;
  assign n6234 = n1011 & n6233 ;
  assign n6230 = \i_tv80_core_IR_reg[0]/P0001  & n1036 ;
  assign n6231 = ~n1014 & ~n1037 ;
  assign n6232 = ~n6230 & n6231 ;
  assign n6235 = n6190 & n6232 ;
  assign n6236 = n6234 & n6235 ;
  assign n6237 = n6229 & n6236 ;
  assign n6238 = \i_tv80_core_IR_reg[5]/P0001  & ~n6237 ;
  assign n6228 = ~n860 & n1006 ;
  assign n6239 = n1468 & ~n6228 ;
  assign n6240 = ~n6238 & n6239 ;
  assign n6241 = \i_tv80_core_ISet_reg[1]/P0001  & ~n6240 ;
  assign n6242 = \i_tv80_core_IR_reg[5]/P0001  & n1430 ;
  assign n6243 = ~n6033 & n6242 ;
  assign n6244 = ~n6241 & ~n6243 ;
  assign n6245 = ~n6227 & n6244 ;
  assign n6246 = n5997 & ~n6245 ;
  assign n6247 = ~n6211 & ~n6246 ;
  assign n6248 = \i_tv80_core_ALU_Op_r_reg[0]/P0001  & n6028 ;
  assign n6249 = ~n1170 & n1376 ;
  assign n6250 = n1388 & n6249 ;
  assign n6251 = n6161 & n6250 ;
  assign n6252 = n6215 & n6251 ;
  assign n6253 = n6214 & n6252 ;
  assign n6254 = \i_tv80_core_IR_reg[3]/P0001  & ~n6253 ;
  assign n6255 = ~\i_tv80_core_IR_reg[3]/P0001  & ~n856 ;
  assign n6256 = ~n857 & ~n6255 ;
  assign n6257 = n915 & n6256 ;
  assign n6258 = ~n6254 & ~n6257 ;
  assign n6259 = n382 & ~n6258 ;
  assign n6260 = ~n1034 & ~n1451 ;
  assign n6261 = ~n6228 & n6260 ;
  assign n6262 = n6232 & n6261 ;
  assign n6263 = n6229 & n6262 ;
  assign n6264 = n6192 & n6263 ;
  assign n6265 = \i_tv80_core_IR_reg[3]/P0001  & ~n6264 ;
  assign n6266 = n1050 & ~n6255 ;
  assign n6267 = ~n1000 & ~n1010 ;
  assign n6268 = ~n6266 & n6267 ;
  assign n6269 = ~n2712 & n6268 ;
  assign n6270 = ~n6265 & n6269 ;
  assign n6271 = \i_tv80_core_ISet_reg[1]/P0001  & ~n6270 ;
  assign n6272 = \i_tv80_core_IR_reg[3]/P0001  & ~n6125 ;
  assign n6273 = n989 & n6033 ;
  assign n6274 = ~n6272 & ~n6273 ;
  assign n6275 = ~n6032 & n6274 ;
  assign n6276 = n1430 & ~n6275 ;
  assign n6277 = ~n6271 & ~n6276 ;
  assign n6278 = ~n6259 & n6277 ;
  assign n6279 = n5997 & ~n6278 ;
  assign n6280 = ~n6248 & ~n6279 ;
  assign n6281 = n4390 & ~n4392 ;
  assign n6282 = reset_n_pad & ~n6281 ;
  assign n6283 = ~n1103 & n6282 ;
  assign n6284 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_RegAddrC_reg[1]/NET0131  ;
  assign n6285 = ~n1277 & ~n2997 ;
  assign n6286 = ~\i_tv80_core_BusAck_reg/P0001  & n6285 ;
  assign n6287 = n1529 & n6286 ;
  assign n6288 = ~n6284 & ~n6287 ;
  assign n6289 = ~n1430 & n4594 ;
  assign n6290 = \i_tv80_core_IR_reg[0]/P0001  & ~n6289 ;
  assign n6291 = n1036 & n2715 ;
  assign n6292 = \i_tv80_core_IR_reg[3]/P0001  & n6291 ;
  assign n6298 = ~n1042 & ~n6292 ;
  assign n6293 = n675 & n1481 ;
  assign n6294 = n856 & n5736 ;
  assign n6295 = ~n6293 & ~n6294 ;
  assign n6296 = n1008 & ~n6295 ;
  assign n6297 = n5737 & n5767 ;
  assign n6299 = ~n6296 & ~n6297 ;
  assign n6300 = n6298 & n6299 ;
  assign n6301 = \i_tv80_core_ISet_reg[1]/P0001  & ~n6300 ;
  assign n6303 = ~n871 & ~n910 ;
  assign n6304 = ~n970 & n974 ;
  assign n6305 = n6303 & ~n6304 ;
  assign n6306 = \i_tv80_core_mcycle_reg[0]/P0001  & ~n6305 ;
  assign n6307 = n915 & n5737 ;
  assign n6308 = ~n5780 & ~n6307 ;
  assign n6309 = ~n6306 & n6308 ;
  assign n6310 = n856 & ~n6309 ;
  assign n6311 = n860 & n1080 ;
  assign n6312 = ~n1171 & ~n1412 ;
  assign n6313 = ~n6311 & n6312 ;
  assign n6314 = \i_tv80_core_IR_reg[0]/P0001  & ~n6313 ;
  assign n6317 = n860 & ~n1404 ;
  assign n6316 = n894 & n956 ;
  assign n6318 = ~n4772 & ~n6316 ;
  assign n6319 = ~n6317 & n6318 ;
  assign n6302 = n860 & ~n2632 ;
  assign n6315 = n2620 & ~n5736 ;
  assign n6320 = ~n6302 & ~n6315 ;
  assign n6321 = n6319 & n6320 ;
  assign n6322 = ~n6314 & n6321 ;
  assign n6323 = ~n6310 & n6322 ;
  assign n6324 = n382 & ~n6323 ;
  assign n6325 = ~n6301 & ~n6324 ;
  assign n6326 = n4594 & ~n6325 ;
  assign n6327 = ~n6290 & ~n6326 ;
  assign n6355 = \i_tv80_core_IR_reg[2]/P0001  & ~n4594 ;
  assign n6343 = ~n2620 & ~n5773 ;
  assign n6363 = ~\i_tv80_core_IR_reg[4]/P0001  & ~n6343 ;
  assign n6364 = n860 & n948 ;
  assign n6365 = ~n6363 & ~n6364 ;
  assign n6366 = \i_tv80_core_IR_reg[5]/P0001  & ~n6365 ;
  assign n6367 = ~n1482 & ~n6303 ;
  assign n6373 = ~n5781 & ~n6030 ;
  assign n6374 = ~n6367 & n6373 ;
  assign n6375 = n6319 & n6374 ;
  assign n6376 = ~n6366 & n6375 ;
  assign n6368 = ~n2626 & ~n2633 ;
  assign n6369 = ~n887 & ~n1335 ;
  assign n6370 = n857 & ~n6369 ;
  assign n6371 = n6313 & ~n6370 ;
  assign n6372 = \i_tv80_core_IR_reg[2]/P0001  & ~n6371 ;
  assign n6377 = n6368 & ~n6372 ;
  assign n6378 = n6376 & n6377 ;
  assign n6379 = n382 & ~n6378 ;
  assign n6329 = n1008 & ~n1482 ;
  assign n6330 = ~n5767 & ~n6329 ;
  assign n6356 = ~\i_tv80_core_IR_reg[4]/P0001  & ~n6330 ;
  assign n6357 = ~n6291 & ~n6356 ;
  assign n6358 = \i_tv80_core_IR_reg[5]/P0001  & ~n6357 ;
  assign n6359 = n857 & n1006 ;
  assign n6360 = n5709 & ~n6359 ;
  assign n6361 = ~n6358 & n6360 ;
  assign n6362 = \i_tv80_core_ISet_reg[1]/P0001  & ~n6361 ;
  assign n6380 = ~n5772 & ~n6362 ;
  assign n6381 = ~n6379 & n6380 ;
  assign n6382 = n4594 & ~n6381 ;
  assign n6383 = ~n6355 & ~n6382 ;
  assign n6339 = n857 & n1490 ;
  assign n6340 = n6313 & ~n6339 ;
  assign n6341 = \i_tv80_core_IR_reg[1]/P0001  & ~n6340 ;
  assign n6338 = ~n6037 & n6114 ;
  assign n6342 = \i_tv80_core_IR_reg[5]/P0001  & ~n2620 ;
  assign n6344 = \i_tv80_core_IR_reg[4]/P0001  & ~n6342 ;
  assign n6345 = ~n6343 & n6344 ;
  assign n6346 = ~n4776 & n6319 ;
  assign n6347 = ~n6345 & n6346 ;
  assign n6348 = n6338 & n6347 ;
  assign n6349 = ~n6341 & n6348 ;
  assign n6350 = n382 & ~n6349 ;
  assign n6331 = ~\i_tv80_core_IR_reg[5]/P0001  & ~n6330 ;
  assign n6332 = ~n6291 & ~n6331 ;
  assign n6333 = \i_tv80_core_IR_reg[4]/P0001  & ~n6332 ;
  assign n6334 = n381 & n1006 ;
  assign n6335 = n5709 & ~n6334 ;
  assign n6336 = ~n6333 & n6335 ;
  assign n6337 = \i_tv80_core_ISet_reg[1]/P0001  & ~n6336 ;
  assign n6351 = ~n5712 & ~n6337 ;
  assign n6352 = ~n6350 & n6351 ;
  assign n6387 = n675 & n5773 ;
  assign n6388 = ~n2619 & ~n6387 ;
  assign n6389 = n6338 & n6388 ;
  assign n6390 = n6368 & n6389 ;
  assign n6391 = n382 & ~n6390 ;
  assign n6385 = n857 & n2994 ;
  assign n6386 = n948 & n6385 ;
  assign n6392 = n675 & ~n6330 ;
  assign n6393 = n673 & n6291 ;
  assign n6394 = ~n6052 & ~n6393 ;
  assign n6395 = ~n6392 & n6394 ;
  assign n6396 = \i_tv80_core_ISet_reg[1]/P0001  & ~n6395 ;
  assign n6397 = ~n6386 & ~n6396 ;
  assign n6398 = ~n6391 & n6397 ;
  assign n6399 = n4594 & ~n6398 ;
  assign n6418 = n6352 & n6399 ;
  assign n6419 = ~n6383 & n6418 ;
  assign n6422 = n6327 & n6419 ;
  assign n6423 = \i_tv80_core_PC_reg[0]/P0001  & n6422 ;
  assign n6328 = \i_tv80_core_IR_reg[1]/P0001  & ~n4594 ;
  assign n6353 = n4594 & ~n6352 ;
  assign n6354 = ~n6328 & ~n6353 ;
  assign n6413 = ~\i_tv80_core_SP_reg[0]/P0001  & n6354 ;
  assign n6409 = n6381 & n6399 ;
  assign n6414 = n6327 & n6409 ;
  assign n6415 = ~n6413 & n6414 ;
  assign n6420 = ~n6327 & n6419 ;
  assign n6421 = \i_tv80_core_PC_reg[8]/P0001  & n6420 ;
  assign n6425 = ~n6415 & ~n6421 ;
  assign n6426 = ~n6423 & n6425 ;
  assign n6384 = ~n6354 & ~n6383 ;
  assign n6400 = n6384 & ~n6399 ;
  assign n6401 = ~n6327 & n6400 ;
  assign n6402 = \i_tv80_core_ACC_reg[0]/P0001  & n6401 ;
  assign n6403 = \i_tv80_core_F_reg[0]/P0001  & n6386 ;
  assign n6410 = n6354 & n6409 ;
  assign n6411 = ~n6327 & n6410 ;
  assign n6412 = \i_tv80_core_SP_reg[8]/P0001  & n6411 ;
  assign n6424 = ~n6403 & ~n6412 ;
  assign n6427 = ~n6402 & n6424 ;
  assign n6406 = n4112 & n6327 ;
  assign n6404 = ~n6384 & ~n6399 ;
  assign n6405 = n5939 & ~n6327 ;
  assign n6407 = n6404 & ~n6405 ;
  assign n6408 = ~n6406 & n6407 ;
  assign n6416 = n6327 & n6400 ;
  assign n6417 = \di_reg_reg[0]/P0001  & n6416 ;
  assign n6428 = ~n6408 & ~n6417 ;
  assign n6429 = n6427 & n6428 ;
  assign n6430 = n6426 & n6429 ;
  assign n6438 = \i_tv80_core_PC_reg[11]/P0001  & n6420 ;
  assign n6434 = \i_tv80_core_SP_reg[11]/P0001  & n6411 ;
  assign n6437 = \i_tv80_core_PC_reg[3]/P0001  & n6422 ;
  assign n6444 = ~n6434 & ~n6437 ;
  assign n6445 = ~n6438 & n6444 ;
  assign n6431 = \i_tv80_core_ACC_reg[3]/P0001  & n6401 ;
  assign n6432 = n6327 & n6410 ;
  assign n6433 = \i_tv80_core_SP_reg[3]/P0001  & n6432 ;
  assign n6435 = \i_tv80_core_F_reg[3]/P0001  & n6386 ;
  assign n6443 = ~n6433 & ~n6435 ;
  assign n6446 = ~n6431 & n6443 ;
  assign n6436 = \di_reg_reg[3]/P0001  & n6416 ;
  assign n6440 = n4015 & n6327 ;
  assign n6439 = n4531 & ~n6327 ;
  assign n6441 = n6404 & ~n6439 ;
  assign n6442 = ~n6440 & n6441 ;
  assign n6447 = ~n6436 & ~n6442 ;
  assign n6448 = n6446 & n6447 ;
  assign n6449 = n6445 & n6448 ;
  assign n6456 = \i_tv80_core_PC_reg[2]/P0001  & n6422 ;
  assign n6452 = \i_tv80_core_SP_reg[10]/P0001  & n6411 ;
  assign n6455 = \i_tv80_core_PC_reg[10]/P0001  & n6420 ;
  assign n6462 = ~n6452 & ~n6455 ;
  assign n6463 = ~n6456 & n6462 ;
  assign n6450 = \di_reg_reg[2]/P0001  & n6416 ;
  assign n6451 = \i_tv80_core_SP_reg[2]/P0001  & n6432 ;
  assign n6453 = \i_tv80_core_F_reg[2]/P0001  & n6386 ;
  assign n6461 = ~n6451 & ~n6453 ;
  assign n6464 = ~n6450 & n6461 ;
  assign n6454 = \i_tv80_core_ACC_reg[2]/P0001  & n6401 ;
  assign n6458 = n3889 & n6327 ;
  assign n6457 = n4688 & ~n6327 ;
  assign n6459 = n6404 & ~n6457 ;
  assign n6460 = ~n6458 & n6459 ;
  assign n6465 = ~n6454 & ~n6460 ;
  assign n6466 = n6464 & n6465 ;
  assign n6467 = n6463 & n6466 ;
  assign n6474 = \i_tv80_core_PC_reg[12]/P0001  & n6420 ;
  assign n6470 = \i_tv80_core_SP_reg[12]/P0001  & n6411 ;
  assign n6473 = \i_tv80_core_PC_reg[4]/P0001  & n6422 ;
  assign n6480 = ~n6470 & ~n6473 ;
  assign n6481 = ~n6474 & n6480 ;
  assign n6468 = \i_tv80_core_ACC_reg[4]/P0001  & n6401 ;
  assign n6469 = \i_tv80_core_SP_reg[4]/P0001  & n6432 ;
  assign n6471 = \i_tv80_core_F_reg[4]/P0001  & n6386 ;
  assign n6479 = ~n6469 & ~n6471 ;
  assign n6482 = ~n6468 & n6479 ;
  assign n6472 = \di_reg_reg[4]/P0001  & n6416 ;
  assign n6476 = n3688 & n6327 ;
  assign n6475 = n4358 & ~n6327 ;
  assign n6477 = n6404 & ~n6475 ;
  assign n6478 = ~n6476 & n6477 ;
  assign n6483 = ~n6472 & ~n6478 ;
  assign n6484 = n6482 & n6483 ;
  assign n6485 = n6481 & n6484 ;
  assign n6492 = \i_tv80_core_PC_reg[13]/P0001  & n6420 ;
  assign n6488 = \i_tv80_core_SP_reg[5]/P0001  & n6432 ;
  assign n6491 = \i_tv80_core_PC_reg[5]/P0001  & n6422 ;
  assign n6498 = ~n6488 & ~n6491 ;
  assign n6499 = ~n6492 & n6498 ;
  assign n6486 = \i_tv80_core_ACC_reg[5]/P0001  & n6401 ;
  assign n6487 = \i_tv80_core_SP_reg[13]/P0001  & n6411 ;
  assign n6489 = \i_tv80_core_F_reg[5]/P0001  & n6386 ;
  assign n6497 = ~n6487 & ~n6489 ;
  assign n6500 = ~n6486 & n6497 ;
  assign n6490 = \di_reg_reg[5]/P0001  & n6416 ;
  assign n6494 = n3630 & n6327 ;
  assign n6493 = n4267 & ~n6327 ;
  assign n6495 = n6404 & ~n6493 ;
  assign n6496 = ~n6494 & n6495 ;
  assign n6501 = ~n6490 & ~n6496 ;
  assign n6502 = n6500 & n6501 ;
  assign n6503 = n6499 & n6502 ;
  assign n6510 = \i_tv80_core_PC_reg[14]/P0001  & n6420 ;
  assign n6506 = \i_tv80_core_SP_reg[14]/P0001  & n6411 ;
  assign n6509 = \i_tv80_core_PC_reg[6]/P0001  & n6422 ;
  assign n6516 = ~n6506 & ~n6509 ;
  assign n6517 = ~n6510 & n6516 ;
  assign n6504 = \di_reg_reg[6]/P0001  & n6416 ;
  assign n6505 = \i_tv80_core_SP_reg[6]/P0001  & n6432 ;
  assign n6507 = \i_tv80_core_F_reg[6]/P0001  & n6386 ;
  assign n6515 = ~n6505 & ~n6507 ;
  assign n6518 = ~n6504 & n6515 ;
  assign n6508 = \i_tv80_core_ACC_reg[6]/P0001  & n6401 ;
  assign n6512 = n3496 & n6327 ;
  assign n6511 = n3543 & ~n6327 ;
  assign n6513 = n6404 & ~n6511 ;
  assign n6514 = ~n6512 & n6513 ;
  assign n6519 = ~n6508 & ~n6514 ;
  assign n6520 = n6518 & n6519 ;
  assign n6521 = n6517 & n6520 ;
  assign n6528 = \i_tv80_core_PC_reg[7]/P0001  & n6422 ;
  assign n6524 = \i_tv80_core_SP_reg[15]/P0001  & n6411 ;
  assign n6527 = \i_tv80_core_PC_reg[15]/P0001  & n6420 ;
  assign n6534 = ~n6524 & ~n6527 ;
  assign n6535 = ~n6528 & n6534 ;
  assign n6522 = \di_reg_reg[7]/P0001  & n6416 ;
  assign n6523 = \i_tv80_core_SP_reg[7]/P0001  & n6432 ;
  assign n6525 = \i_tv80_core_F_reg[7]/P0001  & n6386 ;
  assign n6533 = ~n6523 & ~n6525 ;
  assign n6536 = ~n6522 & n6533 ;
  assign n6526 = \i_tv80_core_ACC_reg[7]/P0001  & n6401 ;
  assign n6530 = n3427 & n6327 ;
  assign n6529 = n2930 & ~n6327 ;
  assign n6531 = n6404 & ~n6529 ;
  assign n6532 = ~n6530 & n6531 ;
  assign n6537 = ~n6526 & ~n6532 ;
  assign n6538 = n6536 & n6537 ;
  assign n6539 = n6535 & n6538 ;
  assign n6546 = \i_tv80_core_PC_reg[9]/P0001  & n6420 ;
  assign n6542 = \i_tv80_core_SP_reg[9]/P0001  & n6411 ;
  assign n6545 = \i_tv80_core_PC_reg[1]/P0001  & n6422 ;
  assign n6552 = ~n6542 & ~n6545 ;
  assign n6553 = ~n6546 & n6552 ;
  assign n6540 = \i_tv80_core_ACC_reg[1]/P0001  & n6401 ;
  assign n6541 = \i_tv80_core_SP_reg[1]/P0001  & n6432 ;
  assign n6543 = \i_tv80_core_F_reg[1]/P0001  & n6386 ;
  assign n6551 = ~n6541 & ~n6543 ;
  assign n6554 = ~n6540 & n6551 ;
  assign n6544 = \di_reg_reg[1]/P0001  & n6416 ;
  assign n6548 = n4059 & n6327 ;
  assign n6547 = n5533 & ~n6327 ;
  assign n6549 = n6404 & ~n6547 ;
  assign n6550 = ~n6548 & n6549 ;
  assign n6555 = ~n6544 & ~n6550 ;
  assign n6556 = n6554 & n6555 ;
  assign n6557 = n6553 & n6556 ;
  assign n6558 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_RegAddrC_reg[0]/P0001  ;
  assign n6559 = ~n1593 & ~n6285 ;
  assign n6560 = ~n862 & ~n6559 ;
  assign n6561 = n1570 & n6285 ;
  assign n6562 = n6560 & ~n6561 ;
  assign n6563 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6562 ;
  assign n6564 = ~n6558 & ~n6563 ;
  assign n6566 = ~\i_tv80_core_mcycle_reg[0]/P0001  & n1404 ;
  assign n6567 = ~n1080 & n6566 ;
  assign n6568 = ~n876 & n919 ;
  assign n6569 = \i_tv80_core_mcycle_reg[0]/P0001  & ~n1350 ;
  assign n6570 = ~n6568 & n6569 ;
  assign n6571 = ~n6567 & ~n6570 ;
  assign n6572 = ~n948 & n2632 ;
  assign n6573 = ~n6571 & n6572 ;
  assign n6574 = n856 & ~n6573 ;
  assign n6575 = ~n910 & n1311 ;
  assign n6576 = n1309 & ~n6575 ;
  assign n6565 = n894 & n1481 ;
  assign n6577 = ~n2629 & ~n6565 ;
  assign n6578 = ~n6576 & n6577 ;
  assign n6579 = ~n6574 & n6578 ;
  assign n6580 = n382 & ~n6579 ;
  assign n6581 = ~\i_tv80_core_mcycle_reg[0]/P0001  & n1034 ;
  assign n6582 = ~n1008 & ~n6581 ;
  assign n6583 = n1309 & ~n6582 ;
  assign n6584 = n857 & n6230 ;
  assign n6585 = ~n2642 & ~n6584 ;
  assign n6586 = ~n2654 & n6585 ;
  assign n6587 = ~n6583 & n6586 ;
  assign n6588 = \i_tv80_core_ISet_reg[1]/P0001  & ~n6587 ;
  assign n6589 = n885 & n5712 ;
  assign n6590 = n956 & ~n989 ;
  assign n6591 = n6589 & n6590 ;
  assign n6592 = ~n6588 & ~n6591 ;
  assign n6593 = ~n6580 & n6592 ;
  assign n6597 = ~n4751 & ~n5773 ;
  assign n6598 = n382 & ~n6597 ;
  assign n6603 = n857 & n2974 ;
  assign n6600 = n940 & n956 ;
  assign n6601 = ~n1481 & ~n6600 ;
  assign n6602 = n1005 & ~n6601 ;
  assign n6604 = ~n5767 & ~n6602 ;
  assign n6605 = ~n6603 & n6604 ;
  assign n6606 = \i_tv80_core_ISet_reg[1]/P0001  & ~n6605 ;
  assign n6596 = n1462 & n4787 ;
  assign n6599 = ~n1156 & ~n4395 ;
  assign n6607 = ~n6596 & ~n6599 ;
  assign n6608 = ~n6606 & n6607 ;
  assign n6609 = ~n6598 & n6608 ;
  assign n6610 = n6593 & n6609 ;
  assign n6611 = ~n4390 & n6610 ;
  assign n6594 = n1634 & ~n6593 ;
  assign n6612 = ~n860 & ~n6594 ;
  assign n6613 = ~n6611 & n6612 ;
  assign n6595 = n4390 & n6594 ;
  assign n6614 = \i_tv80_core_IntCycle_reg/P0001  & ~n6599 ;
  assign n6615 = n860 & ~n6614 ;
  assign n6616 = reset_n_pad & ~n6615 ;
  assign n6617 = ~n6595 & n6616 ;
  assign n6618 = ~n6613 & n6617 ;
  assign n6620 = n4390 & n6610 ;
  assign n6621 = n6612 & ~n6620 ;
  assign n6619 = ~n4390 & n6594 ;
  assign n6622 = ~\i_tv80_core_IntCycle_reg/P0001  & ~n6599 ;
  assign n6623 = n2697 & ~n6622 ;
  assign n6624 = reset_n_pad & ~n6623 ;
  assign n6625 = ~n6619 & n6624 ;
  assign n6626 = ~n6621 & n6625 ;
  assign n6627 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_RegAddrB_r_reg[0]/P0001  ;
  assign n6628 = n1598 & ~n6383 ;
  assign n6629 = n6354 & ~n6628 ;
  assign n6630 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6629 ;
  assign n6631 = ~n6627 & ~n6630 ;
  assign n6632 = n6354 & n6628 ;
  assign n6633 = \i_tv80_core_XY_State_reg[1]/P0001  & n6632 ;
  assign n6634 = \i_tv80_core_Alternate_reg/P0001  & ~n6632 ;
  assign n6635 = ~n6633 & ~n6634 ;
  assign n6639 = n917 & n1114 ;
  assign n6640 = ~n973 & ~n6639 ;
  assign n6641 = ~\i_tv80_core_IR_reg[0]/P0001  & ~n6640 ;
  assign n6642 = ~\i_tv80_core_IR_reg[2]/P0001  & ~n620 ;
  assign n6643 = \i_tv80_core_IR_reg[3]/P0001  & ~n681 ;
  assign n6644 = n6642 & ~n6643 ;
  assign n6645 = ~\i_tv80_core_IR_reg[6]/P0001  & ~n6644 ;
  assign n6646 = n374 & n1015 ;
  assign n6647 = ~n6645 & n6646 ;
  assign n6648 = ~n6641 & ~n6647 ;
  assign n6657 = \i_tv80_core_IR_reg[2]/P0001  & ~n952 ;
  assign n6658 = ~\i_tv80_core_IR_reg[7]/P0001  & n371 ;
  assign n6659 = ~n6657 & ~n6658 ;
  assign n6660 = \i_tv80_core_IR_reg[1]/P0001  & ~n6659 ;
  assign n6661 = ~n867 & ~n6660 ;
  assign n6662 = ~\i_tv80_core_IR_reg[0]/P0001  & ~n6661 ;
  assign n6663 = n628 & n867 ;
  assign n6664 = ~\i_tv80_core_IR_reg[6]/P0001  & n375 ;
  assign n6665 = ~n6663 & ~n6664 ;
  assign n6666 = ~\i_tv80_core_IR_reg[1]/P0001  & ~n6665 ;
  assign n6667 = ~n953 & ~n6666 ;
  assign n6668 = ~\i_tv80_core_IR_reg[2]/P0001  & ~n6667 ;
  assign n6649 = ~n914 & ~n953 ;
  assign n6650 = \i_tv80_core_IR_reg[0]/P0001  & ~n6649 ;
  assign n6654 = ~\i_tv80_core_IR_reg[1]/P0001  & n952 ;
  assign n6651 = \i_tv80_core_IR_reg[1]/P0001  & \i_tv80_core_IR_reg[5]/P0001  ;
  assign n6652 = ~\i_tv80_core_IR_reg[3]/P0001  & n867 ;
  assign n6653 = ~n6651 & n6652 ;
  assign n6655 = \i_tv80_core_IR_reg[7]/P0001  & n993 ;
  assign n6656 = ~n6642 & n6655 ;
  assign n6669 = ~n6653 & ~n6656 ;
  assign n6670 = ~n6654 & n6669 ;
  assign n6671 = ~n1490 & n6670 ;
  assign n6672 = ~n6650 & n6671 ;
  assign n6673 = ~n6668 & n6672 ;
  assign n6674 = ~n6662 & n6673 ;
  assign n6675 = n6648 & ~n6674 ;
  assign n6677 = n944 & ~n1493 ;
  assign n6638 = n971 & n974 ;
  assign n6676 = n6641 & ~n6647 ;
  assign n6637 = \i_tv80_core_NMICycle_reg/P0001  & n929 ;
  assign n6678 = n4748 & ~n6637 ;
  assign n6679 = ~n6676 & n6678 ;
  assign n6680 = ~n6638 & n6679 ;
  assign n6681 = ~n6677 & n6680 ;
  assign n6682 = ~n6675 & n6681 ;
  assign n6683 = n382 & ~n6682 ;
  assign n6684 = ~n876 & ~n885 ;
  assign n6685 = n1108 & n6684 ;
  assign n6686 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6589 ;
  assign n6687 = ~n6685 & n6686 ;
  assign n6688 = ~n6683 & n6687 ;
  assign n6636 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_mcycles_reg[1]/P0001  ;
  assign n6689 = reset_n_pad & ~n6636 ;
  assign n6690 = ~n6688 & n6689 ;
  assign n6692 = n4300 & n5587 ;
  assign n6693 = \i_tv80_core_TmpAddr_reg[0]/P0001  & n4303 ;
  assign n6694 = ~n6692 & ~n6693 ;
  assign n6695 = ~n5674 & n6694 ;
  assign n6696 = ~\di_reg_reg[0]/P0001  & n5674 ;
  assign n6697 = ~n6695 & ~n6696 ;
  assign n6698 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6697 ;
  assign n6691 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_TmpAddr_reg[0]/P0001  ;
  assign n6699 = reset_n_pad & ~n6691 ;
  assign n6700 = ~n6698 & n6699 ;
  assign n6701 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_RegAddrA_r_reg[1]/NET0131  ;
  assign n6702 = ~n6081 & ~n6701 ;
  assign n6703 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_Z16_r_reg/P0001  ;
  assign n6704 = ~\i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_ISet_reg[1]/P0001  ;
  assign n6705 = n1306 & n6704 ;
  assign n6706 = n6245 & n6705 ;
  assign n6707 = ~n6278 & n6706 ;
  assign n6708 = ~n6703 & ~n6707 ;
  assign n6709 = reset_n_pad & ~n6708 ;
  assign n6710 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_RegAddrA_r_reg[0]/NET0131  ;
  assign n6711 = n1598 & ~n5793 ;
  assign n6712 = n5732 & ~n6711 ;
  assign n6713 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6712 ;
  assign n6714 = ~n6710 & ~n6713 ;
  assign n6716 = ~n860 & ~n6610 ;
  assign n6715 = n860 & ~n6622 ;
  assign n6717 = reset_n_pad & ~n6715 ;
  assign n6718 = ~n6716 & n6717 ;
  assign n6719 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6383 ;
  assign n6720 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_RegAddrB_r_reg[1]/P0001  ;
  assign n6721 = ~n6719 & ~n6720 ;
  assign n6722 = n5732 & n6711 ;
  assign n6723 = \i_tv80_core_XY_State_reg[1]/P0001  & n6722 ;
  assign n6724 = \i_tv80_core_Alternate_reg/P0001  & ~n6722 ;
  assign n6725 = ~n6723 & ~n6724 ;
  assign n6726 = n624 & n1111 ;
  assign n6727 = \i_tv80_core_R_reg[0]/P0001  & n5310 ;
  assign n6728 = \i_tv80_core_R_reg[1]/P0001  & n6727 ;
  assign n6729 = \i_tv80_core_R_reg[2]/P0001  & n6728 ;
  assign n6730 = \i_tv80_core_R_reg[3]/P0001  & n6729 ;
  assign n6731 = \i_tv80_core_R_reg[4]/P0001  & n6730 ;
  assign n6732 = ~n6726 & ~n6731 ;
  assign n6733 = ~\i_tv80_core_R_reg[5]/P0001  & ~n6726 ;
  assign n6734 = ~n6732 & ~n6733 ;
  assign n6735 = ~\i_tv80_core_BusAck_reg/P0001  & n6734 ;
  assign n6737 = ~\i_tv80_core_R_reg[6]/P0001  & ~n6726 ;
  assign n6738 = \i_tv80_core_ACC_reg[6]/P0001  & n6726 ;
  assign n6739 = ~n6737 & ~n6738 ;
  assign n6740 = n6735 & n6739 ;
  assign n6736 = ~\i_tv80_core_R_reg[6]/P0001  & ~n6735 ;
  assign n6741 = reset_n_pad & ~n6736 ;
  assign n6742 = ~n6740 & n6741 ;
  assign n6759 = ~\i_tv80_core_F_reg[6]/P0001  & n1339 ;
  assign n6758 = ~\i_tv80_core_F_reg[0]/P0001  & n1374 ;
  assign n6760 = n857 & ~n6758 ;
  assign n6761 = ~n6759 & n6760 ;
  assign n6762 = ~n4748 & ~n6761 ;
  assign n6763 = ~\i_tv80_core_F_reg[0]/P0001  & n857 ;
  assign n6764 = n6676 & ~n6763 ;
  assign n6747 = \i_tv80_core_IR_reg[0]/P0001  & ~\i_tv80_core_IR_reg[6]/P0001  ;
  assign n6748 = n917 & n1038 ;
  assign n6753 = ~n6747 & ~n6748 ;
  assign n6754 = ~n919 & n6753 ;
  assign n6746 = ~n889 & ~n952 ;
  assign n6749 = \i_tv80_core_IR_reg[6]/P0001  & ~n1026 ;
  assign n6750 = ~\i_tv80_core_IR_reg[7]/P0001  & ~n681 ;
  assign n6751 = ~n6749 & n6750 ;
  assign n6752 = ~\i_tv80_core_IR_reg[2]/P0001  & ~n6751 ;
  assign n6755 = ~n6746 & ~n6752 ;
  assign n6756 = n6754 & n6755 ;
  assign n6757 = n6648 & ~n6756 ;
  assign n6765 = \i_tv80_core_F_reg[6]/P0001  & n1338 ;
  assign n6745 = n374 & n867 ;
  assign n6766 = ~n929 & ~n6745 ;
  assign n6767 = ~n6765 & n6766 ;
  assign n6768 = ~n6757 & n6767 ;
  assign n6769 = ~n6764 & n6768 ;
  assign n6770 = ~n6762 & n6769 ;
  assign n6771 = n382 & ~n6770 ;
  assign n6772 = n681 & n1379 ;
  assign n6773 = ~\i_tv80_core_IR_reg[7]/P0001  & ~n853 ;
  assign n6774 = ~n6772 & n6773 ;
  assign n6775 = n1018 & ~n6774 ;
  assign n6776 = \i_tv80_core_ISet_reg[1]/P0001  & ~n6775 ;
  assign n6744 = n1430 & ~n4738 ;
  assign n6777 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6744 ;
  assign n6778 = ~n6776 & n6777 ;
  assign n6779 = ~n6771 & n6778 ;
  assign n6743 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_mcycles_reg[0]/P0001  ;
  assign n6780 = reset_n_pad & ~n6743 ;
  assign n6781 = ~n6779 & n6780 ;
  assign n6784 = ~\i_tv80_core_R_reg[5]/P0001  & ~n6731 ;
  assign n6785 = ~n6734 & ~n6784 ;
  assign n6783 = \i_tv80_core_ACC_reg[5]/P0001  & n6726 ;
  assign n6786 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6783 ;
  assign n6787 = ~n6785 & n6786 ;
  assign n6782 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_R_reg[5]/P0001  ;
  assign n6788 = reset_n_pad & ~n6782 ;
  assign n6789 = ~n6787 & n6788 ;
  assign n6795 = ~\i_tv80_core_BusAck_reg/P0001  & n382 ;
  assign n6796 = ~n971 & n974 ;
  assign n6797 = n852 & n892 ;
  assign n6798 = ~n870 & ~n6797 ;
  assign n6799 = n6648 & ~n6798 ;
  assign n6800 = ~n977 & ~n1617 ;
  assign n6801 = ~n6799 & n6800 ;
  assign n6802 = ~n6796 & n6801 ;
  assign n6803 = n6795 & ~n6802 ;
  assign n6790 = \i_tv80_core_BusAck_reg/P0001  & \i_tv80_core_mcycles_reg[2]/P0001  ;
  assign n6791 = \i_tv80_core_IR_reg[2]/P0001  & ~n681 ;
  assign n6792 = n990 & ~n6791 ;
  assign n6793 = ~n1005 & ~n6792 ;
  assign n6794 = n6704 & ~n6793 ;
  assign n6804 = ~n6790 & ~n6794 ;
  assign n6805 = ~n6803 & n6804 ;
  assign n6806 = reset_n_pad & ~n6805 ;
  assign n6809 = \i_tv80_core_IR_reg[4]/P0001  & n4723 ;
  assign n6810 = n1635 & ~n6809 ;
  assign n6811 = ~n4722 & n6810 ;
  assign n6812 = \i_tv80_core_XY_Ind_reg/P0001  & ~n6811 ;
  assign n6813 = ~\i_tv80_core_BusAck_reg/P0001  & n1113 ;
  assign n6814 = ~n6812 & n6813 ;
  assign n6807 = ~\i_tv80_core_BusAck_reg/P0001  & n862 ;
  assign n6808 = ~\i_tv80_core_XY_Ind_reg/P0001  & ~n6807 ;
  assign n6815 = reset_n_pad & ~n6808 ;
  assign n6816 = ~n6814 & n6815 ;
  assign n6817 = ~n6726 & ~n6729 ;
  assign n6818 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6817 ;
  assign n6820 = ~\i_tv80_core_R_reg[3]/P0001  & ~n6726 ;
  assign n6821 = \i_tv80_core_ACC_reg[3]/P0001  & n6726 ;
  assign n6822 = ~n6820 & ~n6821 ;
  assign n6823 = n6818 & n6822 ;
  assign n6819 = ~\i_tv80_core_R_reg[3]/P0001  & ~n6818 ;
  assign n6824 = reset_n_pad & ~n6819 ;
  assign n6825 = ~n6823 & n6824 ;
  assign n6826 = reset_n_pad & ~n860 ;
  assign n6827 = n6594 & n6826 ;
  assign n6830 = ~\i_tv80_core_R_reg[0]/P0001  & ~n5310 ;
  assign n6831 = ~n6726 & ~n6727 ;
  assign n6832 = ~n6830 & n6831 ;
  assign n6829 = \i_tv80_core_ACC_reg[0]/P0001  & n6726 ;
  assign n6833 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6829 ;
  assign n6834 = ~n6832 & n6833 ;
  assign n6828 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_R_reg[0]/P0001  ;
  assign n6835 = reset_n_pad & ~n6828 ;
  assign n6836 = ~n6834 & n6835 ;
  assign n6839 = ~\i_tv80_core_R_reg[2]/P0001  & ~n6728 ;
  assign n6840 = n6817 & ~n6839 ;
  assign n6838 = \i_tv80_core_ACC_reg[2]/P0001  & n6726 ;
  assign n6841 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6838 ;
  assign n6842 = ~n6840 & n6841 ;
  assign n6837 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_R_reg[2]/P0001  ;
  assign n6843 = reset_n_pad & ~n6837 ;
  assign n6844 = ~n6842 & n6843 ;
  assign n6847 = ~\i_tv80_core_R_reg[4]/P0001  & ~n6730 ;
  assign n6848 = n6732 & ~n6847 ;
  assign n6846 = \i_tv80_core_ACC_reg[4]/P0001  & n6726 ;
  assign n6849 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6846 ;
  assign n6850 = ~n6848 & n6849 ;
  assign n6845 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_R_reg[4]/P0001  ;
  assign n6851 = reset_n_pad & ~n6845 ;
  assign n6852 = ~n6850 & n6851 ;
  assign n6853 = n4722 & ~n6809 ;
  assign n6854 = ~\i_tv80_core_BusAck_reg/P0001  & n5310 ;
  assign n6855 = ~n6853 & n6854 ;
  assign n6856 = \i_tv80_core_XY_State_reg[1]/P0001  & ~n6855 ;
  assign n6857 = n4723 & n6854 ;
  assign n6858 = n675 & n6857 ;
  assign n6859 = ~n6856 & ~n6858 ;
  assign n6860 = reset_n_pad & ~n6859 ;
  assign n6861 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6831 ;
  assign n6863 = ~\i_tv80_core_R_reg[1]/P0001  & ~n6726 ;
  assign n6864 = \i_tv80_core_ACC_reg[1]/P0001  & n6726 ;
  assign n6865 = ~n6863 & ~n6864 ;
  assign n6866 = n6861 & n6865 ;
  assign n6862 = ~\i_tv80_core_R_reg[1]/P0001  & ~n6861 ;
  assign n6867 = reset_n_pad & ~n6862 ;
  assign n6868 = ~n6866 & n6867 ;
  assign n6869 = \i_tv80_core_XY_State_reg[0]/NET0131  & ~n6855 ;
  assign n6870 = n620 & n6857 ;
  assign n6871 = ~n6869 & ~n6870 ;
  assign n6872 = reset_n_pad & ~n6871 ;
  assign n6873 = \i_tv80_core_ISet_reg[0]/NET0131  & ~n6854 ;
  assign n6874 = n5310 & ~n6809 ;
  assign n6875 = ~n862 & ~n6874 ;
  assign n6876 = n1334 & n6795 ;
  assign n6877 = ~n6875 & n6876 ;
  assign n6878 = ~n6873 & ~n6877 ;
  assign n6879 = reset_n_pad & ~n6878 ;
  assign n6880 = ~\i_tv80_core_BusAck_reg/P0001  & n6726 ;
  assign n6882 = ~\i_tv80_core_R_reg[7]/P0001  & ~n6880 ;
  assign n6881 = ~\i_tv80_core_ACC_reg[7]/P0001  & n6880 ;
  assign n6883 = reset_n_pad & ~n6881 ;
  assign n6884 = ~n6882 & n6883 ;
  assign n6886 = n901 & n1575 ;
  assign n6887 = ~\i_tv80_core_IR_reg[0]/P0001  & n645 ;
  assign n6885 = \i_tv80_core_IR_reg[0]/P0001  & ~n675 ;
  assign n6888 = ~n676 & ~n6885 ;
  assign n6889 = ~n6887 & n6888 ;
  assign n6890 = n6886 & n6889 ;
  assign n6892 = ~\i_tv80_core_IR_reg[0]/P0001  & ~n678 ;
  assign n6893 = n6886 & n6892 ;
  assign n6894 = ~n6890 & ~n6893 ;
  assign n6895 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6894 ;
  assign n6896 = ~\i_tv80_core_IStatus_reg[0]/P0001  & ~n6895 ;
  assign n6891 = ~\i_tv80_core_BusAck_reg/P0001  & n6890 ;
  assign n6897 = reset_n_pad & ~n6891 ;
  assign n6898 = ~n6896 & n6897 ;
  assign n6900 = ~\i_tv80_core_IStatus_reg[1]/P0001  & ~n6895 ;
  assign n6899 = ~\i_tv80_core_BusAck_reg/P0001  & n6893 ;
  assign n6901 = reset_n_pad & ~n6899 ;
  assign n6902 = ~n6900 & n6901 ;
  assign n6903 = n862 & n4722 ;
  assign n6904 = ~n5310 & ~n6903 ;
  assign n6905 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6904 ;
  assign n6906 = \i_tv80_core_ISet_reg[1]/P0001  & ~n6905 ;
  assign n6907 = ~\i_tv80_core_BusAck_reg/P0001  & n4724 ;
  assign n6908 = n6874 & n6907 ;
  assign n6909 = ~n6906 & ~n6908 ;
  assign n6910 = reset_n_pad & ~n6909 ;
  assign n6911 = \di[0]_pad  & n1635 ;
  assign n6912 = ~\i_tv80_core_Halt_FF_reg/P0001  & ~\i_tv80_core_NMICycle_reg/P0001  ;
  assign n6913 = ~n1316 & n6912 ;
  assign n6914 = n6911 & n6913 ;
  assign n6915 = \i_tv80_core_IStatus_reg[0]/P0001  & ~\i_tv80_core_IStatus_reg[1]/P0001  ;
  assign n6916 = \i_tv80_core_IntCycle_reg/P0001  & n6915 ;
  assign n6917 = n1635 & n6916 ;
  assign n6918 = ~n6914 & ~n6917 ;
  assign n6919 = n1113 & ~n6918 ;
  assign n6920 = n1430 & n1462 ;
  assign n6921 = n6911 & n6920 ;
  assign n6922 = ~n6919 & ~n6921 ;
  assign n6923 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6922 ;
  assign n6924 = ~n860 & ~n6920 ;
  assign n6925 = ~\i_tv80_core_BusAck_reg/P0001  & n1635 ;
  assign n6926 = ~n6924 & n6925 ;
  assign n6927 = \i_tv80_core_IR_reg[0]/P0001  & ~n6926 ;
  assign n6928 = ~n6923 & ~n6927 ;
  assign n6929 = reset_n_pad & ~n6928 ;
  assign n6930 = \di[1]_pad  & n1635 ;
  assign n6931 = n6913 & n6930 ;
  assign n6932 = ~n6917 & ~n6931 ;
  assign n6933 = n1113 & ~n6932 ;
  assign n6934 = n6920 & n6930 ;
  assign n6935 = ~n6933 & ~n6934 ;
  assign n6936 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6935 ;
  assign n6937 = \i_tv80_core_IR_reg[1]/P0001  & ~n6926 ;
  assign n6938 = ~n6936 & ~n6937 ;
  assign n6939 = reset_n_pad & ~n6938 ;
  assign n6940 = \di[2]_pad  & n1635 ;
  assign n6941 = n6913 & n6940 ;
  assign n6942 = ~n6917 & ~n6941 ;
  assign n6943 = n1113 & ~n6942 ;
  assign n6944 = n6920 & n6940 ;
  assign n6945 = ~n6943 & ~n6944 ;
  assign n6946 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6945 ;
  assign n6947 = \i_tv80_core_IR_reg[2]/P0001  & ~n6926 ;
  assign n6948 = ~n6946 & ~n6947 ;
  assign n6949 = reset_n_pad & ~n6948 ;
  assign n6950 = \di[3]_pad  & n1635 ;
  assign n6951 = n6913 & n6950 ;
  assign n6952 = ~n6917 & ~n6951 ;
  assign n6953 = n1113 & ~n6952 ;
  assign n6954 = n6920 & n6950 ;
  assign n6955 = ~n6953 & ~n6954 ;
  assign n6956 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6955 ;
  assign n6957 = \i_tv80_core_IR_reg[3]/P0001  & ~n6926 ;
  assign n6958 = ~n6956 & ~n6957 ;
  assign n6959 = reset_n_pad & ~n6958 ;
  assign n6960 = \di[4]_pad  & n1635 ;
  assign n6961 = n6913 & n6960 ;
  assign n6962 = ~n6917 & ~n6961 ;
  assign n6963 = n1113 & ~n6962 ;
  assign n6964 = n6920 & n6960 ;
  assign n6965 = ~n6963 & ~n6964 ;
  assign n6966 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6965 ;
  assign n6967 = \i_tv80_core_IR_reg[4]/P0001  & ~n6926 ;
  assign n6968 = ~n6966 & ~n6967 ;
  assign n6969 = reset_n_pad & ~n6968 ;
  assign n6970 = \di[5]_pad  & n1635 ;
  assign n6971 = n6913 & n6970 ;
  assign n6972 = ~n6917 & ~n6971 ;
  assign n6973 = n1113 & ~n6972 ;
  assign n6974 = n6920 & n6970 ;
  assign n6975 = ~n6973 & ~n6974 ;
  assign n6976 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6975 ;
  assign n6977 = \i_tv80_core_IR_reg[5]/P0001  & ~n6926 ;
  assign n6978 = ~n6976 & ~n6977 ;
  assign n6979 = reset_n_pad & ~n6978 ;
  assign n6980 = \di[6]_pad  & n1635 ;
  assign n6981 = n6913 & n6980 ;
  assign n6982 = ~n6917 & ~n6981 ;
  assign n6983 = n1113 & ~n6982 ;
  assign n6984 = n6920 & n6980 ;
  assign n6985 = ~n6983 & ~n6984 ;
  assign n6986 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6985 ;
  assign n6987 = \i_tv80_core_IR_reg[6]/P0001  & ~n6926 ;
  assign n6988 = ~n6986 & ~n6987 ;
  assign n6989 = reset_n_pad & ~n6988 ;
  assign n6990 = \di[7]_pad  & n1635 ;
  assign n6991 = n6913 & n6990 ;
  assign n6992 = ~n6917 & ~n6991 ;
  assign n6993 = n1113 & ~n6992 ;
  assign n6994 = n6920 & n6990 ;
  assign n6995 = ~n6993 & ~n6994 ;
  assign n6996 = ~\i_tv80_core_BusAck_reg/P0001  & ~n6995 ;
  assign n6997 = \i_tv80_core_IR_reg[7]/P0001  & ~n6926 ;
  assign n6998 = ~n6996 & ~n6997 ;
  assign n6999 = reset_n_pad & ~n6998 ;
  assign n7001 = n382 & ~n6114 ;
  assign n7002 = \i_tv80_core_ISet_reg[1]/P0001  & n2712 ;
  assign n7003 = ~\i_tv80_core_BusAck_reg/P0001  & ~n7002 ;
  assign n7004 = ~n7001 & n7003 ;
  assign n7000 = \i_tv80_core_BusAck_reg/P0001  & ~\i_tv80_core_PreserveC_r_reg/P0001  ;
  assign n7005 = reset_n_pad & ~n7000 ;
  assign n7006 = ~n7004 & n7005 ;
  assign n7007 = n382 & n1384 ;
  assign n7008 = n4964 & n7007 ;
  assign n7010 = \i_tv80_core_Alternate_reg/P0001  & n7008 ;
  assign n7009 = ~\i_tv80_core_Alternate_reg/P0001  & ~n7008 ;
  assign n7011 = reset_n_pad & ~n7009 ;
  assign n7012 = ~n7010 & n7011 ;
  assign n7013 = ~\i_tv80_core_BusAck_reg/P0001  & n668 ;
  assign n7014 = n1111 & n7013 ;
  assign n7016 = ~\i_tv80_core_ACC_reg[0]/P0001  & n7014 ;
  assign n7015 = ~\i_tv80_core_I_reg[0]/P0001  & ~n7014 ;
  assign n7017 = reset_n_pad & ~n7015 ;
  assign n7018 = ~n7016 & n7017 ;
  assign n7020 = ~\i_tv80_core_ACC_reg[1]/P0001  & n7014 ;
  assign n7019 = ~\i_tv80_core_I_reg[1]/P0001  & ~n7014 ;
  assign n7021 = reset_n_pad & ~n7019 ;
  assign n7022 = ~n7020 & n7021 ;
  assign n7024 = ~\i_tv80_core_ACC_reg[2]/P0001  & n7014 ;
  assign n7023 = ~\i_tv80_core_I_reg[2]/P0001  & ~n7014 ;
  assign n7025 = reset_n_pad & ~n7023 ;
  assign n7026 = ~n7024 & n7025 ;
  assign n7028 = ~\i_tv80_core_ACC_reg[3]/P0001  & n7014 ;
  assign n7027 = ~\i_tv80_core_I_reg[3]/P0001  & ~n7014 ;
  assign n7029 = reset_n_pad & ~n7027 ;
  assign n7030 = ~n7028 & n7029 ;
  assign n7032 = ~\i_tv80_core_ACC_reg[4]/P0001  & n7014 ;
  assign n7031 = ~\i_tv80_core_I_reg[4]/P0001  & ~n7014 ;
  assign n7033 = reset_n_pad & ~n7031 ;
  assign n7034 = ~n7032 & n7033 ;
  assign n7036 = ~\i_tv80_core_ACC_reg[5]/P0001  & n7014 ;
  assign n7035 = ~\i_tv80_core_I_reg[5]/P0001  & ~n7014 ;
  assign n7037 = reset_n_pad & ~n7035 ;
  assign n7038 = ~n7036 & n7037 ;
  assign n7040 = ~\i_tv80_core_ACC_reg[6]/P0001  & n7014 ;
  assign n7039 = ~\i_tv80_core_I_reg[6]/P0001  & ~n7014 ;
  assign n7041 = reset_n_pad & ~n7039 ;
  assign n7042 = ~n7040 & n7041 ;
  assign n7044 = ~\i_tv80_core_ACC_reg[7]/P0001  & n7014 ;
  assign n7043 = ~\i_tv80_core_I_reg[7]/P0001  & ~n7014 ;
  assign n7045 = reset_n_pad & ~n7043 ;
  assign n7046 = ~n7044 & n7045 ;
  assign n7047 = ~\i_tv80_core_F_reg[6]/P0001  & \i_tv80_core_IR_reg[4]/P0001  ;
  assign n7048 = n1006 & ~n7047 ;
  assign n7049 = \i_tv80_core_F_reg[6]/P0001  & \i_tv80_core_IR_reg[0]/P0001  ;
  assign n7050 = \i_tv80_core_F_reg[2]/P0001  & \i_tv80_core_IR_reg[4]/P0001  ;
  assign n7051 = ~n7049 & n7050 ;
  assign n7052 = n1012 & ~n7051 ;
  assign n7053 = ~n7048 & ~n7052 ;
  assign n7054 = reset_n_pad & n1128 ;
  assign n7055 = ~n7053 & n7054 ;
  assign n7056 = n1117 & n4964 ;
  assign n7058 = \i_tv80_core_Ap_reg[2]/P0001  & ~n7056 ;
  assign n7057 = \i_tv80_core_ACC_reg[2]/P0001  & n7056 ;
  assign n7059 = reset_n_pad & ~n7057 ;
  assign n7060 = ~n7058 & n7059 ;
  assign n7062 = \i_tv80_core_Fp_reg[0]/P0001  & ~n7056 ;
  assign n7061 = \i_tv80_core_F_reg[0]/P0001  & n7056 ;
  assign n7063 = reset_n_pad & ~n7061 ;
  assign n7064 = ~n7062 & n7063 ;
  assign n7066 = \i_tv80_core_Fp_reg[1]/P0001  & ~n7056 ;
  assign n7065 = \i_tv80_core_F_reg[1]/P0001  & n7056 ;
  assign n7067 = reset_n_pad & ~n7065 ;
  assign n7068 = ~n7066 & n7067 ;
  assign n7070 = \i_tv80_core_Fp_reg[2]/P0001  & ~n7056 ;
  assign n7069 = \i_tv80_core_F_reg[2]/P0001  & n7056 ;
  assign n7071 = reset_n_pad & ~n7069 ;
  assign n7072 = ~n7070 & n7071 ;
  assign n7074 = \i_tv80_core_Fp_reg[3]/P0001  & ~n7056 ;
  assign n7073 = \i_tv80_core_F_reg[3]/P0001  & n7056 ;
  assign n7075 = reset_n_pad & ~n7073 ;
  assign n7076 = ~n7074 & n7075 ;
  assign n7078 = \i_tv80_core_Fp_reg[4]/P0001  & ~n7056 ;
  assign n7077 = \i_tv80_core_F_reg[4]/P0001  & n7056 ;
  assign n7079 = reset_n_pad & ~n7077 ;
  assign n7080 = ~n7078 & n7079 ;
  assign n7082 = \i_tv80_core_Fp_reg[5]/P0001  & ~n7056 ;
  assign n7081 = \i_tv80_core_F_reg[5]/P0001  & n7056 ;
  assign n7083 = reset_n_pad & ~n7081 ;
  assign n7084 = ~n7082 & n7083 ;
  assign n7086 = \i_tv80_core_Fp_reg[6]/P0001  & ~n7056 ;
  assign n7085 = \i_tv80_core_F_reg[6]/P0001  & n7056 ;
  assign n7087 = reset_n_pad & ~n7085 ;
  assign n7088 = ~n7086 & n7087 ;
  assign n7090 = \i_tv80_core_Fp_reg[7]/P0001  & ~n7056 ;
  assign n7089 = \i_tv80_core_F_reg[7]/P0001  & n7056 ;
  assign n7091 = reset_n_pad & ~n7089 ;
  assign n7092 = ~n7090 & n7091 ;
  assign n7094 = \i_tv80_core_Ap_reg[0]/P0001  & ~n7056 ;
  assign n7093 = \i_tv80_core_ACC_reg[0]/P0001  & n7056 ;
  assign n7095 = reset_n_pad & ~n7093 ;
  assign n7096 = ~n7094 & n7095 ;
  assign n7098 = \i_tv80_core_Ap_reg[1]/P0001  & ~n7056 ;
  assign n7097 = \i_tv80_core_ACC_reg[1]/P0001  & n7056 ;
  assign n7099 = reset_n_pad & ~n7097 ;
  assign n7100 = ~n7098 & n7099 ;
  assign n7102 = \i_tv80_core_Ap_reg[3]/P0001  & ~n7056 ;
  assign n7101 = \i_tv80_core_ACC_reg[3]/P0001  & n7056 ;
  assign n7103 = reset_n_pad & ~n7101 ;
  assign n7104 = ~n7102 & n7103 ;
  assign n7106 = \i_tv80_core_Ap_reg[4]/P0001  & ~n7056 ;
  assign n7105 = \i_tv80_core_ACC_reg[4]/P0001  & n7056 ;
  assign n7107 = reset_n_pad & ~n7105 ;
  assign n7108 = ~n7106 & n7107 ;
  assign n7110 = \i_tv80_core_Ap_reg[5]/P0001  & ~n7056 ;
  assign n7109 = \i_tv80_core_ACC_reg[5]/P0001  & n7056 ;
  assign n7111 = reset_n_pad & ~n7109 ;
  assign n7112 = ~n7110 & n7111 ;
  assign n7114 = \i_tv80_core_Ap_reg[6]/P0001  & ~n7056 ;
  assign n7113 = \i_tv80_core_ACC_reg[6]/P0001  & n7056 ;
  assign n7115 = reset_n_pad & ~n7113 ;
  assign n7116 = ~n7114 & n7115 ;
  assign n7118 = \i_tv80_core_Ap_reg[7]/P0001  & ~n7056 ;
  assign n7117 = \i_tv80_core_ACC_reg[7]/P0001  & n7056 ;
  assign n7119 = reset_n_pad & ~n7117 ;
  assign n7120 = ~n7118 & n7119 ;
  assign n7121 = \i_tv80_core_XY_State_reg[1]/P0001  & ~n6560 ;
  assign n7122 = \i_tv80_core_Alternate_reg/P0001  & n6560 ;
  assign n7123 = ~n7121 & ~n7122 ;
  assign n7124 = ~n2617 & ~n5310 ;
  assign n7125 = reset_n_pad & ~n7124 ;
  assign n7126 = \i_tv80_core_Arith16_r_reg/P0001  & n6028 ;
  assign n7127 = n382 & n6105 ;
  assign n7128 = n5773 & n7127 ;
  assign n7129 = ~n7126 & ~n7128 ;
  assign n7130 = \di_reg_reg[1]/P0001  & ~n1635 ;
  assign n7131 = ~n6930 & ~n7130 ;
  assign n7132 = reset_n_pad & ~n7131 ;
  assign n7133 = \di_reg_reg[3]/P0001  & ~n1635 ;
  assign n7134 = ~n6950 & ~n7133 ;
  assign n7135 = reset_n_pad & ~n7134 ;
  assign n7136 = \di_reg_reg[5]/P0001  & ~n1635 ;
  assign n7137 = ~n6970 & ~n7136 ;
  assign n7138 = reset_n_pad & ~n7137 ;
  assign n7139 = \di_reg_reg[4]/P0001  & ~n1635 ;
  assign n7140 = ~n6960 & ~n7139 ;
  assign n7141 = reset_n_pad & ~n7140 ;
  assign n7142 = \di_reg_reg[6]/P0001  & ~n1635 ;
  assign n7143 = ~n6980 & ~n7142 ;
  assign n7144 = reset_n_pad & ~n7143 ;
  assign n7145 = \di_reg_reg[7]/P0001  & ~n1635 ;
  assign n7146 = ~n6990 & ~n7145 ;
  assign n7147 = reset_n_pad & ~n7146 ;
  assign n7148 = \di_reg_reg[2]/P0001  & ~n1635 ;
  assign n7149 = ~n6940 & ~n7148 ;
  assign n7150 = reset_n_pad & ~n7149 ;
  assign n7151 = \di_reg_reg[0]/P0001  & ~n1635 ;
  assign n7152 = ~n6911 & ~n7151 ;
  assign n7153 = reset_n_pad & ~n7152 ;
  assign n7154 = \i_tv80_core_Oldnmi_n_reg/P0001  & ~nmi_n_pad ;
  assign n7155 = ~\i_tv80_core_NMI_s_reg/P0001  & ~n7154 ;
  assign n7156 = ~\i_tv80_core_NMICycle_reg/P0001  & reset_n_pad ;
  assign n7157 = ~n7155 & n7156 ;
  assign n7158 = ~busrq_n_pad & reset_n_pad ;
  assign n7159 = ~int_n_pad & reset_n_pad ;
  assign n7160 = nmi_n_pad & reset_n_pad ;
  assign n7161 = ~n3408 & n3410 ;
  assign n7162 = n2731 & ~n7161 ;
  assign n7163 = \i_tv80_core_i_reg_RegsH_reg[7][7]/P0002  & ~n2731 ;
  assign n7164 = ~n7162 & ~n7163 ;
  assign n7165 = n3456 & ~n3691 ;
  assign n7166 = \i_tv80_core_i_reg_RegsH_reg[0][4]/P0001  & ~n3456 ;
  assign n7167 = ~n7165 & ~n7166 ;
  assign n7168 = ~n3691 & n4081 ;
  assign n7169 = \i_tv80_core_i_reg_RegsH_reg[5][4]/P0001  & ~n4081 ;
  assign n7170 = ~n7168 & ~n7169 ;
  assign n7171 = ~n3691 & n4034 ;
  assign n7172 = \i_tv80_core_i_reg_RegsH_reg[2][4]/P0001  & ~n4034 ;
  assign n7173 = ~n7171 & ~n7172 ;
  assign n7174 = ~n3691 & n4088 ;
  assign n7175 = \i_tv80_core_i_reg_RegsH_reg[6][4]/P0001  & ~n4088 ;
  assign n7176 = ~n7174 & ~n7175 ;
  assign n7177 = ~n3503 & n4081 ;
  assign n7178 = \i_tv80_core_i_reg_RegsH_reg[5][6]/P0001  & ~n4081 ;
  assign n7179 = ~n7177 & ~n7178 ;
  assign n7180 = ~n3503 & n3636 ;
  assign n7181 = \i_tv80_core_i_reg_RegsH_reg[1][6]/P0001  & ~n3636 ;
  assign n7182 = ~n7180 & ~n7181 ;
  assign n7183 = ~n3503 & n4088 ;
  assign n7184 = \i_tv80_core_i_reg_RegsH_reg[6][6]/P0001  & ~n4088 ;
  assign n7185 = ~n7183 & ~n7184 ;
  assign n7186 = n3636 & ~n3892 ;
  assign n7187 = \i_tv80_core_i_reg_RegsH_reg[1][2]/P0001  & ~n3636 ;
  assign n7188 = ~n7186 & ~n7187 ;
  assign n7189 = \i_tv80_core_i_reg_RegsH_reg[0][0]/P0001  & ~n3456 ;
  assign n7190 = n3456 & n4124 ;
  assign n7191 = ~n7189 & ~n7190 ;
  assign n7192 = ~n3892 & n4088 ;
  assign n7193 = \i_tv80_core_i_reg_RegsH_reg[6][2]/P0001  & ~n4088 ;
  assign n7194 = ~n7192 & ~n7193 ;
  assign n7195 = ~n3892 & n4034 ;
  assign n7196 = \i_tv80_core_i_reg_RegsH_reg[2][2]/P0001  & ~n4034 ;
  assign n7197 = ~n7195 & ~n7196 ;
  assign n7198 = ~n3632 & n3636 ;
  assign n7199 = \i_tv80_core_i_reg_RegsH_reg[1][5]/P0001  & ~n3636 ;
  assign n7200 = ~n7198 & ~n7199 ;
  assign n7201 = ~n3892 & n4081 ;
  assign n7202 = \i_tv80_core_i_reg_RegsH_reg[5][2]/P0001  & ~n4081 ;
  assign n7203 = ~n7201 & ~n7202 ;
  assign n7204 = n3636 & ~n4062 ;
  assign n7205 = \i_tv80_core_i_reg_RegsH_reg[1][1]/P0001  & ~n3636 ;
  assign n7206 = ~n7204 & ~n7205 ;
  assign n7207 = ~n3632 & n4034 ;
  assign n7208 = \i_tv80_core_i_reg_RegsH_reg[2][5]/P0001  & ~n4034 ;
  assign n7209 = ~n7207 & ~n7208 ;
  assign n7210 = n3456 & ~n4062 ;
  assign n7211 = \i_tv80_core_i_reg_RegsH_reg[0][1]/P0001  & ~n3456 ;
  assign n7212 = ~n7210 & ~n7211 ;
  assign n7213 = ~n2618 & ~n2646 ;
  assign n7214 = n2659 & n7213 ;
  assign n7215 = n2674 & n7214 ;
  assign n7216 = n5512 & n7215 ;
  assign n7217 = n4668 & n7216 ;
  assign n7218 = ~n4511 & n7217 ;
  assign n7219 = ~n4247 & n7218 ;
  assign n7220 = ~n4338 & n7219 ;
  assign n7221 = ~n2889 & n7220 ;
  assign n7222 = ~n3523 & ~n4039 ;
  assign n7223 = n7221 & n7222 ;
  assign n7226 = ~n3648 & n7223 ;
  assign n7227 = ~n3869 & n7226 ;
  assign n7224 = ~n3613 & ~n4021 ;
  assign n7225 = ~n4119 & n7224 ;
  assign n7228 = ~n3407 & n7225 ;
  assign n7229 = n7227 & n7228 ;
  assign n7230 = ~n3480 & n7229 ;
  assign n7231 = \i_tv80_core_Save_ALU_r_reg/P0001  & n384 ;
  assign n7233 = ~n1258 & n7231 ;
  assign n7232 = \i_tv80_core_IncDecZ_reg/P0002  & ~n7231 ;
  assign n7234 = ~n7215 & ~n7232 ;
  assign n7235 = ~n7233 & n7234 ;
  assign n7236 = ~n7230 & ~n7235 ;
  assign n7237 = ~n4062 & n4088 ;
  assign n7238 = \i_tv80_core_i_reg_RegsH_reg[6][1]/P0001  & ~n4088 ;
  assign n7239 = ~n7237 & ~n7238 ;
  assign n7240 = \i_tv80_core_i_reg_RegsH_reg[5][5]/P0001  & ~n4081 ;
  assign n7241 = ~n3615 & n4081 ;
  assign n7242 = ~n7240 & ~n7241 ;
  assign n7243 = ~n3632 & n4088 ;
  assign n7244 = \i_tv80_core_i_reg_RegsH_reg[6][5]/P0001  & ~n4088 ;
  assign n7245 = ~n7243 & ~n7244 ;
  assign n7246 = ~n3503 & n4034 ;
  assign n7247 = \i_tv80_core_i_reg_RegsH_reg[2][6]/P0001  & ~n4034 ;
  assign n7248 = ~n7246 & ~n7247 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g28227/_0_  = ~n1199 ;
  assign \g28233/_0_  = ~n1275 ;
  assign \g28274/_0_  = n1644 ;
  assign \g28275/_0_  = n1701 ;
  assign \g28276/_0_  = n1762 ;
  assign \g28277/_0_  = n1820 ;
  assign \g28278/_0_  = ~n1868 ;
  assign \g28279/_0_  = n1928 ;
  assign \g28280/_0_  = n1999 ;
  assign \g28281/_0_  = n2062 ;
  assign \g28282/_0_  = n2125 ;
  assign \g28283/_0_  = n2188 ;
  assign \g28284/_0_  = n2251 ;
  assign \g28285/_0_  = n2314 ;
  assign \g28286/_0_  = n2373 ;
  assign \g28287/_0_  = n2432 ;
  assign \g28288/_0_  = n2492 ;
  assign \g28289/_0_  = n2554 ;
  assign \g28290/_0_  = n2616 ;
  assign \g28294/_0_  = ~n2936 ;
  assign \g28295/_0_  = ~n2940 ;
  assign \g28296/_0_  = ~n2944 ;
  assign \g28297/_0_  = ~n2948 ;
  assign \g28298/_0_  = ~n2952 ;
  assign \g28299/_0_  = ~n2956 ;
  assign \g28300/_0_  = ~n2960 ;
  assign \g28301/_0_  = ~n2964 ;
  assign \g28349/_0_  = n2988 ;
  assign \g28350/_0_  = ~n3086 ;
  assign \g28351/_0_  = ~n3141 ;
  assign \g28352/_0_  = ~n3169 ;
  assign \g28353/_0_  = ~n3251 ;
  assign \g28354/_0_  = n3432 ;
  assign \g28355/_0_  = n3435 ;
  assign \g28356/_0_  = n3438 ;
  assign \g28357/_0_  = n3441 ;
  assign \g28358/_0_  = n3444 ;
  assign \g28359/_0_  = n3447 ;
  assign \g28360/_0_  = n3450 ;
  assign \g28414/_0_  = ~n3506 ;
  assign \g28417/_0_  = ~n3510 ;
  assign \g28418/_0_  = ~n3514 ;
  assign \g28421/_0_  = ~n3518 ;
  assign \g28422/_0_  = ~n3547 ;
  assign \g28423/_0_  = ~n3550 ;
  assign \g28424/_0_  = ~n3553 ;
  assign \g28425/_0_  = ~n3556 ;
  assign \g28426/_0_  = ~n3559 ;
  assign \g28427/_0_  = ~n3562 ;
  assign \g28428/_0_  = ~n3565 ;
  assign \g28429/_0_  = ~n3568 ;
  assign \g28464/_0_  = ~n3635 ;
  assign \g28466/_0_  = ~n3694 ;
  assign \g28470/_0_  = ~n3697 ;
  assign \g28471/_0_  = ~n3700 ;
  assign \g28472/_0_  = ~n3703 ;
  assign \g28473/_0_  = ~n3706 ;
  assign \g28478/_0_  = ~n3709 ;
  assign \g28479/_0_  = ~n3712 ;
  assign \g28500/_0_  = n3728 ;
  assign \g28501/_0_  = ~n3750 ;
  assign \g28502/_0_  = ~n3789 ;
  assign \g28503/_0_  = ~n3808 ;
  assign \g28507/_0_  = ~n3827 ;
  assign \g28509/_0_  = ~n3865 ;
  assign \g28536/_0_  = ~n3895 ;
  assign \g28539/_0_  = ~n3898 ;
  assign \g28540/_0_  = ~n3901 ;
  assign \g28543/_0_  = ~n3904 ;
  assign \g28555/_0_  = ~n3923 ;
  assign \g28561/_0_  = ~n3942 ;
  assign \g28562/_0_  = ~n3961 ;
  assign \g28563/_0_  = ~n4000 ;
  assign \g28604/_0_  = n4030 ;
  assign \g28606/_0_  = n4033 ;
  assign \g28607/_0_  = ~n4065 ;
  assign \g28608/_0_  = n4068 ;
  assign \g28609/_0_  = ~n4071 ;
  assign \g28610/_0_  = n4074 ;
  assign \g28611/_0_  = ~n4077 ;
  assign \g28612/_0_  = n4080 ;
  assign \g28613/_0_  = ~n4084 ;
  assign \g28614/_0_  = n4087 ;
  assign \g28616/_0_  = n4091 ;
  assign \g28617/_0_  = ~n4094 ;
  assign \g28618/_0_  = n4097 ;
  assign \g28660/_0_  = ~n4128 ;
  assign \g28661/_0_  = ~n4131 ;
  assign \g28662/_0_  = ~n4134 ;
  assign \g28663/_0_  = ~n4137 ;
  assign \g28664/_0_  = ~n4140 ;
  assign \g28665/_0_  = ~n4143 ;
  assign \g28666/_0_  = ~n4146 ;
  assign \g28691/_0_  = ~n4172 ;
  assign \g28693/_0_  = ~n4209 ;
  assign \g28694/_0_  = ~n4242 ;
  assign \g28727/_0_  = ~n4271 ;
  assign \g28728/_0_  = ~n4274 ;
  assign \g28729/_0_  = ~n4277 ;
  assign \g28730/_0_  = ~n4280 ;
  assign \g28731/_0_  = ~n4283 ;
  assign \g28732/_0_  = ~n4286 ;
  assign \g28733/_0_  = ~n4289 ;
  assign \g28734/_0_  = ~n4292 ;
  assign \g28750/_0_  = n4310 ;
  assign \g28759/_0_  = ~n4333 ;
  assign \g28787/_0_  = ~n4362 ;
  assign \g28788/_0_  = ~n4365 ;
  assign \g28789/_0_  = ~n4368 ;
  assign \g28790/_0_  = ~n4371 ;
  assign \g28791/_0_  = ~n4374 ;
  assign \g28792/_0_  = ~n4377 ;
  assign \g28793/_0_  = ~n4380 ;
  assign \g28794/_0_  = ~n4383 ;
  assign \g28810/_0_  = n4406 ;
  assign \g28811/_0_  = n4417 ;
  assign \g28812/_0_  = n4424 ;
  assign \g28813/_0_  = n4440 ;
  assign \g28814/_0_  = ~n4460 ;
  assign \g28835/_0_  = ~n4482 ;
  assign \g28836/_0_  = ~n4506 ;
  assign \g28856/_0_  = ~n4535 ;
  assign \g28857/_0_  = ~n4538 ;
  assign \g28858/_0_  = ~n4541 ;
  assign \g28859/_0_  = ~n4544 ;
  assign \g28860/_0_  = ~n4547 ;
  assign \g28861/_0_  = ~n4550 ;
  assign \g28862/_0_  = ~n4553 ;
  assign \g28863/_0_  = ~n4556 ;
  assign \g28894/_0_  = n4572 ;
  assign \g28898/_0_  = ~n4592 ;
  assign \g28914/_0_  = ~n4608 ;
  assign \g28917/_0_  = ~n4638 ;
  assign \g28922/_0_  = ~n4651 ;
  assign \g28923/_0_  = n4663 ;
  assign \g28953/_0_  = ~n4692 ;
  assign \g28954/_0_  = ~n4695 ;
  assign \g28955/_0_  = ~n4698 ;
  assign \g28956/_0_  = ~n4701 ;
  assign \g28957/_0_  = ~n4704 ;
  assign \g28958/_0_  = ~n4707 ;
  assign \g28959/_0_  = ~n4710 ;
  assign \g28960/_0_  = ~n4713 ;
  assign \g28970/_0_  = n4730 ;
  assign \g28971/_0_  = n4736 ;
  assign \g28972/_0_  = n4811 ;
  assign \g28973/_0_  = n4891 ;
  assign \g28974/_0_  = n4928 ;
  assign \g28975/_0_  = n4962 ;
  assign \g28976/_0_  = n4996 ;
  assign \g28977/_0_  = n5031 ;
  assign \g28978/_0_  = n5071 ;
  assign \g28979/_0_  = n5096 ;
  assign \g28980/_0_  = n5121 ;
  assign \g28981/_0_  = n5148 ;
  assign \g28982/_0_  = n5175 ;
  assign \g28983/_0_  = n5200 ;
  assign \g28984/_0_  = n5225 ;
  assign \g28985/_0_  = n5252 ;
  assign \g28986/_0_  = n5280 ;
  assign \g28987/_0_  = n5308 ;
  assign \g28988/_0_  = ~n5314 ;
  assign \g28993/_0_  = n5324 ;
  assign \g28994/_0_  = ~n5344 ;
  assign \g29029/_0_  = ~n5367 ;
  assign \g29081/_0_  = n5371 ;
  assign \g29082/_0_  = n5381 ;
  assign \g29083/_0_  = n5397 ;
  assign \g29084/_0_  = n5413 ;
  assign \g29085/_0_  = n5429 ;
  assign \g29086/_0_  = n5445 ;
  assign \g29093/_0_  = ~n5465 ;
  assign \g29188/_0_  = n5470 ;
  assign \g29189/_0_  = n5474 ;
  assign \g29190/_0_  = n5478 ;
  assign \g29191/_0_  = n5488 ;
  assign \g29192/_0_  = n5498 ;
  assign \g29193/_0_  = n5508 ;
  assign \g29221/_0_  = ~n5537 ;
  assign \g29222/_0_  = ~n5540 ;
  assign \g29223/_0_  = ~n5543 ;
  assign \g29224/_0_  = ~n5546 ;
  assign \g29225/_0_  = ~n5549 ;
  assign \g29227/_0_  = ~n5552 ;
  assign \g29228/_0_  = ~n5555 ;
  assign \g29229/_0_  = ~n5558 ;
  assign \g29366/_0_  = ~n5578 ;
  assign \g29385/_0_  = ~n5597 ;
  assign \g29387/_0_  = ~n5617 ;
  assign \g29388/_0_  = ~n5637 ;
  assign \g29405/_0_  = ~\i_tv80_core_BusAck_reg/P0001  ;
  assign \g29450/_0_  = n5647 ;
  assign \g29451/_0_  = n5663 ;
  assign \g29472/_0_  = n2710 ;
  assign \g29552/_0_  = n5683 ;
  assign \g29553/_0_  = n5693 ;
  assign \g29559/_0_  = ~n5820 ;
  assign \g29561/_0_  = ~n5834 ;
  assign \g29562/_0_  = ~n5848 ;
  assign \g29563/_0_  = ~n5862 ;
  assign \g29564/_0_  = ~n5876 ;
  assign \g29565/_0_  = ~n5890 ;
  assign \g29566/_0_  = ~n5904 ;
  assign \g29577/_0_  = ~n5918 ;
  assign \g29623/_0_  = ~n5943 ;
  assign \g29624/_0_  = ~n5946 ;
  assign \g29625/_0_  = ~n5949 ;
  assign \g29626/_0_  = ~n5952 ;
  assign \g29627/_0_  = ~n5955 ;
  assign \g29628/_0_  = ~n5958 ;
  assign \g29629/_0_  = ~n5961 ;
  assign \g29630/_0_  = ~n5964 ;
  assign \g29657/_0_  = n5977 ;
  assign \g29658/_0_  = n5987 ;
  assign \g29679/_0_  = n5992 ;
  assign \g29689/_3_  = ~n6001 ;
  assign \g29728/_0_  = n6014 ;
  assign \g29828/_0_  = n6027 ;
  assign \g29909/_3_  = ~n6063 ;
  assign \g29966/_0_  = n6073 ;
  assign \g30036/_3_  = ~n6078 ;
  assign \g30038/_3_  = n6085 ;
  assign \g30040/_3_  = n6090 ;
  assign \g30080/_0_  = n6100 ;
  assign \g30081/_0_  = n6102 ;
  assign \g30107/_0_  = n6103 ;
  assign \g30176/_0_  = ~n6109 ;
  assign \g30189/_3_  = ~n6122 ;
  assign \g30192/_3_  = ~n6132 ;
  assign \g30194/_3_  = ~n6210 ;
  assign \g30354/_0_  = ~n6247 ;
  assign \g30377/_0_  = ~n6280 ;
  assign \g30454/_2_  = n6283 ;
  assign \g30479/_2_  = n6288 ;
  assign \g30490/_0_  = ~n3299 ;
  assign \g30492/_1_  = ~n2754 ;
  assign \g30495/_0_  = ~n2770 ;
  assign \g30497/_1_  = ~n3266 ;
  assign \g30501/_1_  = ~n3357 ;
  assign \g30503/_1_  = ~n2823 ;
  assign \g30509/_1_  = ~n3325 ;
  assign \g30513/_0_  = ~n3401 ;
  assign \g30514/_0_  = ~n2840 ;
  assign \g30517/_0_  = ~n3341 ;
  assign \g30523/_0_  = ~n2788 ;
  assign \g30678/_0_  = ~n6430 ;
  assign \g30982/_0_  = ~n6449 ;
  assign \g30983/_0_  = ~n6467 ;
  assign \g30984/_0_  = ~n6485 ;
  assign \g30985/_0_  = ~n6503 ;
  assign \g30986/_0_  = ~n6521 ;
  assign \g30987/_0_  = ~n6539 ;
  assign \g30988/_0_  = ~n6557 ;
  assign \g30998/_0_  = ~n6564 ;
  assign \g31212/_0_  = ~n6618 ;
  assign \g31235/_0_  = ~n6626 ;
  assign \g31236/_0_  = ~n6631 ;
  assign \g31296/_3_  = ~n6635 ;
  assign \g31303/_0_  = n6690 ;
  assign \g31306/_0_  = n6700 ;
  assign \g31312/_0_  = ~n6702 ;
  assign \g31356/_0_  = n6709 ;
  assign \g31397/_0_  = ~n6714 ;
  assign \g31430/_0_  = ~n6718 ;
  assign \g31440/_3_  = ~n6721 ;
  assign \g31455/_3_  = ~n6725 ;
  assign \g31459/_0_  = n6742 ;
  assign \g31511/_0_  = n6781 ;
  assign \g31512/_0_  = n6789 ;
  assign \g31561/_0_  = n6806 ;
  assign \g31603/_0_  = n6816 ;
  assign \g31604/_0_  = n6825 ;
  assign \g31666/_0_  = ~n6827 ;
  assign \g31794/_0_  = n6836 ;
  assign \g31795/_0_  = n6844 ;
  assign \g31796/_0_  = n6852 ;
  assign \g31854/_0_  = n6860 ;
  assign \g31855/_0_  = n6868 ;
  assign \g31856/_0_  = n6872 ;
  assign \g31871/_0_  = n6879 ;
  assign \g31920/_0_  = n6884 ;
  assign \g31934/_0_  = n6898 ;
  assign \g31935/_0_  = n6902 ;
  assign \g31943/_0_  = n6910 ;
  assign \g32128/_0_  = n6929 ;
  assign \g32129/_0_  = n6939 ;
  assign \g32130/_0_  = n6949 ;
  assign \g32131/_0_  = n6959 ;
  assign \g32132/_0_  = n6969 ;
  assign \g32133/_0_  = n6979 ;
  assign \g32134/_0_  = n6989 ;
  assign \g32135/_0_  = n6999 ;
  assign \g32136/_0_  = n7006 ;
  assign \g32137/_0_  = n7012 ;
  assign \g32140/_0_  = n7018 ;
  assign \g32141/_0_  = n7022 ;
  assign \g32142/_0_  = n7026 ;
  assign \g32143/_0_  = n7030 ;
  assign \g32144/_0_  = n7034 ;
  assign \g32145/_0_  = n7038 ;
  assign \g32146/_0_  = n7042 ;
  assign \g32147/_0_  = n7046 ;
  assign \g32475/_0_  = n7055 ;
  assign \g32639/_0_  = ~n7060 ;
  assign \g32640/_0_  = ~n7064 ;
  assign \g32641/_0_  = ~n7068 ;
  assign \g32642/_0_  = ~n7072 ;
  assign \g32643/_0_  = ~n7076 ;
  assign \g32644/_0_  = ~n7080 ;
  assign \g32645/_0_  = ~n7084 ;
  assign \g32646/_0_  = ~n7088 ;
  assign \g32647/_0_  = ~n7092 ;
  assign \g32648/_0_  = ~n7096 ;
  assign \g32649/_0_  = ~n7100 ;
  assign \g32650/_0_  = ~n7104 ;
  assign \g32651/_0_  = ~n7108 ;
  assign \g32652/_0_  = ~n7112 ;
  assign \g32653/_0_  = ~n7116 ;
  assign \g32654/_0_  = ~n7120 ;
  assign \g32798/_3_  = ~n7123 ;
  assign \g33177/_0_  = ~n7125 ;
  assign \g33187/_0_  = ~n7129 ;
  assign \g33306/_0_  = n7132 ;
  assign \g33307/_0_  = n7135 ;
  assign \g33308/_0_  = n7138 ;
  assign \g33309/_0_  = n7141 ;
  assign \g33310/_0_  = n7144 ;
  assign \g33311/_0_  = n7147 ;
  assign \g33312/_0_  = n7150 ;
  assign \g33313/_0_  = n7153 ;
  assign \g34088/_0_  = n7157 ;
  assign \g35570/_0_  = n7158 ;
  assign \g35594/_0_  = n7159 ;
  assign \g35838/_0_  = n7160 ;
  assign \g37467/_0_  = ~n7164 ;
  assign \g37492/_0_  = ~n7167 ;
  assign \g37503/_0_  = ~n7170 ;
  assign \g37513/_0_  = ~n7173 ;
  assign \g37524/_0_  = ~n7176 ;
  assign \g37727/_0_  = ~n7179 ;
  assign \g37748/_0_  = ~n7182 ;
  assign \g37758/_0_  = ~n7185 ;
  assign \g37767/_0_  = ~n7188 ;
  assign \g37777/_0_  = ~n7191 ;
  assign \g37790/_0_  = ~n7194 ;
  assign \g37809/_0_  = ~n7197 ;
  assign \g37840/_0_  = ~n7200 ;
  assign \g37852/_0_  = ~n7203 ;
  assign \g38312_dup/_0_  = ~n3282 ;
  assign \g38324/_0_  = ~n2856 ;
  assign \g38354/_0_  = ~n2883 ;
  assign \g38781/_1_  = ~n2807 ;
  assign \g38840/_0_  = ~n7206 ;
  assign \g38851/_0_  = ~n7209 ;
  assign \g38866/_0_  = ~n7212 ;
  assign \g38892/_1_  = n7236 ;
  assign \g38932/_0_  = ~n7239 ;
  assign \g38943/_0_  = ~n7242 ;
  assign \g39103/_0_  = ~n7245 ;
  assign \g39113/_2__syn_2  = n3455 ;
  assign \g39127/_0_  = ~n3374 ;
  assign \g44/_0_  = ~n7248 ;
  assign halt_n_pad = ~\i_tv80_core_Halt_FF_reg/P0001  ;
endmodule
